module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 ,
    po6 , po7 , po8 , po9 , po10 ,
    po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 ,
    po21 , po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 , po30 ,
    po31 , po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 ,
    po46 , po47 , po48 , po49 , po50 ,
    po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 ,
    po61 , po62 , po63   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 ;
  wire n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535,
    n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201,
    n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291,
    n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321,
    n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351,
    n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381,
    n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411,
    n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441,
    n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471,
    n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501,
    n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531,
    n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681,
    n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711,
    n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741,
    n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771,
    n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801,
    n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831,
    n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861,
    n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921,
    n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951,
    n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101,
    n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131,
    n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161,
    n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173,
    n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191,
    n2192, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203,
    n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221,
    n2222, n2223, n2224, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311,
    n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341,
    n2342, n2343, n2344, n2345, n2346, n2347,
    n2348, n2349, n2350, n2351, n2352, n2353,
    n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371,
    n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461,
    n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581,
    n2582, n2583, n2584, n2585, n2586, n2587,
    n2588, n2589, n2590, n2591, n2592, n2593,
    n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617,
    n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641,
    n2642, n2643, n2644, n2645, n2646, n2647,
    n2648, n2649, n2650, n2651, n2652, n2653,
    n2654, n2655, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671,
    n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2680, n2681, n2682, n2683,
    n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2697, n2698, n2699, n2700, n2701,
    n2702, n2703, n2704, n2705, n2706, n2707,
    n2708, n2709, n2710, n2711, n2712, n2713,
    n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731,
    n2732, n2733, n2734, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743,
    n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761,
    n2762, n2763, n2764, n2765, n2766, n2767,
    n2768, n2769, n2770, n2771, n2772, n2773,
    n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791,
    n2792, n2793, n2794, n2795, n2796, n2797,
    n2798, n2799, n2800, n2801, n2802, n2803,
    n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821,
    n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851,
    n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2880, n2881,
    n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911,
    n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953,
    n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001,
    n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061,
    n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085,
    n3086, n3087, n3088, n3089, n3090, n3091,
    n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151,
    n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175,
    n3176, n3177, n3178, n3179, n3180, n3181,
    n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211,
    n3212, n3213, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241,
    n3242, n3243, n3244, n3245, n3246, n3247,
    n3248, n3249, n3250, n3251, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271,
    n3272, n3273, n3274, n3275, n3276, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541,
    n3542, n3543, n3544, n3545, n3546, n3547,
    n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565,
    n3566, n3567, n3568, n3569, n3570, n3571,
    n3572, n3573, n3574, n3575, n3576, n3577,
    n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601,
    n3602, n3603, n3604, n3605, n3606, n3607,
    n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631,
    n3632, n3633, n3634, n3635, n3636, n3637,
    n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661,
    n3662, n3663, n3664, n3665, n3666, n3667,
    n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691,
    n3692, n3693, n3694, n3695, n3696, n3697,
    n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721,
    n3722, n3723, n3724, n3725, n3726, n3727,
    n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751,
    n3752, n3753, n3754, n3755, n3756, n3757,
    n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775,
    n3776, n3777, n3778, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787,
    n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805,
    n3806, n3807, n3808, n3809, n3810, n3811,
    n3812, n3813, n3814, n3815, n3816, n3817,
    n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835,
    n3836, n3837, n3838, n3839, n3840, n3841,
    n3842, n3843, n3844, n3845, n3846, n3847,
    n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877,
    n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901,
    n3902, n3903, n3904, n3905, n3906, n3907,
    n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931,
    n3932, n3933, n3934, n3935, n3936, n3937,
    n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961,
    n3962, n3963, n3964, n3965, n3966, n3967,
    n3968, n3969, n3970, n3971, n3972, n3973,
    n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3991,
    n3992, n3993, n3994, n3995, n3996, n3997,
    n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057,
    n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117,
    n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141,
    n4142, n4143, n4144, n4145, n4146, n4147,
    n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171,
    n4172, n4173, n4174, n4175, n4176, n4177,
    n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195,
    n4196, n4197, n4198, n4199, n4200, n4201,
    n4202, n4203, n4204, n4205, n4206, n4207,
    n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219,
    n4220, n4221, n4222, n4223, n4224, n4225,
    n4226, n4227, n4228, n4229, n4230, n4231,
    n4232, n4233, n4234, n4235, n4236, n4237,
    n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249,
    n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4259, n4260, n4261,
    n4262, n4263, n4264, n4265, n4266, n4267,
    n4268, n4269, n4270, n4271, n4272, n4273,
    n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291,
    n4292, n4293, n4294, n4295, n4296, n4297,
    n4298, n4299, n4300, n4301, n4302, n4303,
    n4304, n4305, n4306, n4307, n4308, n4309,
    n4310, n4311, n4312, n4313, n4314, n4315,
    n4316, n4317, n4318, n4319, n4320, n4321,
    n4322, n4323, n4324, n4325, n4326, n4327,
    n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339,
    n4340, n4341, n4342, n4343, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351,
    n4352, n4353, n4354, n4355, n4356, n4357,
    n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369,
    n4370, n4371, n4372, n4373, n4374, n4375,
    n4376, n4377, n4378, n4379, n4380, n4381,
    n4382, n4383, n4384, n4385, n4386, n4387,
    n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399,
    n4400, n4401, n4402, n4403, n4404, n4405,
    n4406, n4407, n4408, n4409, n4410, n4411,
    n4412, n4413, n4414, n4415, n4416, n4417,
    n4418, n4419, n4420, n4421, n4422, n4423,
    n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435,
    n4436, n4437, n4438, n4439, n4440, n4441,
    n4442, n4443, n4444, n4445, n4446, n4447,
    n4448, n4449, n4450, n4451, n4452, n4453,
    n4454, n4455, n4456, n4457, n4458, n4459,
    n4460, n4461, n4462, n4463, n4464, n4465,
    n4466, n4467, n4468, n4469, n4470, n4471,
    n4472, n4473, n4474, n4475, n4476, n4477,
    n4478, n4479, n4480, n4481, n4482, n4483,
    n4484, n4485, n4486, n4487, n4488, n4489,
    n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501,
    n4502, n4503, n4504, n4505, n4506, n4507,
    n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531,
    n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843,
    n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861,
    n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873,
    n4874, n4875, n4876, n4877, n4878, n4879,
    n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891,
    n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137,
    n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161,
    n5162, n5163, n5164, n5165, n5166, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191,
    n5192, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209,
    n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221,
    n5222, n5223, n5224, n5225, n5226, n5227,
    n5228, n5229, n5230, n5231, n5232, n5233,
    n5234, n5235, n5236, n5237, n5238, n5239,
    n5240, n5241, n5242, n5243, n5244, n5245,
    n5246, n5247, n5248, n5249, n5250, n5251,
    n5252, n5253, n5254, n5255, n5256, n5257,
    n5258, n5259, n5260, n5261, n5262, n5263,
    n5264, n5265, n5266, n5267, n5268, n5269,
    n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281,
    n5282, n5283, n5284, n5285, n5286, n5287,
    n5288, n5289, n5290, n5291, n5292, n5293,
    n5294, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5308, n5309, n5310, n5311,
    n5312, n5313, n5314, n5315, n5316, n5317,
    n5318, n5319, n5320, n5321, n5322, n5323,
    n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335,
    n5336, n5337, n5338, n5339, n5340, n5341,
    n5342, n5343, n5344, n5345, n5346, n5347,
    n5348, n5349, n5350, n5351, n5352, n5353,
    n5354, n5355, n5356, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371,
    n5372, n5373, n5374, n5375, n5376, n5377,
    n5378, n5379, n5380, n5381, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389,
    n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401,
    n5402, n5403, n5404, n5405, n5406, n5407,
    n5408, n5409, n5410, n5411, n5412, n5413,
    n5414, n5415, n5416, n5417, n5418, n5419,
    n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431,
    n5432, n5433, n5434, n5435, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443,
    n5444, n5445, n5446, n5447, n5448, n5449,
    n5450, n5451, n5452, n5453, n5454, n5455,
    n5456, n5457, n5458, n5459, n5460, n5461,
    n5462, n5463, n5464, n5465, n5466, n5467,
    n5468, n5469, n5470, n5471, n5472, n5473,
    n5474, n5475, n5476, n5477, n5478, n5479,
    n5480, n5481, n5482, n5483, n5484, n5485,
    n5486, n5487, n5488, n5489, n5490, n5491,
    n5492, n5493, n5494, n5495, n5496, n5497,
    n5498, n5499, n5500, n5501, n5502, n5503,
    n5504, n5505, n5506, n5507, n5508, n5509,
    n5510, n5511, n5512, n5513, n5514, n5515,
    n5516, n5517, n5518, n5519, n5520, n5521,
    n5522, n5523, n5524, n5525, n5526, n5527,
    n5528, n5529, n5530, n5531, n5532, n5533,
    n5534, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551,
    n5552, n5553, n5554, n5555, n5556, n5557,
    n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581,
    n5582, n5583, n5584, n5585, n5586, n5587,
    n5588, n5589, n5590, n5591, n5592, n5593,
    n5594, n5595, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611,
    n5612, n5613, n5614, n5615, n5616, n5617,
    n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5625, n5626, n5627, n5628, n5629,
    n5630, n5631, n5632, n5633, n5634, n5635,
    n5636, n5637, n5638, n5639, n5640, n5641,
    n5642, n5643, n5644, n5645, n5646, n5647,
    n5648, n5649, n5650, n5651, n5652, n5653,
    n5654, n5655, n5656, n5657, n5658, n5659,
    n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5670, n5671,
    n5672, n5673, n5674, n5675, n5676, n5677,
    n5678, n5679, n5680, n5681, n5682, n5683,
    n5684, n5685, n5686, n5687, n5688, n5689,
    n5690, n5691, n5692, n5693, n5694, n5695,
    n5696, n5697, n5698, n5699, n5700, n5701,
    n5702, n5703, n5704, n5705, n5706, n5707,
    n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5716, n5717, n5718, n5719,
    n5720, n5721, n5722, n5723, n5724, n5725,
    n5726, n5727, n5728, n5729, n5730, n5731,
    n5732, n5733, n5734, n5735, n5736, n5737,
    n5738, n5739, n5740, n5741, n5742, n5743,
    n5744, n5745, n5746, n5747, n5748, n5749,
    n5750, n5751, n5752, n5753, n5754, n5755,
    n5756, n5757, n5758, n5759, n5760, n5761,
    n5762, n5763, n5764, n5765, n5766, n5767,
    n5768, n5769, n5770, n5771, n5772, n5773,
    n5774, n5775, n5776, n5777, n5778, n5779,
    n5780, n5781, n5782, n5783, n5784, n5785,
    n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797,
    n5798, n5799, n5800, n5801, n5802, n5803,
    n5804, n5805, n5806, n5807, n5808, n5809,
    n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5817, n5818, n5819, n5820, n5821,
    n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839,
    n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857,
    n5858, n5859, n5860, n5861, n5862, n5863,
    n5864, n5865, n5866, n5867, n5868, n5869,
    n5870, n5871, n5872, n5873, n5874, n5875,
    n5876, n5877, n5878, n5879, n5880, n5881,
    n5882, n5883, n5884, n5885, n5886, n5887,
    n5888, n5889, n5890, n5891, n5892, n5893,
    n5894, n5895, n5896, n5897, n5898, n5899,
    n5900, n5901, n5902, n5903, n5904, n5905,
    n5906, n5907, n5908, n5909, n5910, n5911,
    n5912, n5913, n5914, n5915, n5916, n5917,
    n5918, n5919, n5920, n5921, n5922, n5923,
    n5924, n5925, n5926, n5927, n5928, n5929,
    n5930, n5931, n5932, n5933, n5934, n5935,
    n5936, n5937, n5938, n5939, n5940, n5941,
    n5942, n5943, n5944, n5945, n5946, n5947,
    n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5958, n5959,
    n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977,
    n5978, n5979, n5980, n5981, n5982, n5983,
    n5984, n5985, n5986, n5987, n5988, n5989,
    n5990, n5991, n5992, n5993, n5994, n5995,
    n5996, n5997, n5998, n5999, n6000, n6001,
    n6002, n6003, n6004, n6005, n6006, n6007,
    n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019,
    n6020, n6021, n6022, n6023, n6024, n6025,
    n6026, n6027, n6028, n6029, n6030, n6031,
    n6032, n6033, n6034, n6035, n6036, n6037,
    n6038, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049,
    n6050, n6051, n6052, n6053, n6054, n6055,
    n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067,
    n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079,
    n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097,
    n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151,
    n6152, n6153, n6154, n6155, n6156, n6157,
    n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175,
    n6176, n6177, n6178, n6179, n6180, n6181,
    n6182, n6183, n6184, n6185, n6186, n6187,
    n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6203, n6204, n6205,
    n6206, n6207, n6208, n6209, n6210, n6211,
    n6212, n6213, n6214, n6215, n6216, n6217,
    n6218, n6219, n6220, n6221, n6222, n6223,
    n6224, n6225, n6226, n6227, n6228, n6229,
    n6230, n6231, n6232, n6233, n6234, n6235,
    n6236, n6237, n6238, n6239, n6240, n6241,
    n6242, n6243, n6244, n6245, n6246, n6247,
    n6248, n6249, n6250, n6251, n6252, n6253,
    n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271,
    n6272, n6273, n6274, n6275, n6276, n6277,
    n6278, n6279, n6280, n6281, n6282, n6283,
    n6284, n6285, n6286, n6287, n6288, n6289,
    n6290, n6291, n6292, n6293, n6294, n6295,
    n6296, n6297, n6298, n6299, n6300, n6301,
    n6302, n6303, n6304, n6305, n6306, n6307,
    n6308, n6309, n6310, n6311, n6312, n6313,
    n6314, n6315, n6316, n6317, n6318, n6319,
    n6320, n6321, n6322, n6323, n6324, n6325,
    n6326, n6327, n6328, n6329, n6330, n6331,
    n6332, n6333, n6334, n6335, n6336, n6337,
    n6338, n6339, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349,
    n6350, n6351, n6352, n6353, n6354, n6355,
    n6356, n6357, n6358, n6359, n6360, n6361,
    n6362, n6363, n6364, n6365, n6366, n6367,
    n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379,
    n6380, n6381, n6382, n6383, n6384, n6385,
    n6386, n6387, n6388, n6389, n6390, n6391,
    n6392, n6393, n6394, n6395, n6396, n6397,
    n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409,
    n6410, n6411, n6412, n6413, n6414, n6415,
    n6416, n6417, n6418, n6419, n6420, n6421,
    n6422, n6423, n6424, n6425, n6426, n6427,
    n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6437, n6438, n6439,
    n6440, n6441, n6442, n6443, n6444, n6445,
    n6446, n6447, n6448, n6449, n6450, n6451,
    n6452, n6453, n6454, n6455, n6456, n6457,
    n6458, n6459, n6460, n6461, n6462, n6463,
    n6464, n6465, n6466, n6467, n6468, n6469,
    n6470, n6471, n6472, n6473, n6474, n6475,
    n6476, n6477, n6478, n6479, n6480, n6481,
    n6482, n6483, n6484, n6485, n6486, n6487,
    n6488, n6489, n6490, n6491, n6492, n6493,
    n6494, n6495, n6496, n6497, n6498, n6499,
    n6500, n6501, n6502, n6503, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511,
    n6512, n6513, n6514, n6515, n6516, n6517,
    n6518, n6519, n6520, n6521, n6522, n6523,
    n6524, n6525, n6526, n6527, n6528, n6529,
    n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541,
    n6542, n6543, n6544, n6545, n6546, n6547,
    n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571,
    n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601,
    n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649,
    n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661,
    n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691,
    n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721,
    n6722, n6723, n6724, n6725, n6726, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751,
    n6752, n6753, n6754, n6755, n6756, n6757,
    n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781,
    n6782, n6783, n6784, n6785, n6786, n6787,
    n6788, n6789, n6790, n6791, n6792, n6793,
    n6794, n6795, n6796, n6797, n6798, n6799,
    n6800, n6801, n6802, n6803, n6804, n6805,
    n6806, n6807, n6808, n6809, n6810, n6811,
    n6812, n6813, n6814, n6815, n6816, n6817,
    n6818, n6819, n6820, n6821, n6822, n6823,
    n6824, n6825, n6826, n6827, n6828, n6829,
    n6830, n6831, n6832, n6833, n6834, n6835,
    n6836, n6837, n6838, n6839, n6840, n6841,
    n6842, n6843, n6844, n6845, n6846, n6847,
    n6848, n6849, n6850, n6851, n6852, n6853,
    n6854, n6855, n6856, n6857, n6858, n6859,
    n6860, n6861, n6862, n6863, n6864, n6865,
    n6866, n6867, n6868, n6869, n6870, n6871,
    n6872, n6873, n6874, n6875, n6876, n6877,
    n6878, n6879, n6880, n6881, n6882, n6883,
    n6884, n6885, n6886, n6887, n6888, n6889,
    n6890, n6891, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901,
    n6902, n6903, n6904, n6905, n6906, n6907,
    n6908, n6909, n6910, n6911, n6912, n6913,
    n6914, n6915, n6916, n6917, n6918, n6919,
    n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931,
    n6932, n6933, n6934, n6935, n6936, n6937,
    n6938, n6939, n6940, n6941, n6942, n6943,
    n6944, n6945, n6946, n6947, n6948, n6949,
    n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961,
    n6962, n6963, n6964, n6965, n6966, n6967,
    n6968, n6969, n6970, n6971, n6972, n6973,
    n6974, n6975, n6976, n6977, n6978, n6979,
    n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991,
    n6992, n6993, n6994, n6995, n6996, n6997,
    n6998, n6999, n7000, n7001, n7002, n7003,
    n7004, n7005, n7006, n7007, n7008, n7009,
    n7010, n7011, n7012, n7013, n7014, n7015,
    n7016, n7017, n7018, n7019, n7020, n7021,
    n7022, n7023, n7024, n7025, n7026, n7027,
    n7028, n7029, n7030, n7031, n7032, n7033,
    n7034, n7035, n7036, n7037, n7038, n7039,
    n7040, n7041, n7042, n7043, n7044, n7045,
    n7046, n7047, n7048, n7049, n7050, n7051,
    n7052, n7053, n7054, n7055, n7056, n7057,
    n7058, n7059, n7060, n7061, n7062, n7063,
    n7064, n7065, n7066, n7067, n7068, n7069,
    n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081,
    n7082, n7083, n7084, n7085, n7086, n7087,
    n7088, n7089, n7090, n7091, n7092, n7093,
    n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7101, n7102, n7103, n7104, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111,
    n7112, n7113, n7114, n7115, n7116, n7117,
    n7118, n7119, n7120, n7121, n7122, n7123,
    n7124, n7125, n7126, n7127, n7128, n7129,
    n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141,
    n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153,
    n7154, n7155, n7156, n7157, n7158, n7159,
    n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171,
    n7172, n7173, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7229, n7230, n7231,
    n7232, n7233, n7234, n7235, n7236, n7237,
    n7238, n7239, n7240, n7241, n7242, n7243,
    n7244, n7245, n7246, n7247, n7248, n7249,
    n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7260, n7261,
    n7262, n7263, n7264, n7265, n7266, n7267,
    n7268, n7269, n7270, n7271, n7272, n7273,
    n7274, n7275, n7276, n7277, n7278, n7279,
    n7280, n7281, n7282, n7283, n7284, n7285,
    n7286, n7287, n7288, n7289, n7290, n7291,
    n7292, n7293, n7294, n7295, n7296, n7297,
    n7298, n7299, n7300, n7301, n7302, n7303,
    n7304, n7305, n7306, n7307, n7308, n7309,
    n7310, n7311, n7312, n7313, n7314, n7315,
    n7316, n7317, n7318, n7319, n7320, n7321,
    n7322, n7323, n7324, n7325, n7326, n7327,
    n7328, n7329, n7330, n7331, n7332, n7333,
    n7334, n7335, n7336, n7337, n7338, n7339,
    n7340, n7341, n7342, n7343, n7344, n7345,
    n7346, n7347, n7348, n7349, n7350, n7351,
    n7352, n7353, n7354, n7355, n7356, n7357,
    n7358, n7359, n7360, n7361, n7362, n7363,
    n7364, n7365, n7366, n7367, n7368, n7369,
    n7370, n7371, n7372, n7373, n7374, n7375,
    n7376, n7377, n7378, n7379, n7380, n7381,
    n7382, n7383, n7384, n7385, n7386, n7387,
    n7388, n7389, n7390, n7391, n7392, n7393,
    n7394, n7395, n7396, n7397, n7398, n7399,
    n7400, n7401, n7402, n7403, n7404, n7405,
    n7406, n7407, n7408, n7409, n7410, n7411,
    n7412, n7413, n7414, n7415, n7416, n7417,
    n7418, n7419, n7420, n7421, n7422, n7423,
    n7424, n7425, n7426, n7427, n7428, n7429,
    n7430, n7431, n7432, n7433, n7434, n7435,
    n7436, n7437, n7438, n7439, n7440, n7441,
    n7442, n7443, n7444, n7445, n7446, n7447,
    n7448, n7449, n7450, n7451, n7452, n7453,
    n7454, n7455, n7456, n7457, n7458, n7459,
    n7460, n7461, n7462, n7463, n7464, n7465,
    n7466, n7467, n7468, n7469, n7470, n7471,
    n7472, n7473, n7474, n7475, n7476, n7477,
    n7478, n7479, n7480, n7481, n7482, n7483,
    n7484, n7485, n7486, n7487, n7488, n7489,
    n7490, n7491, n7492, n7493, n7494, n7495,
    n7496, n7497, n7498, n7499, n7500, n7501,
    n7502, n7503, n7504, n7505, n7506, n7507,
    n7508, n7509, n7510, n7511, n7512, n7513,
    n7514, n7515, n7516, n7517, n7518, n7519,
    n7520, n7521, n7522, n7523, n7524, n7525,
    n7526, n7527, n7528, n7529, n7530, n7531,
    n7532, n7533, n7534, n7535, n7536, n7537,
    n7538, n7539, n7540, n7541, n7542, n7543,
    n7544, n7545, n7546, n7547, n7548, n7549,
    n7550, n7551, n7552, n7553, n7554, n7555,
    n7556, n7557, n7558, n7559, n7560, n7561,
    n7562, n7563, n7564, n7565, n7566, n7567,
    n7568, n7569, n7570, n7571, n7572, n7573,
    n7574, n7575, n7576, n7577, n7578, n7579,
    n7580, n7581, n7582, n7583, n7584, n7585,
    n7586, n7587, n7588, n7589, n7590, n7591,
    n7592, n7593, n7594, n7595, n7596, n7597,
    n7598, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7607, n7608, n7609,
    n7610, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621,
    n7622, n7623, n7624, n7625, n7626, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633,
    n7634, n7635, n7636, n7637, n7638, n7639,
    n7640, n7641, n7642, n7643, n7644, n7645,
    n7646, n7647, n7648, n7649, n7650, n7651,
    n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663,
    n7664, n7665, n7666, n7667, n7668, n7669,
    n7670, n7671, n7672, n7673, n7674, n7675,
    n7676, n7677, n7678, n7679, n7680, n7681,
    n7682, n7683, n7684, n7685, n7686, n7687,
    n7688, n7689, n7690, n7691, n7692, n7693,
    n7694, n7695, n7696, n7697, n7698, n7699,
    n7700, n7701, n7702, n7703, n7704, n7705,
    n7706, n7707, n7708, n7709, n7710, n7711,
    n7712, n7713, n7714, n7715, n7716, n7717,
    n7718, n7719, n7720, n7721, n7722, n7723,
    n7724, n7725, n7726, n7727, n7728, n7729,
    n7730, n7731, n7732, n7733, n7734, n7735,
    n7736, n7737, n7738, n7739, n7740, n7741,
    n7742, n7743, n7744, n7745, n7746, n7747,
    n7748, n7749, n7750, n7751, n7752, n7753,
    n7754, n7755, n7756, n7757, n7758, n7759,
    n7760, n7761, n7762, n7763, n7764, n7765,
    n7766, n7767, n7768, n7769, n7770, n7771,
    n7772, n7773, n7774, n7775, n7776, n7777,
    n7778, n7779, n7780, n7781, n7782, n7783,
    n7784, n7785, n7786, n7787, n7788, n7789,
    n7790, n7791, n7792, n7793, n7794, n7795,
    n7796, n7797, n7798, n7799, n7800, n7801,
    n7802, n7803, n7804, n7805, n7806, n7807,
    n7808, n7809, n7810, n7811, n7812, n7813,
    n7814, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825,
    n7826, n7827, n7828, n7829, n7830, n7831,
    n7832, n7833, n7834, n7835, n7836, n7837,
    n7838, n7839, n7840, n7841, n7842, n7843,
    n7844, n7845, n7846, n7847, n7848, n7849,
    n7850, n7851, n7852, n7853, n7854, n7855,
    n7856, n7857, n7858, n7859, n7860, n7861,
    n7862, n7863, n7864, n7865, n7866, n7867,
    n7868, n7869, n7870, n7871, n7872, n7873,
    n7874, n7875, n7876, n7877, n7878, n7879,
    n7880, n7881, n7882, n7883, n7884, n7885,
    n7886, n7887, n7888, n7889, n7890, n7891,
    n7892, n7893, n7894, n7895, n7896, n7897,
    n7898, n7899, n7900, n7901, n7902, n7903,
    n7904, n7905, n7906, n7907, n7908, n7909,
    n7910, n7911, n7912, n7913, n7914, n7915,
    n7916, n7917, n7918, n7919, n7920, n7921,
    n7922, n7923, n7924, n7925, n7926, n7927,
    n7928, n7929, n7930, n7931, n7932, n7933,
    n7934, n7935, n7936, n7937, n7938, n7939,
    n7940, n7941, n7942, n7943, n7944, n7945,
    n7946, n7947, n7948, n7949, n7950, n7951,
    n7952, n7953, n7954, n7955, n7956, n7957,
    n7958, n7959, n7960, n7961, n7962, n7963,
    n7964, n7965, n7966, n7967, n7968, n7969,
    n7970, n7971, n7972, n7973, n7974, n7975,
    n7976, n7977, n7978, n7979, n7980, n7981,
    n7982, n7983, n7984, n7985, n7986, n7987,
    n7988, n7989, n7990, n7991, n7992, n7993,
    n7994, n7995, n7996, n7997, n7998, n7999,
    n8000, n8001, n8002, n8003, n8004, n8005,
    n8006, n8007, n8008, n8009, n8010, n8011,
    n8012, n8013, n8014, n8015, n8016, n8017,
    n8018, n8019, n8020, n8021, n8022, n8023,
    n8024, n8025, n8026, n8027, n8028, n8029,
    n8030, n8031, n8032, n8033, n8034, n8035,
    n8036, n8037, n8038, n8039, n8040, n8041,
    n8042, n8043, n8044, n8045, n8046, n8047,
    n8048, n8049, n8050, n8051, n8052, n8053,
    n8054, n8055, n8056, n8057, n8058, n8059,
    n8060, n8061, n8062, n8063, n8064, n8065,
    n8066, n8067, n8068, n8069, n8070, n8071,
    n8072, n8073, n8074, n8075, n8076, n8077,
    n8078, n8079, n8080, n8081, n8082, n8083,
    n8084, n8085, n8086, n8087, n8088, n8089,
    n8090, n8091, n8092, n8093, n8094, n8095,
    n8096, n8097, n8098, n8099, n8100, n8101,
    n8102, n8103, n8104, n8105, n8106, n8107,
    n8108, n8109, n8110, n8111, n8112, n8113,
    n8114, n8115, n8116, n8117, n8118, n8119,
    n8120, n8121, n8122, n8123, n8124, n8125,
    n8126, n8127, n8128, n8129, n8130, n8131,
    n8132, n8133, n8134, n8135, n8136, n8137,
    n8138, n8139, n8140, n8141, n8142, n8143,
    n8144, n8145, n8146, n8147, n8148, n8149,
    n8150, n8151, n8152, n8153, n8154, n8155,
    n8156, n8157, n8158, n8159, n8160, n8161,
    n8162, n8163, n8164, n8165, n8166, n8167,
    n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8176, n8177, n8178, n8179,
    n8180, n8181, n8182, n8183, n8184, n8185,
    n8186, n8187, n8188, n8189, n8190, n8191,
    n8192, n8193, n8194, n8195, n8196, n8197,
    n8198, n8199, n8200, n8201, n8202, n8203,
    n8204, n8205, n8206, n8207, n8208, n8209,
    n8210, n8211, n8212, n8213, n8214, n8215,
    n8216, n8217, n8218, n8219, n8220, n8221,
    n8222, n8223, n8224, n8225, n8226, n8227,
    n8228, n8229, n8230, n8231, n8232, n8233,
    n8234, n8235, n8236, n8237, n8238, n8239,
    n8240, n8241, n8242, n8243, n8244, n8245,
    n8246, n8247, n8248, n8249, n8250, n8251,
    n8252, n8253, n8254, n8255, n8256, n8257,
    n8258, n8259, n8260, n8261, n8262, n8263,
    n8264, n8265, n8266, n8267, n8268, n8269,
    n8270, n8271, n8272, n8273, n8274, n8275,
    n8276, n8277, n8278, n8279, n8280, n8281,
    n8282, n8283, n8284, n8285, n8286, n8287,
    n8288, n8289, n8290, n8291, n8292, n8293,
    n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8301, n8302, n8303, n8304, n8305,
    n8306, n8307, n8308, n8309, n8310, n8311,
    n8312, n8313, n8314, n8315, n8316, n8317,
    n8318, n8319, n8320, n8321, n8322, n8323,
    n8324, n8325, n8326, n8327, n8328, n8329,
    n8330, n8331, n8332, n8333, n8334, n8335,
    n8336, n8337, n8338, n8339, n8340, n8341,
    n8342, n8343, n8344, n8345, n8346, n8347,
    n8348, n8349, n8350, n8351, n8352, n8353,
    n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8361, n8362, n8363, n8364, n8365,
    n8366, n8367, n8368, n8369, n8370, n8371,
    n8372, n8373, n8374, n8375, n8376, n8377,
    n8378, n8379, n8380, n8381, n8382, n8383,
    n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8392, n8393, n8394, n8395,
    n8396, n8397, n8398, n8399, n8400, n8401,
    n8402, n8403, n8404, n8405, n8406, n8407,
    n8408, n8409, n8410, n8411, n8412, n8413,
    n8414, n8415, n8416, n8417, n8418, n8419,
    n8420, n8421, n8422, n8423, n8424, n8425,
    n8426, n8427, n8428, n8429, n8430, n8431,
    n8432, n8433, n8434, n8435, n8436, n8437,
    n8438, n8439, n8440, n8441, n8442, n8443,
    n8444, n8445, n8446, n8447, n8448, n8449,
    n8450, n8451, n8452, n8453, n8454, n8455,
    n8456, n8457, n8458, n8459, n8460, n8461,
    n8462, n8463, n8464, n8465, n8466, n8467,
    n8468, n8469, n8470, n8471, n8472, n8473,
    n8474, n8475, n8476, n8477, n8478, n8479,
    n8480, n8481, n8482, n8483, n8484, n8485,
    n8486, n8487, n8488, n8489, n8490, n8491,
    n8492, n8493, n8494, n8495, n8496, n8497,
    n8498, n8499, n8500, n8501, n8502, n8503,
    n8504, n8505, n8506, n8507, n8508, n8509,
    n8510, n8511, n8512, n8513, n8514, n8515,
    n8516, n8517, n8518, n8519, n8520, n8521,
    n8522, n8523, n8524, n8525, n8526, n8527,
    n8528, n8529, n8530, n8531, n8532, n8533,
    n8534, n8535, n8536, n8537, n8538, n8539,
    n8540, n8541, n8542, n8543, n8544, n8545,
    n8546, n8547, n8548, n8549, n8550, n8551,
    n8552, n8553, n8554, n8555, n8556, n8557,
    n8558, n8559, n8560, n8561, n8562, n8563,
    n8564, n8565, n8566, n8567, n8568, n8569,
    n8570, n8571, n8572, n8573, n8574, n8575,
    n8576, n8577, n8578, n8579, n8580, n8581,
    n8582, n8583, n8584, n8585, n8586, n8587,
    n8588, n8589, n8590, n8591, n8592, n8593,
    n8594, n8595, n8596, n8597, n8598, n8599,
    n8600, n8601, n8602, n8603, n8604, n8605,
    n8606, n8607, n8608, n8609, n8610, n8611,
    n8612, n8613, n8614, n8615, n8616, n8617,
    n8618, n8619, n8620, n8621, n8622, n8623,
    n8624, n8625, n8626, n8627, n8628, n8629,
    n8630, n8631, n8632, n8633, n8634, n8635,
    n8636, n8637, n8638, n8639, n8640, n8641,
    n8642, n8643, n8644, n8645, n8646, n8647,
    n8648, n8649, n8650, n8651, n8652, n8653,
    n8654, n8655, n8656, n8657, n8658, n8659,
    n8660, n8661, n8662, n8663, n8664, n8665,
    n8666, n8667, n8668, n8669, n8670, n8671,
    n8672, n8673, n8674, n8675, n8676, n8677,
    n8678, n8679, n8680, n8681, n8682, n8683,
    n8684, n8685, n8686, n8687, n8688, n8689,
    n8690, n8691, n8692, n8693, n8694, n8695,
    n8696, n8697, n8698, n8699, n8700, n8701,
    n8702, n8703, n8704, n8705, n8706, n8707,
    n8708, n8709, n8710, n8711, n8712, n8713,
    n8714, n8715, n8716, n8717, n8718, n8719,
    n8720, n8721, n8722, n8723, n8724, n8725,
    n8726, n8727, n8728, n8729, n8730, n8731,
    n8732, n8733, n8734, n8735, n8736, n8737,
    n8738, n8739, n8740, n8741, n8742, n8743,
    n8744, n8745, n8746, n8747, n8748, n8749,
    n8750, n8751, n8752, n8753, n8754, n8755,
    n8756, n8757, n8758, n8759, n8760, n8761,
    n8762, n8763, n8764, n8765, n8766, n8767,
    n8768, n8769, n8770, n8771, n8772, n8773,
    n8774, n8775, n8776, n8777, n8778, n8779,
    n8780, n8781, n8782, n8783, n8784, n8785,
    n8786, n8787, n8788, n8789, n8790, n8791,
    n8792, n8793, n8794, n8795, n8796, n8797,
    n8798, n8799, n8800, n8801, n8802, n8803,
    n8804, n8805, n8806, n8807, n8808, n8809,
    n8810, n8811, n8812, n8813, n8814, n8815,
    n8816, n8817, n8818, n8819, n8820, n8821,
    n8822, n8823, n8824, n8825, n8826, n8827,
    n8828, n8829, n8830, n8831, n8832, n8833,
    n8834, n8835, n8836, n8837, n8838, n8839,
    n8840, n8841, n8842, n8843, n8844, n8845,
    n8846, n8847, n8848, n8849, n8850, n8851,
    n8852, n8853, n8854, n8855, n8856, n8857,
    n8858, n8859, n8860, n8861, n8862, n8863,
    n8864, n8865, n8866, n8867, n8868, n8869,
    n8870, n8871, n8872, n8873, n8874, n8875,
    n8876, n8877, n8878, n8879, n8880, n8881,
    n8882, n8883, n8884, n8885, n8886, n8887,
    n8888, n8889, n8890, n8891, n8892, n8893,
    n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8908, n8909, n8910, n8911,
    n8912, n8913, n8914, n8915, n8916, n8917,
    n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8929,
    n8930, n8931, n8932, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941,
    n8942, n8943, n8944, n8945, n8946, n8947,
    n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959,
    n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971,
    n8972, n8973, n8974, n8975, n8976, n8977,
    n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001,
    n9002, n9003, n9004, n9005, n9006, n9007,
    n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019,
    n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031,
    n9032, n9033, n9034, n9035, n9036, n9037,
    n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121,
    n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151,
    n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271,
    n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289,
    n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301,
    n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319,
    n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331,
    n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349,
    n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361,
    n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373,
    n9374, n9375, n9376, n9377, n9378, n9379,
    n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391,
    n9392, n9393, n9394, n9395, n9396, n9397,
    n9398, n9399, n9400, n9401, n9402, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421,
    n9422, n9423, n9424, n9425, n9426, n9427,
    n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439,
    n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9457,
    n9458, n9459, n9460, n9461, n9462, n9463,
    n9464, n9465, n9466, n9467, n9468, n9469,
    n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481,
    n9482, n9483, n9484, n9485, n9486, n9487,
    n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9496, n9497, n9498, n9499,
    n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511,
    n9512, n9513, n9514, n9515, n9516, n9517,
    n9518, n9519, n9520, n9521, n9522, n9523,
    n9524, n9525, n9526, n9527, n9528, n9529,
    n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541,
    n9542, n9543, n9544, n9545, n9546, n9547,
    n9548, n9549, n9550, n9551, n9552, n9553,
    n9554, n9555, n9556, n9557, n9558, n9559,
    n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571,
    n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583,
    n9584, n9585, n9586, n9587, n9588, n9589,
    n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9597, n9598, n9599, n9600, n9601,
    n9602, n9603, n9604, n9605, n9606, n9607,
    n9608, n9609, n9610, n9611, n9612, n9613,
    n9614, n9615, n9616, n9617, n9618, n9619,
    n9620, n9621, n9622, n9623, n9624, n9625,
    n9626, n9627, n9628, n9629, n9630, n9631,
    n9632, n9633, n9634, n9635, n9636, n9637,
    n9638, n9639, n9640, n9641, n9642, n9643,
    n9644, n9645, n9646, n9647, n9648, n9649,
    n9650, n9651, n9652, n9653, n9654, n9655,
    n9656, n9657, n9658, n9659, n9660, n9661,
    n9662, n9663, n9664, n9665, n9666, n9667,
    n9668, n9669, n9670, n9671, n9672, n9673,
    n9674, n9675, n9676, n9677, n9678, n9679,
    n9680, n9681, n9682, n9683, n9684, n9685,
    n9686, n9687, n9688, n9689, n9690, n9691,
    n9692, n9693, n9694, n9695, n9696, n9697,
    n9698, n9699, n9700, n9701, n9702, n9703,
    n9704, n9705, n9706, n9707, n9708, n9709,
    n9710, n9711, n9712, n9713, n9714, n9715,
    n9716, n9717, n9718, n9719, n9720, n9721,
    n9722, n9723, n9724, n9725, n9726, n9727,
    n9728, n9729, n9730, n9731, n9732, n9733,
    n9734, n9735, n9736, n9737, n9738, n9739,
    n9740, n9741, n9742, n9743, n9744, n9745,
    n9746, n9747, n9748, n9749, n9750, n9751,
    n9752, n9753, n9754, n9755, n9756, n9757,
    n9758, n9759, n9760, n9761, n9762, n9763,
    n9764, n9765, n9766, n9767, n9768, n9769,
    n9770, n9771, n9772, n9773, n9774, n9775,
    n9776, n9777, n9778, n9779, n9780, n9781,
    n9782, n9783, n9784, n9785, n9786, n9787,
    n9788, n9789, n9790, n9791, n9792, n9793,
    n9794, n9795, n9796, n9797, n9798, n9799,
    n9800, n9801, n9802, n9803, n9804, n9805,
    n9806, n9807, n9808, n9809, n9810, n9811,
    n9812, n9813, n9814, n9815, n9816, n9817,
    n9818, n9819, n9820, n9821, n9822, n9823,
    n9824, n9825, n9826, n9827, n9828, n9829,
    n9830, n9831, n9832, n9833, n9834, n9835,
    n9836, n9837, n9838, n9839, n9840, n9841,
    n9842, n9843, n9844, n9845, n9846, n9847,
    n9848, n9849, n9850, n9851, n9852, n9853,
    n9854, n9855, n9856, n9857, n9858, n9859,
    n9860, n9861, n9862, n9863, n9864, n9865,
    n9866, n9867, n9868, n9869, n9870, n9871,
    n9872, n9873, n9874, n9875, n9876, n9877,
    n9878, n9879, n9880, n9881, n9882, n9883,
    n9884, n9885, n9886, n9887, n9888, n9889,
    n9890, n9891, n9892, n9893, n9894, n9895,
    n9896, n9897, n9898, n9899, n9900, n9901,
    n9902, n9903, n9904, n9905, n9906, n9907,
    n9908, n9909, n9910, n9911, n9912, n9913,
    n9914, n9915, n9916, n9917, n9918, n9919,
    n9920, n9921, n9922, n9923, n9924, n9925,
    n9926, n9927, n9928, n9929, n9930, n9931,
    n9932, n9933, n9934, n9935, n9936, n9937,
    n9938, n9939, n9940, n9941, n9942, n9943,
    n9944, n9945, n9946, n9947, n9948, n9949,
    n9950, n9951, n9952, n9953, n9954, n9955,
    n9956, n9957, n9958, n9959, n9960, n9961,
    n9962, n9963, n9964, n9965, n9966, n9967,
    n9968, n9969, n9970, n9971, n9972, n9973,
    n9974, n9975, n9976, n9977, n9978, n9979,
    n9980, n9981, n9982, n9983, n9984, n9985,
    n9986, n9987, n9988, n9989, n9990, n9991,
    n9992, n9993, n9994, n9995, n9996, n9997,
    n9998, n9999, n10000, n10001, n10002, n10003,
    n10004, n10005, n10006, n10007, n10008, n10009,
    n10010, n10011, n10012, n10013, n10014, n10015,
    n10016, n10017, n10018, n10019, n10020, n10021,
    n10022, n10023, n10024, n10025, n10026, n10027,
    n10028, n10029, n10030, n10031, n10032, n10033,
    n10034, n10035, n10036, n10037, n10038, n10039,
    n10040, n10041, n10042, n10043, n10044, n10045,
    n10046, n10047, n10048, n10049, n10050, n10051,
    n10052, n10053, n10054, n10055, n10056, n10057,
    n10058, n10059, n10060, n10061, n10062, n10063,
    n10064, n10065, n10066, n10067, n10068, n10069,
    n10070, n10071, n10072, n10073, n10074, n10075,
    n10076, n10077, n10078, n10079, n10080, n10081,
    n10082, n10083, n10084, n10085, n10086, n10087,
    n10088, n10089, n10090, n10091, n10092, n10093,
    n10094, n10095, n10096, n10097, n10098, n10099,
    n10100, n10101, n10102, n10103, n10104, n10105,
    n10106, n10107, n10108, n10109, n10110, n10111,
    n10112, n10113, n10114, n10115, n10116, n10117,
    n10118, n10119, n10120, n10121, n10122, n10123,
    n10124, n10125, n10126, n10127, n10128, n10129,
    n10130, n10131, n10132, n10133, n10134, n10135,
    n10136, n10137, n10138, n10139, n10140, n10141,
    n10142, n10143, n10144, n10145, n10146, n10147,
    n10148, n10149, n10150, n10151, n10152, n10153,
    n10154, n10155, n10156, n10157, n10158, n10159,
    n10160, n10161, n10162, n10163, n10164, n10165,
    n10166, n10167, n10168, n10169, n10170, n10171,
    n10172, n10173, n10174, n10175, n10176, n10177,
    n10178, n10179, n10180, n10181, n10182, n10183,
    n10184, n10185, n10186, n10187, n10188, n10189,
    n10190, n10191, n10192, n10193, n10194, n10195,
    n10196, n10197, n10198, n10199, n10200, n10201,
    n10202, n10203, n10204, n10205, n10206, n10207,
    n10208, n10209, n10210, n10211, n10212, n10213,
    n10214, n10215, n10216, n10217, n10218, n10219,
    n10220, n10221, n10222, n10223, n10224, n10225,
    n10226, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237,
    n10238, n10239, n10240, n10241, n10242, n10243,
    n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255,
    n10256, n10257, n10258, n10259, n10260, n10261,
    n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273,
    n10274, n10275, n10276, n10277, n10278, n10279,
    n10280, n10281, n10282, n10283, n10284, n10285,
    n10286, n10287, n10288, n10289, n10290, n10291,
    n10292, n10293, n10294, n10295, n10296, n10297,
    n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309,
    n10310, n10311, n10312, n10313, n10314, n10315,
    n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327,
    n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345,
    n10346, n10347, n10348, n10349, n10350, n10351,
    n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363,
    n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10397, n10398, n10399,
    n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411,
    n10412, n10413, n10414, n10415, n10416, n10417,
    n10418, n10419, n10420, n10421, n10422, n10423,
    n10424, n10425, n10426, n10427, n10428, n10429,
    n10430, n10431, n10432, n10433, n10434, n10435,
    n10436, n10437, n10438, n10439, n10440, n10441,
    n10442, n10443, n10444, n10445, n10446, n10447,
    n10448, n10449, n10450, n10451, n10452, n10453,
    n10454, n10455, n10456, n10457, n10458, n10459,
    n10460, n10461, n10462, n10463, n10464, n10465,
    n10466, n10467, n10468, n10469, n10470, n10471,
    n10472, n10473, n10474, n10475, n10476, n10477,
    n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10487, n10488, n10489,
    n10490, n10491, n10492, n10493, n10494, n10495,
    n10496, n10497, n10498, n10499, n10500, n10501,
    n10502, n10503, n10504, n10505, n10506, n10507,
    n10508, n10509, n10510, n10511, n10512, n10513,
    n10514, n10515, n10516, n10517, n10518, n10519,
    n10520, n10521, n10522, n10523, n10524, n10525,
    n10526, n10527, n10528, n10529, n10530, n10531,
    n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543,
    n10544, n10545, n10546, n10547, n10548, n10549,
    n10550, n10551, n10552, n10553, n10554, n10555,
    n10556, n10557, n10558, n10559, n10560, n10561,
    n10562, n10563, n10564, n10565, n10566, n10567,
    n10568, n10569, n10570, n10571, n10572, n10573,
    n10574, n10575, n10576, n10577, n10578, n10579,
    n10580, n10581, n10582, n10583, n10584, n10585,
    n10586, n10587, n10588, n10589, n10590, n10591,
    n10592, n10593, n10594, n10595, n10596, n10597,
    n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10606, n10607, n10608, n10609,
    n10610, n10611, n10612, n10613, n10614, n10615,
    n10616, n10617, n10618, n10619, n10620, n10621,
    n10622, n10623, n10624, n10625, n10626, n10627,
    n10628, n10629, n10630, n10631, n10632, n10633,
    n10634, n10635, n10636, n10637, n10638, n10639,
    n10640, n10641, n10642, n10643, n10644, n10645,
    n10646, n10647, n10648, n10649, n10650, n10651,
    n10652, n10653, n10654, n10655, n10656, n10657,
    n10658, n10659, n10660, n10661, n10662, n10663,
    n10664, n10665, n10666, n10667, n10668, n10669,
    n10670, n10671, n10672, n10673, n10674, n10675,
    n10676, n10677, n10678, n10679, n10680, n10681,
    n10682, n10683, n10684, n10685, n10686, n10687,
    n10688, n10689, n10690, n10691, n10692, n10693,
    n10694, n10695, n10696, n10697, n10698, n10699,
    n10700, n10701, n10702, n10703, n10704, n10705,
    n10706, n10707, n10708, n10709, n10710, n10711,
    n10712, n10713, n10714, n10715, n10716, n10717,
    n10718, n10719, n10720, n10721, n10722, n10723,
    n10724, n10725, n10726, n10727, n10728, n10729,
    n10730, n10731, n10732, n10733, n10734, n10735,
    n10736, n10737, n10738, n10739, n10740, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747,
    n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10759,
    n10760, n10761, n10762, n10763, n10764, n10765,
    n10766, n10767, n10768, n10769, n10770, n10771,
    n10772, n10773, n10774, n10775, n10776, n10777,
    n10778, n10779, n10780, n10781, n10782, n10783,
    n10784, n10785, n10786, n10787, n10788, n10789,
    n10790, n10791, n10792, n10793, n10794, n10795,
    n10796, n10797, n10798, n10799, n10800, n10801,
    n10802, n10803, n10804, n10805, n10806, n10807,
    n10808, n10809, n10810, n10811, n10812, n10813,
    n10814, n10815, n10816, n10817, n10818, n10819,
    n10820, n10821, n10822, n10823, n10824, n10825,
    n10826, n10827, n10828, n10829, n10830, n10831,
    n10832, n10833, n10834, n10835, n10836, n10837,
    n10838, n10839, n10840, n10841, n10842, n10843,
    n10844, n10845, n10846, n10847, n10848, n10849,
    n10850, n10851, n10852, n10853, n10854, n10855,
    n10856, n10857, n10858, n10859, n10860, n10861,
    n10862, n10863, n10864, n10865, n10866, n10867,
    n10868, n10869, n10870, n10871, n10872, n10873,
    n10874, n10875, n10876, n10877, n10878, n10879,
    n10880, n10881, n10882, n10883, n10884, n10885,
    n10886, n10887, n10888, n10889, n10890, n10891,
    n10892, n10893, n10894, n10895, n10896, n10897,
    n10898, n10899, n10900, n10901, n10902, n10903,
    n10904, n10905, n10906, n10907, n10908, n10909,
    n10910, n10911, n10912, n10913, n10914, n10915,
    n10916, n10917, n10918, n10919, n10920, n10921,
    n10922, n10923, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10945,
    n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963,
    n10964, n10965, n10966, n10967, n10968, n10969,
    n10970, n10971, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10981,
    n10982, n10983, n10984, n10985, n10986, n10987,
    n10988, n10989, n10990, n10991, n10992, n10993,
    n10994, n10995, n10996, n10997, n10998, n10999,
    n11000, n11001, n11002, n11003, n11004, n11005,
    n11006, n11007, n11008, n11009, n11010, n11011,
    n11012, n11013, n11014, n11015, n11016, n11017,
    n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11025, n11026, n11027, n11028, n11029,
    n11030, n11031, n11032, n11033, n11034, n11035,
    n11036, n11037, n11038, n11039, n11040, n11041,
    n11042, n11043, n11044, n11045, n11046, n11047,
    n11048, n11049, n11050, n11051, n11052, n11053,
    n11054, n11055, n11056, n11057, n11058, n11059,
    n11060, n11061, n11062, n11063, n11064, n11065,
    n11066, n11067, n11068, n11069, n11070, n11071,
    n11072, n11073, n11074, n11075, n11076, n11077,
    n11078, n11079, n11080, n11081, n11082, n11083,
    n11084, n11085, n11086, n11087, n11088, n11089,
    n11090, n11091, n11092, n11093, n11094, n11095,
    n11096, n11097, n11098, n11099, n11100, n11101,
    n11102, n11103, n11104, n11105, n11106, n11107,
    n11108, n11109, n11110, n11111, n11112, n11113,
    n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125,
    n11126, n11127, n11128, n11129, n11130, n11131,
    n11132, n11133, n11134, n11135, n11136, n11137,
    n11138, n11139, n11140, n11141, n11142, n11143,
    n11144, n11145, n11146, n11147, n11148, n11149,
    n11150, n11151, n11152, n11153, n11154, n11155,
    n11156, n11157, n11158, n11159, n11160, n11161,
    n11162, n11163, n11164, n11165, n11166, n11167,
    n11168, n11169, n11170, n11171, n11172, n11173,
    n11174, n11175, n11176, n11177, n11178, n11179,
    n11180, n11181, n11182, n11183, n11184, n11185,
    n11186, n11187, n11188, n11189, n11190, n11191,
    n11192, n11193, n11194, n11195, n11196, n11197,
    n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209,
    n11210, n11211, n11212, n11213, n11214, n11215,
    n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227,
    n11228, n11229, n11230, n11231, n11232, n11233,
    n11234, n11235, n11236, n11237, n11238, n11239,
    n11240, n11241, n11242, n11243, n11244, n11245,
    n11246, n11247, n11248, n11249, n11250, n11251,
    n11252, n11253, n11254, n11255, n11256, n11257,
    n11258, n11259, n11260, n11261, n11262, n11263,
    n11264, n11265, n11266, n11267, n11268, n11269,
    n11270, n11271, n11272, n11273, n11274, n11275,
    n11276, n11277, n11278, n11279, n11280, n11281,
    n11282, n11283, n11284, n11285, n11286, n11287,
    n11288, n11289, n11290, n11291, n11292, n11293,
    n11294, n11295, n11296, n11297, n11298, n11299,
    n11300, n11301, n11302, n11303, n11304, n11305,
    n11306, n11307, n11308, n11309, n11310, n11311,
    n11312, n11313, n11314, n11315, n11316, n11317,
    n11318, n11319, n11320, n11321, n11322, n11323,
    n11324, n11325, n11326, n11327, n11328, n11329,
    n11330, n11331, n11332, n11333, n11334, n11335,
    n11336, n11337, n11338, n11339, n11340, n11341,
    n11342, n11343, n11344, n11345, n11346, n11347,
    n11348, n11349, n11350, n11351, n11352, n11353,
    n11354, n11355, n11356, n11357, n11358, n11359,
    n11360, n11361, n11362, n11363, n11364, n11365,
    n11366, n11367, n11368, n11369, n11370, n11371,
    n11372, n11373, n11374, n11375, n11376, n11377,
    n11378, n11379, n11380, n11381, n11382, n11383,
    n11384, n11385, n11386, n11387, n11388, n11389,
    n11390, n11391, n11392, n11393, n11394, n11395,
    n11396, n11397, n11398, n11399, n11400, n11401,
    n11402, n11403, n11404, n11405, n11406, n11407,
    n11408, n11409, n11410, n11411, n11412, n11413,
    n11414, n11415, n11416, n11417, n11418, n11419,
    n11420, n11421, n11422, n11423, n11424, n11425,
    n11426, n11427, n11428, n11429, n11430, n11431,
    n11432, n11433, n11434, n11435, n11436, n11437,
    n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449,
    n11450, n11451, n11452, n11453, n11454, n11455,
    n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473,
    n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497,
    n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515,
    n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527,
    n11528, n11529, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545,
    n11546, n11547, n11548, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575,
    n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11590, n11591, n11592, n11593,
    n11594, n11595, n11596, n11597, n11598, n11599,
    n11600, n11601, n11602, n11603, n11604, n11605,
    n11606, n11607, n11608, n11609, n11610, n11611,
    n11612, n11613, n11614, n11615, n11616, n11617,
    n11618, n11619, n11620, n11621, n11622, n11623,
    n11624, n11625, n11626, n11627, n11628, n11629,
    n11630, n11631, n11632, n11633, n11634, n11635,
    n11636, n11637, n11638, n11639, n11640, n11641,
    n11642, n11643, n11644, n11645, n11646, n11647,
    n11648, n11649, n11650, n11651, n11652, n11653,
    n11654, n11655, n11656, n11657, n11658, n11659,
    n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671,
    n11672, n11673, n11674, n11675, n11676, n11677,
    n11678, n11679, n11680, n11681, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11693, n11694, n11695,
    n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11706, n11707,
    n11708, n11709, n11710, n11711, n11712, n11713,
    n11714, n11715, n11716, n11717, n11718, n11719,
    n11720, n11721, n11722, n11723, n11724, n11725,
    n11726, n11727, n11728, n11729, n11730, n11731,
    n11732, n11733, n11734, n11735, n11736, n11737,
    n11738, n11739, n11740, n11741, n11742, n11743,
    n11744, n11745, n11746, n11747, n11748, n11749,
    n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761,
    n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779,
    n11780, n11781, n11782, n11783, n11784, n11785,
    n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797,
    n11798, n11799, n11800, n11801, n11802, n11803,
    n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815,
    n11816, n11817, n11818, n11819, n11820, n11821,
    n11822, n11823, n11824, n11825, n11826, n11827,
    n11828, n11829, n11830, n11831, n11832, n11833,
    n11834, n11835, n11836, n11837, n11838, n11839,
    n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11849, n11850, n11851,
    n11852, n11853, n11854, n11855, n11856, n11857,
    n11858, n11859, n11860, n11861, n11862, n11863,
    n11864, n11865, n11866, n11867, n11868, n11869,
    n11870, n11871, n11872, n11873, n11874, n11875,
    n11876, n11877, n11878, n11879, n11880, n11881,
    n11882, n11883, n11884, n11885, n11886, n11887,
    n11888, n11889, n11890, n11891, n11892, n11893,
    n11894, n11895, n11896, n11897, n11898, n11899,
    n11900, n11901, n11902, n11903, n11904, n11905,
    n11906, n11907, n11908, n11909, n11910, n11911,
    n11912, n11913, n11914, n11915, n11916, n11917,
    n11918, n11919, n11920, n11921, n11922, n11923,
    n11924, n11925, n11926, n11927, n11928, n11929,
    n11930, n11931, n11932, n11933, n11934, n11935,
    n11936, n11937, n11938, n11939, n11940, n11941,
    n11942, n11943, n11944, n11945, n11946, n11947,
    n11948, n11949, n11950, n11951, n11952, n11953,
    n11954, n11955, n11956, n11957, n11958, n11959,
    n11960, n11961, n11962, n11963, n11964, n11965,
    n11966, n11967, n11968, n11969, n11970, n11971,
    n11972, n11973, n11974, n11975, n11976, n11977,
    n11978, n11979, n11980, n11981, n11982, n11983,
    n11984, n11985, n11986, n11987, n11988, n11989,
    n11990, n11991, n11992, n11993, n11994, n11995,
    n11996, n11997, n11998, n11999, n12000, n12001,
    n12002, n12003, n12004, n12005, n12006, n12007,
    n12008, n12009, n12010, n12011, n12012, n12013,
    n12014, n12015, n12016, n12017, n12018, n12019,
    n12020, n12021, n12022, n12023, n12024, n12025,
    n12026, n12027, n12028, n12029, n12030, n12031,
    n12032, n12033, n12034, n12035, n12036, n12037,
    n12038, n12039, n12040, n12041, n12042, n12043,
    n12044, n12045, n12046, n12047, n12048, n12049,
    n12050, n12051, n12052, n12053, n12054, n12055,
    n12056, n12057, n12058, n12059, n12060, n12061,
    n12062, n12063, n12064, n12065, n12066, n12067,
    n12068, n12069, n12070, n12071, n12072, n12073,
    n12074, n12075, n12076, n12077, n12078, n12079,
    n12080, n12081, n12082, n12083, n12084, n12085,
    n12086, n12087, n12088, n12089, n12090, n12091,
    n12092, n12093, n12094, n12095, n12096, n12097,
    n12098, n12099, n12100, n12101, n12102, n12103,
    n12104, n12105, n12106, n12107, n12108, n12109,
    n12110, n12111, n12112, n12113, n12114, n12115,
    n12116, n12117, n12118, n12119, n12120, n12121,
    n12122, n12123, n12124, n12125, n12126, n12127,
    n12128, n12129, n12130, n12131, n12132, n12133,
    n12134, n12135, n12136, n12137, n12138, n12139,
    n12140, n12141, n12142, n12143, n12144, n12145,
    n12146, n12147, n12148, n12149, n12150, n12151,
    n12152, n12153, n12154, n12155, n12156, n12157,
    n12158, n12159, n12160, n12161, n12162, n12163,
    n12164, n12165, n12166, n12167, n12168, n12169,
    n12170, n12171, n12172, n12173, n12174, n12175,
    n12176, n12177, n12178, n12179, n12180, n12181,
    n12182, n12183, n12184, n12185, n12186, n12187,
    n12188, n12189, n12190, n12191, n12192, n12193,
    n12194, n12195, n12196, n12197, n12198, n12199,
    n12200, n12201, n12202, n12203, n12204, n12205,
    n12206, n12207, n12208, n12209, n12210, n12211,
    n12212, n12213, n12214, n12215, n12216, n12217,
    n12218, n12219, n12220, n12221, n12222, n12223,
    n12224, n12225, n12226, n12227, n12228, n12229,
    n12230, n12231, n12232, n12233, n12234, n12235,
    n12236, n12237, n12238, n12239, n12240, n12241,
    n12242, n12243, n12244, n12245, n12246, n12247,
    n12248, n12249, n12250, n12251, n12252, n12253,
    n12254, n12255, n12256, n12257, n12258, n12259,
    n12260, n12261, n12262, n12263, n12264, n12265,
    n12266, n12267, n12268, n12269, n12270, n12271,
    n12272, n12273, n12274, n12275, n12276, n12277,
    n12278, n12279, n12280, n12281, n12282, n12283,
    n12284, n12285, n12286, n12287, n12288, n12289,
    n12290, n12291, n12292, n12293, n12294, n12295,
    n12296, n12297, n12298, n12299, n12300, n12301,
    n12302, n12303, n12304, n12305, n12306, n12307,
    n12308, n12309, n12310, n12311, n12312, n12313,
    n12314, n12315, n12316, n12317, n12318, n12319,
    n12320, n12321, n12322, n12323, n12324, n12325,
    n12326, n12327, n12328, n12329, n12330, n12331,
    n12332, n12333, n12334, n12335, n12336, n12337,
    n12338, n12339, n12340, n12341, n12342, n12343,
    n12344, n12345, n12346, n12347, n12348, n12349,
    n12350, n12351, n12352, n12353, n12354, n12355,
    n12356, n12357, n12358, n12359, n12360, n12361,
    n12362, n12363, n12364, n12365, n12366, n12367,
    n12368, n12369, n12370, n12371, n12372, n12373,
    n12374, n12375, n12376, n12377, n12378, n12379,
    n12380, n12381, n12382, n12383, n12384, n12385,
    n12386, n12387, n12388, n12389, n12390, n12391,
    n12392, n12393, n12394, n12395, n12396, n12397,
    n12398, n12399, n12400, n12401, n12402, n12403,
    n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415,
    n12416, n12417, n12418, n12419, n12420, n12421,
    n12422, n12423, n12424, n12425, n12426, n12427,
    n12428, n12429, n12430, n12431, n12432, n12433,
    n12434, n12435, n12436, n12437, n12438, n12439,
    n12440, n12441, n12442, n12443, n12444, n12445,
    n12446, n12447, n12448, n12449, n12450, n12451,
    n12452, n12453, n12454, n12455, n12456, n12457,
    n12458, n12459, n12460, n12461, n12462, n12463,
    n12464, n12465, n12466, n12467, n12468, n12469,
    n12470, n12471, n12472, n12473, n12474, n12475,
    n12476, n12477, n12478, n12479, n12480, n12481,
    n12482, n12483, n12484, n12485, n12486, n12487,
    n12488, n12489, n12490, n12491, n12492, n12493,
    n12494, n12495, n12496, n12497, n12498, n12499,
    n12500, n12501, n12502, n12503, n12504, n12505,
    n12506, n12507, n12508, n12509, n12510, n12511,
    n12512, n12513, n12514, n12515, n12516, n12517,
    n12518, n12519, n12520, n12521, n12522, n12523,
    n12524, n12525, n12526, n12527, n12528, n12529,
    n12530, n12531, n12532, n12533, n12534, n12535,
    n12536, n12537, n12538, n12539, n12540, n12541,
    n12542, n12543, n12544, n12545, n12546, n12547,
    n12548, n12549, n12550, n12551, n12552, n12553,
    n12554, n12555, n12556, n12557, n12558, n12559,
    n12560, n12561, n12562, n12563, n12564, n12565,
    n12566, n12567, n12568, n12569, n12570, n12571,
    n12572, n12573, n12574, n12575, n12576, n12577,
    n12578, n12579, n12580, n12581, n12582, n12583,
    n12584, n12585, n12586, n12587, n12588, n12589,
    n12590, n12591, n12592, n12593, n12594, n12595,
    n12596, n12597, n12598, n12599, n12600, n12601,
    n12602, n12603, n12604, n12605, n12606, n12607,
    n12608, n12609, n12610, n12611, n12612, n12613,
    n12614, n12615, n12616, n12617, n12618, n12619,
    n12620, n12621, n12622, n12623, n12624, n12625,
    n12626, n12627, n12628, n12629, n12630, n12631,
    n12632, n12633, n12634, n12635, n12636, n12637,
    n12638, n12639, n12640, n12641, n12642, n12643,
    n12644, n12645, n12646, n12647, n12648, n12649,
    n12650, n12651, n12652, n12653, n12654, n12655,
    n12656, n12657, n12658, n12659, n12660, n12661,
    n12662, n12663, n12664, n12665, n12666, n12667,
    n12668, n12669, n12670, n12671, n12672, n12673,
    n12674, n12675, n12676, n12677, n12678, n12679,
    n12680, n12681, n12682, n12683, n12684, n12685,
    n12686, n12687, n12688, n12689, n12690, n12691,
    n12692, n12693, n12694, n12695, n12696, n12697,
    n12698, n12699, n12700, n12701, n12702, n12703,
    n12704, n12705, n12706, n12707, n12708, n12709,
    n12710, n12711, n12712, n12713, n12714, n12715,
    n12716, n12717, n12718, n12719, n12720, n12721,
    n12722, n12723, n12724, n12725, n12726, n12727,
    n12728, n12729, n12730, n12731, n12732, n12733,
    n12734, n12735, n12736, n12737, n12738, n12739,
    n12740, n12741, n12742, n12743, n12744, n12745,
    n12746, n12747, n12748, n12749, n12750, n12751,
    n12752, n12753, n12754, n12755, n12756, n12757,
    n12758, n12759, n12760, n12761, n12762, n12763,
    n12764, n12765, n12766, n12767, n12768, n12769,
    n12770, n12771, n12772, n12773, n12774, n12775,
    n12776, n12777, n12778, n12779, n12780, n12781,
    n12782, n12783, n12784, n12785, n12786, n12787,
    n12788, n12789, n12790, n12791, n12792, n12793,
    n12794, n12795, n12796, n12797, n12798, n12799,
    n12800, n12801, n12802, n12803, n12804, n12805,
    n12806, n12807, n12808, n12809, n12810, n12811,
    n12812, n12813, n12814, n12815, n12816, n12817,
    n12818, n12819, n12820, n12821, n12822, n12823,
    n12824, n12825, n12826, n12827, n12828, n12829,
    n12830, n12831, n12832, n12833, n12834, n12835,
    n12836, n12837, n12838, n12839, n12840, n12841,
    n12842, n12843, n12844, n12845, n12846, n12847,
    n12848, n12849, n12850, n12851, n12852, n12853,
    n12854, n12855, n12856, n12857, n12858, n12859,
    n12860, n12861, n12862, n12863, n12864, n12865,
    n12866, n12867, n12868, n12869, n12870, n12871,
    n12872, n12873, n12874, n12875, n12876, n12877,
    n12878, n12879, n12880, n12881, n12882, n12883,
    n12884, n12885, n12886, n12887, n12888, n12889,
    n12890, n12891, n12892, n12893, n12894, n12895,
    n12896, n12897, n12898, n12899, n12900, n12901,
    n12902, n12903, n12904, n12905, n12906, n12907,
    n12908, n12909, n12910, n12911, n12912, n12913,
    n12914, n12915, n12916, n12917, n12918, n12919,
    n12920, n12921, n12922, n12923, n12924, n12925,
    n12926, n12927, n12928, n12929, n12930, n12931,
    n12932, n12933, n12934, n12935, n12936, n12937,
    n12938, n12939, n12940, n12941, n12942, n12943,
    n12944, n12945, n12946, n12947, n12948, n12949,
    n12950, n12951, n12952, n12953, n12954, n12955,
    n12956, n12957, n12958, n12959, n12960, n12961,
    n12962, n12963, n12964, n12965, n12966, n12967,
    n12968, n12969, n12970, n12971, n12972, n12973,
    n12974, n12975, n12976, n12977, n12978, n12979,
    n12980, n12981, n12982, n12983, n12984, n12985,
    n12986, n12987, n12988, n12989, n12990, n12991,
    n12992, n12993, n12994, n12995, n12996, n12997,
    n12998, n12999, n13000, n13001, n13002, n13003,
    n13004, n13005, n13006, n13007, n13008, n13009,
    n13010, n13011, n13012, n13013, n13014, n13015,
    n13016, n13017, n13018, n13019, n13020, n13021,
    n13022, n13023, n13024, n13025, n13026, n13027,
    n13028, n13029, n13030, n13031, n13032, n13033,
    n13034, n13035, n13036, n13037, n13038, n13039,
    n13040, n13041, n13042, n13043, n13044, n13045,
    n13046, n13047, n13048, n13049, n13050, n13051,
    n13052, n13053, n13054, n13055, n13056, n13057,
    n13058, n13059, n13060, n13061, n13062, n13063,
    n13064, n13065, n13066, n13067, n13068, n13069,
    n13070, n13071, n13072, n13073, n13074, n13075,
    n13076, n13077, n13078, n13079, n13080, n13081,
    n13082, n13083, n13084, n13085, n13086, n13087,
    n13088, n13089, n13090, n13091, n13092, n13093,
    n13094, n13095, n13096, n13097, n13098, n13099,
    n13100, n13101, n13102, n13103, n13104, n13105,
    n13106, n13107, n13108, n13109, n13110, n13111,
    n13112, n13113, n13114, n13115, n13116, n13117,
    n13118, n13119, n13120, n13121, n13122, n13123,
    n13124, n13125, n13126, n13127, n13128, n13129,
    n13130, n13131, n13132, n13133, n13134, n13135,
    n13136, n13137, n13138, n13139, n13140, n13141,
    n13142, n13143, n13144, n13145, n13146, n13147,
    n13148, n13149, n13150, n13151, n13152, n13153,
    n13154, n13155, n13156, n13157, n13158, n13159,
    n13160, n13161, n13162, n13163, n13164, n13165,
    n13166, n13167, n13168, n13169, n13170, n13171,
    n13172, n13173, n13174, n13175, n13176, n13177,
    n13178, n13179, n13180, n13181, n13182, n13183,
    n13184, n13185, n13186, n13187, n13188, n13189,
    n13190, n13191, n13192, n13193, n13194, n13195,
    n13196, n13197, n13198, n13199, n13200, n13201,
    n13202, n13203, n13204, n13205, n13206, n13207,
    n13208, n13209, n13210, n13211, n13212, n13213,
    n13214, n13215, n13216, n13217, n13218, n13219,
    n13220, n13221, n13222, n13223, n13224, n13225,
    n13226, n13227, n13228, n13229, n13230, n13231,
    n13232, n13233, n13234, n13235, n13236, n13237,
    n13238, n13239, n13240, n13241, n13242, n13243,
    n13244, n13245, n13246, n13247, n13248, n13249,
    n13250, n13251, n13252, n13253, n13254, n13255,
    n13256, n13257, n13258, n13259, n13260, n13261,
    n13262, n13263, n13264, n13265, n13266, n13267,
    n13268, n13269, n13270, n13271, n13272, n13273,
    n13274, n13275, n13276, n13277, n13278, n13279,
    n13280, n13281, n13282, n13283, n13284, n13285,
    n13286, n13287, n13288, n13289, n13290, n13291,
    n13292, n13293, n13294, n13295, n13296, n13297,
    n13298, n13299, n13300, n13301, n13302, n13303,
    n13304, n13305, n13306, n13307, n13308, n13309,
    n13310, n13311, n13312, n13313, n13314, n13315,
    n13316, n13317, n13318, n13319, n13320, n13321,
    n13322, n13323, n13324, n13325, n13326, n13327,
    n13328, n13329, n13330, n13331, n13332, n13333,
    n13334, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13342, n13343, n13344, n13345,
    n13346, n13347, n13348, n13349, n13350, n13351,
    n13352, n13353, n13354, n13355, n13356, n13357,
    n13358, n13359, n13360, n13361, n13362, n13363,
    n13364, n13365, n13366, n13367, n13368, n13369,
    n13370, n13371, n13372, n13373, n13374, n13375,
    n13376, n13377, n13378, n13379, n13380, n13381,
    n13382, n13383, n13384, n13385, n13386, n13387,
    n13388, n13389, n13390, n13391, n13392, n13393,
    n13394, n13395, n13396, n13397, n13398, n13399,
    n13400, n13401, n13402, n13403, n13404, n13405,
    n13406, n13407, n13408, n13409, n13410, n13411,
    n13412, n13413, n13414, n13415, n13416, n13417,
    n13418, n13419, n13420, n13421, n13422, n13423,
    n13424, n13425, n13426, n13427, n13428, n13429,
    n13430, n13431, n13432, n13433, n13434, n13435,
    n13436, n13437, n13438, n13439, n13440, n13441,
    n13442, n13443, n13444, n13445, n13446, n13447,
    n13448, n13449, n13450, n13451, n13452, n13453,
    n13454, n13455, n13456, n13457, n13458, n13459,
    n13460, n13461, n13462, n13463, n13464, n13465,
    n13466, n13467, n13468, n13469, n13470, n13471,
    n13472, n13473, n13474, n13475, n13476, n13477,
    n13478, n13479, n13480, n13481, n13482, n13483,
    n13484, n13485, n13486, n13487, n13488, n13489,
    n13490, n13491, n13492, n13493, n13494, n13495,
    n13496, n13497, n13498, n13499, n13500, n13501,
    n13502, n13503, n13504, n13505, n13506, n13507,
    n13508, n13509, n13510, n13511, n13512, n13513,
    n13514, n13515, n13516, n13517, n13518, n13519,
    n13520, n13521, n13522, n13523, n13524, n13525,
    n13526, n13527, n13528, n13529, n13530, n13531,
    n13532, n13533, n13534, n13535, n13536, n13537,
    n13538, n13539, n13540, n13541, n13542, n13543,
    n13544, n13545, n13546, n13547, n13548, n13549,
    n13550, n13551, n13552, n13553, n13554, n13555,
    n13556, n13557, n13558, n13559, n13560, n13561,
    n13562, n13563, n13564, n13565, n13566, n13567,
    n13568, n13569, n13570, n13571, n13572, n13573,
    n13574, n13575, n13576, n13577, n13578, n13579,
    n13580, n13581, n13582, n13583, n13584, n13585,
    n13586, n13587, n13588, n13589, n13590, n13591,
    n13592, n13593, n13594, n13595, n13596, n13597,
    n13598, n13599, n13600, n13601, n13602, n13603,
    n13604, n13605, n13606, n13607, n13608, n13609,
    n13610, n13611, n13612, n13613, n13614, n13615,
    n13616, n13617, n13618, n13619, n13620, n13621,
    n13622, n13623, n13624, n13625, n13626, n13627,
    n13628, n13629, n13630, n13631, n13632, n13633,
    n13634, n13635, n13636, n13637, n13638, n13639,
    n13640, n13641, n13642, n13643, n13644, n13645,
    n13646, n13647, n13648, n13649, n13650, n13651,
    n13652, n13653, n13654, n13655, n13656, n13657,
    n13658, n13659, n13660, n13661, n13662, n13663,
    n13664, n13665, n13666, n13667, n13668, n13669,
    n13670, n13671, n13672, n13673, n13674, n13675,
    n13676, n13677, n13678, n13679, n13680, n13681,
    n13682, n13683, n13684, n13685, n13686, n13687,
    n13688, n13689, n13690, n13691, n13692, n13693,
    n13694, n13695, n13696, n13697, n13698, n13699,
    n13700, n13701, n13702, n13703, n13704, n13705,
    n13706, n13707, n13708, n13709, n13710, n13711,
    n13712, n13713, n13714, n13715, n13716, n13717,
    n13718, n13719, n13720, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729,
    n13730, n13731, n13732, n13733, n13734, n13735,
    n13736, n13737, n13738, n13739, n13740, n13741,
    n13742, n13743, n13744, n13745, n13746, n13747,
    n13748, n13749, n13750, n13751, n13752, n13753,
    n13754, n13755, n13756, n13757, n13758, n13759,
    n13760, n13761, n13762, n13763, n13764, n13765,
    n13766, n13767, n13768, n13769, n13770, n13771,
    n13772, n13773, n13774, n13775, n13776, n13777,
    n13778, n13779, n13780, n13781, n13782, n13783,
    n13784, n13785, n13786, n13787, n13788, n13789,
    n13790, n13791, n13792, n13793, n13794, n13795,
    n13796, n13797, n13798, n13799, n13800, n13801,
    n13802, n13803, n13804, n13805, n13806, n13807,
    n13808, n13809, n13810, n13811, n13812, n13813,
    n13814, n13815, n13816, n13817, n13818, n13819,
    n13820, n13821, n13822, n13823, n13824, n13825,
    n13826, n13827, n13828, n13829, n13830, n13831,
    n13832, n13833, n13834, n13835, n13836, n13837,
    n13838, n13839, n13840, n13841, n13842, n13843,
    n13844, n13845, n13846, n13847, n13848, n13849,
    n13850, n13851, n13852, n13853, n13854, n13855,
    n13856, n13857, n13858, n13859, n13860, n13861,
    n13862, n13863, n13864, n13865, n13866, n13867,
    n13868, n13869, n13870, n13871, n13872, n13873,
    n13874, n13875, n13876, n13877, n13878, n13879,
    n13880, n13881, n13882, n13883, n13884, n13885,
    n13886, n13887, n13888, n13889, n13890, n13891,
    n13892, n13893, n13894, n13895, n13896, n13897,
    n13898, n13899, n13900, n13901, n13902, n13903,
    n13904, n13905, n13906, n13907, n13908, n13909,
    n13910, n13911, n13912, n13913, n13914, n13915,
    n13916, n13917, n13918, n13919, n13920, n13921,
    n13922, n13923, n13924, n13925, n13926, n13927,
    n13928, n13929, n13930, n13931, n13932, n13933,
    n13934, n13935, n13936, n13937, n13938, n13939,
    n13940, n13941, n13942, n13943, n13944, n13945,
    n13946, n13947, n13948, n13949, n13950, n13951,
    n13952, n13953, n13954, n13955, n13956, n13957,
    n13958, n13959, n13960, n13961, n13962, n13963,
    n13964, n13965, n13966, n13967, n13968, n13969,
    n13970, n13971, n13972, n13973, n13974, n13975,
    n13976, n13977, n13978, n13979, n13980, n13981,
    n13982, n13983, n13984, n13985, n13986, n13987,
    n13988, n13989, n13990, n13991, n13992, n13993,
    n13994, n13995, n13996, n13997, n13998, n13999,
    n14000, n14001, n14002, n14003, n14004, n14005,
    n14006, n14007, n14008, n14009, n14010, n14011,
    n14012, n14013, n14014, n14015, n14016, n14017,
    n14018, n14019, n14020, n14021, n14022, n14023,
    n14024, n14025, n14026, n14027, n14028, n14029,
    n14030, n14031, n14032, n14033, n14034, n14035,
    n14036, n14037, n14038, n14039, n14040, n14041,
    n14042, n14043, n14044, n14045, n14046, n14047,
    n14048, n14049, n14050, n14051, n14052, n14053,
    n14054, n14055, n14056, n14057, n14058, n14059,
    n14060, n14061, n14062, n14063, n14064, n14065,
    n14066, n14067, n14068, n14069, n14070, n14071,
    n14072, n14073, n14074, n14075, n14076, n14077,
    n14078, n14079, n14080, n14081, n14082, n14083,
    n14084, n14085, n14086, n14087, n14088, n14089,
    n14090, n14091, n14092, n14093, n14094, n14095,
    n14096, n14097, n14098, n14099, n14100, n14101,
    n14102, n14103, n14104, n14105, n14106, n14107,
    n14108, n14109, n14110, n14111, n14112, n14113,
    n14114, n14115, n14116, n14117, n14118, n14119,
    n14120, n14121, n14122, n14123, n14124, n14125,
    n14126, n14127, n14128, n14129, n14130, n14131,
    n14132, n14133, n14134, n14135, n14136, n14137,
    n14138, n14139, n14140, n14141, n14142, n14143,
    n14144, n14145, n14146, n14147, n14148, n14149,
    n14150, n14151, n14152, n14153, n14154, n14155,
    n14156, n14157, n14158, n14159, n14160, n14161,
    n14162, n14163, n14164, n14165, n14166, n14167,
    n14168, n14169, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14178, n14179,
    n14180, n14181, n14182, n14183, n14184, n14185,
    n14186, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197,
    n14198, n14199, n14200, n14201, n14202, n14203,
    n14204, n14205, n14206, n14207, n14208, n14209,
    n14210, n14211, n14212, n14213, n14214, n14215,
    n14216, n14217, n14218, n14219, n14220, n14221,
    n14222, n14223, n14224, n14225, n14226, n14227,
    n14228, n14229, n14230, n14231, n14232, n14233,
    n14234, n14235, n14236, n14237, n14238, n14239,
    n14240, n14241, n14242, n14243, n14244, n14245,
    n14246, n14247, n14248, n14249, n14250, n14251,
    n14252, n14253, n14254, n14255, n14256, n14257,
    n14258, n14259, n14260, n14261, n14262, n14263,
    n14264, n14265, n14266, n14267, n14268, n14269,
    n14270, n14271, n14272, n14273, n14274, n14275,
    n14276, n14277, n14278, n14279, n14280, n14281,
    n14282, n14283, n14284, n14285, n14286, n14287,
    n14288, n14289, n14290, n14291, n14292, n14293,
    n14294, n14295, n14296, n14297, n14298, n14299,
    n14300, n14301, n14302, n14303, n14304, n14305,
    n14306, n14307, n14308, n14309, n14310, n14311,
    n14312, n14313, n14314, n14315, n14316, n14317,
    n14318, n14319, n14320, n14321, n14322, n14323,
    n14324, n14325, n14326, n14327, n14328, n14329,
    n14330, n14331, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14340, n14341,
    n14342, n14343, n14344, n14345, n14346, n14347,
    n14348, n14349, n14350, n14351, n14352, n14353,
    n14354, n14355, n14356, n14357, n14358, n14359,
    n14360, n14361, n14362, n14363, n14364, n14365,
    n14366, n14367, n14368, n14369, n14370, n14371,
    n14372, n14373, n14374, n14375, n14376, n14377,
    n14378, n14379, n14380, n14381, n14382, n14383,
    n14384, n14385, n14386, n14387, n14388, n14389,
    n14390, n14391, n14392, n14393, n14394, n14395,
    n14396, n14397, n14398, n14399, n14400, n14401,
    n14402, n14403, n14404, n14405, n14406, n14407,
    n14408, n14409, n14410, n14411, n14412, n14413,
    n14414, n14415, n14416, n14417, n14418, n14419,
    n14420, n14421, n14422, n14423, n14424, n14425,
    n14426, n14427, n14428, n14429, n14430, n14431,
    n14432, n14433, n14434, n14435, n14436, n14437,
    n14438, n14439, n14440, n14441, n14442, n14443,
    n14444, n14445, n14446, n14447, n14448, n14449,
    n14450, n14451, n14452, n14453, n14454, n14455,
    n14456, n14457, n14458, n14459, n14460, n14461,
    n14462, n14463, n14464, n14465, n14466, n14467,
    n14468, n14469, n14470, n14471, n14472, n14473,
    n14474, n14475, n14476, n14477, n14478, n14479,
    n14480, n14481, n14482, n14483, n14484, n14485,
    n14486, n14487, n14488, n14489, n14490, n14491,
    n14492, n14493, n14494, n14495, n14496, n14497,
    n14498, n14499, n14500, n14501, n14502, n14503,
    n14504, n14505, n14506, n14507, n14508, n14509,
    n14510, n14511, n14512, n14513, n14514, n14515,
    n14516, n14517, n14518, n14519, n14520, n14521,
    n14522, n14523, n14524, n14525, n14526, n14527,
    n14528, n14529, n14530, n14531, n14532, n14533,
    n14534, n14535, n14536, n14537, n14538, n14539,
    n14540, n14541, n14542, n14543, n14544, n14545,
    n14546, n14547, n14548, n14549, n14550, n14551,
    n14552, n14553, n14554, n14555, n14556, n14557,
    n14558, n14559, n14560, n14561, n14562, n14563,
    n14564, n14565, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14573, n14574, n14575,
    n14576, n14577, n14578, n14579, n14580, n14581,
    n14582, n14583, n14584, n14585, n14586, n14587,
    n14588, n14589, n14590, n14591, n14592, n14593,
    n14594, n14595, n14596, n14597, n14598, n14599,
    n14600, n14601, n14602, n14603, n14604, n14605,
    n14606, n14607, n14608, n14609, n14610, n14611,
    n14612, n14613, n14614, n14615, n14616, n14617,
    n14618, n14619, n14620, n14621, n14622, n14623,
    n14624, n14625, n14626, n14627, n14628, n14629,
    n14630, n14631, n14632, n14633, n14634, n14635,
    n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647,
    n14648, n14649, n14650, n14651, n14652, n14653,
    n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665,
    n14666, n14667, n14668, n14669, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683,
    n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701,
    n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719,
    n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731,
    n14732, n14733, n14734, n14735, n14736, n14737,
    n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749,
    n14750, n14751, n14752, n14753, n14754, n14755,
    n14756, n14757, n14758, n14759, n14760, n14761,
    n14762, n14763, n14764, n14765, n14766, n14767,
    n14768, n14769, n14770, n14771, n14772, n14773,
    n14774, n14775, n14776, n14777, n14778, n14779,
    n14780, n14781, n14782, n14783, n14784, n14785,
    n14786, n14787, n14788, n14789, n14790, n14791,
    n14792, n14793, n14794, n14795, n14796, n14797,
    n14798, n14799, n14800, n14801, n14802, n14803,
    n14804, n14805, n14806, n14807, n14808, n14809,
    n14810, n14811, n14812, n14813, n14814, n14815,
    n14816, n14817, n14818, n14819, n14820, n14821,
    n14822, n14823, n14824, n14825, n14826, n14827,
    n14828, n14829, n14830, n14831, n14832, n14833,
    n14834, n14835, n14836, n14837, n14838, n14839,
    n14840, n14841, n14842, n14843, n14844, n14845,
    n14846, n14847, n14848, n14849, n14850, n14851,
    n14852, n14853, n14854, n14855, n14856, n14857,
    n14858, n14859, n14860, n14861, n14862, n14863,
    n14864, n14865, n14866, n14867, n14868, n14869,
    n14870, n14871, n14872, n14873, n14874, n14875,
    n14876, n14877, n14878, n14879, n14880, n14881,
    n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14890, n14891, n14892, n14893,
    n14894, n14895, n14896, n14897, n14898, n14899,
    n14900, n14901, n14902, n14903, n14904, n14905,
    n14906, n14907, n14908, n14909, n14910, n14911,
    n14912, n14913, n14914, n14915, n14916, n14917,
    n14918, n14919, n14920, n14921, n14922, n14923,
    n14924, n14925, n14926, n14927, n14928, n14929,
    n14930, n14931, n14932, n14933, n14934, n14935,
    n14936, n14937, n14938, n14939, n14940, n14941,
    n14942, n14943, n14944, n14945, n14946, n14947,
    n14948, n14949, n14950, n14951, n14952, n14953,
    n14954, n14955, n14956, n14957, n14958, n14959,
    n14960, n14961, n14962, n14963, n14964, n14965,
    n14966, n14967, n14968, n14969, n14970, n14971,
    n14972, n14973, n14974, n14975, n14976, n14977,
    n14978, n14979, n14980, n14981, n14982, n14983,
    n14984, n14985, n14986, n14987, n14988, n14989,
    n14990, n14991, n14992, n14993, n14994, n14995,
    n14996, n14997, n14998, n14999, n15000, n15001,
    n15002, n15003, n15004, n15005, n15006, n15007,
    n15008, n15009, n15010, n15011, n15012, n15013,
    n15014, n15015, n15016, n15017, n15018, n15019,
    n15020, n15021, n15022, n15023, n15024, n15025,
    n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037,
    n15038, n15039, n15040, n15041, n15042, n15043,
    n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055,
    n15056, n15057, n15058, n15059, n15060, n15061,
    n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073,
    n15074, n15075, n15076, n15077, n15078, n15079,
    n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091,
    n15092, n15093, n15094, n15095, n15096, n15097,
    n15098, n15099, n15100, n15101, n15102, n15103,
    n15104, n15105, n15106, n15107, n15108, n15109,
    n15110, n15111, n15112, n15113, n15114, n15115,
    n15116, n15117, n15118, n15119, n15120, n15121,
    n15122, n15123, n15124, n15125, n15126, n15127,
    n15128, n15129, n15130, n15131, n15132, n15133,
    n15134, n15135, n15136, n15137, n15138, n15139,
    n15140, n15141, n15142, n15143, n15144, n15145,
    n15146, n15147, n15148, n15149, n15150, n15151,
    n15152, n15153, n15154, n15155, n15156, n15157,
    n15158, n15159, n15160, n15161, n15162, n15163,
    n15164, n15165, n15166, n15167, n15168, n15169,
    n15170, n15171, n15172, n15173, n15174, n15175,
    n15176, n15177, n15178, n15179, n15180, n15181,
    n15182, n15183, n15184, n15185, n15186, n15187,
    n15188, n15189, n15190, n15191, n15192, n15193,
    n15194, n15195, n15196, n15197, n15198, n15199,
    n15200, n15201, n15202, n15203, n15204, n15205,
    n15206, n15207, n15208, n15209, n15210, n15211,
    n15212, n15213, n15214, n15215, n15216, n15217,
    n15218, n15219, n15220, n15221, n15222, n15223,
    n15224, n15225, n15226, n15227, n15228, n15229,
    n15230, n15231, n15232, n15233, n15234, n15235,
    n15236, n15237, n15238, n15239, n15240, n15241,
    n15242, n15243, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253,
    n15254, n15255, n15256, n15257, n15258, n15259,
    n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271,
    n15272, n15273, n15274, n15275, n15276, n15277,
    n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289,
    n15290, n15291, n15292, n15293, n15294, n15295,
    n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307,
    n15308, n15309, n15310, n15311, n15312, n15313,
    n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325,
    n15326, n15327, n15328, n15329, n15330, n15331,
    n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343,
    n15344, n15345, n15346, n15347, n15348, n15349,
    n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15357, n15358, n15359, n15360, n15361,
    n15362, n15363, n15364, n15365, n15366, n15367,
    n15368, n15369, n15370, n15371, n15372, n15373,
    n15374, n15375, n15376, n15377, n15378, n15379,
    n15380, n15381, n15382, n15383, n15384, n15385,
    n15386, n15387, n15388, n15389, n15390, n15391,
    n15392, n15393, n15394, n15395, n15396, n15397,
    n15398, n15399, n15400, n15401, n15402, n15403,
    n15404, n15405, n15406, n15407, n15408, n15409,
    n15410, n15411, n15412, n15413, n15414, n15415,
    n15416, n15417, n15418, n15419, n15420, n15421,
    n15422, n15423, n15424, n15425, n15426, n15427,
    n15428, n15429, n15430, n15431, n15432, n15433,
    n15434, n15435, n15436, n15437, n15438, n15439,
    n15440, n15441, n15442, n15443, n15444, n15445,
    n15446, n15447, n15448, n15449, n15450, n15451,
    n15452, n15453, n15454, n15455, n15456, n15457,
    n15458, n15459, n15460, n15461, n15462, n15463,
    n15464, n15465, n15466, n15467, n15468, n15469,
    n15470, n15471, n15472, n15473, n15474, n15475,
    n15476, n15477, n15478, n15479, n15480, n15481,
    n15482, n15483, n15484, n15485, n15486, n15487,
    n15488, n15489, n15490, n15491, n15492, n15493,
    n15494, n15495, n15496, n15497, n15498, n15499,
    n15500, n15501, n15502, n15503, n15504, n15505,
    n15506, n15507, n15508, n15509, n15510, n15511,
    n15512, n15513, n15514, n15515, n15516, n15517,
    n15518, n15519, n15520, n15521, n15522, n15523,
    n15524, n15525, n15526, n15527, n15528, n15529,
    n15530, n15531, n15532, n15533, n15534, n15535,
    n15536, n15537, n15538, n15539, n15540, n15541,
    n15542, n15543, n15544, n15545, n15546, n15547,
    n15548, n15549, n15550, n15551, n15552, n15553,
    n15554, n15555, n15556, n15557, n15558, n15559,
    n15560, n15561, n15562, n15563, n15564, n15565,
    n15566, n15567, n15568, n15569, n15570, n15571,
    n15572, n15573, n15574, n15575, n15576, n15577,
    n15578, n15579, n15580, n15581, n15582, n15583,
    n15584, n15585, n15586, n15587, n15588, n15589,
    n15590, n15591, n15592, n15593, n15594, n15595,
    n15596, n15597, n15598, n15599, n15600, n15601,
    n15602, n15603, n15604, n15605, n15606, n15607,
    n15608, n15609, n15610, n15611, n15612, n15613,
    n15614, n15615, n15616, n15617, n15618, n15619,
    n15620, n15621, n15622, n15623, n15624, n15625,
    n15626, n15627, n15628, n15629, n15630, n15631,
    n15632, n15633, n15634, n15635, n15636, n15637,
    n15638, n15639, n15640, n15641, n15642, n15643,
    n15644, n15645, n15646, n15647, n15648, n15649,
    n15650, n15651, n15652, n15653, n15654, n15655,
    n15656, n15657, n15658, n15659, n15660, n15661,
    n15662, n15663, n15664, n15665, n15666, n15667,
    n15668, n15669, n15670, n15671, n15672, n15673,
    n15674, n15675, n15676, n15677, n15678, n15679,
    n15680, n15681, n15682, n15683, n15684, n15685,
    n15686, n15687, n15688, n15689, n15690, n15691,
    n15692, n15693, n15694, n15695, n15696, n15697,
    n15698, n15699, n15700, n15701, n15702, n15703,
    n15704, n15705, n15706, n15707, n15708, n15709,
    n15710, n15711, n15712, n15713, n15714, n15715,
    n15716, n15717, n15718, n15719, n15720, n15721,
    n15722, n15723, n15724, n15725, n15726, n15727,
    n15728, n15729, n15730, n15731, n15732, n15733,
    n15734, n15735, n15736, n15737, n15738, n15739,
    n15740, n15741, n15742, n15743, n15744, n15745,
    n15746, n15747, n15748, n15749, n15750, n15751,
    n15752, n15753, n15754, n15755, n15756, n15757,
    n15758, n15759, n15760, n15761, n15762, n15763,
    n15764, n15765, n15766, n15767, n15768, n15769,
    n15770, n15771, n15772, n15773, n15774, n15775,
    n15776, n15777, n15778, n15779, n15780, n15781,
    n15782, n15783, n15784, n15785, n15786, n15787,
    n15788, n15789, n15790, n15791, n15792, n15793,
    n15794, n15795, n15796, n15797, n15798, n15799,
    n15800, n15801, n15802, n15803, n15804, n15805,
    n15806, n15807, n15808, n15809, n15810, n15811,
    n15812, n15813, n15814, n15815, n15816, n15817,
    n15818, n15819, n15820, n15821, n15822, n15823,
    n15824, n15825, n15826, n15827, n15828, n15829,
    n15830, n15831, n15832, n15833, n15834, n15835,
    n15836, n15837, n15838, n15839, n15840, n15841,
    n15842, n15843, n15844, n15845, n15846, n15847,
    n15848, n15849, n15850, n15851, n15852, n15853,
    n15854, n15855, n15856, n15857, n15858, n15859,
    n15860, n15861, n15862, n15863, n15864, n15865,
    n15866, n15867, n15868, n15869, n15870, n15871,
    n15872, n15873, n15874, n15875, n15876, n15877,
    n15878, n15879, n15880, n15881, n15882, n15883,
    n15884, n15885, n15886, n15887, n15888, n15889,
    n15890, n15891, n15892, n15893, n15894, n15895,
    n15896, n15897, n15898, n15899, n15900, n15901,
    n15902, n15903, n15904, n15905, n15906, n15907,
    n15908, n15909, n15910, n15911, n15912, n15913,
    n15914, n15915, n15916, n15917, n15918, n15919,
    n15920, n15921, n15922, n15923, n15924, n15925,
    n15926, n15927, n15928, n15929, n15930, n15931,
    n15932, n15933, n15934, n15935, n15936, n15937,
    n15938, n15939, n15940, n15941, n15942, n15943,
    n15944, n15945, n15946, n15947, n15948, n15949,
    n15950, n15951, n15952, n15953, n15954, n15955,
    n15956, n15957, n15958, n15959, n15960, n15961,
    n15962, n15963, n15964, n15965, n15966, n15967,
    n15968, n15969, n15970, n15971, n15972, n15973,
    n15974, n15975, n15976, n15977, n15978, n15979,
    n15980, n15981, n15982, n15983, n15984, n15985,
    n15986, n15987, n15988, n15989, n15990, n15991,
    n15992, n15993, n15994, n15995, n15996, n15997,
    n15998, n15999, n16000, n16001, n16002, n16003,
    n16004, n16005, n16006, n16007, n16008, n16009,
    n16010, n16011, n16012, n16013, n16014, n16015,
    n16016, n16017, n16018, n16019, n16020, n16021,
    n16022, n16023, n16024, n16025, n16026, n16027,
    n16028, n16029, n16030, n16031, n16032, n16033,
    n16034, n16035, n16036, n16037, n16038, n16039,
    n16040, n16041, n16042, n16043, n16044, n16045,
    n16046, n16047, n16048, n16049, n16050, n16051,
    n16052, n16053, n16054, n16055, n16056, n16057,
    n16058, n16059, n16060, n16061, n16062, n16063,
    n16064, n16065, n16066, n16067, n16068, n16069,
    n16070, n16071, n16072, n16073, n16074, n16075,
    n16076, n16077, n16078, n16079, n16080, n16081,
    n16082, n16083, n16084, n16085, n16086, n16087,
    n16088, n16089, n16090, n16091, n16092, n16093,
    n16094, n16095, n16096, n16097, n16098, n16099,
    n16100, n16101, n16102, n16103, n16104, n16105,
    n16106, n16107, n16108, n16109, n16110, n16111,
    n16112, n16113, n16114, n16115, n16116, n16117,
    n16118, n16119, n16120, n16121, n16122, n16123,
    n16124, n16125, n16126, n16127, n16128, n16129,
    n16130, n16131, n16132, n16133, n16134, n16135,
    n16136, n16137, n16138, n16139, n16140, n16141,
    n16142, n16143, n16144, n16145, n16146, n16147,
    n16148, n16149, n16150, n16151, n16152, n16153,
    n16154, n16155, n16156, n16157, n16158, n16159,
    n16160, n16161, n16162, n16163, n16164, n16165,
    n16166, n16167, n16168, n16169, n16170, n16171,
    n16172, n16173, n16174, n16175, n16176, n16177,
    n16178, n16179, n16180, n16181, n16182, n16183,
    n16184, n16185, n16186, n16187, n16188, n16189,
    n16190, n16191, n16192, n16193, n16194, n16195,
    n16196, n16197, n16198, n16199, n16200, n16201,
    n16202, n16203, n16204, n16205, n16206, n16207,
    n16208, n16209, n16210, n16211, n16212, n16213,
    n16214, n16215, n16216, n16217, n16218, n16219,
    n16220, n16221, n16222, n16223, n16224, n16225,
    n16226, n16227, n16228, n16229, n16230, n16231,
    n16232, n16233, n16234, n16235, n16236, n16237,
    n16238, n16239, n16240, n16241, n16242, n16243,
    n16244, n16245, n16246, n16247, n16248, n16249,
    n16250, n16251, n16252, n16253, n16254, n16255,
    n16256, n16257, n16258, n16259, n16260, n16261,
    n16262, n16263, n16264, n16265, n16266, n16267,
    n16268, n16269, n16270, n16271, n16272, n16273,
    n16274, n16275, n16276, n16277, n16278, n16279,
    n16280, n16281, n16282, n16283, n16284, n16285,
    n16286, n16287, n16288, n16289, n16290, n16291,
    n16292, n16293, n16294, n16295, n16296, n16297,
    n16298, n16299, n16300, n16301, n16302, n16303,
    n16304, n16305, n16306, n16307, n16308, n16309,
    n16310, n16311, n16312, n16313, n16314, n16315,
    n16316, n16317, n16318, n16319, n16320, n16321,
    n16322, n16323, n16324, n16325, n16326, n16327,
    n16328, n16329, n16330, n16331, n16332, n16333,
    n16334, n16335, n16336, n16337, n16338, n16339,
    n16340, n16341, n16342, n16343, n16344, n16345,
    n16346, n16347, n16348, n16349, n16350, n16351,
    n16352, n16353, n16354, n16355, n16356, n16357,
    n16358, n16359, n16360, n16361, n16362, n16363,
    n16364, n16365, n16366, n16367, n16368, n16369,
    n16370, n16371, n16372, n16373, n16374, n16375,
    n16376, n16377, n16378, n16379, n16380, n16381,
    n16382, n16383, n16384, n16385, n16386, n16387,
    n16388, n16389, n16390, n16391, n16392, n16393,
    n16394, n16395, n16396, n16397, n16398, n16399,
    n16400, n16401, n16402, n16403, n16404, n16405,
    n16406, n16407, n16408, n16409, n16410, n16411,
    n16412, n16413, n16414, n16415, n16416, n16417,
    n16418, n16419, n16420, n16421, n16422, n16423,
    n16424, n16425, n16426, n16427, n16428, n16429,
    n16430, n16431, n16432, n16433, n16434, n16435,
    n16436, n16437, n16438, n16439, n16440, n16441,
    n16442, n16443, n16444, n16445, n16446, n16447,
    n16448, n16449, n16450, n16451, n16452, n16453,
    n16454, n16455, n16456, n16457, n16458, n16459,
    n16460, n16461, n16462, n16463, n16464, n16465,
    n16466, n16467, n16468, n16469, n16470, n16471,
    n16472, n16473, n16474, n16475, n16476, n16477,
    n16478, n16479, n16480, n16481, n16482, n16483,
    n16484, n16485, n16486, n16487, n16488, n16489,
    n16490, n16491, n16492, n16493, n16494, n16495,
    n16496, n16497, n16498, n16499, n16500, n16501,
    n16502, n16503, n16504, n16505, n16506, n16507,
    n16508, n16509, n16510, n16511, n16512, n16513,
    n16514, n16515, n16516, n16517, n16518, n16519,
    n16520, n16521, n16522, n16523, n16524, n16525,
    n16526, n16527, n16528, n16529, n16530, n16531,
    n16532, n16533, n16534, n16535, n16536, n16537,
    n16538, n16539, n16540, n16541, n16542, n16543,
    n16544, n16545, n16546, n16547, n16548, n16549,
    n16550, n16551, n16552, n16553, n16554, n16555,
    n16556, n16557, n16558, n16559, n16560, n16561,
    n16562, n16563, n16564, n16565, n16566, n16567,
    n16568, n16569, n16570, n16571, n16572, n16573,
    n16574, n16575, n16576, n16577, n16578, n16579,
    n16580, n16581, n16582, n16583, n16584, n16585,
    n16586, n16587, n16588, n16589, n16590, n16591,
    n16592, n16593, n16594, n16595, n16596, n16597,
    n16598, n16599, n16600, n16601, n16602, n16603,
    n16604, n16605, n16606, n16607, n16608, n16609,
    n16610, n16611, n16612, n16613, n16614, n16615,
    n16616, n16617, n16618, n16619, n16620, n16621,
    n16622, n16623, n16624, n16625, n16626, n16627,
    n16628, n16629, n16630, n16631, n16632, n16633,
    n16634, n16635, n16636, n16637, n16638, n16639,
    n16640, n16641, n16642, n16643, n16644, n16645,
    n16646, n16647, n16648, n16649, n16650, n16651,
    n16652, n16653, n16654, n16655, n16656, n16657,
    n16658, n16659, n16660, n16661, n16662, n16663,
    n16664, n16665, n16666, n16667, n16668, n16669,
    n16670, n16671, n16672, n16673, n16674, n16675,
    n16676, n16677, n16678, n16679, n16680, n16681,
    n16682, n16683, n16684, n16685, n16686, n16687,
    n16688, n16689, n16690, n16691, n16692, n16693,
    n16694, n16695, n16696, n16697, n16698, n16699,
    n16700, n16701, n16702, n16703, n16704, n16705,
    n16706, n16707, n16708, n16709, n16710, n16711,
    n16712, n16713, n16714, n16715, n16716, n16717,
    n16718, n16719, n16720, n16721, n16722, n16723,
    n16724, n16725, n16726, n16727, n16728, n16729,
    n16730, n16731, n16732, n16733, n16734, n16735,
    n16736, n16737, n16738, n16739, n16740, n16741,
    n16742, n16743, n16744, n16745, n16746, n16747,
    n16748, n16749, n16750, n16751, n16752, n16753,
    n16754, n16755, n16756, n16757, n16758, n16759,
    n16760, n16761, n16762, n16763, n16764, n16765,
    n16766, n16767, n16768, n16769, n16770, n16771,
    n16772, n16773, n16774, n16775, n16776, n16777,
    n16778, n16779, n16780, n16781, n16782, n16783,
    n16784, n16785, n16786, n16787, n16788, n16789,
    n16790, n16791, n16792, n16793, n16794, n16795,
    n16796, n16797, n16798, n16799, n16800, n16801,
    n16802, n16803, n16804, n16805, n16806, n16807,
    n16808, n16809, n16810, n16811, n16812, n16813,
    n16814, n16815, n16816, n16817, n16818, n16819,
    n16820, n16821, n16822, n16823, n16824, n16825,
    n16826, n16827, n16828, n16829, n16830, n16831,
    n16832, n16833, n16834, n16835, n16836, n16837,
    n16838, n16839, n16840, n16841, n16842, n16843,
    n16844, n16845, n16846, n16847, n16848, n16849,
    n16850, n16851, n16852, n16853, n16854, n16855,
    n16856, n16857, n16858, n16859, n16860, n16861,
    n16862, n16863, n16864, n16865, n16866, n16867,
    n16868, n16869, n16870, n16871, n16872, n16873,
    n16874, n16875, n16876, n16877, n16878, n16879,
    n16880, n16881, n16882, n16883, n16884, n16885,
    n16886, n16887, n16888, n16889, n16890, n16891,
    n16892, n16893, n16894, n16895, n16896, n16897,
    n16898, n16899, n16900, n16901, n16902, n16903,
    n16904, n16905, n16906, n16907, n16908, n16909,
    n16910, n16911, n16912, n16913, n16914, n16915,
    n16916, n16917, n16918, n16919, n16920, n16921,
    n16922, n16923, n16924, n16925, n16926, n16927,
    n16928, n16929, n16930, n16931, n16932, n16933,
    n16934, n16935, n16936, n16937, n16938, n16939,
    n16940, n16941, n16942, n16943, n16944, n16945,
    n16946, n16947, n16948, n16949, n16950, n16951,
    n16952, n16953, n16954, n16955, n16956, n16957,
    n16958, n16959, n16960, n16961, n16962, n16963,
    n16964, n16965, n16966, n16967, n16968, n16969,
    n16970, n16971, n16972, n16973, n16974, n16975,
    n16976, n16977, n16978, n16979, n16980, n16981,
    n16982, n16983, n16984, n16985, n16986, n16987,
    n16988, n16989, n16990, n16991, n16992, n16993,
    n16994, n16995, n16996, n16997, n16998, n16999,
    n17000, n17001, n17002, n17003, n17004, n17005,
    n17006, n17007, n17008, n17009, n17010, n17011,
    n17012, n17013, n17014, n17015, n17016, n17017,
    n17018, n17019, n17020, n17021, n17022, n17023,
    n17024, n17025, n17026, n17027, n17028, n17029,
    n17030, n17031, n17032, n17033, n17034, n17035,
    n17036, n17037, n17038, n17039, n17040, n17041,
    n17042, n17043, n17044, n17045, n17046, n17047,
    n17048, n17049, n17050, n17051, n17052, n17053,
    n17054, n17055, n17056, n17057, n17058, n17059,
    n17060, n17061, n17062, n17063, n17064, n17065,
    n17066, n17067, n17068, n17069, n17070, n17071,
    n17072, n17073, n17074, n17075, n17076, n17077,
    n17078, n17079, n17080, n17081, n17082, n17083,
    n17084, n17085, n17086, n17087, n17088, n17089,
    n17090, n17091, n17092, n17093, n17094, n17095,
    n17096, n17097, n17098, n17099, n17100, n17101,
    n17102, n17103, n17104, n17105, n17106, n17107,
    n17108, n17109, n17110, n17111, n17112, n17113,
    n17114, n17115, n17116, n17117, n17118, n17119,
    n17120, n17121, n17122, n17123, n17124, n17125,
    n17126, n17127, n17128, n17129, n17130, n17131,
    n17132, n17133, n17134, n17135, n17136, n17137,
    n17138, n17139, n17140, n17141, n17142, n17143,
    n17144, n17145, n17146, n17147, n17148, n17149,
    n17150, n17151, n17152, n17153, n17154, n17155,
    n17156, n17157, n17158, n17159, n17160, n17161,
    n17162, n17163, n17164, n17165, n17166, n17167,
    n17168, n17169, n17170, n17171, n17172, n17173,
    n17174, n17175, n17176, n17177, n17178, n17179,
    n17180, n17181, n17182, n17183, n17184, n17185,
    n17186, n17187, n17188, n17189, n17190, n17191,
    n17192, n17193, n17194, n17195, n17196, n17197,
    n17198, n17199, n17200, n17201, n17202, n17203,
    n17204, n17205, n17206, n17207, n17208, n17209,
    n17210, n17211, n17212, n17213, n17214, n17215,
    n17216, n17217, n17218, n17219, n17220, n17221,
    n17222, n17223, n17224, n17225, n17226, n17227,
    n17228, n17229, n17230, n17231, n17232, n17233,
    n17234, n17235, n17236, n17237, n17238, n17239,
    n17240, n17241, n17242, n17243, n17244, n17245,
    n17246, n17247, n17248, n17249, n17250, n17251,
    n17252, n17253, n17254, n17255, n17256, n17257,
    n17258, n17259, n17260, n17261, n17262, n17263,
    n17264, n17265, n17266, n17267, n17268, n17269,
    n17270, n17271, n17272, n17273, n17274, n17275,
    n17276, n17277, n17278, n17279, n17280, n17281,
    n17282, n17283, n17284, n17285, n17286, n17287,
    n17288, n17289, n17290, n17291, n17292, n17293,
    n17294, n17295, n17296, n17297, n17298, n17299,
    n17300, n17301, n17302, n17303, n17304, n17305,
    n17306, n17307, n17308, n17309, n17310, n17311,
    n17312, n17313, n17314, n17315, n17316, n17317,
    n17318, n17319, n17320, n17321, n17322, n17323,
    n17324, n17325, n17326, n17327, n17328, n17329,
    n17330, n17331, n17332, n17333, n17334, n17335,
    n17336, n17337, n17338, n17339, n17340, n17341,
    n17342, n17343, n17344, n17345, n17346, n17347,
    n17348, n17349, n17350, n17351, n17352, n17353,
    n17354, n17355, n17356, n17357, n17358, n17359,
    n17360, n17361, n17362, n17363, n17364, n17365,
    n17366, n17367, n17368, n17369, n17370, n17371,
    n17372, n17373, n17374, n17375, n17376, n17377,
    n17378, n17379, n17380, n17381, n17382, n17383,
    n17384, n17385, n17386, n17387, n17388, n17389,
    n17390, n17391, n17392, n17393, n17394, n17395,
    n17396, n17397, n17398, n17399, n17400, n17401,
    n17402, n17403, n17404, n17405, n17406, n17407,
    n17408, n17409, n17410, n17411, n17412, n17413,
    n17414, n17415, n17416, n17417, n17418, n17419,
    n17420, n17421, n17422, n17423, n17424, n17425,
    n17426, n17427, n17428, n17429, n17430, n17431,
    n17432, n17433, n17434, n17435, n17436, n17437,
    n17438, n17439, n17440, n17441, n17442, n17443,
    n17444, n17445, n17446, n17447, n17448, n17449,
    n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461,
    n17462, n17463, n17464, n17465, n17466, n17467,
    n17468, n17469, n17470, n17471, n17472, n17473,
    n17474, n17475, n17476, n17477, n17478, n17479,
    n17480, n17481, n17482, n17483, n17484, n17485,
    n17486, n17487, n17488, n17489, n17490, n17491,
    n17492, n17493, n17494, n17495, n17496, n17497,
    n17498, n17499, n17500, n17501, n17502, n17503,
    n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515,
    n17516, n17517, n17518, n17519, n17520, n17521,
    n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533,
    n17534, n17535, n17536, n17537, n17538, n17539,
    n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551,
    n17552, n17553, n17554, n17555, n17556, n17557,
    n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569,
    n17570, n17571, n17572, n17573, n17574, n17575,
    n17576, n17577, n17578, n17579, n17580, n17581,
    n17582, n17583, n17584, n17585, n17586, n17587,
    n17588, n17589, n17590, n17591, n17592, n17593,
    n17594, n17595, n17596, n17597, n17598, n17599,
    n17600, n17601, n17602, n17603, n17604, n17605,
    n17606, n17607, n17608, n17609, n17610, n17611,
    n17612, n17613, n17614, n17615, n17616, n17617,
    n17618, n17619, n17620, n17621, n17622, n17623,
    n17624, n17625, n17626, n17627, n17628, n17629,
    n17630, n17631, n17632, n17633, n17634, n17635,
    n17636, n17637, n17638, n17639, n17640, n17641,
    n17642, n17643, n17644, n17645, n17646, n17647,
    n17648, n17649, n17650, n17651, n17652, n17653,
    n17654, n17655, n17656, n17657, n17658, n17659,
    n17660, n17661, n17662, n17663, n17664, n17665,
    n17666, n17667, n17668, n17669, n17670, n17671,
    n17672, n17673, n17674, n17675, n17676, n17677,
    n17678, n17679, n17680, n17681, n17682, n17683,
    n17684, n17685, n17686, n17687, n17688, n17689,
    n17690, n17691, n17692, n17693, n17694, n17695,
    n17696, n17697, n17698, n17699, n17700, n17701,
    n17702, n17703, n17704, n17705, n17706, n17707,
    n17708, n17709, n17710, n17711, n17712, n17713,
    n17714, n17715, n17716, n17717, n17718, n17719,
    n17720, n17721, n17722, n17723, n17724, n17725,
    n17726, n17727, n17728, n17729, n17730, n17731,
    n17732, n17733, n17734, n17735, n17736, n17737,
    n17738, n17739, n17740, n17741, n17742, n17743,
    n17744, n17745, n17746, n17747, n17748, n17749,
    n17750, n17751, n17752, n17753, n17754, n17755,
    n17756, n17757, n17758, n17759, n17760, n17761,
    n17762, n17763, n17764, n17765, n17766, n17767,
    n17768, n17769, n17770, n17771, n17772, n17773,
    n17774, n17775, n17776, n17777, n17778, n17779,
    n17780, n17781, n17782, n17783, n17784, n17785,
    n17786, n17787, n17788, n17789, n17790, n17791,
    n17792, n17793, n17794, n17795, n17796, n17797,
    n17798, n17799, n17800, n17801, n17802, n17803,
    n17804, n17805, n17806, n17807, n17808, n17809,
    n17810, n17811, n17812, n17813, n17814, n17815,
    n17816, n17817, n17818, n17819, n17820, n17821,
    n17822, n17823, n17824, n17825, n17826, n17827,
    n17828, n17829, n17830, n17831, n17832, n17833,
    n17834, n17835, n17836, n17837, n17838, n17839,
    n17840, n17841, n17842, n17843, n17844, n17845,
    n17846, n17847, n17848, n17849, n17850, n17851,
    n17852, n17853, n17854, n17855, n17856, n17857,
    n17858, n17859, n17860, n17861, n17862, n17863,
    n17864, n17865, n17866, n17867, n17868, n17869,
    n17870, n17871, n17872, n17873, n17874, n17875,
    n17876, n17877, n17878, n17879, n17880, n17881,
    n17882, n17883, n17884, n17885, n17886, n17887,
    n17888, n17889, n17890, n17891, n17892, n17893,
    n17894, n17895, n17896, n17897, n17898, n17899,
    n17900, n17901, n17902, n17903, n17904, n17905,
    n17906, n17907, n17908, n17909, n17910, n17911,
    n17912, n17913, n17914, n17915, n17916, n17917,
    n17918, n17919, n17920, n17921, n17922, n17923,
    n17924, n17925, n17926, n17927, n17928, n17929,
    n17930, n17931, n17932, n17933, n17934, n17935,
    n17936, n17937, n17938, n17939, n17940, n17941,
    n17942, n17943, n17944, n17945, n17946, n17947,
    n17948, n17949, n17950, n17951, n17952, n17953,
    n17954, n17955, n17956, n17957, n17958, n17959,
    n17960, n17961, n17962, n17963, n17964, n17965,
    n17966, n17967, n17968, n17969, n17970, n17971,
    n17972, n17973, n17974, n17975, n17976, n17977,
    n17978, n17979, n17980, n17981, n17982, n17983,
    n17984, n17985, n17986, n17987, n17988, n17989,
    n17990, n17991, n17992, n17993, n17994, n17995,
    n17996, n17997, n17998, n17999, n18000, n18001,
    n18002, n18003, n18004, n18005, n18006, n18007,
    n18008, n18009, n18010, n18011, n18012, n18013,
    n18014, n18015, n18016, n18017, n18018, n18019,
    n18020, n18021, n18022, n18023, n18024, n18025,
    n18026, n18027, n18028, n18029, n18030, n18031,
    n18032, n18033, n18034, n18035, n18036, n18037,
    n18038, n18039, n18040, n18041, n18042, n18043,
    n18044, n18045, n18046, n18047, n18048, n18049,
    n18050, n18051, n18052, n18053, n18054, n18055,
    n18056, n18057, n18058, n18059, n18060, n18061,
    n18062, n18063, n18064, n18065, n18066, n18067,
    n18068, n18069, n18070, n18071, n18072, n18073,
    n18074, n18075, n18076, n18077, n18078, n18079,
    n18080, n18081, n18082, n18083, n18084, n18085,
    n18086, n18087, n18088, n18089, n18090, n18091,
    n18092, n18093, n18094, n18095, n18096, n18097,
    n18098, n18099, n18100, n18101, n18102, n18103,
    n18104, n18105, n18106, n18107, n18108, n18109,
    n18110, n18111, n18112, n18113, n18114, n18115,
    n18116, n18117, n18118, n18119, n18120, n18121,
    n18122, n18123, n18124, n18125, n18126, n18127,
    n18128, n18129, n18130, n18131, n18132, n18133,
    n18134, n18135, n18136, n18137, n18138, n18139,
    n18140, n18141, n18142, n18143, n18144, n18145,
    n18146, n18147, n18148, n18149, n18150, n18151,
    n18152, n18153, n18154, n18155, n18156, n18157,
    n18158, n18159, n18160, n18161, n18162, n18163,
    n18164, n18165, n18166, n18167, n18168, n18169,
    n18170, n18171, n18172, n18173, n18174, n18175,
    n18176, n18177, n18178, n18179, n18180, n18181,
    n18182, n18183, n18184, n18185, n18186, n18187,
    n18188, n18189, n18190, n18191, n18192, n18193,
    n18194, n18195, n18196, n18197, n18198, n18199,
    n18200, n18201, n18202, n18203, n18204, n18205,
    n18206, n18207, n18208, n18209, n18210, n18211,
    n18212, n18213, n18214, n18215, n18216, n18217,
    n18218, n18219, n18220, n18221, n18222, n18223,
    n18224, n18225, n18226, n18227, n18228, n18229,
    n18230, n18231, n18232, n18233, n18234, n18235,
    n18236, n18237, n18238, n18239, n18240, n18241,
    n18242, n18243, n18244, n18245, n18246, n18247,
    n18248, n18249, n18250, n18251, n18252, n18253,
    n18254, n18255, n18256, n18257, n18258, n18259,
    n18260, n18261, n18262, n18263, n18264, n18265,
    n18266, n18267, n18268, n18269, n18270, n18271,
    n18272, n18273, n18274, n18275, n18276, n18277,
    n18278, n18279, n18280, n18281, n18282, n18283,
    n18284, n18285, n18286, n18287, n18288, n18289,
    n18290, n18291, n18292, n18293, n18294, n18295,
    n18296, n18297, n18298, n18299, n18300, n18301,
    n18302, n18303, n18304, n18305, n18306, n18307,
    n18308, n18309, n18310, n18311, n18312, n18313,
    n18314, n18315, n18316, n18317, n18318, n18319,
    n18320, n18321, n18322, n18323, n18324, n18325,
    n18326, n18327, n18328, n18329, n18330, n18331,
    n18332, n18333, n18334, n18335, n18336, n18337,
    n18338, n18339, n18340, n18341, n18342, n18343,
    n18344, n18345, n18346, n18347, n18348, n18349,
    n18350, n18351, n18352, n18353, n18354, n18355,
    n18356, n18357, n18358, n18359, n18360, n18361,
    n18362, n18363, n18364, n18365, n18366, n18367,
    n18368, n18369, n18370, n18371, n18372, n18373,
    n18374, n18375, n18376, n18377, n18378, n18379,
    n18380, n18381, n18382, n18383, n18384, n18385,
    n18386, n18387, n18388, n18389, n18390, n18391,
    n18392, n18393, n18394, n18395, n18396, n18397,
    n18398, n18399, n18400, n18401, n18402, n18403,
    n18404, n18405, n18406, n18407, n18408, n18409,
    n18410, n18411, n18412, n18413, n18414, n18415,
    n18416, n18417, n18418, n18419, n18420, n18421,
    n18422, n18423, n18424, n18425, n18426, n18427,
    n18428, n18429, n18430, n18431, n18432, n18433,
    n18434, n18435, n18436, n18437, n18438, n18439,
    n18440, n18441, n18442, n18443, n18444, n18445,
    n18446, n18447, n18448, n18449, n18450, n18451,
    n18452, n18453, n18454, n18455, n18456, n18457,
    n18458, n18459, n18460, n18461, n18462, n18463,
    n18464, n18465, n18466, n18467, n18468, n18469,
    n18470, n18471, n18472, n18473, n18474, n18475,
    n18476, n18477, n18478, n18479, n18480, n18481,
    n18482, n18483, n18484, n18485, n18486, n18487,
    n18488, n18489, n18490, n18491, n18492, n18493,
    n18494, n18495, n18496, n18497, n18498, n18499,
    n18500, n18501, n18502, n18503, n18504, n18505,
    n18506, n18507, n18508, n18509, n18510, n18511,
    n18512, n18513, n18514, n18515, n18516, n18517,
    n18518, n18519, n18520, n18521, n18522, n18523,
    n18524, n18525, n18526, n18527, n18528, n18529,
    n18530, n18531, n18532, n18533, n18534, n18535,
    n18536, n18537, n18538, n18539, n18540, n18541,
    n18542, n18543, n18544, n18545, n18546, n18547,
    n18548, n18549, n18550, n18551, n18552, n18553,
    n18554, n18555, n18556, n18557, n18558, n18559,
    n18560, n18561, n18562, n18563, n18564, n18565,
    n18566, n18567, n18568, n18569, n18570, n18571,
    n18572, n18573, n18574, n18575, n18576, n18577,
    n18578, n18579, n18580, n18581, n18582, n18583,
    n18584, n18585, n18586, n18587, n18588, n18589,
    n18590, n18591, n18592, n18593, n18594, n18595,
    n18596, n18597, n18598, n18599, n18600, n18601,
    n18602, n18603, n18604, n18605, n18606, n18607,
    n18608, n18609, n18610, n18611, n18612, n18613,
    n18614, n18615, n18616, n18617, n18618, n18619,
    n18620, n18621, n18622, n18623, n18624, n18625,
    n18626, n18627, n18628, n18629, n18630, n18631,
    n18632, n18633, n18634, n18635, n18636, n18637,
    n18638, n18639, n18640, n18641, n18642, n18643,
    n18644, n18645, n18646, n18647, n18648, n18649,
    n18650, n18651, n18652, n18653, n18654, n18655,
    n18656, n18657, n18658, n18659, n18660, n18661,
    n18662, n18663, n18664, n18665, n18666, n18667,
    n18668, n18669, n18670, n18671, n18672, n18673,
    n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685,
    n18686, n18687, n18688, n18689, n18690, n18691,
    n18692, n18693, n18694, n18695, n18696, n18697,
    n18698, n18699, n18700, n18701, n18702, n18703,
    n18704, n18705, n18706, n18707, n18708, n18709,
    n18710, n18711, n18712, n18713, n18714, n18715,
    n18716, n18717, n18718, n18719, n18720, n18721,
    n18722, n18723, n18724, n18725, n18726, n18727,
    n18728, n18729, n18730, n18731, n18732, n18733,
    n18734, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18742, n18743, n18744, n18745,
    n18746, n18747, n18748, n18749, n18750, n18751,
    n18752, n18753, n18754, n18755, n18756, n18757,
    n18758, n18759, n18760, n18761, n18762, n18763,
    n18764, n18765, n18766, n18767, n18768, n18769,
    n18770, n18771, n18772, n18773, n18774, n18775,
    n18776, n18777, n18778, n18779, n18780, n18781,
    n18782, n18783, n18784, n18785, n18786, n18787,
    n18788, n18789, n18790, n18791, n18792, n18793,
    n18794, n18795, n18796, n18797, n18798, n18799,
    n18800, n18801, n18802, n18803, n18804, n18805,
    n18806, n18807, n18808, n18809, n18810, n18811,
    n18812, n18813, n18814, n18815, n18816, n18817,
    n18818, n18819, n18820, n18821, n18822, n18823,
    n18824, n18825, n18826, n18827, n18828, n18829,
    n18830, n18831, n18832, n18833, n18834, n18835,
    n18836, n18837, n18838, n18839, n18840, n18841,
    n18842, n18843, n18844, n18845, n18846, n18847,
    n18848, n18849, n18850, n18851, n18852, n18853,
    n18854, n18855, n18856, n18857, n18858, n18859,
    n18860, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18871,
    n18872, n18873, n18874, n18875, n18876, n18877,
    n18878, n18879, n18880, n18881, n18882, n18883,
    n18884, n18885, n18886, n18887, n18888, n18889,
    n18890, n18891, n18892, n18893, n18894, n18895,
    n18896, n18897, n18898, n18899, n18900, n18901,
    n18902, n18903, n18904, n18905, n18906, n18907,
    n18908, n18909, n18910, n18911, n18912, n18913,
    n18914, n18915, n18916, n18917, n18918, n18919,
    n18920, n18921, n18922, n18923, n18924, n18925,
    n18926, n18927, n18928, n18929, n18930, n18931,
    n18932, n18933, n18934, n18935, n18936, n18937,
    n18938, n18939, n18940, n18941, n18942, n18943,
    n18944, n18945, n18946, n18947, n18948, n18949,
    n18950, n18951, n18952, n18953, n18954, n18955,
    n18956, n18957, n18958, n18959, n18960, n18961,
    n18962, n18963, n18964, n18965, n18966, n18967,
    n18968, n18969, n18970, n18971, n18972, n18973,
    n18974, n18975, n18976, n18977, n18978, n18979,
    n18980, n18981, n18982, n18983, n18984, n18985,
    n18986, n18987, n18988, n18989, n18990, n18991,
    n18992, n18993, n18994, n18995, n18996, n18997,
    n18998, n18999, n19000, n19001, n19002, n19003,
    n19004, n19005, n19006, n19007, n19008, n19009,
    n19010, n19011, n19012, n19013, n19014, n19015,
    n19016, n19017, n19018, n19019, n19020, n19021,
    n19022, n19023, n19024, n19025, n19026, n19027,
    n19028, n19029, n19030, n19031, n19032, n19033,
    n19034, n19035, n19036, n19037, n19038, n19039,
    n19040, n19041, n19042, n19043, n19044, n19045,
    n19046, n19047, n19048, n19049, n19050, n19051,
    n19052, n19053, n19054, n19055, n19056, n19057,
    n19058, n19059, n19060, n19061, n19062, n19063,
    n19064, n19065, n19066, n19067, n19068, n19069,
    n19070, n19071, n19072, n19073, n19074, n19075,
    n19076, n19077, n19078, n19079, n19080, n19081,
    n19082, n19083, n19084, n19085, n19086, n19087,
    n19088, n19089, n19090, n19091, n19092, n19093,
    n19094, n19095, n19096, n19097, n19098, n19099,
    n19100, n19101, n19102, n19103, n19104, n19105,
    n19106, n19107, n19108, n19109, n19110, n19111,
    n19112, n19113, n19114, n19115, n19116, n19117,
    n19118, n19119, n19120, n19121, n19122, n19123,
    n19124, n19125, n19126, n19127, n19128, n19129,
    n19130, n19131, n19132, n19133, n19134, n19135,
    n19136, n19137, n19138, n19139, n19140, n19141,
    n19142, n19143, n19144, n19145, n19146, n19147,
    n19148, n19149, n19150, n19151, n19152, n19153,
    n19154, n19155, n19156, n19157, n19158, n19159,
    n19160, n19161, n19162, n19163, n19164, n19165,
    n19166, n19167, n19168, n19169, n19170, n19171,
    n19172, n19173, n19174, n19175, n19176, n19177,
    n19178, n19179, n19180, n19181, n19182, n19183,
    n19184, n19185, n19186, n19187, n19188, n19189,
    n19190, n19191, n19192, n19193, n19194, n19195,
    n19196, n19197, n19198, n19199, n19200, n19201,
    n19202, n19203, n19204, n19205, n19206, n19207,
    n19208, n19209, n19210, n19211, n19212, n19213,
    n19214, n19215, n19216, n19217, n19218, n19219,
    n19220, n19221, n19222, n19223, n19224, n19225,
    n19226, n19227, n19228, n19229, n19230, n19231,
    n19232, n19233, n19234, n19235, n19236, n19237,
    n19238, n19239, n19240, n19241, n19242, n19243,
    n19244, n19245, n19246, n19247, n19248, n19249,
    n19250, n19251, n19252, n19253, n19254, n19255,
    n19256, n19257, n19258, n19259, n19260, n19261,
    n19262, n19263, n19264, n19265, n19266, n19267,
    n19268, n19269, n19270, n19271, n19272, n19273,
    n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19282, n19283, n19284, n19285,
    n19286, n19287, n19288, n19289, n19290, n19291,
    n19292, n19293, n19294, n19295, n19296, n19297,
    n19298, n19299, n19300, n19301, n19302, n19303,
    n19304, n19305, n19306, n19307, n19308, n19309,
    n19310, n19311, n19312, n19313, n19314, n19315,
    n19316, n19317, n19318, n19319, n19320, n19321,
    n19322, n19323, n19324, n19325, n19326, n19327,
    n19328, n19329, n19330, n19331, n19332, n19333,
    n19334, n19335, n19336, n19337, n19338, n19339,
    n19340, n19341, n19342, n19343, n19344, n19345,
    n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357,
    n19358, n19359, n19360, n19361, n19362, n19363,
    n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19372, n19373, n19374, n19375,
    n19376, n19377, n19378, n19379, n19380, n19381,
    n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19391, n19392, n19393,
    n19394, n19395, n19396, n19397, n19398, n19399,
    n19400, n19401, n19402, n19403, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411,
    n19412, n19413, n19414, n19415, n19416, n19417,
    n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429,
    n19430, n19431, n19432, n19433, n19434, n19435,
    n19436, n19437, n19438, n19439, n19440, n19441,
    n19442, n19443, n19444, n19445, n19446, n19447,
    n19448, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459,
    n19460, n19461, n19462, n19463, n19464, n19465,
    n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19477,
    n19478, n19479, n19480, n19481, n19482, n19483,
    n19484, n19485, n19486, n19487, n19488, n19489,
    n19490, n19491, n19492, n19493, n19494, n19495,
    n19496, n19497, n19498, n19499, n19500, n19501,
    n19502, n19503, n19504, n19505, n19506, n19507,
    n19508, n19509, n19510, n19511, n19512, n19513,
    n19514, n19515, n19516, n19517, n19518, n19519,
    n19520, n19521, n19522, n19523, n19524, n19525,
    n19526, n19527, n19528, n19529, n19530, n19531,
    n19532, n19533, n19534, n19535, n19536, n19537,
    n19538, n19539, n19540, n19541, n19542, n19543,
    n19544, n19545, n19546, n19547, n19548, n19549,
    n19550, n19551, n19552, n19553, n19554, n19555,
    n19556, n19557, n19558, n19559, n19560, n19561,
    n19562, n19563, n19564, n19565, n19566, n19567,
    n19568, n19569, n19570, n19571, n19572, n19573,
    n19574, n19575, n19576, n19577, n19578, n19579,
    n19580, n19581, n19582, n19583, n19584, n19585,
    n19586, n19587, n19588, n19589, n19590, n19591,
    n19592, n19593, n19594, n19595, n19596, n19597,
    n19598, n19599, n19600, n19601, n19602, n19603,
    n19604, n19605, n19606, n19607, n19608, n19609,
    n19610, n19611, n19612, n19613, n19614, n19615,
    n19616, n19617, n19618, n19619, n19620, n19621,
    n19622, n19623, n19624, n19625, n19626, n19627,
    n19628, n19629, n19630, n19631, n19632, n19633,
    n19634, n19635, n19636, n19637, n19638, n19639,
    n19640, n19641, n19642, n19643, n19644, n19645,
    n19646, n19647, n19648, n19649, n19650, n19651,
    n19652, n19653, n19654, n19655, n19656, n19657,
    n19658, n19659, n19660, n19661, n19662, n19663,
    n19664, n19665, n19666, n19667, n19668, n19669,
    n19670, n19671, n19672, n19673, n19674, n19675,
    n19676, n19677, n19678, n19679, n19680, n19681,
    n19682, n19683, n19684, n19685, n19686, n19687,
    n19688, n19689, n19690, n19691, n19692, n19693,
    n19694, n19695, n19696, n19697, n19698, n19699,
    n19700, n19701, n19702, n19703, n19704, n19705,
    n19706, n19707, n19708, n19709, n19710, n19711,
    n19712, n19713, n19714, n19715, n19716, n19717,
    n19718, n19719, n19720, n19721, n19722, n19723,
    n19724, n19725, n19726, n19727, n19728, n19729,
    n19730, n19731, n19732, n19733, n19734, n19735,
    n19736, n19737, n19738, n19739, n19740, n19741,
    n19742, n19743, n19744, n19745, n19746, n19747,
    n19748, n19749, n19750, n19751, n19752, n19753,
    n19754, n19755, n19756, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765,
    n19766, n19767, n19768, n19769, n19770, n19771,
    n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783,
    n19784, n19785, n19786, n19787, n19788, n19789,
    n19790, n19791, n19792, n19793, n19794, n19795,
    n19796, n19797, n19798, n19799, n19800, n19801,
    n19802, n19803, n19804, n19805, n19806, n19807,
    n19808, n19809, n19810, n19811, n19812, n19813,
    n19814, n19815, n19816, n19817, n19818, n19819,
    n19820, n19821, n19822, n19823, n19824, n19825,
    n19826, n19827, n19828, n19829, n19830, n19831,
    n19832, n19833, n19834, n19835, n19836, n19837,
    n19838, n19839, n19840, n19841, n19842, n19843,
    n19844, n19845, n19846, n19847, n19848, n19849,
    n19850, n19851, n19852, n19853, n19854, n19855,
    n19856, n19857, n19858, n19859, n19860, n19861,
    n19862, n19863, n19864, n19865, n19866, n19867,
    n19868, n19869, n19870, n19871, n19872, n19873,
    n19874, n19875, n19876, n19877, n19878, n19879,
    n19880, n19881, n19882, n19883, n19884, n19885,
    n19886, n19887, n19888, n19889, n19890, n19891,
    n19892, n19893, n19894, n19895, n19896, n19897,
    n19898, n19899, n19900, n19901, n19902, n19903,
    n19904, n19905, n19906, n19907, n19908, n19909,
    n19910, n19911, n19912, n19913, n19914, n19915,
    n19916, n19917, n19918, n19919, n19920, n19921,
    n19922, n19923, n19924, n19925, n19926, n19927,
    n19928, n19929, n19930, n19931, n19932, n19933,
    n19934, n19935, n19936, n19937, n19938, n19939,
    n19940, n19941, n19942, n19943, n19944, n19945,
    n19946, n19947, n19948, n19949, n19950, n19951,
    n19952, n19953, n19954, n19955, n19956, n19957,
    n19958, n19959, n19960, n19961, n19962, n19963,
    n19964, n19965, n19966, n19967, n19968, n19969,
    n19970, n19971, n19972, n19973, n19974, n19975,
    n19976, n19977, n19978, n19979, n19980, n19981,
    n19982, n19983, n19984, n19985, n19986, n19987,
    n19988, n19989, n19990, n19991, n19992, n19993,
    n19994, n19995, n19996, n19997, n19998, n19999,
    n20000, n20001, n20002, n20003, n20004, n20005,
    n20006, n20007, n20008, n20009, n20010, n20011,
    n20012, n20013, n20014, n20015, n20016, n20017,
    n20018, n20019, n20020, n20021, n20022, n20023,
    n20024, n20025, n20026, n20027, n20028, n20029,
    n20030, n20031, n20032, n20033, n20034, n20035,
    n20036, n20037, n20038, n20039, n20040, n20041,
    n20042, n20043, n20044, n20045, n20046, n20047,
    n20048, n20049, n20050, n20051, n20052, n20053,
    n20054, n20055, n20056, n20057, n20058, n20059,
    n20060, n20061, n20062, n20063, n20064, n20065,
    n20066, n20067, n20068, n20069, n20070, n20071,
    n20072, n20073, n20074, n20075, n20076, n20077,
    n20078, n20079, n20080, n20081, n20082, n20083,
    n20084, n20085, n20086, n20087, n20088, n20089,
    n20090, n20091, n20092, n20093, n20094, n20095,
    n20096, n20097, n20098, n20099, n20100, n20101,
    n20102, n20103, n20104, n20105, n20106, n20107,
    n20108, n20109, n20110, n20111, n20112, n20113,
    n20114, n20115, n20116, n20117, n20118, n20119,
    n20120, n20121, n20122, n20123, n20124, n20125,
    n20126, n20127, n20128, n20129, n20130, n20131,
    n20132, n20133, n20134, n20135, n20136, n20137,
    n20138, n20139, n20140, n20141, n20142, n20143,
    n20144, n20145, n20146, n20147, n20148, n20149,
    n20150, n20151, n20152, n20153, n20154, n20155,
    n20156, n20157, n20158, n20159, n20160, n20161,
    n20162, n20163, n20164, n20165, n20166, n20167,
    n20168, n20169, n20170, n20171, n20172, n20173,
    n20174, n20175, n20176, n20177, n20178, n20179,
    n20180, n20181, n20182, n20183, n20184, n20185,
    n20186, n20187, n20188, n20189, n20190, n20191,
    n20192, n20193, n20194, n20195, n20196, n20197,
    n20198, n20199, n20200, n20201, n20202, n20203,
    n20204, n20205, n20206, n20207, n20208, n20209,
    n20210, n20211, n20212, n20213, n20214, n20215,
    n20216, n20217, n20218, n20219, n20220, n20221,
    n20222, n20223, n20224, n20225, n20226, n20227,
    n20228, n20229, n20230, n20231, n20232, n20233,
    n20234, n20235, n20236, n20237, n20238, n20239,
    n20240, n20241, n20242, n20243, n20244, n20245,
    n20246, n20247, n20248, n20249, n20250, n20251,
    n20252, n20253, n20254, n20255, n20256, n20257,
    n20258, n20259, n20260, n20261, n20262, n20263,
    n20264, n20265, n20266, n20267, n20268, n20269,
    n20270, n20271, n20272, n20273, n20274, n20275,
    n20276, n20277, n20278, n20279, n20280, n20281,
    n20282, n20283, n20284, n20285, n20286, n20287,
    n20288, n20289, n20290, n20291, n20292, n20293,
    n20294, n20295, n20296, n20297, n20298, n20299,
    n20300, n20301, n20302, n20303, n20304, n20305,
    n20306, n20307, n20308, n20309, n20310, n20311,
    n20312, n20313, n20314, n20315, n20316, n20317,
    n20318, n20319, n20320, n20321, n20322, n20323,
    n20324, n20325, n20326, n20327, n20328, n20329,
    n20330, n20331, n20332, n20333, n20334, n20335,
    n20336, n20337, n20338, n20339, n20340, n20341,
    n20342, n20343, n20344, n20345, n20346, n20347,
    n20348, n20349, n20350, n20351, n20352, n20353,
    n20354, n20355, n20356, n20357, n20358, n20359,
    n20360, n20361, n20362, n20363, n20364, n20365,
    n20366, n20367, n20368, n20369, n20370, n20371,
    n20372, n20373, n20374, n20375, n20376, n20377,
    n20378, n20379, n20380, n20381, n20382, n20383,
    n20384, n20385, n20386, n20387, n20388, n20389,
    n20390, n20391, n20392, n20393, n20394, n20395,
    n20396, n20397, n20398, n20399, n20400, n20401,
    n20402, n20403, n20404, n20405, n20406, n20407,
    n20408, n20409, n20410, n20411, n20412, n20413,
    n20414, n20415, n20416, n20417, n20418, n20419,
    n20420, n20421, n20422, n20423, n20424, n20425,
    n20426, n20427, n20428, n20429, n20430, n20431,
    n20432, n20433, n20434, n20435, n20436, n20437,
    n20438, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449,
    n20450, n20451, n20452, n20453, n20454, n20455,
    n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467,
    n20468, n20469, n20470, n20471, n20472, n20473,
    n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485,
    n20486, n20487, n20488, n20489, n20490, n20491,
    n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503,
    n20504, n20505, n20506, n20507, n20508, n20509,
    n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521,
    n20522, n20523, n20524, n20525, n20526, n20527,
    n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539,
    n20540, n20541, n20542, n20543, n20544, n20545,
    n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557,
    n20558, n20559, n20560, n20561, n20562, n20563,
    n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581,
    n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599,
    n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617,
    n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635,
    n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647,
    n20648, n20649, n20650, n20651, n20652, n20653,
    n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665,
    n20666, n20667, n20668, n20669, n20670, n20671,
    n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689,
    n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701,
    n20702, n20703, n20704, n20705, n20706, n20707,
    n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719,
    n20720, n20721, n20722, n20723, n20724, n20725,
    n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737,
    n20738, n20739, n20740, n20741, n20742, n20743,
    n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755,
    n20756, n20757, n20758, n20759, n20760, n20761,
    n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773,
    n20774, n20775, n20776, n20777, n20778, n20779,
    n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791,
    n20792, n20793, n20794, n20795, n20796, n20797,
    n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809,
    n20810, n20811, n20812, n20813, n20814, n20815,
    n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827,
    n20828, n20829, n20830, n20831, n20832, n20833,
    n20834, n20835, n20836, n20837, n20838, n20839,
    n20840, n20841, n20842, n20843, n20844, n20845,
    n20846, n20847, n20848, n20849, n20850, n20851,
    n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863,
    n20864, n20865, n20866, n20867, n20868, n20869,
    n20870, n20871, n20872, n20873, n20874, n20875,
    n20876, n20877, n20878, n20879, n20880, n20881,
    n20882, n20883, n20884, n20885, n20886, n20887,
    n20888, n20889, n20890, n20891, n20892, n20893,
    n20894, n20895, n20896, n20897, n20898, n20899,
    n20900, n20901, n20902, n20903, n20904, n20905,
    n20906, n20907, n20908, n20909, n20910, n20911,
    n20912, n20913, n20914, n20915, n20916, n20917,
    n20918, n20919, n20920, n20921, n20922, n20923,
    n20924, n20925, n20926, n20927, n20928, n20929,
    n20930, n20931, n20932, n20933, n20934, n20935,
    n20936, n20937, n20938, n20939, n20940, n20941,
    n20942, n20943, n20944, n20945, n20946, n20947,
    n20948, n20949, n20950, n20951, n20952, n20953,
    n20954, n20955, n20956, n20957, n20958, n20959,
    n20960, n20961, n20962, n20963, n20964, n20965,
    n20966, n20967, n20968, n20969, n20970, n20971,
    n20972, n20973, n20974, n20975, n20976, n20977,
    n20978, n20979, n20980, n20981, n20982, n20983,
    n20984, n20985, n20986, n20987, n20988, n20989,
    n20990, n20991, n20992, n20993, n20994, n20995,
    n20996, n20997, n20998, n20999, n21000, n21001,
    n21002, n21003, n21004, n21005, n21006, n21007,
    n21008, n21009, n21010, n21011, n21012, n21013,
    n21014, n21015, n21016, n21017, n21018, n21019,
    n21020, n21021, n21022, n21023, n21024, n21025,
    n21026, n21027, n21028, n21029, n21030, n21031,
    n21032, n21033, n21034, n21035, n21036, n21037,
    n21038, n21039, n21040, n21041, n21042, n21043,
    n21044, n21045, n21046, n21047, n21048, n21049,
    n21050, n21051, n21052, n21053, n21054, n21055,
    n21056, n21057, n21058, n21059, n21060, n21061,
    n21062, n21063, n21064, n21065, n21066, n21067,
    n21068, n21069, n21070, n21071, n21072, n21073,
    n21074, n21075, n21076, n21077, n21078, n21079,
    n21080, n21081, n21082, n21083, n21084, n21085,
    n21086, n21087, n21088, n21089, n21090, n21091,
    n21092, n21093, n21094, n21095, n21096, n21097,
    n21098, n21099, n21100, n21101, n21102, n21103,
    n21104, n21105, n21106, n21107, n21108, n21109,
    n21110, n21111, n21112, n21113, n21114, n21115,
    n21116, n21117, n21118, n21119, n21120, n21121,
    n21122, n21123, n21124, n21125, n21126, n21127,
    n21128, n21129, n21130, n21131, n21132, n21133,
    n21134, n21135, n21136, n21137, n21138, n21139,
    n21140, n21141, n21142, n21143, n21144, n21145,
    n21146, n21147, n21148, n21149, n21150, n21151,
    n21152, n21153, n21154, n21155, n21156, n21157,
    n21158, n21159, n21160, n21161, n21162, n21163,
    n21164, n21165, n21166, n21167, n21168, n21169,
    n21170, n21171, n21172, n21173, n21174, n21175,
    n21176, n21177, n21178, n21179, n21180, n21181,
    n21182, n21183, n21184, n21185, n21186, n21187,
    n21188, n21189, n21190, n21191, n21192, n21193,
    n21194, n21195, n21196, n21197, n21198, n21199,
    n21200, n21201, n21202, n21203, n21204, n21205,
    n21206, n21207, n21208, n21209, n21210, n21211,
    n21212, n21213, n21214, n21215, n21216, n21217,
    n21218, n21219, n21220, n21221, n21222, n21223,
    n21224, n21225, n21226, n21227, n21228, n21229,
    n21230, n21231, n21232, n21233, n21234, n21235,
    n21236, n21237, n21238, n21239, n21240, n21241,
    n21242, n21243, n21244, n21245, n21246, n21247,
    n21248, n21249, n21250, n21251, n21252, n21253,
    n21254, n21255, n21256, n21257, n21258, n21259,
    n21260, n21261, n21262, n21263, n21264, n21265,
    n21266, n21267, n21268, n21269, n21270, n21271,
    n21272, n21273, n21274, n21275, n21276, n21277,
    n21278, n21279, n21280, n21281, n21282, n21283,
    n21284, n21285, n21286, n21287, n21288, n21289,
    n21290, n21291, n21292, n21293, n21294, n21295,
    n21296, n21297, n21298, n21299, n21300, n21301,
    n21302, n21303, n21304, n21305, n21306, n21307,
    n21308, n21309, n21310, n21311, n21312, n21313,
    n21314, n21315, n21316, n21317, n21318, n21319,
    n21320, n21321, n21322, n21323, n21324, n21325,
    n21326, n21327, n21328, n21329, n21330, n21331,
    n21332, n21333, n21334, n21335, n21336, n21337,
    n21338, n21339, n21340, n21341, n21342, n21343,
    n21344, n21345, n21346, n21347, n21348, n21349,
    n21350, n21351, n21352, n21353, n21354, n21355,
    n21356, n21357, n21358, n21359, n21360, n21361,
    n21362, n21363, n21364, n21365, n21366, n21367,
    n21368, n21369, n21370, n21371, n21372, n21373,
    n21374, n21375, n21376, n21377, n21378, n21379,
    n21380, n21381, n21382, n21383, n21384, n21385,
    n21386, n21387, n21388, n21389, n21390, n21391,
    n21392, n21393, n21394, n21395, n21396, n21397,
    n21398, n21399, n21400, n21401, n21402, n21403,
    n21404, n21405, n21406, n21407, n21408, n21409,
    n21410, n21411, n21412, n21413, n21414, n21415,
    n21416, n21417, n21418, n21419, n21420, n21421,
    n21422, n21423, n21424, n21425, n21426, n21427,
    n21428, n21429, n21430, n21431, n21432, n21433,
    n21434, n21435, n21436, n21437, n21438, n21439,
    n21440, n21441, n21442, n21443, n21444, n21445,
    n21446, n21447, n21448, n21449, n21450, n21451,
    n21452, n21453, n21454, n21455, n21456, n21457,
    n21458, n21459, n21460, n21461, n21462, n21463,
    n21464, n21465, n21466, n21467, n21468, n21469,
    n21470, n21471, n21472, n21473, n21474, n21475,
    n21476, n21477, n21478, n21479, n21480, n21481,
    n21482, n21483, n21484, n21485, n21486, n21487,
    n21488, n21489, n21490, n21491, n21492, n21493,
    n21494, n21495, n21496, n21497, n21498, n21499,
    n21500, n21501, n21502, n21503, n21504, n21505,
    n21506, n21507, n21508, n21509, n21510, n21511,
    n21512, n21513, n21514, n21515, n21516, n21517,
    n21518, n21519, n21520, n21521, n21522, n21523,
    n21524, n21525, n21526, n21527, n21528, n21529,
    n21530, n21531, n21532, n21533, n21534, n21535,
    n21536, n21537, n21538, n21539, n21540, n21541,
    n21542, n21543, n21544, n21545, n21546, n21547,
    n21548, n21549, n21550, n21551, n21552, n21553,
    n21554, n21555, n21556, n21557, n21558, n21559,
    n21560, n21561, n21562, n21563, n21564, n21565,
    n21566, n21567, n21568, n21569, n21570, n21571,
    n21572, n21573, n21574, n21575, n21576, n21577,
    n21578, n21579, n21580, n21581, n21582, n21583,
    n21584, n21585, n21586, n21587, n21588, n21589,
    n21590, n21591, n21592, n21593, n21594, n21595,
    n21596, n21597, n21598, n21599, n21600, n21601,
    n21602, n21603, n21604, n21605, n21606, n21607,
    n21608, n21609, n21610, n21611, n21612, n21613,
    n21614, n21615, n21616, n21617, n21618, n21619,
    n21620, n21621, n21622, n21623, n21624, n21625,
    n21626, n21627, n21628, n21629, n21630, n21631,
    n21632, n21633, n21634, n21635, n21636, n21637,
    n21638, n21639, n21640, n21641, n21642, n21643,
    n21644, n21645, n21646, n21647, n21648, n21649,
    n21650, n21651, n21652, n21653, n21654, n21655,
    n21656, n21657, n21658, n21659, n21660, n21661,
    n21662, n21663, n21664, n21665, n21666, n21667,
    n21668, n21669, n21670, n21671, n21672, n21673,
    n21674, n21675, n21676, n21677, n21678, n21679,
    n21680, n21681, n21682, n21683, n21684, n21685,
    n21686, n21687, n21688, n21689, n21690, n21691,
    n21692, n21693, n21694, n21695, n21696, n21697,
    n21698, n21699, n21700, n21701, n21702, n21703,
    n21704, n21705, n21706, n21707, n21708, n21709,
    n21710, n21711, n21712, n21713, n21714, n21715,
    n21716, n21717, n21718, n21719, n21720, n21721,
    n21722, n21723, n21724, n21725, n21726, n21727,
    n21728, n21729, n21730, n21731, n21732, n21733,
    n21734, n21735, n21736, n21737, n21738, n21739,
    n21740, n21741, n21742, n21743, n21744, n21745,
    n21746, n21747, n21748, n21749, n21750, n21751,
    n21752, n21753, n21754, n21755, n21756, n21757,
    n21758, n21759, n21760, n21761, n21762, n21763,
    n21764, n21765, n21766, n21767, n21768, n21769,
    n21770, n21771, n21772, n21773, n21774, n21775,
    n21776, n21777, n21778, n21779, n21780, n21781,
    n21782, n21783, n21784, n21785, n21786, n21787,
    n21788, n21789, n21790, n21791, n21792, n21793,
    n21794, n21795, n21796, n21797, n21798, n21799,
    n21800, n21801, n21802, n21803, n21804, n21805,
    n21806, n21807, n21808, n21809, n21810, n21811,
    n21812, n21813, n21814, n21815, n21816, n21817,
    n21818, n21819, n21820, n21821, n21822, n21823,
    n21824, n21825, n21826, n21827, n21828, n21829,
    n21830, n21831, n21832, n21833, n21834, n21835,
    n21836, n21837, n21838, n21839, n21840, n21841,
    n21842, n21843, n21844, n21845, n21846, n21847,
    n21848, n21849, n21850, n21851, n21852, n21853,
    n21854, n21855, n21856, n21857, n21858, n21859,
    n21860, n21861, n21862, n21863, n21864, n21865,
    n21866, n21867, n21868, n21869, n21870, n21871,
    n21872, n21873, n21874, n21875, n21876, n21877,
    n21878, n21879, n21880, n21881, n21882, n21883,
    n21884, n21885, n21886, n21887, n21888, n21889,
    n21890, n21891, n21892, n21893, n21894, n21895,
    n21896, n21897, n21898, n21899, n21900, n21901,
    n21902, n21903, n21904, n21905, n21906, n21907,
    n21908, n21909, n21910, n21911, n21912, n21913,
    n21914, n21915, n21916, n21917, n21918, n21919,
    n21920, n21921, n21922, n21923, n21924, n21925,
    n21926, n21927, n21928, n21929, n21930, n21931,
    n21932, n21933, n21934, n21935, n21936, n21937,
    n21938, n21939, n21940, n21941, n21942, n21943,
    n21944, n21945, n21946, n21947, n21948, n21949,
    n21950, n21951, n21952, n21953, n21954, n21955,
    n21956, n21957, n21958, n21959, n21960, n21961,
    n21962, n21963, n21964, n21965, n21966, n21967,
    n21968, n21969, n21970, n21971, n21972, n21973,
    n21974, n21975, n21976, n21977, n21978, n21979,
    n21980, n21981, n21982, n21983, n21984, n21985,
    n21986, n21987, n21988, n21989, n21990, n21991,
    n21992, n21993, n21994, n21995, n21996, n21997,
    n21998, n21999, n22000, n22001, n22002, n22003,
    n22004, n22005, n22006, n22007, n22008, n22009,
    n22010, n22011, n22012, n22013, n22014, n22015,
    n22016, n22017, n22018, n22019, n22020, n22021,
    n22022, n22023, n22024, n22025, n22026, n22027,
    n22028, n22029, n22030, n22031, n22032, n22033,
    n22034, n22035, n22036, n22037, n22038, n22039,
    n22040, n22041, n22042, n22043, n22044, n22045,
    n22046, n22047, n22048, n22049, n22050, n22051,
    n22052, n22053, n22054, n22055, n22056, n22057,
    n22058, n22059, n22060, n22061, n22062, n22063,
    n22064, n22065, n22066, n22067, n22068, n22069,
    n22070, n22071, n22072, n22073, n22074, n22075,
    n22076, n22077, n22078, n22079, n22080, n22081,
    n22082, n22083, n22084, n22085, n22086, n22087,
    n22088, n22089, n22090, n22091, n22092, n22093,
    n22094, n22095, n22096, n22097, n22098, n22099,
    n22100, n22101, n22102, n22103, n22104, n22105,
    n22106, n22107, n22108, n22109, n22110, n22111,
    n22112, n22113, n22114, n22115, n22116, n22117,
    n22118, n22119, n22120, n22121, n22122, n22123,
    n22124, n22125, n22126, n22127, n22128, n22129,
    n22130, n22131, n22132, n22133, n22134, n22135,
    n22136, n22137, n22138, n22139, n22140, n22141,
    n22142, n22143, n22144, n22145, n22146, n22147,
    n22148, n22149, n22150, n22151, n22152, n22153,
    n22154, n22155, n22156, n22157, n22158, n22159,
    n22160, n22161, n22162, n22163, n22164, n22165,
    n22166, n22167, n22168, n22169, n22170, n22171,
    n22172, n22173, n22174, n22175, n22176, n22177,
    n22178, n22179, n22180, n22181, n22182, n22183,
    n22184, n22185, n22186, n22187, n22188, n22189,
    n22190, n22191, n22192, n22193, n22194, n22195,
    n22196, n22197, n22198, n22199, n22200, n22201,
    n22202, n22203, n22204, n22205, n22206, n22207,
    n22208, n22209, n22210, n22211, n22212, n22213,
    n22214, n22215, n22216, n22217, n22218, n22219,
    n22220, n22221, n22222, n22223, n22224, n22225,
    n22226, n22227, n22228, n22229, n22230, n22231,
    n22232, n22233, n22234, n22235, n22236, n22237,
    n22238, n22239, n22240, n22241, n22242, n22243,
    n22244, n22245, n22246, n22247, n22248, n22249,
    n22250, n22251, n22252, n22253, n22254, n22255,
    n22256, n22257, n22258, n22259, n22260, n22261,
    n22262, n22263, n22264, n22265, n22266, n22267,
    n22268, n22269, n22270, n22271, n22272, n22273,
    n22274, n22275, n22276, n22277, n22278, n22279,
    n22280, n22281, n22282, n22283, n22284, n22285,
    n22286, n22287, n22288, n22289, n22290, n22291,
    n22292, n22293, n22294, n22295, n22296, n22297,
    n22298, n22299, n22300, n22301, n22302, n22303,
    n22304, n22305, n22306, n22307, n22308, n22309,
    n22310, n22311, n22312, n22313, n22314, n22315,
    n22316, n22317, n22318, n22319, n22320, n22321,
    n22322, n22323, n22324, n22325, n22326, n22327,
    n22328, n22329, n22330, n22331, n22332, n22333,
    n22334, n22335, n22336, n22337, n22338, n22339,
    n22340, n22341, n22342, n22343, n22344, n22345,
    n22346, n22347, n22348, n22349, n22350, n22351,
    n22352, n22353, n22354, n22355, n22356, n22357,
    n22358, n22359, n22360, n22361, n22362, n22363,
    n22364, n22365, n22366, n22367, n22368, n22369,
    n22370, n22371, n22372, n22373, n22374, n22375,
    n22376, n22377, n22378, n22379, n22380, n22381,
    n22382, n22383, n22384, n22385, n22386, n22387,
    n22388, n22389, n22390, n22391, n22392, n22393,
    n22394, n22395, n22396, n22397, n22398, n22399,
    n22400, n22401, n22402, n22403, n22404, n22405,
    n22406, n22407, n22408, n22409, n22410, n22411,
    n22412, n22413, n22414, n22415, n22416, n22417,
    n22418, n22419, n22420, n22421, n22422, n22423,
    n22424, n22425, n22426, n22427, n22428, n22429,
    n22430, n22431, n22432, n22433, n22434, n22435,
    n22436, n22437, n22438, n22439, n22440, n22441,
    n22442, n22443, n22444, n22445, n22446, n22447,
    n22448, n22449, n22450, n22451, n22452, n22453,
    n22454, n22455, n22456, n22457, n22458, n22459,
    n22460, n22461, n22462, n22463, n22464, n22465,
    n22466, n22467, n22468, n22469, n22470, n22471,
    n22472, n22473, n22474, n22475, n22476, n22477,
    n22478, n22479, n22480, n22481, n22482, n22483,
    n22484, n22485, n22486, n22487, n22488, n22489,
    n22490, n22491, n22492, n22493, n22494, n22495,
    n22496, n22497, n22498, n22499, n22500, n22501,
    n22502, n22503, n22504, n22505, n22506, n22507,
    n22508, n22509, n22510, n22511, n22512, n22513,
    n22514, n22515, n22516, n22517, n22518, n22519,
    n22520, n22521, n22522, n22523, n22524, n22525,
    n22526, n22527, n22528, n22529, n22530, n22531,
    n22532, n22533, n22534, n22535, n22536, n22537,
    n22538, n22539, n22540, n22541, n22542, n22543,
    n22544, n22545, n22546, n22547, n22548, n22549,
    n22550, n22551, n22552, n22553, n22554, n22555,
    n22556, n22557, n22558, n22559, n22560, n22561,
    n22562, n22563, n22564, n22565, n22566, n22567,
    n22568, n22569, n22570, n22571, n22572, n22573,
    n22574, n22575, n22576, n22577, n22578, n22579,
    n22580, n22581, n22582, n22583, n22584, n22585,
    n22586, n22587, n22588, n22589, n22590, n22591,
    n22592, n22593, n22594, n22595, n22596, n22597,
    n22598, n22599, n22600, n22601, n22602, n22603,
    n22604, n22605, n22606, n22607, n22608, n22609,
    n22610, n22611, n22612, n22613, n22614, n22615,
    n22616, n22617, n22618, n22619, n22620, n22621,
    n22622, n22623, n22624, n22625, n22626, n22627,
    n22628, n22629, n22630, n22631, n22632, n22633,
    n22634, n22635, n22636, n22637, n22638, n22639,
    n22640, n22641, n22642, n22643, n22644, n22645,
    n22646, n22647, n22648, n22649, n22650, n22651,
    n22652, n22653, n22654, n22655, n22656, n22657,
    n22658, n22659, n22660, n22661, n22662, n22663,
    n22664, n22665, n22666, n22667, n22668, n22669,
    n22670, n22671, n22672, n22673, n22674, n22675,
    n22676, n22677, n22678, n22679, n22680, n22681,
    n22682, n22683, n22684, n22685, n22686, n22687,
    n22688, n22689, n22690, n22691, n22692, n22693,
    n22694, n22695, n22696, n22697, n22698, n22699,
    n22700, n22701, n22702, n22703, n22704, n22705,
    n22706, n22707, n22708, n22709, n22710, n22711,
    n22712, n22713, n22714, n22715, n22716, n22717,
    n22718, n22719, n22720, n22721, n22722, n22723,
    n22724, n22725, n22726, n22727, n22728, n22729,
    n22730, n22731, n22732, n22733, n22734, n22735,
    n22736, n22737, n22738, n22739, n22740, n22741,
    n22742, n22743, n22744, n22745, n22746, n22747,
    n22748, n22749, n22750, n22751, n22752, n22753,
    n22754, n22755, n22756, n22757, n22758, n22759,
    n22760, n22761, n22762, n22763, n22764, n22765,
    n22766, n22767, n22768, n22769, n22770, n22771,
    n22772, n22773, n22774, n22775, n22776, n22777,
    n22778, n22779, n22780, n22781, n22782, n22783,
    n22784, n22785, n22786, n22787, n22788, n22789,
    n22790, n22791, n22792, n22793, n22794, n22795,
    n22796, n22797, n22798, n22799, n22800, n22801,
    n22802, n22803, n22804, n22805, n22806, n22807,
    n22808, n22809, n22810, n22811, n22812, n22813,
    n22814, n22815, n22816, n22817, n22818, n22819,
    n22820, n22821, n22822, n22823, n22824, n22825,
    n22826, n22827, n22828, n22829, n22830, n22831,
    n22832, n22833, n22834, n22835, n22836, n22837,
    n22838, n22839, n22840, n22841, n22842, n22843,
    n22844, n22845, n22846, n22847, n22848, n22849,
    n22850, n22851, n22852, n22853, n22854, n22855,
    n22856, n22857, n22858, n22859, n22860, n22861,
    n22862, n22863, n22864, n22865, n22866, n22867,
    n22868, n22869, n22870, n22871, n22872, n22873,
    n22874, n22875, n22876, n22877, n22878, n22879,
    n22880, n22881, n22882, n22883, n22884, n22885,
    n22886, n22887, n22888, n22889, n22890, n22891,
    n22892, n22893, n22894, n22895, n22896, n22897,
    n22898, n22899, n22900, n22901, n22902, n22903,
    n22904, n22905, n22906, n22907, n22908, n22909,
    n22910, n22911, n22912, n22913, n22914, n22915,
    n22916, n22917, n22918, n22919, n22920, n22921,
    n22922, n22923, n22924, n22925, n22926, n22927,
    n22928, n22929, n22930, n22931, n22932, n22933,
    n22934, n22935, n22936, n22937, n22938, n22939,
    n22940, n22941, n22942, n22943, n22944, n22945,
    n22946, n22947, n22948, n22949, n22950, n22951,
    n22952, n22953, n22954, n22955, n22956, n22957,
    n22958, n22959, n22960, n22961, n22962, n22963,
    n22964, n22965, n22966, n22967, n22968, n22969,
    n22970, n22971, n22972, n22973, n22974, n22975,
    n22976, n22977, n22978, n22979, n22980, n22981,
    n22982, n22983, n22984, n22985, n22986, n22987,
    n22988, n22989, n22990, n22991, n22992, n22993,
    n22994, n22995, n22996, n22997, n22998, n22999,
    n23000, n23001, n23002, n23003, n23004, n23005,
    n23006, n23007, n23008, n23009, n23010, n23011,
    n23012, n23013, n23014, n23015, n23016, n23017,
    n23018, n23019, n23020, n23021, n23022, n23023,
    n23024, n23025, n23026, n23027, n23028, n23029,
    n23030, n23031, n23032, n23033, n23034, n23035,
    n23036, n23037, n23038, n23039, n23040, n23041,
    n23042, n23043, n23044, n23045, n23046, n23047,
    n23048, n23049, n23050, n23051, n23052, n23053,
    n23054, n23055, n23056, n23057, n23058, n23059,
    n23060, n23061, n23062, n23063, n23064, n23065,
    n23066, n23067, n23068, n23069, n23070, n23071,
    n23072, n23073, n23074, n23075, n23076, n23077,
    n23078, n23079, n23080, n23081, n23082, n23083,
    n23084, n23085, n23086, n23087, n23088, n23089,
    n23090, n23091, n23092, n23093, n23094, n23095,
    n23096, n23097, n23098, n23099, n23100, n23101,
    n23102, n23103, n23104, n23105, n23106, n23107,
    n23108, n23109, n23110, n23111, n23112, n23113,
    n23114, n23115, n23116, n23117, n23118, n23119,
    n23120, n23121, n23122, n23123, n23124, n23125,
    n23126, n23127, n23128, n23129, n23130, n23131,
    n23132, n23133, n23134, n23135, n23136, n23137,
    n23138, n23139, n23140, n23141, n23142, n23143,
    n23144, n23145, n23146, n23147, n23148, n23149,
    n23150, n23151, n23152, n23153, n23154, n23155,
    n23156, n23157, n23158, n23159, n23160, n23161,
    n23162, n23163, n23164, n23165, n23166, n23167,
    n23168, n23169, n23170, n23171, n23172, n23173,
    n23174, n23175, n23176, n23177, n23178, n23179,
    n23180, n23181, n23182, n23183, n23184, n23185,
    n23186, n23187, n23188, n23189, n23190, n23191,
    n23192, n23193, n23194, n23195, n23196, n23197,
    n23198, n23199, n23200, n23201, n23202, n23203,
    n23204, n23205, n23206, n23207, n23208, n23209,
    n23210, n23211, n23212, n23213, n23214, n23215,
    n23216, n23217, n23218, n23219, n23220, n23221,
    n23222, n23223, n23224, n23225, n23226, n23227,
    n23228, n23229, n23230, n23231, n23232, n23233,
    n23234, n23235, n23236, n23237, n23238, n23239,
    n23240, n23241, n23242, n23243, n23244, n23245,
    n23246, n23247, n23248, n23249, n23250, n23251,
    n23252, n23253, n23254, n23255, n23256, n23257,
    n23258, n23259, n23260, n23261, n23262, n23263,
    n23264, n23265, n23266, n23267, n23268, n23269,
    n23270, n23271, n23272, n23273, n23274, n23275,
    n23276, n23277, n23278, n23279, n23280, n23281,
    n23282, n23283, n23284, n23285, n23286, n23287,
    n23288, n23289, n23290, n23291, n23292, n23293,
    n23294, n23295, n23296, n23297, n23298, n23299,
    n23300, n23301, n23302, n23303, n23304, n23305,
    n23306, n23307, n23308, n23309, n23310, n23311,
    n23312, n23313, n23314, n23315, n23316, n23317,
    n23318, n23319, n23320, n23321, n23322, n23323,
    n23324, n23325, n23326, n23327, n23328, n23329,
    n23330, n23331, n23332, n23333, n23334, n23335,
    n23336, n23337, n23338, n23339, n23340, n23341,
    n23342, n23343, n23344, n23345, n23346, n23347,
    n23348, n23349, n23350, n23351, n23352, n23353,
    n23354, n23355, n23356, n23357, n23358, n23359,
    n23360, n23361, n23362, n23363, n23364, n23365,
    n23366, n23367, n23368, n23369, n23370, n23371,
    n23372, n23373, n23374, n23375, n23376, n23377,
    n23378, n23379, n23380, n23381, n23382, n23383,
    n23384, n23385, n23386, n23387, n23388, n23389,
    n23390, n23391, n23392, n23393, n23394, n23395,
    n23396, n23397, n23398, n23399, n23400, n23401,
    n23402, n23403, n23404, n23405, n23406, n23407,
    n23408, n23409, n23410, n23411, n23412, n23413,
    n23414, n23415, n23416, n23417, n23418, n23419,
    n23420, n23421, n23422, n23423, n23424, n23425,
    n23426, n23427, n23428, n23429, n23430, n23431,
    n23432, n23433, n23434, n23435, n23436, n23437,
    n23438, n23439, n23440, n23441, n23442, n23443,
    n23444, n23445, n23446, n23447, n23448, n23449,
    n23450, n23451, n23452, n23453, n23454, n23455,
    n23456, n23457, n23458, n23459, n23460, n23461,
    n23462, n23463, n23464, n23465, n23466, n23467,
    n23468, n23469, n23470, n23471, n23472, n23473,
    n23474, n23475, n23476, n23477, n23478, n23479,
    n23480, n23481, n23482, n23483, n23484, n23485,
    n23486, n23487, n23488, n23489, n23490, n23491,
    n23492, n23493, n23494, n23495, n23496, n23497,
    n23498, n23499, n23500, n23501, n23502, n23503,
    n23504, n23505, n23506, n23507, n23508, n23509,
    n23510, n23511, n23512, n23513, n23514, n23515,
    n23516, n23517, n23518, n23519, n23520, n23521,
    n23522, n23523, n23524, n23525, n23526, n23527,
    n23528, n23529, n23530, n23531, n23532, n23533,
    n23534, n23535, n23536, n23537, n23538, n23539,
    n23540, n23541, n23542, n23543, n23544, n23545,
    n23546, n23547, n23548, n23549, n23550, n23551,
    n23552, n23553, n23554, n23555, n23556, n23557,
    n23558, n23559, n23560, n23561, n23562, n23563,
    n23564, n23565, n23566, n23567, n23568, n23569,
    n23570, n23571, n23572, n23573, n23574, n23575,
    n23576, n23577, n23578, n23579, n23580, n23581,
    n23582, n23583, n23584, n23585, n23586, n23587,
    n23588, n23589, n23590, n23591, n23592, n23593,
    n23594, n23595, n23596, n23597, n23598, n23599,
    n23600, n23601, n23602, n23603, n23604, n23605,
    n23606, n23607, n23608, n23609, n23610, n23611,
    n23612, n23613, n23614, n23615, n23616, n23617,
    n23618, n23619, n23620, n23621, n23622, n23623,
    n23624, n23625, n23626, n23627, n23628, n23629,
    n23630, n23631, n23632, n23633, n23634, n23635,
    n23636, n23637, n23638, n23639, n23640, n23641,
    n23642, n23643, n23644, n23645, n23646, n23647,
    n23648, n23649, n23650, n23651, n23652, n23653,
    n23654, n23655, n23656, n23657, n23658, n23659,
    n23660, n23661, n23662, n23663, n23664, n23665,
    n23666, n23667, n23668, n23669, n23670, n23671,
    n23672, n23673, n23674, n23675, n23676, n23677,
    n23678, n23679, n23680, n23681, n23682, n23683,
    n23684, n23685, n23686, n23687, n23688, n23689,
    n23690, n23691, n23692, n23693, n23694, n23695,
    n23696, n23697, n23698, n23699, n23700, n23701,
    n23702, n23703, n23704, n23705, n23706, n23707,
    n23708, n23709, n23710, n23711, n23712, n23713,
    n23714, n23715, n23716, n23717, n23718, n23719,
    n23720, n23721, n23722, n23723, n23724, n23725,
    n23726, n23727, n23728, n23729, n23730, n23731,
    n23732, n23733, n23734, n23735, n23736, n23737,
    n23738, n23739, n23740, n23741, n23742, n23743,
    n23744, n23745, n23746, n23747, n23748, n23749,
    n23750, n23751, n23752, n23753, n23754, n23755,
    n23756, n23757, n23758, n23759, n23760, n23761,
    n23762, n23763, n23764, n23765, n23766, n23767,
    n23768, n23769, n23770, n23771, n23772, n23773,
    n23774, n23775, n23776, n23777, n23778, n23779,
    n23780, n23781, n23782, n23783, n23784, n23785,
    n23786, n23787, n23788, n23789, n23790, n23791,
    n23792, n23793, n23794, n23795, n23796, n23797,
    n23798, n23799, n23800, n23801, n23802, n23803,
    n23804, n23805, n23806, n23807, n23808, n23809,
    n23810, n23811, n23812, n23813, n23814, n23815,
    n23816, n23817, n23818, n23819, n23820, n23821,
    n23822, n23823, n23824, n23825, n23826, n23827,
    n23828, n23829, n23830, n23831, n23832, n23833,
    n23834, n23835, n23836, n23837, n23838, n23839,
    n23840, n23841, n23842, n23843, n23844, n23845,
    n23846, n23847, n23848, n23849, n23850, n23851,
    n23852, n23853, n23854, n23855, n23856, n23857,
    n23858, n23859, n23860, n23861, n23862, n23863,
    n23864, n23865, n23866, n23867, n23868, n23869,
    n23870, n23871, n23872, n23873, n23874, n23875,
    n23876, n23877, n23878, n23879, n23880, n23881,
    n23882, n23883, n23884, n23885, n23886, n23887,
    n23888, n23889, n23890, n23891, n23892, n23893,
    n23894, n23895, n23896, n23897, n23898, n23899,
    n23900, n23901, n23902, n23903, n23904, n23905,
    n23906, n23907, n23908, n23909, n23910, n23911,
    n23912, n23913, n23914, n23915, n23916, n23917,
    n23918, n23919, n23920, n23921, n23922, n23923,
    n23924, n23925, n23926, n23927, n23928, n23929,
    n23930, n23931, n23932, n23933, n23934, n23935,
    n23936, n23937, n23938, n23939, n23940, n23941,
    n23942, n23943, n23944, n23945, n23946, n23947,
    n23948, n23949, n23950, n23951, n23952, n23953,
    n23954, n23955, n23956, n23957, n23958, n23959,
    n23960, n23961, n23962, n23963, n23964, n23965,
    n23966, n23967, n23968, n23969, n23970, n23971,
    n23972, n23973, n23974, n23975, n23976, n23977,
    n23978, n23979, n23980, n23981, n23982, n23983,
    n23984, n23985, n23986, n23987, n23988, n23989,
    n23990, n23991, n23992, n23993, n23994, n23995,
    n23996, n23997, n23998, n23999, n24000, n24001,
    n24002, n24003, n24004, n24005, n24006, n24007,
    n24008, n24009, n24010, n24011, n24012, n24013,
    n24014, n24015, n24016, n24017, n24018, n24019,
    n24020, n24021, n24022, n24023, n24024, n24025,
    n24026, n24027, n24028, n24029, n24030, n24031,
    n24032, n24033, n24034, n24035, n24036, n24037,
    n24038, n24039, n24040, n24041, n24042, n24043,
    n24044, n24045, n24046, n24047, n24048, n24049,
    n24050, n24051, n24052, n24053, n24054, n24055,
    n24056, n24057, n24058, n24059, n24060, n24061,
    n24062, n24063, n24064, n24065, n24066, n24067,
    n24068, n24069, n24070, n24071, n24072, n24073,
    n24074, n24075, n24076, n24077, n24078, n24079,
    n24080, n24081, n24082, n24083, n24084, n24085,
    n24086, n24087, n24088, n24089, n24090, n24091,
    n24092, n24093, n24094, n24095, n24096, n24097,
    n24098, n24099, n24100, n24101, n24102, n24103,
    n24104, n24105, n24106, n24107, n24108, n24109,
    n24110, n24111, n24112, n24113, n24114, n24115,
    n24116, n24117, n24118, n24119, n24120, n24121,
    n24122, n24123, n24124, n24125, n24126, n24127,
    n24128, n24129, n24130, n24131, n24132, n24133,
    n24134, n24135, n24136, n24137, n24138, n24139,
    n24140, n24141, n24142, n24143, n24144, n24145,
    n24146, n24147, n24148, n24149, n24150, n24151,
    n24152, n24153, n24154, n24155, n24156, n24157,
    n24158, n24159, n24160, n24161, n24162, n24163,
    n24164, n24165, n24166, n24167, n24168, n24169,
    n24170, n24171, n24172, n24173, n24174, n24175,
    n24176, n24177, n24178, n24179, n24180, n24181,
    n24182, n24183, n24184, n24185, n24186, n24187,
    n24188, n24189, n24190, n24191, n24192, n24193,
    n24194, n24195, n24196, n24197, n24198, n24199,
    n24200, n24201, n24202, n24203, n24204, n24205,
    n24206, n24207, n24208, n24209, n24210, n24211,
    n24212, n24213, n24214, n24215, n24216, n24217,
    n24218, n24219, n24220, n24221, n24222, n24223,
    n24224, n24225, n24226, n24227, n24228, n24229,
    n24230, n24231, n24232, n24233, n24234, n24235,
    n24236, n24237, n24238, n24239, n24240, n24241,
    n24242, n24243, n24244, n24245, n24246, n24247,
    n24248, n24249, n24250, n24251, n24252, n24253,
    n24254, n24255, n24256, n24257, n24258, n24259,
    n24260, n24261, n24262, n24263, n24264, n24265,
    n24266, n24267, n24268, n24269, n24270, n24271,
    n24272, n24273, n24274, n24275, n24276, n24277,
    n24278, n24279, n24280, n24281, n24282, n24283,
    n24284, n24285, n24286, n24287, n24288, n24289,
    n24290, n24291, n24292, n24293, n24294, n24295,
    n24296, n24297, n24298, n24299, n24300, n24301,
    n24302, n24303, n24304, n24305, n24306, n24307,
    n24308, n24309, n24310, n24311, n24312, n24313,
    n24314, n24315, n24316, n24317, n24318, n24319,
    n24320, n24321, n24322, n24323, n24324, n24325,
    n24326, n24327, n24328, n24329, n24330, n24331,
    n24332, n24333, n24334, n24335, n24336, n24337,
    n24338, n24339, n24340, n24341, n24342, n24343,
    n24344, n24345, n24346, n24347, n24348, n24349,
    n24350, n24351, n24352, n24353, n24354, n24355,
    n24356, n24357, n24358, n24359, n24360, n24361,
    n24362, n24363, n24364, n24365, n24366, n24367,
    n24368, n24369, n24370, n24371, n24372, n24373,
    n24374, n24375, n24376, n24377, n24378, n24379,
    n24380, n24381, n24382, n24383, n24384, n24385,
    n24386, n24387, n24388, n24389, n24390, n24391,
    n24392, n24393, n24394, n24395, n24396, n24397,
    n24398, n24399, n24400, n24401, n24402, n24403,
    n24404, n24405, n24406, n24407, n24408, n24409,
    n24410, n24411, n24412, n24413, n24414, n24415,
    n24416, n24417, n24418, n24419, n24420, n24421,
    n24422, n24423, n24424, n24425, n24426, n24427,
    n24428, n24429, n24430, n24431, n24432, n24433,
    n24434, n24435, n24436, n24437, n24438, n24439,
    n24440, n24441, n24442, n24443, n24444, n24445,
    n24446, n24447, n24448, n24449, n24450, n24451,
    n24452, n24453, n24454, n24455, n24456, n24457,
    n24458, n24459, n24460, n24461, n24462, n24463,
    n24464, n24465, n24466, n24467, n24468, n24469,
    n24470, n24471, n24472, n24473, n24474, n24475,
    n24476, n24477, n24478, n24479, n24480, n24481,
    n24482, n24483, n24484, n24485, n24486, n24487,
    n24488, n24489, n24490, n24491, n24492, n24493,
    n24494, n24495, n24496, n24497, n24498, n24499,
    n24500, n24501, n24502, n24503, n24504, n24505,
    n24506, n24507, n24508, n24509, n24510, n24511,
    n24512, n24513, n24514, n24515, n24516, n24517,
    n24518, n24519, n24520, n24521, n24522, n24523,
    n24524, n24525, n24526, n24527, n24528, n24529,
    n24530, n24531, n24532, n24533, n24534, n24535,
    n24536, n24537, n24538, n24539, n24540, n24541,
    n24542, n24543, n24544, n24545, n24546, n24547,
    n24548, n24549, n24550, n24551, n24552, n24553,
    n24554, n24555, n24556, n24557, n24558, n24559,
    n24560, n24561, n24562, n24563, n24564, n24565,
    n24566, n24567, n24568, n24569, n24570, n24571,
    n24572, n24573, n24574, n24575, n24576, n24577,
    n24578, n24579, n24580, n24581, n24582, n24583,
    n24584, n24585, n24586, n24587, n24588, n24589,
    n24590, n24591, n24592, n24593, n24594, n24595,
    n24596, n24597, n24598, n24599, n24600, n24601,
    n24602, n24603, n24604, n24605, n24606, n24607,
    n24608, n24609, n24610, n24611, n24612, n24613,
    n24614, n24615, n24616, n24617, n24618, n24619,
    n24620, n24621, n24622, n24623, n24624, n24625,
    n24626, n24627, n24628, n24629, n24630, n24631,
    n24632, n24633, n24634, n24635, n24636, n24637,
    n24638, n24639, n24640, n24641, n24642, n24643,
    n24644, n24645, n24646, n24647, n24648, n24649,
    n24650, n24651, n24652, n24653, n24654, n24655,
    n24656, n24657, n24658, n24659, n24660, n24661,
    n24662, n24663, n24664, n24665, n24666, n24667,
    n24668, n24669, n24670, n24671, n24672, n24673,
    n24674, n24675, n24676, n24677, n24678, n24679,
    n24680, n24681, n24682, n24683, n24684, n24685,
    n24686, n24687, n24688, n24689, n24690, n24691,
    n24692, n24693, n24694, n24695, n24696, n24697,
    n24698, n24699, n24700, n24701, n24702, n24703,
    n24704, n24705, n24706, n24707, n24708, n24709,
    n24710, n24711, n24712, n24713, n24714, n24715,
    n24716, n24717, n24718, n24719, n24720, n24721,
    n24722, n24723, n24724, n24725, n24726, n24727,
    n24728, n24729, n24730, n24731, n24732, n24733,
    n24734, n24735, n24736, n24737, n24738, n24739,
    n24740, n24741, n24742, n24743, n24744, n24745,
    n24746, n24747, n24748, n24749, n24750, n24751,
    n24752, n24753, n24754, n24755, n24756, n24757,
    n24758, n24759, n24760, n24761, n24762, n24763,
    n24764, n24765, n24766, n24767, n24768, n24769,
    n24770, n24771, n24772, n24773, n24774, n24775,
    n24776, n24777, n24778, n24779, n24780, n24781,
    n24782, n24783, n24784, n24785, n24786, n24787,
    n24788, n24789, n24790, n24791, n24792, n24793,
    n24794, n24795, n24796, n24797, n24798, n24799,
    n24800, n24801, n24802, n24803, n24804, n24805,
    n24806, n24807, n24808, n24809, n24810, n24811,
    n24812, n24813, n24814, n24815, n24816, n24817,
    n24818, n24819, n24820, n24821, n24822, n24823,
    n24824, n24825, n24826, n24827, n24828, n24829,
    n24830, n24831, n24832, n24833, n24834, n24835,
    n24836, n24837, n24838, n24839, n24840, n24841,
    n24842, n24843, n24844, n24845, n24846, n24847,
    n24848, n24849, n24850, n24851, n24852, n24853,
    n24854, n24855, n24856, n24857, n24858, n24859,
    n24860, n24861, n24862, n24863, n24864, n24865,
    n24866, n24867, n24868, n24869, n24870, n24871,
    n24872, n24873, n24874, n24875, n24876, n24877,
    n24878, n24879, n24880, n24881, n24882, n24883,
    n24884, n24885, n24886, n24887, n24888, n24889,
    n24890, n24891, n24892, n24893, n24894, n24895,
    n24896, n24897, n24898, n24899, n24900, n24901,
    n24902, n24903, n24904, n24905, n24906, n24907,
    n24908, n24909, n24910, n24911, n24912, n24913,
    n24914, n24915, n24916, n24917, n24918, n24919,
    n24920, n24921, n24922, n24923, n24924, n24925,
    n24926, n24927, n24928, n24929, n24930, n24931,
    n24932, n24933, n24934, n24935, n24936, n24937,
    n24938, n24939, n24940, n24941, n24942, n24943,
    n24944, n24945, n24946, n24947, n24948, n24949,
    n24950, n24951, n24952, n24953, n24954, n24955,
    n24956, n24957, n24958, n24959, n24960, n24961,
    n24962, n24963, n24964, n24965, n24966, n24967,
    n24968, n24969, n24970, n24971, n24972, n24973,
    n24974, n24975, n24976, n24977, n24978, n24979,
    n24980, n24981, n24982, n24983, n24984, n24985,
    n24986, n24987, n24988, n24989, n24990, n24991,
    n24992, n24993, n24994, n24995, n24996, n24997,
    n24998, n24999, n25000, n25001, n25002, n25003,
    n25004, n25005, n25006, n25007, n25008, n25009,
    n25010, n25011, n25012, n25013, n25014, n25015,
    n25016, n25017, n25018, n25019, n25020, n25021,
    n25022, n25023, n25024, n25025, n25026, n25027,
    n25028, n25029, n25030, n25031, n25032, n25033,
    n25034, n25035, n25036, n25037, n25038, n25039,
    n25040, n25041, n25042, n25043, n25044, n25045,
    n25046, n25047, n25048, n25049, n25050, n25051,
    n25052, n25053, n25054, n25055, n25056, n25057,
    n25058, n25059, n25060, n25061, n25062, n25063,
    n25064, n25065, n25066, n25067, n25068, n25069,
    n25070, n25071, n25072, n25073, n25074, n25075,
    n25076, n25077, n25078, n25079, n25080, n25081,
    n25082, n25083, n25084, n25085, n25086, n25087,
    n25088, n25089, n25090, n25091, n25092, n25093,
    n25094, n25095, n25096, n25097, n25098, n25099,
    n25100, n25101, n25102, n25103, n25104, n25105,
    n25106, n25107, n25108, n25109, n25110, n25111,
    n25112, n25113, n25114, n25115, n25116, n25117,
    n25118, n25119, n25120, n25121, n25122, n25123,
    n25124, n25125, n25126, n25127, n25128, n25129,
    n25130, n25131, n25132, n25133, n25134, n25135,
    n25136, n25137, n25138, n25139, n25140, n25141,
    n25142, n25143, n25144, n25145, n25146, n25147,
    n25148, n25149, n25150, n25151, n25152, n25153,
    n25154, n25155, n25156, n25157, n25158, n25159,
    n25160, n25161, n25162, n25163, n25164, n25165,
    n25166, n25167, n25168, n25169, n25170, n25171,
    n25172, n25173, n25174, n25175, n25176, n25177,
    n25178, n25179, n25180, n25181, n25182, n25183,
    n25184, n25185, n25186, n25187, n25188, n25189,
    n25190, n25191, n25192, n25193, n25194, n25195,
    n25196, n25197, n25198, n25199, n25200, n25201,
    n25202, n25203, n25204, n25205, n25206, n25207,
    n25208, n25209, n25210, n25211, n25212, n25213,
    n25214, n25215, n25216, n25217, n25218, n25219,
    n25220, n25221, n25222, n25223, n25224, n25225,
    n25226, n25227, n25228, n25229, n25230, n25231,
    n25232, n25233, n25234, n25235, n25236, n25237,
    n25238, n25239, n25240, n25241, n25242, n25243,
    n25244, n25245, n25246, n25247, n25248, n25249,
    n25250, n25251, n25252, n25253, n25254, n25255,
    n25256, n25257, n25258, n25259, n25260, n25261,
    n25262, n25263, n25264, n25265, n25266, n25267,
    n25268, n25269, n25270, n25271, n25272, n25273,
    n25274, n25275, n25276, n25277, n25278, n25279,
    n25280, n25281, n25282, n25283, n25284, n25285,
    n25286, n25287, n25288, n25289, n25290, n25291,
    n25292, n25293, n25294, n25295, n25296, n25297,
    n25298, n25299, n25300, n25301, n25302, n25303,
    n25304, n25305, n25306, n25307, n25308, n25309,
    n25310, n25311, n25312, n25313, n25314, n25315,
    n25316, n25317, n25318, n25319, n25320, n25321,
    n25322, n25323, n25324, n25325, n25326, n25327,
    n25328, n25329, n25330, n25331, n25332, n25333,
    n25334, n25335, n25336, n25337, n25338, n25339,
    n25340, n25341, n25342, n25343, n25344, n25345,
    n25346, n25347, n25348, n25349, n25350, n25351,
    n25352, n25353, n25354, n25355, n25356, n25357,
    n25358, n25359, n25360, n25361, n25362, n25363,
    n25364, n25365, n25366, n25367, n25368, n25369,
    n25370, n25371, n25372, n25373, n25374, n25375,
    n25376, n25377, n25378, n25379, n25380, n25381,
    n25382, n25383, n25384, n25385, n25386, n25387,
    n25388, n25389, n25390, n25391, n25392, n25393,
    n25394, n25395, n25396, n25397, n25398, n25399,
    n25400, n25401, n25402, n25403, n25404, n25405,
    n25406, n25407, n25408, n25409, n25410, n25411,
    n25412, n25413, n25414, n25415, n25416, n25417,
    n25418, n25419, n25420, n25421, n25422, n25423,
    n25424, n25425, n25426, n25427, n25428, n25429,
    n25430, n25431, n25432, n25433, n25434, n25435,
    n25436, n25437, n25438, n25439, n25440, n25441,
    n25442, n25443, n25444, n25445, n25446, n25447,
    n25448, n25449, n25450, n25451, n25452, n25453,
    n25454, n25455, n25456, n25457, n25458, n25459,
    n25460, n25461, n25462, n25463, n25464, n25465,
    n25466, n25467, n25468, n25469, n25470, n25471,
    n25472, n25473, n25474, n25475, n25476, n25477,
    n25478, n25479, n25480, n25481, n25482, n25483,
    n25484, n25485, n25486, n25487, n25488, n25489,
    n25490, n25491, n25492, n25493, n25494, n25495,
    n25496, n25497, n25498, n25499, n25500, n25501,
    n25502, n25503, n25504, n25505, n25506, n25507,
    n25508, n25509, n25510, n25511, n25512, n25513,
    n25514, n25515, n25516, n25517, n25518, n25519,
    n25520, n25521, n25522, n25523, n25524, n25525,
    n25526, n25527, n25528, n25529, n25530, n25531,
    n25532, n25533, n25534, n25535, n25536, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543,
    n25544, n25545, n25546, n25547, n25548, n25549,
    n25550, n25551, n25552, n25553, n25554, n25555,
    n25556, n25557, n25558, n25559, n25560, n25561,
    n25562, n25563, n25564, n25565, n25566, n25567,
    n25568, n25569, n25570, n25571, n25572, n25573,
    n25574, n25575, n25576, n25577, n25578, n25579,
    n25580, n25581, n25582, n25583, n25584, n25585,
    n25586, n25587, n25588, n25589, n25590, n25591,
    n25592, n25593, n25594, n25595, n25596, n25597,
    n25598, n25599, n25600, n25601, n25602, n25603,
    n25604, n25605, n25606, n25607, n25608, n25609,
    n25610, n25611, n25612, n25613, n25614, n25615,
    n25616, n25617, n25618, n25619, n25620, n25621,
    n25622, n25623, n25624, n25625, n25626, n25627,
    n25628, n25629, n25630, n25631, n25632, n25633,
    n25634, n25635, n25636, n25637, n25638, n25639,
    n25640, n25641, n25642, n25643, n25644, n25645,
    n25646, n25647, n25648, n25649, n25650, n25651,
    n25652, n25653, n25654, n25655, n25656, n25657,
    n25658, n25659, n25660, n25661, n25662, n25663,
    n25664, n25665, n25666, n25667, n25668, n25669,
    n25670, n25671, n25672, n25673, n25674, n25675,
    n25676, n25677, n25678, n25679, n25680, n25681,
    n25682, n25683, n25684, n25685, n25686, n25687,
    n25688, n25689, n25690, n25691, n25692, n25693,
    n25694, n25695, n25696, n25697, n25698, n25699,
    n25700, n25701, n25702, n25703, n25704, n25705,
    n25706, n25707, n25708, n25709, n25710, n25711,
    n25712, n25713, n25714, n25715, n25716, n25717,
    n25718, n25719, n25720, n25721, n25722, n25723,
    n25724, n25725, n25726, n25727, n25728, n25729,
    n25730, n25731, n25732, n25733, n25734, n25735,
    n25736, n25737, n25738, n25739, n25740, n25741,
    n25742, n25743, n25744, n25745, n25746, n25747,
    n25748, n25749, n25750, n25751, n25752, n25753,
    n25754, n25755, n25756, n25757, n25758, n25759,
    n25760, n25761, n25762, n25763, n25764, n25765,
    n25766, n25767, n25768, n25769, n25770, n25771,
    n25772, n25773, n25774, n25775, n25776, n25777,
    n25778, n25779, n25780, n25781, n25782, n25783,
    n25784, n25785, n25786, n25787, n25788, n25789,
    n25790, n25791, n25792, n25793, n25794, n25795,
    n25796, n25797, n25798, n25799, n25800, n25801,
    n25802, n25803, n25804, n25805, n25806, n25807,
    n25808, n25809, n25810, n25811, n25812, n25813,
    n25814, n25815, n25816, n25817, n25818, n25819,
    n25820, n25821, n25822, n25823, n25824, n25825,
    n25826, n25827, n25828, n25829, n25830, n25831,
    n25832, n25833, n25834, n25835, n25836, n25837,
    n25838, n25839, n25840, n25841, n25842, n25843,
    n25844, n25845, n25846, n25847, n25848, n25849,
    n25850, n25851, n25852, n25853, n25854, n25855,
    n25856, n25857, n25858, n25859, n25860, n25861,
    n25862, n25863, n25864, n25865, n25866, n25867,
    n25868, n25869, n25870, n25871, n25872, n25873,
    n25874, n25875, n25876, n25877, n25878, n25879,
    n25880, n25881, n25882, n25883, n25884, n25885,
    n25886, n25887, n25888, n25889, n25890, n25891,
    n25892, n25893, n25894, n25895, n25896, n25897,
    n25898, n25899, n25900, n25901, n25902, n25903,
    n25904, n25905, n25906, n25907, n25908, n25909,
    n25910, n25911, n25912, n25913, n25914, n25915,
    n25916, n25917, n25918, n25919, n25920, n25921,
    n25922, n25923, n25924, n25925, n25926, n25927,
    n25928, n25929, n25930, n25931, n25932, n25933,
    n25934, n25935, n25936, n25937, n25938, n25939,
    n25940, n25941, n25942, n25943, n25944, n25945,
    n25946, n25947, n25948, n25949, n25950, n25951,
    n25952, n25953, n25954, n25955, n25956, n25957,
    n25958, n25959, n25960, n25961, n25962, n25963,
    n25964, n25965, n25966, n25967, n25968, n25969,
    n25970, n25971, n25972, n25973, n25974, n25975,
    n25976, n25977, n25978, n25979, n25980, n25981,
    n25982, n25983, n25984, n25985, n25986, n25987,
    n25988, n25989, n25990, n25991, n25992, n25993,
    n25994, n25995, n25996, n25997, n25998, n25999,
    n26000, n26001, n26002, n26003, n26004, n26005,
    n26006, n26007, n26008, n26009, n26010, n26011,
    n26012, n26013, n26014, n26015, n26016, n26017,
    n26018, n26019, n26020, n26021, n26022, n26023,
    n26024, n26025, n26026, n26027, n26028, n26029,
    n26030, n26031, n26032, n26033, n26034, n26035,
    n26036, n26037, n26038, n26039, n26040, n26041,
    n26042, n26043, n26044, n26045, n26046, n26047,
    n26048, n26049, n26050, n26051, n26052, n26053,
    n26054, n26055, n26056, n26057, n26058, n26059,
    n26060, n26061, n26062, n26063, n26064, n26065,
    n26066, n26067, n26068, n26069, n26070, n26071,
    n26072, n26073, n26074, n26075, n26076, n26077,
    n26078, n26079, n26080, n26081, n26082, n26083,
    n26084, n26085, n26086, n26087, n26088, n26089,
    n26090, n26091, n26092, n26093, n26094, n26095,
    n26096, n26097, n26098, n26099, n26100, n26101,
    n26102, n26103, n26104, n26105, n26106, n26107,
    n26108, n26109, n26110, n26111, n26112, n26113,
    n26114, n26115, n26116, n26117, n26118, n26119,
    n26120, n26121, n26122, n26123, n26124, n26125,
    n26126, n26127, n26128, n26129, n26130, n26131,
    n26132, n26133, n26134, n26135, n26136, n26137,
    n26138, n26139, n26140, n26141, n26142, n26143,
    n26144, n26145, n26146, n26147, n26148, n26149,
    n26150, n26151, n26152, n26153, n26154, n26155,
    n26156, n26157, n26158, n26159, n26160, n26161,
    n26162, n26163, n26164, n26165, n26166, n26167,
    n26168, n26169, n26170, n26171, n26172, n26173,
    n26174, n26175, n26176, n26177, n26178, n26179,
    n26180, n26181, n26182, n26183, n26184, n26185,
    n26186, n26187, n26188, n26189, n26190, n26191,
    n26192, n26193, n26194, n26195, n26196, n26197,
    n26198, n26199, n26200, n26201, n26202, n26203,
    n26204, n26205, n26206, n26207, n26208, n26209,
    n26210, n26211, n26212, n26213, n26214, n26215,
    n26216, n26217, n26218, n26219, n26220, n26221,
    n26222, n26223, n26224, n26225, n26226, n26227,
    n26228, n26229, n26230, n26231, n26232, n26233,
    n26234, n26235, n26236, n26237, n26238, n26239,
    n26240, n26241, n26242, n26243, n26244, n26245,
    n26246, n26247, n26248, n26249, n26250, n26251,
    n26252, n26253, n26254, n26255, n26256, n26257,
    n26258, n26259, n26260, n26261, n26262, n26263,
    n26264, n26265, n26266, n26267, n26268, n26269,
    n26270, n26271, n26272, n26273, n26274, n26275,
    n26276, n26277, n26278, n26279, n26280, n26281,
    n26282, n26283, n26284, n26285, n26286, n26287,
    n26288, n26289, n26290, n26291, n26292, n26293,
    n26294, n26295, n26296, n26297, n26298, n26299,
    n26300, n26301, n26302, n26303, n26304, n26305,
    n26306, n26307, n26308, n26309, n26310, n26311,
    n26312, n26313, n26314, n26315, n26316, n26317,
    n26318, n26319, n26320, n26321, n26322, n26323,
    n26324, n26325, n26326, n26327, n26328, n26329,
    n26330, n26331, n26332, n26333, n26334, n26335,
    n26336, n26337, n26338, n26339, n26340, n26341,
    n26342, n26343, n26344, n26345, n26346, n26347,
    n26348, n26349, n26350, n26351, n26352, n26353,
    n26354, n26355, n26356, n26357, n26358, n26359,
    n26360, n26361, n26362, n26363, n26364, n26365,
    n26366, n26367, n26368, n26369, n26370, n26371,
    n26372, n26373, n26374, n26375, n26376, n26377,
    n26378, n26379, n26380, n26381, n26382, n26383,
    n26384, n26385, n26386, n26387, n26388, n26389,
    n26390, n26391, n26392, n26393, n26394, n26395,
    n26396, n26397, n26398, n26399, n26400, n26401,
    n26402, n26403, n26404, n26405, n26406, n26407,
    n26408, n26409, n26410, n26411, n26412, n26413,
    n26414, n26415, n26416, n26417, n26418, n26419,
    n26420, n26421, n26422, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26431,
    n26432, n26433, n26434, n26435, n26436, n26437,
    n26438, n26439, n26440, n26441, n26442, n26443,
    n26444, n26445, n26446, n26447, n26448, n26449,
    n26450, n26451, n26452, n26453, n26454, n26455,
    n26456, n26457, n26458, n26459, n26460, n26461,
    n26462, n26463, n26464, n26465, n26466, n26467,
    n26468, n26469, n26470, n26471, n26472, n26473,
    n26474, n26475, n26476, n26477, n26478, n26479,
    n26480, n26481, n26482, n26483, n26484, n26485,
    n26486, n26487, n26488, n26489, n26490, n26491,
    n26492, n26493, n26494, n26495, n26496, n26497,
    n26498, n26499, n26500, n26501, n26502, n26503,
    n26504, n26505, n26506, n26507, n26508, n26509,
    n26510, n26511, n26512, n26513, n26514, n26515,
    n26516, n26517, n26518, n26519, n26520, n26521,
    n26522, n26523, n26524, n26525, n26526, n26527,
    n26528, n26529, n26530, n26531, n26532, n26533,
    n26534, n26535, n26536, n26537, n26538, n26539,
    n26540, n26541, n26542, n26543, n26544, n26545,
    n26546, n26547, n26548, n26549, n26550, n26551,
    n26552, n26553, n26554, n26555, n26556, n26557,
    n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26571, n26572, n26573, n26574, n26575,
    n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587,
    n26588, n26589, n26590, n26591, n26592, n26593,
    n26594, n26595, n26596, n26597, n26598, n26599,
    n26600, n26601, n26602, n26603, n26604, n26605,
    n26606, n26607, n26608, n26609, n26610, n26611,
    n26612, n26613, n26614, n26615, n26616, n26617,
    n26618, n26619, n26620, n26621, n26622, n26623,
    n26624, n26625, n26626, n26627, n26628, n26629,
    n26630, n26631, n26632, n26633, n26634, n26635,
    n26636, n26637, n26638, n26639, n26640, n26641,
    n26642, n26643, n26644, n26645, n26646, n26647,
    n26648, n26649, n26650, n26651, n26652, n26653,
    n26654, n26655, n26656, n26657, n26658, n26659,
    n26660, n26661, n26662, n26663, n26664, n26665,
    n26666, n26667, n26668, n26669, n26670, n26671,
    n26672, n26673, n26674, n26675, n26676, n26677,
    n26678, n26679, n26680, n26681, n26682, n26683,
    n26684, n26685, n26686, n26687, n26688, n26689,
    n26690, n26691, n26692, n26693, n26694, n26695,
    n26696, n26697, n26698, n26699, n26700, n26701,
    n26702, n26703, n26704, n26705, n26706, n26707,
    n26708, n26709, n26710, n26711, n26712, n26713,
    n26714, n26715, n26716, n26717, n26718, n26719,
    n26720, n26721, n26722, n26723, n26724, n26725,
    n26726, n26727, n26728, n26729, n26730, n26731,
    n26732, n26733, n26734, n26735, n26736, n26737,
    n26738, n26739, n26740, n26741, n26742, n26743,
    n26744, n26745, n26746, n26747, n26748, n26749,
    n26750, n26751, n26752, n26753, n26754, n26755,
    n26756, n26757, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767,
    n26768, n26769, n26770, n26771, n26772, n26773,
    n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785,
    n26786, n26787, n26788, n26789, n26790, n26791,
    n26792, n26793, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26802, n26803,
    n26804, n26805, n26806, n26807, n26808, n26809,
    n26810, n26811, n26812, n26813, n26814, n26815,
    n26816, n26817, n26818, n26819, n26820, n26821,
    n26822, n26823, n26824, n26825, n26826, n26827,
    n26828, n26829, n26830, n26831, n26832, n26833,
    n26834, n26835, n26836, n26837, n26838, n26839,
    n26840, n26841, n26842, n26843, n26844, n26845,
    n26846, n26847, n26848, n26849, n26850, n26851,
    n26852, n26853, n26854, n26855, n26856, n26857,
    n26858, n26859, n26860, n26861, n26862, n26863,
    n26864, n26865, n26866, n26867, n26868, n26869,
    n26870, n26871, n26872, n26873, n26874, n26875,
    n26876, n26877, n26878, n26879, n26880, n26881,
    n26882, n26883, n26884, n26885, n26886, n26887,
    n26888, n26889, n26890, n26891, n26892, n26893,
    n26894, n26895, n26896, n26897, n26898, n26899,
    n26900, n26901, n26902, n26903, n26904, n26905,
    n26906, n26907, n26908, n26909, n26910, n26911,
    n26912, n26913, n26914, n26915, n26916, n26917,
    n26918, n26919, n26920, n26921, n26922, n26923,
    n26924, n26925, n26926, n26927, n26928, n26929,
    n26930, n26931, n26932, n26933, n26934, n26935,
    n26936, n26937, n26938, n26939, n26940, n26941,
    n26942, n26943, n26944, n26945, n26946, n26947,
    n26948, n26949, n26950, n26951, n26952, n26953,
    n26954, n26955, n26956, n26957, n26958, n26959,
    n26960, n26961, n26962, n26963, n26964, n26965,
    n26966, n26967, n26968, n26969, n26970, n26971,
    n26972, n26973, n26974, n26975, n26976, n26977,
    n26978, n26979, n26980, n26981, n26982, n26983,
    n26984, n26985, n26986, n26987, n26988, n26989,
    n26990, n26991, n26992, n26993, n26994, n26995,
    n26996, n26997, n26998, n26999, n27000, n27001,
    n27002, n27003, n27004, n27005, n27006, n27007,
    n27008, n27009, n27010, n27011, n27012, n27013,
    n27014, n27015, n27016, n27017, n27018, n27019,
    n27020, n27021, n27022, n27023, n27024, n27025,
    n27026, n27027, n27028, n27029, n27030, n27031,
    n27032, n27033, n27034, n27035, n27036, n27037,
    n27038, n27039, n27040, n27041, n27042, n27043,
    n27044, n27045, n27046, n27047, n27048, n27049,
    n27050, n27051, n27052, n27053, n27054, n27055,
    n27056, n27057, n27058, n27059, n27060, n27061,
    n27062, n27063, n27064, n27065, n27066, n27067,
    n27068, n27069, n27070, n27071, n27072, n27073,
    n27074, n27075, n27076, n27077, n27078, n27079,
    n27080, n27081, n27082, n27083, n27084, n27085,
    n27086, n27087, n27088, n27089, n27090, n27091,
    n27092, n27093, n27094, n27095, n27096, n27097,
    n27098, n27099, n27100, n27101, n27102, n27103,
    n27104, n27105, n27106, n27107, n27108, n27109,
    n27110, n27111, n27112, n27113, n27114, n27115,
    n27116, n27117, n27118, n27119, n27120, n27121,
    n27122, n27123, n27124, n27125, n27126, n27127,
    n27128, n27129, n27130, n27131, n27132, n27133,
    n27134, n27135, n27136, n27137, n27138, n27139,
    n27140, n27141, n27142, n27143, n27144, n27145,
    n27146, n27147, n27148, n27149, n27150, n27151,
    n27152, n27153, n27154, n27155, n27156, n27157,
    n27158, n27159, n27160, n27161, n27162, n27163,
    n27164, n27165, n27166, n27167, n27168, n27169,
    n27170, n27171, n27172, n27173, n27174, n27175,
    n27176, n27177, n27178, n27179, n27180, n27181,
    n27182, n27183, n27184, n27185, n27186, n27187,
    n27188, n27189, n27190, n27191, n27192, n27193,
    n27194, n27195, n27196, n27197, n27198, n27199,
    n27200, n27201, n27202, n27203, n27204, n27205,
    n27206, n27207, n27208, n27209, n27210, n27211,
    n27212, n27213, n27214, n27215, n27216, n27217,
    n27218, n27219, n27220, n27221, n27222, n27223,
    n27224, n27225, n27226, n27227, n27228, n27229,
    n27230, n27231, n27232, n27233, n27234, n27235,
    n27236, n27237, n27238, n27239, n27240, n27241,
    n27242, n27243, n27244, n27245, n27246, n27247,
    n27248, n27249, n27250, n27251, n27252, n27253,
    n27254, n27255, n27256, n27257, n27258, n27259,
    n27260, n27261, n27262, n27263, n27264, n27265,
    n27266, n27267, n27268, n27269, n27270, n27271,
    n27272, n27273, n27274, n27275, n27276, n27277,
    n27278, n27279, n27280, n27281, n27282, n27283,
    n27284, n27285, n27286, n27287, n27288, n27289,
    n27290, n27291, n27292, n27293, n27294, n27295,
    n27296, n27297, n27298, n27299, n27300, n27301,
    n27302, n27303, n27304, n27305, n27306, n27307,
    n27308, n27309, n27310, n27311, n27312, n27313,
    n27314, n27315, n27316, n27317, n27318, n27319,
    n27320, n27321, n27322, n27323, n27324, n27325,
    n27326, n27327, n27328, n27329, n27330, n27331,
    n27332, n27333, n27334, n27335, n27336, n27337,
    n27338, n27339, n27340, n27341, n27342, n27343,
    n27344, n27345, n27346, n27347, n27348, n27349,
    n27350, n27351, n27352, n27353, n27354, n27355,
    n27356, n27357, n27358, n27359, n27360, n27361,
    n27362, n27363, n27364, n27365, n27366, n27367,
    n27368, n27369, n27370, n27371, n27372, n27373,
    n27374, n27375, n27376, n27377, n27378, n27379,
    n27380, n27381, n27382, n27383, n27384, n27385,
    n27386, n27387, n27388, n27389, n27390, n27391,
    n27392, n27393, n27394, n27395, n27396, n27397,
    n27398, n27399, n27400, n27401, n27402, n27403,
    n27404, n27405, n27406, n27407, n27408, n27409,
    n27410, n27411, n27412, n27413, n27414, n27415,
    n27416, n27417, n27418, n27419, n27420, n27421,
    n27422, n27423, n27424, n27425, n27426, n27427,
    n27428, n27429, n27430, n27431, n27432, n27433,
    n27434, n27435, n27436, n27437, n27438, n27439,
    n27440, n27441, n27442, n27443, n27444, n27445,
    n27446, n27447, n27448, n27449, n27450, n27451,
    n27452, n27453, n27454, n27455, n27456, n27457,
    n27458, n27459, n27460, n27461, n27462, n27463,
    n27464, n27465, n27466, n27467, n27468, n27469,
    n27470, n27471, n27472, n27473, n27474, n27475,
    n27476, n27477, n27478, n27479, n27480, n27481,
    n27482, n27483, n27484, n27485, n27486, n27487,
    n27488, n27489, n27490, n27491, n27492, n27493,
    n27494, n27495, n27496, n27497, n27498, n27499,
    n27500, n27501, n27502, n27503, n27504, n27505,
    n27506, n27507, n27508, n27509, n27510, n27511,
    n27512, n27513, n27514, n27515, n27516, n27517,
    n27518, n27519, n27520, n27521, n27522, n27523,
    n27524, n27525, n27526, n27527, n27528, n27529,
    n27530, n27531, n27532, n27533, n27534, n27535,
    n27536, n27537, n27538, n27539, n27540, n27541,
    n27542, n27543, n27544, n27545, n27546, n27547,
    n27548, n27549, n27550, n27551, n27552, n27553,
    n27554, n27555, n27556, n27557, n27558, n27559,
    n27560, n27561, n27562, n27563, n27564, n27565,
    n27566, n27567, n27568, n27569, n27570, n27571,
    n27572, n27573, n27574, n27575, n27576, n27577,
    n27578, n27579, n27580, n27581, n27582, n27583,
    n27584, n27585, n27586, n27587, n27588, n27589,
    n27590, n27591, n27592, n27593, n27594, n27595,
    n27596, n27597, n27598, n27599, n27600, n27601,
    n27602, n27603, n27604, n27605, n27606, n27607,
    n27608, n27609, n27610, n27611, n27612, n27613,
    n27614, n27615, n27616, n27617, n27618, n27619,
    n27620, n27621, n27622, n27623, n27624, n27625,
    n27626, n27627, n27628, n27629, n27630, n27631,
    n27632, n27633, n27634, n27635, n27636, n27637,
    n27638, n27639, n27640, n27641, n27642, n27643,
    n27644, n27645, n27646, n27647, n27648, n27649,
    n27650, n27651, n27652, n27653, n27654, n27655,
    n27656, n27657, n27658, n27659, n27660, n27661,
    n27662, n27663, n27664, n27665, n27666, n27667,
    n27668, n27669, n27670, n27671, n27672, n27673,
    n27674, n27675, n27676, n27677, n27678, n27679,
    n27680, n27681, n27682, n27683, n27684, n27685,
    n27686, n27687, n27688, n27689, n27690, n27691,
    n27692, n27693, n27694, n27695, n27696, n27697,
    n27698, n27699, n27700, n27701, n27702, n27703,
    n27704, n27705, n27706, n27707, n27708, n27709,
    n27710, n27711, n27712, n27713, n27714, n27715,
    n27716, n27717, n27718, n27719, n27720, n27721,
    n27722, n27723, n27724, n27725, n27726, n27727,
    n27728, n27729, n27730, n27731, n27732, n27733,
    n27734, n27735, n27736, n27737, n27738, n27739,
    n27740, n27741, n27742, n27743, n27744, n27745,
    n27746, n27747, n27748, n27749, n27750, n27751,
    n27752, n27753, n27754, n27755, n27756, n27757,
    n27758, n27759, n27760, n27761, n27762, n27763,
    n27764, n27765, n27766, n27767, n27768, n27769,
    n27770, n27771, n27772, n27773, n27774, n27775,
    n27776, n27777, n27778, n27779, n27780, n27781,
    n27782, n27783, n27784, n27785, n27786, n27787,
    n27788, n27789, n27790, n27791, n27792, n27793,
    n27794, n27795, n27796, n27797, n27798, n27799,
    n27800, n27801, n27802, n27803, n27804, n27805,
    n27806, n27807, n27808, n27809, n27810, n27811,
    n27812, n27813, n27814, n27815, n27816, n27817,
    n27818, n27819, n27820, n27821, n27822, n27823,
    n27824, n27825, n27826, n27827, n27828, n27829,
    n27830, n27831, n27832, n27833, n27834, n27835,
    n27836, n27837, n27838, n27839, n27840, n27841,
    n27842, n27843, n27844, n27845, n27846, n27847,
    n27848, n27849, n27850, n27851, n27852, n27853,
    n27854, n27855, n27856, n27857, n27858, n27859,
    n27860, n27861, n27862, n27863, n27864, n27865,
    n27866, n27867, n27868, n27869, n27870, n27871,
    n27872, n27873, n27874, n27875, n27876, n27877,
    n27878, n27879, n27880, n27881, n27882, n27883,
    n27884, n27885, n27886, n27887, n27888, n27889,
    n27890, n27891, n27892, n27893, n27894, n27895,
    n27896, n27897, n27898, n27899, n27900, n27901,
    n27902, n27903, n27904, n27905, n27906, n27907,
    n27908, n27909, n27910, n27911, n27912, n27913,
    n27914, n27915, n27916, n27917, n27918, n27919,
    n27920, n27921, n27922, n27923, n27924, n27925,
    n27926, n27927, n27928, n27929, n27930, n27931,
    n27932, n27933, n27934, n27935, n27936, n27937,
    n27938, n27939, n27940, n27941, n27942, n27943,
    n27944, n27945, n27946, n27947, n27948, n27949,
    n27950, n27951, n27952, n27953, n27954, n27955,
    n27956, n27957, n27958, n27959, n27960, n27961,
    n27962, n27963, n27964, n27965, n27966, n27967,
    n27968, n27969, n27970, n27971, n27972, n27973,
    n27974, n27975, n27976, n27977, n27978, n27979,
    n27980, n27981, n27982, n27983, n27984, n27985,
    n27986, n27987, n27988, n27989, n27990, n27991,
    n27992, n27993, n27994, n27995, n27996, n27997,
    n27998, n27999, n28000, n28001, n28002, n28003,
    n28004, n28005, n28006, n28007, n28008, n28009,
    n28010, n28011, n28012, n28013, n28014, n28015,
    n28016, n28017, n28018, n28019, n28020, n28021,
    n28022, n28023, n28024, n28025, n28026, n28027,
    n28028, n28029, n28030, n28031, n28032, n28033,
    n28034, n28035, n28036, n28037, n28038, n28039,
    n28040, n28041, n28042, n28043, n28044, n28045,
    n28046, n28047, n28048, n28049, n28050, n28051,
    n28052, n28053, n28054, n28055, n28056, n28057,
    n28058, n28059, n28060, n28061, n28062, n28063,
    n28064, n28065, n28066, n28067, n28068, n28069,
    n28070, n28071, n28072, n28073, n28074, n28075,
    n28076, n28077, n28078, n28079, n28080, n28081,
    n28082, n28083, n28084, n28085, n28086, n28087,
    n28088, n28089, n28090, n28091, n28092, n28093,
    n28094, n28095, n28096, n28097, n28098, n28099,
    n28100, n28101, n28102, n28103, n28104, n28105,
    n28106, n28107, n28108, n28109, n28110, n28111,
    n28112, n28113, n28114, n28115, n28116, n28117,
    n28118, n28119, n28120, n28121, n28122, n28123,
    n28124, n28125, n28126, n28127, n28128, n28129,
    n28130, n28131, n28132, n28133, n28134, n28135,
    n28136, n28137, n28138, n28139, n28140, n28141,
    n28142, n28143, n28144, n28145, n28146, n28147,
    n28148, n28149, n28150, n28151, n28152, n28153,
    n28154, n28155, n28156, n28157, n28158, n28159,
    n28160, n28161, n28162, n28163, n28164, n28165,
    n28166, n28167, n28168, n28169, n28170, n28171,
    n28172, n28173, n28174, n28175, n28176, n28177,
    n28178, n28179, n28180, n28181, n28182, n28183,
    n28184, n28185, n28186, n28187, n28188, n28189,
    n28190, n28191, n28192, n28193, n28194, n28195,
    n28196, n28197, n28198, n28199, n28200, n28201,
    n28202, n28203, n28204, n28205, n28206, n28207,
    n28208, n28209, n28210, n28211, n28212, n28213,
    n28214, n28215, n28216, n28217, n28218, n28219,
    n28220, n28221, n28222, n28223, n28224, n28225,
    n28226, n28227, n28228, n28229, n28230, n28231,
    n28232, n28233, n28234, n28235, n28236, n28237,
    n28238, n28239, n28240, n28241, n28242, n28243,
    n28244, n28245, n28246, n28247, n28248, n28249,
    n28250, n28251, n28252, n28253, n28254, n28255,
    n28256, n28257, n28258, n28259, n28260, n28261,
    n28262, n28263, n28264, n28265, n28266, n28267,
    n28268, n28269, n28270, n28271, n28272, n28273,
    n28274, n28275, n28276, n28277, n28278, n28279,
    n28280, n28281, n28282, n28283, n28284, n28285,
    n28286, n28287, n28288, n28289, n28290, n28291,
    n28292, n28293, n28294, n28295, n28296, n28297,
    n28298, n28299, n28300, n28301, n28302, n28303,
    n28304, n28305, n28306, n28307, n28308, n28309,
    n28310, n28311, n28312, n28313, n28314, n28315,
    n28316, n28317, n28318, n28319, n28320, n28321,
    n28322, n28323, n28324, n28325, n28326, n28327,
    n28328, n28329, n28330, n28331, n28332, n28333,
    n28334, n28335, n28336, n28337, n28338, n28339,
    n28340, n28341, n28342, n28343, n28344, n28345,
    n28346, n28347, n28348, n28349, n28350, n28351,
    n28352, n28353, n28354, n28355, n28356, n28357,
    n28358, n28359, n28360, n28361, n28362, n28363,
    n28364, n28365, n28366, n28367, n28368, n28369,
    n28370, n28371, n28372, n28373, n28374, n28375,
    n28376, n28377, n28378, n28379, n28380, n28381,
    n28382, n28383, n28384, n28385, n28386, n28387,
    n28388, n28389, n28390, n28391, n28392, n28393,
    n28394, n28395, n28396, n28397, n28398, n28399,
    n28400, n28401, n28402, n28403, n28404, n28405,
    n28406, n28407, n28408, n28409, n28410, n28411,
    n28412, n28413, n28414, n28415, n28416, n28417,
    n28418, n28419, n28420, n28421, n28422, n28423,
    n28424, n28425, n28426, n28427, n28428, n28429,
    n28430, n28431, n28432, n28433, n28434, n28435,
    n28436, n28437, n28438, n28439, n28440, n28441,
    n28442, n28443, n28444, n28445, n28446, n28447,
    n28448, n28449, n28450, n28451, n28452, n28453,
    n28454, n28455, n28456, n28457, n28458, n28459,
    n28460, n28461, n28462, n28463, n28464, n28465,
    n28466, n28467, n28468, n28469, n28470, n28471,
    n28472, n28473, n28474, n28475, n28476, n28477,
    n28478, n28479, n28480, n28481, n28482, n28483,
    n28484, n28485, n28486, n28487, n28488, n28489,
    n28490, n28491, n28492, n28493, n28494, n28495,
    n28496, n28497, n28498, n28499, n28500, n28501,
    n28502, n28503, n28504, n28505, n28506, n28507,
    n28508, n28509, n28510, n28511, n28512, n28513,
    n28514, n28515, n28516, n28517, n28518, n28519,
    n28520, n28521, n28522, n28523, n28524, n28525,
    n28526, n28527, n28528, n28529, n28530, n28531,
    n28532, n28533, n28534, n28535, n28536, n28537,
    n28538, n28539, n28540, n28541, n28542, n28543,
    n28544, n28545, n28546, n28547, n28548, n28549,
    n28550, n28551, n28552, n28553, n28554, n28555,
    n28556, n28557, n28558, n28559, n28560, n28561,
    n28562, n28563, n28564, n28565, n28566, n28567,
    n28568, n28569, n28570, n28571, n28572, n28573,
    n28574, n28575, n28576, n28577, n28578, n28579,
    n28580, n28581, n28582, n28583, n28584, n28585,
    n28586, n28587, n28588, n28589, n28590, n28591,
    n28592, n28593, n28594, n28595, n28596, n28597,
    n28598, n28599, n28600, n28601, n28602, n28603,
    n28604, n28605, n28606, n28607, n28608, n28609,
    n28610, n28611, n28612, n28613, n28614, n28615,
    n28616, n28617, n28618, n28619, n28620, n28621,
    n28622, n28623, n28624, n28625, n28626, n28627,
    n28628, n28629, n28630, n28631, n28632, n28633,
    n28634, n28635, n28636, n28637, n28638, n28639,
    n28640, n28641, n28642, n28643, n28644, n28645,
    n28646, n28647, n28648, n28649, n28650, n28651,
    n28652, n28653, n28654, n28655, n28656, n28657,
    n28658, n28659, n28660, n28661, n28662, n28663,
    n28664, n28665, n28666, n28667, n28668, n28669,
    n28670, n28671, n28672, n28673, n28674, n28675,
    n28676, n28677, n28678, n28679, n28680, n28681,
    n28682, n28683, n28684, n28685, n28686, n28687,
    n28688, n28689, n28690, n28691, n28692, n28693,
    n28694, n28695, n28696, n28697, n28698, n28699,
    n28700, n28701, n28702, n28703, n28704, n28705,
    n28706, n28707, n28708, n28709, n28710, n28711,
    n28712, n28713, n28714, n28715, n28716, n28717,
    n28718, n28719, n28720, n28721, n28722, n28723,
    n28724, n28725, n28726, n28727, n28728, n28729,
    n28730, n28731, n28732, n28733, n28734, n28735,
    n28736, n28737, n28738, n28739, n28740, n28741,
    n28742, n28743, n28744, n28745, n28746, n28747,
    n28748, n28749, n28750, n28751, n28752, n28753,
    n28754, n28755, n28756, n28757, n28758, n28759,
    n28760, n28761, n28762, n28763, n28764, n28765,
    n28766, n28767, n28768, n28769, n28770, n28771,
    n28772, n28773, n28774, n28775, n28776, n28777,
    n28778, n28779, n28780, n28781, n28782, n28783,
    n28784, n28785, n28786, n28787, n28788, n28789,
    n28790, n28791, n28792, n28793, n28794, n28795,
    n28796, n28797, n28798, n28799, n28800, n28801,
    n28802, n28803, n28804, n28805, n28806, n28807,
    n28808, n28809, n28810, n28811, n28812, n28813,
    n28814, n28815, n28816, n28817, n28818, n28819,
    n28820, n28821, n28822, n28823, n28824, n28825,
    n28826, n28827, n28828, n28829, n28830, n28831,
    n28832, n28833, n28834, n28835, n28836, n28837,
    n28838, n28839, n28840, n28841, n28842, n28843,
    n28844, n28845, n28846, n28847, n28848, n28849,
    n28850, n28851, n28852, n28853, n28854, n28855,
    n28856, n28857, n28858, n28859, n28860, n28861,
    n28862, n28863, n28864, n28865, n28866, n28867,
    n28868, n28869, n28870, n28871, n28872, n28873,
    n28874, n28875, n28876, n28877, n28878, n28879,
    n28880, n28881, n28882, n28883, n28884, n28885,
    n28886, n28887, n28888, n28889, n28890, n28891,
    n28892, n28893, n28894, n28895, n28896, n28897,
    n28898, n28899, n28900, n28901, n28902, n28903,
    n28904, n28905, n28906, n28907, n28908, n28909,
    n28910, n28911, n28912, n28913, n28914, n28915,
    n28916, n28917, n28918, n28919, n28920, n28921,
    n28922, n28923, n28924, n28925, n28926, n28927,
    n28928, n28929, n28930, n28931, n28932, n28933,
    n28934, n28935, n28936, n28937, n28938, n28939,
    n28940, n28941, n28942, n28943, n28944, n28945,
    n28946, n28947, n28948, n28949, n28950, n28951,
    n28952, n28953, n28954, n28955, n28956, n28957,
    n28958, n28959, n28960, n28961, n28962, n28963,
    n28964, n28965, n28966, n28967, n28968, n28969,
    n28970, n28971, n28972, n28973, n28974, n28975,
    n28976, n28977, n28978, n28979, n28980, n28981,
    n28982, n28983, n28984, n28985, n28986, n28987,
    n28988, n28989, n28990, n28991, n28992, n28993,
    n28994, n28995, n28996, n28997, n28998, n28999,
    n29000, n29001, n29002, n29003, n29004, n29005,
    n29006, n29007, n29008, n29009, n29010, n29011,
    n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023,
    n29024, n29025, n29026, n29027, n29028, n29029,
    n29030, n29031, n29032, n29033, n29034, n29035,
    n29036, n29037, n29038, n29039, n29040, n29041,
    n29042, n29043, n29044, n29045, n29046, n29047,
    n29048, n29049, n29050, n29051, n29052, n29053,
    n29054, n29055, n29056, n29057, n29058, n29059,
    n29060, n29061, n29062, n29063, n29064, n29065,
    n29066, n29067, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077,
    n29078, n29079, n29080, n29081, n29082, n29083,
    n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095,
    n29096, n29097, n29098, n29099, n29100, n29101,
    n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113,
    n29114, n29115, n29116, n29117, n29118, n29119,
    n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131,
    n29132, n29133, n29134, n29135, n29136, n29137,
    n29138, n29139, n29140, n29141, n29142, n29143,
    n29144, n29145, n29146, n29147, n29148, n29149,
    n29150, n29151, n29152, n29153, n29154, n29155,
    n29156, n29157, n29158, n29159, n29160, n29161,
    n29162, n29163, n29164, n29165, n29166, n29167,
    n29168, n29169, n29170, n29171, n29172, n29173,
    n29174, n29175, n29176, n29177, n29178, n29179,
    n29180, n29181, n29182, n29183, n29184, n29185,
    n29186, n29187, n29188, n29189, n29190, n29191,
    n29192, n29193, n29194, n29195, n29196, n29197,
    n29198, n29199, n29200, n29201, n29202, n29203,
    n29204, n29205, n29206, n29207, n29208, n29209,
    n29210, n29211, n29212, n29213, n29214, n29215,
    n29216, n29217, n29218, n29219, n29220, n29221,
    n29222, n29223, n29224, n29225, n29226, n29227,
    n29228, n29229, n29230, n29231, n29232, n29233,
    n29234, n29235, n29236, n29237, n29238, n29239,
    n29240, n29241, n29242, n29243, n29244, n29245,
    n29246, n29247, n29248, n29249, n29250, n29251,
    n29252, n29253, n29254, n29255, n29256, n29257,
    n29258, n29259, n29260, n29261, n29262, n29263,
    n29264, n29265, n29266, n29267, n29268, n29269,
    n29270, n29271, n29272, n29273, n29274, n29275,
    n29276, n29277, n29278, n29279, n29280, n29281,
    n29282, n29283, n29284, n29285, n29286, n29287,
    n29288, n29289, n29290, n29291, n29292, n29293,
    n29294, n29295, n29296, n29297, n29298, n29299,
    n29300, n29301, n29302, n29303, n29304, n29305,
    n29306, n29307, n29308, n29309, n29310, n29311,
    n29312, n29313, n29314, n29315, n29316, n29317,
    n29318, n29319, n29320, n29321, n29322, n29323,
    n29324, n29325, n29326, n29327, n29328, n29329,
    n29330, n29331, n29332, n29333, n29334, n29335,
    n29336, n29337, n29338, n29339, n29340, n29341,
    n29342, n29343, n29344, n29345, n29346, n29347,
    n29348, n29349, n29350, n29351, n29352, n29353,
    n29354, n29355, n29356, n29357, n29358, n29359,
    n29360, n29361, n29362, n29363, n29364, n29365,
    n29366, n29367, n29368, n29369, n29370, n29371,
    n29372, n29373, n29374, n29375, n29376, n29377,
    n29378, n29379, n29380, n29381, n29382, n29383,
    n29384, n29385, n29386, n29387, n29388, n29389,
    n29390, n29391, n29392, n29393, n29394, n29395,
    n29396, n29397, n29398, n29399, n29400, n29401,
    n29402, n29403, n29404, n29405, n29406, n29407,
    n29408, n29409, n29410, n29411, n29412, n29413,
    n29414, n29415, n29416, n29417, n29418, n29419,
    n29420, n29421, n29422, n29423, n29424, n29425,
    n29426, n29427, n29428, n29429, n29430, n29431,
    n29432, n29433, n29434, n29435, n29436, n29437,
    n29438, n29439, n29440, n29441, n29442, n29443,
    n29444, n29445, n29446, n29447, n29448, n29449,
    n29450, n29451, n29452, n29453, n29454, n29455,
    n29456, n29457, n29458, n29459, n29460, n29461,
    n29462, n29463, n29464, n29465, n29466, n29467,
    n29468, n29469, n29470, n29471, n29472, n29473,
    n29474, n29475, n29476, n29477, n29478, n29479,
    n29480, n29481, n29482, n29483, n29484, n29485,
    n29486, n29487, n29488, n29489, n29490, n29491,
    n29492, n29493, n29494, n29495, n29496, n29497,
    n29498, n29499, n29500, n29501, n29502, n29503,
    n29504, n29505, n29506, n29507, n29508, n29509,
    n29510, n29511, n29512, n29513, n29514, n29515,
    n29516, n29517, n29518, n29519, n29520, n29521,
    n29522, n29523, n29524, n29525, n29526, n29527,
    n29528, n29529, n29530, n29531, n29532, n29533,
    n29534, n29535, n29536, n29537, n29538, n29539,
    n29540, n29541, n29542, n29543, n29544, n29545,
    n29546, n29547, n29548, n29549, n29550, n29551,
    n29552, n29553, n29554, n29555, n29556, n29557,
    n29558, n29559, n29560, n29561, n29562, n29563,
    n29564, n29565, n29566, n29567, n29568, n29569,
    n29570, n29571, n29572, n29573, n29574, n29575,
    n29576, n29577, n29578, n29579, n29580, n29581,
    n29582, n29583, n29584, n29585, n29586, n29587,
    n29588, n29589, n29590, n29591, n29592, n29593,
    n29594, n29595, n29596, n29597, n29598, n29599,
    n29600, n29601, n29602, n29603, n29604, n29605,
    n29606, n29607, n29608, n29609, n29610, n29611,
    n29612, n29613, n29614, n29615, n29616, n29617,
    n29618, n29619, n29620, n29621, n29622, n29623,
    n29624, n29625, n29626, n29627, n29628, n29629,
    n29630, n29631, n29632, n29633, n29634, n29635,
    n29636, n29637, n29638, n29639, n29640, n29641,
    n29642, n29643, n29644, n29645, n29646, n29647,
    n29648, n29649, n29650, n29651, n29652, n29653,
    n29654, n29655, n29656, n29657, n29658, n29659,
    n29660, n29661, n29662, n29663, n29664, n29665,
    n29666, n29667, n29668, n29669, n29670, n29671,
    n29672, n29673, n29674, n29675, n29676, n29677,
    n29678, n29679, n29680, n29681, n29682, n29683,
    n29684, n29685, n29686, n29687, n29688, n29689,
    n29690, n29691, n29692, n29693, n29694, n29695,
    n29696, n29697, n29698, n29699, n29700, n29701,
    n29702, n29703, n29704, n29705, n29706, n29707,
    n29708, n29709, n29710, n29711, n29712, n29713,
    n29714, n29715, n29716, n29717, n29718, n29719,
    n29720, n29721, n29722, n29723, n29724, n29725,
    n29726, n29727, n29728, n29729, n29730, n29731,
    n29732, n29733, n29734, n29735, n29736, n29737,
    n29738, n29739, n29740, n29741, n29742, n29743,
    n29744, n29745, n29746, n29747, n29748, n29749,
    n29750, n29751, n29752, n29753, n29754, n29755,
    n29756, n29757, n29758, n29759, n29760, n29761,
    n29762, n29763, n29764, n29765, n29766, n29767,
    n29768, n29769, n29770, n29771, n29772, n29773,
    n29774, n29775, n29776, n29777, n29778, n29779,
    n29780, n29781, n29782, n29783, n29784, n29785,
    n29786, n29787, n29788, n29789, n29790, n29791,
    n29792, n29793, n29794, n29795, n29796, n29797,
    n29798, n29799, n29800, n29801, n29802, n29803,
    n29804, n29805, n29806, n29807, n29808, n29809,
    n29810, n29811, n29812, n29813, n29814, n29815,
    n29816, n29817, n29818, n29819, n29820, n29821,
    n29822, n29823, n29824, n29825, n29826, n29827,
    n29828, n29829, n29830, n29831, n29832, n29833,
    n29834, n29835, n29836, n29837, n29838, n29839,
    n29840, n29841, n29842, n29843, n29844, n29845,
    n29846, n29847, n29848, n29849, n29850, n29851,
    n29852, n29853, n29854, n29855, n29856, n29857,
    n29858, n29859, n29860, n29861, n29862, n29863,
    n29864, n29865, n29866, n29867, n29868, n29869,
    n29870, n29871, n29872, n29873, n29874, n29875,
    n29876, n29877, n29878, n29879, n29880, n29881,
    n29882, n29883, n29884, n29885, n29886, n29887,
    n29888, n29889, n29890, n29891, n29892, n29893,
    n29894, n29895, n29896, n29897, n29898, n29899,
    n29900, n29901, n29902, n29903, n29904, n29905,
    n29906, n29907, n29908, n29909, n29910, n29911,
    n29912, n29913, n29914, n29915, n29916, n29917,
    n29918, n29919, n29920, n29921, n29922, n29923,
    n29924, n29925, n29926, n29927, n29928, n29929,
    n29930, n29931, n29932, n29933, n29934, n29935,
    n29936, n29937, n29938, n29939, n29940, n29941,
    n29942, n29943, n29944, n29945, n29946, n29947,
    n29948, n29949, n29950, n29951, n29952, n29953,
    n29954, n29955, n29956, n29957, n29958, n29959,
    n29960, n29961, n29962, n29963, n29964, n29965,
    n29966, n29967, n29968, n29969, n29970, n29971,
    n29972, n29973, n29974, n29975, n29976, n29977,
    n29978, n29979, n29980, n29981, n29982, n29983,
    n29984, n29985, n29986, n29987, n29988, n29989,
    n29990, n29991, n29992, n29993, n29994, n29995,
    n29996, n29997, n29998, n29999, n30000, n30001,
    n30002, n30003, n30004, n30005, n30006, n30007,
    n30008, n30009, n30010, n30011, n30012, n30013,
    n30014, n30015, n30016, n30017, n30018, n30019,
    n30020, n30021, n30022, n30023, n30024, n30025,
    n30026, n30027, n30028, n30029, n30030, n30031,
    n30032, n30033, n30034, n30035, n30036, n30037,
    n30038, n30039, n30040, n30041, n30042, n30043,
    n30044, n30045, n30046, n30047, n30048, n30049,
    n30050, n30051, n30052, n30053, n30054, n30055,
    n30056, n30057, n30058, n30059, n30060, n30061,
    n30062, n30063, n30064, n30065, n30066, n30067,
    n30068, n30069, n30070, n30071, n30072, n30073,
    n30074, n30075, n30076, n30077, n30078, n30079,
    n30080, n30081, n30082, n30083, n30084, n30085,
    n30086, n30087, n30088, n30089, n30090, n30091,
    n30092, n30093, n30094, n30095, n30096, n30097,
    n30098, n30099, n30100, n30101, n30102, n30103,
    n30104, n30105, n30106, n30107, n30108, n30109,
    n30110, n30111, n30112, n30113, n30114, n30115,
    n30116, n30117, n30118, n30119, n30120, n30121,
    n30122, n30123, n30124, n30125, n30126, n30127,
    n30128, n30129, n30130, n30131, n30132, n30133,
    n30134, n30135, n30136, n30137, n30138, n30139,
    n30140, n30141, n30142, n30143, n30144, n30145,
    n30146, n30147, n30148, n30149, n30150, n30151,
    n30152, n30153, n30154, n30155, n30156, n30157,
    n30158, n30159, n30160, n30161, n30162, n30163,
    n30164, n30165, n30166, n30167, n30168, n30169,
    n30170, n30171, n30172, n30173, n30174, n30175,
    n30176, n30177, n30178, n30179, n30180, n30181,
    n30182, n30183, n30184, n30185, n30186, n30187,
    n30188, n30189, n30190, n30191, n30192, n30193,
    n30194, n30195, n30196, n30197, n30198, n30199,
    n30200, n30201, n30202, n30203, n30204, n30205,
    n30206, n30207, n30208, n30209, n30210, n30211,
    n30212, n30213, n30214, n30215, n30216, n30217,
    n30218, n30219, n30220, n30221, n30222, n30223,
    n30224, n30225, n30226, n30227, n30228, n30229,
    n30230, n30231, n30232, n30233, n30234, n30235,
    n30236, n30237, n30238, n30239, n30240, n30241,
    n30242, n30243, n30244, n30245, n30246, n30247,
    n30248, n30249, n30250, n30251, n30252, n30253,
    n30254, n30255, n30256, n30257, n30258, n30259,
    n30260, n30261, n30262, n30263, n30264, n30265,
    n30266, n30267, n30268, n30269, n30270, n30271,
    n30272, n30273, n30274, n30275, n30276, n30277,
    n30278, n30279, n30280, n30281, n30282, n30283,
    n30284, n30285, n30286, n30287, n30288, n30289,
    n30290, n30291, n30292, n30293, n30294, n30295,
    n30296, n30297, n30298, n30299, n30300, n30301,
    n30302, n30303, n30304, n30305, n30306, n30307,
    n30308, n30309, n30310, n30311, n30312, n30313,
    n30314, n30315, n30316, n30317, n30318, n30319,
    n30320, n30321, n30322, n30323, n30324, n30325,
    n30326, n30327, n30328, n30329, n30330, n30331,
    n30332, n30333, n30334, n30335, n30336, n30337,
    n30338, n30339, n30340, n30341, n30342, n30343,
    n30344, n30345, n30346, n30347, n30348, n30349,
    n30350, n30351, n30352, n30353, n30354, n30355,
    n30356, n30357, n30358, n30359, n30360, n30361,
    n30362, n30363, n30364, n30365, n30366, n30367,
    n30368, n30369, n30370, n30371, n30372, n30373,
    n30374, n30375, n30376, n30377, n30378, n30379,
    n30380, n30381, n30382, n30383, n30384, n30385,
    n30386, n30387, n30388, n30389, n30390, n30391,
    n30392, n30393, n30394, n30395, n30396, n30397,
    n30398, n30399, n30400, n30401, n30402, n30403,
    n30404, n30405, n30406, n30407, n30408, n30409,
    n30410, n30411, n30412, n30413, n30414, n30415,
    n30416, n30417, n30418, n30419, n30420, n30421,
    n30422, n30423, n30424, n30425, n30426, n30427,
    n30428, n30429, n30430, n30431, n30432, n30433,
    n30434, n30435, n30436, n30437, n30438, n30439,
    n30440, n30441, n30442, n30443, n30444, n30445,
    n30446, n30447, n30448, n30449, n30450, n30451,
    n30452, n30453, n30454, n30455, n30456, n30457,
    n30458, n30459, n30460, n30461, n30462, n30463,
    n30464, n30465, n30466, n30467, n30468, n30469,
    n30470, n30471, n30472, n30473, n30474, n30475,
    n30476, n30477, n30478, n30479, n30480, n30481,
    n30482, n30483, n30484, n30485, n30486, n30487,
    n30488, n30489, n30490, n30491, n30492, n30493,
    n30494, n30495, n30496, n30497, n30498, n30499,
    n30500, n30501, n30502, n30503, n30504, n30505,
    n30506, n30507, n30508, n30509, n30510, n30511,
    n30512, n30513, n30514, n30515, n30516, n30517,
    n30518, n30519, n30520, n30521, n30522, n30523,
    n30524, n30525, n30526, n30527, n30528, n30529,
    n30530, n30531, n30532, n30533, n30534, n30535,
    n30536, n30537, n30538, n30539, n30540, n30541,
    n30542, n30543, n30544, n30545, n30546, n30547,
    n30548, n30549, n30550, n30551, n30552, n30553,
    n30554, n30555, n30556, n30557, n30558, n30559,
    n30560, n30561, n30562, n30563, n30564, n30565,
    n30566, n30567, n30568, n30569, n30570, n30571,
    n30572, n30573, n30574, n30575, n30576, n30577,
    n30578, n30579, n30580, n30581, n30582, n30583,
    n30584, n30585, n30586, n30587, n30588, n30589,
    n30590, n30591, n30592, n30593, n30594, n30595,
    n30596, n30597, n30598, n30599, n30600, n30601,
    n30602, n30603, n30604, n30605, n30606, n30607,
    n30608, n30609, n30610, n30611, n30612, n30613,
    n30614, n30615, n30616, n30617, n30618, n30619,
    n30620, n30621, n30622, n30623, n30624, n30625,
    n30626, n30627, n30628, n30629, n30630, n30631,
    n30632, n30633, n30634, n30635, n30636, n30637,
    n30638, n30639, n30640, n30641, n30642, n30643,
    n30644, n30645, n30646, n30647, n30648, n30649,
    n30650, n30651, n30652, n30653, n30654, n30655,
    n30656, n30657, n30658, n30659, n30660, n30661,
    n30662, n30663, n30664, n30665, n30666, n30667,
    n30668, n30669, n30670, n30671, n30672, n30673,
    n30674, n30675, n30676, n30677, n30678, n30679,
    n30680, n30681, n30682, n30683, n30684, n30685,
    n30686, n30687, n30688, n30689, n30690, n30691,
    n30692, n30693, n30694, n30695, n30696, n30697,
    n30698, n30699, n30700, n30701, n30702, n30703,
    n30704, n30705, n30706, n30707, n30708, n30709,
    n30710, n30711, n30712, n30713, n30714, n30715,
    n30716, n30717, n30718, n30719, n30720, n30721,
    n30722, n30723, n30724, n30725, n30726, n30727,
    n30728, n30729, n30730, n30731, n30732, n30733,
    n30734, n30735, n30736, n30737, n30738, n30739,
    n30740, n30741, n30742, n30743, n30744, n30745,
    n30746, n30747, n30748, n30749, n30750, n30751,
    n30752, n30753, n30754, n30755, n30756, n30757,
    n30758, n30759, n30760, n30761, n30762, n30763,
    n30764, n30765, n30766, n30767, n30768, n30769,
    n30770, n30771, n30772, n30773, n30774, n30775,
    n30776, n30777, n30778, n30779, n30780, n30781,
    n30782, n30783, n30784, n30785, n30786, n30787,
    n30788, n30789, n30790, n30791, n30792, n30793,
    n30794, n30795, n30796, n30797, n30798, n30799,
    n30800, n30801, n30802, n30803, n30804, n30805,
    n30806, n30807, n30808, n30809, n30810, n30811,
    n30812, n30813, n30814, n30815, n30816, n30817,
    n30818, n30819, n30820, n30821, n30822, n30823,
    n30824, n30825, n30826, n30827, n30828, n30829,
    n30830, n30831, n30832, n30833, n30834, n30835,
    n30836, n30837, n30838, n30839, n30840, n30841,
    n30842, n30843, n30844, n30845, n30846, n30847,
    n30848, n30849, n30850, n30851, n30852, n30853,
    n30854, n30855, n30856, n30857, n30858, n30859,
    n30860, n30861, n30862, n30863, n30864, n30865,
    n30866, n30867, n30868, n30869, n30870, n30871,
    n30872, n30873, n30874, n30875, n30876, n30877,
    n30878, n30879, n30880, n30881, n30882, n30883,
    n30884, n30885, n30886, n30887, n30888, n30889,
    n30890, n30891, n30892, n30893, n30894, n30895,
    n30896, n30897, n30898, n30899, n30900, n30901,
    n30902, n30903, n30904, n30905, n30906, n30907,
    n30908, n30909, n30910, n30911, n30912, n30913,
    n30914, n30915, n30916, n30917, n30918, n30919,
    n30920, n30921, n30922, n30923, n30924, n30925,
    n30926, n30927, n30928, n30929, n30930, n30931,
    n30932, n30933, n30934, n30935, n30936, n30937,
    n30938, n30939, n30940, n30941, n30942, n30943,
    n30944, n30945, n30946, n30947, n30948, n30949,
    n30950, n30951, n30952, n30953, n30954, n30955,
    n30956, n30957, n30958, n30959, n30960, n30961,
    n30962, n30963, n30964, n30965, n30966, n30967,
    n30968, n30969, n30970, n30971, n30972, n30973,
    n30974, n30975, n30976, n30977, n30978, n30979,
    n30980, n30981, n30982, n30983, n30984, n30985,
    n30986, n30987, n30988, n30989, n30990, n30991,
    n30992, n30993, n30994, n30995, n30996, n30997,
    n30998, n30999, n31000, n31001, n31002, n31003,
    n31004, n31005, n31006, n31007, n31008, n31009,
    n31010, n31011, n31012, n31013, n31014, n31015,
    n31016, n31017, n31018, n31019, n31020, n31021,
    n31022, n31023, n31024, n31025, n31026, n31027,
    n31028, n31029, n31030, n31031, n31032, n31033,
    n31034, n31035, n31036, n31037, n31038, n31039,
    n31040, n31041, n31042, n31043, n31044, n31045,
    n31046, n31047, n31048, n31049, n31050, n31051,
    n31052, n31053, n31054, n31055, n31056, n31057,
    n31058, n31059, n31060, n31061, n31062, n31063,
    n31064, n31065, n31066, n31067, n31068, n31069,
    n31070, n31071, n31072, n31073, n31074, n31075,
    n31076, n31077, n31078, n31079, n31080, n31081,
    n31082, n31083, n31084, n31085, n31086, n31087,
    n31088, n31089, n31090, n31091, n31092, n31093,
    n31094, n31095, n31096, n31097, n31098, n31099,
    n31100, n31101, n31102, n31103, n31104, n31105,
    n31106, n31107, n31108, n31109, n31110, n31111,
    n31112, n31113, n31114, n31115, n31116, n31117,
    n31118, n31119, n31120, n31121, n31122, n31123,
    n31124, n31125, n31126, n31127, n31128, n31129,
    n31130, n31131, n31132, n31133, n31134, n31135,
    n31136, n31137, n31138, n31139, n31140, n31141,
    n31142, n31143, n31144, n31145, n31146, n31147,
    n31148, n31149, n31150, n31151, n31152, n31153,
    n31154, n31155, n31156, n31157, n31158, n31159,
    n31160, n31161, n31162, n31163, n31164, n31165,
    n31166, n31167, n31168, n31169, n31170, n31171,
    n31172, n31173, n31174, n31175, n31176, n31177,
    n31178, n31179, n31180, n31181, n31182, n31183,
    n31184, n31185, n31186, n31187, n31188, n31189,
    n31190, n31191, n31192, n31193, n31194, n31195,
    n31196, n31197, n31198, n31199, n31200, n31201,
    n31202, n31203, n31204, n31205, n31206, n31207,
    n31208, n31209, n31210, n31211, n31212, n31213,
    n31214, n31215, n31216, n31217, n31218, n31219,
    n31220, n31221, n31222, n31223, n31224, n31225,
    n31226, n31227, n31228, n31229, n31230, n31231,
    n31232, n31233, n31234, n31235, n31236, n31237,
    n31238, n31239, n31240, n31241, n31242, n31243,
    n31244, n31245, n31246, n31247, n31248, n31249,
    n31250, n31251, n31252, n31253, n31254, n31255,
    n31256, n31257, n31258, n31259, n31260, n31261,
    n31262, n31263, n31264, n31265, n31266, n31267,
    n31268, n31269, n31270, n31271, n31272, n31273,
    n31274, n31275, n31276, n31277, n31278, n31279,
    n31280, n31281, n31282, n31283, n31284, n31285,
    n31286, n31287, n31288, n31289, n31290, n31291,
    n31292, n31293, n31294, n31295, n31296, n31297,
    n31298, n31299, n31300, n31301, n31302, n31303,
    n31304, n31305, n31306, n31307, n31308, n31309,
    n31310, n31311, n31312, n31313, n31314, n31315,
    n31316, n31317, n31318, n31319, n31320, n31321,
    n31322, n31323, n31324, n31325, n31326, n31327,
    n31328, n31329, n31330, n31331, n31332, n31333,
    n31334, n31335, n31336, n31337, n31338, n31339,
    n31340, n31341, n31342, n31343, n31344, n31345,
    n31346, n31347, n31348, n31349, n31350, n31351,
    n31352, n31353, n31354, n31355, n31356, n31357,
    n31358, n31359, n31360, n31361, n31362, n31363,
    n31364, n31365, n31366, n31367, n31368, n31369,
    n31370, n31371, n31372, n31373, n31374, n31375,
    n31376, n31377, n31378, n31379, n31380, n31381,
    n31382, n31383, n31384, n31385, n31386, n31387,
    n31388, n31389, n31390, n31391, n31392, n31393,
    n31394, n31395, n31396, n31397, n31398, n31399,
    n31400, n31401, n31402, n31403, n31404, n31405,
    n31406, n31407, n31408, n31409, n31410, n31411,
    n31412, n31413, n31414, n31415, n31416, n31417,
    n31418, n31419, n31420, n31421, n31422, n31423,
    n31424, n31425, n31426, n31427, n31428, n31429,
    n31430, n31431, n31432, n31433, n31434, n31435,
    n31436, n31437, n31438, n31439, n31440, n31441,
    n31442, n31443, n31444, n31445, n31446, n31447,
    n31448, n31449, n31450, n31451, n31452, n31453,
    n31454, n31455, n31456, n31457, n31458, n31459,
    n31460, n31461, n31462, n31463, n31464, n31465,
    n31466, n31467, n31468, n31469, n31470, n31471,
    n31472, n31473, n31474, n31475, n31476, n31477,
    n31478, n31479, n31480, n31481, n31482, n31483,
    n31484, n31485, n31486, n31487, n31488, n31489,
    n31490, n31491, n31492, n31493, n31494, n31495,
    n31496, n31497, n31498, n31499, n31500, n31501,
    n31502, n31503, n31504, n31505, n31506, n31507,
    n31508, n31509, n31510, n31511, n31512, n31513,
    n31514, n31515, n31516, n31517, n31518, n31519,
    n31520, n31521, n31522, n31523, n31524, n31525,
    n31526, n31527, n31528, n31529, n31530, n31531,
    n31532, n31533, n31534, n31535, n31536, n31537,
    n31538, n31539, n31540, n31541, n31542, n31543,
    n31544, n31545, n31546, n31547, n31548, n31549,
    n31550, n31551, n31552, n31553, n31554, n31555,
    n31556, n31557, n31558, n31559, n31560, n31561,
    n31562, n31563, n31564, n31565, n31566, n31567,
    n31568, n31569, n31570, n31571, n31572, n31573,
    n31574, n31575, n31576, n31577, n31578, n31579,
    n31580, n31581, n31582, n31583, n31584, n31585,
    n31586, n31587, n31588, n31589, n31590, n31591,
    n31592, n31593, n31594, n31595, n31596, n31597,
    n31598, n31599, n31600, n31601, n31602, n31603,
    n31604, n31605, n31606, n31607, n31608, n31609,
    n31610, n31611, n31612, n31613, n31614, n31615,
    n31616, n31617, n31618, n31619, n31620, n31621,
    n31622, n31623, n31624, n31625, n31626, n31627,
    n31628, n31629, n31630, n31631, n31632, n31633,
    n31634, n31635, n31636, n31637, n31638, n31639,
    n31640, n31641, n31642, n31643, n31644, n31645,
    n31646, n31647, n31648, n31649, n31650, n31651,
    n31652, n31653, n31654, n31655, n31656, n31657,
    n31658, n31659, n31660, n31661, n31662, n31663,
    n31664, n31665, n31666, n31667, n31668, n31669,
    n31670, n31671, n31672, n31673, n31674, n31675,
    n31676, n31677, n31678, n31679, n31680, n31681,
    n31682, n31683, n31684, n31685, n31686, n31687,
    n31688, n31689, n31690, n31691, n31692, n31693,
    n31694, n31695, n31696, n31697, n31698, n31699,
    n31700, n31701, n31702, n31703, n31704, n31705,
    n31706, n31707, n31708, n31709, n31710, n31711,
    n31712, n31713, n31714, n31715, n31716, n31717,
    n31718, n31719, n31720, n31721, n31722, n31723,
    n31724, n31725, n31726, n31727, n31728, n31729,
    n31730, n31731, n31732, n31733, n31734, n31735,
    n31736, n31737, n31738, n31739, n31740, n31741,
    n31742, n31743, n31744, n31745, n31746, n31747,
    n31748, n31749, n31750, n31751, n31752, n31753,
    n31754, n31755, n31756, n31757, n31758, n31759,
    n31760, n31761, n31762, n31763, n31764, n31765,
    n31766, n31767, n31768, n31769, n31770, n31771,
    n31772, n31773, n31774, n31775, n31776, n31777,
    n31778, n31779, n31780, n31781, n31782, n31783,
    n31784, n31785, n31786, n31787, n31788, n31789,
    n31790, n31791, n31792, n31793, n31794, n31795,
    n31796, n31797, n31798, n31799, n31800, n31801,
    n31802, n31803, n31804, n31805, n31806, n31807,
    n31808, n31809, n31810, n31811, n31812, n31813,
    n31814, n31815, n31816, n31817, n31818, n31819,
    n31820, n31821, n31822, n31823, n31824, n31825,
    n31826, n31827, n31828, n31829, n31830, n31831,
    n31832, n31833, n31834, n31835, n31836, n31837,
    n31838, n31839, n31840, n31841, n31842, n31843,
    n31844, n31845, n31846, n31847, n31848, n31849,
    n31850, n31851, n31852, n31853, n31854, n31855,
    n31856, n31857, n31858, n31859, n31860, n31861,
    n31862, n31863, n31864, n31865, n31866, n31867,
    n31868, n31869, n31870, n31871, n31872, n31873,
    n31874, n31875, n31876, n31877, n31878, n31879,
    n31880, n31881, n31882, n31883, n31884, n31885,
    n31886, n31887, n31888, n31889, n31890, n31891,
    n31892, n31893, n31894, n31895, n31896, n31897,
    n31898, n31899, n31900, n31901, n31902, n31903,
    n31904, n31905, n31906, n31907, n31908, n31909,
    n31910, n31911, n31912, n31913, n31914, n31915,
    n31916, n31917, n31918, n31919, n31920, n31921,
    n31922, n31923, n31924, n31925, n31926, n31927,
    n31928, n31929, n31930, n31931, n31932, n31933,
    n31934, n31935, n31936, n31937, n31938, n31939,
    n31940, n31941, n31942, n31943, n31944, n31945,
    n31946, n31947, n31948, n31949, n31950, n31951,
    n31952, n31953, n31954, n31955, n31956, n31957,
    n31958, n31959, n31960, n31961, n31962, n31963,
    n31964, n31965, n31966, n31967, n31968, n31969,
    n31970, n31971, n31972, n31973, n31974, n31975,
    n31976, n31977, n31978, n31979, n31980, n31981,
    n31982, n31983, n31984, n31985, n31986, n31987,
    n31988, n31989, n31990, n31991, n31992, n31993,
    n31994, n31995, n31996, n31997, n31998, n31999,
    n32000, n32001, n32002, n32003, n32004, n32005,
    n32006, n32007, n32008, n32009, n32010, n32011,
    n32012, n32013, n32014, n32015, n32016, n32017,
    n32018, n32019, n32020, n32021, n32022, n32023,
    n32024, n32025, n32026, n32027, n32028, n32029,
    n32030, n32031, n32032, n32033, n32034, n32035,
    n32036, n32037, n32038, n32039, n32040, n32041,
    n32042, n32043, n32044, n32045, n32046, n32047,
    n32048, n32049, n32050, n32051, n32052, n32053,
    n32054, n32055, n32056, n32057, n32058, n32059,
    n32060, n32061, n32062, n32063, n32064, n32065,
    n32066, n32067, n32068, n32069, n32070, n32071,
    n32072, n32073, n32074, n32075, n32076, n32077,
    n32078, n32079, n32080, n32081, n32082, n32083,
    n32084, n32085, n32086, n32087, n32088, n32089,
    n32090, n32091, n32092, n32093, n32094, n32095,
    n32096, n32097, n32098, n32099, n32100, n32101,
    n32102, n32103, n32104, n32105, n32106, n32107,
    n32108, n32109, n32110, n32111, n32112, n32113,
    n32114, n32115, n32116, n32117, n32118, n32119,
    n32120, n32121, n32122, n32123, n32124, n32125,
    n32126, n32127, n32128, n32129, n32130, n32131,
    n32132, n32133, n32134, n32135, n32136, n32137,
    n32138, n32139, n32140, n32141, n32142, n32143,
    n32144, n32145, n32146, n32147, n32148, n32149,
    n32150, n32151, n32152, n32153, n32154, n32155,
    n32156, n32157, n32158, n32159, n32160, n32161,
    n32162, n32163, n32164, n32165, n32166, n32167,
    n32168, n32169, n32170, n32171, n32172, n32173,
    n32174, n32175, n32176, n32177, n32178, n32179,
    n32180, n32181, n32182, n32183, n32184, n32185,
    n32186, n32187, n32188, n32189, n32190, n32191,
    n32192, n32193, n32194, n32195, n32196, n32197,
    n32198, n32199, n32200, n32201, n32202, n32203,
    n32204, n32205, n32206, n32207, n32208, n32209,
    n32210, n32211, n32212, n32213, n32214, n32215,
    n32216, n32217, n32218, n32219, n32220, n32221,
    n32222, n32223, n32224, n32225, n32226, n32227,
    n32228, n32229, n32230, n32231, n32232, n32233,
    n32234, n32235, n32236, n32237, n32238, n32239,
    n32240, n32241, n32242, n32243, n32244, n32245,
    n32246, n32247, n32248, n32249, n32250, n32251,
    n32252, n32253, n32254, n32255, n32256, n32257,
    n32258, n32259, n32260, n32261, n32262, n32263,
    n32264, n32265, n32266, n32267, n32268, n32269,
    n32270, n32271, n32272, n32273, n32274, n32275,
    n32276, n32277, n32278, n32279, n32280, n32281,
    n32282, n32283, n32284, n32285, n32286, n32287,
    n32288, n32289, n32290, n32291, n32292, n32293,
    n32294, n32295, n32296, n32297, n32298, n32299,
    n32300, n32301, n32302, n32303, n32304, n32305,
    n32306, n32307, n32308, n32309, n32310, n32311,
    n32312, n32313, n32314, n32315, n32316, n32317,
    n32318, n32319, n32320, n32321, n32322, n32323,
    n32324, n32325, n32326, n32327, n32328, n32329,
    n32330, n32331, n32332, n32333, n32334, n32335,
    n32336, n32337, n32338, n32339, n32340, n32341,
    n32342, n32343, n32344, n32345, n32346, n32347,
    n32348, n32349, n32350, n32351, n32352, n32353,
    n32354, n32355, n32356, n32357, n32358, n32359,
    n32360, n32361, n32362, n32363, n32364, n32365,
    n32366, n32367, n32368, n32369, n32370, n32371,
    n32372, n32373, n32374, n32375, n32376, n32377,
    n32378, n32379, n32380, n32381, n32382, n32383,
    n32384, n32385, n32386, n32387, n32388, n32389,
    n32390, n32391, n32392, n32393, n32394, n32395,
    n32396, n32397, n32398, n32399, n32400, n32401,
    n32402, n32403, n32404, n32405, n32406, n32407,
    n32408, n32409, n32410, n32411, n32412, n32413,
    n32414, n32415, n32416, n32417, n32418, n32419,
    n32420, n32421, n32422, n32423, n32424, n32425,
    n32426, n32427, n32428, n32429, n32430, n32431,
    n32432, n32433, n32434, n32435, n32436, n32437,
    n32438, n32439, n32440, n32441, n32442, n32443,
    n32444, n32445, n32446, n32447, n32448, n32449,
    n32450, n32451, n32452, n32453, n32454, n32455,
    n32456, n32457, n32458, n32459, n32460, n32461,
    n32462, n32463, n32464, n32465, n32466, n32467,
    n32468, n32469, n32470, n32471, n32472, n32473,
    n32474, n32475, n32476, n32477, n32478, n32479,
    n32480, n32481, n32482, n32483, n32484, n32485,
    n32486, n32487, n32488, n32489, n32490, n32491,
    n32492, n32493, n32494, n32495, n32496, n32497,
    n32498, n32499, n32500, n32501, n32502, n32503,
    n32504, n32505, n32506, n32507, n32508, n32509,
    n32510, n32511, n32512, n32513, n32514, n32515,
    n32516, n32517, n32518, n32519, n32520, n32521,
    n32522, n32523, n32524, n32525, n32526, n32527,
    n32528, n32529, n32530, n32531, n32532, n32533,
    n32534, n32535, n32536, n32537, n32538, n32539,
    n32540, n32541, n32542, n32543, n32544, n32545,
    n32546, n32547, n32548, n32549, n32550, n32551,
    n32552, n32553, n32554, n32555, n32556, n32557,
    n32558, n32559, n32560, n32561, n32562, n32563,
    n32564, n32565, n32566, n32567, n32568, n32569,
    n32570, n32571, n32572, n32573, n32574, n32575,
    n32576, n32577, n32578, n32579, n32580, n32581,
    n32582, n32583, n32584, n32585, n32586, n32587,
    n32588, n32589, n32590, n32591, n32592, n32593,
    n32594, n32595, n32596, n32597, n32598, n32599,
    n32600, n32601, n32602, n32603, n32604, n32605,
    n32606, n32607, n32608, n32609, n32610, n32611,
    n32612, n32613, n32614, n32615, n32616, n32617,
    n32618, n32619, n32620, n32621, n32622, n32623,
    n32624, n32625, n32626, n32627, n32628, n32629,
    n32630, n32631, n32632, n32633, n32634, n32635,
    n32636, n32637, n32638, n32639, n32640, n32641,
    n32642, n32643, n32644, n32645, n32646, n32647,
    n32648, n32649, n32650, n32651, n32652, n32653,
    n32654, n32655, n32656, n32657, n32658, n32659,
    n32660, n32661, n32662, n32663, n32664, n32665,
    n32666, n32667, n32668, n32669, n32670, n32671,
    n32672, n32673, n32674, n32675, n32676, n32677,
    n32678, n32679, n32680, n32681, n32682, n32683,
    n32684, n32685, n32686, n32687, n32688, n32689,
    n32690, n32691, n32692, n32693, n32694, n32695,
    n32696, n32697, n32698, n32699, n32700, n32701,
    n32702, n32703, n32704, n32705, n32706, n32707,
    n32708, n32709, n32710, n32711, n32712, n32713,
    n32714, n32715, n32716, n32717, n32718, n32719,
    n32720, n32721, n32722, n32723, n32724, n32725,
    n32726, n32727, n32728, n32729, n32730, n32731,
    n32732, n32733, n32734, n32735, n32736, n32737,
    n32738, n32739, n32740, n32741, n32742, n32743,
    n32744, n32745, n32746, n32747, n32748, n32749,
    n32750, n32751, n32752, n32753, n32754, n32755,
    n32756, n32757, n32758, n32759, n32760, n32761,
    n32762, n32763, n32764, n32765, n32766, n32767,
    n32768, n32769, n32770, n32771, n32772, n32773,
    n32774, n32775, n32776, n32777, n32778, n32779,
    n32780, n32781, n32782, n32783, n32784, n32785,
    n32786, n32787, n32788, n32789, n32790, n32791,
    n32792, n32793, n32794, n32795, n32796, n32797,
    n32798, n32799, n32800, n32801, n32802, n32803,
    n32804, n32805, n32806, n32807, n32808, n32809,
    n32810, n32811, n32812, n32813, n32814, n32815,
    n32816, n32817, n32818, n32819, n32820, n32821,
    n32822, n32823, n32824, n32825, n32826, n32827,
    n32828, n32829, n32830, n32831, n32832, n32833,
    n32834, n32835, n32836, n32837, n32838, n32839,
    n32840, n32841, n32842, n32843, n32844, n32845,
    n32846, n32847, n32848, n32849, n32850, n32851,
    n32852, n32853, n32854, n32855, n32856, n32857,
    n32858, n32859, n32860, n32861, n32862, n32863,
    n32864, n32865, n32866, n32867, n32868, n32869,
    n32870, n32871, n32872, n32873, n32874, n32875,
    n32876, n32877, n32878, n32879, n32880, n32881,
    n32882, n32883, n32884, n32885, n32886, n32887,
    n32888, n32889, n32890, n32891, n32892, n32893,
    n32894, n32895, n32896, n32897, n32898, n32899,
    n32900, n32901, n32902, n32903, n32904, n32905,
    n32906, n32907, n32908, n32909, n32910, n32911,
    n32912, n32913, n32914, n32915, n32916, n32917,
    n32918, n32919, n32920, n32921, n32922, n32923,
    n32924, n32925, n32926, n32927, n32928, n32929,
    n32930, n32931, n32932, n32933, n32934, n32935,
    n32936, n32937, n32938, n32939, n32940, n32941,
    n32942, n32943, n32944, n32945, n32946, n32947,
    n32948, n32949, n32950, n32951, n32952, n32953,
    n32954, n32955, n32956, n32957, n32958, n32959,
    n32960, n32961, n32962, n32963, n32964, n32965,
    n32966, n32967, n32968, n32969, n32970, n32971,
    n32972, n32973, n32974, n32975, n32976, n32977,
    n32978, n32979, n32980, n32981, n32982, n32983,
    n32984, n32985, n32986, n32987, n32988, n32989,
    n32990, n32991, n32992, n32993, n32994, n32995,
    n32996, n32997, n32998, n32999, n33000, n33001,
    n33002, n33003, n33004, n33005, n33006, n33007,
    n33008, n33009, n33010, n33011, n33012, n33013,
    n33014, n33015, n33016, n33017, n33018, n33019,
    n33020, n33021, n33022, n33023, n33024, n33025,
    n33026, n33027, n33028, n33029, n33030, n33031,
    n33032, n33033, n33034, n33035, n33036, n33037,
    n33038, n33039, n33040, n33041, n33042, n33043,
    n33044, n33045, n33046, n33047, n33048, n33049,
    n33050, n33051, n33052, n33053, n33054, n33055,
    n33056, n33057, n33058, n33059, n33060, n33061,
    n33062, n33063, n33064, n33065, n33066, n33067,
    n33068, n33069, n33070, n33071, n33072, n33073,
    n33074, n33075, n33076, n33077, n33078, n33079,
    n33080, n33081, n33082, n33083, n33084, n33085,
    n33086, n33087, n33088, n33089, n33090, n33091,
    n33092, n33093, n33094, n33095, n33096, n33097,
    n33098, n33099, n33100, n33101, n33102, n33103,
    n33104, n33105, n33106, n33107, n33108, n33109,
    n33110, n33111, n33112, n33113, n33114, n33115,
    n33116, n33117, n33118, n33119, n33120, n33121,
    n33122, n33123, n33124, n33125, n33126, n33127,
    n33128, n33129, n33130, n33131, n33132, n33133,
    n33134, n33135, n33136, n33137, n33138, n33139,
    n33140, n33141, n33142, n33143, n33144, n33145,
    n33146, n33147, n33148, n33149, n33150, n33151,
    n33152, n33153, n33154, n33155, n33156, n33157,
    n33158, n33159, n33160, n33161, n33162, n33163,
    n33164, n33165, n33166, n33167, n33168, n33169,
    n33170, n33171, n33172, n33173, n33174, n33175,
    n33176, n33177, n33178, n33179, n33180, n33181,
    n33182, n33183, n33184, n33185, n33186, n33187,
    n33188, n33189, n33190, n33191, n33192, n33193,
    n33194, n33195, n33196, n33197, n33198, n33199,
    n33200, n33201, n33202, n33203, n33204, n33205,
    n33206, n33207, n33208, n33209, n33210, n33211,
    n33212, n33213, n33214, n33215, n33216, n33217,
    n33218, n33219, n33220, n33221, n33222, n33223,
    n33224, n33225, n33226, n33227, n33228, n33229,
    n33230, n33231, n33232, n33233, n33234, n33235,
    n33236, n33237, n33238, n33239, n33240, n33241,
    n33242, n33243, n33244, n33245, n33246, n33247,
    n33248, n33249, n33250, n33251, n33252, n33253,
    n33254, n33255, n33256, n33257, n33258, n33259,
    n33260, n33261, n33262, n33263, n33264, n33265,
    n33266, n33267, n33268, n33269, n33270, n33271,
    n33272, n33273, n33274, n33275, n33276, n33277,
    n33278, n33279, n33280, n33281, n33282, n33283,
    n33284, n33285, n33286, n33287, n33288, n33289,
    n33290, n33291, n33292, n33293, n33294, n33295,
    n33296, n33297, n33298, n33299, n33300, n33301,
    n33302, n33303, n33304, n33305, n33306, n33307,
    n33308, n33309, n33310, n33311, n33312, n33313,
    n33314, n33315, n33316, n33317, n33318, n33319,
    n33320, n33321, n33322, n33323, n33324, n33325,
    n33326, n33327, n33328, n33329, n33330, n33331,
    n33332, n33333, n33334, n33335, n33336, n33337,
    n33338, n33339, n33340, n33341, n33342, n33343,
    n33344, n33345, n33346, n33347, n33348, n33349,
    n33350, n33351, n33352, n33353, n33354, n33355,
    n33356, n33357, n33358, n33359, n33360, n33361,
    n33362, n33363, n33364, n33365, n33366, n33367,
    n33368, n33369, n33370, n33371, n33372, n33373,
    n33374, n33375, n33376, n33377, n33378, n33379,
    n33380, n33381, n33382, n33383, n33384, n33385,
    n33386, n33387, n33388, n33389, n33390, n33391,
    n33392, n33393, n33394, n33395, n33396, n33397,
    n33398, n33399, n33400, n33401, n33402, n33403,
    n33404, n33405, n33406, n33407, n33408, n33409,
    n33410, n33411, n33412, n33413, n33414, n33415,
    n33416, n33417, n33418, n33419, n33420, n33421,
    n33422, n33423, n33424, n33425, n33426, n33427,
    n33428, n33429, n33430, n33431, n33432, n33433,
    n33434, n33435, n33436, n33437, n33438, n33439,
    n33440, n33441, n33442, n33443, n33444, n33445,
    n33446, n33447, n33448, n33449, n33450, n33451,
    n33452, n33453, n33454, n33455, n33456, n33457,
    n33458, n33459, n33460, n33461, n33462, n33463,
    n33464, n33465, n33466, n33467, n33468, n33469,
    n33470, n33471, n33472, n33473, n33474, n33475,
    n33476, n33477, n33478, n33479, n33480, n33481,
    n33482, n33483, n33484, n33485, n33486, n33487,
    n33488, n33489, n33490, n33491, n33492, n33493,
    n33494, n33495, n33496, n33497, n33498, n33499,
    n33500, n33501, n33502, n33503, n33504, n33505,
    n33506, n33507, n33508, n33509, n33510, n33511,
    n33512, n33513, n33514, n33515, n33516, n33517,
    n33518, n33519, n33520, n33521, n33522, n33523,
    n33524, n33525, n33526, n33527, n33528, n33529,
    n33530, n33531, n33532, n33533, n33534, n33535,
    n33536, n33537, n33538, n33539, n33540, n33541,
    n33542, n33543, n33544, n33545, n33546, n33547,
    n33548, n33549, n33550, n33551, n33552, n33553,
    n33554, n33555, n33556, n33557, n33558, n33559,
    n33560, n33561, n33562, n33563, n33564, n33565,
    n33566, n33567, n33568, n33569, n33570, n33571,
    n33572, n33573, n33574, n33575, n33576, n33577,
    n33578, n33579, n33580, n33581, n33582, n33583,
    n33584, n33585, n33586, n33587, n33588, n33589,
    n33590, n33591, n33592, n33593, n33594, n33595,
    n33596, n33597, n33598, n33599, n33600, n33601,
    n33602, n33603, n33604, n33605, n33606, n33607,
    n33608, n33609, n33610, n33611, n33612, n33613,
    n33614, n33615, n33616, n33617, n33618, n33619,
    n33620, n33621, n33622, n33623, n33624, n33625,
    n33626, n33627, n33628, n33629, n33630, n33631,
    n33632, n33633, n33634, n33635, n33636, n33637,
    n33638, n33639, n33640, n33641, n33642, n33643,
    n33644, n33645, n33646, n33647, n33648, n33649,
    n33650, n33651, n33652, n33653, n33654, n33655,
    n33656, n33657, n33658, n33659, n33660, n33661,
    n33662, n33663, n33664, n33665, n33666, n33667,
    n33668, n33669, n33670, n33671, n33672, n33673,
    n33674, n33675, n33676, n33677, n33678, n33679,
    n33680, n33681, n33682, n33683, n33684, n33685,
    n33686, n33687, n33688, n33689, n33690, n33691,
    n33692, n33693, n33694, n33695, n33696, n33697,
    n33698, n33699, n33700, n33701, n33702, n33703,
    n33704, n33705, n33706, n33707, n33708, n33709,
    n33710, n33711, n33712, n33713, n33714, n33715,
    n33716, n33717, n33718, n33719, n33720, n33721,
    n33722, n33723, n33724, n33725, n33726, n33727,
    n33728, n33729, n33730, n33731, n33732, n33733,
    n33734, n33735, n33736, n33737, n33738, n33739,
    n33740, n33741, n33742, n33743, n33744, n33745,
    n33746, n33747, n33748, n33749, n33750, n33751,
    n33752, n33753, n33754, n33755, n33756, n33757,
    n33758, n33759, n33760, n33761, n33762, n33763,
    n33764, n33765, n33766, n33767, n33768, n33769,
    n33770, n33771, n33772, n33773, n33774, n33775,
    n33776, n33777, n33778, n33779, n33780, n33781,
    n33782, n33783, n33784, n33785, n33786, n33787,
    n33788, n33789, n33790, n33791, n33792, n33793,
    n33794, n33795, n33796, n33797, n33798, n33799,
    n33800, n33801, n33802, n33803, n33804, n33805,
    n33806, n33807, n33808, n33809, n33810, n33811,
    n33812, n33813, n33814, n33815, n33816, n33817,
    n33818, n33819, n33820, n33821, n33822, n33823,
    n33824, n33825, n33826, n33827, n33828, n33829,
    n33830, n33831, n33832, n33833, n33834, n33835,
    n33836, n33837, n33838, n33839, n33840, n33841,
    n33842, n33843, n33844, n33845, n33846, n33847,
    n33848, n33849, n33850, n33851, n33852, n33853,
    n33854, n33855, n33856, n33857, n33858, n33859,
    n33860, n33861, n33862, n33863, n33864, n33865,
    n33866, n33867, n33868, n33869, n33870, n33871,
    n33872, n33873, n33874, n33875, n33876, n33877,
    n33878, n33879, n33880, n33881, n33882, n33883,
    n33884, n33885, n33886, n33887, n33888, n33889,
    n33890, n33891, n33892, n33893, n33894, n33895,
    n33896, n33897, n33898, n33899, n33900, n33901,
    n33902, n33903, n33904, n33905, n33906, n33907,
    n33908, n33909, n33910, n33911, n33912, n33913,
    n33914, n33915, n33916, n33917, n33918, n33919,
    n33920, n33921, n33922, n33923, n33924, n33925,
    n33926, n33927, n33928, n33929, n33930, n33931,
    n33932, n33933, n33934, n33935, n33936, n33937,
    n33938, n33939, n33940, n33941, n33942, n33943,
    n33944, n33945, n33946, n33947, n33948, n33949,
    n33950, n33951, n33952, n33953, n33954, n33955,
    n33956, n33957, n33958, n33959, n33960, n33961,
    n33962, n33963, n33964, n33965, n33966, n33967,
    n33968, n33969, n33970, n33971, n33972, n33973,
    n33974, n33975, n33976, n33977, n33978, n33979,
    n33980, n33981, n33982, n33983, n33984, n33985,
    n33986, n33987, n33988, n33989, n33990, n33991,
    n33992, n33993, n33994, n33995, n33996, n33997,
    n33998, n33999, n34000, n34001, n34002, n34003,
    n34004, n34005, n34006, n34007, n34008, n34009,
    n34010, n34011, n34012, n34013, n34014, n34015,
    n34016, n34017, n34018, n34019, n34020, n34021,
    n34022, n34023, n34024, n34025, n34026, n34027,
    n34028, n34029, n34030, n34031, n34032, n34033,
    n34034, n34035, n34036, n34037, n34038, n34039,
    n34040, n34041, n34042, n34043, n34044, n34045,
    n34046, n34047, n34048, n34049, n34050, n34051,
    n34052, n34053, n34054, n34055, n34056, n34057,
    n34058, n34059, n34060, n34061, n34062, n34063,
    n34064, n34065, n34066, n34067, n34068, n34069,
    n34070, n34071, n34072, n34073, n34074, n34075,
    n34076, n34077, n34078, n34079, n34080, n34081,
    n34082, n34083, n34084, n34085, n34086, n34087,
    n34088, n34089, n34090, n34091, n34092, n34093,
    n34094, n34095, n34096, n34097, n34098, n34099,
    n34100, n34101, n34102, n34103, n34104, n34105,
    n34106, n34107, n34108, n34109, n34110, n34111,
    n34112, n34113, n34114, n34115, n34116, n34117,
    n34118, n34119, n34120, n34121, n34122, n34123,
    n34124, n34125, n34126, n34127, n34128, n34129,
    n34130, n34131, n34132, n34133, n34134, n34135,
    n34136, n34137, n34138, n34139, n34140, n34141,
    n34142, n34143, n34144, n34145, n34146, n34147,
    n34148, n34149, n34150, n34151, n34152, n34153,
    n34154, n34155, n34156, n34157, n34158, n34159,
    n34160, n34161, n34162, n34163, n34164, n34165,
    n34166, n34167, n34168, n34169, n34170, n34171,
    n34172, n34173, n34174, n34175, n34176, n34177,
    n34178, n34179, n34180, n34181, n34182, n34183,
    n34184, n34185, n34186, n34187, n34188, n34189,
    n34190, n34191, n34192, n34193, n34194, n34195,
    n34196, n34197, n34198, n34199, n34200, n34201,
    n34202, n34203, n34204, n34205, n34206, n34207,
    n34208, n34209, n34210, n34211, n34212, n34213,
    n34214, n34215, n34216, n34217, n34218, n34219,
    n34220, n34221, n34222, n34223, n34224, n34225,
    n34226, n34227, n34228, n34229, n34230, n34231,
    n34232, n34233, n34234, n34235, n34236, n34237,
    n34238, n34239, n34240, n34241, n34242, n34243,
    n34244, n34245, n34246, n34247, n34248, n34249,
    n34250, n34251, n34252, n34253, n34254, n34255,
    n34256, n34257, n34258, n34259, n34260, n34261,
    n34262, n34263, n34264, n34265, n34266, n34267,
    n34268, n34269, n34270, n34271, n34272, n34273,
    n34274, n34275, n34276, n34277, n34278, n34279,
    n34280, n34281, n34282, n34283, n34284, n34285,
    n34286, n34287, n34288, n34289, n34290, n34291,
    n34292, n34293, n34294, n34295, n34296, n34297,
    n34298, n34299, n34300, n34301, n34302, n34303,
    n34304, n34305, n34306, n34307, n34308, n34309,
    n34310, n34311, n34312, n34313, n34314, n34315,
    n34316, n34317, n34318, n34319, n34320, n34321,
    n34322, n34323, n34324, n34325, n34326, n34327,
    n34328, n34329, n34330, n34331, n34332, n34333,
    n34334, n34335, n34336, n34337, n34338, n34339,
    n34340, n34341, n34342, n34343, n34344, n34345,
    n34346, n34347, n34348, n34349, n34350, n34351,
    n34352, n34353, n34354, n34355, n34356, n34357,
    n34358, n34359, n34360, n34361, n34362, n34363,
    n34364, n34365, n34366, n34367, n34368, n34369,
    n34370, n34371, n34372, n34373, n34374, n34375,
    n34376, n34377, n34378, n34379, n34380, n34381,
    n34382, n34383, n34384, n34385, n34386, n34387,
    n34388, n34389, n34390, n34391, n34392, n34393,
    n34394, n34395, n34396, n34397, n34398, n34399,
    n34400, n34401, n34402, n34403, n34404, n34405,
    n34406, n34407, n34408, n34409, n34410, n34411,
    n34412, n34413, n34414, n34415, n34416, n34417,
    n34418, n34419, n34420, n34421, n34422, n34423,
    n34424, n34425, n34426, n34427, n34428, n34429,
    n34430, n34431, n34432, n34433, n34434, n34435,
    n34436, n34437, n34438, n34439, n34440, n34441,
    n34442, n34443, n34444, n34445, n34446, n34447,
    n34448, n34449, n34450, n34451, n34452, n34453,
    n34454, n34455, n34456, n34457, n34458, n34459,
    n34460, n34461, n34462, n34463, n34464, n34465,
    n34466, n34467, n34468, n34469, n34470, n34471,
    n34472, n34473, n34474, n34475, n34476, n34477,
    n34478, n34479, n34480, n34481, n34482, n34483,
    n34484, n34485, n34486, n34487, n34488, n34489,
    n34490, n34491, n34492, n34493, n34494, n34495,
    n34496, n34497, n34498, n34499, n34500, n34501,
    n34502, n34503, n34504, n34505, n34506, n34507,
    n34508, n34509, n34510, n34511, n34512, n34513,
    n34514, n34515, n34516, n34517, n34518, n34519,
    n34520, n34521, n34522, n34523, n34524, n34525,
    n34526, n34527, n34528, n34529, n34530, n34531,
    n34532, n34533, n34534, n34535, n34536, n34537,
    n34538, n34539, n34540, n34541, n34542, n34543,
    n34544, n34545, n34546, n34547, n34548, n34549,
    n34550, n34551, n34552, n34553, n34554, n34555,
    n34556, n34557, n34558, n34559, n34560, n34561,
    n34562, n34563, n34564, n34565, n34566, n34567,
    n34568, n34569, n34570, n34571, n34572, n34573,
    n34574, n34575, n34576, n34577, n34578, n34579,
    n34580, n34581, n34582, n34583, n34584, n34585,
    n34586, n34587, n34588, n34589, n34590, n34591,
    n34592, n34593, n34594, n34595, n34596, n34597,
    n34598, n34599, n34600, n34601, n34602, n34603,
    n34604, n34605, n34606, n34607, n34608, n34609,
    n34610, n34611, n34612, n34613, n34614, n34615,
    n34616, n34617, n34618, n34619, n34620, n34621,
    n34622, n34623, n34624, n34625, n34626, n34627,
    n34628, n34629, n34630, n34631, n34632, n34633,
    n34634, n34635, n34636, n34637, n34638, n34639,
    n34640, n34641, n34642, n34643, n34644, n34645,
    n34646, n34647, n34648, n34649, n34650, n34651,
    n34652, n34653, n34654, n34655, n34656, n34657,
    n34658, n34659, n34660, n34661, n34662, n34663,
    n34664, n34665, n34666, n34667, n34668, n34669,
    n34670, n34671, n34672, n34673, n34674, n34675,
    n34676, n34677, n34678, n34679, n34680, n34681,
    n34682, n34683, n34684, n34685, n34686, n34687,
    n34688, n34689, n34690, n34691, n34692, n34693,
    n34694, n34695, n34696, n34697, n34698, n34699,
    n34700, n34701, n34702, n34703, n34704, n34705,
    n34706, n34707, n34708, n34709, n34710, n34711,
    n34712, n34713, n34714, n34715, n34716, n34717,
    n34718, n34719, n34720, n34721, n34722, n34723,
    n34724, n34725, n34726, n34727, n34728, n34729,
    n34730, n34731, n34732, n34733, n34734, n34735,
    n34736, n34737, n34738, n34739, n34740, n34741,
    n34742, n34743, n34744, n34745, n34746, n34747,
    n34748, n34749, n34750, n34751, n34752, n34753,
    n34754, n34755, n34756, n34757, n34758, n34759,
    n34760, n34761, n34762, n34763, n34764, n34765,
    n34766, n34767, n34768, n34769, n34770, n34771,
    n34772, n34773, n34774, n34775, n34776, n34777,
    n34778, n34779, n34780, n34781, n34782, n34783,
    n34784, n34785, n34786, n34787, n34788, n34789,
    n34790, n34791, n34792, n34793, n34794, n34795,
    n34796, n34797, n34798, n34799, n34800, n34801,
    n34802, n34803, n34804, n34805, n34806, n34807,
    n34808, n34809, n34810, n34811, n34812, n34813,
    n34814, n34815, n34816, n34817, n34818, n34819,
    n34820, n34821, n34822, n34823, n34824, n34825,
    n34826, n34827, n34828, n34829, n34830, n34831,
    n34832, n34833, n34834, n34835, n34836, n34837,
    n34838, n34839, n34840, n34841, n34842, n34843,
    n34844, n34845, n34846, n34847, n34848, n34849,
    n34850, n34851, n34852, n34853, n34854, n34855,
    n34856, n34857, n34858, n34859, n34860, n34861,
    n34862, n34863, n34864, n34865, n34866, n34867,
    n34868, n34869, n34870, n34871, n34872, n34873,
    n34874, n34875, n34876, n34877, n34878, n34879,
    n34880, n34881, n34882, n34883, n34884, n34885,
    n34886, n34887, n34888, n34889, n34890, n34891,
    n34892, n34893, n34894, n34895, n34896, n34897,
    n34898, n34899, n34900, n34901, n34902, n34903,
    n34904, n34905, n34906, n34907, n34908, n34909,
    n34910, n34911, n34912, n34913, n34914, n34915,
    n34916, n34917, n34918, n34919, n34920, n34921,
    n34922, n34923, n34924, n34925, n34926, n34927,
    n34928, n34929, n34930, n34931, n34932, n34933,
    n34934, n34935, n34936, n34937, n34938, n34939,
    n34940, n34941, n34942, n34943, n34944, n34945,
    n34946, n34947, n34948, n34949, n34950, n34951,
    n34952, n34953, n34954, n34955, n34956, n34957,
    n34958, n34959, n34960, n34961, n34962, n34963,
    n34964, n34965, n34966, n34967, n34968, n34969,
    n34970, n34971, n34972, n34973, n34974, n34975,
    n34976, n34977, n34978, n34979, n34980, n34981,
    n34982, n34983, n34984, n34985, n34986, n34987,
    n34988, n34989, n34990, n34991, n34992, n34993,
    n34994, n34995, n34996, n34997, n34998, n34999,
    n35000, n35001, n35002, n35003, n35004, n35005,
    n35006, n35007, n35008, n35009, n35010, n35011,
    n35012, n35013, n35014, n35015, n35016, n35017,
    n35018, n35019, n35020, n35021, n35022, n35023,
    n35024, n35025, n35026, n35027, n35028, n35029,
    n35030, n35031, n35032, n35033, n35034, n35035,
    n35036, n35037, n35038, n35039, n35040, n35041,
    n35042, n35043, n35044, n35045, n35046, n35047,
    n35048, n35049, n35050, n35051, n35052, n35053,
    n35054, n35055, n35056, n35057, n35058, n35059,
    n35060, n35061, n35062, n35063, n35064, n35065,
    n35066, n35067, n35068, n35069, n35070, n35071,
    n35072, n35073, n35074, n35075, n35076, n35077,
    n35078, n35079, n35080, n35081, n35082, n35083,
    n35084, n35085, n35086, n35087, n35088, n35089,
    n35090, n35091, n35092, n35093, n35094, n35095,
    n35096, n35097, n35098, n35099, n35100, n35101,
    n35102, n35103, n35104, n35105, n35106, n35107,
    n35108, n35109, n35110, n35111, n35112, n35113,
    n35114, n35115, n35116, n35117, n35118, n35119,
    n35120, n35121, n35122, n35123, n35124, n35125,
    n35126, n35127, n35128, n35129, n35130, n35131,
    n35132, n35133, n35134, n35135, n35136, n35137,
    n35138, n35139, n35140, n35141, n35142, n35143,
    n35144, n35145, n35146, n35147, n35148, n35149,
    n35150, n35151, n35152, n35153, n35154, n35155,
    n35156, n35157, n35158, n35159, n35160, n35161,
    n35162, n35163, n35164, n35165, n35166, n35167,
    n35168, n35169, n35170, n35171, n35172, n35173,
    n35174, n35175, n35176, n35177, n35178, n35179,
    n35180, n35181, n35182, n35183, n35184, n35185,
    n35186, n35187, n35188, n35189, n35190, n35191,
    n35192, n35193, n35194, n35195, n35196, n35197,
    n35198, n35199, n35200, n35201, n35202, n35203,
    n35204, n35205, n35206, n35207, n35208, n35209,
    n35210, n35211, n35212, n35213, n35214, n35215,
    n35216, n35217, n35218, n35219, n35220, n35221,
    n35222, n35223, n35224, n35225, n35226, n35227,
    n35228, n35229, n35230, n35231, n35232, n35233,
    n35234, n35235, n35236, n35237, n35238, n35239,
    n35240, n35241, n35242, n35243, n35244, n35245,
    n35246, n35247, n35248, n35249, n35250, n35251,
    n35252, n35253, n35254, n35255, n35256, n35257,
    n35258, n35259, n35260, n35261, n35262, n35263,
    n35264, n35265, n35266, n35267, n35268, n35269,
    n35270, n35271, n35272, n35273, n35274, n35275,
    n35276, n35277, n35278, n35279, n35280, n35281,
    n35282, n35283, n35284, n35285, n35286, n35287,
    n35288, n35289, n35290, n35291, n35292, n35293,
    n35294, n35295, n35296, n35297, n35298, n35299,
    n35300, n35301, n35302, n35303, n35304, n35305,
    n35306, n35307, n35308, n35309, n35310, n35311,
    n35312, n35313, n35314, n35315, n35316, n35317,
    n35318, n35319, n35320, n35321, n35322, n35323,
    n35324, n35325, n35326, n35327, n35328, n35329,
    n35330, n35331, n35332, n35333, n35334, n35335,
    n35336, n35337, n35338, n35339, n35340, n35341,
    n35342, n35343, n35344, n35345, n35346, n35347,
    n35348, n35349, n35350, n35351, n35352, n35353,
    n35354, n35355, n35356, n35357, n35358, n35359,
    n35360, n35361, n35362, n35363, n35364, n35365,
    n35366, n35367, n35368, n35369, n35370, n35371,
    n35372, n35373, n35374, n35375, n35376, n35377,
    n35378, n35379, n35380, n35381, n35382, n35383,
    n35384, n35385, n35386, n35387, n35388, n35389,
    n35390, n35391, n35392, n35393, n35394, n35395,
    n35396, n35397, n35398, n35399, n35400, n35401,
    n35402, n35403, n35404, n35405, n35406, n35407,
    n35408, n35409, n35410, n35411, n35412, n35413,
    n35414, n35415, n35416, n35417, n35418, n35419,
    n35420, n35421, n35422, n35423, n35424, n35425,
    n35426, n35427, n35428, n35429, n35430, n35431,
    n35432, n35433, n35434, n35435, n35436, n35437,
    n35438, n35439, n35440, n35441, n35442, n35443,
    n35444, n35445, n35446, n35447, n35448, n35449,
    n35450, n35451, n35452, n35453, n35454, n35455,
    n35456, n35457, n35458, n35459, n35460, n35461,
    n35462, n35463, n35464, n35465, n35466, n35467,
    n35468, n35469, n35470, n35471, n35472, n35473,
    n35474, n35475, n35476, n35477, n35478, n35479,
    n35480, n35481, n35482, n35483, n35484, n35485,
    n35486, n35487, n35488, n35489, n35490, n35491,
    n35492, n35493, n35494, n35495, n35496, n35497,
    n35498, n35499, n35500, n35501, n35502, n35503,
    n35504, n35505, n35506, n35507, n35508, n35509,
    n35510, n35511, n35512, n35513, n35514, n35515,
    n35516, n35517, n35518, n35519, n35520, n35521,
    n35522, n35523, n35524, n35525, n35526, n35527,
    n35528, n35529, n35530, n35531, n35532, n35533,
    n35534, n35535, n35536, n35537, n35538, n35539,
    n35540, n35541, n35542, n35543, n35544, n35545,
    n35546, n35547, n35548, n35549, n35550, n35551,
    n35552, n35553, n35554, n35555, n35556, n35557,
    n35558, n35559, n35560, n35561, n35562, n35563,
    n35564, n35565, n35566, n35567, n35568, n35569,
    n35570, n35571, n35572, n35573, n35574, n35575,
    n35576, n35577, n35578, n35579, n35580, n35581,
    n35582, n35583, n35584, n35585, n35586, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593,
    n35594, n35595, n35596, n35597, n35598, n35599,
    n35600, n35601, n35602, n35603, n35604, n35605,
    n35606, n35607, n35608, n35609, n35610, n35611,
    n35612, n35613, n35614, n35615, n35616, n35617,
    n35618, n35619, n35620, n35621, n35622, n35623,
    n35624, n35625, n35626, n35627, n35628, n35629,
    n35630, n35631, n35632, n35633, n35634, n35635,
    n35636, n35637, n35638, n35639, n35640, n35641,
    n35642, n35643, n35644, n35645, n35646, n35647,
    n35648, n35649, n35650, n35651, n35652, n35653,
    n35654, n35655, n35656, n35657, n35658, n35659,
    n35660, n35661, n35662, n35663, n35664, n35665,
    n35666, n35667, n35668, n35669, n35670, n35671,
    n35672, n35673, n35674, n35675, n35676, n35677,
    n35678, n35679, n35680, n35681, n35682, n35683,
    n35684, n35685, n35686, n35687, n35688, n35689,
    n35690, n35691, n35692, n35693, n35694, n35695,
    n35696, n35697, n35698, n35699, n35700, n35701,
    n35702, n35703, n35704, n35705, n35706, n35707,
    n35708, n35709, n35710, n35711, n35712, n35713,
    n35714, n35715, n35716, n35717, n35718, n35719,
    n35720, n35721, n35722, n35723, n35724, n35725,
    n35726, n35727, n35728, n35729, n35730, n35731,
    n35732, n35733, n35734, n35735, n35736, n35737,
    n35738, n35739, n35740, n35741, n35742, n35743,
    n35744, n35745, n35746, n35747, n35748, n35749,
    n35750, n35751, n35752, n35753, n35754, n35755,
    n35756, n35757, n35758, n35759, n35760, n35761,
    n35762, n35763, n35764, n35765, n35766, n35767,
    n35768, n35769, n35770, n35771, n35772, n35773,
    n35774, n35775, n35776, n35777, n35778, n35779,
    n35780, n35781, n35782, n35783, n35784, n35785,
    n35786, n35787, n35788, n35789, n35790, n35791,
    n35792, n35793, n35794, n35795, n35796, n35797,
    n35798, n35799, n35800, n35801, n35802, n35803,
    n35804, n35805, n35806, n35807, n35808, n35809,
    n35810, n35811, n35812, n35813, n35814, n35815,
    n35816, n35817;
  assign n193 = ~pi126  & ~pi127 ;
  assign n194 = pi126  & pi127 ;
  assign n195 = ~pi124  & ~pi125 ;
  assign n196 = ~pi126  & ~n195;
  assign n197 = ~n194 & ~n196;
  assign n198 = ~pi124  & ~n197;
  assign n199 = pi125  & ~n198;
  assign n200 = n195 & ~n197;
  assign n201 = n194 & n195;
  assign n202 = ~n199 & ~n31780;
  assign n203 = pi124  & ~n197;
  assign n204 = ~pi122  & ~pi123 ;
  assign n205 = ~pi124  & n204;
  assign n206 = ~n203 & ~n205;
  assign n207 = n202 & ~n206;
  assign n208 = n193 & ~n207;
  assign n209 = ~n202 & n206;
  assign n210 = pi126  & n195;
  assign n211 = pi127  & ~n196;
  assign n212 = ~n210 & n211;
  assign n213 = ~n209 & ~n212;
  assign n214 = ~n208 & n213;
  assign n215 = pi122  & ~n214;
  assign n216 = ~pi120  & ~pi121 ;
  assign n217 = ~pi122  & n216;
  assign n218 = ~n194 & ~n217;
  assign n219 = ~n196 & n218;
  assign n220 = ~pi122  & ~n216;
  assign n221 = pi122  & n214;
  assign n222 = ~n220 & ~n221;
  assign n223 = ~n215 & ~n217;
  assign n224 = n197 & ~n31781;
  assign n225 = ~n215 & n219;
  assign n226 = ~n197 & n31781;
  assign n227 = ~pi122  & ~n214;
  assign n228 = ~pi123  & n227;
  assign n229 = n204 & ~n214;
  assign n230 = pi123  & ~n227;
  assign n231 = ~n31783 & ~n230;
  assign n232 = ~n226 & ~n231;
  assign n233 = ~n31782 & n231;
  assign n234 = ~n226 & ~n233;
  assign n235 = ~n31782 & ~n232;
  assign n236 = ~n197 & ~n212;
  assign n237 = ~n209 & n236;
  assign n238 = ~n197 & n214;
  assign n239 = ~n208 & n237;
  assign n240 = ~n31783 & ~n31785;
  assign n241 = pi124  & ~n240;
  assign n242 = ~pi124  & ~n31785;
  assign n243 = ~pi124  & n240;
  assign n244 = ~n31783 & n242;
  assign n245 = ~n241 & ~n31786;
  assign n246 = n207 & ~n214;
  assign n247 = n207 & n212;
  assign n248 = ~n209 & ~n31787;
  assign n249 = ~n245 & n248;
  assign n250 = ~n31784 & ~n245;
  assign n251 = n248 & n250;
  assign n252 = ~n31784 & n249;
  assign n253 = n193 & ~n31788;
  assign n254 = n31784 & n245;
  assign n255 = ~n193 & ~n207;
  assign n256 = ~n209 & n255;
  assign n257 = n206 & ~n212;
  assign n258 = n202 & ~n214;
  assign n259 = n206 & ~n258;
  assign n260 = n255 & ~n259;
  assign n261 = n256 & ~n257;
  assign n262 = ~n254 & ~n31789;
  assign n263 = ~n253 & n262;
  assign n264 = pi120  & ~n263;
  assign n265 = ~pi118  & ~pi119 ;
  assign n266 = ~pi120  & n265;
  assign n267 = ~n264 & ~n266;
  assign n268 = ~n214 & ~n267;
  assign n269 = ~pi120  & ~n263;
  assign n270 = pi121  & ~n269;
  assign n271 = ~pi121  & n269;
  assign n272 = n216 & ~n263;
  assign n273 = ~n270 & ~n31790;
  assign n274 = ~n212 & ~n266;
  assign n275 = ~n209 & n274;
  assign n276 = ~n208 & n275;
  assign n277 = n214 & n267;
  assign n278 = ~n264 & n276;
  assign n279 = n273 & ~n31791;
  assign n280 = ~n268 & ~n279;
  assign n281 = ~n197 & ~n280;
  assign n282 = n197 & ~n268;
  assign n283 = ~n279 & n282;
  assign n284 = ~n214 & ~n31789;
  assign n285 = ~n214 & ~n256;
  assign n286 = ~n254 & n31792;
  assign n287 = ~n253 & n286;
  assign n288 = ~n31790 & ~n287;
  assign n289 = pi122  & ~n288;
  assign n290 = ~pi122  & ~n287;
  assign n291 = ~pi122  & n288;
  assign n292 = ~n31790 & n290;
  assign n293 = ~n289 & ~n31793;
  assign n294 = ~n283 & ~n293;
  assign n295 = ~n281 & ~n294;
  assign n296 = ~n31782 & ~n226;
  assign n297 = ~n263 & n296;
  assign n298 = n231 & ~n297;
  assign n299 = ~n231 & n296;
  assign n300 = ~n231 & n297;
  assign n301 = ~n263 & n299;
  assign n302 = ~n298 & ~n31794;
  assign n303 = n250 & ~n263;
  assign n304 = ~n254 & ~n303;
  assign n305 = ~n302 & n304;
  assign n306 = ~n295 & n305;
  assign n307 = n193 & ~n306;
  assign n308 = ~n281 & n302;
  assign n309 = ~n294 & n308;
  assign n310 = n295 & n302;
  assign n311 = ~n245 & n263;
  assign n312 = ~n193 & ~n250;
  assign n313 = ~n254 & n312;
  assign n314 = ~n263 & ~n313;
  assign n315 = n31784 & ~n263;
  assign n316 = ~n245 & ~n315;
  assign n317 = ~n193 & ~n254;
  assign n318 = ~n316 & n317;
  assign n319 = ~n311 & ~n314;
  assign n320 = ~n31795 & ~n31796;
  assign n321 = ~n307 & n320;
  assign n322 = pi118  & ~n321;
  assign n323 = ~pi116  & ~pi117 ;
  assign n324 = ~pi118  & n323;
  assign n325 = ~n322 & ~n324;
  assign n326 = ~n263 & ~n325;
  assign n327 = ~n202 & ~n212;
  assign n328 = ~n209 & n327;
  assign n329 = ~n202 & n214;
  assign n330 = ~n208 & n328;
  assign n331 = ~n324 & ~n31797;
  assign n332 = ~n31789 & n331;
  assign n333 = ~n254 & n332;
  assign n334 = ~n253 & n333;
  assign n335 = n263 & n325;
  assign n336 = ~n322 & n334;
  assign n337 = ~pi118  & ~n321;
  assign n338 = pi119  & ~n337;
  assign n339 = ~pi119  & n337;
  assign n340 = n265 & ~n321;
  assign n341 = ~n338 & ~n31799;
  assign n342 = ~n31798 & n341;
  assign n343 = ~n326 & ~n342;
  assign n344 = ~n214 & ~n343;
  assign n345 = ~n31795 & n314;
  assign n346 = ~n307 & n345;
  assign n347 = ~n31799 & ~n346;
  assign n348 = pi120  & ~n347;
  assign n349 = ~pi120  & ~n346;
  assign n350 = ~pi120  & n347;
  assign n351 = ~n31799 & n349;
  assign n352 = ~n348 & ~n31800;
  assign n353 = n214 & ~n326;
  assign n354 = n214 & n343;
  assign n355 = ~n342 & n353;
  assign n356 = ~n352 & ~n31801;
  assign n357 = ~n344 & ~n356;
  assign n358 = ~n197 & ~n357;
  assign n359 = n197 & ~n344;
  assign n360 = ~n356 & n359;
  assign n361 = ~n268 & ~n31791;
  assign n362 = ~n321 & n361;
  assign n363 = n273 & ~n362;
  assign n364 = ~n273 & ~n31791;
  assign n365 = ~n268 & n364;
  assign n366 = ~n273 & n362;
  assign n367 = ~n321 & n365;
  assign n368 = ~n363 & ~n31802;
  assign n369 = ~n360 & ~n368;
  assign n370 = ~n358 & ~n369;
  assign n371 = ~n281 & ~n283;
  assign n372 = ~n321 & n371;
  assign n373 = ~n293 & ~n372;
  assign n374 = ~n283 & n293;
  assign n375 = ~n281 & n374;
  assign n376 = n293 & n372;
  assign n377 = ~n321 & n375;
  assign n378 = ~n373 & ~n31803;
  assign n379 = ~n295 & ~n302;
  assign n380 = ~n321 & n379;
  assign n381 = ~n31795 & ~n380;
  assign n382 = ~n378 & n381;
  assign n383 = ~n370 & n382;
  assign n384 = n193 & ~n383;
  assign n385 = ~n358 & n378;
  assign n386 = n370 & n378;
  assign n387 = ~n369 & n385;
  assign n388 = n295 & ~n321;
  assign n389 = ~n302 & ~n388;
  assign n390 = ~n193 & ~n31795;
  assign n391 = ~n389 & n390;
  assign n392 = ~n31804 & ~n391;
  assign n393 = ~n384 & n392;
  assign n394 = pi116  & ~n393;
  assign n395 = ~pi114  & ~pi115 ;
  assign n396 = ~pi116  & n395;
  assign n397 = ~n394 & ~n396;
  assign n398 = ~n321 & ~n397;
  assign n399 = ~pi116  & ~n393;
  assign n400 = pi117  & ~n399;
  assign n401 = ~pi117  & n399;
  assign n402 = n323 & ~n393;
  assign n403 = ~n400 & ~n31805;
  assign n404 = ~n31786 & ~n31797;
  assign n405 = ~n241 & n404;
  assign n406 = ~n31789 & n405;
  assign n407 = ~n254 & n406;
  assign n408 = ~n253 & n407;
  assign n409 = ~n396 & ~n408;
  assign n410 = ~n31796 & n409;
  assign n411 = ~n31795 & n410;
  assign n412 = ~n307 & n411;
  assign n413 = n321 & n397;
  assign n414 = ~n394 & n412;
  assign n415 = n403 & ~n31806;
  assign n416 = ~n398 & ~n415;
  assign n417 = ~n263 & ~n416;
  assign n418 = n263 & ~n398;
  assign n419 = ~n415 & n418;
  assign n420 = ~n321 & ~n391;
  assign n421 = ~n31804 & n420;
  assign n422 = ~n384 & n421;
  assign n423 = ~n31805 & ~n422;
  assign n424 = pi118  & ~n423;
  assign n425 = ~pi118  & ~n422;
  assign n426 = ~pi118  & n423;
  assign n427 = ~n31805 & n425;
  assign n428 = ~n424 & ~n31807;
  assign n429 = ~n419 & ~n428;
  assign n430 = ~n417 & ~n429;
  assign n431 = ~n214 & ~n430;
  assign n432 = n214 & ~n417;
  assign n433 = ~n429 & n432;
  assign n434 = n214 & n430;
  assign n435 = ~n326 & ~n31798;
  assign n436 = ~n393 & n435;
  assign n437 = n341 & ~n436;
  assign n438 = ~n341 & n435;
  assign n439 = ~n341 & n436;
  assign n440 = ~n393 & n438;
  assign n441 = ~n437 & ~n31809;
  assign n442 = ~n31808 & ~n441;
  assign n443 = ~n431 & ~n442;
  assign n444 = ~n197 & ~n443;
  assign n445 = n197 & ~n431;
  assign n446 = ~n442 & n445;
  assign n447 = ~n344 & ~n31801;
  assign n448 = ~n344 & ~n393;
  assign n449 = ~n31801 & n448;
  assign n450 = ~n393 & n447;
  assign n451 = n352 & ~n31810;
  assign n452 = n356 & n448;
  assign n453 = n352 & ~n31801;
  assign n454 = ~n344 & n453;
  assign n455 = ~n393 & n454;
  assign n456 = ~n352 & ~n31810;
  assign n457 = ~n455 & ~n456;
  assign n458 = ~n451 & ~n452;
  assign n459 = ~n446 & ~n31811;
  assign n460 = ~n444 & ~n459;
  assign n461 = ~n358 & ~n360;
  assign n462 = ~n393 & n461;
  assign n463 = ~n368 & ~n462;
  assign n464 = ~n358 & n368;
  assign n465 = ~n360 & n464;
  assign n466 = n368 & n462;
  assign n467 = ~n393 & n465;
  assign n468 = n368 & ~n462;
  assign n469 = ~n368 & n462;
  assign n470 = ~n468 & ~n469;
  assign n471 = ~n463 & ~n31812;
  assign n472 = ~n370 & ~n378;
  assign n473 = ~n378 & ~n393;
  assign n474 = ~n370 & n473;
  assign n475 = ~n393 & n472;
  assign n476 = ~n31804 & ~n31814;
  assign n477 = n31813 & n476;
  assign n478 = ~n460 & n477;
  assign n479 = n193 & ~n478;
  assign n480 = ~n444 & ~n31813;
  assign n481 = ~n459 & n480;
  assign n482 = n460 & ~n31813;
  assign n483 = n370 & ~n473;
  assign n484 = ~n193 & ~n472;
  assign n485 = ~n483 & n484;
  assign n486 = ~n31815 & ~n485;
  assign n487 = ~n479 & n486;
  assign n488 = pi114  & ~n487;
  assign n489 = ~pi112  & ~pi113 ;
  assign n490 = ~pi114  & n489;
  assign n491 = ~n488 & ~n490;
  assign n492 = ~n393 & ~n491;
  assign n493 = ~n31794 & ~n408;
  assign n494 = ~n298 & n493;
  assign n495 = ~n31796 & n494;
  assign n496 = ~n31795 & n495;
  assign n497 = n302 & n321;
  assign n498 = ~n307 & n496;
  assign n499 = ~n490 & ~n31816;
  assign n500 = ~n391 & n499;
  assign n501 = ~n31804 & n500;
  assign n502 = ~n384 & n501;
  assign n503 = n393 & n491;
  assign n504 = ~n488 & n502;
  assign n505 = ~pi114  & ~n487;
  assign n506 = pi115  & ~n505;
  assign n507 = ~pi115  & n505;
  assign n508 = n395 & ~n487;
  assign n509 = ~n506 & ~n31818;
  assign n510 = ~n31817 & n509;
  assign n511 = ~n492 & ~n510;
  assign n512 = ~n321 & ~n511;
  assign n513 = ~n393 & ~n485;
  assign n514 = ~n31815 & n513;
  assign n515 = ~n479 & n514;
  assign n516 = ~n31818 & ~n515;
  assign n517 = pi116  & ~n516;
  assign n518 = ~pi116  & ~n515;
  assign n519 = ~pi116  & n516;
  assign n520 = ~n31818 & n518;
  assign n521 = ~n517 & ~n31819;
  assign n522 = n321 & ~n492;
  assign n523 = n321 & n511;
  assign n524 = ~n510 & n522;
  assign n525 = ~n521 & ~n31820;
  assign n526 = ~n512 & ~n525;
  assign n527 = ~n263 & ~n526;
  assign n528 = n263 & ~n512;
  assign n529 = ~n525 & n528;
  assign n530 = ~n398 & ~n31806;
  assign n531 = ~n487 & n530;
  assign n532 = n403 & ~n531;
  assign n533 = ~n403 & n530;
  assign n534 = ~n403 & n531;
  assign n535 = ~n487 & n533;
  assign n536 = ~n532 & ~n31821;
  assign n537 = ~n529 & ~n536;
  assign n538 = ~n527 & ~n537;
  assign n539 = ~n214 & ~n538;
  assign n540 = ~n417 & ~n419;
  assign n541 = ~n487 & n540;
  assign n542 = ~n428 & ~n541;
  assign n543 = ~n419 & n428;
  assign n544 = ~n417 & n543;
  assign n545 = n428 & n541;
  assign n546 = ~n487 & n544;
  assign n547 = ~n542 & ~n31822;
  assign n548 = n214 & ~n527;
  assign n549 = n214 & n538;
  assign n550 = ~n537 & n548;
  assign n551 = ~n547 & ~n31823;
  assign n552 = ~n539 & ~n551;
  assign n553 = ~n197 & ~n552;
  assign n554 = n197 & ~n539;
  assign n555 = ~n551 & n554;
  assign n556 = ~n431 & ~n31808;
  assign n557 = ~n487 & n556;
  assign n558 = ~n441 & ~n557;
  assign n559 = ~n431 & n441;
  assign n560 = ~n31808 & n559;
  assign n561 = n441 & n557;
  assign n562 = ~n487 & n560;
  assign n563 = n441 & ~n557;
  assign n564 = ~n441 & n557;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~n558 & ~n31824;
  assign n567 = ~n555 & n31825;
  assign n568 = ~n553 & ~n567;
  assign n569 = ~n444 & ~n446;
  assign n570 = ~n487 & n569;
  assign n571 = ~n31811 & ~n570;
  assign n572 = ~n446 & n31811;
  assign n573 = ~n444 & n572;
  assign n574 = n31811 & n570;
  assign n575 = ~n487 & n573;
  assign n576 = ~n571 & ~n31826;
  assign n577 = ~n460 & n31813;
  assign n578 = n31813 & ~n487;
  assign n579 = ~n460 & n578;
  assign n580 = ~n487 & n577;
  assign n581 = ~n31815 & ~n31827;
  assign n582 = ~n576 & n581;
  assign n583 = ~n568 & n582;
  assign n584 = n193 & ~n583;
  assign n585 = ~n553 & n576;
  assign n586 = n568 & n576;
  assign n587 = ~n567 & n585;
  assign n588 = n460 & ~n578;
  assign n589 = ~n193 & ~n577;
  assign n590 = ~n588 & n589;
  assign n591 = ~n31828 & ~n590;
  assign n592 = ~n584 & n591;
  assign n593 = pi112  & ~n592;
  assign n594 = ~pi110  & ~pi111 ;
  assign n595 = ~pi112  & n594;
  assign n596 = ~n593 & ~n595;
  assign n597 = ~n487 & ~n596;
  assign n598 = ~pi112  & ~n592;
  assign n599 = pi113  & ~n598;
  assign n600 = ~pi113  & n598;
  assign n601 = n489 & ~n592;
  assign n602 = ~n599 & ~n31829;
  assign n603 = ~n31803 & ~n31816;
  assign n604 = ~n373 & n603;
  assign n605 = ~n391 & n604;
  assign n606 = ~n31804 & n605;
  assign n607 = n378 & n393;
  assign n608 = ~n384 & n606;
  assign n609 = ~n595 & ~n31830;
  assign n610 = ~n485 & n609;
  assign n611 = ~n31815 & n610;
  assign n612 = ~n479 & n611;
  assign n613 = n487 & n596;
  assign n614 = ~n593 & n612;
  assign n615 = n602 & ~n31831;
  assign n616 = ~n597 & ~n615;
  assign n617 = ~n393 & ~n616;
  assign n618 = n393 & ~n597;
  assign n619 = ~n615 & n618;
  assign n620 = ~n487 & ~n590;
  assign n621 = ~n31828 & n620;
  assign n622 = ~n584 & n621;
  assign n623 = ~n31829 & ~n622;
  assign n624 = pi114  & ~n623;
  assign n625 = ~pi114  & ~n622;
  assign n626 = ~pi114  & n623;
  assign n627 = ~n31829 & n625;
  assign n628 = ~n624 & ~n31832;
  assign n629 = ~n619 & ~n628;
  assign n630 = ~n617 & ~n629;
  assign n631 = ~n321 & ~n630;
  assign n632 = n321 & ~n617;
  assign n633 = ~n629 & n632;
  assign n634 = n321 & n630;
  assign n635 = ~n492 & ~n31817;
  assign n636 = ~n592 & n635;
  assign n637 = n509 & ~n636;
  assign n638 = ~n509 & n635;
  assign n639 = ~n509 & n636;
  assign n640 = ~n592 & n638;
  assign n641 = ~n637 & ~n31834;
  assign n642 = ~n31833 & ~n641;
  assign n643 = ~n631 & ~n642;
  assign n644 = ~n263 & ~n643;
  assign n645 = n263 & ~n631;
  assign n646 = ~n642 & n645;
  assign n647 = ~n512 & ~n31820;
  assign n648 = ~n512 & ~n592;
  assign n649 = ~n31820 & n648;
  assign n650 = ~n592 & n647;
  assign n651 = n521 & ~n31835;
  assign n652 = n525 & n648;
  assign n653 = n521 & ~n31820;
  assign n654 = ~n512 & n653;
  assign n655 = ~n592 & n654;
  assign n656 = ~n521 & ~n31835;
  assign n657 = ~n655 & ~n656;
  assign n658 = ~n651 & ~n652;
  assign n659 = ~n646 & ~n31836;
  assign n660 = ~n644 & ~n659;
  assign n661 = ~n214 & ~n660;
  assign n662 = n214 & ~n644;
  assign n663 = ~n659 & n662;
  assign n664 = n214 & n660;
  assign n665 = ~n527 & ~n529;
  assign n666 = ~n592 & n665;
  assign n667 = ~n536 & ~n666;
  assign n668 = ~n527 & n536;
  assign n669 = ~n529 & n668;
  assign n670 = n536 & n666;
  assign n671 = ~n592 & n669;
  assign n672 = n536 & ~n666;
  assign n673 = ~n536 & n666;
  assign n674 = ~n672 & ~n673;
  assign n675 = ~n667 & ~n31838;
  assign n676 = ~n31837 & n31839;
  assign n677 = ~n661 & ~n676;
  assign n678 = ~n197 & ~n677;
  assign n679 = n197 & ~n661;
  assign n680 = ~n676 & n679;
  assign n681 = ~n539 & ~n31823;
  assign n682 = ~n539 & ~n592;
  assign n683 = ~n31823 & n682;
  assign n684 = ~n592 & n681;
  assign n685 = n547 & ~n31840;
  assign n686 = n551 & n682;
  assign n687 = n547 & ~n31823;
  assign n688 = ~n539 & n687;
  assign n689 = ~n592 & n688;
  assign n690 = ~n547 & ~n31840;
  assign n691 = ~n689 & ~n690;
  assign n692 = ~n685 & ~n686;
  assign n693 = ~n680 & ~n31841;
  assign n694 = ~n678 & ~n693;
  assign n695 = ~n553 & ~n555;
  assign n696 = ~n592 & n695;
  assign n697 = ~n31825 & ~n696;
  assign n698 = n31825 & n696;
  assign n699 = ~n553 & ~n31825;
  assign n700 = ~n555 & n699;
  assign n701 = ~n592 & n700;
  assign n702 = n31825 & ~n696;
  assign n703 = ~n701 & ~n702;
  assign n704 = ~n697 & ~n698;
  assign n705 = ~n568 & ~n576;
  assign n706 = ~n576 & ~n592;
  assign n707 = ~n568 & n706;
  assign n708 = ~n592 & n705;
  assign n709 = ~n31828 & ~n31843;
  assign n710 = ~n31842 & n709;
  assign n711 = ~n694 & n710;
  assign n712 = n193 & ~n711;
  assign n713 = ~n678 & n31842;
  assign n714 = ~n693 & n713;
  assign n715 = n694 & n31842;
  assign n716 = n568 & ~n706;
  assign n717 = ~n193 & ~n705;
  assign n718 = ~n716 & n717;
  assign n719 = ~n31844 & ~n718;
  assign n720 = ~n712 & n719;
  assign n721 = pi110  & ~n720;
  assign n722 = ~pi108  & ~pi109 ;
  assign n723 = ~pi110  & n722;
  assign n724 = ~n721 & ~n723;
  assign n725 = ~n592 & ~n724;
  assign n726 = ~n31812 & ~n31830;
  assign n727 = ~n463 & n726;
  assign n728 = ~n485 & n727;
  assign n729 = ~n31815 & n728;
  assign n730 = ~n31813 & n487;
  assign n731 = ~n479 & n729;
  assign n732 = ~n723 & ~n31845;
  assign n733 = ~n590 & n732;
  assign n734 = ~n31828 & n733;
  assign n735 = ~n584 & n734;
  assign n736 = n592 & n724;
  assign n737 = ~n721 & n735;
  assign n738 = ~pi110  & ~n720;
  assign n739 = pi111  & ~n738;
  assign n740 = ~pi111  & n738;
  assign n741 = n594 & ~n720;
  assign n742 = ~n739 & ~n31847;
  assign n743 = ~n31846 & n742;
  assign n744 = ~n725 & ~n743;
  assign n745 = ~n487 & ~n744;
  assign n746 = ~n592 & ~n718;
  assign n747 = ~n31844 & n746;
  assign n748 = ~n712 & n747;
  assign n749 = ~n31847 & ~n748;
  assign n750 = pi112  & ~n749;
  assign n751 = ~pi112  & ~n748;
  assign n752 = ~pi112  & n749;
  assign n753 = ~n31847 & n751;
  assign n754 = ~n750 & ~n31848;
  assign n755 = n487 & ~n725;
  assign n756 = n487 & n744;
  assign n757 = ~n743 & n755;
  assign n758 = ~n754 & ~n31849;
  assign n759 = ~n745 & ~n758;
  assign n760 = ~n393 & ~n759;
  assign n761 = n393 & ~n745;
  assign n762 = ~n758 & n761;
  assign n763 = ~n597 & ~n31831;
  assign n764 = ~n720 & n763;
  assign n765 = n602 & ~n764;
  assign n766 = ~n602 & ~n31831;
  assign n767 = ~n597 & n766;
  assign n768 = ~n602 & n764;
  assign n769 = ~n720 & n767;
  assign n770 = ~n765 & ~n31850;
  assign n771 = ~n762 & ~n770;
  assign n772 = ~n760 & ~n771;
  assign n773 = ~n321 & ~n772;
  assign n774 = ~n617 & ~n619;
  assign n775 = ~n720 & n774;
  assign n776 = ~n628 & ~n775;
  assign n777 = ~n619 & n628;
  assign n778 = ~n617 & n777;
  assign n779 = n628 & n775;
  assign n780 = ~n720 & n778;
  assign n781 = ~n776 & ~n31851;
  assign n782 = n321 & ~n760;
  assign n783 = n321 & n772;
  assign n784 = ~n771 & n782;
  assign n785 = ~n781 & ~n31852;
  assign n786 = ~n773 & ~n785;
  assign n787 = ~n263 & ~n786;
  assign n788 = n263 & ~n773;
  assign n789 = ~n785 & n788;
  assign n790 = ~n631 & ~n31833;
  assign n791 = ~n720 & n790;
  assign n792 = ~n641 & ~n791;
  assign n793 = ~n631 & n641;
  assign n794 = ~n31833 & n793;
  assign n795 = n641 & n791;
  assign n796 = ~n720 & n794;
  assign n797 = n641 & ~n791;
  assign n798 = ~n641 & n791;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~n792 & ~n31853;
  assign n801 = ~n789 & n31854;
  assign n802 = ~n787 & ~n801;
  assign n803 = ~n214 & ~n802;
  assign n804 = ~n644 & ~n646;
  assign n805 = ~n720 & n804;
  assign n806 = ~n31836 & ~n805;
  assign n807 = ~n646 & n31836;
  assign n808 = ~n644 & n807;
  assign n809 = n31836 & n805;
  assign n810 = ~n720 & n808;
  assign n811 = ~n806 & ~n31855;
  assign n812 = n214 & ~n787;
  assign n813 = n214 & n802;
  assign n814 = ~n801 & n812;
  assign n815 = ~n811 & ~n31856;
  assign n816 = ~n803 & ~n815;
  assign n817 = ~n197 & ~n816;
  assign n818 = n197 & ~n803;
  assign n819 = ~n815 & n818;
  assign n820 = ~n661 & ~n31837;
  assign n821 = ~n720 & n820;
  assign n822 = ~n31839 & ~n821;
  assign n823 = n31839 & n821;
  assign n824 = ~n661 & ~n31839;
  assign n825 = ~n31837 & n824;
  assign n826 = ~n720 & n825;
  assign n827 = n31839 & ~n821;
  assign n828 = ~n826 & ~n827;
  assign n829 = ~n822 & ~n823;
  assign n830 = ~n819 & ~n31857;
  assign n831 = ~n817 & ~n830;
  assign n832 = ~n678 & ~n680;
  assign n833 = ~n720 & n832;
  assign n834 = ~n31841 & ~n833;
  assign n835 = ~n680 & n31841;
  assign n836 = ~n678 & n835;
  assign n837 = n31841 & n833;
  assign n838 = ~n720 & n836;
  assign n839 = ~n834 & ~n31858;
  assign n840 = ~n694 & ~n31842;
  assign n841 = ~n31842 & ~n720;
  assign n842 = ~n694 & n841;
  assign n843 = ~n720 & n840;
  assign n844 = ~n31844 & ~n31859;
  assign n845 = ~n839 & n844;
  assign n846 = ~n831 & n845;
  assign n847 = n193 & ~n846;
  assign n848 = ~n817 & n839;
  assign n849 = n831 & n839;
  assign n850 = ~n830 & n848;
  assign n851 = n694 & ~n841;
  assign n852 = ~n193 & ~n840;
  assign n853 = ~n851 & n852;
  assign n854 = ~n31860 & ~n853;
  assign n855 = ~n847 & n854;
  assign n856 = pi108  & ~n855;
  assign n857 = ~pi106  & ~pi107 ;
  assign n858 = ~pi108  & n857;
  assign n859 = ~n856 & ~n858;
  assign n860 = ~n720 & ~n859;
  assign n861 = ~pi108  & ~n855;
  assign n862 = pi109  & ~n861;
  assign n863 = ~pi109  & n861;
  assign n864 = n722 & ~n855;
  assign n865 = ~n862 & ~n31861;
  assign n866 = ~n31826 & ~n31845;
  assign n867 = ~n571 & n866;
  assign n868 = ~n590 & n867;
  assign n869 = ~n31828 & n868;
  assign n870 = n576 & n592;
  assign n871 = ~n584 & n869;
  assign n872 = ~n858 & ~n31862;
  assign n873 = ~n718 & n872;
  assign n874 = ~n31844 & n873;
  assign n875 = ~n712 & n874;
  assign n876 = n720 & n859;
  assign n877 = ~n856 & n875;
  assign n878 = n865 & ~n31863;
  assign n879 = ~n860 & ~n878;
  assign n880 = ~n592 & ~n879;
  assign n881 = n592 & ~n860;
  assign n882 = ~n878 & n881;
  assign n883 = ~n720 & ~n853;
  assign n884 = ~n31860 & n883;
  assign n885 = ~n847 & n884;
  assign n886 = ~n31861 & ~n885;
  assign n887 = pi110  & ~n886;
  assign n888 = ~pi110  & ~n885;
  assign n889 = ~pi110  & n886;
  assign n890 = ~n31861 & n888;
  assign n891 = ~n887 & ~n31864;
  assign n892 = ~n882 & ~n891;
  assign n893 = ~n880 & ~n892;
  assign n894 = ~n487 & ~n893;
  assign n895 = n487 & ~n880;
  assign n896 = ~n892 & n895;
  assign n897 = n487 & n893;
  assign n898 = ~n725 & ~n31846;
  assign n899 = ~n855 & n898;
  assign n900 = n742 & ~n899;
  assign n901 = ~n742 & n898;
  assign n902 = ~n742 & n899;
  assign n903 = ~n855 & n901;
  assign n904 = ~n900 & ~n31866;
  assign n905 = ~n31865 & ~n904;
  assign n906 = ~n894 & ~n905;
  assign n907 = ~n393 & ~n906;
  assign n908 = n393 & ~n894;
  assign n909 = ~n905 & n908;
  assign n910 = ~n745 & ~n31849;
  assign n911 = ~n745 & ~n855;
  assign n912 = ~n31849 & n911;
  assign n913 = ~n855 & n910;
  assign n914 = n754 & ~n31867;
  assign n915 = n758 & n911;
  assign n916 = n754 & ~n31849;
  assign n917 = ~n745 & n916;
  assign n918 = ~n855 & n917;
  assign n919 = ~n754 & ~n31867;
  assign n920 = ~n918 & ~n919;
  assign n921 = ~n914 & ~n915;
  assign n922 = ~n909 & ~n31868;
  assign n923 = ~n907 & ~n922;
  assign n924 = ~n321 & ~n923;
  assign n925 = n321 & ~n907;
  assign n926 = ~n922 & n925;
  assign n927 = n321 & n923;
  assign n928 = ~n760 & ~n762;
  assign n929 = ~n855 & n928;
  assign n930 = ~n770 & ~n929;
  assign n931 = ~n760 & n770;
  assign n932 = ~n762 & n931;
  assign n933 = n770 & n929;
  assign n934 = ~n855 & n932;
  assign n935 = n770 & ~n929;
  assign n936 = ~n770 & n929;
  assign n937 = ~n935 & ~n936;
  assign n938 = ~n930 & ~n31870;
  assign n939 = ~n31869 & n31871;
  assign n940 = ~n924 & ~n939;
  assign n941 = ~n263 & ~n940;
  assign n942 = n263 & ~n924;
  assign n943 = ~n939 & n942;
  assign n944 = ~n773 & ~n31852;
  assign n945 = ~n773 & ~n855;
  assign n946 = ~n31852 & n945;
  assign n947 = ~n855 & n944;
  assign n948 = n781 & ~n31872;
  assign n949 = n785 & n945;
  assign n950 = n781 & ~n31852;
  assign n951 = ~n773 & n950;
  assign n952 = ~n855 & n951;
  assign n953 = ~n781 & ~n31872;
  assign n954 = ~n952 & ~n953;
  assign n955 = ~n948 & ~n949;
  assign n956 = ~n943 & ~n31873;
  assign n957 = ~n941 & ~n956;
  assign n958 = ~n214 & ~n957;
  assign n959 = n214 & ~n941;
  assign n960 = ~n956 & n959;
  assign n961 = n214 & n957;
  assign n962 = ~n787 & ~n789;
  assign n963 = ~n855 & n962;
  assign n964 = ~n31854 & ~n963;
  assign n965 = n31854 & n963;
  assign n966 = ~n787 & ~n31854;
  assign n967 = ~n789 & n966;
  assign n968 = ~n855 & n967;
  assign n969 = n31854 & ~n963;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~n964 & ~n965;
  assign n972 = ~n31874 & ~n31875;
  assign n973 = ~n958 & ~n972;
  assign n974 = ~n197 & ~n973;
  assign n975 = n197 & ~n958;
  assign n976 = ~n972 & n975;
  assign n977 = ~n803 & ~n31856;
  assign n978 = ~n803 & ~n855;
  assign n979 = ~n31856 & n978;
  assign n980 = ~n855 & n977;
  assign n981 = n811 & ~n31876;
  assign n982 = n815 & n978;
  assign n983 = n811 & ~n31856;
  assign n984 = ~n803 & n983;
  assign n985 = ~n855 & n984;
  assign n986 = ~n811 & ~n31876;
  assign n987 = ~n985 & ~n986;
  assign n988 = ~n981 & ~n982;
  assign n989 = ~n976 & ~n31877;
  assign n990 = ~n974 & ~n989;
  assign n991 = ~n817 & ~n819;
  assign n992 = ~n855 & n991;
  assign n993 = ~n31857 & n992;
  assign n994 = n31857 & ~n992;
  assign n995 = ~n817 & n31857;
  assign n996 = ~n819 & n995;
  assign n997 = ~n855 & n996;
  assign n998 = ~n31857 & ~n992;
  assign n999 = ~n997 & ~n998;
  assign n1000 = ~n993 & ~n994;
  assign n1001 = ~n831 & ~n839;
  assign n1002 = ~n839 & ~n855;
  assign n1003 = ~n831 & n1002;
  assign n1004 = ~n855 & n1001;
  assign n1005 = ~n31860 & ~n31879;
  assign n1006 = ~n31878 & n1005;
  assign n1007 = ~n990 & n1006;
  assign n1008 = n193 & ~n1007;
  assign n1009 = ~n974 & n31878;
  assign n1010 = ~n989 & n1009;
  assign n1011 = n990 & n31878;
  assign n1012 = n831 & ~n1002;
  assign n1013 = ~n193 & ~n1001;
  assign n1014 = ~n1012 & n1013;
  assign n1015 = ~n31880 & ~n1014;
  assign n1016 = ~n1008 & n1015;
  assign n1017 = pi106  & ~n1016;
  assign n1018 = ~pi104  & ~pi105 ;
  assign n1019 = ~pi106  & n1018;
  assign n1020 = ~n1017 & ~n1019;
  assign n1021 = ~n855 & ~n1020;
  assign n1022 = ~n701 & ~n31862;
  assign n1023 = ~n702 & n1022;
  assign n1024 = ~n718 & n1023;
  assign n1025 = ~n31844 & n1024;
  assign n1026 = n31842 & n720;
  assign n1027 = ~n712 & n1025;
  assign n1028 = ~n1019 & ~n31881;
  assign n1029 = ~n853 & n1028;
  assign n1030 = ~n31860 & n1029;
  assign n1031 = ~n847 & n1030;
  assign n1032 = n855 & n1020;
  assign n1033 = ~n1017 & n1031;
  assign n1034 = ~pi106  & ~n1016;
  assign n1035 = pi107  & ~n1034;
  assign n1036 = ~pi107  & n1034;
  assign n1037 = n857 & ~n1016;
  assign n1038 = ~n1035 & ~n31883;
  assign n1039 = ~n31882 & n1038;
  assign n1040 = ~n1021 & ~n1039;
  assign n1041 = ~n720 & ~n1040;
  assign n1042 = ~n855 & ~n1014;
  assign n1043 = ~n31880 & n1042;
  assign n1044 = ~n1008 & n1043;
  assign n1045 = ~n31883 & ~n1044;
  assign n1046 = pi108  & ~n1045;
  assign n1047 = ~pi108  & ~n1044;
  assign n1048 = ~pi108  & n1045;
  assign n1049 = ~n31883 & n1047;
  assign n1050 = ~n1046 & ~n31884;
  assign n1051 = n720 & ~n1021;
  assign n1052 = n720 & n1040;
  assign n1053 = ~n1039 & n1051;
  assign n1054 = ~n1050 & ~n31885;
  assign n1055 = ~n1041 & ~n1054;
  assign n1056 = ~n592 & ~n1055;
  assign n1057 = n592 & ~n1041;
  assign n1058 = ~n1054 & n1057;
  assign n1059 = ~n860 & ~n31863;
  assign n1060 = ~n1016 & n1059;
  assign n1061 = n865 & ~n1060;
  assign n1062 = ~n865 & n1059;
  assign n1063 = ~n865 & n1060;
  assign n1064 = ~n1016 & n1062;
  assign n1065 = ~n1061 & ~n31886;
  assign n1066 = ~n1058 & ~n1065;
  assign n1067 = ~n1056 & ~n1066;
  assign n1068 = ~n487 & ~n1067;
  assign n1069 = ~n880 & ~n882;
  assign n1070 = ~n1016 & n1069;
  assign n1071 = ~n891 & ~n1070;
  assign n1072 = ~n882 & n891;
  assign n1073 = ~n880 & n1072;
  assign n1074 = n891 & n1070;
  assign n1075 = ~n1016 & n1073;
  assign n1076 = ~n1071 & ~n31887;
  assign n1077 = n487 & ~n1056;
  assign n1078 = n487 & n1067;
  assign n1079 = ~n1066 & n1077;
  assign n1080 = ~n1076 & ~n31888;
  assign n1081 = ~n1068 & ~n1080;
  assign n1082 = ~n393 & ~n1081;
  assign n1083 = n393 & ~n1068;
  assign n1084 = ~n1080 & n1083;
  assign n1085 = ~n894 & ~n31865;
  assign n1086 = ~n1016 & n1085;
  assign n1087 = ~n904 & ~n1086;
  assign n1088 = ~n894 & n904;
  assign n1089 = ~n31865 & n1088;
  assign n1090 = n904 & n1086;
  assign n1091 = ~n1016 & n1089;
  assign n1092 = n904 & ~n1086;
  assign n1093 = ~n904 & n1086;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = ~n1087 & ~n31889;
  assign n1096 = ~n1084 & n31890;
  assign n1097 = ~n1082 & ~n1096;
  assign n1098 = ~n321 & ~n1097;
  assign n1099 = ~n907 & ~n909;
  assign n1100 = ~n1016 & n1099;
  assign n1101 = ~n31868 & ~n1100;
  assign n1102 = ~n909 & n31868;
  assign n1103 = ~n907 & n1102;
  assign n1104 = n31868 & n1100;
  assign n1105 = ~n1016 & n1103;
  assign n1106 = ~n1101 & ~n31891;
  assign n1107 = n321 & ~n1082;
  assign n1108 = n321 & n1097;
  assign n1109 = ~n1096 & n1107;
  assign n1110 = ~n1106 & ~n31892;
  assign n1111 = ~n1098 & ~n1110;
  assign n1112 = ~n263 & ~n1111;
  assign n1113 = n263 & ~n1098;
  assign n1114 = ~n1110 & n1113;
  assign n1115 = ~n924 & ~n31869;
  assign n1116 = ~n1016 & n1115;
  assign n1117 = ~n31871 & ~n1116;
  assign n1118 = n31871 & n1116;
  assign n1119 = ~n924 & ~n31871;
  assign n1120 = ~n31869 & n1119;
  assign n1121 = ~n1016 & n1120;
  assign n1122 = n31871 & ~n1116;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = ~n1117 & ~n1118;
  assign n1125 = ~n1114 & ~n31893;
  assign n1126 = ~n1112 & ~n1125;
  assign n1127 = ~n214 & ~n1126;
  assign n1128 = ~n941 & ~n943;
  assign n1129 = ~n1016 & n1128;
  assign n1130 = ~n31873 & ~n1129;
  assign n1131 = ~n943 & n31873;
  assign n1132 = ~n941 & n1131;
  assign n1133 = n31873 & n1129;
  assign n1134 = ~n1016 & n1132;
  assign n1135 = ~n1130 & ~n31894;
  assign n1136 = n214 & ~n1112;
  assign n1137 = n214 & n1126;
  assign n1138 = ~n1125 & n1136;
  assign n1139 = ~n1135 & ~n31895;
  assign n1140 = ~n1127 & ~n1139;
  assign n1141 = ~n197 & ~n1140;
  assign n1142 = n197 & ~n1127;
  assign n1143 = ~n1139 & n1142;
  assign n1144 = ~n958 & ~n31874;
  assign n1145 = ~n1016 & n1144;
  assign n1146 = ~n31875 & n1145;
  assign n1147 = n31875 & ~n1145;
  assign n1148 = ~n958 & n31875;
  assign n1149 = ~n31874 & n1148;
  assign n1150 = ~n1016 & n1149;
  assign n1151 = ~n31875 & ~n1145;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = ~n1146 & ~n1147;
  assign n1154 = ~n1143 & ~n31896;
  assign n1155 = ~n1141 & ~n1154;
  assign n1156 = ~n974 & ~n976;
  assign n1157 = ~n1016 & n1156;
  assign n1158 = ~n31877 & ~n1157;
  assign n1159 = ~n976 & n31877;
  assign n1160 = ~n974 & n1159;
  assign n1161 = n31877 & n1157;
  assign n1162 = ~n1016 & n1160;
  assign n1163 = ~n1158 & ~n31897;
  assign n1164 = ~n990 & ~n31878;
  assign n1165 = ~n31878 & ~n1016;
  assign n1166 = ~n990 & n1165;
  assign n1167 = ~n1016 & n1164;
  assign n1168 = ~n31880 & ~n31898;
  assign n1169 = ~n1163 & n1168;
  assign n1170 = ~n1155 & n1169;
  assign n1171 = n193 & ~n1170;
  assign n1172 = ~n1141 & n1163;
  assign n1173 = n1155 & n1163;
  assign n1174 = ~n1154 & n1172;
  assign n1175 = n990 & ~n1165;
  assign n1176 = ~n193 & ~n1164;
  assign n1177 = ~n1175 & n1176;
  assign n1178 = ~n31899 & ~n1177;
  assign n1179 = ~n1171 & n1178;
  assign n1180 = pi104  & ~n1179;
  assign n1181 = ~pi102  & ~pi103 ;
  assign n1182 = ~pi104  & n1181;
  assign n1183 = ~n1180 & ~n1182;
  assign n1184 = ~n1016 & ~n1183;
  assign n1185 = ~pi104  & ~n1179;
  assign n1186 = pi105  & ~n1185;
  assign n1187 = ~pi105  & n1185;
  assign n1188 = n1018 & ~n1179;
  assign n1189 = ~n1186 & ~n31900;
  assign n1190 = ~n31858 & ~n31881;
  assign n1191 = ~n834 & n1190;
  assign n1192 = ~n853 & n1191;
  assign n1193 = ~n31860 & n1192;
  assign n1194 = n839 & n855;
  assign n1195 = ~n847 & n1193;
  assign n1196 = ~n1182 & ~n31901;
  assign n1197 = ~n1014 & n1196;
  assign n1198 = ~n31880 & n1197;
  assign n1199 = ~n1008 & n1198;
  assign n1200 = n1016 & n1183;
  assign n1201 = ~n1180 & n1199;
  assign n1202 = n1189 & ~n31902;
  assign n1203 = ~n1184 & ~n1202;
  assign n1204 = ~n855 & ~n1203;
  assign n1205 = n855 & ~n1184;
  assign n1206 = ~n1202 & n1205;
  assign n1207 = ~n1016 & ~n1177;
  assign n1208 = ~n31899 & n1207;
  assign n1209 = ~n1171 & n1208;
  assign n1210 = ~n31900 & ~n1209;
  assign n1211 = pi106  & ~n1210;
  assign n1212 = ~pi106  & ~n1209;
  assign n1213 = ~pi106  & n1210;
  assign n1214 = ~n31900 & n1212;
  assign n1215 = ~n1211 & ~n31903;
  assign n1216 = ~n1206 & ~n1215;
  assign n1217 = ~n1204 & ~n1216;
  assign n1218 = ~n720 & ~n1217;
  assign n1219 = n720 & ~n1204;
  assign n1220 = ~n1216 & n1219;
  assign n1221 = n720 & n1217;
  assign n1222 = ~n1021 & ~n31882;
  assign n1223 = ~n1179 & n1222;
  assign n1224 = n1038 & ~n1223;
  assign n1225 = ~n1038 & n1222;
  assign n1226 = ~n1038 & n1223;
  assign n1227 = ~n1179 & n1225;
  assign n1228 = ~n1224 & ~n31905;
  assign n1229 = ~n31904 & ~n1228;
  assign n1230 = ~n1218 & ~n1229;
  assign n1231 = ~n592 & ~n1230;
  assign n1232 = n592 & ~n1218;
  assign n1233 = ~n1229 & n1232;
  assign n1234 = ~n1041 & ~n31885;
  assign n1235 = ~n1041 & ~n1179;
  assign n1236 = ~n31885 & n1235;
  assign n1237 = ~n1179 & n1234;
  assign n1238 = n1050 & ~n31906;
  assign n1239 = n1054 & n1235;
  assign n1240 = n1050 & ~n31885;
  assign n1241 = ~n1041 & n1240;
  assign n1242 = ~n1179 & n1241;
  assign n1243 = ~n1050 & ~n31906;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = ~n1238 & ~n1239;
  assign n1246 = ~n1233 & ~n31907;
  assign n1247 = ~n1231 & ~n1246;
  assign n1248 = ~n487 & ~n1247;
  assign n1249 = n487 & ~n1231;
  assign n1250 = ~n1246 & n1249;
  assign n1251 = n487 & n1247;
  assign n1252 = ~n1056 & ~n1058;
  assign n1253 = ~n1179 & n1252;
  assign n1254 = ~n1065 & ~n1253;
  assign n1255 = ~n1056 & n1065;
  assign n1256 = ~n1058 & n1255;
  assign n1257 = n1065 & n1253;
  assign n1258 = ~n1179 & n1256;
  assign n1259 = n1065 & ~n1253;
  assign n1260 = ~n1065 & n1253;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = ~n1254 & ~n31909;
  assign n1263 = ~n31908 & n31910;
  assign n1264 = ~n1248 & ~n1263;
  assign n1265 = ~n393 & ~n1264;
  assign n1266 = n393 & ~n1248;
  assign n1267 = ~n1263 & n1266;
  assign n1268 = ~n1068 & ~n31888;
  assign n1269 = ~n1068 & ~n1179;
  assign n1270 = ~n31888 & n1269;
  assign n1271 = ~n1179 & n1268;
  assign n1272 = n1076 & ~n31911;
  assign n1273 = n1080 & n1269;
  assign n1274 = n1076 & ~n31888;
  assign n1275 = ~n1068 & n1274;
  assign n1276 = ~n1179 & n1275;
  assign n1277 = ~n1076 & ~n31911;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = ~n1272 & ~n1273;
  assign n1280 = ~n1267 & ~n31912;
  assign n1281 = ~n1265 & ~n1280;
  assign n1282 = ~n321 & ~n1281;
  assign n1283 = n321 & ~n1265;
  assign n1284 = ~n1280 & n1283;
  assign n1285 = n321 & n1281;
  assign n1286 = ~n1082 & ~n1084;
  assign n1287 = ~n1179 & n1286;
  assign n1288 = ~n31890 & ~n1287;
  assign n1289 = n31890 & n1287;
  assign n1290 = ~n1082 & ~n31890;
  assign n1291 = ~n1084 & n1290;
  assign n1292 = ~n1179 & n1291;
  assign n1293 = n31890 & ~n1287;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = ~n1288 & ~n1289;
  assign n1296 = ~n31913 & ~n31914;
  assign n1297 = ~n1282 & ~n1296;
  assign n1298 = ~n263 & ~n1297;
  assign n1299 = n263 & ~n1282;
  assign n1300 = ~n1296 & n1299;
  assign n1301 = ~n1098 & ~n31892;
  assign n1302 = ~n1098 & ~n1179;
  assign n1303 = ~n31892 & n1302;
  assign n1304 = ~n1179 & n1301;
  assign n1305 = n1106 & ~n31915;
  assign n1306 = n1110 & n1302;
  assign n1307 = n1106 & ~n31892;
  assign n1308 = ~n1098 & n1307;
  assign n1309 = ~n1179 & n1308;
  assign n1310 = ~n1106 & ~n31915;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = ~n1305 & ~n1306;
  assign n1313 = ~n1300 & ~n31916;
  assign n1314 = ~n1298 & ~n1313;
  assign n1315 = ~n214 & ~n1314;
  assign n1316 = n214 & ~n1298;
  assign n1317 = ~n1313 & n1316;
  assign n1318 = n214 & n1314;
  assign n1319 = ~n1112 & ~n1114;
  assign n1320 = ~n1179 & n1319;
  assign n1321 = ~n31893 & n1320;
  assign n1322 = n31893 & ~n1320;
  assign n1323 = ~n1112 & n31893;
  assign n1324 = ~n1114 & n1323;
  assign n1325 = ~n1179 & n1324;
  assign n1326 = ~n31893 & ~n1320;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = ~n1321 & ~n1322;
  assign n1329 = ~n31917 & ~n31918;
  assign n1330 = ~n1315 & ~n1329;
  assign n1331 = ~n197 & ~n1330;
  assign n1332 = n197 & ~n1315;
  assign n1333 = ~n1329 & n1332;
  assign n1334 = ~n1127 & ~n31895;
  assign n1335 = ~n1127 & ~n1179;
  assign n1336 = ~n31895 & n1335;
  assign n1337 = ~n1179 & n1334;
  assign n1338 = n1135 & ~n31919;
  assign n1339 = n1139 & n1335;
  assign n1340 = n1135 & ~n31895;
  assign n1341 = ~n1127 & n1340;
  assign n1342 = ~n1179 & n1341;
  assign n1343 = ~n1135 & ~n31919;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = ~n1338 & ~n1339;
  assign n1346 = ~n1333 & ~n31920;
  assign n1347 = ~n1331 & ~n1346;
  assign n1348 = ~n1141 & ~n1143;
  assign n1349 = ~n1179 & n1348;
  assign n1350 = ~n31896 & n1349;
  assign n1351 = n31896 & ~n1349;
  assign n1352 = ~n31896 & ~n1349;
  assign n1353 = ~n1141 & n31896;
  assign n1354 = ~n1143 & n1353;
  assign n1355 = n31896 & n1349;
  assign n1356 = ~n1179 & n1354;
  assign n1357 = ~n1352 & ~n31921;
  assign n1358 = ~n1350 & ~n1351;
  assign n1359 = ~n1155 & ~n1163;
  assign n1360 = ~n1163 & ~n1179;
  assign n1361 = ~n1155 & n1360;
  assign n1362 = ~n1179 & n1359;
  assign n1363 = ~n31899 & ~n31923;
  assign n1364 = ~n31922 & n1363;
  assign n1365 = ~n1347 & n1364;
  assign n1366 = n193 & ~n1365;
  assign n1367 = ~n1331 & n31922;
  assign n1368 = ~n1346 & n1367;
  assign n1369 = n1347 & n31922;
  assign n1370 = n1155 & ~n1360;
  assign n1371 = ~n193 & ~n1359;
  assign n1372 = ~n1370 & n1371;
  assign n1373 = ~n31924 & ~n1372;
  assign n1374 = ~n1366 & n1373;
  assign n1375 = pi102  & ~n1374;
  assign n1376 = ~pi100  & ~pi101 ;
  assign n1377 = ~pi102  & n1376;
  assign n1378 = ~n1375 & ~n1377;
  assign n1379 = ~n1179 & ~n1378;
  assign n1380 = ~n997 & ~n31901;
  assign n1381 = ~n998 & n1380;
  assign n1382 = ~n1014 & n1381;
  assign n1383 = ~n31880 & n1382;
  assign n1384 = n31878 & n1016;
  assign n1385 = ~n1008 & n1383;
  assign n1386 = ~n1377 & ~n31925;
  assign n1387 = ~n1177 & n1386;
  assign n1388 = ~n31899 & n1387;
  assign n1389 = ~n1171 & n1388;
  assign n1390 = n1179 & n1378;
  assign n1391 = ~n1375 & n1389;
  assign n1392 = ~pi102  & ~n1374;
  assign n1393 = pi103  & ~n1392;
  assign n1394 = ~pi103  & n1392;
  assign n1395 = n1181 & ~n1374;
  assign n1396 = ~n1393 & ~n31927;
  assign n1397 = ~n31926 & n1396;
  assign n1398 = ~n1379 & ~n1397;
  assign n1399 = ~n1016 & ~n1398;
  assign n1400 = ~n1179 & ~n1372;
  assign n1401 = ~n31924 & n1400;
  assign n1402 = ~n1366 & n1401;
  assign n1403 = ~n31927 & ~n1402;
  assign n1404 = pi104  & ~n1403;
  assign n1405 = ~pi104  & ~n1402;
  assign n1406 = ~pi104  & n1403;
  assign n1407 = ~n31927 & n1405;
  assign n1408 = ~n1404 & ~n31928;
  assign n1409 = n1016 & ~n1379;
  assign n1410 = n1016 & n1398;
  assign n1411 = ~n1397 & n1409;
  assign n1412 = ~n1408 & ~n31929;
  assign n1413 = ~n1399 & ~n1412;
  assign n1414 = ~n855 & ~n1413;
  assign n1415 = n855 & ~n1399;
  assign n1416 = ~n1412 & n1415;
  assign n1417 = ~n1184 & ~n31902;
  assign n1418 = ~n1374 & n1417;
  assign n1419 = n1189 & ~n1418;
  assign n1420 = ~n1189 & n1417;
  assign n1421 = ~n1189 & n1418;
  assign n1422 = ~n1374 & n1420;
  assign n1423 = ~n1419 & ~n31930;
  assign n1424 = ~n1416 & ~n1423;
  assign n1425 = ~n1414 & ~n1424;
  assign n1426 = ~n720 & ~n1425;
  assign n1427 = ~n1204 & ~n1206;
  assign n1428 = ~n1374 & n1427;
  assign n1429 = ~n1215 & ~n1428;
  assign n1430 = ~n1206 & n1215;
  assign n1431 = ~n1204 & n1430;
  assign n1432 = n1215 & n1428;
  assign n1433 = ~n1374 & n1431;
  assign n1434 = ~n1429 & ~n31931;
  assign n1435 = n720 & ~n1414;
  assign n1436 = n720 & n1425;
  assign n1437 = ~n1424 & n1435;
  assign n1438 = ~n1434 & ~n31932;
  assign n1439 = ~n1426 & ~n1438;
  assign n1440 = ~n592 & ~n1439;
  assign n1441 = n592 & ~n1426;
  assign n1442 = ~n1438 & n1441;
  assign n1443 = ~n1218 & ~n31904;
  assign n1444 = ~n1374 & n1443;
  assign n1445 = ~n1228 & ~n1444;
  assign n1446 = ~n1218 & n1228;
  assign n1447 = ~n31904 & n1446;
  assign n1448 = n1228 & n1444;
  assign n1449 = ~n1374 & n1447;
  assign n1450 = n1228 & ~n1444;
  assign n1451 = ~n1228 & n1444;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = ~n1445 & ~n31933;
  assign n1454 = ~n1442 & n31934;
  assign n1455 = ~n1440 & ~n1454;
  assign n1456 = ~n487 & ~n1455;
  assign n1457 = ~n1231 & ~n1233;
  assign n1458 = ~n1374 & n1457;
  assign n1459 = ~n31907 & ~n1458;
  assign n1460 = ~n1233 & n31907;
  assign n1461 = ~n1231 & n1460;
  assign n1462 = n31907 & n1458;
  assign n1463 = ~n1374 & n1461;
  assign n1464 = ~n1459 & ~n31935;
  assign n1465 = n487 & ~n1440;
  assign n1466 = n487 & n1455;
  assign n1467 = ~n1454 & n1465;
  assign n1468 = ~n1464 & ~n31936;
  assign n1469 = ~n1456 & ~n1468;
  assign n1470 = ~n393 & ~n1469;
  assign n1471 = n393 & ~n1456;
  assign n1472 = ~n1468 & n1471;
  assign n1473 = ~n1248 & ~n31908;
  assign n1474 = ~n1374 & n1473;
  assign n1475 = ~n31910 & ~n1474;
  assign n1476 = n31910 & n1474;
  assign n1477 = ~n1248 & ~n31910;
  assign n1478 = ~n31908 & n1477;
  assign n1479 = ~n1374 & n1478;
  assign n1480 = n31910 & ~n1474;
  assign n1481 = ~n1479 & ~n1480;
  assign n1482 = ~n1475 & ~n1476;
  assign n1483 = ~n1472 & ~n31937;
  assign n1484 = ~n1470 & ~n1483;
  assign n1485 = ~n321 & ~n1484;
  assign n1486 = ~n1265 & ~n1267;
  assign n1487 = ~n1374 & n1486;
  assign n1488 = ~n31912 & ~n1487;
  assign n1489 = ~n1267 & n31912;
  assign n1490 = ~n1265 & n1489;
  assign n1491 = n31912 & n1487;
  assign n1492 = ~n1374 & n1490;
  assign n1493 = ~n1488 & ~n31938;
  assign n1494 = n321 & ~n1470;
  assign n1495 = n321 & n1484;
  assign n1496 = ~n1483 & n1494;
  assign n1497 = ~n1493 & ~n31939;
  assign n1498 = ~n1485 & ~n1497;
  assign n1499 = ~n263 & ~n1498;
  assign n1500 = n263 & ~n1485;
  assign n1501 = ~n1497 & n1500;
  assign n1502 = ~n1282 & ~n31913;
  assign n1503 = ~n1374 & n1502;
  assign n1504 = ~n31914 & n1503;
  assign n1505 = n31914 & ~n1503;
  assign n1506 = ~n1282 & n31914;
  assign n1507 = ~n31913 & n1506;
  assign n1508 = ~n1374 & n1507;
  assign n1509 = ~n31914 & ~n1503;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = ~n1504 & ~n1505;
  assign n1512 = ~n1501 & ~n31940;
  assign n1513 = ~n1499 & ~n1512;
  assign n1514 = ~n214 & ~n1513;
  assign n1515 = ~n1298 & ~n1300;
  assign n1516 = ~n1374 & n1515;
  assign n1517 = ~n31916 & ~n1516;
  assign n1518 = ~n1300 & n31916;
  assign n1519 = ~n1298 & n1518;
  assign n1520 = n31916 & n1516;
  assign n1521 = ~n1374 & n1519;
  assign n1522 = ~n1517 & ~n31941;
  assign n1523 = n214 & ~n1499;
  assign n1524 = n214 & n1513;
  assign n1525 = ~n1512 & n1523;
  assign n1526 = ~n1522 & ~n31942;
  assign n1527 = ~n1514 & ~n1526;
  assign n1528 = ~n197 & ~n1527;
  assign n1529 = n197 & ~n1514;
  assign n1530 = ~n1526 & n1529;
  assign n1531 = ~n1315 & ~n31917;
  assign n1532 = ~n1374 & n1531;
  assign n1533 = ~n31918 & ~n1532;
  assign n1534 = ~n1315 & n31918;
  assign n1535 = ~n31917 & n1534;
  assign n1536 = n31918 & n1532;
  assign n1537 = ~n1374 & n1535;
  assign n1538 = n31918 & ~n1532;
  assign n1539 = ~n31918 & n1532;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = ~n1533 & ~n31943;
  assign n1542 = ~n1530 & n31944;
  assign n1543 = ~n1528 & ~n1542;
  assign n1544 = ~n1331 & ~n1333;
  assign n1545 = ~n1374 & n1544;
  assign n1546 = ~n31920 & ~n1545;
  assign n1547 = ~n1333 & n31920;
  assign n1548 = ~n1331 & n1547;
  assign n1549 = n31920 & n1545;
  assign n1550 = ~n1374 & n1548;
  assign n1551 = ~n1546 & ~n31945;
  assign n1552 = ~n1347 & ~n31922;
  assign n1553 = ~n31922 & ~n1374;
  assign n1554 = ~n1347 & n1553;
  assign n1555 = ~n1374 & n1552;
  assign n1556 = ~n31924 & ~n31946;
  assign n1557 = ~n1551 & n1556;
  assign n1558 = ~n1543 & n1557;
  assign n1559 = n193 & ~n1558;
  assign n1560 = ~n1528 & n1551;
  assign n1561 = n1543 & n1551;
  assign n1562 = ~n1542 & n1560;
  assign n1563 = n1347 & ~n1553;
  assign n1564 = ~n193 & ~n1552;
  assign n1565 = ~n1563 & n1564;
  assign n1566 = ~n31947 & ~n1565;
  assign n1567 = ~n1559 & n1566;
  assign n1568 = pi100  & ~n1567;
  assign n1569 = ~pi98  & ~pi99 ;
  assign n1570 = ~pi100  & n1569;
  assign n1571 = ~n1568 & ~n1570;
  assign n1572 = ~n1374 & ~n1571;
  assign n1573 = ~pi100  & ~n1567;
  assign n1574 = pi101  & ~n1573;
  assign n1575 = ~pi101  & n1573;
  assign n1576 = n1376 & ~n1567;
  assign n1577 = ~n1574 & ~n31948;
  assign n1578 = ~n31897 & ~n31925;
  assign n1579 = ~n1158 & n1578;
  assign n1580 = ~n1177 & n1579;
  assign n1581 = ~n31899 & n1580;
  assign n1582 = n1163 & n1179;
  assign n1583 = ~n1171 & n1581;
  assign n1584 = ~n1570 & ~n31949;
  assign n1585 = ~n1372 & n1584;
  assign n1586 = ~n31924 & n1585;
  assign n1587 = ~n1366 & n1586;
  assign n1588 = n1374 & n1571;
  assign n1589 = ~n1568 & n1587;
  assign n1590 = n1577 & ~n31950;
  assign n1591 = ~n1572 & ~n1590;
  assign n1592 = ~n1179 & ~n1591;
  assign n1593 = n1179 & ~n1572;
  assign n1594 = ~n1590 & n1593;
  assign n1595 = ~n1374 & ~n1565;
  assign n1596 = ~n31947 & n1595;
  assign n1597 = ~n1559 & n1596;
  assign n1598 = ~n31948 & ~n1597;
  assign n1599 = pi102  & ~n1598;
  assign n1600 = ~pi102  & ~n1597;
  assign n1601 = ~pi102  & n1598;
  assign n1602 = ~n31948 & n1600;
  assign n1603 = ~n1599 & ~n31951;
  assign n1604 = ~n1594 & ~n1603;
  assign n1605 = ~n1592 & ~n1604;
  assign n1606 = ~n1016 & ~n1605;
  assign n1607 = n1016 & ~n1592;
  assign n1608 = ~n1604 & n1607;
  assign n1609 = n1016 & n1605;
  assign n1610 = ~n1379 & ~n31926;
  assign n1611 = ~n1567 & n1610;
  assign n1612 = n1396 & ~n1611;
  assign n1613 = ~n1396 & n1610;
  assign n1614 = ~n1396 & n1611;
  assign n1615 = ~n1567 & n1613;
  assign n1616 = ~n1612 & ~n31953;
  assign n1617 = ~n31952 & ~n1616;
  assign n1618 = ~n1606 & ~n1617;
  assign n1619 = ~n855 & ~n1618;
  assign n1620 = n855 & ~n1606;
  assign n1621 = ~n1617 & n1620;
  assign n1622 = ~n1399 & ~n31929;
  assign n1623 = ~n1399 & ~n1567;
  assign n1624 = ~n31929 & n1623;
  assign n1625 = ~n1567 & n1622;
  assign n1626 = n1408 & ~n31954;
  assign n1627 = n1412 & n1623;
  assign n1628 = n1408 & ~n31929;
  assign n1629 = ~n1399 & n1628;
  assign n1630 = ~n1567 & n1629;
  assign n1631 = ~n1408 & ~n31954;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = ~n1626 & ~n1627;
  assign n1634 = ~n1621 & ~n31955;
  assign n1635 = ~n1619 & ~n1634;
  assign n1636 = ~n720 & ~n1635;
  assign n1637 = n720 & ~n1619;
  assign n1638 = ~n1634 & n1637;
  assign n1639 = n720 & n1635;
  assign n1640 = ~n1414 & ~n1416;
  assign n1641 = ~n1567 & n1640;
  assign n1642 = ~n1423 & ~n1641;
  assign n1643 = ~n1414 & n1423;
  assign n1644 = ~n1416 & n1643;
  assign n1645 = n1423 & n1641;
  assign n1646 = ~n1567 & n1644;
  assign n1647 = n1423 & ~n1641;
  assign n1648 = ~n1423 & n1641;
  assign n1649 = ~n1647 & ~n1648;
  assign n1650 = ~n1642 & ~n31957;
  assign n1651 = ~n31956 & n31958;
  assign n1652 = ~n1636 & ~n1651;
  assign n1653 = ~n592 & ~n1652;
  assign n1654 = n592 & ~n1636;
  assign n1655 = ~n1651 & n1654;
  assign n1656 = ~n1426 & ~n31932;
  assign n1657 = ~n1426 & ~n1567;
  assign n1658 = ~n31932 & n1657;
  assign n1659 = ~n1567 & n1656;
  assign n1660 = n1434 & ~n31959;
  assign n1661 = n1438 & n1657;
  assign n1662 = n1434 & ~n31932;
  assign n1663 = ~n1426 & n1662;
  assign n1664 = ~n1567 & n1663;
  assign n1665 = ~n1434 & ~n31959;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = ~n1660 & ~n1661;
  assign n1668 = ~n1655 & ~n31960;
  assign n1669 = ~n1653 & ~n1668;
  assign n1670 = ~n487 & ~n1669;
  assign n1671 = n487 & ~n1653;
  assign n1672 = ~n1668 & n1671;
  assign n1673 = n487 & n1669;
  assign n1674 = ~n1440 & ~n1442;
  assign n1675 = ~n1567 & n1674;
  assign n1676 = ~n31934 & ~n1675;
  assign n1677 = n31934 & n1675;
  assign n1678 = ~n1440 & ~n31934;
  assign n1679 = ~n1442 & n1678;
  assign n1680 = ~n1567 & n1679;
  assign n1681 = n31934 & ~n1675;
  assign n1682 = ~n1680 & ~n1681;
  assign n1683 = ~n1676 & ~n1677;
  assign n1684 = ~n31961 & ~n31962;
  assign n1685 = ~n1670 & ~n1684;
  assign n1686 = ~n393 & ~n1685;
  assign n1687 = n393 & ~n1670;
  assign n1688 = ~n1684 & n1687;
  assign n1689 = ~n1456 & ~n31936;
  assign n1690 = ~n1456 & ~n1567;
  assign n1691 = ~n31936 & n1690;
  assign n1692 = ~n1567 & n1689;
  assign n1693 = n1464 & ~n31963;
  assign n1694 = n1468 & n1690;
  assign n1695 = n1464 & ~n31936;
  assign n1696 = ~n1456 & n1695;
  assign n1697 = ~n1567 & n1696;
  assign n1698 = ~n1464 & ~n31963;
  assign n1699 = ~n1697 & ~n1698;
  assign n1700 = ~n1693 & ~n1694;
  assign n1701 = ~n1688 & ~n31964;
  assign n1702 = ~n1686 & ~n1701;
  assign n1703 = ~n321 & ~n1702;
  assign n1704 = n321 & ~n1686;
  assign n1705 = ~n1701 & n1704;
  assign n1706 = n321 & n1702;
  assign n1707 = ~n1470 & ~n1472;
  assign n1708 = ~n1567 & n1707;
  assign n1709 = ~n31937 & n1708;
  assign n1710 = n31937 & ~n1708;
  assign n1711 = ~n1470 & n31937;
  assign n1712 = ~n1472 & n1711;
  assign n1713 = ~n1567 & n1712;
  assign n1714 = ~n31937 & ~n1708;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = ~n1709 & ~n1710;
  assign n1717 = ~n31965 & ~n31966;
  assign n1718 = ~n1703 & ~n1717;
  assign n1719 = ~n263 & ~n1718;
  assign n1720 = n263 & ~n1703;
  assign n1721 = ~n1717 & n1720;
  assign n1722 = ~n1485 & ~n31939;
  assign n1723 = ~n1485 & ~n1567;
  assign n1724 = ~n31939 & n1723;
  assign n1725 = ~n1567 & n1722;
  assign n1726 = n1493 & ~n31967;
  assign n1727 = n1497 & n1723;
  assign n1728 = n1493 & ~n31939;
  assign n1729 = ~n1485 & n1728;
  assign n1730 = ~n1567 & n1729;
  assign n1731 = ~n1493 & ~n31967;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = ~n1726 & ~n1727;
  assign n1734 = ~n1721 & ~n31968;
  assign n1735 = ~n1719 & ~n1734;
  assign n1736 = ~n214 & ~n1735;
  assign n1737 = n214 & ~n1719;
  assign n1738 = ~n1734 & n1737;
  assign n1739 = n214 & n1735;
  assign n1740 = ~n1499 & ~n1501;
  assign n1741 = ~n1567 & n1740;
  assign n1742 = ~n31940 & n1741;
  assign n1743 = n31940 & ~n1741;
  assign n1744 = ~n31940 & ~n1741;
  assign n1745 = ~n1499 & n31940;
  assign n1746 = ~n1501 & n1745;
  assign n1747 = n31940 & n1741;
  assign n1748 = ~n1567 & n1746;
  assign n1749 = ~n1744 & ~n31970;
  assign n1750 = ~n1742 & ~n1743;
  assign n1751 = ~n31969 & ~n31971;
  assign n1752 = ~n1736 & ~n1751;
  assign n1753 = ~n197 & ~n1752;
  assign n1754 = n197 & ~n1736;
  assign n1755 = ~n1751 & n1754;
  assign n1756 = ~n1514 & ~n31942;
  assign n1757 = ~n1514 & ~n1567;
  assign n1758 = ~n31942 & n1757;
  assign n1759 = ~n1567 & n1756;
  assign n1760 = n1522 & ~n31972;
  assign n1761 = n1526 & n1757;
  assign n1762 = n1522 & ~n31942;
  assign n1763 = ~n1514 & n1762;
  assign n1764 = ~n1567 & n1763;
  assign n1765 = ~n1522 & ~n31972;
  assign n1766 = ~n1764 & ~n1765;
  assign n1767 = ~n1760 & ~n1761;
  assign n1768 = ~n1755 & ~n31973;
  assign n1769 = ~n1753 & ~n1768;
  assign n1770 = ~n1528 & ~n1530;
  assign n1771 = ~n1567 & n1770;
  assign n1772 = ~n31944 & ~n1771;
  assign n1773 = n31944 & n1771;
  assign n1774 = n31944 & ~n1771;
  assign n1775 = ~n1528 & ~n31944;
  assign n1776 = ~n1530 & n1775;
  assign n1777 = ~n31944 & n1771;
  assign n1778 = ~n1567 & n1776;
  assign n1779 = ~n1774 & ~n31974;
  assign n1780 = ~n1772 & ~n1773;
  assign n1781 = ~n1543 & ~n1551;
  assign n1782 = ~n1551 & ~n1567;
  assign n1783 = ~n1543 & n1782;
  assign n1784 = ~n1567 & n1781;
  assign n1785 = ~n31947 & ~n31976;
  assign n1786 = ~n31975 & n1785;
  assign n1787 = ~n1769 & n1786;
  assign n1788 = n193 & ~n1787;
  assign n1789 = ~n1753 & n31975;
  assign n1790 = ~n1768 & n1789;
  assign n1791 = n1769 & n31975;
  assign n1792 = n1543 & ~n1782;
  assign n1793 = ~n193 & ~n1781;
  assign n1794 = ~n1792 & n1793;
  assign n1795 = ~n31977 & ~n1794;
  assign n1796 = ~n1788 & n1795;
  assign n1797 = pi98  & ~n1796;
  assign n1798 = ~pi96  & ~pi97 ;
  assign n1799 = ~pi98  & n1798;
  assign n1800 = ~n1797 & ~n1799;
  assign n1801 = ~n1567 & ~n1800;
  assign n1802 = ~n31921 & ~n31949;
  assign n1803 = ~n1352 & n1802;
  assign n1804 = ~n1372 & n1803;
  assign n1805 = ~n31924 & n1804;
  assign n1806 = n31922 & n1374;
  assign n1807 = ~n1366 & n1805;
  assign n1808 = ~n1799 & ~n31978;
  assign n1809 = ~n1565 & n1808;
  assign n1810 = ~n31947 & n1809;
  assign n1811 = ~n1559 & n1810;
  assign n1812 = n1567 & n1800;
  assign n1813 = ~n1797 & n1811;
  assign n1814 = ~pi98  & ~n1796;
  assign n1815 = pi99  & ~n1814;
  assign n1816 = ~pi99  & n1814;
  assign n1817 = n1569 & ~n1796;
  assign n1818 = ~n1815 & ~n31980;
  assign n1819 = ~n31979 & n1818;
  assign n1820 = ~n1801 & ~n1819;
  assign n1821 = ~n1374 & ~n1820;
  assign n1822 = ~n1567 & ~n1794;
  assign n1823 = ~n31977 & n1822;
  assign n1824 = ~n1788 & n1823;
  assign n1825 = ~n31980 & ~n1824;
  assign n1826 = pi100  & ~n1825;
  assign n1827 = ~pi100  & ~n1824;
  assign n1828 = ~pi100  & n1825;
  assign n1829 = ~n31980 & n1827;
  assign n1830 = ~n1826 & ~n31981;
  assign n1831 = n1374 & ~n1801;
  assign n1832 = n1374 & n1820;
  assign n1833 = ~n1819 & n1831;
  assign n1834 = ~n1830 & ~n31982;
  assign n1835 = ~n1821 & ~n1834;
  assign n1836 = ~n1179 & ~n1835;
  assign n1837 = n1179 & ~n1821;
  assign n1838 = ~n1834 & n1837;
  assign n1839 = ~n1572 & ~n31950;
  assign n1840 = ~n1796 & n1839;
  assign n1841 = n1577 & ~n1840;
  assign n1842 = ~n1577 & n1839;
  assign n1843 = ~n1577 & n1840;
  assign n1844 = ~n1796 & n1842;
  assign n1845 = ~n1841 & ~n31983;
  assign n1846 = ~n1838 & ~n1845;
  assign n1847 = ~n1836 & ~n1846;
  assign n1848 = ~n1016 & ~n1847;
  assign n1849 = ~n1592 & ~n1594;
  assign n1850 = ~n1796 & n1849;
  assign n1851 = ~n1603 & ~n1850;
  assign n1852 = ~n1594 & n1603;
  assign n1853 = ~n1592 & n1852;
  assign n1854 = n1603 & n1850;
  assign n1855 = ~n1796 & n1853;
  assign n1856 = ~n1851 & ~n31984;
  assign n1857 = n1016 & ~n1836;
  assign n1858 = n1016 & n1847;
  assign n1859 = ~n1846 & n1857;
  assign n1860 = ~n1856 & ~n31985;
  assign n1861 = ~n1848 & ~n1860;
  assign n1862 = ~n855 & ~n1861;
  assign n1863 = n855 & ~n1848;
  assign n1864 = ~n1860 & n1863;
  assign n1865 = ~n1606 & ~n31952;
  assign n1866 = ~n1796 & n1865;
  assign n1867 = ~n1616 & ~n1866;
  assign n1868 = ~n1606 & n1616;
  assign n1869 = ~n31952 & n1868;
  assign n1870 = n1616 & n1866;
  assign n1871 = ~n1796 & n1869;
  assign n1872 = n1616 & ~n1866;
  assign n1873 = ~n1616 & n1866;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = ~n1867 & ~n31986;
  assign n1876 = ~n1864 & n31987;
  assign n1877 = ~n1862 & ~n1876;
  assign n1878 = ~n720 & ~n1877;
  assign n1879 = ~n1619 & ~n1621;
  assign n1880 = ~n1796 & n1879;
  assign n1881 = ~n31955 & ~n1880;
  assign n1882 = ~n1621 & n31955;
  assign n1883 = ~n1619 & n1882;
  assign n1884 = n31955 & n1880;
  assign n1885 = ~n1796 & n1883;
  assign n1886 = ~n1881 & ~n31988;
  assign n1887 = n720 & ~n1862;
  assign n1888 = n720 & n1877;
  assign n1889 = ~n1876 & n1887;
  assign n1890 = ~n1886 & ~n31989;
  assign n1891 = ~n1878 & ~n1890;
  assign n1892 = ~n592 & ~n1891;
  assign n1893 = n592 & ~n1878;
  assign n1894 = ~n1890 & n1893;
  assign n1895 = ~n1636 & ~n31956;
  assign n1896 = ~n1796 & n1895;
  assign n1897 = ~n31958 & ~n1896;
  assign n1898 = n31958 & n1896;
  assign n1899 = ~n1636 & ~n31958;
  assign n1900 = ~n31956 & n1899;
  assign n1901 = ~n1796 & n1900;
  assign n1902 = n31958 & ~n1896;
  assign n1903 = ~n1901 & ~n1902;
  assign n1904 = ~n1897 & ~n1898;
  assign n1905 = ~n1894 & ~n31990;
  assign n1906 = ~n1892 & ~n1905;
  assign n1907 = ~n487 & ~n1906;
  assign n1908 = ~n1653 & ~n1655;
  assign n1909 = ~n1796 & n1908;
  assign n1910 = ~n31960 & ~n1909;
  assign n1911 = ~n1655 & n31960;
  assign n1912 = ~n1653 & n1911;
  assign n1913 = n31960 & n1909;
  assign n1914 = ~n1796 & n1912;
  assign n1915 = ~n1910 & ~n31991;
  assign n1916 = n487 & ~n1892;
  assign n1917 = n487 & n1906;
  assign n1918 = ~n1905 & n1916;
  assign n1919 = ~n1915 & ~n31992;
  assign n1920 = ~n1907 & ~n1919;
  assign n1921 = ~n393 & ~n1920;
  assign n1922 = n393 & ~n1907;
  assign n1923 = ~n1919 & n1922;
  assign n1924 = ~n1670 & ~n31961;
  assign n1925 = ~n1796 & n1924;
  assign n1926 = ~n31962 & n1925;
  assign n1927 = n31962 & ~n1925;
  assign n1928 = ~n1670 & n31962;
  assign n1929 = ~n31961 & n1928;
  assign n1930 = ~n1796 & n1929;
  assign n1931 = ~n31962 & ~n1925;
  assign n1932 = ~n1930 & ~n1931;
  assign n1933 = ~n1926 & ~n1927;
  assign n1934 = ~n1923 & ~n31993;
  assign n1935 = ~n1921 & ~n1934;
  assign n1936 = ~n321 & ~n1935;
  assign n1937 = ~n1686 & ~n1688;
  assign n1938 = ~n1796 & n1937;
  assign n1939 = ~n31964 & ~n1938;
  assign n1940 = ~n1688 & n31964;
  assign n1941 = ~n1686 & n1940;
  assign n1942 = n31964 & n1938;
  assign n1943 = ~n1796 & n1941;
  assign n1944 = ~n1939 & ~n31994;
  assign n1945 = n321 & ~n1921;
  assign n1946 = n321 & n1935;
  assign n1947 = ~n1934 & n1945;
  assign n1948 = ~n1944 & ~n31995;
  assign n1949 = ~n1936 & ~n1948;
  assign n1950 = ~n263 & ~n1949;
  assign n1951 = n263 & ~n1936;
  assign n1952 = ~n1948 & n1951;
  assign n1953 = ~n1703 & ~n31965;
  assign n1954 = ~n1796 & n1953;
  assign n1955 = ~n31966 & n1954;
  assign n1956 = n31966 & ~n1954;
  assign n1957 = ~n31966 & ~n1954;
  assign n1958 = ~n1703 & n31966;
  assign n1959 = ~n31965 & n1958;
  assign n1960 = n31966 & n1954;
  assign n1961 = ~n1796 & n1959;
  assign n1962 = ~n1957 & ~n31996;
  assign n1963 = ~n1955 & ~n1956;
  assign n1964 = ~n1952 & ~n31997;
  assign n1965 = ~n1950 & ~n1964;
  assign n1966 = ~n214 & ~n1965;
  assign n1967 = ~n1719 & ~n1721;
  assign n1968 = ~n1796 & n1967;
  assign n1969 = ~n31968 & ~n1968;
  assign n1970 = ~n1721 & n31968;
  assign n1971 = ~n1719 & n1970;
  assign n1972 = n31968 & n1968;
  assign n1973 = ~n1796 & n1971;
  assign n1974 = ~n1969 & ~n31998;
  assign n1975 = n214 & ~n1950;
  assign n1976 = n214 & n1965;
  assign n1977 = ~n1964 & n1975;
  assign n1978 = ~n1974 & ~n31999;
  assign n1979 = ~n1966 & ~n1978;
  assign n1980 = ~n197 & ~n1979;
  assign n1981 = n197 & ~n1966;
  assign n1982 = ~n1978 & n1981;
  assign n1983 = ~n1736 & ~n31969;
  assign n1984 = ~n1736 & ~n1796;
  assign n1985 = ~n31969 & n1984;
  assign n1986 = ~n1796 & n1983;
  assign n1987 = n31971 & ~n32000;
  assign n1988 = n1751 & n1984;
  assign n1989 = ~n31971 & n32000;
  assign n1990 = ~n1736 & n31971;
  assign n1991 = ~n31969 & n1990;
  assign n1992 = ~n1796 & n1991;
  assign n1993 = ~n31971 & ~n32000;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = ~n1987 & ~n32001;
  assign n1996 = ~n1982 & ~n32002;
  assign n1997 = ~n1980 & ~n1996;
  assign n1998 = ~n1753 & ~n1755;
  assign n1999 = ~n1796 & n1998;
  assign n2000 = ~n31973 & ~n1999;
  assign n2001 = ~n1755 & n31973;
  assign n2002 = ~n1753 & n2001;
  assign n2003 = n31973 & n1999;
  assign n2004 = ~n1796 & n2002;
  assign n2005 = ~n2000 & ~n32003;
  assign n2006 = ~n1769 & ~n31975;
  assign n2007 = ~n31975 & ~n1796;
  assign n2008 = ~n1769 & n2007;
  assign n2009 = ~n1796 & n2006;
  assign n2010 = ~n31977 & ~n32004;
  assign n2011 = ~n2005 & n2010;
  assign n2012 = ~n1997 & n2011;
  assign n2013 = n193 & ~n2012;
  assign n2014 = ~n1980 & n2005;
  assign n2015 = n1997 & n2005;
  assign n2016 = ~n1996 & n2014;
  assign n2017 = n1769 & ~n2007;
  assign n2018 = ~n193 & ~n2006;
  assign n2019 = ~n2017 & n2018;
  assign n2020 = ~n32005 & ~n2019;
  assign n2021 = ~n2013 & n2020;
  assign n2022 = pi96  & ~n2021;
  assign n2023 = ~pi94  & ~pi95 ;
  assign n2024 = ~pi96  & n2023;
  assign n2025 = ~n2022 & ~n2024;
  assign n2026 = ~n1796 & ~n2025;
  assign n2027 = ~pi96  & ~n2021;
  assign n2028 = pi97  & ~n2027;
  assign n2029 = ~pi97  & n2027;
  assign n2030 = n1798 & ~n2021;
  assign n2031 = ~n2028 & ~n32006;
  assign n2032 = ~n31945 & ~n31978;
  assign n2033 = ~n1546 & n2032;
  assign n2034 = ~n1565 & n2033;
  assign n2035 = ~n31947 & n2034;
  assign n2036 = n1551 & n1567;
  assign n2037 = ~n1559 & n2035;
  assign n2038 = ~n2024 & ~n32007;
  assign n2039 = ~n1794 & n2038;
  assign n2040 = ~n31977 & n2039;
  assign n2041 = ~n1788 & n2040;
  assign n2042 = n1796 & n2025;
  assign n2043 = ~n2022 & n2041;
  assign n2044 = n2031 & ~n32008;
  assign n2045 = ~n2026 & ~n2044;
  assign n2046 = ~n1567 & ~n2045;
  assign n2047 = n1567 & ~n2026;
  assign n2048 = ~n2044 & n2047;
  assign n2049 = ~n1796 & ~n2019;
  assign n2050 = ~n32005 & n2049;
  assign n2051 = ~n2013 & n2050;
  assign n2052 = ~n32006 & ~n2051;
  assign n2053 = pi98  & ~n2052;
  assign n2054 = ~pi98  & ~n2051;
  assign n2055 = ~pi98  & n2052;
  assign n2056 = ~n32006 & n2054;
  assign n2057 = ~n2053 & ~n32009;
  assign n2058 = ~n2048 & ~n2057;
  assign n2059 = ~n2046 & ~n2058;
  assign n2060 = ~n1374 & ~n2059;
  assign n2061 = n1374 & ~n2046;
  assign n2062 = ~n2058 & n2061;
  assign n2063 = n1374 & n2059;
  assign n2064 = ~n1801 & ~n31979;
  assign n2065 = ~n2021 & n2064;
  assign n2066 = n1818 & ~n2065;
  assign n2067 = ~n1818 & n2064;
  assign n2068 = ~n1818 & n2065;
  assign n2069 = ~n2021 & n2067;
  assign n2070 = ~n2066 & ~n32011;
  assign n2071 = ~n32010 & ~n2070;
  assign n2072 = ~n2060 & ~n2071;
  assign n2073 = ~n1179 & ~n2072;
  assign n2074 = n1179 & ~n2060;
  assign n2075 = ~n2071 & n2074;
  assign n2076 = ~n1821 & ~n31982;
  assign n2077 = ~n1821 & ~n2021;
  assign n2078 = ~n31982 & n2077;
  assign n2079 = ~n2021 & n2076;
  assign n2080 = n1830 & ~n32012;
  assign n2081 = n1834 & n2077;
  assign n2082 = n1830 & ~n31982;
  assign n2083 = ~n1821 & n2082;
  assign n2084 = ~n2021 & n2083;
  assign n2085 = ~n1830 & ~n32012;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = ~n2080 & ~n2081;
  assign n2088 = ~n2075 & ~n32013;
  assign n2089 = ~n2073 & ~n2088;
  assign n2090 = ~n1016 & ~n2089;
  assign n2091 = n1016 & ~n2073;
  assign n2092 = ~n2088 & n2091;
  assign n2093 = n1016 & n2089;
  assign n2094 = ~n1836 & ~n1838;
  assign n2095 = ~n2021 & n2094;
  assign n2096 = ~n1845 & ~n2095;
  assign n2097 = ~n1836 & n1845;
  assign n2098 = ~n1838 & n2097;
  assign n2099 = n1845 & n2095;
  assign n2100 = ~n2021 & n2098;
  assign n2101 = n1845 & ~n2095;
  assign n2102 = ~n1845 & n2095;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = ~n2096 & ~n32015;
  assign n2105 = ~n32014 & n32016;
  assign n2106 = ~n2090 & ~n2105;
  assign n2107 = ~n855 & ~n2106;
  assign n2108 = n855 & ~n2090;
  assign n2109 = ~n2105 & n2108;
  assign n2110 = ~n1848 & ~n31985;
  assign n2111 = ~n1848 & ~n2021;
  assign n2112 = ~n31985 & n2111;
  assign n2113 = ~n2021 & n2110;
  assign n2114 = n1856 & ~n32017;
  assign n2115 = n1860 & n2111;
  assign n2116 = n1856 & ~n31985;
  assign n2117 = ~n1848 & n2116;
  assign n2118 = ~n2021 & n2117;
  assign n2119 = ~n1856 & ~n32017;
  assign n2120 = ~n2118 & ~n2119;
  assign n2121 = ~n2114 & ~n2115;
  assign n2122 = ~n2109 & ~n32018;
  assign n2123 = ~n2107 & ~n2122;
  assign n2124 = ~n720 & ~n2123;
  assign n2125 = n720 & ~n2107;
  assign n2126 = ~n2122 & n2125;
  assign n2127 = n720 & n2123;
  assign n2128 = ~n1862 & ~n1864;
  assign n2129 = ~n2021 & n2128;
  assign n2130 = ~n31987 & ~n2129;
  assign n2131 = n31987 & n2129;
  assign n2132 = ~n1862 & ~n31987;
  assign n2133 = ~n1864 & n2132;
  assign n2134 = ~n2021 & n2133;
  assign n2135 = n31987 & ~n2129;
  assign n2136 = ~n2134 & ~n2135;
  assign n2137 = ~n2130 & ~n2131;
  assign n2138 = ~n32019 & ~n32020;
  assign n2139 = ~n2124 & ~n2138;
  assign n2140 = ~n592 & ~n2139;
  assign n2141 = n592 & ~n2124;
  assign n2142 = ~n2138 & n2141;
  assign n2143 = ~n1878 & ~n31989;
  assign n2144 = ~n1878 & ~n2021;
  assign n2145 = ~n31989 & n2144;
  assign n2146 = ~n2021 & n2143;
  assign n2147 = n1886 & ~n32021;
  assign n2148 = n1890 & n2144;
  assign n2149 = n1886 & ~n31989;
  assign n2150 = ~n1878 & n2149;
  assign n2151 = ~n2021 & n2150;
  assign n2152 = ~n1886 & ~n32021;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = ~n2147 & ~n2148;
  assign n2155 = ~n2142 & ~n32022;
  assign n2156 = ~n2140 & ~n2155;
  assign n2157 = ~n487 & ~n2156;
  assign n2158 = n487 & ~n2140;
  assign n2159 = ~n2155 & n2158;
  assign n2160 = n487 & n2156;
  assign n2161 = ~n1892 & ~n1894;
  assign n2162 = ~n2021 & n2161;
  assign n2163 = ~n31990 & n2162;
  assign n2164 = n31990 & ~n2162;
  assign n2165 = ~n1892 & n31990;
  assign n2166 = ~n1894 & n2165;
  assign n2167 = ~n2021 & n2166;
  assign n2168 = ~n31990 & ~n2162;
  assign n2169 = ~n2167 & ~n2168;
  assign n2170 = ~n2163 & ~n2164;
  assign n2171 = ~n32023 & ~n32024;
  assign n2172 = ~n2157 & ~n2171;
  assign n2173 = ~n393 & ~n2172;
  assign n2174 = n393 & ~n2157;
  assign n2175 = ~n2171 & n2174;
  assign n2176 = ~n1907 & ~n31992;
  assign n2177 = ~n1907 & ~n2021;
  assign n2178 = ~n31992 & n2177;
  assign n2179 = ~n2021 & n2176;
  assign n2180 = n1915 & ~n32025;
  assign n2181 = n1919 & n2177;
  assign n2182 = n1915 & ~n31992;
  assign n2183 = ~n1907 & n2182;
  assign n2184 = ~n2021 & n2183;
  assign n2185 = ~n1915 & ~n32025;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = ~n2180 & ~n2181;
  assign n2188 = ~n2175 & ~n32026;
  assign n2189 = ~n2173 & ~n2188;
  assign n2190 = ~n321 & ~n2189;
  assign n2191 = n321 & ~n2173;
  assign n2192 = ~n2188 & n2191;
  assign n2193 = n321 & n2189;
  assign n2194 = ~n1921 & ~n1923;
  assign n2195 = ~n2021 & n2194;
  assign n2196 = ~n31993 & n2195;
  assign n2197 = n31993 & ~n2195;
  assign n2198 = ~n31993 & ~n2195;
  assign n2199 = ~n1921 & n31993;
  assign n2200 = ~n1923 & n2199;
  assign n2201 = n31993 & n2195;
  assign n2202 = ~n2021 & n2200;
  assign n2203 = ~n2198 & ~n32028;
  assign n2204 = ~n2196 & ~n2197;
  assign n2205 = ~n32027 & ~n32029;
  assign n2206 = ~n2190 & ~n2205;
  assign n2207 = ~n263 & ~n2206;
  assign n2208 = n263 & ~n2190;
  assign n2209 = ~n2205 & n2208;
  assign n2210 = ~n1936 & ~n31995;
  assign n2211 = ~n1936 & ~n2021;
  assign n2212 = ~n31995 & n2211;
  assign n2213 = ~n2021 & n2210;
  assign n2214 = n1944 & ~n32030;
  assign n2215 = n1948 & n2211;
  assign n2216 = n1944 & ~n31995;
  assign n2217 = ~n1936 & n2216;
  assign n2218 = ~n2021 & n2217;
  assign n2219 = ~n1944 & ~n32030;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = ~n2214 & ~n2215;
  assign n2222 = ~n2209 & ~n32031;
  assign n2223 = ~n2207 & ~n2222;
  assign n2224 = ~n214 & ~n2223;
  assign n2225 = n214 & ~n2207;
  assign n2226 = ~n2222 & n2225;
  assign n2227 = n214 & n2223;
  assign n2228 = ~n1950 & ~n1952;
  assign n2229 = ~n1950 & ~n2021;
  assign n2230 = ~n1952 & n2229;
  assign n2231 = ~n2021 & n2228;
  assign n2232 = n31997 & ~n32033;
  assign n2233 = n1964 & n2229;
  assign n2234 = ~n31997 & n32033;
  assign n2235 = ~n1950 & n31997;
  assign n2236 = ~n1952 & n2235;
  assign n2237 = ~n2021 & n2236;
  assign n2238 = ~n31997 & ~n32033;
  assign n2239 = ~n2237 & ~n2238;
  assign n2240 = ~n2232 & ~n32034;
  assign n2241 = ~n32032 & ~n32035;
  assign n2242 = ~n2224 & ~n2241;
  assign n2243 = ~n197 & ~n2242;
  assign n2244 = n197 & ~n2224;
  assign n2245 = ~n2241 & n2244;
  assign n2246 = ~n1966 & ~n31999;
  assign n2247 = ~n1966 & ~n2021;
  assign n2248 = ~n31999 & n2247;
  assign n2249 = ~n2021 & n2246;
  assign n2250 = n1974 & ~n32036;
  assign n2251 = n1978 & n2247;
  assign n2252 = n1974 & ~n31999;
  assign n2253 = ~n1966 & n2252;
  assign n2254 = ~n2021 & n2253;
  assign n2255 = ~n1974 & ~n32036;
  assign n2256 = ~n2254 & ~n2255;
  assign n2257 = ~n2250 & ~n2251;
  assign n2258 = ~n2245 & ~n32037;
  assign n2259 = ~n2243 & ~n2258;
  assign n2260 = ~n1980 & ~n1982;
  assign n2261 = ~n2021 & n2260;
  assign n2262 = ~n32002 & ~n2261;
  assign n2263 = ~n1980 & n32002;
  assign n2264 = ~n1982 & n2263;
  assign n2265 = n32002 & n2261;
  assign n2266 = ~n2021 & n2264;
  assign n2267 = ~n2262 & ~n32038;
  assign n2268 = ~n1997 & ~n2005;
  assign n2269 = ~n2005 & ~n2021;
  assign n2270 = ~n1997 & n2269;
  assign n2271 = ~n2021 & n2268;
  assign n2272 = ~n32005 & ~n32039;
  assign n2273 = ~n2267 & n2272;
  assign n2274 = ~n2259 & n2273;
  assign n2275 = n193 & ~n2274;
  assign n2276 = ~n2243 & n2267;
  assign n2277 = ~n2258 & n2276;
  assign n2278 = n2259 & n2267;
  assign n2279 = n1997 & ~n2269;
  assign n2280 = ~n193 & ~n2268;
  assign n2281 = ~n2279 & n2280;
  assign n2282 = ~n32040 & ~n2281;
  assign n2283 = ~n2275 & n2282;
  assign n2284 = pi94  & ~n2283;
  assign n2285 = ~pi92  & ~pi93 ;
  assign n2286 = ~pi94  & n2285;
  assign n2287 = ~n2284 & ~n2286;
  assign n2288 = ~n2021 & ~n2287;
  assign n2289 = ~n31974 & ~n32007;
  assign n2290 = ~n1774 & n2289;
  assign n2291 = ~n1794 & n2290;
  assign n2292 = ~n31977 & n2291;
  assign n2293 = n31975 & n1796;
  assign n2294 = ~n1788 & n2292;
  assign n2295 = ~n2286 & ~n32041;
  assign n2296 = ~n2019 & n2295;
  assign n2297 = ~n32005 & n2296;
  assign n2298 = ~n2013 & n2297;
  assign n2299 = n2021 & n2287;
  assign n2300 = ~n2284 & n2298;
  assign n2301 = ~pi94  & ~n2283;
  assign n2302 = pi95  & ~n2301;
  assign n2303 = ~pi95  & n2301;
  assign n2304 = n2023 & ~n2283;
  assign n2305 = ~n2302 & ~n32043;
  assign n2306 = ~n32042 & n2305;
  assign n2307 = ~n2288 & ~n2306;
  assign n2308 = ~n1796 & ~n2307;
  assign n2309 = ~n2021 & ~n2281;
  assign n2310 = ~n32040 & n2309;
  assign n2311 = ~n2275 & n2310;
  assign n2312 = ~n32043 & ~n2311;
  assign n2313 = pi96  & ~n2312;
  assign n2314 = ~pi96  & ~n2311;
  assign n2315 = ~pi96  & n2312;
  assign n2316 = ~n32043 & n2314;
  assign n2317 = ~n2313 & ~n32044;
  assign n2318 = n1796 & ~n2288;
  assign n2319 = n1796 & n2307;
  assign n2320 = ~n2306 & n2318;
  assign n2321 = ~n2317 & ~n32045;
  assign n2322 = ~n2308 & ~n2321;
  assign n2323 = ~n1567 & ~n2322;
  assign n2324 = n1567 & ~n2308;
  assign n2325 = ~n2321 & n2324;
  assign n2326 = ~n2026 & ~n32008;
  assign n2327 = ~n2283 & n2326;
  assign n2328 = n2031 & ~n2327;
  assign n2329 = ~n2031 & ~n32008;
  assign n2330 = ~n2026 & n2329;
  assign n2331 = ~n2031 & n2327;
  assign n2332 = ~n2283 & n2330;
  assign n2333 = ~n2328 & ~n32046;
  assign n2334 = ~n2325 & ~n2333;
  assign n2335 = ~n2323 & ~n2334;
  assign n2336 = ~n1374 & ~n2335;
  assign n2337 = ~n2046 & ~n2048;
  assign n2338 = ~n2283 & n2337;
  assign n2339 = ~n2057 & ~n2338;
  assign n2340 = ~n2048 & n2057;
  assign n2341 = ~n2046 & n2340;
  assign n2342 = n2057 & n2338;
  assign n2343 = ~n2283 & n2341;
  assign n2344 = ~n2339 & ~n32047;
  assign n2345 = n1374 & ~n2323;
  assign n2346 = n1374 & n2335;
  assign n2347 = ~n2334 & n2345;
  assign n2348 = ~n2344 & ~n32048;
  assign n2349 = ~n2336 & ~n2348;
  assign n2350 = ~n1179 & ~n2349;
  assign n2351 = n1179 & ~n2336;
  assign n2352 = ~n2348 & n2351;
  assign n2353 = ~n2060 & ~n32010;
  assign n2354 = ~n2283 & n2353;
  assign n2355 = ~n2070 & ~n2354;
  assign n2356 = ~n2060 & n2070;
  assign n2357 = ~n32010 & n2356;
  assign n2358 = n2070 & n2354;
  assign n2359 = ~n2283 & n2357;
  assign n2360 = n2070 & ~n2354;
  assign n2361 = ~n2070 & n2354;
  assign n2362 = ~n2360 & ~n2361;
  assign n2363 = ~n2355 & ~n32049;
  assign n2364 = ~n2352 & n32050;
  assign n2365 = ~n2350 & ~n2364;
  assign n2366 = ~n1016 & ~n2365;
  assign n2367 = ~n2073 & ~n2075;
  assign n2368 = ~n2283 & n2367;
  assign n2369 = ~n32013 & ~n2368;
  assign n2370 = ~n2075 & n32013;
  assign n2371 = ~n2073 & n2370;
  assign n2372 = n32013 & n2368;
  assign n2373 = ~n2283 & n2371;
  assign n2374 = ~n2369 & ~n32051;
  assign n2375 = n1016 & ~n2350;
  assign n2376 = n1016 & n2365;
  assign n2377 = ~n2364 & n2375;
  assign n2378 = ~n2374 & ~n32052;
  assign n2379 = ~n2366 & ~n2378;
  assign n2380 = ~n855 & ~n2379;
  assign n2381 = n855 & ~n2366;
  assign n2382 = ~n2378 & n2381;
  assign n2383 = ~n2090 & ~n32014;
  assign n2384 = ~n2283 & n2383;
  assign n2385 = ~n32016 & ~n2384;
  assign n2386 = n32016 & n2384;
  assign n2387 = ~n2090 & ~n32016;
  assign n2388 = ~n32014 & n2387;
  assign n2389 = ~n2283 & n2388;
  assign n2390 = n32016 & ~n2384;
  assign n2391 = ~n2389 & ~n2390;
  assign n2392 = ~n2385 & ~n2386;
  assign n2393 = ~n2382 & ~n32053;
  assign n2394 = ~n2380 & ~n2393;
  assign n2395 = ~n720 & ~n2394;
  assign n2396 = ~n2107 & ~n2109;
  assign n2397 = ~n2283 & n2396;
  assign n2398 = ~n32018 & ~n2397;
  assign n2399 = ~n2109 & n32018;
  assign n2400 = ~n2107 & n2399;
  assign n2401 = n32018 & n2397;
  assign n2402 = ~n2283 & n2400;
  assign n2403 = ~n2398 & ~n32054;
  assign n2404 = n720 & ~n2380;
  assign n2405 = n720 & n2394;
  assign n2406 = ~n2393 & n2404;
  assign n2407 = ~n2403 & ~n32055;
  assign n2408 = ~n2395 & ~n2407;
  assign n2409 = ~n592 & ~n2408;
  assign n2410 = n592 & ~n2395;
  assign n2411 = ~n2407 & n2410;
  assign n2412 = ~n2124 & ~n32019;
  assign n2413 = ~n2283 & n2412;
  assign n2414 = ~n32020 & n2413;
  assign n2415 = n32020 & ~n2413;
  assign n2416 = ~n2124 & n32020;
  assign n2417 = ~n32019 & n2416;
  assign n2418 = ~n2283 & n2417;
  assign n2419 = ~n32020 & ~n2413;
  assign n2420 = ~n2418 & ~n2419;
  assign n2421 = ~n2414 & ~n2415;
  assign n2422 = ~n2411 & ~n32056;
  assign n2423 = ~n2409 & ~n2422;
  assign n2424 = ~n487 & ~n2423;
  assign n2425 = ~n2140 & ~n2142;
  assign n2426 = ~n2283 & n2425;
  assign n2427 = ~n32022 & ~n2426;
  assign n2428 = ~n2142 & n32022;
  assign n2429 = ~n2140 & n2428;
  assign n2430 = n32022 & n2426;
  assign n2431 = ~n2283 & n2429;
  assign n2432 = ~n2427 & ~n32057;
  assign n2433 = n487 & ~n2409;
  assign n2434 = n487 & n2423;
  assign n2435 = ~n2422 & n2433;
  assign n2436 = ~n2432 & ~n32058;
  assign n2437 = ~n2424 & ~n2436;
  assign n2438 = ~n393 & ~n2437;
  assign n2439 = n393 & ~n2424;
  assign n2440 = ~n2436 & n2439;
  assign n2441 = ~n2157 & ~n32023;
  assign n2442 = ~n2283 & n2441;
  assign n2443 = ~n32024 & n2442;
  assign n2444 = n32024 & ~n2442;
  assign n2445 = ~n32024 & ~n2442;
  assign n2446 = ~n2157 & n32024;
  assign n2447 = ~n32023 & n2446;
  assign n2448 = n32024 & n2442;
  assign n2449 = ~n2283 & n2447;
  assign n2450 = ~n2445 & ~n32059;
  assign n2451 = ~n2443 & ~n2444;
  assign n2452 = ~n2440 & ~n32060;
  assign n2453 = ~n2438 & ~n2452;
  assign n2454 = ~n321 & ~n2453;
  assign n2455 = ~n2173 & ~n2175;
  assign n2456 = ~n2283 & n2455;
  assign n2457 = ~n32026 & ~n2456;
  assign n2458 = ~n2175 & n32026;
  assign n2459 = ~n2173 & n2458;
  assign n2460 = n32026 & n2456;
  assign n2461 = ~n2283 & n2459;
  assign n2462 = ~n2457 & ~n32061;
  assign n2463 = n321 & ~n2438;
  assign n2464 = n321 & n2453;
  assign n2465 = ~n2452 & n2463;
  assign n2466 = ~n2462 & ~n32062;
  assign n2467 = ~n2454 & ~n2466;
  assign n2468 = ~n263 & ~n2467;
  assign n2469 = n263 & ~n2454;
  assign n2470 = ~n2466 & n2469;
  assign n2471 = ~n2190 & ~n32027;
  assign n2472 = ~n2190 & ~n2283;
  assign n2473 = ~n32027 & n2472;
  assign n2474 = ~n2283 & n2471;
  assign n2475 = n32029 & ~n32063;
  assign n2476 = n2205 & n2472;
  assign n2477 = ~n32029 & n32063;
  assign n2478 = ~n2190 & n32029;
  assign n2479 = ~n32027 & n2478;
  assign n2480 = ~n2283 & n2479;
  assign n2481 = ~n32029 & ~n32063;
  assign n2482 = ~n2480 & ~n2481;
  assign n2483 = ~n2475 & ~n32064;
  assign n2484 = ~n2470 & ~n32065;
  assign n2485 = ~n2468 & ~n2484;
  assign n2486 = ~n214 & ~n2485;
  assign n2487 = ~n2207 & ~n2209;
  assign n2488 = ~n2283 & n2487;
  assign n2489 = ~n32031 & ~n2488;
  assign n2490 = ~n2209 & n32031;
  assign n2491 = ~n2207 & n2490;
  assign n2492 = n32031 & n2488;
  assign n2493 = ~n2283 & n2491;
  assign n2494 = ~n2489 & ~n32066;
  assign n2495 = n214 & ~n2468;
  assign n2496 = n214 & n2485;
  assign n2497 = ~n2484 & n2495;
  assign n2498 = ~n2494 & ~n32067;
  assign n2499 = ~n2486 & ~n2498;
  assign n2500 = ~n197 & ~n2499;
  assign n2501 = ~n2224 & ~n32032;
  assign n2502 = ~n2283 & n2501;
  assign n2503 = ~n32035 & ~n2502;
  assign n2504 = ~n2224 & n32035;
  assign n2505 = ~n32032 & n2504;
  assign n2506 = n32035 & n2502;
  assign n2507 = ~n2283 & n2505;
  assign n2508 = ~n2503 & ~n32068;
  assign n2509 = n197 & ~n2486;
  assign n2510 = ~n2498 & n2509;
  assign n2511 = ~n2508 & ~n2510;
  assign n2512 = ~n2500 & ~n2511;
  assign n2513 = ~n2243 & ~n2245;
  assign n2514 = ~n2283 & n2513;
  assign n2515 = ~n32037 & ~n2514;
  assign n2516 = ~n2245 & n32037;
  assign n2517 = ~n2243 & n2516;
  assign n2518 = n32037 & n2514;
  assign n2519 = ~n2283 & n2517;
  assign n2520 = ~n2515 & ~n32069;
  assign n2521 = ~n2259 & ~n2267;
  assign n2522 = ~n2267 & ~n2283;
  assign n2523 = ~n2259 & n2522;
  assign n2524 = ~n2283 & n2521;
  assign n2525 = ~n32040 & ~n32070;
  assign n2526 = ~n2520 & n2525;
  assign n2527 = ~n2512 & n2526;
  assign n2528 = n193 & ~n2527;
  assign n2529 = ~n2500 & n2520;
  assign n2530 = n2512 & n2520;
  assign n2531 = ~n2511 & n2529;
  assign n2532 = n2259 & ~n2522;
  assign n2533 = ~n193 & ~n2521;
  assign n2534 = ~n2532 & n2533;
  assign n2535 = ~n32071 & ~n2534;
  assign n2536 = ~n2528 & n2535;
  assign n2537 = pi92  & ~n2536;
  assign n2538 = ~pi90  & ~pi91 ;
  assign n2539 = ~pi92  & n2538;
  assign n2540 = ~n2537 & ~n2539;
  assign n2541 = ~n2283 & ~n2540;
  assign n2542 = ~pi92  & ~n2536;
  assign n2543 = pi93  & ~n2542;
  assign n2544 = ~pi93  & n2542;
  assign n2545 = n2285 & ~n2536;
  assign n2546 = ~n2543 & ~n32072;
  assign n2547 = ~n32003 & ~n32041;
  assign n2548 = ~n2000 & n2547;
  assign n2549 = ~n2019 & n2548;
  assign n2550 = ~n32005 & n2549;
  assign n2551 = n2005 & n2021;
  assign n2552 = ~n2013 & n2550;
  assign n2553 = ~n2539 & ~n32073;
  assign n2554 = ~n2281 & n2553;
  assign n2555 = ~n32040 & n2554;
  assign n2556 = ~n2275 & n2555;
  assign n2557 = n2283 & n2540;
  assign n2558 = ~n2537 & n2556;
  assign n2559 = n2546 & ~n32074;
  assign n2560 = ~n2541 & ~n2559;
  assign n2561 = ~n2021 & ~n2560;
  assign n2562 = n2021 & ~n2541;
  assign n2563 = ~n2559 & n2562;
  assign n2564 = ~n2283 & ~n2534;
  assign n2565 = ~n32071 & n2564;
  assign n2566 = ~n2528 & n2565;
  assign n2567 = ~n32072 & ~n2566;
  assign n2568 = pi94  & ~n2567;
  assign n2569 = ~pi94  & ~n2566;
  assign n2570 = ~pi94  & n2567;
  assign n2571 = ~n32072 & n2569;
  assign n2572 = ~n2568 & ~n32075;
  assign n2573 = ~n2563 & ~n2572;
  assign n2574 = ~n2561 & ~n2573;
  assign n2575 = ~n1796 & ~n2574;
  assign n2576 = n1796 & ~n2561;
  assign n2577 = ~n2573 & n2576;
  assign n2578 = n1796 & n2574;
  assign n2579 = ~n2288 & ~n32042;
  assign n2580 = ~n2536 & n2579;
  assign n2581 = n2305 & ~n2580;
  assign n2582 = ~n2305 & n2579;
  assign n2583 = ~n2305 & n2580;
  assign n2584 = ~n2536 & n2582;
  assign n2585 = ~n2581 & ~n32077;
  assign n2586 = ~n32076 & ~n2585;
  assign n2587 = ~n2575 & ~n2586;
  assign n2588 = ~n1567 & ~n2587;
  assign n2589 = n1567 & ~n2575;
  assign n2590 = ~n2586 & n2589;
  assign n2591 = ~n2308 & ~n32045;
  assign n2592 = ~n2308 & ~n2536;
  assign n2593 = ~n32045 & n2592;
  assign n2594 = ~n2536 & n2591;
  assign n2595 = n2317 & ~n32078;
  assign n2596 = n2321 & n2592;
  assign n2597 = n2317 & ~n32045;
  assign n2598 = ~n2308 & n2597;
  assign n2599 = ~n2536 & n2598;
  assign n2600 = ~n2317 & ~n32078;
  assign n2601 = ~n2599 & ~n2600;
  assign n2602 = ~n2595 & ~n2596;
  assign n2603 = ~n2590 & ~n32079;
  assign n2604 = ~n2588 & ~n2603;
  assign n2605 = ~n1374 & ~n2604;
  assign n2606 = n1374 & ~n2588;
  assign n2607 = ~n2603 & n2606;
  assign n2608 = n1374 & n2604;
  assign n2609 = ~n2323 & ~n2325;
  assign n2610 = ~n2536 & n2609;
  assign n2611 = ~n2333 & ~n2610;
  assign n2612 = ~n2323 & n2333;
  assign n2613 = ~n2325 & n2612;
  assign n2614 = n2333 & n2610;
  assign n2615 = ~n2536 & n2613;
  assign n2616 = n2333 & ~n2610;
  assign n2617 = ~n2333 & n2610;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = ~n2611 & ~n32081;
  assign n2620 = ~n32080 & n32082;
  assign n2621 = ~n2605 & ~n2620;
  assign n2622 = ~n1179 & ~n2621;
  assign n2623 = n1179 & ~n2605;
  assign n2624 = ~n2620 & n2623;
  assign n2625 = ~n2336 & ~n32048;
  assign n2626 = ~n2336 & ~n2536;
  assign n2627 = ~n32048 & n2626;
  assign n2628 = ~n2536 & n2625;
  assign n2629 = n2344 & ~n32083;
  assign n2630 = n2348 & n2626;
  assign n2631 = n2344 & ~n32048;
  assign n2632 = ~n2336 & n2631;
  assign n2633 = ~n2536 & n2632;
  assign n2634 = ~n2344 & ~n32083;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = ~n2629 & ~n2630;
  assign n2637 = ~n2624 & ~n32084;
  assign n2638 = ~n2622 & ~n2637;
  assign n2639 = ~n1016 & ~n2638;
  assign n2640 = n1016 & ~n2622;
  assign n2641 = ~n2637 & n2640;
  assign n2642 = n1016 & n2638;
  assign n2643 = ~n2350 & ~n2352;
  assign n2644 = ~n2536 & n2643;
  assign n2645 = ~n32050 & ~n2644;
  assign n2646 = n32050 & n2644;
  assign n2647 = ~n2350 & ~n32050;
  assign n2648 = ~n2352 & n2647;
  assign n2649 = ~n2536 & n2648;
  assign n2650 = n32050 & ~n2644;
  assign n2651 = ~n2649 & ~n2650;
  assign n2652 = ~n2645 & ~n2646;
  assign n2653 = ~n32085 & ~n32086;
  assign n2654 = ~n2639 & ~n2653;
  assign n2655 = ~n855 & ~n2654;
  assign n2656 = n855 & ~n2639;
  assign n2657 = ~n2653 & n2656;
  assign n2658 = ~n2366 & ~n32052;
  assign n2659 = ~n2366 & ~n2536;
  assign n2660 = ~n32052 & n2659;
  assign n2661 = ~n2536 & n2658;
  assign n2662 = n2374 & ~n32087;
  assign n2663 = n2378 & n2659;
  assign n2664 = n2374 & ~n32052;
  assign n2665 = ~n2366 & n2664;
  assign n2666 = ~n2536 & n2665;
  assign n2667 = ~n2374 & ~n32087;
  assign n2668 = ~n2666 & ~n2667;
  assign n2669 = ~n2662 & ~n2663;
  assign n2670 = ~n2657 & ~n32088;
  assign n2671 = ~n2655 & ~n2670;
  assign n2672 = ~n720 & ~n2671;
  assign n2673 = n720 & ~n2655;
  assign n2674 = ~n2670 & n2673;
  assign n2675 = n720 & n2671;
  assign n2676 = ~n2380 & ~n2382;
  assign n2677 = ~n2536 & n2676;
  assign n2678 = ~n32053 & n2677;
  assign n2679 = n32053 & ~n2677;
  assign n2680 = ~n2380 & n32053;
  assign n2681 = ~n2382 & n2680;
  assign n2682 = ~n2536 & n2681;
  assign n2683 = ~n32053 & ~n2677;
  assign n2684 = ~n2682 & ~n2683;
  assign n2685 = ~n2678 & ~n2679;
  assign n2686 = ~n32089 & ~n32090;
  assign n2687 = ~n2672 & ~n2686;
  assign n2688 = ~n592 & ~n2687;
  assign n2689 = n592 & ~n2672;
  assign n2690 = ~n2686 & n2689;
  assign n2691 = ~n2395 & ~n32055;
  assign n2692 = ~n2395 & ~n2536;
  assign n2693 = ~n32055 & n2692;
  assign n2694 = ~n2536 & n2691;
  assign n2695 = n2403 & ~n32091;
  assign n2696 = n2407 & n2692;
  assign n2697 = n2403 & ~n32055;
  assign n2698 = ~n2395 & n2697;
  assign n2699 = ~n2536 & n2698;
  assign n2700 = ~n2403 & ~n32091;
  assign n2701 = ~n2699 & ~n2700;
  assign n2702 = ~n2695 & ~n2696;
  assign n2703 = ~n2690 & ~n32092;
  assign n2704 = ~n2688 & ~n2703;
  assign n2705 = ~n487 & ~n2704;
  assign n2706 = n487 & ~n2688;
  assign n2707 = ~n2703 & n2706;
  assign n2708 = n487 & n2704;
  assign n2709 = ~n2409 & ~n2411;
  assign n2710 = ~n2536 & n2709;
  assign n2711 = ~n32056 & n2710;
  assign n2712 = n32056 & ~n2710;
  assign n2713 = ~n32056 & ~n2710;
  assign n2714 = ~n2409 & n32056;
  assign n2715 = ~n2411 & n2714;
  assign n2716 = n32056 & n2710;
  assign n2717 = ~n2536 & n2715;
  assign n2718 = ~n2713 & ~n32094;
  assign n2719 = ~n2711 & ~n2712;
  assign n2720 = ~n32093 & ~n32095;
  assign n2721 = ~n2705 & ~n2720;
  assign n2722 = ~n393 & ~n2721;
  assign n2723 = n393 & ~n2705;
  assign n2724 = ~n2720 & n2723;
  assign n2725 = ~n2424 & ~n32058;
  assign n2726 = ~n2424 & ~n2536;
  assign n2727 = ~n32058 & n2726;
  assign n2728 = ~n2536 & n2725;
  assign n2729 = n2432 & ~n32096;
  assign n2730 = n2436 & n2726;
  assign n2731 = n2432 & ~n32058;
  assign n2732 = ~n2424 & n2731;
  assign n2733 = ~n2536 & n2732;
  assign n2734 = ~n2432 & ~n32096;
  assign n2735 = ~n2733 & ~n2734;
  assign n2736 = ~n2729 & ~n2730;
  assign n2737 = ~n2724 & ~n32097;
  assign n2738 = ~n2722 & ~n2737;
  assign n2739 = ~n321 & ~n2738;
  assign n2740 = n321 & ~n2722;
  assign n2741 = ~n2737 & n2740;
  assign n2742 = n321 & n2738;
  assign n2743 = ~n2438 & ~n2440;
  assign n2744 = ~n2438 & ~n2536;
  assign n2745 = ~n2440 & n2744;
  assign n2746 = ~n2536 & n2743;
  assign n2747 = n32060 & ~n32099;
  assign n2748 = n2452 & n2744;
  assign n2749 = ~n32060 & n32099;
  assign n2750 = ~n2438 & n32060;
  assign n2751 = ~n2440 & n2750;
  assign n2752 = ~n2536 & n2751;
  assign n2753 = ~n32060 & ~n32099;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = ~n2747 & ~n32100;
  assign n2756 = ~n32098 & ~n32101;
  assign n2757 = ~n2739 & ~n2756;
  assign n2758 = ~n263 & ~n2757;
  assign n2759 = n263 & ~n2739;
  assign n2760 = ~n2756 & n2759;
  assign n2761 = ~n2454 & ~n32062;
  assign n2762 = ~n2454 & ~n2536;
  assign n2763 = ~n32062 & n2762;
  assign n2764 = ~n2536 & n2761;
  assign n2765 = n2462 & ~n32102;
  assign n2766 = n2466 & n2762;
  assign n2767 = n2462 & ~n32062;
  assign n2768 = ~n2454 & n2767;
  assign n2769 = ~n2536 & n2768;
  assign n2770 = ~n2462 & ~n32102;
  assign n2771 = ~n2769 & ~n2770;
  assign n2772 = ~n2765 & ~n2766;
  assign n2773 = ~n2760 & ~n32103;
  assign n2774 = ~n2758 & ~n2773;
  assign n2775 = ~n214 & ~n2774;
  assign n2776 = ~n2468 & ~n2470;
  assign n2777 = ~n2536 & n2776;
  assign n2778 = ~n32065 & ~n2777;
  assign n2779 = ~n2468 & n32065;
  assign n2780 = ~n2470 & n2779;
  assign n2781 = n32065 & n2777;
  assign n2782 = ~n2536 & n2780;
  assign n2783 = ~n2778 & ~n32104;
  assign n2784 = n214 & ~n2758;
  assign n2785 = ~n2773 & n2784;
  assign n2786 = n214 & n2774;
  assign n2787 = ~n2783 & ~n32105;
  assign n2788 = ~n2775 & ~n2787;
  assign n2789 = ~n197 & ~n2788;
  assign n2790 = n197 & ~n2775;
  assign n2791 = ~n2787 & n2790;
  assign n2792 = ~n2486 & ~n32067;
  assign n2793 = ~n2486 & ~n2536;
  assign n2794 = ~n32067 & n2793;
  assign n2795 = ~n2536 & n2792;
  assign n2796 = n2494 & ~n32106;
  assign n2797 = n2498 & n2793;
  assign n2798 = n2494 & ~n32067;
  assign n2799 = ~n2486 & n2798;
  assign n2800 = ~n2536 & n2799;
  assign n2801 = ~n2494 & ~n32106;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = ~n2796 & ~n2797;
  assign n2804 = ~n2791 & ~n32107;
  assign n2805 = ~n2789 & ~n2804;
  assign n2806 = ~n2500 & ~n2510;
  assign n2807 = ~n2500 & ~n2536;
  assign n2808 = ~n2510 & n2807;
  assign n2809 = ~n2536 & n2806;
  assign n2810 = n2508 & ~n32108;
  assign n2811 = n2511 & n2807;
  assign n2812 = ~n2500 & n2508;
  assign n2813 = ~n2510 & n2812;
  assign n2814 = ~n2536 & n2813;
  assign n2815 = ~n2508 & ~n32108;
  assign n2816 = ~n2814 & ~n2815;
  assign n2817 = ~n2810 & ~n2811;
  assign n2818 = ~n2512 & ~n2520;
  assign n2819 = ~n2520 & ~n2536;
  assign n2820 = ~n2512 & n2819;
  assign n2821 = ~n2536 & n2818;
  assign n2822 = ~n32071 & ~n32110;
  assign n2823 = ~n32109 & n2822;
  assign n2824 = ~n2805 & n2823;
  assign n2825 = n193 & ~n2824;
  assign n2826 = ~n2789 & n32109;
  assign n2827 = ~n2804 & n2826;
  assign n2828 = n2805 & n32109;
  assign n2829 = n2512 & ~n2819;
  assign n2830 = ~n193 & ~n2818;
  assign n2831 = ~n2829 & n2830;
  assign n2832 = ~n32111 & ~n2831;
  assign n2833 = ~n2825 & n2832;
  assign n2834 = pi90  & ~n2833;
  assign n2835 = ~pi88  & ~pi89 ;
  assign n2836 = ~pi90  & n2835;
  assign n2837 = ~n2834 & ~n2836;
  assign n2838 = ~n2536 & ~n2837;
  assign n2839 = ~n32038 & ~n32073;
  assign n2840 = ~n2262 & n2839;
  assign n2841 = ~n2281 & n2840;
  assign n2842 = ~n32040 & n2841;
  assign n2843 = n2267 & n2283;
  assign n2844 = ~n2275 & n2842;
  assign n2845 = ~n2836 & ~n32112;
  assign n2846 = ~n2534 & n2845;
  assign n2847 = ~n32071 & n2846;
  assign n2848 = ~n2528 & n2847;
  assign n2849 = n2536 & n2837;
  assign n2850 = ~n2834 & n2848;
  assign n2851 = ~pi90  & ~n2833;
  assign n2852 = pi91  & ~n2851;
  assign n2853 = ~pi91  & n2851;
  assign n2854 = n2538 & ~n2833;
  assign n2855 = ~n2852 & ~n32114;
  assign n2856 = ~n32113 & n2855;
  assign n2857 = ~n2838 & ~n2856;
  assign n2858 = ~n2283 & ~n2857;
  assign n2859 = ~n2536 & ~n2831;
  assign n2860 = ~n32111 & n2859;
  assign n2861 = ~n2825 & n2860;
  assign n2862 = ~n32114 & ~n2861;
  assign n2863 = pi92  & ~n2862;
  assign n2864 = ~pi92  & ~n2861;
  assign n2865 = ~pi92  & n2862;
  assign n2866 = ~n32114 & n2864;
  assign n2867 = ~n2863 & ~n32115;
  assign n2868 = n2283 & ~n2838;
  assign n2869 = n2283 & n2857;
  assign n2870 = ~n2856 & n2868;
  assign n2871 = ~n2867 & ~n32116;
  assign n2872 = ~n2858 & ~n2871;
  assign n2873 = ~n2021 & ~n2872;
  assign n2874 = n2021 & ~n2858;
  assign n2875 = ~n2871 & n2874;
  assign n2876 = ~n2541 & ~n32074;
  assign n2877 = ~n2833 & n2876;
  assign n2878 = n2546 & ~n2877;
  assign n2879 = ~n2546 & n2876;
  assign n2880 = ~n2546 & n2877;
  assign n2881 = ~n2833 & n2879;
  assign n2882 = ~n2878 & ~n32117;
  assign n2883 = ~n2875 & ~n2882;
  assign n2884 = ~n2873 & ~n2883;
  assign n2885 = ~n1796 & ~n2884;
  assign n2886 = ~n2561 & ~n2563;
  assign n2887 = ~n2833 & n2886;
  assign n2888 = ~n2572 & ~n2887;
  assign n2889 = ~n2563 & n2572;
  assign n2890 = ~n2561 & n2889;
  assign n2891 = n2572 & n2887;
  assign n2892 = ~n2833 & n2890;
  assign n2893 = ~n2888 & ~n32118;
  assign n2894 = n1796 & ~n2873;
  assign n2895 = n1796 & n2884;
  assign n2896 = ~n2883 & n2894;
  assign n2897 = ~n2893 & ~n32119;
  assign n2898 = ~n2885 & ~n2897;
  assign n2899 = ~n1567 & ~n2898;
  assign n2900 = n1567 & ~n2885;
  assign n2901 = ~n2897 & n2900;
  assign n2902 = ~n2575 & ~n32076;
  assign n2903 = ~n2833 & n2902;
  assign n2904 = ~n2585 & ~n2903;
  assign n2905 = ~n2575 & n2585;
  assign n2906 = ~n32076 & n2905;
  assign n2907 = n2585 & n2903;
  assign n2908 = ~n2833 & n2906;
  assign n2909 = n2585 & ~n2903;
  assign n2910 = ~n2585 & n2903;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912 = ~n2904 & ~n32120;
  assign n2913 = ~n2901 & n32121;
  assign n2914 = ~n2899 & ~n2913;
  assign n2915 = ~n1374 & ~n2914;
  assign n2916 = ~n2588 & ~n2590;
  assign n2917 = ~n2833 & n2916;
  assign n2918 = ~n32079 & ~n2917;
  assign n2919 = ~n2590 & n32079;
  assign n2920 = ~n2588 & n2919;
  assign n2921 = n32079 & n2917;
  assign n2922 = ~n2833 & n2920;
  assign n2923 = ~n2918 & ~n32122;
  assign n2924 = n1374 & ~n2899;
  assign n2925 = n1374 & n2914;
  assign n2926 = ~n2913 & n2924;
  assign n2927 = ~n2923 & ~n32123;
  assign n2928 = ~n2915 & ~n2927;
  assign n2929 = ~n1179 & ~n2928;
  assign n2930 = n1179 & ~n2915;
  assign n2931 = ~n2927 & n2930;
  assign n2932 = ~n2605 & ~n32080;
  assign n2933 = ~n2833 & n2932;
  assign n2934 = ~n32082 & ~n2933;
  assign n2935 = n32082 & n2933;
  assign n2936 = ~n2605 & ~n32082;
  assign n2937 = ~n32080 & n2936;
  assign n2938 = ~n2833 & n2937;
  assign n2939 = n32082 & ~n2933;
  assign n2940 = ~n2938 & ~n2939;
  assign n2941 = ~n2934 & ~n2935;
  assign n2942 = ~n2931 & ~n32124;
  assign n2943 = ~n2929 & ~n2942;
  assign n2944 = ~n1016 & ~n2943;
  assign n2945 = ~n2622 & ~n2624;
  assign n2946 = ~n2833 & n2945;
  assign n2947 = ~n32084 & ~n2946;
  assign n2948 = ~n2624 & n32084;
  assign n2949 = ~n2622 & n2948;
  assign n2950 = n32084 & n2946;
  assign n2951 = ~n2833 & n2949;
  assign n2952 = ~n2947 & ~n32125;
  assign n2953 = n1016 & ~n2929;
  assign n2954 = n1016 & n2943;
  assign n2955 = ~n2942 & n2953;
  assign n2956 = ~n2952 & ~n32126;
  assign n2957 = ~n2944 & ~n2956;
  assign n2958 = ~n855 & ~n2957;
  assign n2959 = n855 & ~n2944;
  assign n2960 = ~n2956 & n2959;
  assign n2961 = ~n2639 & ~n32085;
  assign n2962 = ~n2833 & n2961;
  assign n2963 = ~n32086 & n2962;
  assign n2964 = n32086 & ~n2962;
  assign n2965 = ~n2639 & n32086;
  assign n2966 = ~n32085 & n2965;
  assign n2967 = ~n2833 & n2966;
  assign n2968 = ~n32086 & ~n2962;
  assign n2969 = ~n2967 & ~n2968;
  assign n2970 = ~n2963 & ~n2964;
  assign n2971 = ~n2960 & ~n32127;
  assign n2972 = ~n2958 & ~n2971;
  assign n2973 = ~n720 & ~n2972;
  assign n2974 = ~n2655 & ~n2657;
  assign n2975 = ~n2833 & n2974;
  assign n2976 = ~n32088 & ~n2975;
  assign n2977 = ~n2657 & n32088;
  assign n2978 = ~n2655 & n2977;
  assign n2979 = n32088 & n2975;
  assign n2980 = ~n2833 & n2978;
  assign n2981 = ~n2976 & ~n32128;
  assign n2982 = n720 & ~n2958;
  assign n2983 = n720 & n2972;
  assign n2984 = ~n2971 & n2982;
  assign n2985 = ~n2981 & ~n32129;
  assign n2986 = ~n2973 & ~n2985;
  assign n2987 = ~n592 & ~n2986;
  assign n2988 = n592 & ~n2973;
  assign n2989 = ~n2985 & n2988;
  assign n2990 = ~n2672 & ~n32089;
  assign n2991 = ~n2833 & n2990;
  assign n2992 = ~n32090 & n2991;
  assign n2993 = n32090 & ~n2991;
  assign n2994 = ~n32090 & ~n2991;
  assign n2995 = ~n2672 & n32090;
  assign n2996 = ~n32089 & n2995;
  assign n2997 = n32090 & n2991;
  assign n2998 = ~n2833 & n2996;
  assign n2999 = ~n2994 & ~n32130;
  assign n3000 = ~n2992 & ~n2993;
  assign n3001 = ~n2989 & ~n32131;
  assign n3002 = ~n2987 & ~n3001;
  assign n3003 = ~n487 & ~n3002;
  assign n3004 = ~n2688 & ~n2690;
  assign n3005 = ~n2833 & n3004;
  assign n3006 = ~n32092 & ~n3005;
  assign n3007 = ~n2690 & n32092;
  assign n3008 = ~n2688 & n3007;
  assign n3009 = n32092 & n3005;
  assign n3010 = ~n2833 & n3008;
  assign n3011 = ~n3006 & ~n32132;
  assign n3012 = n487 & ~n2987;
  assign n3013 = n487 & n3002;
  assign n3014 = ~n3001 & n3012;
  assign n3015 = ~n3011 & ~n32133;
  assign n3016 = ~n3003 & ~n3015;
  assign n3017 = ~n393 & ~n3016;
  assign n3018 = n393 & ~n3003;
  assign n3019 = ~n3015 & n3018;
  assign n3020 = ~n2705 & ~n32093;
  assign n3021 = ~n2705 & ~n2833;
  assign n3022 = ~n32093 & n3021;
  assign n3023 = ~n2833 & n3020;
  assign n3024 = n32095 & ~n32134;
  assign n3025 = n2720 & n3021;
  assign n3026 = ~n32095 & n32134;
  assign n3027 = ~n2705 & n32095;
  assign n3028 = ~n32093 & n3027;
  assign n3029 = ~n2833 & n3028;
  assign n3030 = ~n32095 & ~n32134;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = ~n3024 & ~n32135;
  assign n3033 = ~n3019 & ~n32136;
  assign n3034 = ~n3017 & ~n3033;
  assign n3035 = ~n321 & ~n3034;
  assign n3036 = ~n2722 & ~n2724;
  assign n3037 = ~n2833 & n3036;
  assign n3038 = ~n32097 & ~n3037;
  assign n3039 = ~n2724 & n32097;
  assign n3040 = ~n2722 & n3039;
  assign n3041 = n32097 & n3037;
  assign n3042 = ~n2833 & n3040;
  assign n3043 = ~n3038 & ~n32137;
  assign n3044 = n321 & ~n3017;
  assign n3045 = n321 & n3034;
  assign n3046 = ~n3033 & n3044;
  assign n3047 = ~n3043 & ~n32138;
  assign n3048 = ~n3035 & ~n3047;
  assign n3049 = ~n263 & ~n3048;
  assign n3050 = ~n2739 & ~n32098;
  assign n3051 = ~n2833 & n3050;
  assign n3052 = ~n32101 & ~n3051;
  assign n3053 = ~n2739 & n32101;
  assign n3054 = ~n32098 & n3053;
  assign n3055 = n32101 & n3051;
  assign n3056 = ~n2833 & n3054;
  assign n3057 = ~n3052 & ~n32139;
  assign n3058 = n263 & ~n3035;
  assign n3059 = ~n3047 & n3058;
  assign n3060 = ~n3057 & ~n3059;
  assign n3061 = ~n3049 & ~n3060;
  assign n3062 = ~n214 & ~n3061;
  assign n3063 = ~n2758 & ~n2760;
  assign n3064 = ~n2833 & n3063;
  assign n3065 = ~n32103 & ~n3064;
  assign n3066 = ~n2760 & n32103;
  assign n3067 = ~n2758 & n3066;
  assign n3068 = n32103 & n3064;
  assign n3069 = ~n2833 & n3067;
  assign n3070 = ~n3065 & ~n32140;
  assign n3071 = n214 & ~n3049;
  assign n3072 = n214 & n3061;
  assign n3073 = ~n3060 & n3071;
  assign n3074 = ~n3070 & ~n32141;
  assign n3075 = ~n3062 & ~n3074;
  assign n3076 = ~n197 & ~n3075;
  assign n3077 = n197 & ~n3062;
  assign n3078 = ~n3074 & n3077;
  assign n3079 = ~n2775 & ~n32105;
  assign n3080 = ~n2775 & ~n2833;
  assign n3081 = ~n32105 & n3080;
  assign n3082 = ~n2833 & n3079;
  assign n3083 = n2783 & ~n32142;
  assign n3084 = n2787 & n3080;
  assign n3085 = ~n2775 & n2783;
  assign n3086 = ~n32105 & n3085;
  assign n3087 = ~n2833 & n3086;
  assign n3088 = ~n2783 & ~n32142;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090 = ~n3083 & ~n3084;
  assign n3091 = ~n3078 & ~n32143;
  assign n3092 = ~n3076 & ~n3091;
  assign n3093 = ~n2789 & ~n2791;
  assign n3094 = ~n2833 & n3093;
  assign n3095 = ~n32107 & ~n3094;
  assign n3096 = ~n2791 & n32107;
  assign n3097 = ~n2789 & n3096;
  assign n3098 = n32107 & n3094;
  assign n3099 = ~n2833 & n3097;
  assign n3100 = ~n3095 & ~n32144;
  assign n3101 = ~n2805 & ~n32109;
  assign n3102 = ~n32109 & ~n2833;
  assign n3103 = ~n2805 & n3102;
  assign n3104 = ~n2833 & n3101;
  assign n3105 = ~n32111 & ~n32145;
  assign n3106 = ~n3100 & n3105;
  assign n3107 = ~n3092 & n3106;
  assign n3108 = n193 & ~n3107;
  assign n3109 = ~n3076 & n3100;
  assign n3110 = n3092 & n3100;
  assign n3111 = ~n3091 & n3109;
  assign n3112 = n2805 & ~n3102;
  assign n3113 = ~n193 & ~n3101;
  assign n3114 = ~n3112 & n3113;
  assign n3115 = ~n32146 & ~n3114;
  assign n3116 = ~n3108 & n3115;
  assign n3117 = pi88  & ~n3116;
  assign n3118 = ~pi86  & ~pi87 ;
  assign n3119 = ~pi88  & n3118;
  assign n3120 = ~n3117 & ~n3119;
  assign n3121 = ~n2833 & ~n3120;
  assign n3122 = ~pi88  & ~n3116;
  assign n3123 = pi89  & ~n3122;
  assign n3124 = ~pi89  & n3122;
  assign n3125 = n2835 & ~n3116;
  assign n3126 = ~n3123 & ~n32147;
  assign n3127 = ~n32069 & ~n32112;
  assign n3128 = ~n2515 & n3127;
  assign n3129 = ~n2534 & n3128;
  assign n3130 = ~n32071 & n3129;
  assign n3131 = n2520 & n2536;
  assign n3132 = ~n2528 & n3130;
  assign n3133 = ~n3119 & ~n32148;
  assign n3134 = ~n2831 & n3133;
  assign n3135 = ~n32111 & n3134;
  assign n3136 = ~n2825 & n3135;
  assign n3137 = n2833 & n3120;
  assign n3138 = ~n3117 & n3136;
  assign n3139 = n3126 & ~n32149;
  assign n3140 = ~n3121 & ~n3139;
  assign n3141 = ~n2536 & ~n3140;
  assign n3142 = n2536 & ~n3121;
  assign n3143 = ~n3139 & n3142;
  assign n3144 = ~n2833 & ~n3114;
  assign n3145 = ~n32146 & n3144;
  assign n3146 = ~n3108 & n3145;
  assign n3147 = ~n32147 & ~n3146;
  assign n3148 = pi90  & ~n3147;
  assign n3149 = ~pi90  & ~n3146;
  assign n3150 = ~pi90  & n3147;
  assign n3151 = ~n32147 & n3149;
  assign n3152 = ~n3148 & ~n32150;
  assign n3153 = ~n3143 & ~n3152;
  assign n3154 = ~n3141 & ~n3153;
  assign n3155 = ~n2283 & ~n3154;
  assign n3156 = n2283 & ~n3141;
  assign n3157 = ~n3153 & n3156;
  assign n3158 = n2283 & n3154;
  assign n3159 = ~n2838 & ~n32113;
  assign n3160 = ~n3116 & n3159;
  assign n3161 = n2855 & ~n3160;
  assign n3162 = ~n2855 & n3159;
  assign n3163 = ~n2855 & n3160;
  assign n3164 = ~n3116 & n3162;
  assign n3165 = ~n3161 & ~n32152;
  assign n3166 = ~n32151 & ~n3165;
  assign n3167 = ~n3155 & ~n3166;
  assign n3168 = ~n2021 & ~n3167;
  assign n3169 = n2021 & ~n3155;
  assign n3170 = ~n3166 & n3169;
  assign n3171 = ~n2858 & ~n32116;
  assign n3172 = ~n2858 & ~n3116;
  assign n3173 = ~n32116 & n3172;
  assign n3174 = ~n3116 & n3171;
  assign n3175 = n2867 & ~n32153;
  assign n3176 = n2871 & n3172;
  assign n3177 = n2867 & ~n32116;
  assign n3178 = ~n2858 & n3177;
  assign n3179 = ~n3116 & n3178;
  assign n3180 = ~n2867 & ~n32153;
  assign n3181 = ~n3179 & ~n3180;
  assign n3182 = ~n3175 & ~n3176;
  assign n3183 = ~n3170 & ~n32154;
  assign n3184 = ~n3168 & ~n3183;
  assign n3185 = ~n1796 & ~n3184;
  assign n3186 = n1796 & ~n3168;
  assign n3187 = ~n3183 & n3186;
  assign n3188 = n1796 & n3184;
  assign n3189 = ~n2873 & ~n2875;
  assign n3190 = ~n3116 & n3189;
  assign n3191 = ~n2882 & ~n3190;
  assign n3192 = ~n2873 & n2882;
  assign n3193 = ~n2875 & n3192;
  assign n3194 = n2882 & n3190;
  assign n3195 = ~n3116 & n3193;
  assign n3196 = n2882 & ~n3190;
  assign n3197 = ~n2882 & n3190;
  assign n3198 = ~n3196 & ~n3197;
  assign n3199 = ~n3191 & ~n32156;
  assign n3200 = ~n32155 & n32157;
  assign n3201 = ~n3185 & ~n3200;
  assign n3202 = ~n1567 & ~n3201;
  assign n3203 = n1567 & ~n3185;
  assign n3204 = ~n3200 & n3203;
  assign n3205 = ~n2885 & ~n32119;
  assign n3206 = ~n2885 & ~n3116;
  assign n3207 = ~n32119 & n3206;
  assign n3208 = ~n3116 & n3205;
  assign n3209 = n2893 & ~n32158;
  assign n3210 = n2897 & n3206;
  assign n3211 = n2893 & ~n32119;
  assign n3212 = ~n2885 & n3211;
  assign n3213 = ~n3116 & n3212;
  assign n3214 = ~n2893 & ~n32158;
  assign n3215 = ~n3213 & ~n3214;
  assign n3216 = ~n3209 & ~n3210;
  assign n3217 = ~n3204 & ~n32159;
  assign n3218 = ~n3202 & ~n3217;
  assign n3219 = ~n1374 & ~n3218;
  assign n3220 = n1374 & ~n3202;
  assign n3221 = ~n3217 & n3220;
  assign n3222 = n1374 & n3218;
  assign n3223 = ~n2899 & ~n2901;
  assign n3224 = ~n3116 & n3223;
  assign n3225 = ~n32121 & ~n3224;
  assign n3226 = n32121 & n3224;
  assign n3227 = ~n2899 & ~n32121;
  assign n3228 = ~n2901 & n3227;
  assign n3229 = ~n3116 & n3228;
  assign n3230 = n32121 & ~n3224;
  assign n3231 = ~n3229 & ~n3230;
  assign n3232 = ~n3225 & ~n3226;
  assign n3233 = ~n32160 & ~n32161;
  assign n3234 = ~n3219 & ~n3233;
  assign n3235 = ~n1179 & ~n3234;
  assign n3236 = n1179 & ~n3219;
  assign n3237 = ~n3233 & n3236;
  assign n3238 = ~n2915 & ~n32123;
  assign n3239 = ~n2915 & ~n3116;
  assign n3240 = ~n32123 & n3239;
  assign n3241 = ~n3116 & n3238;
  assign n3242 = n2923 & ~n32162;
  assign n3243 = n2927 & n3239;
  assign n3244 = n2923 & ~n32123;
  assign n3245 = ~n2915 & n3244;
  assign n3246 = ~n3116 & n3245;
  assign n3247 = ~n2923 & ~n32162;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = ~n3242 & ~n3243;
  assign n3250 = ~n3237 & ~n32163;
  assign n3251 = ~n3235 & ~n3250;
  assign n3252 = ~n1016 & ~n3251;
  assign n3253 = n1016 & ~n3235;
  assign n3254 = ~n3250 & n3253;
  assign n3255 = n1016 & n3251;
  assign n3256 = ~n2929 & ~n2931;
  assign n3257 = ~n3116 & n3256;
  assign n3258 = ~n32124 & n3257;
  assign n3259 = n32124 & ~n3257;
  assign n3260 = ~n2929 & n32124;
  assign n3261 = ~n2931 & n3260;
  assign n3262 = ~n3116 & n3261;
  assign n3263 = ~n32124 & ~n3257;
  assign n3264 = ~n3262 & ~n3263;
  assign n3265 = ~n3258 & ~n3259;
  assign n3266 = ~n32164 & ~n32165;
  assign n3267 = ~n3252 & ~n3266;
  assign n3268 = ~n855 & ~n3267;
  assign n3269 = n855 & ~n3252;
  assign n3270 = ~n3266 & n3269;
  assign n3271 = ~n2944 & ~n32126;
  assign n3272 = ~n2944 & ~n3116;
  assign n3273 = ~n32126 & n3272;
  assign n3274 = ~n3116 & n3271;
  assign n3275 = n2952 & ~n32166;
  assign n3276 = n2956 & n3272;
  assign n3277 = n2952 & ~n32126;
  assign n3278 = ~n2944 & n3277;
  assign n3279 = ~n3116 & n3278;
  assign n3280 = ~n2952 & ~n32166;
  assign n3281 = ~n3279 & ~n3280;
  assign n3282 = ~n3275 & ~n3276;
  assign n3283 = ~n3270 & ~n32167;
  assign n3284 = ~n3268 & ~n3283;
  assign n3285 = ~n720 & ~n3284;
  assign n3286 = n720 & ~n3268;
  assign n3287 = ~n3283 & n3286;
  assign n3288 = n720 & n3284;
  assign n3289 = ~n2958 & ~n2960;
  assign n3290 = ~n3116 & n3289;
  assign n3291 = ~n32127 & n3290;
  assign n3292 = n32127 & ~n3290;
  assign n3293 = ~n32127 & ~n3290;
  assign n3294 = ~n2958 & n32127;
  assign n3295 = ~n2960 & n3294;
  assign n3296 = n32127 & n3290;
  assign n3297 = ~n3116 & n3295;
  assign n3298 = ~n3293 & ~n32169;
  assign n3299 = ~n3291 & ~n3292;
  assign n3300 = ~n32168 & ~n32170;
  assign n3301 = ~n3285 & ~n3300;
  assign n3302 = ~n592 & ~n3301;
  assign n3303 = n592 & ~n3285;
  assign n3304 = ~n3300 & n3303;
  assign n3305 = ~n2973 & ~n32129;
  assign n3306 = ~n2973 & ~n3116;
  assign n3307 = ~n32129 & n3306;
  assign n3308 = ~n3116 & n3305;
  assign n3309 = n2981 & ~n32171;
  assign n3310 = n2985 & n3306;
  assign n3311 = n2981 & ~n32129;
  assign n3312 = ~n2973 & n3311;
  assign n3313 = ~n3116 & n3312;
  assign n3314 = ~n2981 & ~n32171;
  assign n3315 = ~n3313 & ~n3314;
  assign n3316 = ~n3309 & ~n3310;
  assign n3317 = ~n3304 & ~n32172;
  assign n3318 = ~n3302 & ~n3317;
  assign n3319 = ~n487 & ~n3318;
  assign n3320 = n487 & ~n3302;
  assign n3321 = ~n3317 & n3320;
  assign n3322 = n487 & n3318;
  assign n3323 = ~n2987 & ~n2989;
  assign n3324 = ~n2987 & ~n3116;
  assign n3325 = ~n2989 & n3324;
  assign n3326 = ~n3116 & n3323;
  assign n3327 = n32131 & ~n32174;
  assign n3328 = n3001 & n3324;
  assign n3329 = ~n32131 & n32174;
  assign n3330 = ~n2987 & n32131;
  assign n3331 = ~n2989 & n3330;
  assign n3332 = ~n3116 & n3331;
  assign n3333 = ~n32131 & ~n32174;
  assign n3334 = ~n3332 & ~n3333;
  assign n3335 = ~n3327 & ~n32175;
  assign n3336 = ~n32173 & ~n32176;
  assign n3337 = ~n3319 & ~n3336;
  assign n3338 = ~n393 & ~n3337;
  assign n3339 = n393 & ~n3319;
  assign n3340 = ~n3336 & n3339;
  assign n3341 = ~n3003 & ~n32133;
  assign n3342 = ~n3003 & ~n3116;
  assign n3343 = ~n32133 & n3342;
  assign n3344 = ~n3116 & n3341;
  assign n3345 = n3011 & ~n32177;
  assign n3346 = n3015 & n3342;
  assign n3347 = n3011 & ~n32133;
  assign n3348 = ~n3003 & n3347;
  assign n3349 = ~n3116 & n3348;
  assign n3350 = ~n3011 & ~n32177;
  assign n3351 = ~n3349 & ~n3350;
  assign n3352 = ~n3345 & ~n3346;
  assign n3353 = ~n3340 & ~n32178;
  assign n3354 = ~n3338 & ~n3353;
  assign n3355 = ~n321 & ~n3354;
  assign n3356 = ~n3017 & ~n3019;
  assign n3357 = ~n3116 & n3356;
  assign n3358 = ~n32136 & ~n3357;
  assign n3359 = ~n3017 & n32136;
  assign n3360 = ~n3019 & n3359;
  assign n3361 = n32136 & n3357;
  assign n3362 = ~n3116 & n3360;
  assign n3363 = ~n3358 & ~n32179;
  assign n3364 = n321 & ~n3338;
  assign n3365 = ~n3353 & n3364;
  assign n3366 = n321 & n3354;
  assign n3367 = ~n3363 & ~n32180;
  assign n3368 = ~n3355 & ~n3367;
  assign n3369 = ~n263 & ~n3368;
  assign n3370 = n263 & ~n3355;
  assign n3371 = ~n3367 & n3370;
  assign n3372 = ~n3035 & ~n32138;
  assign n3373 = ~n3035 & ~n3116;
  assign n3374 = ~n32138 & n3373;
  assign n3375 = ~n3116 & n3372;
  assign n3376 = n3043 & ~n32181;
  assign n3377 = n3047 & n3373;
  assign n3378 = n3043 & ~n32138;
  assign n3379 = ~n3035 & n3378;
  assign n3380 = ~n3116 & n3379;
  assign n3381 = ~n3043 & ~n32181;
  assign n3382 = ~n3380 & ~n3381;
  assign n3383 = ~n3376 & ~n3377;
  assign n3384 = ~n3371 & ~n32182;
  assign n3385 = ~n3369 & ~n3384;
  assign n3386 = ~n214 & ~n3385;
  assign n3387 = n214 & ~n3369;
  assign n3388 = ~n3384 & n3387;
  assign n3389 = n214 & n3385;
  assign n3390 = ~n3049 & ~n3059;
  assign n3391 = ~n3049 & ~n3116;
  assign n3392 = ~n3059 & n3391;
  assign n3393 = ~n3116 & n3390;
  assign n3394 = n3057 & ~n32184;
  assign n3395 = n3060 & n3391;
  assign n3396 = ~n3049 & n3057;
  assign n3397 = ~n3059 & n3396;
  assign n3398 = ~n3116 & n3397;
  assign n3399 = ~n3057 & ~n32184;
  assign n3400 = ~n3398 & ~n3399;
  assign n3401 = ~n3394 & ~n3395;
  assign n3402 = ~n32183 & ~n32185;
  assign n3403 = ~n3386 & ~n3402;
  assign n3404 = ~n197 & ~n3403;
  assign n3405 = n197 & ~n3386;
  assign n3406 = ~n3402 & n3405;
  assign n3407 = ~n3062 & ~n32141;
  assign n3408 = ~n3062 & ~n3116;
  assign n3409 = ~n32141 & n3408;
  assign n3410 = ~n3116 & n3407;
  assign n3411 = n3070 & ~n32186;
  assign n3412 = n3074 & n3408;
  assign n3413 = n3070 & ~n32141;
  assign n3414 = ~n3062 & n3413;
  assign n3415 = ~n3116 & n3414;
  assign n3416 = ~n3070 & ~n32186;
  assign n3417 = ~n3415 & ~n3416;
  assign n3418 = ~n3411 & ~n3412;
  assign n3419 = ~n3406 & ~n32187;
  assign n3420 = ~n3404 & ~n3419;
  assign n3421 = ~n3076 & ~n3078;
  assign n3422 = ~n3116 & n3421;
  assign n3423 = ~n32143 & ~n3422;
  assign n3424 = ~n3076 & n32143;
  assign n3425 = ~n3078 & n3424;
  assign n3426 = n32143 & n3422;
  assign n3427 = ~n3116 & n3425;
  assign n3428 = ~n3423 & ~n32188;
  assign n3429 = ~n3092 & ~n3100;
  assign n3430 = ~n3100 & ~n3116;
  assign n3431 = ~n3092 & n3430;
  assign n3432 = ~n3116 & n3429;
  assign n3433 = ~n32146 & ~n32189;
  assign n3434 = ~n3428 & n3433;
  assign n3435 = ~n3420 & n3434;
  assign n3436 = n193 & ~n3435;
  assign n3437 = ~n3404 & n3428;
  assign n3438 = ~n3419 & n3437;
  assign n3439 = n3420 & n3428;
  assign n3440 = n3092 & ~n3430;
  assign n3441 = ~n193 & ~n3429;
  assign n3442 = ~n3440 & n3441;
  assign n3443 = ~n32190 & ~n3442;
  assign n3444 = ~n3436 & n3443;
  assign n3445 = pi86  & ~n3444;
  assign n3446 = ~pi84  & ~pi85 ;
  assign n3447 = ~pi86  & n3446;
  assign n3448 = ~n3445 & ~n3447;
  assign n3449 = ~n3116 & ~n3448;
  assign n3450 = ~n2814 & ~n32148;
  assign n3451 = ~n2815 & n3450;
  assign n3452 = ~n2831 & n3451;
  assign n3453 = ~n32111 & n3452;
  assign n3454 = n32109 & n2833;
  assign n3455 = ~n2825 & n3453;
  assign n3456 = ~n3447 & ~n32191;
  assign n3457 = ~n3114 & n3456;
  assign n3458 = ~n32146 & n3457;
  assign n3459 = ~n3108 & n3458;
  assign n3460 = n3116 & n3448;
  assign n3461 = ~n3445 & n3459;
  assign n3462 = ~pi86  & ~n3444;
  assign n3463 = pi87  & ~n3462;
  assign n3464 = ~pi87  & n3462;
  assign n3465 = n3118 & ~n3444;
  assign n3466 = ~n3463 & ~n32193;
  assign n3467 = ~n32192 & n3466;
  assign n3468 = ~n3449 & ~n3467;
  assign n3469 = ~n2833 & ~n3468;
  assign n3470 = ~n3116 & ~n3442;
  assign n3471 = ~n32190 & n3470;
  assign n3472 = ~n3436 & n3471;
  assign n3473 = ~n32193 & ~n3472;
  assign n3474 = pi88  & ~n3473;
  assign n3475 = ~pi88  & ~n3472;
  assign n3476 = ~pi88  & n3473;
  assign n3477 = ~n32193 & n3475;
  assign n3478 = ~n3474 & ~n32194;
  assign n3479 = n2833 & ~n3449;
  assign n3480 = n2833 & n3468;
  assign n3481 = ~n3467 & n3479;
  assign n3482 = ~n3478 & ~n32195;
  assign n3483 = ~n3469 & ~n3482;
  assign n3484 = ~n2536 & ~n3483;
  assign n3485 = n2536 & ~n3469;
  assign n3486 = ~n3482 & n3485;
  assign n3487 = ~n3121 & ~n32149;
  assign n3488 = ~n3444 & n3487;
  assign n3489 = n3126 & ~n3488;
  assign n3490 = ~n3126 & n3487;
  assign n3491 = ~n3126 & n3488;
  assign n3492 = ~n3444 & n3490;
  assign n3493 = ~n3489 & ~n32196;
  assign n3494 = ~n3486 & ~n3493;
  assign n3495 = ~n3484 & ~n3494;
  assign n3496 = ~n2283 & ~n3495;
  assign n3497 = ~n3141 & ~n3143;
  assign n3498 = ~n3444 & n3497;
  assign n3499 = ~n3152 & ~n3498;
  assign n3500 = ~n3143 & n3152;
  assign n3501 = ~n3141 & n3500;
  assign n3502 = n3152 & n3498;
  assign n3503 = ~n3444 & n3501;
  assign n3504 = ~n3499 & ~n32197;
  assign n3505 = n2283 & ~n3484;
  assign n3506 = n2283 & n3495;
  assign n3507 = ~n3494 & n3505;
  assign n3508 = ~n3504 & ~n32198;
  assign n3509 = ~n3496 & ~n3508;
  assign n3510 = ~n2021 & ~n3509;
  assign n3511 = n2021 & ~n3496;
  assign n3512 = ~n3508 & n3511;
  assign n3513 = ~n3155 & ~n32151;
  assign n3514 = ~n3444 & n3513;
  assign n3515 = ~n3165 & ~n3514;
  assign n3516 = ~n3155 & n3165;
  assign n3517 = ~n32151 & n3516;
  assign n3518 = n3165 & n3514;
  assign n3519 = ~n3444 & n3517;
  assign n3520 = n3165 & ~n3514;
  assign n3521 = ~n3165 & n3514;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = ~n3515 & ~n32199;
  assign n3524 = ~n3512 & n32200;
  assign n3525 = ~n3510 & ~n3524;
  assign n3526 = ~n1796 & ~n3525;
  assign n3527 = ~n3168 & ~n3170;
  assign n3528 = ~n3444 & n3527;
  assign n3529 = ~n32154 & ~n3528;
  assign n3530 = ~n3170 & n32154;
  assign n3531 = ~n3168 & n3530;
  assign n3532 = n32154 & n3528;
  assign n3533 = ~n3444 & n3531;
  assign n3534 = ~n3529 & ~n32201;
  assign n3535 = n1796 & ~n3510;
  assign n3536 = n1796 & n3525;
  assign n3537 = ~n3524 & n3535;
  assign n3538 = ~n3534 & ~n32202;
  assign n3539 = ~n3526 & ~n3538;
  assign n3540 = ~n1567 & ~n3539;
  assign n3541 = n1567 & ~n3526;
  assign n3542 = ~n3538 & n3541;
  assign n3543 = ~n3185 & ~n32155;
  assign n3544 = ~n3444 & n3543;
  assign n3545 = ~n32157 & ~n3544;
  assign n3546 = n32157 & n3544;
  assign n3547 = ~n3185 & ~n32157;
  assign n3548 = ~n32155 & n3547;
  assign n3549 = ~n3444 & n3548;
  assign n3550 = n32157 & ~n3544;
  assign n3551 = ~n3549 & ~n3550;
  assign n3552 = ~n3545 & ~n3546;
  assign n3553 = ~n3542 & ~n32203;
  assign n3554 = ~n3540 & ~n3553;
  assign n3555 = ~n1374 & ~n3554;
  assign n3556 = ~n3202 & ~n3204;
  assign n3557 = ~n3444 & n3556;
  assign n3558 = ~n32159 & ~n3557;
  assign n3559 = ~n3204 & n32159;
  assign n3560 = ~n3202 & n3559;
  assign n3561 = n32159 & n3557;
  assign n3562 = ~n3444 & n3560;
  assign n3563 = ~n3558 & ~n32204;
  assign n3564 = n1374 & ~n3540;
  assign n3565 = n1374 & n3554;
  assign n3566 = ~n3553 & n3564;
  assign n3567 = ~n3563 & ~n32205;
  assign n3568 = ~n3555 & ~n3567;
  assign n3569 = ~n1179 & ~n3568;
  assign n3570 = n1179 & ~n3555;
  assign n3571 = ~n3567 & n3570;
  assign n3572 = ~n3219 & ~n32160;
  assign n3573 = ~n3444 & n3572;
  assign n3574 = ~n32161 & n3573;
  assign n3575 = n32161 & ~n3573;
  assign n3576 = ~n3219 & n32161;
  assign n3577 = ~n32160 & n3576;
  assign n3578 = ~n3444 & n3577;
  assign n3579 = ~n32161 & ~n3573;
  assign n3580 = ~n3578 & ~n3579;
  assign n3581 = ~n3574 & ~n3575;
  assign n3582 = ~n3571 & ~n32206;
  assign n3583 = ~n3569 & ~n3582;
  assign n3584 = ~n1016 & ~n3583;
  assign n3585 = ~n3235 & ~n3237;
  assign n3586 = ~n3444 & n3585;
  assign n3587 = ~n32163 & ~n3586;
  assign n3588 = ~n3237 & n32163;
  assign n3589 = ~n3235 & n3588;
  assign n3590 = n32163 & n3586;
  assign n3591 = ~n3444 & n3589;
  assign n3592 = ~n3587 & ~n32207;
  assign n3593 = n1016 & ~n3569;
  assign n3594 = n1016 & n3583;
  assign n3595 = ~n3582 & n3593;
  assign n3596 = ~n3592 & ~n32208;
  assign n3597 = ~n3584 & ~n3596;
  assign n3598 = ~n855 & ~n3597;
  assign n3599 = n855 & ~n3584;
  assign n3600 = ~n3596 & n3599;
  assign n3601 = ~n3252 & ~n32164;
  assign n3602 = ~n3444 & n3601;
  assign n3603 = ~n32165 & ~n3602;
  assign n3604 = ~n3252 & n32165;
  assign n3605 = ~n32164 & n3604;
  assign n3606 = n32165 & n3602;
  assign n3607 = ~n3444 & n3605;
  assign n3608 = n32165 & ~n3602;
  assign n3609 = ~n32165 & n3602;
  assign n3610 = ~n3608 & ~n3609;
  assign n3611 = ~n3603 & ~n32209;
  assign n3612 = ~n3600 & n32210;
  assign n3613 = ~n3598 & ~n3612;
  assign n3614 = ~n720 & ~n3613;
  assign n3615 = ~n3268 & ~n3270;
  assign n3616 = ~n3444 & n3615;
  assign n3617 = ~n32167 & ~n3616;
  assign n3618 = ~n3270 & n32167;
  assign n3619 = ~n3268 & n3618;
  assign n3620 = n32167 & n3616;
  assign n3621 = ~n3444 & n3619;
  assign n3622 = ~n3617 & ~n32211;
  assign n3623 = n720 & ~n3598;
  assign n3624 = n720 & n3613;
  assign n3625 = ~n3612 & n3623;
  assign n3626 = ~n3622 & ~n32212;
  assign n3627 = ~n3614 & ~n3626;
  assign n3628 = ~n592 & ~n3627;
  assign n3629 = n592 & ~n3614;
  assign n3630 = ~n3626 & n3629;
  assign n3631 = ~n3285 & ~n32168;
  assign n3632 = ~n3285 & ~n3444;
  assign n3633 = ~n32168 & n3632;
  assign n3634 = ~n3444 & n3631;
  assign n3635 = n32170 & ~n32213;
  assign n3636 = n3300 & n3632;
  assign n3637 = ~n32170 & n32213;
  assign n3638 = ~n3285 & n32170;
  assign n3639 = ~n32168 & n3638;
  assign n3640 = ~n3444 & n3639;
  assign n3641 = ~n32170 & ~n32213;
  assign n3642 = ~n3640 & ~n3641;
  assign n3643 = ~n3635 & ~n32214;
  assign n3644 = ~n3630 & ~n32215;
  assign n3645 = ~n3628 & ~n3644;
  assign n3646 = ~n487 & ~n3645;
  assign n3647 = ~n3302 & ~n3304;
  assign n3648 = ~n3444 & n3647;
  assign n3649 = ~n32172 & ~n3648;
  assign n3650 = ~n3304 & n32172;
  assign n3651 = ~n3302 & n3650;
  assign n3652 = n32172 & n3648;
  assign n3653 = ~n3444 & n3651;
  assign n3654 = ~n3649 & ~n32216;
  assign n3655 = n487 & ~n3628;
  assign n3656 = n487 & n3645;
  assign n3657 = ~n3644 & n3655;
  assign n3658 = ~n3654 & ~n32217;
  assign n3659 = ~n3646 & ~n3658;
  assign n3660 = ~n393 & ~n3659;
  assign n3661 = ~n3319 & ~n32173;
  assign n3662 = ~n3444 & n3661;
  assign n3663 = ~n32176 & ~n3662;
  assign n3664 = ~n3319 & n32176;
  assign n3665 = ~n32173 & n3664;
  assign n3666 = n32176 & n3662;
  assign n3667 = ~n3444 & n3665;
  assign n3668 = ~n3663 & ~n32218;
  assign n3669 = n393 & ~n3646;
  assign n3670 = ~n3658 & n3669;
  assign n3671 = ~n3668 & ~n3670;
  assign n3672 = ~n3660 & ~n3671;
  assign n3673 = ~n321 & ~n3672;
  assign n3674 = ~n3338 & ~n3340;
  assign n3675 = ~n3444 & n3674;
  assign n3676 = ~n32178 & ~n3675;
  assign n3677 = ~n3340 & n32178;
  assign n3678 = ~n3338 & n3677;
  assign n3679 = n32178 & n3675;
  assign n3680 = ~n3444 & n3678;
  assign n3681 = ~n3676 & ~n32219;
  assign n3682 = n321 & ~n3660;
  assign n3683 = n321 & n3672;
  assign n3684 = ~n3671 & n3682;
  assign n3685 = ~n3681 & ~n32220;
  assign n3686 = ~n3673 & ~n3685;
  assign n3687 = ~n263 & ~n3686;
  assign n3688 = n263 & ~n3673;
  assign n3689 = ~n3685 & n3688;
  assign n3690 = ~n3355 & ~n32180;
  assign n3691 = ~n3355 & ~n3444;
  assign n3692 = ~n32180 & n3691;
  assign n3693 = ~n3444 & n3690;
  assign n3694 = n3363 & ~n32221;
  assign n3695 = n3367 & n3691;
  assign n3696 = ~n3355 & n3363;
  assign n3697 = ~n32180 & n3696;
  assign n3698 = ~n3444 & n3697;
  assign n3699 = ~n3363 & ~n32221;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = ~n3694 & ~n3695;
  assign n3702 = ~n3689 & ~n32222;
  assign n3703 = ~n3687 & ~n3702;
  assign n3704 = ~n214 & ~n3703;
  assign n3705 = ~n3369 & ~n3371;
  assign n3706 = ~n3444 & n3705;
  assign n3707 = ~n32182 & ~n3706;
  assign n3708 = ~n3371 & n32182;
  assign n3709 = ~n3369 & n3708;
  assign n3710 = n32182 & n3706;
  assign n3711 = ~n3444 & n3709;
  assign n3712 = ~n3707 & ~n32223;
  assign n3713 = n214 & ~n3687;
  assign n3714 = n214 & n3703;
  assign n3715 = ~n3702 & n3713;
  assign n3716 = ~n3712 & ~n32224;
  assign n3717 = ~n3704 & ~n3716;
  assign n3718 = ~n197 & ~n3717;
  assign n3719 = ~n3386 & ~n32183;
  assign n3720 = ~n3444 & n3719;
  assign n3721 = ~n32185 & ~n3720;
  assign n3722 = ~n3386 & n32185;
  assign n3723 = ~n32183 & n3722;
  assign n3724 = n32185 & n3720;
  assign n3725 = ~n3444 & n3723;
  assign n3726 = ~n3721 & ~n32225;
  assign n3727 = n197 & ~n3704;
  assign n3728 = ~n3716 & n3727;
  assign n3729 = ~n3726 & ~n3728;
  assign n3730 = ~n3718 & ~n3729;
  assign n3731 = ~n3404 & ~n3406;
  assign n3732 = ~n3444 & n3731;
  assign n3733 = ~n32187 & ~n3732;
  assign n3734 = ~n3406 & n32187;
  assign n3735 = ~n3404 & n3734;
  assign n3736 = n32187 & n3732;
  assign n3737 = ~n3444 & n3735;
  assign n3738 = ~n3733 & ~n32226;
  assign n3739 = ~n3420 & ~n3428;
  assign n3740 = ~n3428 & ~n3444;
  assign n3741 = ~n3420 & n3740;
  assign n3742 = ~n3444 & n3739;
  assign n3743 = ~n32190 & ~n32227;
  assign n3744 = ~n3738 & n3743;
  assign n3745 = ~n3730 & n3744;
  assign n3746 = n193 & ~n3745;
  assign n3747 = ~n3718 & n3738;
  assign n3748 = n3730 & n3738;
  assign n3749 = ~n3729 & n3747;
  assign n3750 = n3420 & ~n3740;
  assign n3751 = ~n193 & ~n3739;
  assign n3752 = ~n3750 & n3751;
  assign n3753 = ~n32228 & ~n3752;
  assign n3754 = ~n3746 & n3753;
  assign n3755 = pi84  & ~n3754;
  assign n3756 = ~pi82  & ~pi83 ;
  assign n3757 = ~pi84  & n3756;
  assign n3758 = ~n3755 & ~n3757;
  assign n3759 = ~n3444 & ~n3758;
  assign n3760 = ~pi84  & ~n3754;
  assign n3761 = pi85  & ~n3760;
  assign n3762 = ~pi85  & n3760;
  assign n3763 = n3446 & ~n3754;
  assign n3764 = ~n3761 & ~n32229;
  assign n3765 = ~n32144 & ~n32191;
  assign n3766 = ~n3095 & n3765;
  assign n3767 = ~n3114 & n3766;
  assign n3768 = ~n32146 & n3767;
  assign n3769 = n3100 & n3116;
  assign n3770 = ~n3108 & n3768;
  assign n3771 = ~n3757 & ~n32230;
  assign n3772 = ~n3442 & n3771;
  assign n3773 = ~n32190 & n3772;
  assign n3774 = ~n3436 & n3773;
  assign n3775 = n3444 & n3758;
  assign n3776 = ~n3755 & n3774;
  assign n3777 = n3764 & ~n32231;
  assign n3778 = ~n3759 & ~n3777;
  assign n3779 = ~n3116 & ~n3778;
  assign n3780 = n3116 & ~n3759;
  assign n3781 = ~n3777 & n3780;
  assign n3782 = ~n3444 & ~n3752;
  assign n3783 = ~n32228 & n3782;
  assign n3784 = ~n3746 & n3783;
  assign n3785 = ~n32229 & ~n3784;
  assign n3786 = pi86  & ~n3785;
  assign n3787 = ~pi86  & ~n3784;
  assign n3788 = ~pi86  & n3785;
  assign n3789 = ~n32229 & n3787;
  assign n3790 = ~n3786 & ~n32232;
  assign n3791 = ~n3781 & ~n3790;
  assign n3792 = ~n3779 & ~n3791;
  assign n3793 = ~n2833 & ~n3792;
  assign n3794 = n2833 & ~n3779;
  assign n3795 = ~n3791 & n3794;
  assign n3796 = n2833 & n3792;
  assign n3797 = ~n3449 & ~n32192;
  assign n3798 = ~n3754 & n3797;
  assign n3799 = n3466 & ~n3798;
  assign n3800 = ~n3466 & n3797;
  assign n3801 = ~n3466 & n3798;
  assign n3802 = ~n3754 & n3800;
  assign n3803 = ~n3799 & ~n32234;
  assign n3804 = ~n32233 & ~n3803;
  assign n3805 = ~n3793 & ~n3804;
  assign n3806 = ~n2536 & ~n3805;
  assign n3807 = n2536 & ~n3793;
  assign n3808 = ~n3804 & n3807;
  assign n3809 = ~n3469 & ~n32195;
  assign n3810 = ~n3469 & ~n3754;
  assign n3811 = ~n32195 & n3810;
  assign n3812 = ~n3754 & n3809;
  assign n3813 = n3478 & ~n32235;
  assign n3814 = n3482 & n3810;
  assign n3815 = n3478 & ~n32195;
  assign n3816 = ~n3469 & n3815;
  assign n3817 = ~n3754 & n3816;
  assign n3818 = ~n3478 & ~n32235;
  assign n3819 = ~n3817 & ~n3818;
  assign n3820 = ~n3813 & ~n3814;
  assign n3821 = ~n3808 & ~n32236;
  assign n3822 = ~n3806 & ~n3821;
  assign n3823 = ~n2283 & ~n3822;
  assign n3824 = n2283 & ~n3806;
  assign n3825 = ~n3821 & n3824;
  assign n3826 = n2283 & n3822;
  assign n3827 = ~n3484 & ~n3486;
  assign n3828 = ~n3754 & n3827;
  assign n3829 = ~n3493 & ~n3828;
  assign n3830 = ~n3484 & n3493;
  assign n3831 = ~n3486 & n3830;
  assign n3832 = n3493 & n3828;
  assign n3833 = ~n3754 & n3831;
  assign n3834 = n3493 & ~n3828;
  assign n3835 = ~n3493 & n3828;
  assign n3836 = ~n3834 & ~n3835;
  assign n3837 = ~n3829 & ~n32238;
  assign n3838 = ~n32237 & n32239;
  assign n3839 = ~n3823 & ~n3838;
  assign n3840 = ~n2021 & ~n3839;
  assign n3841 = n2021 & ~n3823;
  assign n3842 = ~n3838 & n3841;
  assign n3843 = ~n3496 & ~n32198;
  assign n3844 = ~n3496 & ~n3754;
  assign n3845 = ~n32198 & n3844;
  assign n3846 = ~n3754 & n3843;
  assign n3847 = n3504 & ~n32240;
  assign n3848 = n3508 & n3844;
  assign n3849 = n3504 & ~n32198;
  assign n3850 = ~n3496 & n3849;
  assign n3851 = ~n3754 & n3850;
  assign n3852 = ~n3504 & ~n32240;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = ~n3847 & ~n3848;
  assign n3855 = ~n3842 & ~n32241;
  assign n3856 = ~n3840 & ~n3855;
  assign n3857 = ~n1796 & ~n3856;
  assign n3858 = n1796 & ~n3840;
  assign n3859 = ~n3855 & n3858;
  assign n3860 = n1796 & n3856;
  assign n3861 = ~n3510 & ~n3512;
  assign n3862 = ~n3754 & n3861;
  assign n3863 = ~n32200 & ~n3862;
  assign n3864 = n32200 & n3862;
  assign n3865 = ~n3510 & ~n32200;
  assign n3866 = ~n3512 & n3865;
  assign n3867 = ~n3754 & n3866;
  assign n3868 = n32200 & ~n3862;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = ~n3863 & ~n3864;
  assign n3871 = ~n32242 & ~n32243;
  assign n3872 = ~n3857 & ~n3871;
  assign n3873 = ~n1567 & ~n3872;
  assign n3874 = n1567 & ~n3857;
  assign n3875 = ~n3871 & n3874;
  assign n3876 = ~n3526 & ~n32202;
  assign n3877 = ~n3526 & ~n3754;
  assign n3878 = ~n32202 & n3877;
  assign n3879 = ~n3754 & n3876;
  assign n3880 = n3534 & ~n32244;
  assign n3881 = n3538 & n3877;
  assign n3882 = n3534 & ~n32202;
  assign n3883 = ~n3526 & n3882;
  assign n3884 = ~n3754 & n3883;
  assign n3885 = ~n3534 & ~n32244;
  assign n3886 = ~n3884 & ~n3885;
  assign n3887 = ~n3880 & ~n3881;
  assign n3888 = ~n3875 & ~n32245;
  assign n3889 = ~n3873 & ~n3888;
  assign n3890 = ~n1374 & ~n3889;
  assign n3891 = n1374 & ~n3873;
  assign n3892 = ~n3888 & n3891;
  assign n3893 = n1374 & n3889;
  assign n3894 = ~n3540 & ~n3542;
  assign n3895 = ~n3754 & n3894;
  assign n3896 = ~n32203 & n3895;
  assign n3897 = n32203 & ~n3895;
  assign n3898 = ~n3540 & n32203;
  assign n3899 = ~n3542 & n3898;
  assign n3900 = ~n3754 & n3899;
  assign n3901 = ~n32203 & ~n3895;
  assign n3902 = ~n3900 & ~n3901;
  assign n3903 = ~n3896 & ~n3897;
  assign n3904 = ~n32246 & ~n32247;
  assign n3905 = ~n3890 & ~n3904;
  assign n3906 = ~n1179 & ~n3905;
  assign n3907 = n1179 & ~n3890;
  assign n3908 = ~n3904 & n3907;
  assign n3909 = ~n3555 & ~n32205;
  assign n3910 = ~n3555 & ~n3754;
  assign n3911 = ~n32205 & n3910;
  assign n3912 = ~n3754 & n3909;
  assign n3913 = n3563 & ~n32248;
  assign n3914 = n3567 & n3910;
  assign n3915 = n3563 & ~n32205;
  assign n3916 = ~n3555 & n3915;
  assign n3917 = ~n3754 & n3916;
  assign n3918 = ~n3563 & ~n32248;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~n3913 & ~n3914;
  assign n3921 = ~n3908 & ~n32249;
  assign n3922 = ~n3906 & ~n3921;
  assign n3923 = ~n1016 & ~n3922;
  assign n3924 = n1016 & ~n3906;
  assign n3925 = ~n3921 & n3924;
  assign n3926 = n1016 & n3922;
  assign n3927 = ~n3569 & ~n3571;
  assign n3928 = ~n3754 & n3927;
  assign n3929 = ~n32206 & n3928;
  assign n3930 = n32206 & ~n3928;
  assign n3931 = ~n32206 & ~n3928;
  assign n3932 = ~n3569 & n32206;
  assign n3933 = ~n3571 & n3932;
  assign n3934 = n32206 & n3928;
  assign n3935 = ~n3754 & n3933;
  assign n3936 = ~n3931 & ~n32251;
  assign n3937 = ~n3929 & ~n3930;
  assign n3938 = ~n32250 & ~n32252;
  assign n3939 = ~n3923 & ~n3938;
  assign n3940 = ~n855 & ~n3939;
  assign n3941 = n855 & ~n3923;
  assign n3942 = ~n3938 & n3941;
  assign n3943 = ~n3584 & ~n32208;
  assign n3944 = ~n3584 & ~n3754;
  assign n3945 = ~n32208 & n3944;
  assign n3946 = ~n3754 & n3943;
  assign n3947 = n3592 & ~n32253;
  assign n3948 = n3596 & n3944;
  assign n3949 = n3592 & ~n32208;
  assign n3950 = ~n3584 & n3949;
  assign n3951 = ~n3754 & n3950;
  assign n3952 = ~n3592 & ~n32253;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = ~n3947 & ~n3948;
  assign n3955 = ~n3942 & ~n32254;
  assign n3956 = ~n3940 & ~n3955;
  assign n3957 = ~n720 & ~n3956;
  assign n3958 = n720 & ~n3940;
  assign n3959 = ~n3955 & n3958;
  assign n3960 = n720 & n3956;
  assign n3961 = ~n3598 & ~n3600;
  assign n3962 = ~n3754 & n3961;
  assign n3963 = ~n32210 & ~n3962;
  assign n3964 = n32210 & n3962;
  assign n3965 = n32210 & ~n3962;
  assign n3966 = ~n3598 & ~n32210;
  assign n3967 = ~n3600 & n3966;
  assign n3968 = ~n32210 & n3962;
  assign n3969 = ~n3754 & n3967;
  assign n3970 = ~n3965 & ~n32256;
  assign n3971 = ~n3963 & ~n3964;
  assign n3972 = ~n32255 & ~n32257;
  assign n3973 = ~n3957 & ~n3972;
  assign n3974 = ~n592 & ~n3973;
  assign n3975 = n592 & ~n3957;
  assign n3976 = ~n3972 & n3975;
  assign n3977 = ~n3614 & ~n32212;
  assign n3978 = ~n3614 & ~n3754;
  assign n3979 = ~n32212 & n3978;
  assign n3980 = ~n3754 & n3977;
  assign n3981 = n3622 & ~n32258;
  assign n3982 = n3626 & n3978;
  assign n3983 = n3622 & ~n32212;
  assign n3984 = ~n3614 & n3983;
  assign n3985 = ~n3754 & n3984;
  assign n3986 = ~n3622 & ~n32258;
  assign n3987 = ~n3985 & ~n3986;
  assign n3988 = ~n3981 & ~n3982;
  assign n3989 = ~n3976 & ~n32259;
  assign n3990 = ~n3974 & ~n3989;
  assign n3991 = ~n487 & ~n3990;
  assign n3992 = ~n3628 & ~n3630;
  assign n3993 = ~n3754 & n3992;
  assign n3994 = ~n32215 & ~n3993;
  assign n3995 = ~n3628 & n32215;
  assign n3996 = ~n3630 & n3995;
  assign n3997 = n32215 & n3993;
  assign n3998 = ~n3754 & n3996;
  assign n3999 = ~n3994 & ~n32260;
  assign n4000 = n487 & ~n3974;
  assign n4001 = ~n3989 & n4000;
  assign n4002 = n487 & n3990;
  assign n4003 = ~n3999 & ~n32261;
  assign n4004 = ~n3991 & ~n4003;
  assign n4005 = ~n393 & ~n4004;
  assign n4006 = n393 & ~n3991;
  assign n4007 = ~n4003 & n4006;
  assign n4008 = ~n3646 & ~n32217;
  assign n4009 = ~n3646 & ~n3754;
  assign n4010 = ~n32217 & n4009;
  assign n4011 = ~n3754 & n4008;
  assign n4012 = n3654 & ~n32262;
  assign n4013 = n3658 & n4009;
  assign n4014 = n3654 & ~n32217;
  assign n4015 = ~n3646 & n4014;
  assign n4016 = ~n3754 & n4015;
  assign n4017 = ~n3654 & ~n32262;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = ~n4012 & ~n4013;
  assign n4020 = ~n4007 & ~n32263;
  assign n4021 = ~n4005 & ~n4020;
  assign n4022 = ~n321 & ~n4021;
  assign n4023 = n321 & ~n4005;
  assign n4024 = ~n4020 & n4023;
  assign n4025 = n321 & n4021;
  assign n4026 = ~n3660 & ~n3670;
  assign n4027 = ~n3660 & ~n3754;
  assign n4028 = ~n3670 & n4027;
  assign n4029 = ~n3754 & n4026;
  assign n4030 = n3668 & ~n32265;
  assign n4031 = n3671 & n4027;
  assign n4032 = ~n3660 & n3668;
  assign n4033 = ~n3670 & n4032;
  assign n4034 = ~n3754 & n4033;
  assign n4035 = ~n3668 & ~n32265;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = ~n4030 & ~n4031;
  assign n4038 = ~n32264 & ~n32266;
  assign n4039 = ~n4022 & ~n4038;
  assign n4040 = ~n263 & ~n4039;
  assign n4041 = n263 & ~n4022;
  assign n4042 = ~n4038 & n4041;
  assign n4043 = ~n3673 & ~n32220;
  assign n4044 = ~n3673 & ~n3754;
  assign n4045 = ~n32220 & n4044;
  assign n4046 = ~n3754 & n4043;
  assign n4047 = n3681 & ~n32267;
  assign n4048 = n3685 & n4044;
  assign n4049 = n3681 & ~n32220;
  assign n4050 = ~n3673 & n4049;
  assign n4051 = ~n3754 & n4050;
  assign n4052 = ~n3681 & ~n32267;
  assign n4053 = ~n4051 & ~n4052;
  assign n4054 = ~n4047 & ~n4048;
  assign n4055 = ~n4042 & ~n32268;
  assign n4056 = ~n4040 & ~n4055;
  assign n4057 = ~n214 & ~n4056;
  assign n4058 = ~n3687 & ~n3689;
  assign n4059 = ~n3754 & n4058;
  assign n4060 = ~n32222 & ~n4059;
  assign n4061 = ~n3687 & n32222;
  assign n4062 = ~n3689 & n4061;
  assign n4063 = n32222 & n4059;
  assign n4064 = ~n3754 & n4062;
  assign n4065 = ~n4060 & ~n32269;
  assign n4066 = n214 & ~n4040;
  assign n4067 = ~n4055 & n4066;
  assign n4068 = n214 & n4056;
  assign n4069 = ~n4065 & ~n32270;
  assign n4070 = ~n4057 & ~n4069;
  assign n4071 = ~n197 & ~n4070;
  assign n4072 = n197 & ~n4057;
  assign n4073 = ~n4069 & n4072;
  assign n4074 = ~n3704 & ~n32224;
  assign n4075 = ~n3704 & ~n3754;
  assign n4076 = ~n32224 & n4075;
  assign n4077 = ~n3754 & n4074;
  assign n4078 = n3712 & ~n32271;
  assign n4079 = n3716 & n4075;
  assign n4080 = n3712 & ~n32224;
  assign n4081 = ~n3704 & n4080;
  assign n4082 = ~n3754 & n4081;
  assign n4083 = ~n3712 & ~n32271;
  assign n4084 = ~n4082 & ~n4083;
  assign n4085 = ~n4078 & ~n4079;
  assign n4086 = ~n4073 & ~n32272;
  assign n4087 = ~n4071 & ~n4086;
  assign n4088 = ~n3718 & ~n3728;
  assign n4089 = ~n3718 & ~n3754;
  assign n4090 = ~n3728 & n4089;
  assign n4091 = ~n3754 & n4088;
  assign n4092 = n3726 & ~n32273;
  assign n4093 = n3729 & n4089;
  assign n4094 = ~n3718 & n3726;
  assign n4095 = ~n3728 & n4094;
  assign n4096 = ~n3754 & n4095;
  assign n4097 = ~n3726 & ~n32273;
  assign n4098 = ~n4096 & ~n4097;
  assign n4099 = ~n4092 & ~n4093;
  assign n4100 = ~n3730 & ~n3738;
  assign n4101 = ~n3738 & ~n3754;
  assign n4102 = ~n3730 & n4101;
  assign n4103 = ~n3754 & n4100;
  assign n4104 = ~n32228 & ~n32275;
  assign n4105 = ~n32274 & n4104;
  assign n4106 = ~n4087 & n4105;
  assign n4107 = n193 & ~n4106;
  assign n4108 = ~n4071 & n32274;
  assign n4109 = ~n4086 & n4108;
  assign n4110 = n4087 & n32274;
  assign n4111 = n3730 & ~n4101;
  assign n4112 = ~n193 & ~n4100;
  assign n4113 = ~n4111 & n4112;
  assign n4114 = ~n32276 & ~n4113;
  assign n4115 = ~n4107 & n4114;
  assign n4116 = pi82  & ~n4115;
  assign n4117 = ~pi80  & ~pi81 ;
  assign n4118 = ~pi82  & n4117;
  assign n4119 = ~n4116 & ~n4118;
  assign n4120 = ~n3754 & ~n4119;
  assign n4121 = ~n32188 & ~n32230;
  assign n4122 = ~n3423 & n4121;
  assign n4123 = ~n3442 & n4122;
  assign n4124 = ~n32190 & n4123;
  assign n4125 = n3428 & n3444;
  assign n4126 = ~n3436 & n4124;
  assign n4127 = ~n4118 & ~n32277;
  assign n4128 = ~n3752 & n4127;
  assign n4129 = ~n32228 & n4128;
  assign n4130 = ~n3746 & n4129;
  assign n4131 = n3754 & n4119;
  assign n4132 = ~n4116 & n4130;
  assign n4133 = ~pi82  & ~n4115;
  assign n4134 = pi83  & ~n4133;
  assign n4135 = ~pi83  & n4133;
  assign n4136 = n3756 & ~n4115;
  assign n4137 = ~n4134 & ~n32279;
  assign n4138 = ~n32278 & n4137;
  assign n4139 = ~n4120 & ~n4138;
  assign n4140 = ~n3444 & ~n4139;
  assign n4141 = ~n3754 & ~n4113;
  assign n4142 = ~n32276 & n4141;
  assign n4143 = ~n4107 & n4142;
  assign n4144 = ~n32279 & ~n4143;
  assign n4145 = pi84  & ~n4144;
  assign n4146 = ~pi84  & ~n4143;
  assign n4147 = ~pi84  & n4144;
  assign n4148 = ~n32279 & n4146;
  assign n4149 = ~n4145 & ~n32280;
  assign n4150 = n3444 & ~n4120;
  assign n4151 = n3444 & n4139;
  assign n4152 = ~n4138 & n4150;
  assign n4153 = ~n4149 & ~n32281;
  assign n4154 = ~n4140 & ~n4153;
  assign n4155 = ~n3116 & ~n4154;
  assign n4156 = n3116 & ~n4140;
  assign n4157 = ~n4153 & n4156;
  assign n4158 = ~n3759 & ~n32231;
  assign n4159 = ~n4115 & n4158;
  assign n4160 = n3764 & ~n4159;
  assign n4161 = ~n3764 & n4158;
  assign n4162 = ~n3764 & n4159;
  assign n4163 = ~n4115 & n4161;
  assign n4164 = ~n4160 & ~n32282;
  assign n4165 = ~n4157 & ~n4164;
  assign n4166 = ~n4155 & ~n4165;
  assign n4167 = ~n2833 & ~n4166;
  assign n4168 = ~n3779 & ~n3781;
  assign n4169 = ~n4115 & n4168;
  assign n4170 = ~n3790 & ~n4169;
  assign n4171 = ~n3781 & n3790;
  assign n4172 = ~n3779 & n4171;
  assign n4173 = n3790 & n4169;
  assign n4174 = ~n4115 & n4172;
  assign n4175 = ~n4170 & ~n32283;
  assign n4176 = n2833 & ~n4155;
  assign n4177 = n2833 & n4166;
  assign n4178 = ~n4165 & n4176;
  assign n4179 = ~n4175 & ~n32284;
  assign n4180 = ~n4167 & ~n4179;
  assign n4181 = ~n2536 & ~n4180;
  assign n4182 = n2536 & ~n4167;
  assign n4183 = ~n4179 & n4182;
  assign n4184 = ~n3793 & ~n32233;
  assign n4185 = ~n4115 & n4184;
  assign n4186 = ~n3803 & ~n4185;
  assign n4187 = ~n3793 & n3803;
  assign n4188 = ~n32233 & n4187;
  assign n4189 = n3803 & n4185;
  assign n4190 = ~n4115 & n4188;
  assign n4191 = n3803 & ~n4185;
  assign n4192 = ~n3803 & n4185;
  assign n4193 = ~n4191 & ~n4192;
  assign n4194 = ~n4186 & ~n32285;
  assign n4195 = ~n4183 & n32286;
  assign n4196 = ~n4181 & ~n4195;
  assign n4197 = ~n2283 & ~n4196;
  assign n4198 = ~n3806 & ~n3808;
  assign n4199 = ~n4115 & n4198;
  assign n4200 = ~n32236 & ~n4199;
  assign n4201 = ~n3808 & n32236;
  assign n4202 = ~n3806 & n4201;
  assign n4203 = n32236 & n4199;
  assign n4204 = ~n4115 & n4202;
  assign n4205 = ~n4200 & ~n32287;
  assign n4206 = n2283 & ~n4181;
  assign n4207 = n2283 & n4196;
  assign n4208 = ~n4195 & n4206;
  assign n4209 = ~n4205 & ~n32288;
  assign n4210 = ~n4197 & ~n4209;
  assign n4211 = ~n2021 & ~n4210;
  assign n4212 = n2021 & ~n4197;
  assign n4213 = ~n4209 & n4212;
  assign n4214 = ~n3823 & ~n32237;
  assign n4215 = ~n4115 & n4214;
  assign n4216 = ~n32239 & ~n4215;
  assign n4217 = n32239 & n4215;
  assign n4218 = ~n3823 & ~n32239;
  assign n4219 = ~n32237 & n4218;
  assign n4220 = ~n4115 & n4219;
  assign n4221 = n32239 & ~n4215;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = ~n4216 & ~n4217;
  assign n4224 = ~n4213 & ~n32289;
  assign n4225 = ~n4211 & ~n4224;
  assign n4226 = ~n1796 & ~n4225;
  assign n4227 = ~n3840 & ~n3842;
  assign n4228 = ~n4115 & n4227;
  assign n4229 = ~n32241 & ~n4228;
  assign n4230 = ~n3842 & n32241;
  assign n4231 = ~n3840 & n4230;
  assign n4232 = n32241 & n4228;
  assign n4233 = ~n4115 & n4231;
  assign n4234 = ~n4229 & ~n32290;
  assign n4235 = n1796 & ~n4211;
  assign n4236 = n1796 & n4225;
  assign n4237 = ~n4224 & n4235;
  assign n4238 = ~n4234 & ~n32291;
  assign n4239 = ~n4226 & ~n4238;
  assign n4240 = ~n1567 & ~n4239;
  assign n4241 = n1567 & ~n4226;
  assign n4242 = ~n4238 & n4241;
  assign n4243 = ~n3857 & ~n32242;
  assign n4244 = ~n4115 & n4243;
  assign n4245 = ~n32243 & n4244;
  assign n4246 = n32243 & ~n4244;
  assign n4247 = ~n3857 & n32243;
  assign n4248 = ~n32242 & n4247;
  assign n4249 = ~n4115 & n4248;
  assign n4250 = ~n32243 & ~n4244;
  assign n4251 = ~n4249 & ~n4250;
  assign n4252 = ~n4245 & ~n4246;
  assign n4253 = ~n4242 & ~n32292;
  assign n4254 = ~n4240 & ~n4253;
  assign n4255 = ~n1374 & ~n4254;
  assign n4256 = ~n3873 & ~n3875;
  assign n4257 = ~n4115 & n4256;
  assign n4258 = ~n32245 & ~n4257;
  assign n4259 = ~n3875 & n32245;
  assign n4260 = ~n3873 & n4259;
  assign n4261 = n32245 & n4257;
  assign n4262 = ~n4115 & n4260;
  assign n4263 = ~n4258 & ~n32293;
  assign n4264 = n1374 & ~n4240;
  assign n4265 = n1374 & n4254;
  assign n4266 = ~n4253 & n4264;
  assign n4267 = ~n4263 & ~n32294;
  assign n4268 = ~n4255 & ~n4267;
  assign n4269 = ~n1179 & ~n4268;
  assign n4270 = n1179 & ~n4255;
  assign n4271 = ~n4267 & n4270;
  assign n4272 = ~n3890 & ~n32246;
  assign n4273 = ~n4115 & n4272;
  assign n4274 = ~n32247 & n4273;
  assign n4275 = n32247 & ~n4273;
  assign n4276 = ~n32247 & ~n4273;
  assign n4277 = ~n3890 & n32247;
  assign n4278 = ~n32246 & n4277;
  assign n4279 = n32247 & n4273;
  assign n4280 = ~n4115 & n4278;
  assign n4281 = ~n4276 & ~n32295;
  assign n4282 = ~n4274 & ~n4275;
  assign n4283 = ~n4271 & ~n32296;
  assign n4284 = ~n4269 & ~n4283;
  assign n4285 = ~n1016 & ~n4284;
  assign n4286 = ~n3906 & ~n3908;
  assign n4287 = ~n4115 & n4286;
  assign n4288 = ~n32249 & ~n4287;
  assign n4289 = ~n3908 & n32249;
  assign n4290 = ~n3906 & n4289;
  assign n4291 = n32249 & n4287;
  assign n4292 = ~n4115 & n4290;
  assign n4293 = ~n4288 & ~n32297;
  assign n4294 = n1016 & ~n4269;
  assign n4295 = n1016 & n4284;
  assign n4296 = ~n4283 & n4294;
  assign n4297 = ~n4293 & ~n32298;
  assign n4298 = ~n4285 & ~n4297;
  assign n4299 = ~n855 & ~n4298;
  assign n4300 = n855 & ~n4285;
  assign n4301 = ~n4297 & n4300;
  assign n4302 = ~n3923 & ~n32250;
  assign n4303 = ~n3923 & ~n4115;
  assign n4304 = ~n32250 & n4303;
  assign n4305 = ~n4115 & n4302;
  assign n4306 = n32252 & ~n32299;
  assign n4307 = n3938 & n4303;
  assign n4308 = ~n32252 & n32299;
  assign n4309 = ~n3923 & n32252;
  assign n4310 = ~n32250 & n4309;
  assign n4311 = ~n4115 & n4310;
  assign n4312 = ~n32252 & ~n32299;
  assign n4313 = ~n4311 & ~n4312;
  assign n4314 = ~n4306 & ~n32300;
  assign n4315 = ~n4301 & ~n32301;
  assign n4316 = ~n4299 & ~n4315;
  assign n4317 = ~n720 & ~n4316;
  assign n4318 = ~n3940 & ~n3942;
  assign n4319 = ~n4115 & n4318;
  assign n4320 = ~n32254 & ~n4319;
  assign n4321 = ~n3942 & n32254;
  assign n4322 = ~n3940 & n4321;
  assign n4323 = n32254 & n4319;
  assign n4324 = ~n4115 & n4322;
  assign n4325 = ~n4320 & ~n32302;
  assign n4326 = n720 & ~n4299;
  assign n4327 = n720 & n4316;
  assign n4328 = ~n4315 & n4326;
  assign n4329 = ~n4325 & ~n32303;
  assign n4330 = ~n4317 & ~n4329;
  assign n4331 = ~n592 & ~n4330;
  assign n4332 = n592 & ~n4317;
  assign n4333 = ~n4329 & n4332;
  assign n4334 = ~n3957 & ~n32255;
  assign n4335 = ~n3957 & ~n4115;
  assign n4336 = ~n32255 & n4335;
  assign n4337 = ~n4115 & n4334;
  assign n4338 = ~n32257 & ~n32304;
  assign n4339 = ~n3957 & n32257;
  assign n4340 = ~n32255 & n4339;
  assign n4341 = n32257 & n32304;
  assign n4342 = ~n4115 & n4340;
  assign n4343 = n32257 & ~n32304;
  assign n4344 = n3972 & n4335;
  assign n4345 = ~n4343 & ~n4344;
  assign n4346 = ~n4338 & ~n32305;
  assign n4347 = ~n4333 & n32306;
  assign n4348 = ~n4331 & ~n4347;
  assign n4349 = ~n487 & ~n4348;
  assign n4350 = ~n3974 & ~n3976;
  assign n4351 = ~n4115 & n4350;
  assign n4352 = ~n32259 & ~n4351;
  assign n4353 = ~n3976 & n32259;
  assign n4354 = ~n3974 & n4353;
  assign n4355 = n32259 & n4351;
  assign n4356 = ~n4115 & n4354;
  assign n4357 = ~n4352 & ~n32307;
  assign n4358 = n487 & ~n4331;
  assign n4359 = n487 & n4348;
  assign n4360 = ~n4347 & n4358;
  assign n4361 = ~n4357 & ~n32308;
  assign n4362 = ~n4349 & ~n4361;
  assign n4363 = ~n393 & ~n4362;
  assign n4364 = n393 & ~n4349;
  assign n4365 = ~n4361 & n4364;
  assign n4366 = ~n3991 & ~n32261;
  assign n4367 = ~n3991 & ~n4115;
  assign n4368 = ~n32261 & n4367;
  assign n4369 = ~n4115 & n4366;
  assign n4370 = n3999 & ~n32309;
  assign n4371 = n4003 & n4367;
  assign n4372 = ~n3991 & n3999;
  assign n4373 = ~n32261 & n4372;
  assign n4374 = ~n4115 & n4373;
  assign n4375 = ~n3999 & ~n32309;
  assign n4376 = ~n4374 & ~n4375;
  assign n4377 = ~n4370 & ~n4371;
  assign n4378 = ~n4365 & ~n32310;
  assign n4379 = ~n4363 & ~n4378;
  assign n4380 = ~n321 & ~n4379;
  assign n4381 = ~n4005 & ~n4007;
  assign n4382 = ~n4115 & n4381;
  assign n4383 = ~n32263 & ~n4382;
  assign n4384 = ~n4007 & n32263;
  assign n4385 = ~n4005 & n4384;
  assign n4386 = n32263 & n4382;
  assign n4387 = ~n4115 & n4385;
  assign n4388 = ~n4383 & ~n32311;
  assign n4389 = n321 & ~n4363;
  assign n4390 = n321 & n4379;
  assign n4391 = ~n4378 & n4389;
  assign n4392 = ~n4388 & ~n32312;
  assign n4393 = ~n4380 & ~n4392;
  assign n4394 = ~n263 & ~n4393;
  assign n4395 = ~n4022 & ~n32264;
  assign n4396 = ~n4115 & n4395;
  assign n4397 = ~n32266 & ~n4396;
  assign n4398 = ~n4022 & n32266;
  assign n4399 = ~n32264 & n4398;
  assign n4400 = n32266 & n4396;
  assign n4401 = ~n4115 & n4399;
  assign n4402 = ~n4397 & ~n32313;
  assign n4403 = n263 & ~n4380;
  assign n4404 = ~n4392 & n4403;
  assign n4405 = ~n4402 & ~n4404;
  assign n4406 = ~n4394 & ~n4405;
  assign n4407 = ~n214 & ~n4406;
  assign n4408 = ~n4040 & ~n4042;
  assign n4409 = ~n4115 & n4408;
  assign n4410 = ~n32268 & ~n4409;
  assign n4411 = ~n4042 & n32268;
  assign n4412 = ~n4040 & n4411;
  assign n4413 = n32268 & n4409;
  assign n4414 = ~n4115 & n4412;
  assign n4415 = ~n4410 & ~n32314;
  assign n4416 = n214 & ~n4394;
  assign n4417 = n214 & n4406;
  assign n4418 = ~n4405 & n4416;
  assign n4419 = ~n4415 & ~n32315;
  assign n4420 = ~n4407 & ~n4419;
  assign n4421 = ~n197 & ~n4420;
  assign n4422 = n197 & ~n4407;
  assign n4423 = ~n4419 & n4422;
  assign n4424 = ~n4057 & ~n32270;
  assign n4425 = ~n4057 & ~n4115;
  assign n4426 = ~n32270 & n4425;
  assign n4427 = ~n4115 & n4424;
  assign n4428 = n4065 & ~n32316;
  assign n4429 = n4069 & n4425;
  assign n4430 = ~n4057 & n4065;
  assign n4431 = ~n32270 & n4430;
  assign n4432 = ~n4115 & n4431;
  assign n4433 = ~n4065 & ~n32316;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = ~n4428 & ~n4429;
  assign n4436 = ~n4423 & ~n32317;
  assign n4437 = ~n4421 & ~n4436;
  assign n4438 = ~n4071 & ~n4073;
  assign n4439 = ~n4115 & n4438;
  assign n4440 = ~n32272 & ~n4439;
  assign n4441 = ~n4073 & n32272;
  assign n4442 = ~n4071 & n4441;
  assign n4443 = n32272 & n4439;
  assign n4444 = ~n4115 & n4442;
  assign n4445 = ~n4440 & ~n32318;
  assign n4446 = ~n4087 & ~n32274;
  assign n4447 = ~n32274 & ~n4115;
  assign n4448 = ~n4087 & n4447;
  assign n4449 = ~n4115 & n4446;
  assign n4450 = ~n32276 & ~n32319;
  assign n4451 = ~n4445 & n4450;
  assign n4452 = ~n4437 & n4451;
  assign n4453 = n193 & ~n4452;
  assign n4454 = ~n4421 & n4445;
  assign n4455 = n4437 & n4445;
  assign n4456 = ~n4436 & n4454;
  assign n4457 = n4087 & ~n4447;
  assign n4458 = ~n193 & ~n4446;
  assign n4459 = ~n4457 & n4458;
  assign n4460 = ~n32320 & ~n4459;
  assign n4461 = ~n4453 & n4460;
  assign n4462 = pi80  & ~n4461;
  assign n4463 = ~pi78  & ~pi79 ;
  assign n4464 = ~pi80  & n4463;
  assign n4465 = ~n4462 & ~n4464;
  assign n4466 = ~n4115 & ~n4465;
  assign n4467 = ~pi80  & ~n4461;
  assign n4468 = pi81  & ~n4467;
  assign n4469 = ~pi81  & n4467;
  assign n4470 = n4117 & ~n4461;
  assign n4471 = ~n4468 & ~n32321;
  assign n4472 = ~n32226 & ~n32277;
  assign n4473 = ~n3733 & n4472;
  assign n4474 = ~n3752 & n4473;
  assign n4475 = ~n32228 & n4474;
  assign n4476 = n3738 & n3754;
  assign n4477 = ~n3746 & n4475;
  assign n4478 = ~n4464 & ~n32322;
  assign n4479 = ~n4113 & n4478;
  assign n4480 = ~n32276 & n4479;
  assign n4481 = ~n4107 & n4480;
  assign n4482 = n4115 & n4465;
  assign n4483 = ~n4462 & n4481;
  assign n4484 = n4471 & ~n32323;
  assign n4485 = ~n4466 & ~n4484;
  assign n4486 = ~n3754 & ~n4485;
  assign n4487 = n3754 & ~n4466;
  assign n4488 = ~n4484 & n4487;
  assign n4489 = ~n4115 & ~n4459;
  assign n4490 = ~n32320 & n4489;
  assign n4491 = ~n4453 & n4490;
  assign n4492 = ~n32321 & ~n4491;
  assign n4493 = pi82  & ~n4492;
  assign n4494 = ~pi82  & ~n4491;
  assign n4495 = ~pi82  & n4492;
  assign n4496 = ~n32321 & n4494;
  assign n4497 = ~n4493 & ~n32324;
  assign n4498 = ~n4488 & ~n4497;
  assign n4499 = ~n4486 & ~n4498;
  assign n4500 = ~n3444 & ~n4499;
  assign n4501 = n3444 & ~n4486;
  assign n4502 = ~n4498 & n4501;
  assign n4503 = n3444 & n4499;
  assign n4504 = ~n4120 & ~n32278;
  assign n4505 = ~n4461 & n4504;
  assign n4506 = n4137 & ~n4505;
  assign n4507 = ~n4137 & n4504;
  assign n4508 = ~n4137 & n4505;
  assign n4509 = ~n4461 & n4507;
  assign n4510 = ~n4506 & ~n32326;
  assign n4511 = ~n32325 & ~n4510;
  assign n4512 = ~n4500 & ~n4511;
  assign n4513 = ~n3116 & ~n4512;
  assign n4514 = n3116 & ~n4500;
  assign n4515 = ~n4511 & n4514;
  assign n4516 = ~n4140 & ~n32281;
  assign n4517 = ~n4140 & ~n4461;
  assign n4518 = ~n32281 & n4517;
  assign n4519 = ~n4461 & n4516;
  assign n4520 = n4149 & ~n32327;
  assign n4521 = n4153 & n4517;
  assign n4522 = n4149 & ~n32281;
  assign n4523 = ~n4140 & n4522;
  assign n4524 = ~n4461 & n4523;
  assign n4525 = ~n4149 & ~n32327;
  assign n4526 = ~n4524 & ~n4525;
  assign n4527 = ~n4520 & ~n4521;
  assign n4528 = ~n4515 & ~n32328;
  assign n4529 = ~n4513 & ~n4528;
  assign n4530 = ~n2833 & ~n4529;
  assign n4531 = n2833 & ~n4513;
  assign n4532 = ~n4528 & n4531;
  assign n4533 = n2833 & n4529;
  assign n4534 = ~n4155 & ~n4157;
  assign n4535 = ~n4461 & n4534;
  assign n4536 = ~n4164 & ~n4535;
  assign n4537 = ~n4155 & n4164;
  assign n4538 = ~n4157 & n4537;
  assign n4539 = n4164 & n4535;
  assign n4540 = ~n4461 & n4538;
  assign n4541 = n4164 & ~n4535;
  assign n4542 = ~n4164 & n4535;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = ~n4536 & ~n32330;
  assign n4545 = ~n32329 & n32331;
  assign n4546 = ~n4530 & ~n4545;
  assign n4547 = ~n2536 & ~n4546;
  assign n4548 = n2536 & ~n4530;
  assign n4549 = ~n4545 & n4548;
  assign n4550 = ~n4167 & ~n32284;
  assign n4551 = ~n4167 & ~n4461;
  assign n4552 = ~n32284 & n4551;
  assign n4553 = ~n4461 & n4550;
  assign n4554 = n4175 & ~n32332;
  assign n4555 = n4179 & n4551;
  assign n4556 = n4175 & ~n32284;
  assign n4557 = ~n4167 & n4556;
  assign n4558 = ~n4461 & n4557;
  assign n4559 = ~n4175 & ~n32332;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = ~n4554 & ~n4555;
  assign n4562 = ~n4549 & ~n32333;
  assign n4563 = ~n4547 & ~n4562;
  assign n4564 = ~n2283 & ~n4563;
  assign n4565 = n2283 & ~n4547;
  assign n4566 = ~n4562 & n4565;
  assign n4567 = n2283 & n4563;
  assign n4568 = ~n4181 & ~n4183;
  assign n4569 = ~n4461 & n4568;
  assign n4570 = ~n32286 & ~n4569;
  assign n4571 = n32286 & n4569;
  assign n4572 = ~n4181 & ~n32286;
  assign n4573 = ~n4183 & n4572;
  assign n4574 = ~n4461 & n4573;
  assign n4575 = n32286 & ~n4569;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = ~n4570 & ~n4571;
  assign n4578 = ~n32334 & ~n32335;
  assign n4579 = ~n4564 & ~n4578;
  assign n4580 = ~n2021 & ~n4579;
  assign n4581 = n2021 & ~n4564;
  assign n4582 = ~n4578 & n4581;
  assign n4583 = ~n4197 & ~n32288;
  assign n4584 = ~n4197 & ~n4461;
  assign n4585 = ~n32288 & n4584;
  assign n4586 = ~n4461 & n4583;
  assign n4587 = n4205 & ~n32336;
  assign n4588 = n4209 & n4584;
  assign n4589 = n4205 & ~n32288;
  assign n4590 = ~n4197 & n4589;
  assign n4591 = ~n4461 & n4590;
  assign n4592 = ~n4205 & ~n32336;
  assign n4593 = ~n4591 & ~n4592;
  assign n4594 = ~n4587 & ~n4588;
  assign n4595 = ~n4582 & ~n32337;
  assign n4596 = ~n4580 & ~n4595;
  assign n4597 = ~n1796 & ~n4596;
  assign n4598 = n1796 & ~n4580;
  assign n4599 = ~n4595 & n4598;
  assign n4600 = n1796 & n4596;
  assign n4601 = ~n4211 & ~n4213;
  assign n4602 = ~n4461 & n4601;
  assign n4603 = ~n32289 & n4602;
  assign n4604 = n32289 & ~n4602;
  assign n4605 = ~n4211 & n32289;
  assign n4606 = ~n4213 & n4605;
  assign n4607 = ~n4461 & n4606;
  assign n4608 = ~n32289 & ~n4602;
  assign n4609 = ~n4607 & ~n4608;
  assign n4610 = ~n4603 & ~n4604;
  assign n4611 = ~n32338 & ~n32339;
  assign n4612 = ~n4597 & ~n4611;
  assign n4613 = ~n1567 & ~n4612;
  assign n4614 = n1567 & ~n4597;
  assign n4615 = ~n4611 & n4614;
  assign n4616 = ~n4226 & ~n32291;
  assign n4617 = ~n4226 & ~n4461;
  assign n4618 = ~n32291 & n4617;
  assign n4619 = ~n4461 & n4616;
  assign n4620 = n4234 & ~n32340;
  assign n4621 = n4238 & n4617;
  assign n4622 = n4234 & ~n32291;
  assign n4623 = ~n4226 & n4622;
  assign n4624 = ~n4461 & n4623;
  assign n4625 = ~n4234 & ~n32340;
  assign n4626 = ~n4624 & ~n4625;
  assign n4627 = ~n4620 & ~n4621;
  assign n4628 = ~n4615 & ~n32341;
  assign n4629 = ~n4613 & ~n4628;
  assign n4630 = ~n1374 & ~n4629;
  assign n4631 = n1374 & ~n4613;
  assign n4632 = ~n4628 & n4631;
  assign n4633 = n1374 & n4629;
  assign n4634 = ~n4240 & ~n4242;
  assign n4635 = ~n4461 & n4634;
  assign n4636 = ~n32292 & n4635;
  assign n4637 = n32292 & ~n4635;
  assign n4638 = ~n32292 & ~n4635;
  assign n4639 = ~n4240 & n32292;
  assign n4640 = ~n4242 & n4639;
  assign n4641 = n32292 & n4635;
  assign n4642 = ~n4461 & n4640;
  assign n4643 = ~n4638 & ~n32343;
  assign n4644 = ~n4636 & ~n4637;
  assign n4645 = ~n32342 & ~n32344;
  assign n4646 = ~n4630 & ~n4645;
  assign n4647 = ~n1179 & ~n4646;
  assign n4648 = n1179 & ~n4630;
  assign n4649 = ~n4645 & n4648;
  assign n4650 = ~n4255 & ~n32294;
  assign n4651 = ~n4255 & ~n4461;
  assign n4652 = ~n32294 & n4651;
  assign n4653 = ~n4461 & n4650;
  assign n4654 = n4263 & ~n32345;
  assign n4655 = n4267 & n4651;
  assign n4656 = n4263 & ~n32294;
  assign n4657 = ~n4255 & n4656;
  assign n4658 = ~n4461 & n4657;
  assign n4659 = ~n4263 & ~n32345;
  assign n4660 = ~n4658 & ~n4659;
  assign n4661 = ~n4654 & ~n4655;
  assign n4662 = ~n4649 & ~n32346;
  assign n4663 = ~n4647 & ~n4662;
  assign n4664 = ~n1016 & ~n4663;
  assign n4665 = n1016 & ~n4647;
  assign n4666 = ~n4662 & n4665;
  assign n4667 = n1016 & n4663;
  assign n4668 = ~n4269 & ~n4271;
  assign n4669 = ~n4269 & ~n4461;
  assign n4670 = ~n4271 & n4669;
  assign n4671 = ~n4461 & n4668;
  assign n4672 = n32296 & ~n32348;
  assign n4673 = n4283 & n4669;
  assign n4674 = ~n32296 & n32348;
  assign n4675 = ~n4269 & n32296;
  assign n4676 = ~n4271 & n4675;
  assign n4677 = ~n4461 & n4676;
  assign n4678 = ~n32296 & ~n32348;
  assign n4679 = ~n4677 & ~n4678;
  assign n4680 = ~n4672 & ~n32349;
  assign n4681 = ~n32347 & ~n32350;
  assign n4682 = ~n4664 & ~n4681;
  assign n4683 = ~n855 & ~n4682;
  assign n4684 = n855 & ~n4664;
  assign n4685 = ~n4681 & n4684;
  assign n4686 = ~n4285 & ~n32298;
  assign n4687 = ~n4285 & ~n4461;
  assign n4688 = ~n32298 & n4687;
  assign n4689 = ~n4461 & n4686;
  assign n4690 = n4293 & ~n32351;
  assign n4691 = n4297 & n4687;
  assign n4692 = n4293 & ~n32298;
  assign n4693 = ~n4285 & n4692;
  assign n4694 = ~n4461 & n4693;
  assign n4695 = ~n4293 & ~n32351;
  assign n4696 = ~n4694 & ~n4695;
  assign n4697 = ~n4690 & ~n4691;
  assign n4698 = ~n4685 & ~n32352;
  assign n4699 = ~n4683 & ~n4698;
  assign n4700 = ~n720 & ~n4699;
  assign n4701 = ~n4299 & ~n4301;
  assign n4702 = ~n4461 & n4701;
  assign n4703 = ~n32301 & ~n4702;
  assign n4704 = ~n4299 & n32301;
  assign n4705 = ~n4301 & n4704;
  assign n4706 = n32301 & n4702;
  assign n4707 = ~n4461 & n4705;
  assign n4708 = ~n4703 & ~n32353;
  assign n4709 = n720 & ~n4683;
  assign n4710 = ~n4698 & n4709;
  assign n4711 = n720 & n4699;
  assign n4712 = ~n4708 & ~n32354;
  assign n4713 = ~n4700 & ~n4712;
  assign n4714 = ~n592 & ~n4713;
  assign n4715 = n592 & ~n4700;
  assign n4716 = ~n4712 & n4715;
  assign n4717 = ~n4317 & ~n32303;
  assign n4718 = ~n4317 & ~n4461;
  assign n4719 = ~n32303 & n4718;
  assign n4720 = ~n4461 & n4717;
  assign n4721 = n4325 & ~n32355;
  assign n4722 = n4329 & n4718;
  assign n4723 = n4325 & ~n32303;
  assign n4724 = ~n4317 & n4723;
  assign n4725 = ~n4461 & n4724;
  assign n4726 = ~n4325 & ~n32355;
  assign n4727 = ~n4725 & ~n4726;
  assign n4728 = ~n4721 & ~n4722;
  assign n4729 = ~n4716 & ~n32356;
  assign n4730 = ~n4714 & ~n4729;
  assign n4731 = ~n487 & ~n4730;
  assign n4732 = ~n4331 & ~n4333;
  assign n4733 = ~n4461 & n4732;
  assign n4734 = n32306 & ~n4733;
  assign n4735 = ~n4331 & ~n32306;
  assign n4736 = ~n4333 & n4735;
  assign n4737 = ~n32306 & n4733;
  assign n4738 = ~n4461 & n4736;
  assign n4739 = ~n4734 & ~n32357;
  assign n4740 = n487 & ~n4714;
  assign n4741 = ~n4729 & n4740;
  assign n4742 = n487 & n4730;
  assign n4743 = ~n4739 & ~n32358;
  assign n4744 = ~n4731 & ~n4743;
  assign n4745 = ~n393 & ~n4744;
  assign n4746 = n393 & ~n4731;
  assign n4747 = ~n4743 & n4746;
  assign n4748 = ~n4349 & ~n32308;
  assign n4749 = ~n4349 & ~n4461;
  assign n4750 = ~n32308 & n4749;
  assign n4751 = ~n4461 & n4748;
  assign n4752 = n4357 & ~n32359;
  assign n4753 = n4361 & n4749;
  assign n4754 = n4357 & ~n32308;
  assign n4755 = ~n4349 & n4754;
  assign n4756 = ~n4461 & n4755;
  assign n4757 = ~n4357 & ~n32359;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = ~n4752 & ~n4753;
  assign n4760 = ~n4747 & ~n32360;
  assign n4761 = ~n4745 & ~n4760;
  assign n4762 = ~n321 & ~n4761;
  assign n4763 = ~n4363 & ~n4365;
  assign n4764 = ~n4461 & n4763;
  assign n4765 = ~n32310 & ~n4764;
  assign n4766 = ~n4363 & n32310;
  assign n4767 = ~n4365 & n4766;
  assign n4768 = n32310 & n4764;
  assign n4769 = ~n4461 & n4767;
  assign n4770 = ~n4765 & ~n32361;
  assign n4771 = n321 & ~n4745;
  assign n4772 = ~n4760 & n4771;
  assign n4773 = n321 & n4761;
  assign n4774 = ~n4770 & ~n32362;
  assign n4775 = ~n4762 & ~n4774;
  assign n4776 = ~n263 & ~n4775;
  assign n4777 = n263 & ~n4762;
  assign n4778 = ~n4774 & n4777;
  assign n4779 = ~n4380 & ~n32312;
  assign n4780 = ~n4380 & ~n4461;
  assign n4781 = ~n32312 & n4780;
  assign n4782 = ~n4461 & n4779;
  assign n4783 = n4388 & ~n32363;
  assign n4784 = n4392 & n4780;
  assign n4785 = n4388 & ~n32312;
  assign n4786 = ~n4380 & n4785;
  assign n4787 = ~n4461 & n4786;
  assign n4788 = ~n4388 & ~n32363;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = ~n4783 & ~n4784;
  assign n4791 = ~n4778 & ~n32364;
  assign n4792 = ~n4776 & ~n4791;
  assign n4793 = ~n214 & ~n4792;
  assign n4794 = n214 & ~n4776;
  assign n4795 = ~n4791 & n4794;
  assign n4796 = n214 & n4792;
  assign n4797 = ~n4394 & ~n4404;
  assign n4798 = ~n4394 & ~n4461;
  assign n4799 = ~n4404 & n4798;
  assign n4800 = ~n4461 & n4797;
  assign n4801 = n4402 & ~n32366;
  assign n4802 = n4405 & n4798;
  assign n4803 = ~n4394 & n4402;
  assign n4804 = ~n4404 & n4803;
  assign n4805 = ~n4461 & n4804;
  assign n4806 = ~n4402 & ~n32366;
  assign n4807 = ~n4805 & ~n4806;
  assign n4808 = ~n4801 & ~n4802;
  assign n4809 = ~n32365 & ~n32367;
  assign n4810 = ~n4793 & ~n4809;
  assign n4811 = ~n197 & ~n4810;
  assign n4812 = n197 & ~n4793;
  assign n4813 = ~n4809 & n4812;
  assign n4814 = ~n4407 & ~n32315;
  assign n4815 = ~n4407 & ~n4461;
  assign n4816 = ~n32315 & n4815;
  assign n4817 = ~n4461 & n4814;
  assign n4818 = n4415 & ~n32368;
  assign n4819 = n4419 & n4815;
  assign n4820 = n4415 & ~n32315;
  assign n4821 = ~n4407 & n4820;
  assign n4822 = ~n4461 & n4821;
  assign n4823 = ~n4415 & ~n32368;
  assign n4824 = ~n4822 & ~n4823;
  assign n4825 = ~n4818 & ~n4819;
  assign n4826 = ~n4813 & ~n32369;
  assign n4827 = ~n4811 & ~n4826;
  assign n4828 = ~n4421 & ~n4423;
  assign n4829 = ~n4461 & n4828;
  assign n4830 = ~n32317 & ~n4829;
  assign n4831 = ~n4421 & n32317;
  assign n4832 = ~n4423 & n4831;
  assign n4833 = n32317 & n4829;
  assign n4834 = ~n4461 & n4832;
  assign n4835 = ~n4830 & ~n32370;
  assign n4836 = ~n4437 & ~n4445;
  assign n4837 = ~n4445 & ~n4461;
  assign n4838 = ~n4437 & n4837;
  assign n4839 = ~n4461 & n4836;
  assign n4840 = ~n32320 & ~n32371;
  assign n4841 = ~n4835 & n4840;
  assign n4842 = ~n4827 & n4841;
  assign n4843 = n193 & ~n4842;
  assign n4844 = ~n4811 & n4835;
  assign n4845 = ~n4826 & n4844;
  assign n4846 = n4827 & n4835;
  assign n4847 = n4437 & ~n4837;
  assign n4848 = ~n193 & ~n4836;
  assign n4849 = ~n4847 & n4848;
  assign n4850 = ~n32372 & ~n4849;
  assign n4851 = ~n4843 & n4850;
  assign n4852 = pi78  & ~n4851;
  assign n4853 = ~pi76  & ~pi77 ;
  assign n4854 = ~pi78  & n4853;
  assign n4855 = ~n4852 & ~n4854;
  assign n4856 = ~n4461 & ~n4855;
  assign n4857 = ~n4096 & ~n32322;
  assign n4858 = ~n4097 & n4857;
  assign n4859 = ~n4113 & n4858;
  assign n4860 = ~n32276 & n4859;
  assign n4861 = n32274 & n4115;
  assign n4862 = ~n4107 & n4860;
  assign n4863 = ~n4854 & ~n32373;
  assign n4864 = ~n4459 & n4863;
  assign n4865 = ~n32320 & n4864;
  assign n4866 = ~n4453 & n4865;
  assign n4867 = n4461 & n4855;
  assign n4868 = ~n4852 & n4866;
  assign n4869 = ~pi78  & ~n4851;
  assign n4870 = pi79  & ~n4869;
  assign n4871 = ~pi79  & n4869;
  assign n4872 = n4463 & ~n4851;
  assign n4873 = ~n4870 & ~n32375;
  assign n4874 = ~n32374 & n4873;
  assign n4875 = ~n4856 & ~n4874;
  assign n4876 = ~n4115 & ~n4875;
  assign n4877 = ~n4461 & ~n4849;
  assign n4878 = ~n32372 & n4877;
  assign n4879 = ~n4843 & n4878;
  assign n4880 = ~n32375 & ~n4879;
  assign n4881 = pi80  & ~n4880;
  assign n4882 = ~pi80  & ~n4879;
  assign n4883 = ~pi80  & n4880;
  assign n4884 = ~n32375 & n4882;
  assign n4885 = ~n4881 & ~n32376;
  assign n4886 = n4115 & ~n4856;
  assign n4887 = n4115 & n4875;
  assign n4888 = ~n4874 & n4886;
  assign n4889 = ~n4885 & ~n32377;
  assign n4890 = ~n4876 & ~n4889;
  assign n4891 = ~n3754 & ~n4890;
  assign n4892 = n3754 & ~n4876;
  assign n4893 = ~n4889 & n4892;
  assign n4894 = ~n4466 & ~n32323;
  assign n4895 = ~n4851 & n4894;
  assign n4896 = n4471 & ~n4895;
  assign n4897 = ~n4471 & n4894;
  assign n4898 = ~n4471 & n4895;
  assign n4899 = ~n4851 & n4897;
  assign n4900 = ~n4896 & ~n32378;
  assign n4901 = ~n4893 & ~n4900;
  assign n4902 = ~n4891 & ~n4901;
  assign n4903 = ~n3444 & ~n4902;
  assign n4904 = ~n4486 & ~n4488;
  assign n4905 = ~n4851 & n4904;
  assign n4906 = ~n4497 & ~n4905;
  assign n4907 = ~n4488 & n4497;
  assign n4908 = ~n4486 & n4907;
  assign n4909 = n4497 & n4905;
  assign n4910 = ~n4851 & n4908;
  assign n4911 = ~n4906 & ~n32379;
  assign n4912 = n3444 & ~n4891;
  assign n4913 = n3444 & n4902;
  assign n4914 = ~n4901 & n4912;
  assign n4915 = ~n4911 & ~n32380;
  assign n4916 = ~n4903 & ~n4915;
  assign n4917 = ~n3116 & ~n4916;
  assign n4918 = n3116 & ~n4903;
  assign n4919 = ~n4915 & n4918;
  assign n4920 = ~n4500 & ~n32325;
  assign n4921 = ~n4851 & n4920;
  assign n4922 = ~n4510 & ~n4921;
  assign n4923 = ~n4500 & n4510;
  assign n4924 = ~n32325 & n4923;
  assign n4925 = n4510 & n4921;
  assign n4926 = ~n4851 & n4924;
  assign n4927 = n4510 & ~n4921;
  assign n4928 = ~n4510 & n4921;
  assign n4929 = ~n4927 & ~n4928;
  assign n4930 = ~n4922 & ~n32381;
  assign n4931 = ~n4919 & n32382;
  assign n4932 = ~n4917 & ~n4931;
  assign n4933 = ~n2833 & ~n4932;
  assign n4934 = ~n4513 & ~n4515;
  assign n4935 = ~n4851 & n4934;
  assign n4936 = ~n32328 & ~n4935;
  assign n4937 = ~n4515 & n32328;
  assign n4938 = ~n4513 & n4937;
  assign n4939 = n32328 & n4935;
  assign n4940 = ~n4851 & n4938;
  assign n4941 = ~n4936 & ~n32383;
  assign n4942 = n2833 & ~n4917;
  assign n4943 = n2833 & n4932;
  assign n4944 = ~n4931 & n4942;
  assign n4945 = ~n4941 & ~n32384;
  assign n4946 = ~n4933 & ~n4945;
  assign n4947 = ~n2536 & ~n4946;
  assign n4948 = n2536 & ~n4933;
  assign n4949 = ~n4945 & n4948;
  assign n4950 = ~n4530 & ~n32329;
  assign n4951 = ~n4851 & n4950;
  assign n4952 = ~n32331 & ~n4951;
  assign n4953 = n32331 & n4951;
  assign n4954 = ~n4530 & ~n32331;
  assign n4955 = ~n32329 & n4954;
  assign n4956 = ~n4851 & n4955;
  assign n4957 = n32331 & ~n4951;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = ~n4952 & ~n4953;
  assign n4960 = ~n4949 & ~n32385;
  assign n4961 = ~n4947 & ~n4960;
  assign n4962 = ~n2283 & ~n4961;
  assign n4963 = ~n4547 & ~n4549;
  assign n4964 = ~n4851 & n4963;
  assign n4965 = ~n32333 & ~n4964;
  assign n4966 = ~n4549 & n32333;
  assign n4967 = ~n4547 & n4966;
  assign n4968 = n32333 & n4964;
  assign n4969 = ~n4851 & n4967;
  assign n4970 = ~n4965 & ~n32386;
  assign n4971 = n2283 & ~n4947;
  assign n4972 = n2283 & n4961;
  assign n4973 = ~n4960 & n4971;
  assign n4974 = ~n4970 & ~n32387;
  assign n4975 = ~n4962 & ~n4974;
  assign n4976 = ~n2021 & ~n4975;
  assign n4977 = n2021 & ~n4962;
  assign n4978 = ~n4974 & n4977;
  assign n4979 = ~n4564 & ~n32334;
  assign n4980 = ~n4851 & n4979;
  assign n4981 = ~n32335 & n4980;
  assign n4982 = n32335 & ~n4980;
  assign n4983 = ~n4564 & n32335;
  assign n4984 = ~n32334 & n4983;
  assign n4985 = ~n4851 & n4984;
  assign n4986 = ~n32335 & ~n4980;
  assign n4987 = ~n4985 & ~n4986;
  assign n4988 = ~n4981 & ~n4982;
  assign n4989 = ~n4978 & ~n32388;
  assign n4990 = ~n4976 & ~n4989;
  assign n4991 = ~n1796 & ~n4990;
  assign n4992 = ~n4580 & ~n4582;
  assign n4993 = ~n4851 & n4992;
  assign n4994 = ~n32337 & ~n4993;
  assign n4995 = ~n4582 & n32337;
  assign n4996 = ~n4580 & n4995;
  assign n4997 = n32337 & n4993;
  assign n4998 = ~n4851 & n4996;
  assign n4999 = ~n4994 & ~n32389;
  assign n5000 = n1796 & ~n4976;
  assign n5001 = n1796 & n4990;
  assign n5002 = ~n4989 & n5000;
  assign n5003 = ~n4999 & ~n32390;
  assign n5004 = ~n4991 & ~n5003;
  assign n5005 = ~n1567 & ~n5004;
  assign n5006 = n1567 & ~n4991;
  assign n5007 = ~n5003 & n5006;
  assign n5008 = ~n4597 & ~n32338;
  assign n5009 = ~n4851 & n5008;
  assign n5010 = ~n32339 & n5009;
  assign n5011 = n32339 & ~n5009;
  assign n5012 = ~n32339 & ~n5009;
  assign n5013 = ~n4597 & n32339;
  assign n5014 = ~n32338 & n5013;
  assign n5015 = n32339 & n5009;
  assign n5016 = ~n4851 & n5014;
  assign n5017 = ~n5012 & ~n32391;
  assign n5018 = ~n5010 & ~n5011;
  assign n5019 = ~n5007 & ~n32392;
  assign n5020 = ~n5005 & ~n5019;
  assign n5021 = ~n1374 & ~n5020;
  assign n5022 = ~n4613 & ~n4615;
  assign n5023 = ~n4851 & n5022;
  assign n5024 = ~n32341 & ~n5023;
  assign n5025 = ~n4615 & n32341;
  assign n5026 = ~n4613 & n5025;
  assign n5027 = n32341 & n5023;
  assign n5028 = ~n4851 & n5026;
  assign n5029 = ~n5024 & ~n32393;
  assign n5030 = n1374 & ~n5005;
  assign n5031 = n1374 & n5020;
  assign n5032 = ~n5019 & n5030;
  assign n5033 = ~n5029 & ~n32394;
  assign n5034 = ~n5021 & ~n5033;
  assign n5035 = ~n1179 & ~n5034;
  assign n5036 = n1179 & ~n5021;
  assign n5037 = ~n5033 & n5036;
  assign n5038 = ~n4630 & ~n32342;
  assign n5039 = ~n4630 & ~n4851;
  assign n5040 = ~n32342 & n5039;
  assign n5041 = ~n4851 & n5038;
  assign n5042 = n32344 & ~n32395;
  assign n5043 = n4645 & n5039;
  assign n5044 = ~n32344 & n32395;
  assign n5045 = ~n4630 & n32344;
  assign n5046 = ~n32342 & n5045;
  assign n5047 = ~n4851 & n5046;
  assign n5048 = ~n32344 & ~n32395;
  assign n5049 = ~n5047 & ~n5048;
  assign n5050 = ~n5042 & ~n32396;
  assign n5051 = ~n5037 & ~n32397;
  assign n5052 = ~n5035 & ~n5051;
  assign n5053 = ~n1016 & ~n5052;
  assign n5054 = ~n4647 & ~n4649;
  assign n5055 = ~n4851 & n5054;
  assign n5056 = ~n32346 & ~n5055;
  assign n5057 = ~n4649 & n32346;
  assign n5058 = ~n4647 & n5057;
  assign n5059 = n32346 & n5055;
  assign n5060 = ~n4851 & n5058;
  assign n5061 = ~n5056 & ~n32398;
  assign n5062 = n1016 & ~n5035;
  assign n5063 = n1016 & n5052;
  assign n5064 = ~n5051 & n5062;
  assign n5065 = ~n5061 & ~n32399;
  assign n5066 = ~n5053 & ~n5065;
  assign n5067 = ~n855 & ~n5066;
  assign n5068 = ~n4664 & ~n32347;
  assign n5069 = ~n4851 & n5068;
  assign n5070 = ~n32350 & ~n5069;
  assign n5071 = ~n4664 & n32350;
  assign n5072 = ~n32347 & n5071;
  assign n5073 = n32350 & n5069;
  assign n5074 = ~n4851 & n5072;
  assign n5075 = ~n5070 & ~n32400;
  assign n5076 = n855 & ~n5053;
  assign n5077 = ~n5065 & n5076;
  assign n5078 = ~n5075 & ~n5077;
  assign n5079 = ~n5067 & ~n5078;
  assign n5080 = ~n720 & ~n5079;
  assign n5081 = ~n4683 & ~n4685;
  assign n5082 = ~n4851 & n5081;
  assign n5083 = ~n32352 & ~n5082;
  assign n5084 = ~n4685 & n32352;
  assign n5085 = ~n4683 & n5084;
  assign n5086 = n32352 & n5082;
  assign n5087 = ~n4851 & n5085;
  assign n5088 = ~n5083 & ~n32401;
  assign n5089 = n720 & ~n5067;
  assign n5090 = n720 & n5079;
  assign n5091 = ~n5078 & n5089;
  assign n5092 = ~n5088 & ~n32402;
  assign n5093 = ~n5080 & ~n5092;
  assign n5094 = ~n592 & ~n5093;
  assign n5095 = n592 & ~n5080;
  assign n5096 = ~n5092 & n5095;
  assign n5097 = ~n4700 & ~n32354;
  assign n5098 = ~n4700 & ~n4851;
  assign n5099 = ~n32354 & n5098;
  assign n5100 = ~n4851 & n5097;
  assign n5101 = n4708 & ~n32403;
  assign n5102 = n4712 & n5098;
  assign n5103 = ~n4700 & n4708;
  assign n5104 = ~n32354 & n5103;
  assign n5105 = ~n4851 & n5104;
  assign n5106 = ~n4708 & ~n32403;
  assign n5107 = ~n5105 & ~n5106;
  assign n5108 = ~n5101 & ~n5102;
  assign n5109 = ~n5096 & ~n32404;
  assign n5110 = ~n5094 & ~n5109;
  assign n5111 = ~n487 & ~n5110;
  assign n5112 = ~n4714 & ~n4716;
  assign n5113 = ~n4851 & n5112;
  assign n5114 = ~n32356 & ~n5113;
  assign n5115 = ~n4716 & n32356;
  assign n5116 = ~n4714 & n5115;
  assign n5117 = n32356 & n5113;
  assign n5118 = ~n4851 & n5116;
  assign n5119 = ~n5114 & ~n32405;
  assign n5120 = n487 & ~n5094;
  assign n5121 = n487 & n5110;
  assign n5122 = ~n5109 & n5120;
  assign n5123 = ~n5119 & ~n32406;
  assign n5124 = ~n5111 & ~n5123;
  assign n5125 = ~n393 & ~n5124;
  assign n5126 = n393 & ~n5111;
  assign n5127 = ~n5123 & n5126;
  assign n5128 = ~n4731 & ~n32358;
  assign n5129 = ~n4731 & ~n4851;
  assign n5130 = ~n32358 & n5129;
  assign n5131 = ~n4851 & n5128;
  assign n5132 = n4739 & ~n32407;
  assign n5133 = n4743 & n5129;
  assign n5134 = ~n4731 & n4739;
  assign n5135 = ~n32358 & n5134;
  assign n5136 = ~n4851 & n5135;
  assign n5137 = ~n4739 & ~n32407;
  assign n5138 = ~n5136 & ~n5137;
  assign n5139 = ~n5132 & ~n5133;
  assign n5140 = ~n5127 & ~n32408;
  assign n5141 = ~n5125 & ~n5140;
  assign n5142 = ~n321 & ~n5141;
  assign n5143 = ~n4745 & ~n4747;
  assign n5144 = ~n4851 & n5143;
  assign n5145 = ~n32360 & ~n5144;
  assign n5146 = ~n4747 & n32360;
  assign n5147 = ~n4745 & n5146;
  assign n5148 = n32360 & n5144;
  assign n5149 = ~n4851 & n5147;
  assign n5150 = ~n5145 & ~n32409;
  assign n5151 = n321 & ~n5125;
  assign n5152 = n321 & n5141;
  assign n5153 = ~n5140 & n5151;
  assign n5154 = ~n5150 & ~n32410;
  assign n5155 = ~n5142 & ~n5154;
  assign n5156 = ~n263 & ~n5155;
  assign n5157 = n263 & ~n5142;
  assign n5158 = ~n5154 & n5157;
  assign n5159 = ~n4762 & ~n32362;
  assign n5160 = ~n4762 & ~n4851;
  assign n5161 = ~n32362 & n5160;
  assign n5162 = ~n4851 & n5159;
  assign n5163 = n4770 & ~n32411;
  assign n5164 = n4774 & n5160;
  assign n5165 = ~n4762 & n4770;
  assign n5166 = ~n32362 & n5165;
  assign n5167 = ~n4851 & n5166;
  assign n5168 = ~n4770 & ~n32411;
  assign n5169 = ~n5167 & ~n5168;
  assign n5170 = ~n5163 & ~n5164;
  assign n5171 = ~n5158 & ~n32412;
  assign n5172 = ~n5156 & ~n5171;
  assign n5173 = ~n214 & ~n5172;
  assign n5174 = ~n4776 & ~n4778;
  assign n5175 = ~n4851 & n5174;
  assign n5176 = ~n32364 & ~n5175;
  assign n5177 = ~n4778 & n32364;
  assign n5178 = ~n4776 & n5177;
  assign n5179 = n32364 & n5175;
  assign n5180 = ~n4851 & n5178;
  assign n5181 = ~n5176 & ~n32413;
  assign n5182 = n214 & ~n5156;
  assign n5183 = n214 & n5172;
  assign n5184 = ~n5171 & n5182;
  assign n5185 = ~n5181 & ~n32414;
  assign n5186 = ~n5173 & ~n5185;
  assign n5187 = ~n197 & ~n5186;
  assign n5188 = ~n4793 & ~n32365;
  assign n5189 = ~n4851 & n5188;
  assign n5190 = ~n32367 & ~n5189;
  assign n5191 = ~n4793 & n32367;
  assign n5192 = ~n32365 & n5191;
  assign n5193 = n32367 & n5189;
  assign n5194 = ~n4851 & n5192;
  assign n5195 = ~n5190 & ~n32415;
  assign n5196 = n197 & ~n5173;
  assign n5197 = ~n5185 & n5196;
  assign n5198 = ~n5195 & ~n5197;
  assign n5199 = ~n5187 & ~n5198;
  assign n5200 = ~n4811 & ~n4813;
  assign n5201 = ~n4851 & n5200;
  assign n5202 = ~n32369 & ~n5201;
  assign n5203 = ~n4813 & n32369;
  assign n5204 = ~n4811 & n5203;
  assign n5205 = n32369 & n5201;
  assign n5206 = ~n4851 & n5204;
  assign n5207 = ~n5202 & ~n32416;
  assign n5208 = ~n4827 & ~n4835;
  assign n5209 = ~n4835 & ~n4851;
  assign n5210 = ~n4827 & n5209;
  assign n5211 = ~n4851 & n5208;
  assign n5212 = ~n32372 & ~n32417;
  assign n5213 = ~n5207 & n5212;
  assign n5214 = ~n5199 & n5213;
  assign n5215 = n193 & ~n5214;
  assign n5216 = ~n5187 & n5207;
  assign n5217 = n5199 & n5207;
  assign n5218 = ~n5198 & n5216;
  assign n5219 = n4827 & ~n5209;
  assign n5220 = ~n193 & ~n5208;
  assign n5221 = ~n5219 & n5220;
  assign n5222 = ~n32418 & ~n5221;
  assign n5223 = ~n5215 & n5222;
  assign n5224 = pi76  & ~n5223;
  assign n5225 = ~pi74  & ~pi75 ;
  assign n5226 = ~pi76  & n5225;
  assign n5227 = ~n5224 & ~n5226;
  assign n5228 = ~n4851 & ~n5227;
  assign n5229 = ~pi76  & ~n5223;
  assign n5230 = pi77  & ~n5229;
  assign n5231 = ~pi77  & n5229;
  assign n5232 = n4853 & ~n5223;
  assign n5233 = ~n5230 & ~n32419;
  assign n5234 = ~n32318 & ~n32373;
  assign n5235 = ~n4440 & n5234;
  assign n5236 = ~n4459 & n5235;
  assign n5237 = ~n32320 & n5236;
  assign n5238 = n4445 & n4461;
  assign n5239 = ~n4453 & n5237;
  assign n5240 = ~n5226 & ~n32420;
  assign n5241 = ~n4849 & n5240;
  assign n5242 = ~n32372 & n5241;
  assign n5243 = ~n4843 & n5242;
  assign n5244 = n4851 & n5227;
  assign n5245 = ~n5224 & n5243;
  assign n5246 = n5233 & ~n32421;
  assign n5247 = ~n5228 & ~n5246;
  assign n5248 = ~n4461 & ~n5247;
  assign n5249 = n4461 & ~n5228;
  assign n5250 = ~n5246 & n5249;
  assign n5251 = ~n4851 & ~n5221;
  assign n5252 = ~n32418 & n5251;
  assign n5253 = ~n5215 & n5252;
  assign n5254 = ~n32419 & ~n5253;
  assign n5255 = pi78  & ~n5254;
  assign n5256 = ~pi78  & ~n5253;
  assign n5257 = ~pi78  & n5254;
  assign n5258 = ~n32419 & n5256;
  assign n5259 = ~n5255 & ~n32422;
  assign n5260 = ~n5250 & ~n5259;
  assign n5261 = ~n5248 & ~n5260;
  assign n5262 = ~n4115 & ~n5261;
  assign n5263 = n4115 & ~n5248;
  assign n5264 = ~n5260 & n5263;
  assign n5265 = n4115 & n5261;
  assign n5266 = ~n4856 & ~n32374;
  assign n5267 = ~n5223 & n5266;
  assign n5268 = n4873 & ~n5267;
  assign n5269 = ~n4873 & n5266;
  assign n5270 = ~n4873 & n5267;
  assign n5271 = ~n5223 & n5269;
  assign n5272 = ~n5268 & ~n32424;
  assign n5273 = ~n32423 & ~n5272;
  assign n5274 = ~n5262 & ~n5273;
  assign n5275 = ~n3754 & ~n5274;
  assign n5276 = n3754 & ~n5262;
  assign n5277 = ~n5273 & n5276;
  assign n5278 = ~n4876 & ~n32377;
  assign n5279 = ~n4876 & ~n5223;
  assign n5280 = ~n32377 & n5279;
  assign n5281 = ~n5223 & n5278;
  assign n5282 = n4885 & ~n32425;
  assign n5283 = n4889 & n5279;
  assign n5284 = n4885 & ~n32377;
  assign n5285 = ~n4876 & n5284;
  assign n5286 = ~n5223 & n5285;
  assign n5287 = ~n4885 & ~n32425;
  assign n5288 = ~n5286 & ~n5287;
  assign n5289 = ~n5282 & ~n5283;
  assign n5290 = ~n5277 & ~n32426;
  assign n5291 = ~n5275 & ~n5290;
  assign n5292 = ~n3444 & ~n5291;
  assign n5293 = n3444 & ~n5275;
  assign n5294 = ~n5290 & n5293;
  assign n5295 = n3444 & n5291;
  assign n5296 = ~n4891 & ~n4893;
  assign n5297 = ~n5223 & n5296;
  assign n5298 = ~n4900 & ~n5297;
  assign n5299 = ~n4891 & n4900;
  assign n5300 = ~n4893 & n5299;
  assign n5301 = n4900 & n5297;
  assign n5302 = ~n5223 & n5300;
  assign n5303 = n4900 & ~n5297;
  assign n5304 = ~n4900 & n5297;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = ~n5298 & ~n32428;
  assign n5307 = ~n32427 & n32429;
  assign n5308 = ~n5292 & ~n5307;
  assign n5309 = ~n3116 & ~n5308;
  assign n5310 = n3116 & ~n5292;
  assign n5311 = ~n5307 & n5310;
  assign n5312 = ~n4903 & ~n32380;
  assign n5313 = ~n4903 & ~n5223;
  assign n5314 = ~n32380 & n5313;
  assign n5315 = ~n5223 & n5312;
  assign n5316 = n4911 & ~n32430;
  assign n5317 = n4915 & n5313;
  assign n5318 = n4911 & ~n32380;
  assign n5319 = ~n4903 & n5318;
  assign n5320 = ~n5223 & n5319;
  assign n5321 = ~n4911 & ~n32430;
  assign n5322 = ~n5320 & ~n5321;
  assign n5323 = ~n5316 & ~n5317;
  assign n5324 = ~n5311 & ~n32431;
  assign n5325 = ~n5309 & ~n5324;
  assign n5326 = ~n2833 & ~n5325;
  assign n5327 = n2833 & ~n5309;
  assign n5328 = ~n5324 & n5327;
  assign n5329 = n2833 & n5325;
  assign n5330 = ~n4917 & ~n4919;
  assign n5331 = ~n5223 & n5330;
  assign n5332 = ~n32382 & ~n5331;
  assign n5333 = n32382 & n5331;
  assign n5334 = ~n4917 & ~n32382;
  assign n5335 = ~n4919 & n5334;
  assign n5336 = ~n5223 & n5335;
  assign n5337 = n32382 & ~n5331;
  assign n5338 = ~n5336 & ~n5337;
  assign n5339 = ~n5332 & ~n5333;
  assign n5340 = ~n32432 & ~n32433;
  assign n5341 = ~n5326 & ~n5340;
  assign n5342 = ~n2536 & ~n5341;
  assign n5343 = n2536 & ~n5326;
  assign n5344 = ~n5340 & n5343;
  assign n5345 = ~n4933 & ~n32384;
  assign n5346 = ~n4933 & ~n5223;
  assign n5347 = ~n32384 & n5346;
  assign n5348 = ~n5223 & n5345;
  assign n5349 = n4941 & ~n32434;
  assign n5350 = n4945 & n5346;
  assign n5351 = n4941 & ~n32384;
  assign n5352 = ~n4933 & n5351;
  assign n5353 = ~n5223 & n5352;
  assign n5354 = ~n4941 & ~n32434;
  assign n5355 = ~n5353 & ~n5354;
  assign n5356 = ~n5349 & ~n5350;
  assign n5357 = ~n5344 & ~n32435;
  assign n5358 = ~n5342 & ~n5357;
  assign n5359 = ~n2283 & ~n5358;
  assign n5360 = n2283 & ~n5342;
  assign n5361 = ~n5357 & n5360;
  assign n5362 = n2283 & n5358;
  assign n5363 = ~n4947 & ~n4949;
  assign n5364 = ~n5223 & n5363;
  assign n5365 = ~n32385 & n5364;
  assign n5366 = n32385 & ~n5364;
  assign n5367 = ~n4947 & n32385;
  assign n5368 = ~n4949 & n5367;
  assign n5369 = ~n5223 & n5368;
  assign n5370 = ~n32385 & ~n5364;
  assign n5371 = ~n5369 & ~n5370;
  assign n5372 = ~n5365 & ~n5366;
  assign n5373 = ~n32436 & ~n32437;
  assign n5374 = ~n5359 & ~n5373;
  assign n5375 = ~n2021 & ~n5374;
  assign n5376 = n2021 & ~n5359;
  assign n5377 = ~n5373 & n5376;
  assign n5378 = ~n4962 & ~n32387;
  assign n5379 = ~n4962 & ~n5223;
  assign n5380 = ~n32387 & n5379;
  assign n5381 = ~n5223 & n5378;
  assign n5382 = n4970 & ~n32438;
  assign n5383 = n4974 & n5379;
  assign n5384 = n4970 & ~n32387;
  assign n5385 = ~n4962 & n5384;
  assign n5386 = ~n5223 & n5385;
  assign n5387 = ~n4970 & ~n32438;
  assign n5388 = ~n5386 & ~n5387;
  assign n5389 = ~n5382 & ~n5383;
  assign n5390 = ~n5377 & ~n32439;
  assign n5391 = ~n5375 & ~n5390;
  assign n5392 = ~n1796 & ~n5391;
  assign n5393 = n1796 & ~n5375;
  assign n5394 = ~n5390 & n5393;
  assign n5395 = n1796 & n5391;
  assign n5396 = ~n4976 & ~n4978;
  assign n5397 = ~n5223 & n5396;
  assign n5398 = ~n32388 & n5397;
  assign n5399 = n32388 & ~n5397;
  assign n5400 = ~n32388 & ~n5397;
  assign n5401 = ~n4976 & n32388;
  assign n5402 = ~n4978 & n5401;
  assign n5403 = n32388 & n5397;
  assign n5404 = ~n5223 & n5402;
  assign n5405 = ~n5400 & ~n32441;
  assign n5406 = ~n5398 & ~n5399;
  assign n5407 = ~n32440 & ~n32442;
  assign n5408 = ~n5392 & ~n5407;
  assign n5409 = ~n1567 & ~n5408;
  assign n5410 = n1567 & ~n5392;
  assign n5411 = ~n5407 & n5410;
  assign n5412 = ~n4991 & ~n32390;
  assign n5413 = ~n4991 & ~n5223;
  assign n5414 = ~n32390 & n5413;
  assign n5415 = ~n5223 & n5412;
  assign n5416 = n4999 & ~n32443;
  assign n5417 = n5003 & n5413;
  assign n5418 = n4999 & ~n32390;
  assign n5419 = ~n4991 & n5418;
  assign n5420 = ~n5223 & n5419;
  assign n5421 = ~n4999 & ~n32443;
  assign n5422 = ~n5420 & ~n5421;
  assign n5423 = ~n5416 & ~n5417;
  assign n5424 = ~n5411 & ~n32444;
  assign n5425 = ~n5409 & ~n5424;
  assign n5426 = ~n1374 & ~n5425;
  assign n5427 = n1374 & ~n5409;
  assign n5428 = ~n5424 & n5427;
  assign n5429 = n1374 & n5425;
  assign n5430 = ~n5005 & ~n5007;
  assign n5431 = ~n5005 & ~n5223;
  assign n5432 = ~n5007 & n5431;
  assign n5433 = ~n5223 & n5430;
  assign n5434 = n32392 & ~n32446;
  assign n5435 = n5019 & n5431;
  assign n5436 = ~n32392 & n32446;
  assign n5437 = ~n5005 & n32392;
  assign n5438 = ~n5007 & n5437;
  assign n5439 = ~n5223 & n5438;
  assign n5440 = ~n32392 & ~n32446;
  assign n5441 = ~n5439 & ~n5440;
  assign n5442 = ~n5434 & ~n32447;
  assign n5443 = ~n32445 & ~n32448;
  assign n5444 = ~n5426 & ~n5443;
  assign n5445 = ~n1179 & ~n5444;
  assign n5446 = n1179 & ~n5426;
  assign n5447 = ~n5443 & n5446;
  assign n5448 = ~n5021 & ~n32394;
  assign n5449 = ~n5021 & ~n5223;
  assign n5450 = ~n32394 & n5449;
  assign n5451 = ~n5223 & n5448;
  assign n5452 = n5029 & ~n32449;
  assign n5453 = n5033 & n5449;
  assign n5454 = n5029 & ~n32394;
  assign n5455 = ~n5021 & n5454;
  assign n5456 = ~n5223 & n5455;
  assign n5457 = ~n5029 & ~n32449;
  assign n5458 = ~n5456 & ~n5457;
  assign n5459 = ~n5452 & ~n5453;
  assign n5460 = ~n5447 & ~n32450;
  assign n5461 = ~n5445 & ~n5460;
  assign n5462 = ~n1016 & ~n5461;
  assign n5463 = ~n5035 & ~n5037;
  assign n5464 = ~n5223 & n5463;
  assign n5465 = ~n32397 & ~n5464;
  assign n5466 = ~n5035 & n32397;
  assign n5467 = ~n5037 & n5466;
  assign n5468 = n32397 & n5464;
  assign n5469 = ~n5223 & n5467;
  assign n5470 = ~n5465 & ~n32451;
  assign n5471 = n1016 & ~n5445;
  assign n5472 = ~n5460 & n5471;
  assign n5473 = n1016 & n5461;
  assign n5474 = ~n5470 & ~n32452;
  assign n5475 = ~n5462 & ~n5474;
  assign n5476 = ~n855 & ~n5475;
  assign n5477 = n855 & ~n5462;
  assign n5478 = ~n5474 & n5477;
  assign n5479 = ~n5053 & ~n32399;
  assign n5480 = ~n5053 & ~n5223;
  assign n5481 = ~n32399 & n5480;
  assign n5482 = ~n5223 & n5479;
  assign n5483 = n5061 & ~n32453;
  assign n5484 = n5065 & n5480;
  assign n5485 = n5061 & ~n32399;
  assign n5486 = ~n5053 & n5485;
  assign n5487 = ~n5223 & n5486;
  assign n5488 = ~n5061 & ~n32453;
  assign n5489 = ~n5487 & ~n5488;
  assign n5490 = ~n5483 & ~n5484;
  assign n5491 = ~n5478 & ~n32454;
  assign n5492 = ~n5476 & ~n5491;
  assign n5493 = ~n720 & ~n5492;
  assign n5494 = n720 & ~n5476;
  assign n5495 = ~n5491 & n5494;
  assign n5496 = n720 & n5492;
  assign n5497 = ~n5067 & ~n5077;
  assign n5498 = ~n5067 & ~n5223;
  assign n5499 = ~n5077 & n5498;
  assign n5500 = ~n5223 & n5497;
  assign n5501 = n5075 & ~n32456;
  assign n5502 = n5078 & n5498;
  assign n5503 = ~n5067 & n5075;
  assign n5504 = ~n5077 & n5503;
  assign n5505 = ~n5223 & n5504;
  assign n5506 = ~n5075 & ~n32456;
  assign n5507 = ~n5505 & ~n5506;
  assign n5508 = ~n5501 & ~n5502;
  assign n5509 = ~n32455 & ~n32457;
  assign n5510 = ~n5493 & ~n5509;
  assign n5511 = ~n592 & ~n5510;
  assign n5512 = n592 & ~n5493;
  assign n5513 = ~n5509 & n5512;
  assign n5514 = ~n5080 & ~n32402;
  assign n5515 = ~n5080 & ~n5223;
  assign n5516 = ~n32402 & n5515;
  assign n5517 = ~n5223 & n5514;
  assign n5518 = n5088 & ~n32458;
  assign n5519 = n5092 & n5515;
  assign n5520 = n5088 & ~n32402;
  assign n5521 = ~n5080 & n5520;
  assign n5522 = ~n5223 & n5521;
  assign n5523 = ~n5088 & ~n32458;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = ~n5518 & ~n5519;
  assign n5526 = ~n5513 & ~n32459;
  assign n5527 = ~n5511 & ~n5526;
  assign n5528 = ~n487 & ~n5527;
  assign n5529 = ~n5094 & ~n5096;
  assign n5530 = ~n5223 & n5529;
  assign n5531 = ~n32404 & ~n5530;
  assign n5532 = ~n5094 & n32404;
  assign n5533 = ~n5096 & n5532;
  assign n5534 = n32404 & n5530;
  assign n5535 = ~n5223 & n5533;
  assign n5536 = ~n5531 & ~n32460;
  assign n5537 = n487 & ~n5511;
  assign n5538 = ~n5526 & n5537;
  assign n5539 = n487 & n5527;
  assign n5540 = ~n5536 & ~n32461;
  assign n5541 = ~n5528 & ~n5540;
  assign n5542 = ~n393 & ~n5541;
  assign n5543 = n393 & ~n5528;
  assign n5544 = ~n5540 & n5543;
  assign n5545 = ~n5111 & ~n32406;
  assign n5546 = ~n5111 & ~n5223;
  assign n5547 = ~n32406 & n5546;
  assign n5548 = ~n5223 & n5545;
  assign n5549 = n5119 & ~n32462;
  assign n5550 = n5123 & n5546;
  assign n5551 = n5119 & ~n32406;
  assign n5552 = ~n5111 & n5551;
  assign n5553 = ~n5223 & n5552;
  assign n5554 = ~n5119 & ~n32462;
  assign n5555 = ~n5553 & ~n5554;
  assign n5556 = ~n5549 & ~n5550;
  assign n5557 = ~n5544 & ~n32463;
  assign n5558 = ~n5542 & ~n5557;
  assign n5559 = ~n321 & ~n5558;
  assign n5560 = ~n5125 & ~n5127;
  assign n5561 = ~n5223 & n5560;
  assign n5562 = ~n32408 & ~n5561;
  assign n5563 = ~n5125 & n32408;
  assign n5564 = ~n5127 & n5563;
  assign n5565 = n32408 & n5561;
  assign n5566 = ~n5223 & n5564;
  assign n5567 = ~n5562 & ~n32464;
  assign n5568 = n321 & ~n5542;
  assign n5569 = ~n5557 & n5568;
  assign n5570 = n321 & n5558;
  assign n5571 = ~n5567 & ~n32465;
  assign n5572 = ~n5559 & ~n5571;
  assign n5573 = ~n263 & ~n5572;
  assign n5574 = n263 & ~n5559;
  assign n5575 = ~n5571 & n5574;
  assign n5576 = ~n5142 & ~n32410;
  assign n5577 = ~n5142 & ~n5223;
  assign n5578 = ~n32410 & n5577;
  assign n5579 = ~n5223 & n5576;
  assign n5580 = n5150 & ~n32466;
  assign n5581 = n5154 & n5577;
  assign n5582 = n5150 & ~n32410;
  assign n5583 = ~n5142 & n5582;
  assign n5584 = ~n5223 & n5583;
  assign n5585 = ~n5150 & ~n32466;
  assign n5586 = ~n5584 & ~n5585;
  assign n5587 = ~n5580 & ~n5581;
  assign n5588 = ~n5575 & ~n32467;
  assign n5589 = ~n5573 & ~n5588;
  assign n5590 = ~n214 & ~n5589;
  assign n5591 = ~n5156 & ~n5158;
  assign n5592 = ~n5223 & n5591;
  assign n5593 = ~n32412 & ~n5592;
  assign n5594 = ~n5156 & n32412;
  assign n5595 = ~n5158 & n5594;
  assign n5596 = n32412 & n5592;
  assign n5597 = ~n5223 & n5595;
  assign n5598 = ~n5593 & ~n32468;
  assign n5599 = n214 & ~n5573;
  assign n5600 = ~n5588 & n5599;
  assign n5601 = n214 & n5589;
  assign n5602 = ~n5598 & ~n32469;
  assign n5603 = ~n5590 & ~n5602;
  assign n5604 = ~n197 & ~n5603;
  assign n5605 = n197 & ~n5590;
  assign n5606 = ~n5602 & n5605;
  assign n5607 = ~n5173 & ~n32414;
  assign n5608 = ~n5173 & ~n5223;
  assign n5609 = ~n32414 & n5608;
  assign n5610 = ~n5223 & n5607;
  assign n5611 = n5181 & ~n32470;
  assign n5612 = n5185 & n5608;
  assign n5613 = n5181 & ~n32414;
  assign n5614 = ~n5173 & n5613;
  assign n5615 = ~n5223 & n5614;
  assign n5616 = ~n5181 & ~n32470;
  assign n5617 = ~n5615 & ~n5616;
  assign n5618 = ~n5611 & ~n5612;
  assign n5619 = ~n5606 & ~n32471;
  assign n5620 = ~n5604 & ~n5619;
  assign n5621 = ~n5187 & ~n5197;
  assign n5622 = ~n5187 & ~n5223;
  assign n5623 = ~n5197 & n5622;
  assign n5624 = ~n5223 & n5621;
  assign n5625 = n5195 & ~n32472;
  assign n5626 = n5198 & n5622;
  assign n5627 = ~n5187 & n5195;
  assign n5628 = ~n5197 & n5627;
  assign n5629 = ~n5223 & n5628;
  assign n5630 = ~n5195 & ~n32472;
  assign n5631 = ~n5629 & ~n5630;
  assign n5632 = ~n5625 & ~n5626;
  assign n5633 = ~n5199 & ~n5207;
  assign n5634 = ~n5207 & ~n5223;
  assign n5635 = ~n5199 & n5634;
  assign n5636 = ~n5223 & n5633;
  assign n5637 = ~n32418 & ~n32474;
  assign n5638 = ~n32473 & n5637;
  assign n5639 = ~n5620 & n5638;
  assign n5640 = n193 & ~n5639;
  assign n5641 = ~n5604 & n32473;
  assign n5642 = ~n5619 & n5641;
  assign n5643 = n5620 & n32473;
  assign n5644 = n5199 & ~n5634;
  assign n5645 = ~n193 & ~n5633;
  assign n5646 = ~n5644 & n5645;
  assign n5647 = ~n32475 & ~n5646;
  assign n5648 = ~n5640 & n5647;
  assign n5649 = pi74  & ~n5648;
  assign n5650 = ~pi72  & ~pi73 ;
  assign n5651 = ~pi74  & n5650;
  assign n5652 = ~n5649 & ~n5651;
  assign n5653 = ~n5223 & ~n5652;
  assign n5654 = ~n32370 & ~n32420;
  assign n5655 = ~n4830 & n5654;
  assign n5656 = ~n4849 & n5655;
  assign n5657 = ~n32372 & n5656;
  assign n5658 = n4835 & n4851;
  assign n5659 = ~n4843 & n5657;
  assign n5660 = ~n5651 & ~n32476;
  assign n5661 = ~n5221 & n5660;
  assign n5662 = ~n32418 & n5661;
  assign n5663 = ~n5215 & n5662;
  assign n5664 = n5223 & n5652;
  assign n5665 = ~n5649 & n5663;
  assign n5666 = ~pi74  & ~n5648;
  assign n5667 = pi75  & ~n5666;
  assign n5668 = ~pi75  & n5666;
  assign n5669 = n5225 & ~n5648;
  assign n5670 = ~n5667 & ~n32478;
  assign n5671 = ~n32477 & n5670;
  assign n5672 = ~n5653 & ~n5671;
  assign n5673 = ~n4851 & ~n5672;
  assign n5674 = ~n5223 & ~n5646;
  assign n5675 = ~n32475 & n5674;
  assign n5676 = ~n5640 & n5675;
  assign n5677 = ~n32478 & ~n5676;
  assign n5678 = pi76  & ~n5677;
  assign n5679 = ~pi76  & ~n5676;
  assign n5680 = ~pi76  & n5677;
  assign n5681 = ~n32478 & n5679;
  assign n5682 = ~n5678 & ~n32479;
  assign n5683 = n4851 & ~n5653;
  assign n5684 = n4851 & n5672;
  assign n5685 = ~n5671 & n5683;
  assign n5686 = ~n5682 & ~n32480;
  assign n5687 = ~n5673 & ~n5686;
  assign n5688 = ~n4461 & ~n5687;
  assign n5689 = n4461 & ~n5673;
  assign n5690 = ~n5686 & n5689;
  assign n5691 = ~n5228 & ~n32421;
  assign n5692 = ~n5648 & n5691;
  assign n5693 = n5233 & ~n5692;
  assign n5694 = ~n5233 & n5691;
  assign n5695 = ~n5233 & n5692;
  assign n5696 = ~n5648 & n5694;
  assign n5697 = ~n5693 & ~n32481;
  assign n5698 = ~n5690 & ~n5697;
  assign n5699 = ~n5688 & ~n5698;
  assign n5700 = ~n4115 & ~n5699;
  assign n5701 = ~n5248 & ~n5250;
  assign n5702 = ~n5648 & n5701;
  assign n5703 = ~n5259 & ~n5702;
  assign n5704 = ~n5250 & n5259;
  assign n5705 = ~n5248 & n5704;
  assign n5706 = n5259 & n5702;
  assign n5707 = ~n5648 & n5705;
  assign n5708 = ~n5703 & ~n32482;
  assign n5709 = n4115 & ~n5688;
  assign n5710 = n4115 & n5699;
  assign n5711 = ~n5698 & n5709;
  assign n5712 = ~n5708 & ~n32483;
  assign n5713 = ~n5700 & ~n5712;
  assign n5714 = ~n3754 & ~n5713;
  assign n5715 = n3754 & ~n5700;
  assign n5716 = ~n5712 & n5715;
  assign n5717 = ~n5262 & ~n32423;
  assign n5718 = ~n5648 & n5717;
  assign n5719 = ~n5272 & ~n5718;
  assign n5720 = ~n5262 & n5272;
  assign n5721 = ~n32423 & n5720;
  assign n5722 = n5272 & n5718;
  assign n5723 = ~n5648 & n5721;
  assign n5724 = n5272 & ~n5718;
  assign n5725 = ~n5272 & n5718;
  assign n5726 = ~n5724 & ~n5725;
  assign n5727 = ~n5719 & ~n32484;
  assign n5728 = ~n5716 & n32485;
  assign n5729 = ~n5714 & ~n5728;
  assign n5730 = ~n3444 & ~n5729;
  assign n5731 = ~n5275 & ~n5277;
  assign n5732 = ~n5648 & n5731;
  assign n5733 = ~n32426 & ~n5732;
  assign n5734 = ~n5277 & n32426;
  assign n5735 = ~n5275 & n5734;
  assign n5736 = n32426 & n5732;
  assign n5737 = ~n5648 & n5735;
  assign n5738 = ~n5733 & ~n32486;
  assign n5739 = n3444 & ~n5714;
  assign n5740 = n3444 & n5729;
  assign n5741 = ~n5728 & n5739;
  assign n5742 = ~n5738 & ~n32487;
  assign n5743 = ~n5730 & ~n5742;
  assign n5744 = ~n3116 & ~n5743;
  assign n5745 = n3116 & ~n5730;
  assign n5746 = ~n5742 & n5745;
  assign n5747 = ~n5292 & ~n32427;
  assign n5748 = ~n5648 & n5747;
  assign n5749 = ~n32429 & ~n5748;
  assign n5750 = n32429 & n5748;
  assign n5751 = ~n5292 & ~n32429;
  assign n5752 = ~n32427 & n5751;
  assign n5753 = ~n5648 & n5752;
  assign n5754 = n32429 & ~n5748;
  assign n5755 = ~n5753 & ~n5754;
  assign n5756 = ~n5749 & ~n5750;
  assign n5757 = ~n5746 & ~n32488;
  assign n5758 = ~n5744 & ~n5757;
  assign n5759 = ~n2833 & ~n5758;
  assign n5760 = ~n5309 & ~n5311;
  assign n5761 = ~n5648 & n5760;
  assign n5762 = ~n32431 & ~n5761;
  assign n5763 = ~n5311 & n32431;
  assign n5764 = ~n5309 & n5763;
  assign n5765 = n32431 & n5761;
  assign n5766 = ~n5648 & n5764;
  assign n5767 = ~n5762 & ~n32489;
  assign n5768 = n2833 & ~n5744;
  assign n5769 = n2833 & n5758;
  assign n5770 = ~n5757 & n5768;
  assign n5771 = ~n5767 & ~n32490;
  assign n5772 = ~n5759 & ~n5771;
  assign n5773 = ~n2536 & ~n5772;
  assign n5774 = n2536 & ~n5759;
  assign n5775 = ~n5771 & n5774;
  assign n5776 = ~n5326 & ~n32432;
  assign n5777 = ~n5648 & n5776;
  assign n5778 = ~n32433 & n5777;
  assign n5779 = n32433 & ~n5777;
  assign n5780 = ~n5326 & n32433;
  assign n5781 = ~n32432 & n5780;
  assign n5782 = ~n5648 & n5781;
  assign n5783 = ~n32433 & ~n5777;
  assign n5784 = ~n5782 & ~n5783;
  assign n5785 = ~n5778 & ~n5779;
  assign n5786 = ~n5775 & ~n32491;
  assign n5787 = ~n5773 & ~n5786;
  assign n5788 = ~n2283 & ~n5787;
  assign n5789 = ~n5342 & ~n5344;
  assign n5790 = ~n5648 & n5789;
  assign n5791 = ~n32435 & ~n5790;
  assign n5792 = ~n5344 & n32435;
  assign n5793 = ~n5342 & n5792;
  assign n5794 = n32435 & n5790;
  assign n5795 = ~n5648 & n5793;
  assign n5796 = ~n5791 & ~n32492;
  assign n5797 = n2283 & ~n5773;
  assign n5798 = n2283 & n5787;
  assign n5799 = ~n5786 & n5797;
  assign n5800 = ~n5796 & ~n32493;
  assign n5801 = ~n5788 & ~n5800;
  assign n5802 = ~n2021 & ~n5801;
  assign n5803 = n2021 & ~n5788;
  assign n5804 = ~n5800 & n5803;
  assign n5805 = ~n5359 & ~n32436;
  assign n5806 = ~n5648 & n5805;
  assign n5807 = ~n32437 & n5806;
  assign n5808 = n32437 & ~n5806;
  assign n5809 = ~n32437 & ~n5806;
  assign n5810 = ~n5359 & n32437;
  assign n5811 = ~n32436 & n5810;
  assign n5812 = n32437 & n5806;
  assign n5813 = ~n5648 & n5811;
  assign n5814 = ~n5809 & ~n32494;
  assign n5815 = ~n5807 & ~n5808;
  assign n5816 = ~n5804 & ~n32495;
  assign n5817 = ~n5802 & ~n5816;
  assign n5818 = ~n1796 & ~n5817;
  assign n5819 = ~n5375 & ~n5377;
  assign n5820 = ~n5648 & n5819;
  assign n5821 = ~n32439 & ~n5820;
  assign n5822 = ~n5377 & n32439;
  assign n5823 = ~n5375 & n5822;
  assign n5824 = n32439 & n5820;
  assign n5825 = ~n5648 & n5823;
  assign n5826 = ~n5821 & ~n32496;
  assign n5827 = n1796 & ~n5802;
  assign n5828 = n1796 & n5817;
  assign n5829 = ~n5816 & n5827;
  assign n5830 = ~n5826 & ~n32497;
  assign n5831 = ~n5818 & ~n5830;
  assign n5832 = ~n1567 & ~n5831;
  assign n5833 = n1567 & ~n5818;
  assign n5834 = ~n5830 & n5833;
  assign n5835 = ~n5392 & ~n32440;
  assign n5836 = ~n5392 & ~n5648;
  assign n5837 = ~n32440 & n5836;
  assign n5838 = ~n5648 & n5835;
  assign n5839 = n32442 & ~n32498;
  assign n5840 = n5407 & n5836;
  assign n5841 = ~n32442 & n32498;
  assign n5842 = ~n5392 & n32442;
  assign n5843 = ~n32440 & n5842;
  assign n5844 = ~n5648 & n5843;
  assign n5845 = ~n32442 & ~n32498;
  assign n5846 = ~n5844 & ~n5845;
  assign n5847 = ~n5839 & ~n32499;
  assign n5848 = ~n5834 & ~n32500;
  assign n5849 = ~n5832 & ~n5848;
  assign n5850 = ~n1374 & ~n5849;
  assign n5851 = ~n5409 & ~n5411;
  assign n5852 = ~n5648 & n5851;
  assign n5853 = ~n32444 & ~n5852;
  assign n5854 = ~n5411 & n32444;
  assign n5855 = ~n5409 & n5854;
  assign n5856 = n32444 & n5852;
  assign n5857 = ~n5648 & n5855;
  assign n5858 = ~n5853 & ~n32501;
  assign n5859 = n1374 & ~n5832;
  assign n5860 = n1374 & n5849;
  assign n5861 = ~n5848 & n5859;
  assign n5862 = ~n5858 & ~n32502;
  assign n5863 = ~n5850 & ~n5862;
  assign n5864 = ~n1179 & ~n5863;
  assign n5865 = ~n5426 & ~n32445;
  assign n5866 = ~n5648 & n5865;
  assign n5867 = ~n32448 & ~n5866;
  assign n5868 = ~n5426 & n32448;
  assign n5869 = ~n32445 & n5868;
  assign n5870 = n32448 & n5866;
  assign n5871 = ~n5648 & n5869;
  assign n5872 = ~n5867 & ~n32503;
  assign n5873 = n1179 & ~n5850;
  assign n5874 = ~n5862 & n5873;
  assign n5875 = ~n5872 & ~n5874;
  assign n5876 = ~n5864 & ~n5875;
  assign n5877 = ~n1016 & ~n5876;
  assign n5878 = ~n5445 & ~n5447;
  assign n5879 = ~n5648 & n5878;
  assign n5880 = ~n32450 & ~n5879;
  assign n5881 = ~n5447 & n32450;
  assign n5882 = ~n5445 & n5881;
  assign n5883 = n32450 & n5879;
  assign n5884 = ~n5648 & n5882;
  assign n5885 = ~n5880 & ~n32504;
  assign n5886 = n1016 & ~n5864;
  assign n5887 = n1016 & n5876;
  assign n5888 = ~n5875 & n5886;
  assign n5889 = ~n5885 & ~n32505;
  assign n5890 = ~n5877 & ~n5889;
  assign n5891 = ~n855 & ~n5890;
  assign n5892 = n855 & ~n5877;
  assign n5893 = ~n5889 & n5892;
  assign n5894 = ~n5462 & ~n32452;
  assign n5895 = ~n5462 & ~n5648;
  assign n5896 = ~n32452 & n5895;
  assign n5897 = ~n5648 & n5894;
  assign n5898 = n5470 & ~n32506;
  assign n5899 = n5474 & n5895;
  assign n5900 = ~n5462 & n5470;
  assign n5901 = ~n32452 & n5900;
  assign n5902 = ~n5648 & n5901;
  assign n5903 = ~n5470 & ~n32506;
  assign n5904 = ~n5902 & ~n5903;
  assign n5905 = ~n5898 & ~n5899;
  assign n5906 = ~n5893 & ~n32507;
  assign n5907 = ~n5891 & ~n5906;
  assign n5908 = ~n720 & ~n5907;
  assign n5909 = ~n5476 & ~n5478;
  assign n5910 = ~n5648 & n5909;
  assign n5911 = ~n32454 & ~n5910;
  assign n5912 = ~n5478 & n32454;
  assign n5913 = ~n5476 & n5912;
  assign n5914 = n32454 & n5910;
  assign n5915 = ~n5648 & n5913;
  assign n5916 = ~n5911 & ~n32508;
  assign n5917 = n720 & ~n5891;
  assign n5918 = n720 & n5907;
  assign n5919 = ~n5906 & n5917;
  assign n5920 = ~n5916 & ~n32509;
  assign n5921 = ~n5908 & ~n5920;
  assign n5922 = ~n592 & ~n5921;
  assign n5923 = ~n5493 & ~n32455;
  assign n5924 = ~n5648 & n5923;
  assign n5925 = ~n32457 & ~n5924;
  assign n5926 = ~n5493 & n32457;
  assign n5927 = ~n32455 & n5926;
  assign n5928 = n32457 & n5924;
  assign n5929 = ~n5648 & n5927;
  assign n5930 = ~n5925 & ~n32510;
  assign n5931 = n592 & ~n5908;
  assign n5932 = ~n5920 & n5931;
  assign n5933 = ~n5930 & ~n5932;
  assign n5934 = ~n5922 & ~n5933;
  assign n5935 = ~n487 & ~n5934;
  assign n5936 = ~n5511 & ~n5513;
  assign n5937 = ~n5648 & n5936;
  assign n5938 = ~n32459 & ~n5937;
  assign n5939 = ~n5513 & n32459;
  assign n5940 = ~n5511 & n5939;
  assign n5941 = n32459 & n5937;
  assign n5942 = ~n5648 & n5940;
  assign n5943 = ~n5938 & ~n32511;
  assign n5944 = n487 & ~n5922;
  assign n5945 = n487 & n5934;
  assign n5946 = ~n5933 & n5944;
  assign n5947 = ~n5943 & ~n32512;
  assign n5948 = ~n5935 & ~n5947;
  assign n5949 = ~n393 & ~n5948;
  assign n5950 = n393 & ~n5935;
  assign n5951 = ~n5947 & n5950;
  assign n5952 = ~n5528 & ~n32461;
  assign n5953 = ~n5528 & ~n5648;
  assign n5954 = ~n32461 & n5953;
  assign n5955 = ~n5648 & n5952;
  assign n5956 = n5536 & ~n32513;
  assign n5957 = n5540 & n5953;
  assign n5958 = ~n5528 & n5536;
  assign n5959 = ~n32461 & n5958;
  assign n5960 = ~n5648 & n5959;
  assign n5961 = ~n5536 & ~n32513;
  assign n5962 = ~n5960 & ~n5961;
  assign n5963 = ~n5956 & ~n5957;
  assign n5964 = ~n5951 & ~n32514;
  assign n5965 = ~n5949 & ~n5964;
  assign n5966 = ~n321 & ~n5965;
  assign n5967 = ~n5542 & ~n5544;
  assign n5968 = ~n5648 & n5967;
  assign n5969 = ~n32463 & ~n5968;
  assign n5970 = ~n5544 & n32463;
  assign n5971 = ~n5542 & n5970;
  assign n5972 = n32463 & n5968;
  assign n5973 = ~n5648 & n5971;
  assign n5974 = ~n5969 & ~n32515;
  assign n5975 = n321 & ~n5949;
  assign n5976 = n321 & n5965;
  assign n5977 = ~n5964 & n5975;
  assign n5978 = ~n5974 & ~n32516;
  assign n5979 = ~n5966 & ~n5978;
  assign n5980 = ~n263 & ~n5979;
  assign n5981 = n263 & ~n5966;
  assign n5982 = ~n5978 & n5981;
  assign n5983 = ~n5559 & ~n32465;
  assign n5984 = ~n5559 & ~n5648;
  assign n5985 = ~n32465 & n5984;
  assign n5986 = ~n5648 & n5983;
  assign n5987 = n5567 & ~n32517;
  assign n5988 = n5571 & n5984;
  assign n5989 = ~n5559 & n5567;
  assign n5990 = ~n32465 & n5989;
  assign n5991 = ~n5648 & n5990;
  assign n5992 = ~n5567 & ~n32517;
  assign n5993 = ~n5991 & ~n5992;
  assign n5994 = ~n5987 & ~n5988;
  assign n5995 = ~n5982 & ~n32518;
  assign n5996 = ~n5980 & ~n5995;
  assign n5997 = ~n214 & ~n5996;
  assign n5998 = ~n5573 & ~n5575;
  assign n5999 = ~n5648 & n5998;
  assign n6000 = ~n32467 & ~n5999;
  assign n6001 = ~n5575 & n32467;
  assign n6002 = ~n5573 & n6001;
  assign n6003 = n32467 & n5999;
  assign n6004 = ~n5648 & n6002;
  assign n6005 = ~n6000 & ~n32519;
  assign n6006 = n214 & ~n5980;
  assign n6007 = n214 & n5996;
  assign n6008 = ~n5995 & n6006;
  assign n6009 = ~n6005 & ~n32520;
  assign n6010 = ~n5997 & ~n6009;
  assign n6011 = ~n197 & ~n6010;
  assign n6012 = n197 & ~n5997;
  assign n6013 = ~n6009 & n6012;
  assign n6014 = ~n5590 & ~n32469;
  assign n6015 = ~n5590 & ~n5648;
  assign n6016 = ~n32469 & n6015;
  assign n6017 = ~n5648 & n6014;
  assign n6018 = n5598 & ~n32521;
  assign n6019 = n5602 & n6015;
  assign n6020 = ~n5590 & n5598;
  assign n6021 = ~n32469 & n6020;
  assign n6022 = ~n5648 & n6021;
  assign n6023 = ~n5598 & ~n32521;
  assign n6024 = ~n6022 & ~n6023;
  assign n6025 = ~n6018 & ~n6019;
  assign n6026 = ~n6013 & ~n32522;
  assign n6027 = ~n6011 & ~n6026;
  assign n6028 = ~n5604 & ~n5606;
  assign n6029 = ~n5648 & n6028;
  assign n6030 = ~n32471 & ~n6029;
  assign n6031 = ~n5606 & n32471;
  assign n6032 = ~n5604 & n6031;
  assign n6033 = n32471 & n6029;
  assign n6034 = ~n5648 & n6032;
  assign n6035 = ~n6030 & ~n32523;
  assign n6036 = ~n5620 & ~n32473;
  assign n6037 = ~n32473 & ~n5648;
  assign n6038 = ~n5620 & n6037;
  assign n6039 = ~n5648 & n6036;
  assign n6040 = ~n32475 & ~n32524;
  assign n6041 = ~n6035 & n6040;
  assign n6042 = ~n6027 & n6041;
  assign n6043 = n193 & ~n6042;
  assign n6044 = ~n6011 & n6035;
  assign n6045 = n6027 & n6035;
  assign n6046 = ~n6026 & n6044;
  assign n6047 = n5620 & ~n6037;
  assign n6048 = ~n193 & ~n6036;
  assign n6049 = ~n6047 & n6048;
  assign n6050 = ~n32525 & ~n6049;
  assign n6051 = ~n6043 & n6050;
  assign n6052 = pi72  & ~n6051;
  assign n6053 = ~pi70  & ~pi71 ;
  assign n6054 = ~pi72  & n6053;
  assign n6055 = ~n6052 & ~n6054;
  assign n6056 = ~n5648 & ~n6055;
  assign n6057 = ~pi72  & ~n6051;
  assign n6058 = pi73  & ~n6057;
  assign n6059 = ~pi73  & n6057;
  assign n6060 = n5650 & ~n6051;
  assign n6061 = ~n6058 & ~n32526;
  assign n6062 = ~n32416 & ~n32476;
  assign n6063 = ~n5202 & n6062;
  assign n6064 = ~n5221 & n6063;
  assign n6065 = ~n32418 & n6064;
  assign n6066 = n5207 & n5223;
  assign n6067 = ~n5215 & n6065;
  assign n6068 = ~n6054 & ~n32527;
  assign n6069 = ~n5646 & n6068;
  assign n6070 = ~n32475 & n6069;
  assign n6071 = ~n5640 & n6070;
  assign n6072 = n5648 & n6055;
  assign n6073 = ~n6052 & n6071;
  assign n6074 = n6061 & ~n32528;
  assign n6075 = ~n6056 & ~n6074;
  assign n6076 = ~n5223 & ~n6075;
  assign n6077 = n5223 & ~n6056;
  assign n6078 = ~n6074 & n6077;
  assign n6079 = ~n5648 & ~n6049;
  assign n6080 = ~n32525 & n6079;
  assign n6081 = ~n6043 & n6080;
  assign n6082 = ~n32526 & ~n6081;
  assign n6083 = pi74  & ~n6082;
  assign n6084 = ~pi74  & ~n6081;
  assign n6085 = ~pi74  & n6082;
  assign n6086 = ~n32526 & n6084;
  assign n6087 = ~n6083 & ~n32529;
  assign n6088 = ~n6078 & ~n6087;
  assign n6089 = ~n6076 & ~n6088;
  assign n6090 = ~n4851 & ~n6089;
  assign n6091 = n4851 & ~n6076;
  assign n6092 = ~n6088 & n6091;
  assign n6093 = n4851 & n6089;
  assign n6094 = ~n5653 & ~n32477;
  assign n6095 = ~n6051 & n6094;
  assign n6096 = n5670 & ~n6095;
  assign n6097 = ~n5670 & n6094;
  assign n6098 = ~n5670 & n6095;
  assign n6099 = ~n6051 & n6097;
  assign n6100 = ~n6096 & ~n32531;
  assign n6101 = ~n32530 & ~n6100;
  assign n6102 = ~n6090 & ~n6101;
  assign n6103 = ~n4461 & ~n6102;
  assign n6104 = n4461 & ~n6090;
  assign n6105 = ~n6101 & n6104;
  assign n6106 = ~n5673 & ~n32480;
  assign n6107 = ~n5673 & ~n6051;
  assign n6108 = ~n32480 & n6107;
  assign n6109 = ~n6051 & n6106;
  assign n6110 = n5682 & ~n32532;
  assign n6111 = n5686 & n6107;
  assign n6112 = n5682 & ~n32480;
  assign n6113 = ~n5673 & n6112;
  assign n6114 = ~n6051 & n6113;
  assign n6115 = ~n5682 & ~n32532;
  assign n6116 = ~n6114 & ~n6115;
  assign n6117 = ~n6110 & ~n6111;
  assign n6118 = ~n6105 & ~n32533;
  assign n6119 = ~n6103 & ~n6118;
  assign n6120 = ~n4115 & ~n6119;
  assign n6121 = n4115 & ~n6103;
  assign n6122 = ~n6118 & n6121;
  assign n6123 = n4115 & n6119;
  assign n6124 = ~n5688 & ~n5690;
  assign n6125 = ~n6051 & n6124;
  assign n6126 = ~n5697 & ~n6125;
  assign n6127 = ~n5688 & n5697;
  assign n6128 = ~n5690 & n6127;
  assign n6129 = n5697 & n6125;
  assign n6130 = ~n6051 & n6128;
  assign n6131 = n5697 & ~n6125;
  assign n6132 = ~n5697 & n6125;
  assign n6133 = ~n6131 & ~n6132;
  assign n6134 = ~n6126 & ~n32535;
  assign n6135 = ~n32534 & n32536;
  assign n6136 = ~n6120 & ~n6135;
  assign n6137 = ~n3754 & ~n6136;
  assign n6138 = n3754 & ~n6120;
  assign n6139 = ~n6135 & n6138;
  assign n6140 = ~n5700 & ~n32483;
  assign n6141 = ~n5700 & ~n6051;
  assign n6142 = ~n32483 & n6141;
  assign n6143 = ~n6051 & n6140;
  assign n6144 = n5708 & ~n32537;
  assign n6145 = n5712 & n6141;
  assign n6146 = n5708 & ~n32483;
  assign n6147 = ~n5700 & n6146;
  assign n6148 = ~n6051 & n6147;
  assign n6149 = ~n5708 & ~n32537;
  assign n6150 = ~n6148 & ~n6149;
  assign n6151 = ~n6144 & ~n6145;
  assign n6152 = ~n6139 & ~n32538;
  assign n6153 = ~n6137 & ~n6152;
  assign n6154 = ~n3444 & ~n6153;
  assign n6155 = n3444 & ~n6137;
  assign n6156 = ~n6152 & n6155;
  assign n6157 = n3444 & n6153;
  assign n6158 = ~n5714 & ~n5716;
  assign n6159 = ~n6051 & n6158;
  assign n6160 = ~n32485 & ~n6159;
  assign n6161 = n32485 & n6159;
  assign n6162 = ~n5714 & ~n32485;
  assign n6163 = ~n5716 & n6162;
  assign n6164 = ~n6051 & n6163;
  assign n6165 = n32485 & ~n6159;
  assign n6166 = ~n6164 & ~n6165;
  assign n6167 = ~n6160 & ~n6161;
  assign n6168 = ~n32539 & ~n32540;
  assign n6169 = ~n6154 & ~n6168;
  assign n6170 = ~n3116 & ~n6169;
  assign n6171 = n3116 & ~n6154;
  assign n6172 = ~n6168 & n6171;
  assign n6173 = ~n5730 & ~n32487;
  assign n6174 = ~n5730 & ~n6051;
  assign n6175 = ~n32487 & n6174;
  assign n6176 = ~n6051 & n6173;
  assign n6177 = n5738 & ~n32541;
  assign n6178 = n5742 & n6174;
  assign n6179 = n5738 & ~n32487;
  assign n6180 = ~n5730 & n6179;
  assign n6181 = ~n6051 & n6180;
  assign n6182 = ~n5738 & ~n32541;
  assign n6183 = ~n6181 & ~n6182;
  assign n6184 = ~n6177 & ~n6178;
  assign n6185 = ~n6172 & ~n32542;
  assign n6186 = ~n6170 & ~n6185;
  assign n6187 = ~n2833 & ~n6186;
  assign n6188 = n2833 & ~n6170;
  assign n6189 = ~n6185 & n6188;
  assign n6190 = n2833 & n6186;
  assign n6191 = ~n5744 & ~n5746;
  assign n6192 = ~n6051 & n6191;
  assign n6193 = ~n32488 & n6192;
  assign n6194 = n32488 & ~n6192;
  assign n6195 = ~n5744 & n32488;
  assign n6196 = ~n5746 & n6195;
  assign n6197 = ~n6051 & n6196;
  assign n6198 = ~n32488 & ~n6192;
  assign n6199 = ~n6197 & ~n6198;
  assign n6200 = ~n6193 & ~n6194;
  assign n6201 = ~n32543 & ~n32544;
  assign n6202 = ~n6187 & ~n6201;
  assign n6203 = ~n2536 & ~n6202;
  assign n6204 = n2536 & ~n6187;
  assign n6205 = ~n6201 & n6204;
  assign n6206 = ~n5759 & ~n32490;
  assign n6207 = ~n5759 & ~n6051;
  assign n6208 = ~n32490 & n6207;
  assign n6209 = ~n6051 & n6206;
  assign n6210 = n5767 & ~n32545;
  assign n6211 = n5771 & n6207;
  assign n6212 = n5767 & ~n32490;
  assign n6213 = ~n5759 & n6212;
  assign n6214 = ~n6051 & n6213;
  assign n6215 = ~n5767 & ~n32545;
  assign n6216 = ~n6214 & ~n6215;
  assign n6217 = ~n6210 & ~n6211;
  assign n6218 = ~n6205 & ~n32546;
  assign n6219 = ~n6203 & ~n6218;
  assign n6220 = ~n2283 & ~n6219;
  assign n6221 = n2283 & ~n6203;
  assign n6222 = ~n6218 & n6221;
  assign n6223 = n2283 & n6219;
  assign n6224 = ~n5773 & ~n5775;
  assign n6225 = ~n6051 & n6224;
  assign n6226 = ~n32491 & n6225;
  assign n6227 = n32491 & ~n6225;
  assign n6228 = ~n32491 & ~n6225;
  assign n6229 = ~n5773 & n32491;
  assign n6230 = ~n5775 & n6229;
  assign n6231 = n32491 & n6225;
  assign n6232 = ~n6051 & n6230;
  assign n6233 = ~n6228 & ~n32548;
  assign n6234 = ~n6226 & ~n6227;
  assign n6235 = ~n32547 & ~n32549;
  assign n6236 = ~n6220 & ~n6235;
  assign n6237 = ~n2021 & ~n6236;
  assign n6238 = n2021 & ~n6220;
  assign n6239 = ~n6235 & n6238;
  assign n6240 = ~n5788 & ~n32493;
  assign n6241 = ~n5788 & ~n6051;
  assign n6242 = ~n32493 & n6241;
  assign n6243 = ~n6051 & n6240;
  assign n6244 = n5796 & ~n32550;
  assign n6245 = n5800 & n6241;
  assign n6246 = n5796 & ~n32493;
  assign n6247 = ~n5788 & n6246;
  assign n6248 = ~n6051 & n6247;
  assign n6249 = ~n5796 & ~n32550;
  assign n6250 = ~n6248 & ~n6249;
  assign n6251 = ~n6244 & ~n6245;
  assign n6252 = ~n6239 & ~n32551;
  assign n6253 = ~n6237 & ~n6252;
  assign n6254 = ~n1796 & ~n6253;
  assign n6255 = n1796 & ~n6237;
  assign n6256 = ~n6252 & n6255;
  assign n6257 = n1796 & n6253;
  assign n6258 = ~n5802 & ~n5804;
  assign n6259 = ~n5802 & ~n6051;
  assign n6260 = ~n5804 & n6259;
  assign n6261 = ~n6051 & n6258;
  assign n6262 = n32495 & ~n32553;
  assign n6263 = n5816 & n6259;
  assign n6264 = ~n32495 & n32553;
  assign n6265 = ~n5802 & n32495;
  assign n6266 = ~n5804 & n6265;
  assign n6267 = ~n6051 & n6266;
  assign n6268 = ~n32495 & ~n32553;
  assign n6269 = ~n6267 & ~n6268;
  assign n6270 = ~n6262 & ~n32554;
  assign n6271 = ~n32552 & ~n32555;
  assign n6272 = ~n6254 & ~n6271;
  assign n6273 = ~n1567 & ~n6272;
  assign n6274 = n1567 & ~n6254;
  assign n6275 = ~n6271 & n6274;
  assign n6276 = ~n5818 & ~n32497;
  assign n6277 = ~n5818 & ~n6051;
  assign n6278 = ~n32497 & n6277;
  assign n6279 = ~n6051 & n6276;
  assign n6280 = n5826 & ~n32556;
  assign n6281 = n5830 & n6277;
  assign n6282 = n5826 & ~n32497;
  assign n6283 = ~n5818 & n6282;
  assign n6284 = ~n6051 & n6283;
  assign n6285 = ~n5826 & ~n32556;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = ~n6280 & ~n6281;
  assign n6288 = ~n6275 & ~n32557;
  assign n6289 = ~n6273 & ~n6288;
  assign n6290 = ~n1374 & ~n6289;
  assign n6291 = ~n5832 & ~n5834;
  assign n6292 = ~n6051 & n6291;
  assign n6293 = ~n32500 & ~n6292;
  assign n6294 = ~n5832 & n32500;
  assign n6295 = ~n5834 & n6294;
  assign n6296 = n32500 & n6292;
  assign n6297 = ~n6051 & n6295;
  assign n6298 = ~n6293 & ~n32558;
  assign n6299 = n1374 & ~n6273;
  assign n6300 = ~n6288 & n6299;
  assign n6301 = n1374 & n6289;
  assign n6302 = ~n6298 & ~n32559;
  assign n6303 = ~n6290 & ~n6302;
  assign n6304 = ~n1179 & ~n6303;
  assign n6305 = n1179 & ~n6290;
  assign n6306 = ~n6302 & n6305;
  assign n6307 = ~n5850 & ~n32502;
  assign n6308 = ~n5850 & ~n6051;
  assign n6309 = ~n32502 & n6308;
  assign n6310 = ~n6051 & n6307;
  assign n6311 = n5858 & ~n32560;
  assign n6312 = n5862 & n6308;
  assign n6313 = n5858 & ~n32502;
  assign n6314 = ~n5850 & n6313;
  assign n6315 = ~n6051 & n6314;
  assign n6316 = ~n5858 & ~n32560;
  assign n6317 = ~n6315 & ~n6316;
  assign n6318 = ~n6311 & ~n6312;
  assign n6319 = ~n6306 & ~n32561;
  assign n6320 = ~n6304 & ~n6319;
  assign n6321 = ~n1016 & ~n6320;
  assign n6322 = n1016 & ~n6304;
  assign n6323 = ~n6319 & n6322;
  assign n6324 = n1016 & n6320;
  assign n6325 = ~n5864 & ~n5874;
  assign n6326 = ~n5864 & ~n6051;
  assign n6327 = ~n5874 & n6326;
  assign n6328 = ~n6051 & n6325;
  assign n6329 = n5872 & ~n32563;
  assign n6330 = n5875 & n6326;
  assign n6331 = ~n5864 & n5872;
  assign n6332 = ~n5874 & n6331;
  assign n6333 = ~n6051 & n6332;
  assign n6334 = ~n5872 & ~n32563;
  assign n6335 = ~n6333 & ~n6334;
  assign n6336 = ~n6329 & ~n6330;
  assign n6337 = ~n32562 & ~n32564;
  assign n6338 = ~n6321 & ~n6337;
  assign n6339 = ~n855 & ~n6338;
  assign n6340 = n855 & ~n6321;
  assign n6341 = ~n6337 & n6340;
  assign n6342 = ~n5877 & ~n32505;
  assign n6343 = ~n5877 & ~n6051;
  assign n6344 = ~n32505 & n6343;
  assign n6345 = ~n6051 & n6342;
  assign n6346 = n5885 & ~n32565;
  assign n6347 = n5889 & n6343;
  assign n6348 = n5885 & ~n32505;
  assign n6349 = ~n5877 & n6348;
  assign n6350 = ~n6051 & n6349;
  assign n6351 = ~n5885 & ~n32565;
  assign n6352 = ~n6350 & ~n6351;
  assign n6353 = ~n6346 & ~n6347;
  assign n6354 = ~n6341 & ~n32566;
  assign n6355 = ~n6339 & ~n6354;
  assign n6356 = ~n720 & ~n6355;
  assign n6357 = ~n5891 & ~n5893;
  assign n6358 = ~n6051 & n6357;
  assign n6359 = ~n32507 & ~n6358;
  assign n6360 = ~n5891 & n32507;
  assign n6361 = ~n5893 & n6360;
  assign n6362 = n32507 & n6358;
  assign n6363 = ~n6051 & n6361;
  assign n6364 = ~n6359 & ~n32567;
  assign n6365 = n720 & ~n6339;
  assign n6366 = ~n6354 & n6365;
  assign n6367 = n720 & n6355;
  assign n6368 = ~n6364 & ~n32568;
  assign n6369 = ~n6356 & ~n6368;
  assign n6370 = ~n592 & ~n6369;
  assign n6371 = n592 & ~n6356;
  assign n6372 = ~n6368 & n6371;
  assign n6373 = ~n5908 & ~n32509;
  assign n6374 = ~n5908 & ~n6051;
  assign n6375 = ~n32509 & n6374;
  assign n6376 = ~n6051 & n6373;
  assign n6377 = n5916 & ~n32569;
  assign n6378 = n5920 & n6374;
  assign n6379 = n5916 & ~n32509;
  assign n6380 = ~n5908 & n6379;
  assign n6381 = ~n6051 & n6380;
  assign n6382 = ~n5916 & ~n32569;
  assign n6383 = ~n6381 & ~n6382;
  assign n6384 = ~n6377 & ~n6378;
  assign n6385 = ~n6372 & ~n32570;
  assign n6386 = ~n6370 & ~n6385;
  assign n6387 = ~n487 & ~n6386;
  assign n6388 = n487 & ~n6370;
  assign n6389 = ~n6385 & n6388;
  assign n6390 = n487 & n6386;
  assign n6391 = ~n5922 & ~n5932;
  assign n6392 = ~n5922 & ~n6051;
  assign n6393 = ~n5932 & n6392;
  assign n6394 = ~n6051 & n6391;
  assign n6395 = n5930 & ~n32572;
  assign n6396 = n5933 & n6392;
  assign n6397 = ~n5922 & n5930;
  assign n6398 = ~n5932 & n6397;
  assign n6399 = ~n6051 & n6398;
  assign n6400 = ~n5930 & ~n32572;
  assign n6401 = ~n6399 & ~n6400;
  assign n6402 = ~n6395 & ~n6396;
  assign n6403 = ~n32571 & ~n32573;
  assign n6404 = ~n6387 & ~n6403;
  assign n6405 = ~n393 & ~n6404;
  assign n6406 = n393 & ~n6387;
  assign n6407 = ~n6403 & n6406;
  assign n6408 = ~n5935 & ~n32512;
  assign n6409 = ~n5935 & ~n6051;
  assign n6410 = ~n32512 & n6409;
  assign n6411 = ~n6051 & n6408;
  assign n6412 = n5943 & ~n32574;
  assign n6413 = n5947 & n6409;
  assign n6414 = n5943 & ~n32512;
  assign n6415 = ~n5935 & n6414;
  assign n6416 = ~n6051 & n6415;
  assign n6417 = ~n5943 & ~n32574;
  assign n6418 = ~n6416 & ~n6417;
  assign n6419 = ~n6412 & ~n6413;
  assign n6420 = ~n6407 & ~n32575;
  assign n6421 = ~n6405 & ~n6420;
  assign n6422 = ~n321 & ~n6421;
  assign n6423 = ~n5949 & ~n5951;
  assign n6424 = ~n6051 & n6423;
  assign n6425 = ~n32514 & ~n6424;
  assign n6426 = ~n5949 & n32514;
  assign n6427 = ~n5951 & n6426;
  assign n6428 = n32514 & n6424;
  assign n6429 = ~n6051 & n6427;
  assign n6430 = ~n6425 & ~n32576;
  assign n6431 = n321 & ~n6405;
  assign n6432 = ~n6420 & n6431;
  assign n6433 = n321 & n6421;
  assign n6434 = ~n6430 & ~n32577;
  assign n6435 = ~n6422 & ~n6434;
  assign n6436 = ~n263 & ~n6435;
  assign n6437 = n263 & ~n6422;
  assign n6438 = ~n6434 & n6437;
  assign n6439 = ~n5966 & ~n32516;
  assign n6440 = ~n5966 & ~n6051;
  assign n6441 = ~n32516 & n6440;
  assign n6442 = ~n6051 & n6439;
  assign n6443 = n5974 & ~n32578;
  assign n6444 = n5978 & n6440;
  assign n6445 = n5974 & ~n32516;
  assign n6446 = ~n5966 & n6445;
  assign n6447 = ~n6051 & n6446;
  assign n6448 = ~n5974 & ~n32578;
  assign n6449 = ~n6447 & ~n6448;
  assign n6450 = ~n6443 & ~n6444;
  assign n6451 = ~n6438 & ~n32579;
  assign n6452 = ~n6436 & ~n6451;
  assign n6453 = ~n214 & ~n6452;
  assign n6454 = ~n5980 & ~n5982;
  assign n6455 = ~n6051 & n6454;
  assign n6456 = ~n32518 & ~n6455;
  assign n6457 = ~n5980 & n32518;
  assign n6458 = ~n5982 & n6457;
  assign n6459 = n32518 & n6455;
  assign n6460 = ~n6051 & n6458;
  assign n6461 = ~n6456 & ~n32580;
  assign n6462 = n214 & ~n6436;
  assign n6463 = ~n6451 & n6462;
  assign n6464 = n214 & n6452;
  assign n6465 = ~n6461 & ~n32581;
  assign n6466 = ~n6453 & ~n6465;
  assign n6467 = ~n197 & ~n6466;
  assign n6468 = n197 & ~n6453;
  assign n6469 = ~n6465 & n6468;
  assign n6470 = ~n5997 & ~n32520;
  assign n6471 = ~n5997 & ~n6051;
  assign n6472 = ~n32520 & n6471;
  assign n6473 = ~n6051 & n6470;
  assign n6474 = n6005 & ~n32582;
  assign n6475 = n6009 & n6471;
  assign n6476 = n6005 & ~n32520;
  assign n6477 = ~n5997 & n6476;
  assign n6478 = ~n6051 & n6477;
  assign n6479 = ~n6005 & ~n32582;
  assign n6480 = ~n6478 & ~n6479;
  assign n6481 = ~n6474 & ~n6475;
  assign n6482 = ~n6469 & ~n32583;
  assign n6483 = ~n6467 & ~n6482;
  assign n6484 = ~n6011 & ~n6013;
  assign n6485 = ~n6051 & n6484;
  assign n6486 = ~n32522 & ~n6485;
  assign n6487 = ~n6011 & n32522;
  assign n6488 = ~n6013 & n6487;
  assign n6489 = n32522 & n6485;
  assign n6490 = ~n6051 & n6488;
  assign n6491 = ~n6486 & ~n32584;
  assign n6492 = ~n6027 & ~n6035;
  assign n6493 = ~n6035 & ~n6051;
  assign n6494 = ~n6027 & n6493;
  assign n6495 = ~n6051 & n6492;
  assign n6496 = ~n32525 & ~n32585;
  assign n6497 = ~n6491 & n6496;
  assign n6498 = ~n6483 & n6497;
  assign n6499 = n193 & ~n6498;
  assign n6500 = ~n6467 & n6491;
  assign n6501 = ~n6482 & n6500;
  assign n6502 = n6483 & n6491;
  assign n6503 = n6027 & ~n6493;
  assign n6504 = ~n193 & ~n6492;
  assign n6505 = ~n6503 & n6504;
  assign n6506 = ~n32586 & ~n6505;
  assign n6507 = ~n6499 & n6506;
  assign n6508 = pi70  & ~n6507;
  assign n6509 = ~pi68  & ~pi69 ;
  assign n6510 = ~pi70  & n6509;
  assign n6511 = ~n6508 & ~n6510;
  assign n6512 = ~n6051 & ~n6511;
  assign n6513 = ~n5629 & ~n32527;
  assign n6514 = ~n5630 & n6513;
  assign n6515 = ~n5646 & n6514;
  assign n6516 = ~n32475 & n6515;
  assign n6517 = n32473 & n5648;
  assign n6518 = ~n5640 & n6516;
  assign n6519 = ~n6510 & ~n32587;
  assign n6520 = ~n6049 & n6519;
  assign n6521 = ~n32525 & n6520;
  assign n6522 = ~n6043 & n6521;
  assign n6523 = n6051 & n6511;
  assign n6524 = ~n6508 & n6522;
  assign n6525 = ~pi70  & ~n6507;
  assign n6526 = pi71  & ~n6525;
  assign n6527 = ~pi71  & n6525;
  assign n6528 = n6053 & ~n6507;
  assign n6529 = ~n6526 & ~n32589;
  assign n6530 = ~n32588 & n6529;
  assign n6531 = ~n6512 & ~n6530;
  assign n6532 = ~n5648 & ~n6531;
  assign n6533 = ~n6051 & ~n6505;
  assign n6534 = ~n32586 & n6533;
  assign n6535 = ~n6499 & n6534;
  assign n6536 = ~n32589 & ~n6535;
  assign n6537 = pi72  & ~n6536;
  assign n6538 = ~pi72  & ~n6535;
  assign n6539 = ~pi72  & n6536;
  assign n6540 = ~n32589 & n6538;
  assign n6541 = ~n6537 & ~n32590;
  assign n6542 = n5648 & ~n6512;
  assign n6543 = n5648 & n6531;
  assign n6544 = ~n6530 & n6542;
  assign n6545 = ~n6541 & ~n32591;
  assign n6546 = ~n6532 & ~n6545;
  assign n6547 = ~n5223 & ~n6546;
  assign n6548 = n5223 & ~n6532;
  assign n6549 = ~n6545 & n6548;
  assign n6550 = ~n6056 & ~n32528;
  assign n6551 = ~n6507 & n6550;
  assign n6552 = n6061 & ~n6551;
  assign n6553 = ~n6061 & n6550;
  assign n6554 = ~n6061 & n6551;
  assign n6555 = ~n6507 & n6553;
  assign n6556 = ~n6552 & ~n32592;
  assign n6557 = ~n6549 & ~n6556;
  assign n6558 = ~n6547 & ~n6557;
  assign n6559 = ~n4851 & ~n6558;
  assign n6560 = ~n6076 & ~n6078;
  assign n6561 = ~n6507 & n6560;
  assign n6562 = ~n6087 & ~n6561;
  assign n6563 = ~n6078 & n6087;
  assign n6564 = ~n6076 & n6563;
  assign n6565 = n6087 & n6561;
  assign n6566 = ~n6507 & n6564;
  assign n6567 = ~n6562 & ~n32593;
  assign n6568 = n4851 & ~n6547;
  assign n6569 = n4851 & n6558;
  assign n6570 = ~n6557 & n6568;
  assign n6571 = ~n6567 & ~n32594;
  assign n6572 = ~n6559 & ~n6571;
  assign n6573 = ~n4461 & ~n6572;
  assign n6574 = n4461 & ~n6559;
  assign n6575 = ~n6571 & n6574;
  assign n6576 = ~n6090 & ~n32530;
  assign n6577 = ~n6507 & n6576;
  assign n6578 = ~n6100 & ~n6577;
  assign n6579 = ~n6090 & n6100;
  assign n6580 = ~n32530 & n6579;
  assign n6581 = n6100 & n6577;
  assign n6582 = ~n6507 & n6580;
  assign n6583 = n6100 & ~n6577;
  assign n6584 = ~n6100 & n6577;
  assign n6585 = ~n6583 & ~n6584;
  assign n6586 = ~n6578 & ~n32595;
  assign n6587 = ~n6575 & n32596;
  assign n6588 = ~n6573 & ~n6587;
  assign n6589 = ~n4115 & ~n6588;
  assign n6590 = ~n6103 & ~n6105;
  assign n6591 = ~n6507 & n6590;
  assign n6592 = ~n32533 & ~n6591;
  assign n6593 = ~n6105 & n32533;
  assign n6594 = ~n6103 & n6593;
  assign n6595 = n32533 & n6591;
  assign n6596 = ~n6507 & n6594;
  assign n6597 = ~n6592 & ~n32597;
  assign n6598 = n4115 & ~n6573;
  assign n6599 = n4115 & n6588;
  assign n6600 = ~n6587 & n6598;
  assign n6601 = ~n6597 & ~n32598;
  assign n6602 = ~n6589 & ~n6601;
  assign n6603 = ~n3754 & ~n6602;
  assign n6604 = n3754 & ~n6589;
  assign n6605 = ~n6601 & n6604;
  assign n6606 = ~n6120 & ~n32534;
  assign n6607 = ~n6507 & n6606;
  assign n6608 = ~n32536 & ~n6607;
  assign n6609 = n32536 & n6607;
  assign n6610 = ~n6120 & ~n32536;
  assign n6611 = ~n32534 & n6610;
  assign n6612 = ~n6507 & n6611;
  assign n6613 = n32536 & ~n6607;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = ~n6608 & ~n6609;
  assign n6616 = ~n6605 & ~n32599;
  assign n6617 = ~n6603 & ~n6616;
  assign n6618 = ~n3444 & ~n6617;
  assign n6619 = ~n6137 & ~n6139;
  assign n6620 = ~n6507 & n6619;
  assign n6621 = ~n32538 & ~n6620;
  assign n6622 = ~n6139 & n32538;
  assign n6623 = ~n6137 & n6622;
  assign n6624 = n32538 & n6620;
  assign n6625 = ~n6507 & n6623;
  assign n6626 = ~n6621 & ~n32600;
  assign n6627 = n3444 & ~n6603;
  assign n6628 = n3444 & n6617;
  assign n6629 = ~n6616 & n6627;
  assign n6630 = ~n6626 & ~n32601;
  assign n6631 = ~n6618 & ~n6630;
  assign n6632 = ~n3116 & ~n6631;
  assign n6633 = n3116 & ~n6618;
  assign n6634 = ~n6630 & n6633;
  assign n6635 = ~n6154 & ~n32539;
  assign n6636 = ~n6507 & n6635;
  assign n6637 = ~n32540 & n6636;
  assign n6638 = n32540 & ~n6636;
  assign n6639 = ~n6154 & n32540;
  assign n6640 = ~n32539 & n6639;
  assign n6641 = ~n6507 & n6640;
  assign n6642 = ~n32540 & ~n6636;
  assign n6643 = ~n6641 & ~n6642;
  assign n6644 = ~n6637 & ~n6638;
  assign n6645 = ~n6634 & ~n32602;
  assign n6646 = ~n6632 & ~n6645;
  assign n6647 = ~n2833 & ~n6646;
  assign n6648 = ~n6170 & ~n6172;
  assign n6649 = ~n6507 & n6648;
  assign n6650 = ~n32542 & ~n6649;
  assign n6651 = ~n6172 & n32542;
  assign n6652 = ~n6170 & n6651;
  assign n6653 = n32542 & n6649;
  assign n6654 = ~n6507 & n6652;
  assign n6655 = ~n6650 & ~n32603;
  assign n6656 = n2833 & ~n6632;
  assign n6657 = n2833 & n6646;
  assign n6658 = ~n6645 & n6656;
  assign n6659 = ~n6655 & ~n32604;
  assign n6660 = ~n6647 & ~n6659;
  assign n6661 = ~n2536 & ~n6660;
  assign n6662 = n2536 & ~n6647;
  assign n6663 = ~n6659 & n6662;
  assign n6664 = ~n6187 & ~n32543;
  assign n6665 = ~n6507 & n6664;
  assign n6666 = ~n32544 & n6665;
  assign n6667 = n32544 & ~n6665;
  assign n6668 = ~n32544 & ~n6665;
  assign n6669 = ~n6187 & n32544;
  assign n6670 = ~n32543 & n6669;
  assign n6671 = n32544 & n6665;
  assign n6672 = ~n6507 & n6670;
  assign n6673 = ~n6668 & ~n32605;
  assign n6674 = ~n6666 & ~n6667;
  assign n6675 = ~n6663 & ~n32606;
  assign n6676 = ~n6661 & ~n6675;
  assign n6677 = ~n2283 & ~n6676;
  assign n6678 = ~n6203 & ~n6205;
  assign n6679 = ~n6507 & n6678;
  assign n6680 = ~n32546 & ~n6679;
  assign n6681 = ~n6205 & n32546;
  assign n6682 = ~n6203 & n6681;
  assign n6683 = n32546 & n6679;
  assign n6684 = ~n6507 & n6682;
  assign n6685 = ~n6680 & ~n32607;
  assign n6686 = n2283 & ~n6661;
  assign n6687 = n2283 & n6676;
  assign n6688 = ~n6675 & n6686;
  assign n6689 = ~n6685 & ~n32608;
  assign n6690 = ~n6677 & ~n6689;
  assign n6691 = ~n2021 & ~n6690;
  assign n6692 = n2021 & ~n6677;
  assign n6693 = ~n6689 & n6692;
  assign n6694 = ~n6220 & ~n32547;
  assign n6695 = ~n6220 & ~n6507;
  assign n6696 = ~n32547 & n6695;
  assign n6697 = ~n6507 & n6694;
  assign n6698 = n32549 & ~n32609;
  assign n6699 = n6235 & n6695;
  assign n6700 = ~n32549 & n32609;
  assign n6701 = ~n6220 & n32549;
  assign n6702 = ~n32547 & n6701;
  assign n6703 = ~n6507 & n6702;
  assign n6704 = ~n32549 & ~n32609;
  assign n6705 = ~n6703 & ~n6704;
  assign n6706 = ~n6698 & ~n32610;
  assign n6707 = ~n6693 & ~n32611;
  assign n6708 = ~n6691 & ~n6707;
  assign n6709 = ~n1796 & ~n6708;
  assign n6710 = ~n6237 & ~n6239;
  assign n6711 = ~n6507 & n6710;
  assign n6712 = ~n32551 & ~n6711;
  assign n6713 = ~n6239 & n32551;
  assign n6714 = ~n6237 & n6713;
  assign n6715 = n32551 & n6711;
  assign n6716 = ~n6507 & n6714;
  assign n6717 = ~n6712 & ~n32612;
  assign n6718 = n1796 & ~n6691;
  assign n6719 = n1796 & n6708;
  assign n6720 = ~n6707 & n6718;
  assign n6721 = ~n6717 & ~n32613;
  assign n6722 = ~n6709 & ~n6721;
  assign n6723 = ~n1567 & ~n6722;
  assign n6724 = ~n6254 & ~n32552;
  assign n6725 = ~n6507 & n6724;
  assign n6726 = ~n32555 & ~n6725;
  assign n6727 = ~n6254 & n32555;
  assign n6728 = ~n32552 & n6727;
  assign n6729 = n32555 & n6725;
  assign n6730 = ~n6507 & n6728;
  assign n6731 = ~n6726 & ~n32614;
  assign n6732 = n1567 & ~n6709;
  assign n6733 = ~n6721 & n6732;
  assign n6734 = ~n6731 & ~n6733;
  assign n6735 = ~n6723 & ~n6734;
  assign n6736 = ~n1374 & ~n6735;
  assign n6737 = ~n6273 & ~n6275;
  assign n6738 = ~n6507 & n6737;
  assign n6739 = ~n32557 & ~n6738;
  assign n6740 = ~n6275 & n32557;
  assign n6741 = ~n6273 & n6740;
  assign n6742 = n32557 & n6738;
  assign n6743 = ~n6507 & n6741;
  assign n6744 = ~n6739 & ~n32615;
  assign n6745 = n1374 & ~n6723;
  assign n6746 = n1374 & n6735;
  assign n6747 = ~n6734 & n6745;
  assign n6748 = ~n6744 & ~n32616;
  assign n6749 = ~n6736 & ~n6748;
  assign n6750 = ~n1179 & ~n6749;
  assign n6751 = n1179 & ~n6736;
  assign n6752 = ~n6748 & n6751;
  assign n6753 = ~n6290 & ~n32559;
  assign n6754 = ~n6290 & ~n6507;
  assign n6755 = ~n32559 & n6754;
  assign n6756 = ~n6507 & n6753;
  assign n6757 = n6298 & ~n32617;
  assign n6758 = n6302 & n6754;
  assign n6759 = ~n6290 & n6298;
  assign n6760 = ~n32559 & n6759;
  assign n6761 = ~n6507 & n6760;
  assign n6762 = ~n6298 & ~n32617;
  assign n6763 = ~n6761 & ~n6762;
  assign n6764 = ~n6757 & ~n6758;
  assign n6765 = ~n6752 & ~n32618;
  assign n6766 = ~n6750 & ~n6765;
  assign n6767 = ~n1016 & ~n6766;
  assign n6768 = ~n6304 & ~n6306;
  assign n6769 = ~n6507 & n6768;
  assign n6770 = ~n32561 & ~n6769;
  assign n6771 = ~n6306 & n32561;
  assign n6772 = ~n6304 & n6771;
  assign n6773 = n32561 & n6769;
  assign n6774 = ~n6507 & n6772;
  assign n6775 = ~n6770 & ~n32619;
  assign n6776 = n1016 & ~n6750;
  assign n6777 = n1016 & n6766;
  assign n6778 = ~n6765 & n6776;
  assign n6779 = ~n6775 & ~n32620;
  assign n6780 = ~n6767 & ~n6779;
  assign n6781 = ~n855 & ~n6780;
  assign n6782 = ~n6321 & ~n32562;
  assign n6783 = ~n6507 & n6782;
  assign n6784 = ~n32564 & ~n6783;
  assign n6785 = ~n6321 & n32564;
  assign n6786 = ~n32562 & n6785;
  assign n6787 = n32564 & n6783;
  assign n6788 = ~n6507 & n6786;
  assign n6789 = ~n6784 & ~n32621;
  assign n6790 = n855 & ~n6767;
  assign n6791 = ~n6779 & n6790;
  assign n6792 = ~n6789 & ~n6791;
  assign n6793 = ~n6781 & ~n6792;
  assign n6794 = ~n720 & ~n6793;
  assign n6795 = ~n6339 & ~n6341;
  assign n6796 = ~n6507 & n6795;
  assign n6797 = ~n32566 & ~n6796;
  assign n6798 = ~n6341 & n32566;
  assign n6799 = ~n6339 & n6798;
  assign n6800 = n32566 & n6796;
  assign n6801 = ~n6507 & n6799;
  assign n6802 = ~n6797 & ~n32622;
  assign n6803 = n720 & ~n6781;
  assign n6804 = n720 & n6793;
  assign n6805 = ~n6792 & n6803;
  assign n6806 = ~n6802 & ~n32623;
  assign n6807 = ~n6794 & ~n6806;
  assign n6808 = ~n592 & ~n6807;
  assign n6809 = n592 & ~n6794;
  assign n6810 = ~n6806 & n6809;
  assign n6811 = ~n6356 & ~n32568;
  assign n6812 = ~n6356 & ~n6507;
  assign n6813 = ~n32568 & n6812;
  assign n6814 = ~n6507 & n6811;
  assign n6815 = n6364 & ~n32624;
  assign n6816 = n6368 & n6812;
  assign n6817 = ~n6356 & n6364;
  assign n6818 = ~n32568 & n6817;
  assign n6819 = ~n6507 & n6818;
  assign n6820 = ~n6364 & ~n32624;
  assign n6821 = ~n6819 & ~n6820;
  assign n6822 = ~n6815 & ~n6816;
  assign n6823 = ~n6810 & ~n32625;
  assign n6824 = ~n6808 & ~n6823;
  assign n6825 = ~n487 & ~n6824;
  assign n6826 = ~n6370 & ~n6372;
  assign n6827 = ~n6507 & n6826;
  assign n6828 = ~n32570 & ~n6827;
  assign n6829 = ~n6372 & n32570;
  assign n6830 = ~n6370 & n6829;
  assign n6831 = n32570 & n6827;
  assign n6832 = ~n6507 & n6830;
  assign n6833 = ~n6828 & ~n32626;
  assign n6834 = n487 & ~n6808;
  assign n6835 = n487 & n6824;
  assign n6836 = ~n6823 & n6834;
  assign n6837 = ~n6833 & ~n32627;
  assign n6838 = ~n6825 & ~n6837;
  assign n6839 = ~n393 & ~n6838;
  assign n6840 = ~n6387 & ~n32571;
  assign n6841 = ~n6507 & n6840;
  assign n6842 = ~n32573 & ~n6841;
  assign n6843 = ~n6387 & n32573;
  assign n6844 = ~n32571 & n6843;
  assign n6845 = n32573 & n6841;
  assign n6846 = ~n6507 & n6844;
  assign n6847 = ~n6842 & ~n32628;
  assign n6848 = n393 & ~n6825;
  assign n6849 = ~n6837 & n6848;
  assign n6850 = ~n6847 & ~n6849;
  assign n6851 = ~n6839 & ~n6850;
  assign n6852 = ~n321 & ~n6851;
  assign n6853 = ~n6405 & ~n6407;
  assign n6854 = ~n6507 & n6853;
  assign n6855 = ~n32575 & ~n6854;
  assign n6856 = ~n6407 & n32575;
  assign n6857 = ~n6405 & n6856;
  assign n6858 = n32575 & n6854;
  assign n6859 = ~n6507 & n6857;
  assign n6860 = ~n6855 & ~n32629;
  assign n6861 = n321 & ~n6839;
  assign n6862 = n321 & n6851;
  assign n6863 = ~n6850 & n6861;
  assign n6864 = ~n6860 & ~n32630;
  assign n6865 = ~n6852 & ~n6864;
  assign n6866 = ~n263 & ~n6865;
  assign n6867 = n263 & ~n6852;
  assign n6868 = ~n6864 & n6867;
  assign n6869 = ~n6422 & ~n32577;
  assign n6870 = ~n6422 & ~n6507;
  assign n6871 = ~n32577 & n6870;
  assign n6872 = ~n6507 & n6869;
  assign n6873 = n6430 & ~n32631;
  assign n6874 = n6434 & n6870;
  assign n6875 = ~n6422 & n6430;
  assign n6876 = ~n32577 & n6875;
  assign n6877 = ~n6507 & n6876;
  assign n6878 = ~n6430 & ~n32631;
  assign n6879 = ~n6877 & ~n6878;
  assign n6880 = ~n6873 & ~n6874;
  assign n6881 = ~n6868 & ~n32632;
  assign n6882 = ~n6866 & ~n6881;
  assign n6883 = ~n214 & ~n6882;
  assign n6884 = ~n6436 & ~n6438;
  assign n6885 = ~n6507 & n6884;
  assign n6886 = ~n32579 & ~n6885;
  assign n6887 = ~n6438 & n32579;
  assign n6888 = ~n6436 & n6887;
  assign n6889 = n32579 & n6885;
  assign n6890 = ~n6507 & n6888;
  assign n6891 = ~n6886 & ~n32633;
  assign n6892 = n214 & ~n6866;
  assign n6893 = n214 & n6882;
  assign n6894 = ~n6881 & n6892;
  assign n6895 = ~n6891 & ~n32634;
  assign n6896 = ~n6883 & ~n6895;
  assign n6897 = ~n197 & ~n6896;
  assign n6898 = n197 & ~n6883;
  assign n6899 = ~n6895 & n6898;
  assign n6900 = ~n6453 & ~n32581;
  assign n6901 = ~n6453 & ~n6507;
  assign n6902 = ~n32581 & n6901;
  assign n6903 = ~n6507 & n6900;
  assign n6904 = n6461 & ~n32635;
  assign n6905 = n6465 & n6901;
  assign n6906 = ~n6453 & n6461;
  assign n6907 = ~n32581 & n6906;
  assign n6908 = ~n6507 & n6907;
  assign n6909 = ~n6461 & ~n32635;
  assign n6910 = ~n6908 & ~n6909;
  assign n6911 = ~n6904 & ~n6905;
  assign n6912 = ~n6899 & ~n32636;
  assign n6913 = ~n6897 & ~n6912;
  assign n6914 = ~n6467 & ~n6469;
  assign n6915 = ~n6507 & n6914;
  assign n6916 = ~n32583 & ~n6915;
  assign n6917 = ~n6469 & n32583;
  assign n6918 = ~n6467 & n6917;
  assign n6919 = n32583 & n6915;
  assign n6920 = ~n6507 & n6918;
  assign n6921 = ~n6916 & ~n32637;
  assign n6922 = ~n6483 & ~n6491;
  assign n6923 = ~n6491 & ~n6507;
  assign n6924 = ~n6483 & n6923;
  assign n6925 = ~n6507 & n6922;
  assign n6926 = ~n32586 & ~n32638;
  assign n6927 = ~n6921 & n6926;
  assign n6928 = ~n6913 & n6927;
  assign n6929 = n193 & ~n6928;
  assign n6930 = ~n6897 & n6921;
  assign n6931 = n6913 & n6921;
  assign n6932 = ~n6912 & n6930;
  assign n6933 = n6483 & ~n6923;
  assign n6934 = ~n193 & ~n6922;
  assign n6935 = ~n6933 & n6934;
  assign n6936 = ~n32639 & ~n6935;
  assign n6937 = ~n6929 & n6936;
  assign n6938 = pi68  & ~n6937;
  assign n6939 = ~pi66  & ~pi67 ;
  assign n6940 = ~pi68  & n6939;
  assign n6941 = ~n6938 & ~n6940;
  assign n6942 = ~n6507 & ~n6941;
  assign n6943 = ~pi68  & ~n6937;
  assign n6944 = pi69  & ~n6943;
  assign n6945 = ~pi69  & n6943;
  assign n6946 = n6509 & ~n6937;
  assign n6947 = ~n6944 & ~n32640;
  assign n6948 = ~n32523 & ~n32587;
  assign n6949 = ~n6030 & n6948;
  assign n6950 = ~n6049 & n6949;
  assign n6951 = ~n32525 & n6950;
  assign n6952 = n6035 & n6051;
  assign n6953 = ~n6043 & n6951;
  assign n6954 = ~n6940 & ~n32641;
  assign n6955 = ~n6505 & n6954;
  assign n6956 = ~n32586 & n6955;
  assign n6957 = ~n6499 & n6956;
  assign n6958 = n6507 & n6941;
  assign n6959 = ~n6938 & n6957;
  assign n6960 = n6947 & ~n32642;
  assign n6961 = ~n6942 & ~n6960;
  assign n6962 = ~n6051 & ~n6961;
  assign n6963 = n6051 & ~n6942;
  assign n6964 = ~n6960 & n6963;
  assign n6965 = ~n6507 & ~n6935;
  assign n6966 = ~n32639 & n6965;
  assign n6967 = ~n6929 & n6966;
  assign n6968 = ~n32640 & ~n6967;
  assign n6969 = pi70  & ~n6968;
  assign n6970 = ~pi70  & ~n6967;
  assign n6971 = ~pi70  & n6968;
  assign n6972 = ~n32640 & n6970;
  assign n6973 = ~n6969 & ~n32643;
  assign n6974 = ~n6964 & ~n6973;
  assign n6975 = ~n6962 & ~n6974;
  assign n6976 = ~n5648 & ~n6975;
  assign n6977 = n5648 & ~n6962;
  assign n6978 = ~n6974 & n6977;
  assign n6979 = n5648 & n6975;
  assign n6980 = ~n6512 & ~n32588;
  assign n6981 = ~n6937 & n6980;
  assign n6982 = n6529 & ~n6981;
  assign n6983 = ~n6529 & n6980;
  assign n6984 = ~n6529 & n6981;
  assign n6985 = ~n6937 & n6983;
  assign n6986 = ~n6982 & ~n32645;
  assign n6987 = ~n32644 & ~n6986;
  assign n6988 = ~n6976 & ~n6987;
  assign n6989 = ~n5223 & ~n6988;
  assign n6990 = n5223 & ~n6976;
  assign n6991 = ~n6987 & n6990;
  assign n6992 = ~n6532 & ~n32591;
  assign n6993 = ~n6532 & ~n6937;
  assign n6994 = ~n32591 & n6993;
  assign n6995 = ~n6937 & n6992;
  assign n6996 = n6541 & ~n32646;
  assign n6997 = n6545 & n6993;
  assign n6998 = n6541 & ~n32591;
  assign n6999 = ~n6532 & n6998;
  assign n7000 = ~n6937 & n6999;
  assign n7001 = ~n6541 & ~n32646;
  assign n7002 = ~n7000 & ~n7001;
  assign n7003 = ~n6996 & ~n6997;
  assign n7004 = ~n6991 & ~n32647;
  assign n7005 = ~n6989 & ~n7004;
  assign n7006 = ~n4851 & ~n7005;
  assign n7007 = n4851 & ~n6989;
  assign n7008 = ~n7004 & n7007;
  assign n7009 = n4851 & n7005;
  assign n7010 = ~n6547 & ~n6549;
  assign n7011 = ~n6937 & n7010;
  assign n7012 = ~n6556 & ~n7011;
  assign n7013 = ~n6547 & n6556;
  assign n7014 = ~n6549 & n7013;
  assign n7015 = n6556 & n7011;
  assign n7016 = ~n6937 & n7014;
  assign n7017 = n6556 & ~n7011;
  assign n7018 = ~n6556 & n7011;
  assign n7019 = ~n7017 & ~n7018;
  assign n7020 = ~n7012 & ~n32649;
  assign n7021 = ~n32648 & n32650;
  assign n7022 = ~n7006 & ~n7021;
  assign n7023 = ~n4461 & ~n7022;
  assign n7024 = n4461 & ~n7006;
  assign n7025 = ~n7021 & n7024;
  assign n7026 = ~n6559 & ~n32594;
  assign n7027 = ~n6559 & ~n6937;
  assign n7028 = ~n32594 & n7027;
  assign n7029 = ~n6937 & n7026;
  assign n7030 = n6567 & ~n32651;
  assign n7031 = n6571 & n7027;
  assign n7032 = n6567 & ~n32594;
  assign n7033 = ~n6559 & n7032;
  assign n7034 = ~n6937 & n7033;
  assign n7035 = ~n6567 & ~n32651;
  assign n7036 = ~n7034 & ~n7035;
  assign n7037 = ~n7030 & ~n7031;
  assign n7038 = ~n7025 & ~n32652;
  assign n7039 = ~n7023 & ~n7038;
  assign n7040 = ~n4115 & ~n7039;
  assign n7041 = n4115 & ~n7023;
  assign n7042 = ~n7038 & n7041;
  assign n7043 = n4115 & n7039;
  assign n7044 = ~n6573 & ~n6575;
  assign n7045 = ~n6937 & n7044;
  assign n7046 = ~n32596 & ~n7045;
  assign n7047 = n32596 & n7045;
  assign n7048 = ~n6573 & ~n32596;
  assign n7049 = ~n6575 & n7048;
  assign n7050 = ~n6937 & n7049;
  assign n7051 = n32596 & ~n7045;
  assign n7052 = ~n7050 & ~n7051;
  assign n7053 = ~n7046 & ~n7047;
  assign n7054 = ~n32653 & ~n32654;
  assign n7055 = ~n7040 & ~n7054;
  assign n7056 = ~n3754 & ~n7055;
  assign n7057 = n3754 & ~n7040;
  assign n7058 = ~n7054 & n7057;
  assign n7059 = ~n6589 & ~n32598;
  assign n7060 = ~n6589 & ~n6937;
  assign n7061 = ~n32598 & n7060;
  assign n7062 = ~n6937 & n7059;
  assign n7063 = n6597 & ~n32655;
  assign n7064 = n6601 & n7060;
  assign n7065 = n6597 & ~n32598;
  assign n7066 = ~n6589 & n7065;
  assign n7067 = ~n6937 & n7066;
  assign n7068 = ~n6597 & ~n32655;
  assign n7069 = ~n7067 & ~n7068;
  assign n7070 = ~n7063 & ~n7064;
  assign n7071 = ~n7058 & ~n32656;
  assign n7072 = ~n7056 & ~n7071;
  assign n7073 = ~n3444 & ~n7072;
  assign n7074 = n3444 & ~n7056;
  assign n7075 = ~n7071 & n7074;
  assign n7076 = n3444 & n7072;
  assign n7077 = ~n6603 & ~n6605;
  assign n7078 = ~n6937 & n7077;
  assign n7079 = ~n32599 & n7078;
  assign n7080 = n32599 & ~n7078;
  assign n7081 = ~n6603 & n32599;
  assign n7082 = ~n6605 & n7081;
  assign n7083 = ~n6937 & n7082;
  assign n7084 = ~n32599 & ~n7078;
  assign n7085 = ~n7083 & ~n7084;
  assign n7086 = ~n7079 & ~n7080;
  assign n7087 = ~n32657 & ~n32658;
  assign n7088 = ~n7073 & ~n7087;
  assign n7089 = ~n3116 & ~n7088;
  assign n7090 = n3116 & ~n7073;
  assign n7091 = ~n7087 & n7090;
  assign n7092 = ~n6618 & ~n32601;
  assign n7093 = ~n6618 & ~n6937;
  assign n7094 = ~n32601 & n7093;
  assign n7095 = ~n6937 & n7092;
  assign n7096 = n6626 & ~n32659;
  assign n7097 = n6630 & n7093;
  assign n7098 = n6626 & ~n32601;
  assign n7099 = ~n6618 & n7098;
  assign n7100 = ~n6937 & n7099;
  assign n7101 = ~n6626 & ~n32659;
  assign n7102 = ~n7100 & ~n7101;
  assign n7103 = ~n7096 & ~n7097;
  assign n7104 = ~n7091 & ~n32660;
  assign n7105 = ~n7089 & ~n7104;
  assign n7106 = ~n2833 & ~n7105;
  assign n7107 = n2833 & ~n7089;
  assign n7108 = ~n7104 & n7107;
  assign n7109 = n2833 & n7105;
  assign n7110 = ~n6632 & ~n6634;
  assign n7111 = ~n6937 & n7110;
  assign n7112 = ~n32602 & n7111;
  assign n7113 = n32602 & ~n7111;
  assign n7114 = ~n32602 & ~n7111;
  assign n7115 = ~n6632 & n32602;
  assign n7116 = ~n6634 & n7115;
  assign n7117 = n32602 & n7111;
  assign n7118 = ~n6937 & n7116;
  assign n7119 = ~n7114 & ~n32662;
  assign n7120 = ~n7112 & ~n7113;
  assign n7121 = ~n32661 & ~n32663;
  assign n7122 = ~n7106 & ~n7121;
  assign n7123 = ~n2536 & ~n7122;
  assign n7124 = n2536 & ~n7106;
  assign n7125 = ~n7121 & n7124;
  assign n7126 = ~n6647 & ~n32604;
  assign n7127 = ~n6647 & ~n6937;
  assign n7128 = ~n32604 & n7127;
  assign n7129 = ~n6937 & n7126;
  assign n7130 = n6655 & ~n32664;
  assign n7131 = n6659 & n7127;
  assign n7132 = n6655 & ~n32604;
  assign n7133 = ~n6647 & n7132;
  assign n7134 = ~n6937 & n7133;
  assign n7135 = ~n6655 & ~n32664;
  assign n7136 = ~n7134 & ~n7135;
  assign n7137 = ~n7130 & ~n7131;
  assign n7138 = ~n7125 & ~n32665;
  assign n7139 = ~n7123 & ~n7138;
  assign n7140 = ~n2283 & ~n7139;
  assign n7141 = n2283 & ~n7123;
  assign n7142 = ~n7138 & n7141;
  assign n7143 = n2283 & n7139;
  assign n7144 = ~n6661 & ~n6663;
  assign n7145 = ~n6661 & ~n6937;
  assign n7146 = ~n6663 & n7145;
  assign n7147 = ~n6937 & n7144;
  assign n7148 = n32606 & ~n32667;
  assign n7149 = n6675 & n7145;
  assign n7150 = ~n32606 & n32667;
  assign n7151 = ~n6661 & n32606;
  assign n7152 = ~n6663 & n7151;
  assign n7153 = ~n6937 & n7152;
  assign n7154 = ~n32606 & ~n32667;
  assign n7155 = ~n7153 & ~n7154;
  assign n7156 = ~n7148 & ~n32668;
  assign n7157 = ~n32666 & ~n32669;
  assign n7158 = ~n7140 & ~n7157;
  assign n7159 = ~n2021 & ~n7158;
  assign n7160 = n2021 & ~n7140;
  assign n7161 = ~n7157 & n7160;
  assign n7162 = ~n6677 & ~n32608;
  assign n7163 = ~n6677 & ~n6937;
  assign n7164 = ~n32608 & n7163;
  assign n7165 = ~n6937 & n7162;
  assign n7166 = n6685 & ~n32670;
  assign n7167 = n6689 & n7163;
  assign n7168 = n6685 & ~n32608;
  assign n7169 = ~n6677 & n7168;
  assign n7170 = ~n6937 & n7169;
  assign n7171 = ~n6685 & ~n32670;
  assign n7172 = ~n7170 & ~n7171;
  assign n7173 = ~n7166 & ~n7167;
  assign n7174 = ~n7161 & ~n32671;
  assign n7175 = ~n7159 & ~n7174;
  assign n7176 = ~n1796 & ~n7175;
  assign n7177 = ~n6691 & ~n6693;
  assign n7178 = ~n6937 & n7177;
  assign n7179 = ~n32611 & ~n7178;
  assign n7180 = ~n6691 & n32611;
  assign n7181 = ~n6693 & n7180;
  assign n7182 = n32611 & n7178;
  assign n7183 = ~n6937 & n7181;
  assign n7184 = ~n7179 & ~n32672;
  assign n7185 = n1796 & ~n7159;
  assign n7186 = ~n7174 & n7185;
  assign n7187 = n1796 & n7175;
  assign n7188 = ~n7184 & ~n32673;
  assign n7189 = ~n7176 & ~n7188;
  assign n7190 = ~n1567 & ~n7189;
  assign n7191 = n1567 & ~n7176;
  assign n7192 = ~n7188 & n7191;
  assign n7193 = ~n6709 & ~n32613;
  assign n7194 = ~n6709 & ~n6937;
  assign n7195 = ~n32613 & n7194;
  assign n7196 = ~n6937 & n7193;
  assign n7197 = n6717 & ~n32674;
  assign n7198 = n6721 & n7194;
  assign n7199 = n6717 & ~n32613;
  assign n7200 = ~n6709 & n7199;
  assign n7201 = ~n6937 & n7200;
  assign n7202 = ~n6717 & ~n32674;
  assign n7203 = ~n7201 & ~n7202;
  assign n7204 = ~n7197 & ~n7198;
  assign n7205 = ~n7192 & ~n32675;
  assign n7206 = ~n7190 & ~n7205;
  assign n7207 = ~n1374 & ~n7206;
  assign n7208 = n1374 & ~n7190;
  assign n7209 = ~n7205 & n7208;
  assign n7210 = n1374 & n7206;
  assign n7211 = ~n6723 & ~n6733;
  assign n7212 = ~n6723 & ~n6937;
  assign n7213 = ~n6733 & n7212;
  assign n7214 = ~n6937 & n7211;
  assign n7215 = n6731 & ~n32677;
  assign n7216 = n6734 & n7212;
  assign n7217 = ~n6723 & n6731;
  assign n7218 = ~n6733 & n7217;
  assign n7219 = ~n6937 & n7218;
  assign n7220 = ~n6731 & ~n32677;
  assign n7221 = ~n7219 & ~n7220;
  assign n7222 = ~n7215 & ~n7216;
  assign n7223 = ~n32676 & ~n32678;
  assign n7224 = ~n7207 & ~n7223;
  assign n7225 = ~n1179 & ~n7224;
  assign n7226 = n1179 & ~n7207;
  assign n7227 = ~n7223 & n7226;
  assign n7228 = ~n6736 & ~n32616;
  assign n7229 = ~n6736 & ~n6937;
  assign n7230 = ~n32616 & n7229;
  assign n7231 = ~n6937 & n7228;
  assign n7232 = n6744 & ~n32679;
  assign n7233 = n6748 & n7229;
  assign n7234 = n6744 & ~n32616;
  assign n7235 = ~n6736 & n7234;
  assign n7236 = ~n6937 & n7235;
  assign n7237 = ~n6744 & ~n32679;
  assign n7238 = ~n7236 & ~n7237;
  assign n7239 = ~n7232 & ~n7233;
  assign n7240 = ~n7227 & ~n32680;
  assign n7241 = ~n7225 & ~n7240;
  assign n7242 = ~n1016 & ~n7241;
  assign n7243 = ~n6750 & ~n6752;
  assign n7244 = ~n6937 & n7243;
  assign n7245 = ~n32618 & ~n7244;
  assign n7246 = ~n6750 & n32618;
  assign n7247 = ~n6752 & n7246;
  assign n7248 = n32618 & n7244;
  assign n7249 = ~n6937 & n7247;
  assign n7250 = ~n7245 & ~n32681;
  assign n7251 = n1016 & ~n7225;
  assign n7252 = ~n7240 & n7251;
  assign n7253 = n1016 & n7241;
  assign n7254 = ~n7250 & ~n32682;
  assign n7255 = ~n7242 & ~n7254;
  assign n7256 = ~n855 & ~n7255;
  assign n7257 = n855 & ~n7242;
  assign n7258 = ~n7254 & n7257;
  assign n7259 = ~n6767 & ~n32620;
  assign n7260 = ~n6767 & ~n6937;
  assign n7261 = ~n32620 & n7260;
  assign n7262 = ~n6937 & n7259;
  assign n7263 = n6775 & ~n32683;
  assign n7264 = n6779 & n7260;
  assign n7265 = n6775 & ~n32620;
  assign n7266 = ~n6767 & n7265;
  assign n7267 = ~n6937 & n7266;
  assign n7268 = ~n6775 & ~n32683;
  assign n7269 = ~n7267 & ~n7268;
  assign n7270 = ~n7263 & ~n7264;
  assign n7271 = ~n7258 & ~n32684;
  assign n7272 = ~n7256 & ~n7271;
  assign n7273 = ~n720 & ~n7272;
  assign n7274 = n720 & ~n7256;
  assign n7275 = ~n7271 & n7274;
  assign n7276 = n720 & n7272;
  assign n7277 = ~n6781 & ~n6791;
  assign n7278 = ~n6781 & ~n6937;
  assign n7279 = ~n6791 & n7278;
  assign n7280 = ~n6937 & n7277;
  assign n7281 = n6789 & ~n32686;
  assign n7282 = n6792 & n7278;
  assign n7283 = ~n6781 & n6789;
  assign n7284 = ~n6791 & n7283;
  assign n7285 = ~n6937 & n7284;
  assign n7286 = ~n6789 & ~n32686;
  assign n7287 = ~n7285 & ~n7286;
  assign n7288 = ~n7281 & ~n7282;
  assign n7289 = ~n32685 & ~n32687;
  assign n7290 = ~n7273 & ~n7289;
  assign n7291 = ~n592 & ~n7290;
  assign n7292 = n592 & ~n7273;
  assign n7293 = ~n7289 & n7292;
  assign n7294 = ~n6794 & ~n32623;
  assign n7295 = ~n6794 & ~n6937;
  assign n7296 = ~n32623 & n7295;
  assign n7297 = ~n6937 & n7294;
  assign n7298 = n6802 & ~n32688;
  assign n7299 = n6806 & n7295;
  assign n7300 = n6802 & ~n32623;
  assign n7301 = ~n6794 & n7300;
  assign n7302 = ~n6937 & n7301;
  assign n7303 = ~n6802 & ~n32688;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = ~n7298 & ~n7299;
  assign n7306 = ~n7293 & ~n32689;
  assign n7307 = ~n7291 & ~n7306;
  assign n7308 = ~n487 & ~n7307;
  assign n7309 = ~n6808 & ~n6810;
  assign n7310 = ~n6937 & n7309;
  assign n7311 = ~n32625 & ~n7310;
  assign n7312 = ~n6808 & n32625;
  assign n7313 = ~n6810 & n7312;
  assign n7314 = n32625 & n7310;
  assign n7315 = ~n6937 & n7313;
  assign n7316 = ~n7311 & ~n32690;
  assign n7317 = n487 & ~n7291;
  assign n7318 = ~n7306 & n7317;
  assign n7319 = n487 & n7307;
  assign n7320 = ~n7316 & ~n32691;
  assign n7321 = ~n7308 & ~n7320;
  assign n7322 = ~n393 & ~n7321;
  assign n7323 = n393 & ~n7308;
  assign n7324 = ~n7320 & n7323;
  assign n7325 = ~n6825 & ~n32627;
  assign n7326 = ~n6825 & ~n6937;
  assign n7327 = ~n32627 & n7326;
  assign n7328 = ~n6937 & n7325;
  assign n7329 = n6833 & ~n32692;
  assign n7330 = n6837 & n7326;
  assign n7331 = n6833 & ~n32627;
  assign n7332 = ~n6825 & n7331;
  assign n7333 = ~n6937 & n7332;
  assign n7334 = ~n6833 & ~n32692;
  assign n7335 = ~n7333 & ~n7334;
  assign n7336 = ~n7329 & ~n7330;
  assign n7337 = ~n7324 & ~n32693;
  assign n7338 = ~n7322 & ~n7337;
  assign n7339 = ~n321 & ~n7338;
  assign n7340 = n321 & ~n7322;
  assign n7341 = ~n7337 & n7340;
  assign n7342 = n321 & n7338;
  assign n7343 = ~n6839 & ~n6849;
  assign n7344 = ~n6839 & ~n6937;
  assign n7345 = ~n6849 & n7344;
  assign n7346 = ~n6937 & n7343;
  assign n7347 = n6847 & ~n32695;
  assign n7348 = n6850 & n7344;
  assign n7349 = ~n6839 & n6847;
  assign n7350 = ~n6849 & n7349;
  assign n7351 = ~n6937 & n7350;
  assign n7352 = ~n6847 & ~n32695;
  assign n7353 = ~n7351 & ~n7352;
  assign n7354 = ~n7347 & ~n7348;
  assign n7355 = ~n32694 & ~n32696;
  assign n7356 = ~n7339 & ~n7355;
  assign n7357 = ~n263 & ~n7356;
  assign n7358 = n263 & ~n7339;
  assign n7359 = ~n7355 & n7358;
  assign n7360 = ~n6852 & ~n32630;
  assign n7361 = ~n6852 & ~n6937;
  assign n7362 = ~n32630 & n7361;
  assign n7363 = ~n6937 & n7360;
  assign n7364 = n6860 & ~n32697;
  assign n7365 = n6864 & n7361;
  assign n7366 = n6860 & ~n32630;
  assign n7367 = ~n6852 & n7366;
  assign n7368 = ~n6937 & n7367;
  assign n7369 = ~n6860 & ~n32697;
  assign n7370 = ~n7368 & ~n7369;
  assign n7371 = ~n7364 & ~n7365;
  assign n7372 = ~n7359 & ~n32698;
  assign n7373 = ~n7357 & ~n7372;
  assign n7374 = ~n214 & ~n7373;
  assign n7375 = ~n6866 & ~n6868;
  assign n7376 = ~n6937 & n7375;
  assign n7377 = ~n32632 & ~n7376;
  assign n7378 = ~n6866 & n32632;
  assign n7379 = ~n6868 & n7378;
  assign n7380 = n32632 & n7376;
  assign n7381 = ~n6937 & n7379;
  assign n7382 = ~n7377 & ~n32699;
  assign n7383 = n214 & ~n7357;
  assign n7384 = ~n7372 & n7383;
  assign n7385 = n214 & n7373;
  assign n7386 = ~n7382 & ~n32700;
  assign n7387 = ~n7374 & ~n7386;
  assign n7388 = ~n197 & ~n7387;
  assign n7389 = n197 & ~n7374;
  assign n7390 = ~n7386 & n7389;
  assign n7391 = ~n6883 & ~n32634;
  assign n7392 = ~n6883 & ~n6937;
  assign n7393 = ~n32634 & n7392;
  assign n7394 = ~n6937 & n7391;
  assign n7395 = n6891 & ~n32701;
  assign n7396 = n6895 & n7392;
  assign n7397 = n6891 & ~n32634;
  assign n7398 = ~n6883 & n7397;
  assign n7399 = ~n6937 & n7398;
  assign n7400 = ~n6891 & ~n32701;
  assign n7401 = ~n7399 & ~n7400;
  assign n7402 = ~n7395 & ~n7396;
  assign n7403 = ~n7390 & ~n32702;
  assign n7404 = ~n7388 & ~n7403;
  assign n7405 = ~n6897 & ~n6899;
  assign n7406 = ~n6937 & n7405;
  assign n7407 = ~n32636 & ~n7406;
  assign n7408 = ~n6897 & n32636;
  assign n7409 = ~n6899 & n7408;
  assign n7410 = n32636 & n7406;
  assign n7411 = ~n6937 & n7409;
  assign n7412 = ~n7407 & ~n32703;
  assign n7413 = ~n6913 & ~n6921;
  assign n7414 = ~n6921 & ~n6937;
  assign n7415 = ~n6913 & n7414;
  assign n7416 = ~n6937 & n7413;
  assign n7417 = ~n32639 & ~n32704;
  assign n7418 = ~n7412 & n7417;
  assign n7419 = ~n7404 & n7418;
  assign n7420 = n193 & ~n7419;
  assign n7421 = ~n7388 & n7412;
  assign n7422 = ~n7403 & n7421;
  assign n7423 = n7404 & n7412;
  assign n7424 = n6913 & ~n7414;
  assign n7425 = ~n193 & ~n7413;
  assign n7426 = ~n7424 & n7425;
  assign n7427 = ~n32705 & ~n7426;
  assign n7428 = ~n7420 & n7427;
  assign n7429 = pi66  & ~n7428;
  assign n7430 = ~pi64  & ~pi65 ;
  assign n7431 = ~pi66  & n7430;
  assign n7432 = ~n7429 & ~n7431;
  assign n7433 = ~n6937 & ~n7432;
  assign n7434 = ~n32584 & ~n32641;
  assign n7435 = ~n6486 & n7434;
  assign n7436 = ~n6505 & n7435;
  assign n7437 = ~n32586 & n7436;
  assign n7438 = n6491 & n6507;
  assign n7439 = ~n6499 & n7437;
  assign n7440 = ~n7431 & ~n32706;
  assign n7441 = ~n6935 & n7440;
  assign n7442 = ~n32639 & n7441;
  assign n7443 = ~n6929 & n7442;
  assign n7444 = n6937 & n7432;
  assign n7445 = ~n7429 & n7443;
  assign n7446 = ~pi66  & ~n7428;
  assign n7447 = pi67  & ~n7446;
  assign n7448 = ~pi67  & n7446;
  assign n7449 = n6939 & ~n7428;
  assign n7450 = ~n7447 & ~n32708;
  assign n7451 = ~n32707 & n7450;
  assign n7452 = ~n7433 & ~n7451;
  assign n7453 = ~n6507 & ~n7452;
  assign n7454 = ~n6937 & ~n7426;
  assign n7455 = ~n32705 & n7454;
  assign n7456 = ~n7420 & n7455;
  assign n7457 = ~n32708 & ~n7456;
  assign n7458 = pi68  & ~n7457;
  assign n7459 = ~pi68  & ~n7456;
  assign n7460 = ~pi68  & n7457;
  assign n7461 = ~n32708 & n7459;
  assign n7462 = ~n7458 & ~n32709;
  assign n7463 = n6507 & ~n7433;
  assign n7464 = n6507 & n7452;
  assign n7465 = ~n7451 & n7463;
  assign n7466 = ~n7462 & ~n32710;
  assign n7467 = ~n7453 & ~n7466;
  assign n7468 = ~n6051 & ~n7467;
  assign n7469 = n6051 & ~n7453;
  assign n7470 = ~n7466 & n7469;
  assign n7471 = ~n6942 & ~n32642;
  assign n7472 = ~n7428 & n7471;
  assign n7473 = n6947 & ~n7472;
  assign n7474 = ~n6947 & n7471;
  assign n7475 = ~n6947 & n7472;
  assign n7476 = ~n7428 & n7474;
  assign n7477 = ~n7473 & ~n32711;
  assign n7478 = ~n7470 & ~n7477;
  assign n7479 = ~n7468 & ~n7478;
  assign n7480 = ~n5648 & ~n7479;
  assign n7481 = ~n6962 & ~n6964;
  assign n7482 = ~n7428 & n7481;
  assign n7483 = ~n6973 & ~n7482;
  assign n7484 = ~n6964 & n6973;
  assign n7485 = ~n6962 & n7484;
  assign n7486 = n6973 & n7482;
  assign n7487 = ~n7428 & n7485;
  assign n7488 = ~n7483 & ~n32712;
  assign n7489 = n5648 & ~n7468;
  assign n7490 = n5648 & n7479;
  assign n7491 = ~n7478 & n7489;
  assign n7492 = ~n7488 & ~n32713;
  assign n7493 = ~n7480 & ~n7492;
  assign n7494 = ~n5223 & ~n7493;
  assign n7495 = n5223 & ~n7480;
  assign n7496 = ~n7492 & n7495;
  assign n7497 = ~n6976 & ~n32644;
  assign n7498 = ~n7428 & n7497;
  assign n7499 = ~n6986 & ~n7498;
  assign n7500 = ~n6976 & n6986;
  assign n7501 = ~n32644 & n7500;
  assign n7502 = n6986 & n7498;
  assign n7503 = ~n7428 & n7501;
  assign n7504 = n6986 & ~n7498;
  assign n7505 = ~n6986 & n7498;
  assign n7506 = ~n7504 & ~n7505;
  assign n7507 = ~n7499 & ~n32714;
  assign n7508 = ~n7496 & n32715;
  assign n7509 = ~n7494 & ~n7508;
  assign n7510 = ~n4851 & ~n7509;
  assign n7511 = ~n6989 & ~n6991;
  assign n7512 = ~n7428 & n7511;
  assign n7513 = ~n32647 & ~n7512;
  assign n7514 = ~n6991 & n32647;
  assign n7515 = ~n6989 & n7514;
  assign n7516 = n32647 & n7512;
  assign n7517 = ~n7428 & n7515;
  assign n7518 = ~n7513 & ~n32716;
  assign n7519 = n4851 & ~n7494;
  assign n7520 = n4851 & n7509;
  assign n7521 = ~n7508 & n7519;
  assign n7522 = ~n7518 & ~n32717;
  assign n7523 = ~n7510 & ~n7522;
  assign n7524 = ~n4461 & ~n7523;
  assign n7525 = n4461 & ~n7510;
  assign n7526 = ~n7522 & n7525;
  assign n7527 = ~n7006 & ~n32648;
  assign n7528 = ~n7428 & n7527;
  assign n7529 = ~n32650 & ~n7528;
  assign n7530 = n32650 & n7528;
  assign n7531 = ~n7006 & ~n32650;
  assign n7532 = ~n32648 & n7531;
  assign n7533 = ~n7428 & n7532;
  assign n7534 = n32650 & ~n7528;
  assign n7535 = ~n7533 & ~n7534;
  assign n7536 = ~n7529 & ~n7530;
  assign n7537 = ~n7526 & ~n32718;
  assign n7538 = ~n7524 & ~n7537;
  assign n7539 = ~n4115 & ~n7538;
  assign n7540 = ~n7023 & ~n7025;
  assign n7541 = ~n7428 & n7540;
  assign n7542 = ~n32652 & ~n7541;
  assign n7543 = ~n7025 & n32652;
  assign n7544 = ~n7023 & n7543;
  assign n7545 = n32652 & n7541;
  assign n7546 = ~n7428 & n7544;
  assign n7547 = ~n7542 & ~n32719;
  assign n7548 = n4115 & ~n7524;
  assign n7549 = n4115 & n7538;
  assign n7550 = ~n7537 & n7548;
  assign n7551 = ~n7547 & ~n32720;
  assign n7552 = ~n7539 & ~n7551;
  assign n7553 = ~n3754 & ~n7552;
  assign n7554 = n3754 & ~n7539;
  assign n7555 = ~n7551 & n7554;
  assign n7556 = ~n7040 & ~n32653;
  assign n7557 = ~n7428 & n7556;
  assign n7558 = ~n32654 & n7557;
  assign n7559 = n32654 & ~n7557;
  assign n7560 = ~n7040 & n32654;
  assign n7561 = ~n32653 & n7560;
  assign n7562 = ~n7428 & n7561;
  assign n7563 = ~n32654 & ~n7557;
  assign n7564 = ~n7562 & ~n7563;
  assign n7565 = ~n7558 & ~n7559;
  assign n7566 = ~n7555 & ~n32721;
  assign n7567 = ~n7553 & ~n7566;
  assign n7568 = ~n3444 & ~n7567;
  assign n7569 = ~n7056 & ~n7058;
  assign n7570 = ~n7428 & n7569;
  assign n7571 = ~n32656 & ~n7570;
  assign n7572 = ~n7058 & n32656;
  assign n7573 = ~n7056 & n7572;
  assign n7574 = n32656 & n7570;
  assign n7575 = ~n7428 & n7573;
  assign n7576 = ~n7571 & ~n32722;
  assign n7577 = n3444 & ~n7553;
  assign n7578 = n3444 & n7567;
  assign n7579 = ~n7566 & n7577;
  assign n7580 = ~n7576 & ~n32723;
  assign n7581 = ~n7568 & ~n7580;
  assign n7582 = ~n3116 & ~n7581;
  assign n7583 = n3116 & ~n7568;
  assign n7584 = ~n7580 & n7583;
  assign n7585 = ~n7073 & ~n32657;
  assign n7586 = ~n7428 & n7585;
  assign n7587 = ~n32658 & n7586;
  assign n7588 = n32658 & ~n7586;
  assign n7589 = ~n32658 & ~n7586;
  assign n7590 = ~n7073 & n32658;
  assign n7591 = ~n32657 & n7590;
  assign n7592 = n32658 & n7586;
  assign n7593 = ~n7428 & n7591;
  assign n7594 = ~n7589 & ~n32724;
  assign n7595 = ~n7587 & ~n7588;
  assign n7596 = ~n7584 & ~n32725;
  assign n7597 = ~n7582 & ~n7596;
  assign n7598 = ~n2833 & ~n7597;
  assign n7599 = ~n7089 & ~n7091;
  assign n7600 = ~n7428 & n7599;
  assign n7601 = ~n32660 & ~n7600;
  assign n7602 = ~n7091 & n32660;
  assign n7603 = ~n7089 & n7602;
  assign n7604 = n32660 & n7600;
  assign n7605 = ~n7428 & n7603;
  assign n7606 = ~n7601 & ~n32726;
  assign n7607 = n2833 & ~n7582;
  assign n7608 = n2833 & n7597;
  assign n7609 = ~n7596 & n7607;
  assign n7610 = ~n7606 & ~n32727;
  assign n7611 = ~n7598 & ~n7610;
  assign n7612 = ~n2536 & ~n7611;
  assign n7613 = n2536 & ~n7598;
  assign n7614 = ~n7610 & n7613;
  assign n7615 = ~n7106 & ~n32661;
  assign n7616 = ~n7106 & ~n7428;
  assign n7617 = ~n32661 & n7616;
  assign n7618 = ~n7428 & n7615;
  assign n7619 = n32663 & ~n32728;
  assign n7620 = n7121 & n7616;
  assign n7621 = ~n32663 & n32728;
  assign n7622 = ~n7106 & n32663;
  assign n7623 = ~n32661 & n7622;
  assign n7624 = ~n7428 & n7623;
  assign n7625 = ~n32663 & ~n32728;
  assign n7626 = ~n7624 & ~n7625;
  assign n7627 = ~n7619 & ~n32729;
  assign n7628 = ~n7614 & ~n32730;
  assign n7629 = ~n7612 & ~n7628;
  assign n7630 = ~n2283 & ~n7629;
  assign n7631 = ~n7123 & ~n7125;
  assign n7632 = ~n7428 & n7631;
  assign n7633 = ~n32665 & ~n7632;
  assign n7634 = ~n7125 & n32665;
  assign n7635 = ~n7123 & n7634;
  assign n7636 = n32665 & n7632;
  assign n7637 = ~n7428 & n7635;
  assign n7638 = ~n7633 & ~n32731;
  assign n7639 = n2283 & ~n7612;
  assign n7640 = n2283 & n7629;
  assign n7641 = ~n7628 & n7639;
  assign n7642 = ~n7638 & ~n32732;
  assign n7643 = ~n7630 & ~n7642;
  assign n7644 = ~n2021 & ~n7643;
  assign n7645 = ~n7140 & ~n32666;
  assign n7646 = ~n7428 & n7645;
  assign n7647 = ~n32669 & ~n7646;
  assign n7648 = ~n7140 & n32669;
  assign n7649 = ~n32666 & n7648;
  assign n7650 = n32669 & n7646;
  assign n7651 = ~n7428 & n7649;
  assign n7652 = ~n7647 & ~n32733;
  assign n7653 = n2021 & ~n7630;
  assign n7654 = ~n7642 & n7653;
  assign n7655 = ~n7652 & ~n7654;
  assign n7656 = ~n7644 & ~n7655;
  assign n7657 = ~n1796 & ~n7656;
  assign n7658 = ~n7159 & ~n7161;
  assign n7659 = ~n7428 & n7658;
  assign n7660 = ~n32671 & ~n7659;
  assign n7661 = ~n7161 & n32671;
  assign n7662 = ~n7159 & n7661;
  assign n7663 = n32671 & n7659;
  assign n7664 = ~n7428 & n7662;
  assign n7665 = ~n7660 & ~n32734;
  assign n7666 = n1796 & ~n7644;
  assign n7667 = n1796 & n7656;
  assign n7668 = ~n7655 & n7666;
  assign n7669 = ~n7665 & ~n32735;
  assign n7670 = ~n7657 & ~n7669;
  assign n7671 = ~n1567 & ~n7670;
  assign n7672 = n1567 & ~n7657;
  assign n7673 = ~n7669 & n7672;
  assign n7674 = ~n7176 & ~n32673;
  assign n7675 = ~n7176 & ~n7428;
  assign n7676 = ~n32673 & n7675;
  assign n7677 = ~n7428 & n7674;
  assign n7678 = n7184 & ~n32736;
  assign n7679 = n7188 & n7675;
  assign n7680 = ~n7176 & n7184;
  assign n7681 = ~n32673 & n7680;
  assign n7682 = ~n7428 & n7681;
  assign n7683 = ~n7184 & ~n32736;
  assign n7684 = ~n7682 & ~n7683;
  assign n7685 = ~n7678 & ~n7679;
  assign n7686 = ~n7673 & ~n32737;
  assign n7687 = ~n7671 & ~n7686;
  assign n7688 = ~n1374 & ~n7687;
  assign n7689 = ~n7190 & ~n7192;
  assign n7690 = ~n7428 & n7689;
  assign n7691 = ~n32675 & ~n7690;
  assign n7692 = ~n7192 & n32675;
  assign n7693 = ~n7190 & n7692;
  assign n7694 = n32675 & n7690;
  assign n7695 = ~n7428 & n7693;
  assign n7696 = ~n7691 & ~n32738;
  assign n7697 = n1374 & ~n7671;
  assign n7698 = n1374 & n7687;
  assign n7699 = ~n7686 & n7697;
  assign n7700 = ~n7696 & ~n32739;
  assign n7701 = ~n7688 & ~n7700;
  assign n7702 = ~n1179 & ~n7701;
  assign n7703 = ~n7207 & ~n32676;
  assign n7704 = ~n7428 & n7703;
  assign n7705 = ~n32678 & ~n7704;
  assign n7706 = ~n7207 & n32678;
  assign n7707 = ~n32676 & n7706;
  assign n7708 = n32678 & n7704;
  assign n7709 = ~n7428 & n7707;
  assign n7710 = ~n7705 & ~n32740;
  assign n7711 = n1179 & ~n7688;
  assign n7712 = ~n7700 & n7711;
  assign n7713 = ~n7710 & ~n7712;
  assign n7714 = ~n7702 & ~n7713;
  assign n7715 = ~n1016 & ~n7714;
  assign n7716 = ~n7225 & ~n7227;
  assign n7717 = ~n7428 & n7716;
  assign n7718 = ~n32680 & ~n7717;
  assign n7719 = ~n7227 & n32680;
  assign n7720 = ~n7225 & n7719;
  assign n7721 = n32680 & n7717;
  assign n7722 = ~n7428 & n7720;
  assign n7723 = ~n7718 & ~n32741;
  assign n7724 = n1016 & ~n7702;
  assign n7725 = n1016 & n7714;
  assign n7726 = ~n7713 & n7724;
  assign n7727 = ~n7723 & ~n32742;
  assign n7728 = ~n7715 & ~n7727;
  assign n7729 = ~n855 & ~n7728;
  assign n7730 = n855 & ~n7715;
  assign n7731 = ~n7727 & n7730;
  assign n7732 = ~n7242 & ~n32682;
  assign n7733 = ~n7242 & ~n7428;
  assign n7734 = ~n32682 & n7733;
  assign n7735 = ~n7428 & n7732;
  assign n7736 = n7250 & ~n32743;
  assign n7737 = n7254 & n7733;
  assign n7738 = ~n7242 & n7250;
  assign n7739 = ~n32682 & n7738;
  assign n7740 = ~n7428 & n7739;
  assign n7741 = ~n7250 & ~n32743;
  assign n7742 = ~n7740 & ~n7741;
  assign n7743 = ~n7736 & ~n7737;
  assign n7744 = ~n7731 & ~n32744;
  assign n7745 = ~n7729 & ~n7744;
  assign n7746 = ~n720 & ~n7745;
  assign n7747 = ~n7256 & ~n7258;
  assign n7748 = ~n7428 & n7747;
  assign n7749 = ~n32684 & ~n7748;
  assign n7750 = ~n7258 & n32684;
  assign n7751 = ~n7256 & n7750;
  assign n7752 = n32684 & n7748;
  assign n7753 = ~n7428 & n7751;
  assign n7754 = ~n7749 & ~n32745;
  assign n7755 = n720 & ~n7729;
  assign n7756 = n720 & n7745;
  assign n7757 = ~n7744 & n7755;
  assign n7758 = ~n7754 & ~n32746;
  assign n7759 = ~n7746 & ~n7758;
  assign n7760 = ~n592 & ~n7759;
  assign n7761 = ~n7273 & ~n32685;
  assign n7762 = ~n7428 & n7761;
  assign n7763 = ~n32687 & ~n7762;
  assign n7764 = ~n7273 & n32687;
  assign n7765 = ~n32685 & n7764;
  assign n7766 = n32687 & n7762;
  assign n7767 = ~n7428 & n7765;
  assign n7768 = ~n7763 & ~n32747;
  assign n7769 = n592 & ~n7746;
  assign n7770 = ~n7758 & n7769;
  assign n7771 = ~n7768 & ~n7770;
  assign n7772 = ~n7760 & ~n7771;
  assign n7773 = ~n487 & ~n7772;
  assign n7774 = ~n7291 & ~n7293;
  assign n7775 = ~n7428 & n7774;
  assign n7776 = ~n32689 & ~n7775;
  assign n7777 = ~n7293 & n32689;
  assign n7778 = ~n7291 & n7777;
  assign n7779 = n32689 & n7775;
  assign n7780 = ~n7428 & n7778;
  assign n7781 = ~n7776 & ~n32748;
  assign n7782 = n487 & ~n7760;
  assign n7783 = n487 & n7772;
  assign n7784 = ~n7771 & n7782;
  assign n7785 = ~n7781 & ~n32749;
  assign n7786 = ~n7773 & ~n7785;
  assign n7787 = ~n393 & ~n7786;
  assign n7788 = n393 & ~n7773;
  assign n7789 = ~n7785 & n7788;
  assign n7790 = ~n7308 & ~n32691;
  assign n7791 = ~n7308 & ~n7428;
  assign n7792 = ~n32691 & n7791;
  assign n7793 = ~n7428 & n7790;
  assign n7794 = n7316 & ~n32750;
  assign n7795 = n7320 & n7791;
  assign n7796 = ~n7308 & n7316;
  assign n7797 = ~n32691 & n7796;
  assign n7798 = ~n7428 & n7797;
  assign n7799 = ~n7316 & ~n32750;
  assign n7800 = ~n7798 & ~n7799;
  assign n7801 = ~n7794 & ~n7795;
  assign n7802 = ~n7789 & ~n32751;
  assign n7803 = ~n7787 & ~n7802;
  assign n7804 = ~n321 & ~n7803;
  assign n7805 = ~n7322 & ~n7324;
  assign n7806 = ~n7428 & n7805;
  assign n7807 = ~n32693 & ~n7806;
  assign n7808 = ~n7324 & n32693;
  assign n7809 = ~n7322 & n7808;
  assign n7810 = n32693 & n7806;
  assign n7811 = ~n7428 & n7809;
  assign n7812 = ~n7807 & ~n32752;
  assign n7813 = n321 & ~n7787;
  assign n7814 = n321 & n7803;
  assign n7815 = ~n7802 & n7813;
  assign n7816 = ~n7812 & ~n32753;
  assign n7817 = ~n7804 & ~n7816;
  assign n7818 = ~n263 & ~n7817;
  assign n7819 = ~n7339 & ~n32694;
  assign n7820 = ~n7428 & n7819;
  assign n7821 = ~n32696 & ~n7820;
  assign n7822 = ~n7339 & n32696;
  assign n7823 = ~n32694 & n7822;
  assign n7824 = n32696 & n7820;
  assign n7825 = ~n7428 & n7823;
  assign n7826 = ~n7821 & ~n32754;
  assign n7827 = n263 & ~n7804;
  assign n7828 = ~n7816 & n7827;
  assign n7829 = ~n7826 & ~n7828;
  assign n7830 = ~n7818 & ~n7829;
  assign n7831 = ~n214 & ~n7830;
  assign n7832 = ~n7357 & ~n7359;
  assign n7833 = ~n7428 & n7832;
  assign n7834 = ~n32698 & ~n7833;
  assign n7835 = ~n7359 & n32698;
  assign n7836 = ~n7357 & n7835;
  assign n7837 = n32698 & n7833;
  assign n7838 = ~n7428 & n7836;
  assign n7839 = ~n7834 & ~n32755;
  assign n7840 = n214 & ~n7818;
  assign n7841 = n214 & n7830;
  assign n7842 = ~n7829 & n7840;
  assign n7843 = ~n7839 & ~n32756;
  assign n7844 = ~n7831 & ~n7843;
  assign n7845 = ~n197 & ~n7844;
  assign n7846 = n197 & ~n7831;
  assign n7847 = ~n7843 & n7846;
  assign n7848 = ~n7374 & ~n32700;
  assign n7849 = ~n7374 & ~n7428;
  assign n7850 = ~n32700 & n7849;
  assign n7851 = ~n7428 & n7848;
  assign n7852 = n7382 & ~n32757;
  assign n7853 = n7386 & n7849;
  assign n7854 = ~n7374 & n7382;
  assign n7855 = ~n32700 & n7854;
  assign n7856 = ~n7428 & n7855;
  assign n7857 = ~n7382 & ~n32757;
  assign n7858 = ~n7856 & ~n7857;
  assign n7859 = ~n7852 & ~n7853;
  assign n7860 = ~n7847 & ~n32758;
  assign n7861 = ~n7845 & ~n7860;
  assign n7862 = ~n7388 & ~n7390;
  assign n7863 = ~n7428 & n7862;
  assign n7864 = ~n32702 & ~n7863;
  assign n7865 = ~n7390 & n32702;
  assign n7866 = ~n7388 & n7865;
  assign n7867 = n32702 & n7863;
  assign n7868 = ~n7428 & n7866;
  assign n7869 = ~n7864 & ~n32759;
  assign n7870 = ~n7404 & ~n7412;
  assign n7871 = ~n7412 & ~n7428;
  assign n7872 = ~n7404 & n7871;
  assign n7873 = ~n7428 & n7870;
  assign n7874 = ~n32705 & ~n32760;
  assign n7875 = ~n7869 & n7874;
  assign n7876 = ~n7861 & n7875;
  assign n7877 = n193 & ~n7876;
  assign n7878 = ~n7845 & n7869;
  assign n7879 = n7861 & n7869;
  assign n7880 = ~n7860 & n7878;
  assign n7881 = n7404 & ~n7871;
  assign n7882 = ~n193 & ~n7870;
  assign n7883 = ~n7881 & n7882;
  assign n7884 = ~n32761 & ~n7883;
  assign n7885 = ~n7877 & n7884;
  assign n7886 = pi64  & ~n7885;
  assign n7887 = ~pi62  & ~pi63 ;
  assign n7888 = ~pi64  & n7887;
  assign n7889 = ~n7886 & ~n7888;
  assign n7890 = ~n7428 & ~n7889;
  assign n7891 = ~pi64  & ~n7885;
  assign n7892 = pi65  & ~n7891;
  assign n7893 = ~pi65  & n7891;
  assign n7894 = n7430 & ~n7885;
  assign n7895 = ~n7892 & ~n32762;
  assign n7896 = ~n32637 & ~n32706;
  assign n7897 = ~n6916 & n7896;
  assign n7898 = ~n6935 & n7897;
  assign n7899 = ~n32639 & n7898;
  assign n7900 = n6921 & n6937;
  assign n7901 = ~n6929 & n7899;
  assign n7902 = ~n7888 & ~n32763;
  assign n7903 = ~n7426 & n7902;
  assign n7904 = ~n32705 & n7903;
  assign n7905 = ~n7420 & n7904;
  assign n7906 = n7428 & n7889;
  assign n7907 = ~n7886 & n7905;
  assign n7908 = n7895 & ~n32764;
  assign n7909 = ~n7890 & ~n7908;
  assign n7910 = ~n6937 & ~n7909;
  assign n7911 = n6937 & ~n7890;
  assign n7912 = ~n7908 & n7911;
  assign n7913 = ~n7428 & ~n7883;
  assign n7914 = ~n32761 & n7913;
  assign n7915 = ~n7877 & n7914;
  assign n7916 = ~n32762 & ~n7915;
  assign n7917 = pi66  & ~n7916;
  assign n7918 = ~pi66  & ~n7915;
  assign n7919 = ~pi66  & n7916;
  assign n7920 = ~n32762 & n7918;
  assign n7921 = ~n7917 & ~n32765;
  assign n7922 = ~n7912 & ~n7921;
  assign n7923 = ~n7910 & ~n7922;
  assign n7924 = ~n6507 & ~n7923;
  assign n7925 = n6507 & ~n7910;
  assign n7926 = ~n7922 & n7925;
  assign n7927 = n6507 & n7923;
  assign n7928 = ~n7433 & ~n32707;
  assign n7929 = ~n7885 & n7928;
  assign n7930 = n7450 & ~n7929;
  assign n7931 = ~n7450 & n7928;
  assign n7932 = ~n7450 & n7929;
  assign n7933 = ~n7885 & n7931;
  assign n7934 = ~n7930 & ~n32767;
  assign n7935 = ~n32766 & ~n7934;
  assign n7936 = ~n7924 & ~n7935;
  assign n7937 = ~n6051 & ~n7936;
  assign n7938 = n6051 & ~n7924;
  assign n7939 = ~n7935 & n7938;
  assign n7940 = ~n7453 & ~n32710;
  assign n7941 = ~n7453 & ~n7885;
  assign n7942 = ~n32710 & n7941;
  assign n7943 = ~n7885 & n7940;
  assign n7944 = n7462 & ~n32768;
  assign n7945 = n7466 & n7941;
  assign n7946 = n7462 & ~n32710;
  assign n7947 = ~n7453 & n7946;
  assign n7948 = ~n7885 & n7947;
  assign n7949 = ~n7462 & ~n32768;
  assign n7950 = ~n7948 & ~n7949;
  assign n7951 = ~n7944 & ~n7945;
  assign n7952 = ~n7939 & ~n32769;
  assign n7953 = ~n7937 & ~n7952;
  assign n7954 = ~n5648 & ~n7953;
  assign n7955 = n5648 & ~n7937;
  assign n7956 = ~n7952 & n7955;
  assign n7957 = n5648 & n7953;
  assign n7958 = ~n7468 & ~n7470;
  assign n7959 = ~n7885 & n7958;
  assign n7960 = ~n7477 & ~n7959;
  assign n7961 = ~n7468 & n7477;
  assign n7962 = ~n7470 & n7961;
  assign n7963 = n7477 & n7959;
  assign n7964 = ~n7885 & n7962;
  assign n7965 = n7477 & ~n7959;
  assign n7966 = ~n7477 & n7959;
  assign n7967 = ~n7965 & ~n7966;
  assign n7968 = ~n7960 & ~n32771;
  assign n7969 = ~n32770 & n32772;
  assign n7970 = ~n7954 & ~n7969;
  assign n7971 = ~n5223 & ~n7970;
  assign n7972 = n5223 & ~n7954;
  assign n7973 = ~n7969 & n7972;
  assign n7974 = ~n7480 & ~n32713;
  assign n7975 = ~n7480 & ~n7885;
  assign n7976 = ~n32713 & n7975;
  assign n7977 = ~n7885 & n7974;
  assign n7978 = n7488 & ~n32773;
  assign n7979 = n7492 & n7975;
  assign n7980 = n7488 & ~n32713;
  assign n7981 = ~n7480 & n7980;
  assign n7982 = ~n7885 & n7981;
  assign n7983 = ~n7488 & ~n32773;
  assign n7984 = ~n7982 & ~n7983;
  assign n7985 = ~n7978 & ~n7979;
  assign n7986 = ~n7973 & ~n32774;
  assign n7987 = ~n7971 & ~n7986;
  assign n7988 = ~n4851 & ~n7987;
  assign n7989 = n4851 & ~n7971;
  assign n7990 = ~n7986 & n7989;
  assign n7991 = n4851 & n7987;
  assign n7992 = ~n7494 & ~n7496;
  assign n7993 = ~n7885 & n7992;
  assign n7994 = ~n32715 & ~n7993;
  assign n7995 = n32715 & n7993;
  assign n7996 = ~n7494 & ~n32715;
  assign n7997 = ~n7496 & n7996;
  assign n7998 = ~n7885 & n7997;
  assign n7999 = n32715 & ~n7993;
  assign n8000 = ~n7998 & ~n7999;
  assign n8001 = ~n7994 & ~n7995;
  assign n8002 = ~n32775 & ~n32776;
  assign n8003 = ~n7988 & ~n8002;
  assign n8004 = ~n4461 & ~n8003;
  assign n8005 = n4461 & ~n7988;
  assign n8006 = ~n8002 & n8005;
  assign n8007 = ~n7510 & ~n32717;
  assign n8008 = ~n7510 & ~n7885;
  assign n8009 = ~n32717 & n8008;
  assign n8010 = ~n7885 & n8007;
  assign n8011 = n7518 & ~n32777;
  assign n8012 = n7522 & n8008;
  assign n8013 = n7518 & ~n32717;
  assign n8014 = ~n7510 & n8013;
  assign n8015 = ~n7885 & n8014;
  assign n8016 = ~n7518 & ~n32777;
  assign n8017 = ~n8015 & ~n8016;
  assign n8018 = ~n8011 & ~n8012;
  assign n8019 = ~n8006 & ~n32778;
  assign n8020 = ~n8004 & ~n8019;
  assign n8021 = ~n4115 & ~n8020;
  assign n8022 = n4115 & ~n8004;
  assign n8023 = ~n8019 & n8022;
  assign n8024 = n4115 & n8020;
  assign n8025 = ~n7524 & ~n7526;
  assign n8026 = ~n7885 & n8025;
  assign n8027 = ~n32718 & n8026;
  assign n8028 = n32718 & ~n8026;
  assign n8029 = ~n7524 & n32718;
  assign n8030 = ~n7526 & n8029;
  assign n8031 = ~n7885 & n8030;
  assign n8032 = ~n32718 & ~n8026;
  assign n8033 = ~n8031 & ~n8032;
  assign n8034 = ~n8027 & ~n8028;
  assign n8035 = ~n32779 & ~n32780;
  assign n8036 = ~n8021 & ~n8035;
  assign n8037 = ~n3754 & ~n8036;
  assign n8038 = n3754 & ~n8021;
  assign n8039 = ~n8035 & n8038;
  assign n8040 = ~n7539 & ~n32720;
  assign n8041 = ~n7539 & ~n7885;
  assign n8042 = ~n32720 & n8041;
  assign n8043 = ~n7885 & n8040;
  assign n8044 = n7547 & ~n32781;
  assign n8045 = n7551 & n8041;
  assign n8046 = n7547 & ~n32720;
  assign n8047 = ~n7539 & n8046;
  assign n8048 = ~n7885 & n8047;
  assign n8049 = ~n7547 & ~n32781;
  assign n8050 = ~n8048 & ~n8049;
  assign n8051 = ~n8044 & ~n8045;
  assign n8052 = ~n8039 & ~n32782;
  assign n8053 = ~n8037 & ~n8052;
  assign n8054 = ~n3444 & ~n8053;
  assign n8055 = n3444 & ~n8037;
  assign n8056 = ~n8052 & n8055;
  assign n8057 = n3444 & n8053;
  assign n8058 = ~n7553 & ~n7555;
  assign n8059 = ~n7885 & n8058;
  assign n8060 = ~n32721 & n8059;
  assign n8061 = n32721 & ~n8059;
  assign n8062 = ~n32721 & ~n8059;
  assign n8063 = ~n7553 & n32721;
  assign n8064 = ~n7555 & n8063;
  assign n8065 = n32721 & n8059;
  assign n8066 = ~n7885 & n8064;
  assign n8067 = ~n8062 & ~n32784;
  assign n8068 = ~n8060 & ~n8061;
  assign n8069 = ~n32783 & ~n32785;
  assign n8070 = ~n8054 & ~n8069;
  assign n8071 = ~n3116 & ~n8070;
  assign n8072 = n3116 & ~n8054;
  assign n8073 = ~n8069 & n8072;
  assign n8074 = ~n7568 & ~n32723;
  assign n8075 = ~n7568 & ~n7885;
  assign n8076 = ~n32723 & n8075;
  assign n8077 = ~n7885 & n8074;
  assign n8078 = n7576 & ~n32786;
  assign n8079 = n7580 & n8075;
  assign n8080 = n7576 & ~n32723;
  assign n8081 = ~n7568 & n8080;
  assign n8082 = ~n7885 & n8081;
  assign n8083 = ~n7576 & ~n32786;
  assign n8084 = ~n8082 & ~n8083;
  assign n8085 = ~n8078 & ~n8079;
  assign n8086 = ~n8073 & ~n32787;
  assign n8087 = ~n8071 & ~n8086;
  assign n8088 = ~n2833 & ~n8087;
  assign n8089 = n2833 & ~n8071;
  assign n8090 = ~n8086 & n8089;
  assign n8091 = n2833 & n8087;
  assign n8092 = ~n7582 & ~n7584;
  assign n8093 = ~n7582 & ~n7885;
  assign n8094 = ~n7584 & n8093;
  assign n8095 = ~n7885 & n8092;
  assign n8096 = n32725 & ~n32789;
  assign n8097 = n7596 & n8093;
  assign n8098 = ~n32725 & n32789;
  assign n8099 = ~n7582 & n32725;
  assign n8100 = ~n7584 & n8099;
  assign n8101 = ~n7885 & n8100;
  assign n8102 = ~n32725 & ~n32789;
  assign n8103 = ~n8101 & ~n8102;
  assign n8104 = ~n8096 & ~n32790;
  assign n8105 = ~n32788 & ~n32791;
  assign n8106 = ~n8088 & ~n8105;
  assign n8107 = ~n2536 & ~n8106;
  assign n8108 = n2536 & ~n8088;
  assign n8109 = ~n8105 & n8108;
  assign n8110 = ~n7598 & ~n32727;
  assign n8111 = ~n7598 & ~n7885;
  assign n8112 = ~n32727 & n8111;
  assign n8113 = ~n7885 & n8110;
  assign n8114 = n7606 & ~n32792;
  assign n8115 = n7610 & n8111;
  assign n8116 = n7606 & ~n32727;
  assign n8117 = ~n7598 & n8116;
  assign n8118 = ~n7885 & n8117;
  assign n8119 = ~n7606 & ~n32792;
  assign n8120 = ~n8118 & ~n8119;
  assign n8121 = ~n8114 & ~n8115;
  assign n8122 = ~n8109 & ~n32793;
  assign n8123 = ~n8107 & ~n8122;
  assign n8124 = ~n2283 & ~n8123;
  assign n8125 = ~n7612 & ~n7614;
  assign n8126 = ~n7885 & n8125;
  assign n8127 = ~n32730 & ~n8126;
  assign n8128 = ~n7612 & n32730;
  assign n8129 = ~n7614 & n8128;
  assign n8130 = n32730 & n8126;
  assign n8131 = ~n7885 & n8129;
  assign n8132 = ~n8127 & ~n32794;
  assign n8133 = n2283 & ~n8107;
  assign n8134 = ~n8122 & n8133;
  assign n8135 = n2283 & n8123;
  assign n8136 = ~n8132 & ~n32795;
  assign n8137 = ~n8124 & ~n8136;
  assign n8138 = ~n2021 & ~n8137;
  assign n8139 = n2021 & ~n8124;
  assign n8140 = ~n8136 & n8139;
  assign n8141 = ~n7630 & ~n32732;
  assign n8142 = ~n7630 & ~n7885;
  assign n8143 = ~n32732 & n8142;
  assign n8144 = ~n7885 & n8141;
  assign n8145 = n7638 & ~n32796;
  assign n8146 = n7642 & n8142;
  assign n8147 = n7638 & ~n32732;
  assign n8148 = ~n7630 & n8147;
  assign n8149 = ~n7885 & n8148;
  assign n8150 = ~n7638 & ~n32796;
  assign n8151 = ~n8149 & ~n8150;
  assign n8152 = ~n8145 & ~n8146;
  assign n8153 = ~n8140 & ~n32797;
  assign n8154 = ~n8138 & ~n8153;
  assign n8155 = ~n1796 & ~n8154;
  assign n8156 = n1796 & ~n8138;
  assign n8157 = ~n8153 & n8156;
  assign n8158 = n1796 & n8154;
  assign n8159 = ~n7644 & ~n7654;
  assign n8160 = ~n7644 & ~n7885;
  assign n8161 = ~n7654 & n8160;
  assign n8162 = ~n7885 & n8159;
  assign n8163 = n7652 & ~n32799;
  assign n8164 = n7655 & n8160;
  assign n8165 = ~n7644 & n7652;
  assign n8166 = ~n7654 & n8165;
  assign n8167 = ~n7885 & n8166;
  assign n8168 = ~n7652 & ~n32799;
  assign n8169 = ~n8167 & ~n8168;
  assign n8170 = ~n8163 & ~n8164;
  assign n8171 = ~n32798 & ~n32800;
  assign n8172 = ~n8155 & ~n8171;
  assign n8173 = ~n1567 & ~n8172;
  assign n8174 = n1567 & ~n8155;
  assign n8175 = ~n8171 & n8174;
  assign n8176 = ~n7657 & ~n32735;
  assign n8177 = ~n7657 & ~n7885;
  assign n8178 = ~n32735 & n8177;
  assign n8179 = ~n7885 & n8176;
  assign n8180 = n7665 & ~n32801;
  assign n8181 = n7669 & n8177;
  assign n8182 = n7665 & ~n32735;
  assign n8183 = ~n7657 & n8182;
  assign n8184 = ~n7885 & n8183;
  assign n8185 = ~n7665 & ~n32801;
  assign n8186 = ~n8184 & ~n8185;
  assign n8187 = ~n8180 & ~n8181;
  assign n8188 = ~n8175 & ~n32802;
  assign n8189 = ~n8173 & ~n8188;
  assign n8190 = ~n1374 & ~n8189;
  assign n8191 = ~n7671 & ~n7673;
  assign n8192 = ~n7885 & n8191;
  assign n8193 = ~n32737 & ~n8192;
  assign n8194 = ~n7671 & n32737;
  assign n8195 = ~n7673 & n8194;
  assign n8196 = n32737 & n8192;
  assign n8197 = ~n7885 & n8195;
  assign n8198 = ~n8193 & ~n32803;
  assign n8199 = n1374 & ~n8173;
  assign n8200 = ~n8188 & n8199;
  assign n8201 = n1374 & n8189;
  assign n8202 = ~n8198 & ~n32804;
  assign n8203 = ~n8190 & ~n8202;
  assign n8204 = ~n1179 & ~n8203;
  assign n8205 = n1179 & ~n8190;
  assign n8206 = ~n8202 & n8205;
  assign n8207 = ~n7688 & ~n32739;
  assign n8208 = ~n7688 & ~n7885;
  assign n8209 = ~n32739 & n8208;
  assign n8210 = ~n7885 & n8207;
  assign n8211 = n7696 & ~n32805;
  assign n8212 = n7700 & n8208;
  assign n8213 = n7696 & ~n32739;
  assign n8214 = ~n7688 & n8213;
  assign n8215 = ~n7885 & n8214;
  assign n8216 = ~n7696 & ~n32805;
  assign n8217 = ~n8215 & ~n8216;
  assign n8218 = ~n8211 & ~n8212;
  assign n8219 = ~n8206 & ~n32806;
  assign n8220 = ~n8204 & ~n8219;
  assign n8221 = ~n1016 & ~n8220;
  assign n8222 = n1016 & ~n8204;
  assign n8223 = ~n8219 & n8222;
  assign n8224 = n1016 & n8220;
  assign n8225 = ~n7702 & ~n7712;
  assign n8226 = ~n7702 & ~n7885;
  assign n8227 = ~n7712 & n8226;
  assign n8228 = ~n7885 & n8225;
  assign n8229 = n7710 & ~n32808;
  assign n8230 = n7713 & n8226;
  assign n8231 = ~n7702 & n7710;
  assign n8232 = ~n7712 & n8231;
  assign n8233 = ~n7885 & n8232;
  assign n8234 = ~n7710 & ~n32808;
  assign n8235 = ~n8233 & ~n8234;
  assign n8236 = ~n8229 & ~n8230;
  assign n8237 = ~n32807 & ~n32809;
  assign n8238 = ~n8221 & ~n8237;
  assign n8239 = ~n855 & ~n8238;
  assign n8240 = n855 & ~n8221;
  assign n8241 = ~n8237 & n8240;
  assign n8242 = ~n7715 & ~n32742;
  assign n8243 = ~n7715 & ~n7885;
  assign n8244 = ~n32742 & n8243;
  assign n8245 = ~n7885 & n8242;
  assign n8246 = n7723 & ~n32810;
  assign n8247 = n7727 & n8243;
  assign n8248 = n7723 & ~n32742;
  assign n8249 = ~n7715 & n8248;
  assign n8250 = ~n7885 & n8249;
  assign n8251 = ~n7723 & ~n32810;
  assign n8252 = ~n8250 & ~n8251;
  assign n8253 = ~n8246 & ~n8247;
  assign n8254 = ~n8241 & ~n32811;
  assign n8255 = ~n8239 & ~n8254;
  assign n8256 = ~n720 & ~n8255;
  assign n8257 = ~n7729 & ~n7731;
  assign n8258 = ~n7885 & n8257;
  assign n8259 = ~n32744 & ~n8258;
  assign n8260 = ~n7729 & n32744;
  assign n8261 = ~n7731 & n8260;
  assign n8262 = n32744 & n8258;
  assign n8263 = ~n7885 & n8261;
  assign n8264 = ~n8259 & ~n32812;
  assign n8265 = n720 & ~n8239;
  assign n8266 = ~n8254 & n8265;
  assign n8267 = n720 & n8255;
  assign n8268 = ~n8264 & ~n32813;
  assign n8269 = ~n8256 & ~n8268;
  assign n8270 = ~n592 & ~n8269;
  assign n8271 = n592 & ~n8256;
  assign n8272 = ~n8268 & n8271;
  assign n8273 = ~n7746 & ~n32746;
  assign n8274 = ~n7746 & ~n7885;
  assign n8275 = ~n32746 & n8274;
  assign n8276 = ~n7885 & n8273;
  assign n8277 = n7754 & ~n32814;
  assign n8278 = n7758 & n8274;
  assign n8279 = n7754 & ~n32746;
  assign n8280 = ~n7746 & n8279;
  assign n8281 = ~n7885 & n8280;
  assign n8282 = ~n7754 & ~n32814;
  assign n8283 = ~n8281 & ~n8282;
  assign n8284 = ~n8277 & ~n8278;
  assign n8285 = ~n8272 & ~n32815;
  assign n8286 = ~n8270 & ~n8285;
  assign n8287 = ~n487 & ~n8286;
  assign n8288 = n487 & ~n8270;
  assign n8289 = ~n8285 & n8288;
  assign n8290 = n487 & n8286;
  assign n8291 = ~n7760 & ~n7770;
  assign n8292 = ~n7760 & ~n7885;
  assign n8293 = ~n7770 & n8292;
  assign n8294 = ~n7885 & n8291;
  assign n8295 = n7768 & ~n32817;
  assign n8296 = n7771 & n8292;
  assign n8297 = ~n7760 & n7768;
  assign n8298 = ~n7770 & n8297;
  assign n8299 = ~n7885 & n8298;
  assign n8300 = ~n7768 & ~n32817;
  assign n8301 = ~n8299 & ~n8300;
  assign n8302 = ~n8295 & ~n8296;
  assign n8303 = ~n32816 & ~n32818;
  assign n8304 = ~n8287 & ~n8303;
  assign n8305 = ~n393 & ~n8304;
  assign n8306 = n393 & ~n8287;
  assign n8307 = ~n8303 & n8306;
  assign n8308 = ~n7773 & ~n32749;
  assign n8309 = ~n7773 & ~n7885;
  assign n8310 = ~n32749 & n8309;
  assign n8311 = ~n7885 & n8308;
  assign n8312 = n7781 & ~n32819;
  assign n8313 = n7785 & n8309;
  assign n8314 = n7781 & ~n32749;
  assign n8315 = ~n7773 & n8314;
  assign n8316 = ~n7885 & n8315;
  assign n8317 = ~n7781 & ~n32819;
  assign n8318 = ~n8316 & ~n8317;
  assign n8319 = ~n8312 & ~n8313;
  assign n8320 = ~n8307 & ~n32820;
  assign n8321 = ~n8305 & ~n8320;
  assign n8322 = ~n321 & ~n8321;
  assign n8323 = ~n7787 & ~n7789;
  assign n8324 = ~n7885 & n8323;
  assign n8325 = ~n32751 & ~n8324;
  assign n8326 = ~n7787 & n32751;
  assign n8327 = ~n7789 & n8326;
  assign n8328 = n32751 & n8324;
  assign n8329 = ~n7885 & n8327;
  assign n8330 = ~n8325 & ~n32821;
  assign n8331 = n321 & ~n8305;
  assign n8332 = ~n8320 & n8331;
  assign n8333 = n321 & n8321;
  assign n8334 = ~n8330 & ~n32822;
  assign n8335 = ~n8322 & ~n8334;
  assign n8336 = ~n263 & ~n8335;
  assign n8337 = n263 & ~n8322;
  assign n8338 = ~n8334 & n8337;
  assign n8339 = ~n7804 & ~n32753;
  assign n8340 = ~n7804 & ~n7885;
  assign n8341 = ~n32753 & n8340;
  assign n8342 = ~n7885 & n8339;
  assign n8343 = n7812 & ~n32823;
  assign n8344 = n7816 & n8340;
  assign n8345 = n7812 & ~n32753;
  assign n8346 = ~n7804 & n8345;
  assign n8347 = ~n7885 & n8346;
  assign n8348 = ~n7812 & ~n32823;
  assign n8349 = ~n8347 & ~n8348;
  assign n8350 = ~n8343 & ~n8344;
  assign n8351 = ~n8338 & ~n32824;
  assign n8352 = ~n8336 & ~n8351;
  assign n8353 = ~n214 & ~n8352;
  assign n8354 = n214 & ~n8336;
  assign n8355 = ~n8351 & n8354;
  assign n8356 = n214 & n8352;
  assign n8357 = ~n7818 & ~n7828;
  assign n8358 = ~n7818 & ~n7885;
  assign n8359 = ~n7828 & n8358;
  assign n8360 = ~n7885 & n8357;
  assign n8361 = n7826 & ~n32826;
  assign n8362 = n7829 & n8358;
  assign n8363 = ~n7818 & n7826;
  assign n8364 = ~n7828 & n8363;
  assign n8365 = ~n7885 & n8364;
  assign n8366 = ~n7826 & ~n32826;
  assign n8367 = ~n8365 & ~n8366;
  assign n8368 = ~n8361 & ~n8362;
  assign n8369 = ~n32825 & ~n32827;
  assign n8370 = ~n8353 & ~n8369;
  assign n8371 = ~n197 & ~n8370;
  assign n8372 = n197 & ~n8353;
  assign n8373 = ~n8369 & n8372;
  assign n8374 = ~n7831 & ~n32756;
  assign n8375 = ~n7831 & ~n7885;
  assign n8376 = ~n32756 & n8375;
  assign n8377 = ~n7885 & n8374;
  assign n8378 = n7839 & ~n32828;
  assign n8379 = n7843 & n8375;
  assign n8380 = n7839 & ~n32756;
  assign n8381 = ~n7831 & n8380;
  assign n8382 = ~n7885 & n8381;
  assign n8383 = ~n7839 & ~n32828;
  assign n8384 = ~n8382 & ~n8383;
  assign n8385 = ~n8378 & ~n8379;
  assign n8386 = ~n8373 & ~n32829;
  assign n8387 = ~n8371 & ~n8386;
  assign n8388 = ~n7845 & ~n7847;
  assign n8389 = ~n7885 & n8388;
  assign n8390 = ~n32758 & ~n8389;
  assign n8391 = ~n7845 & n32758;
  assign n8392 = ~n7847 & n8391;
  assign n8393 = n32758 & n8389;
  assign n8394 = ~n7885 & n8392;
  assign n8395 = ~n8390 & ~n32830;
  assign n8396 = ~n7861 & ~n7869;
  assign n8397 = ~n7869 & ~n7885;
  assign n8398 = ~n7861 & n8397;
  assign n8399 = ~n7885 & n8396;
  assign n8400 = ~n32761 & ~n32831;
  assign n8401 = ~n8395 & n8400;
  assign n8402 = ~n8387 & n8401;
  assign n8403 = n193 & ~n8402;
  assign n8404 = ~n8371 & n8395;
  assign n8405 = ~n8386 & n8404;
  assign n8406 = n8387 & n8395;
  assign n8407 = n7861 & ~n8397;
  assign n8408 = ~n193 & ~n8396;
  assign n8409 = ~n8407 & n8408;
  assign n8410 = ~n32832 & ~n8409;
  assign n8411 = ~n8403 & n8410;
  assign n8412 = pi62  & ~n8411;
  assign n8413 = ~pi60  & ~pi61 ;
  assign n8414 = ~pi62  & n8413;
  assign n8415 = ~n8412 & ~n8414;
  assign n8416 = ~n7885 & ~n8415;
  assign n8417 = ~pi62  & ~n8411;
  assign n8418 = ~pi63  & n8417;
  assign n8419 = n7887 & ~n8411;
  assign n8420 = pi63  & ~n8417;
  assign n8421 = ~n32833 & ~n8420;
  assign n8422 = ~n32703 & ~n32763;
  assign n8423 = ~n7407 & n8422;
  assign n8424 = ~n7426 & n8423;
  assign n8425 = ~n32705 & n8424;
  assign n8426 = n7412 & n7428;
  assign n8427 = ~n7420 & n8425;
  assign n8428 = ~n8414 & ~n32834;
  assign n8429 = ~n7883 & n8428;
  assign n8430 = ~n32761 & n8429;
  assign n8431 = ~n7877 & n8430;
  assign n8432 = n7885 & n8415;
  assign n8433 = ~n8412 & n8431;
  assign n8434 = n8421 & ~n32835;
  assign n8435 = ~n8416 & ~n8434;
  assign n8436 = ~n7428 & ~n8435;
  assign n8437 = ~n7885 & ~n8409;
  assign n8438 = ~n32832 & n8437;
  assign n8439 = ~n8403 & n8438;
  assign n8440 = ~n32833 & ~n8439;
  assign n8441 = pi64  & ~n8440;
  assign n8442 = ~pi64  & ~n8439;
  assign n8443 = ~pi64  & n8440;
  assign n8444 = ~n32833 & n8442;
  assign n8445 = ~n8441 & ~n32836;
  assign n8446 = n7428 & ~n8416;
  assign n8447 = n7428 & n8435;
  assign n8448 = ~n8434 & n8446;
  assign n8449 = ~n8445 & ~n32837;
  assign n8450 = ~n8436 & ~n8449;
  assign n8451 = ~n6937 & ~n8450;
  assign n8452 = n6937 & ~n8436;
  assign n8453 = ~n8449 & n8452;
  assign n8454 = ~n7890 & ~n32764;
  assign n8455 = ~n8411 & n8454;
  assign n8456 = n7895 & ~n8455;
  assign n8457 = ~n7895 & ~n32764;
  assign n8458 = ~n7890 & n8457;
  assign n8459 = ~n7895 & n8455;
  assign n8460 = ~n8411 & n8458;
  assign n8461 = ~n8456 & ~n32838;
  assign n8462 = ~n8453 & ~n8461;
  assign n8463 = ~n8451 & ~n8462;
  assign n8464 = ~n6507 & ~n8463;
  assign n8465 = ~n7910 & ~n7912;
  assign n8466 = ~n8411 & n8465;
  assign n8467 = ~n7921 & ~n8466;
  assign n8468 = ~n7912 & n7921;
  assign n8469 = ~n7910 & n8468;
  assign n8470 = n7921 & n8466;
  assign n8471 = ~n8411 & n8469;
  assign n8472 = ~n8467 & ~n32839;
  assign n8473 = n6507 & ~n8451;
  assign n8474 = n6507 & n8463;
  assign n8475 = ~n8462 & n8473;
  assign n8476 = ~n8472 & ~n32840;
  assign n8477 = ~n8464 & ~n8476;
  assign n8478 = ~n6051 & ~n8477;
  assign n8479 = n6051 & ~n8464;
  assign n8480 = ~n8476 & n8479;
  assign n8481 = ~n7924 & ~n32766;
  assign n8482 = ~n8411 & n8481;
  assign n8483 = ~n7934 & ~n8482;
  assign n8484 = ~n7924 & n7934;
  assign n8485 = ~n32766 & n8484;
  assign n8486 = n7934 & n8482;
  assign n8487 = ~n8411 & n8485;
  assign n8488 = n7934 & ~n8482;
  assign n8489 = ~n7934 & n8482;
  assign n8490 = ~n8488 & ~n8489;
  assign n8491 = ~n8483 & ~n32841;
  assign n8492 = ~n8480 & n32842;
  assign n8493 = ~n8478 & ~n8492;
  assign n8494 = ~n5648 & ~n8493;
  assign n8495 = ~n7937 & ~n7939;
  assign n8496 = ~n8411 & n8495;
  assign n8497 = ~n32769 & ~n8496;
  assign n8498 = ~n7939 & n32769;
  assign n8499 = ~n7937 & n8498;
  assign n8500 = n32769 & n8496;
  assign n8501 = ~n8411 & n8499;
  assign n8502 = ~n8497 & ~n32843;
  assign n8503 = n5648 & ~n8478;
  assign n8504 = n5648 & n8493;
  assign n8505 = ~n8492 & n8503;
  assign n8506 = ~n8502 & ~n32844;
  assign n8507 = ~n8494 & ~n8506;
  assign n8508 = ~n5223 & ~n8507;
  assign n8509 = n5223 & ~n8494;
  assign n8510 = ~n8506 & n8509;
  assign n8511 = ~n7954 & ~n32770;
  assign n8512 = ~n8411 & n8511;
  assign n8513 = ~n32772 & ~n8512;
  assign n8514 = n32772 & n8512;
  assign n8515 = ~n7954 & ~n32772;
  assign n8516 = ~n32770 & n8515;
  assign n8517 = ~n8411 & n8516;
  assign n8518 = n32772 & ~n8512;
  assign n8519 = ~n8517 & ~n8518;
  assign n8520 = ~n8513 & ~n8514;
  assign n8521 = ~n8510 & ~n32845;
  assign n8522 = ~n8508 & ~n8521;
  assign n8523 = ~n4851 & ~n8522;
  assign n8524 = ~n7971 & ~n7973;
  assign n8525 = ~n8411 & n8524;
  assign n8526 = ~n32774 & ~n8525;
  assign n8527 = ~n7973 & n32774;
  assign n8528 = ~n7971 & n8527;
  assign n8529 = n32774 & n8525;
  assign n8530 = ~n8411 & n8528;
  assign n8531 = ~n8526 & ~n32846;
  assign n8532 = n4851 & ~n8508;
  assign n8533 = n4851 & n8522;
  assign n8534 = ~n8521 & n8532;
  assign n8535 = ~n8531 & ~n32847;
  assign n8536 = ~n8523 & ~n8535;
  assign n8537 = ~n4461 & ~n8536;
  assign n8538 = n4461 & ~n8523;
  assign n8539 = ~n8535 & n8538;
  assign n8540 = ~n7988 & ~n32775;
  assign n8541 = ~n8411 & n8540;
  assign n8542 = ~n32776 & n8541;
  assign n8543 = n32776 & ~n8541;
  assign n8544 = ~n7988 & n32776;
  assign n8545 = ~n32775 & n8544;
  assign n8546 = ~n8411 & n8545;
  assign n8547 = ~n32776 & ~n8541;
  assign n8548 = ~n8546 & ~n8547;
  assign n8549 = ~n8542 & ~n8543;
  assign n8550 = ~n8539 & ~n32848;
  assign n8551 = ~n8537 & ~n8550;
  assign n8552 = ~n4115 & ~n8551;
  assign n8553 = ~n8004 & ~n8006;
  assign n8554 = ~n8411 & n8553;
  assign n8555 = ~n32778 & ~n8554;
  assign n8556 = ~n8006 & n32778;
  assign n8557 = ~n8004 & n8556;
  assign n8558 = n32778 & n8554;
  assign n8559 = ~n8411 & n8557;
  assign n8560 = ~n8555 & ~n32849;
  assign n8561 = n4115 & ~n8537;
  assign n8562 = n4115 & n8551;
  assign n8563 = ~n8550 & n8561;
  assign n8564 = ~n8560 & ~n32850;
  assign n8565 = ~n8552 & ~n8564;
  assign n8566 = ~n3754 & ~n8565;
  assign n8567 = n3754 & ~n8552;
  assign n8568 = ~n8564 & n8567;
  assign n8569 = ~n8021 & ~n32779;
  assign n8570 = ~n8411 & n8569;
  assign n8571 = ~n32780 & n8570;
  assign n8572 = n32780 & ~n8570;
  assign n8573 = ~n32780 & ~n8570;
  assign n8574 = ~n8021 & n32780;
  assign n8575 = ~n32779 & n8574;
  assign n8576 = n32780 & n8570;
  assign n8577 = ~n8411 & n8575;
  assign n8578 = ~n8573 & ~n32851;
  assign n8579 = ~n8571 & ~n8572;
  assign n8580 = ~n8568 & ~n32852;
  assign n8581 = ~n8566 & ~n8580;
  assign n8582 = ~n3444 & ~n8581;
  assign n8583 = ~n8037 & ~n8039;
  assign n8584 = ~n8411 & n8583;
  assign n8585 = ~n32782 & ~n8584;
  assign n8586 = ~n8039 & n32782;
  assign n8587 = ~n8037 & n8586;
  assign n8588 = n32782 & n8584;
  assign n8589 = ~n8411 & n8587;
  assign n8590 = ~n8585 & ~n32853;
  assign n8591 = n3444 & ~n8566;
  assign n8592 = n3444 & n8581;
  assign n8593 = ~n8580 & n8591;
  assign n8594 = ~n8590 & ~n32854;
  assign n8595 = ~n8582 & ~n8594;
  assign n8596 = ~n3116 & ~n8595;
  assign n8597 = n3116 & ~n8582;
  assign n8598 = ~n8594 & n8597;
  assign n8599 = ~n8054 & ~n32783;
  assign n8600 = ~n8054 & ~n8411;
  assign n8601 = ~n32783 & n8600;
  assign n8602 = ~n8411 & n8599;
  assign n8603 = n32785 & ~n32855;
  assign n8604 = n8069 & n8600;
  assign n8605 = ~n32785 & n32855;
  assign n8606 = ~n8054 & n32785;
  assign n8607 = ~n32783 & n8606;
  assign n8608 = ~n8411 & n8607;
  assign n8609 = ~n32785 & ~n32855;
  assign n8610 = ~n8608 & ~n8609;
  assign n8611 = ~n8603 & ~n32856;
  assign n8612 = ~n8598 & ~n32857;
  assign n8613 = ~n8596 & ~n8612;
  assign n8614 = ~n2833 & ~n8613;
  assign n8615 = ~n8071 & ~n8073;
  assign n8616 = ~n8411 & n8615;
  assign n8617 = ~n32787 & ~n8616;
  assign n8618 = ~n8073 & n32787;
  assign n8619 = ~n8071 & n8618;
  assign n8620 = n32787 & n8616;
  assign n8621 = ~n8411 & n8619;
  assign n8622 = ~n8617 & ~n32858;
  assign n8623 = n2833 & ~n8596;
  assign n8624 = n2833 & n8613;
  assign n8625 = ~n8612 & n8623;
  assign n8626 = ~n8622 & ~n32859;
  assign n8627 = ~n8614 & ~n8626;
  assign n8628 = ~n2536 & ~n8627;
  assign n8629 = ~n8088 & ~n32788;
  assign n8630 = ~n8411 & n8629;
  assign n8631 = ~n32791 & ~n8630;
  assign n8632 = ~n8088 & n32791;
  assign n8633 = ~n32788 & n8632;
  assign n8634 = n32791 & n8630;
  assign n8635 = ~n8411 & n8633;
  assign n8636 = ~n8631 & ~n32860;
  assign n8637 = n2536 & ~n8614;
  assign n8638 = ~n8626 & n8637;
  assign n8639 = ~n8636 & ~n8638;
  assign n8640 = ~n8628 & ~n8639;
  assign n8641 = ~n2283 & ~n8640;
  assign n8642 = ~n8107 & ~n8109;
  assign n8643 = ~n8411 & n8642;
  assign n8644 = ~n32793 & ~n8643;
  assign n8645 = ~n8109 & n32793;
  assign n8646 = ~n8107 & n8645;
  assign n8647 = n32793 & n8643;
  assign n8648 = ~n8411 & n8646;
  assign n8649 = ~n8644 & ~n32861;
  assign n8650 = n2283 & ~n8628;
  assign n8651 = n2283 & n8640;
  assign n8652 = ~n8639 & n8650;
  assign n8653 = ~n8649 & ~n32862;
  assign n8654 = ~n8641 & ~n8653;
  assign n8655 = ~n2021 & ~n8654;
  assign n8656 = n2021 & ~n8641;
  assign n8657 = ~n8653 & n8656;
  assign n8658 = ~n8124 & ~n32795;
  assign n8659 = ~n8124 & ~n8411;
  assign n8660 = ~n32795 & n8659;
  assign n8661 = ~n8411 & n8658;
  assign n8662 = n8132 & ~n32863;
  assign n8663 = n8136 & n8659;
  assign n8664 = ~n8124 & n8132;
  assign n8665 = ~n32795 & n8664;
  assign n8666 = ~n8411 & n8665;
  assign n8667 = ~n8132 & ~n32863;
  assign n8668 = ~n8666 & ~n8667;
  assign n8669 = ~n8662 & ~n8663;
  assign n8670 = ~n8657 & ~n32864;
  assign n8671 = ~n8655 & ~n8670;
  assign n8672 = ~n1796 & ~n8671;
  assign n8673 = ~n8138 & ~n8140;
  assign n8674 = ~n8411 & n8673;
  assign n8675 = ~n32797 & ~n8674;
  assign n8676 = ~n8140 & n32797;
  assign n8677 = ~n8138 & n8676;
  assign n8678 = n32797 & n8674;
  assign n8679 = ~n8411 & n8677;
  assign n8680 = ~n8675 & ~n32865;
  assign n8681 = n1796 & ~n8655;
  assign n8682 = n1796 & n8671;
  assign n8683 = ~n8670 & n8681;
  assign n8684 = ~n8680 & ~n32866;
  assign n8685 = ~n8672 & ~n8684;
  assign n8686 = ~n1567 & ~n8685;
  assign n8687 = ~n8155 & ~n32798;
  assign n8688 = ~n8411 & n8687;
  assign n8689 = ~n32800 & ~n8688;
  assign n8690 = ~n8155 & n32800;
  assign n8691 = ~n32798 & n8690;
  assign n8692 = n32800 & n8688;
  assign n8693 = ~n8411 & n8691;
  assign n8694 = ~n8689 & ~n32867;
  assign n8695 = n1567 & ~n8672;
  assign n8696 = ~n8684 & n8695;
  assign n8697 = ~n8694 & ~n8696;
  assign n8698 = ~n8686 & ~n8697;
  assign n8699 = ~n1374 & ~n8698;
  assign n8700 = ~n8173 & ~n8175;
  assign n8701 = ~n8411 & n8700;
  assign n8702 = ~n32802 & ~n8701;
  assign n8703 = ~n8175 & n32802;
  assign n8704 = ~n8173 & n8703;
  assign n8705 = n32802 & n8701;
  assign n8706 = ~n8411 & n8704;
  assign n8707 = ~n8702 & ~n32868;
  assign n8708 = n1374 & ~n8686;
  assign n8709 = n1374 & n8698;
  assign n8710 = ~n8697 & n8708;
  assign n8711 = ~n8707 & ~n32869;
  assign n8712 = ~n8699 & ~n8711;
  assign n8713 = ~n1179 & ~n8712;
  assign n8714 = n1179 & ~n8699;
  assign n8715 = ~n8711 & n8714;
  assign n8716 = ~n8190 & ~n32804;
  assign n8717 = ~n8190 & ~n8411;
  assign n8718 = ~n32804 & n8717;
  assign n8719 = ~n8411 & n8716;
  assign n8720 = n8198 & ~n32870;
  assign n8721 = n8202 & n8717;
  assign n8722 = ~n8190 & n8198;
  assign n8723 = ~n32804 & n8722;
  assign n8724 = ~n8411 & n8723;
  assign n8725 = ~n8198 & ~n32870;
  assign n8726 = ~n8724 & ~n8725;
  assign n8727 = ~n8720 & ~n8721;
  assign n8728 = ~n8715 & ~n32871;
  assign n8729 = ~n8713 & ~n8728;
  assign n8730 = ~n1016 & ~n8729;
  assign n8731 = ~n8204 & ~n8206;
  assign n8732 = ~n8411 & n8731;
  assign n8733 = ~n32806 & ~n8732;
  assign n8734 = ~n8206 & n32806;
  assign n8735 = ~n8204 & n8734;
  assign n8736 = n32806 & n8732;
  assign n8737 = ~n8411 & n8735;
  assign n8738 = ~n8733 & ~n32872;
  assign n8739 = n1016 & ~n8713;
  assign n8740 = n1016 & n8729;
  assign n8741 = ~n8728 & n8739;
  assign n8742 = ~n8738 & ~n32873;
  assign n8743 = ~n8730 & ~n8742;
  assign n8744 = ~n855 & ~n8743;
  assign n8745 = ~n8221 & ~n32807;
  assign n8746 = ~n8411 & n8745;
  assign n8747 = ~n32809 & ~n8746;
  assign n8748 = ~n8221 & n32809;
  assign n8749 = ~n32807 & n8748;
  assign n8750 = n32809 & n8746;
  assign n8751 = ~n8411 & n8749;
  assign n8752 = ~n8747 & ~n32874;
  assign n8753 = n855 & ~n8730;
  assign n8754 = ~n8742 & n8753;
  assign n8755 = ~n8752 & ~n8754;
  assign n8756 = ~n8744 & ~n8755;
  assign n8757 = ~n720 & ~n8756;
  assign n8758 = ~n8239 & ~n8241;
  assign n8759 = ~n8411 & n8758;
  assign n8760 = ~n32811 & ~n8759;
  assign n8761 = ~n8241 & n32811;
  assign n8762 = ~n8239 & n8761;
  assign n8763 = n32811 & n8759;
  assign n8764 = ~n8411 & n8762;
  assign n8765 = ~n8760 & ~n32875;
  assign n8766 = n720 & ~n8744;
  assign n8767 = n720 & n8756;
  assign n8768 = ~n8755 & n8766;
  assign n8769 = ~n8765 & ~n32876;
  assign n8770 = ~n8757 & ~n8769;
  assign n8771 = ~n592 & ~n8770;
  assign n8772 = n592 & ~n8757;
  assign n8773 = ~n8769 & n8772;
  assign n8774 = ~n8256 & ~n32813;
  assign n8775 = ~n8256 & ~n8411;
  assign n8776 = ~n32813 & n8775;
  assign n8777 = ~n8411 & n8774;
  assign n8778 = n8264 & ~n32877;
  assign n8779 = n8268 & n8775;
  assign n8780 = ~n8256 & n8264;
  assign n8781 = ~n32813 & n8780;
  assign n8782 = ~n8411 & n8781;
  assign n8783 = ~n8264 & ~n32877;
  assign n8784 = ~n8782 & ~n8783;
  assign n8785 = ~n8778 & ~n8779;
  assign n8786 = ~n8773 & ~n32878;
  assign n8787 = ~n8771 & ~n8786;
  assign n8788 = ~n487 & ~n8787;
  assign n8789 = ~n8270 & ~n8272;
  assign n8790 = ~n8411 & n8789;
  assign n8791 = ~n32815 & ~n8790;
  assign n8792 = ~n8272 & n32815;
  assign n8793 = ~n8270 & n8792;
  assign n8794 = n32815 & n8790;
  assign n8795 = ~n8411 & n8793;
  assign n8796 = ~n8791 & ~n32879;
  assign n8797 = n487 & ~n8771;
  assign n8798 = n487 & n8787;
  assign n8799 = ~n8786 & n8797;
  assign n8800 = ~n8796 & ~n32880;
  assign n8801 = ~n8788 & ~n8800;
  assign n8802 = ~n393 & ~n8801;
  assign n8803 = ~n8287 & ~n32816;
  assign n8804 = ~n8411 & n8803;
  assign n8805 = ~n32818 & ~n8804;
  assign n8806 = ~n8287 & n32818;
  assign n8807 = ~n32816 & n8806;
  assign n8808 = n32818 & n8804;
  assign n8809 = ~n8411 & n8807;
  assign n8810 = ~n8805 & ~n32881;
  assign n8811 = n393 & ~n8788;
  assign n8812 = ~n8800 & n8811;
  assign n8813 = ~n8810 & ~n8812;
  assign n8814 = ~n8802 & ~n8813;
  assign n8815 = ~n321 & ~n8814;
  assign n8816 = ~n8305 & ~n8307;
  assign n8817 = ~n8411 & n8816;
  assign n8818 = ~n32820 & ~n8817;
  assign n8819 = ~n8307 & n32820;
  assign n8820 = ~n8305 & n8819;
  assign n8821 = n32820 & n8817;
  assign n8822 = ~n8411 & n8820;
  assign n8823 = ~n8818 & ~n32882;
  assign n8824 = n321 & ~n8802;
  assign n8825 = n321 & n8814;
  assign n8826 = ~n8813 & n8824;
  assign n8827 = ~n8823 & ~n32883;
  assign n8828 = ~n8815 & ~n8827;
  assign n8829 = ~n263 & ~n8828;
  assign n8830 = n263 & ~n8815;
  assign n8831 = ~n8827 & n8830;
  assign n8832 = ~n8322 & ~n32822;
  assign n8833 = ~n8322 & ~n8411;
  assign n8834 = ~n32822 & n8833;
  assign n8835 = ~n8411 & n8832;
  assign n8836 = n8330 & ~n32884;
  assign n8837 = n8334 & n8833;
  assign n8838 = ~n8322 & n8330;
  assign n8839 = ~n32822 & n8838;
  assign n8840 = ~n8411 & n8839;
  assign n8841 = ~n8330 & ~n32884;
  assign n8842 = ~n8840 & ~n8841;
  assign n8843 = ~n8836 & ~n8837;
  assign n8844 = ~n8831 & ~n32885;
  assign n8845 = ~n8829 & ~n8844;
  assign n8846 = ~n214 & ~n8845;
  assign n8847 = ~n8336 & ~n8338;
  assign n8848 = ~n8411 & n8847;
  assign n8849 = ~n32824 & ~n8848;
  assign n8850 = ~n8338 & n32824;
  assign n8851 = ~n8336 & n8850;
  assign n8852 = n32824 & n8848;
  assign n8853 = ~n8411 & n8851;
  assign n8854 = ~n8849 & ~n32886;
  assign n8855 = n214 & ~n8829;
  assign n8856 = n214 & n8845;
  assign n8857 = ~n8844 & n8855;
  assign n8858 = ~n8854 & ~n32887;
  assign n8859 = ~n8846 & ~n8858;
  assign n8860 = ~n197 & ~n8859;
  assign n8861 = ~n8353 & ~n32825;
  assign n8862 = ~n8411 & n8861;
  assign n8863 = ~n32827 & ~n8862;
  assign n8864 = ~n8353 & n32827;
  assign n8865 = ~n32825 & n8864;
  assign n8866 = n32827 & n8862;
  assign n8867 = ~n8411 & n8865;
  assign n8868 = ~n8863 & ~n32888;
  assign n8869 = n197 & ~n8846;
  assign n8870 = ~n8858 & n8869;
  assign n8871 = ~n8868 & ~n8870;
  assign n8872 = ~n8860 & ~n8871;
  assign n8873 = ~n8371 & ~n8373;
  assign n8874 = ~n8411 & n8873;
  assign n8875 = ~n32829 & ~n8874;
  assign n8876 = ~n8373 & n32829;
  assign n8877 = ~n8371 & n8876;
  assign n8878 = n32829 & n8874;
  assign n8879 = ~n8411 & n8877;
  assign n8880 = ~n8875 & ~n32889;
  assign n8881 = ~n8387 & ~n8395;
  assign n8882 = ~n8395 & ~n8411;
  assign n8883 = ~n8387 & n8882;
  assign n8884 = ~n8411 & n8881;
  assign n8885 = ~n32832 & ~n32890;
  assign n8886 = ~n8880 & n8885;
  assign n8887 = ~n8872 & n8886;
  assign n8888 = n193 & ~n8887;
  assign n8889 = ~n8860 & n8880;
  assign n8890 = n8872 & n8880;
  assign n8891 = ~n8871 & n8889;
  assign n8892 = n8387 & ~n8882;
  assign n8893 = ~n193 & ~n8881;
  assign n8894 = ~n8892 & n8893;
  assign n8895 = ~n32891 & ~n8894;
  assign n8896 = ~n8888 & n8895;
  assign n8897 = pi60  & ~n8896;
  assign n8898 = ~pi58  & ~pi59 ;
  assign n8899 = ~pi60  & n8898;
  assign n8900 = ~n8897 & ~n8899;
  assign n8901 = ~n8411 & ~n8900;
  assign n8902 = ~pi60  & ~n8896;
  assign n8903 = pi61  & ~n8902;
  assign n8904 = ~pi61  & n8902;
  assign n8905 = n8413 & ~n8896;
  assign n8906 = ~n8903 & ~n32892;
  assign n8907 = ~n32759 & ~n32834;
  assign n8908 = ~n7864 & n8907;
  assign n8909 = ~n7883 & n8908;
  assign n8910 = ~n32761 & n8909;
  assign n8911 = n7869 & n7885;
  assign n8912 = ~n7877 & n8910;
  assign n8913 = ~n8899 & ~n32893;
  assign n8914 = ~n8409 & n8913;
  assign n8915 = ~n32832 & n8914;
  assign n8916 = ~n8403 & n8915;
  assign n8917 = n8411 & n8900;
  assign n8918 = ~n8897 & n8916;
  assign n8919 = n8906 & ~n32894;
  assign n8920 = ~n8901 & ~n8919;
  assign n8921 = ~n7885 & ~n8920;
  assign n8922 = n7885 & ~n8901;
  assign n8923 = ~n8919 & n8922;
  assign n8924 = ~n8411 & ~n8894;
  assign n8925 = ~n32891 & n8924;
  assign n8926 = ~n8888 & n8925;
  assign n8927 = ~n32892 & ~n8926;
  assign n8928 = pi62  & ~n8927;
  assign n8929 = ~pi62  & ~n8926;
  assign n8930 = ~pi62  & n8927;
  assign n8931 = ~n32892 & n8929;
  assign n8932 = ~n8928 & ~n32895;
  assign n8933 = ~n8923 & ~n8932;
  assign n8934 = ~n8921 & ~n8933;
  assign n8935 = ~n7428 & ~n8934;
  assign n8936 = ~n8416 & ~n32835;
  assign n8937 = ~n8896 & n8936;
  assign n8938 = n8421 & ~n8937;
  assign n8939 = ~n8421 & n8936;
  assign n8940 = ~n8421 & n8937;
  assign n8941 = ~n8896 & n8939;
  assign n8942 = ~n8938 & ~n32896;
  assign n8943 = n7428 & ~n8921;
  assign n8944 = ~n8933 & n8943;
  assign n8945 = n7428 & n8934;
  assign n8946 = ~n8942 & ~n32897;
  assign n8947 = ~n8935 & ~n8946;
  assign n8948 = ~n6937 & ~n8947;
  assign n8949 = n6937 & ~n8935;
  assign n8950 = ~n8946 & n8949;
  assign n8951 = ~n8436 & ~n32837;
  assign n8952 = ~n8436 & ~n8896;
  assign n8953 = ~n32837 & n8952;
  assign n8954 = ~n8896 & n8951;
  assign n8955 = n8445 & ~n32898;
  assign n8956 = n8449 & n8952;
  assign n8957 = n8445 & ~n32837;
  assign n8958 = ~n8436 & n8957;
  assign n8959 = ~n8896 & n8958;
  assign n8960 = ~n8445 & ~n32898;
  assign n8961 = ~n8959 & ~n8960;
  assign n8962 = ~n8955 & ~n8956;
  assign n8963 = ~n8950 & ~n32899;
  assign n8964 = ~n8948 & ~n8963;
  assign n8965 = ~n6507 & ~n8964;
  assign n8966 = n6507 & ~n8948;
  assign n8967 = ~n8963 & n8966;
  assign n8968 = n6507 & n8964;
  assign n8969 = ~n8451 & ~n8453;
  assign n8970 = ~n8896 & n8969;
  assign n8971 = ~n8461 & ~n8970;
  assign n8972 = ~n8451 & n8461;
  assign n8973 = ~n8453 & n8972;
  assign n8974 = n8461 & n8970;
  assign n8975 = ~n8896 & n8973;
  assign n8976 = n8461 & ~n8970;
  assign n8977 = ~n8461 & n8970;
  assign n8978 = ~n8976 & ~n8977;
  assign n8979 = ~n8971 & ~n32901;
  assign n8980 = ~n32900 & n32902;
  assign n8981 = ~n8965 & ~n8980;
  assign n8982 = ~n6051 & ~n8981;
  assign n8983 = n6051 & ~n8965;
  assign n8984 = ~n8980 & n8983;
  assign n8985 = ~n8464 & ~n32840;
  assign n8986 = ~n8464 & ~n8896;
  assign n8987 = ~n32840 & n8986;
  assign n8988 = ~n8896 & n8985;
  assign n8989 = n8472 & ~n32903;
  assign n8990 = n8476 & n8986;
  assign n8991 = n8472 & ~n32840;
  assign n8992 = ~n8464 & n8991;
  assign n8993 = ~n8896 & n8992;
  assign n8994 = ~n8472 & ~n32903;
  assign n8995 = ~n8993 & ~n8994;
  assign n8996 = ~n8989 & ~n8990;
  assign n8997 = ~n8984 & ~n32904;
  assign n8998 = ~n8982 & ~n8997;
  assign n8999 = ~n5648 & ~n8998;
  assign n9000 = n5648 & ~n8982;
  assign n9001 = ~n8997 & n9000;
  assign n9002 = n5648 & n8998;
  assign n9003 = ~n8478 & ~n8480;
  assign n9004 = ~n8896 & n9003;
  assign n9005 = ~n32842 & ~n9004;
  assign n9006 = n32842 & n9004;
  assign n9007 = ~n8478 & ~n32842;
  assign n9008 = ~n8480 & n9007;
  assign n9009 = ~n8896 & n9008;
  assign n9010 = n32842 & ~n9004;
  assign n9011 = ~n9009 & ~n9010;
  assign n9012 = ~n9005 & ~n9006;
  assign n9013 = ~n32905 & ~n32906;
  assign n9014 = ~n8999 & ~n9013;
  assign n9015 = ~n5223 & ~n9014;
  assign n9016 = n5223 & ~n8999;
  assign n9017 = ~n9013 & n9016;
  assign n9018 = ~n8494 & ~n32844;
  assign n9019 = ~n8494 & ~n8896;
  assign n9020 = ~n32844 & n9019;
  assign n9021 = ~n8896 & n9018;
  assign n9022 = n8502 & ~n32907;
  assign n9023 = n8506 & n9019;
  assign n9024 = n8502 & ~n32844;
  assign n9025 = ~n8494 & n9024;
  assign n9026 = ~n8896 & n9025;
  assign n9027 = ~n8502 & ~n32907;
  assign n9028 = ~n9026 & ~n9027;
  assign n9029 = ~n9022 & ~n9023;
  assign n9030 = ~n9017 & ~n32908;
  assign n9031 = ~n9015 & ~n9030;
  assign n9032 = ~n4851 & ~n9031;
  assign n9033 = n4851 & ~n9015;
  assign n9034 = ~n9030 & n9033;
  assign n9035 = n4851 & n9031;
  assign n9036 = ~n8508 & ~n8510;
  assign n9037 = ~n8896 & n9036;
  assign n9038 = ~n32845 & n9037;
  assign n9039 = n32845 & ~n9037;
  assign n9040 = ~n8508 & n32845;
  assign n9041 = ~n8510 & n9040;
  assign n9042 = ~n8896 & n9041;
  assign n9043 = ~n32845 & ~n9037;
  assign n9044 = ~n9042 & ~n9043;
  assign n9045 = ~n9038 & ~n9039;
  assign n9046 = ~n32909 & ~n32910;
  assign n9047 = ~n9032 & ~n9046;
  assign n9048 = ~n4461 & ~n9047;
  assign n9049 = n4461 & ~n9032;
  assign n9050 = ~n9046 & n9049;
  assign n9051 = ~n8523 & ~n32847;
  assign n9052 = ~n8523 & ~n8896;
  assign n9053 = ~n32847 & n9052;
  assign n9054 = ~n8896 & n9051;
  assign n9055 = n8531 & ~n32911;
  assign n9056 = n8535 & n9052;
  assign n9057 = n8531 & ~n32847;
  assign n9058 = ~n8523 & n9057;
  assign n9059 = ~n8896 & n9058;
  assign n9060 = ~n8531 & ~n32911;
  assign n9061 = ~n9059 & ~n9060;
  assign n9062 = ~n9055 & ~n9056;
  assign n9063 = ~n9050 & ~n32912;
  assign n9064 = ~n9048 & ~n9063;
  assign n9065 = ~n4115 & ~n9064;
  assign n9066 = n4115 & ~n9048;
  assign n9067 = ~n9063 & n9066;
  assign n9068 = n4115 & n9064;
  assign n9069 = ~n8537 & ~n8539;
  assign n9070 = ~n8896 & n9069;
  assign n9071 = ~n32848 & n9070;
  assign n9072 = n32848 & ~n9070;
  assign n9073 = ~n32848 & ~n9070;
  assign n9074 = ~n8537 & n32848;
  assign n9075 = ~n8539 & n9074;
  assign n9076 = n32848 & n9070;
  assign n9077 = ~n8896 & n9075;
  assign n9078 = ~n9073 & ~n32914;
  assign n9079 = ~n9071 & ~n9072;
  assign n9080 = ~n32913 & ~n32915;
  assign n9081 = ~n9065 & ~n9080;
  assign n9082 = ~n3754 & ~n9081;
  assign n9083 = n3754 & ~n9065;
  assign n9084 = ~n9080 & n9083;
  assign n9085 = ~n8552 & ~n32850;
  assign n9086 = ~n8552 & ~n8896;
  assign n9087 = ~n32850 & n9086;
  assign n9088 = ~n8896 & n9085;
  assign n9089 = n8560 & ~n32916;
  assign n9090 = n8564 & n9086;
  assign n9091 = n8560 & ~n32850;
  assign n9092 = ~n8552 & n9091;
  assign n9093 = ~n8896 & n9092;
  assign n9094 = ~n8560 & ~n32916;
  assign n9095 = ~n9093 & ~n9094;
  assign n9096 = ~n9089 & ~n9090;
  assign n9097 = ~n9084 & ~n32917;
  assign n9098 = ~n9082 & ~n9097;
  assign n9099 = ~n3444 & ~n9098;
  assign n9100 = n3444 & ~n9082;
  assign n9101 = ~n9097 & n9100;
  assign n9102 = n3444 & n9098;
  assign n9103 = ~n8566 & ~n8568;
  assign n9104 = ~n8566 & ~n8896;
  assign n9105 = ~n8568 & n9104;
  assign n9106 = ~n8896 & n9103;
  assign n9107 = n32852 & ~n32919;
  assign n9108 = n8580 & n9104;
  assign n9109 = ~n32852 & n32919;
  assign n9110 = ~n8566 & n32852;
  assign n9111 = ~n8568 & n9110;
  assign n9112 = ~n8896 & n9111;
  assign n9113 = ~n32852 & ~n32919;
  assign n9114 = ~n9112 & ~n9113;
  assign n9115 = ~n9107 & ~n32920;
  assign n9116 = ~n32918 & ~n32921;
  assign n9117 = ~n9099 & ~n9116;
  assign n9118 = ~n3116 & ~n9117;
  assign n9119 = n3116 & ~n9099;
  assign n9120 = ~n9116 & n9119;
  assign n9121 = ~n8582 & ~n32854;
  assign n9122 = ~n8582 & ~n8896;
  assign n9123 = ~n32854 & n9122;
  assign n9124 = ~n8896 & n9121;
  assign n9125 = n8590 & ~n32922;
  assign n9126 = n8594 & n9122;
  assign n9127 = n8590 & ~n32854;
  assign n9128 = ~n8582 & n9127;
  assign n9129 = ~n8896 & n9128;
  assign n9130 = ~n8590 & ~n32922;
  assign n9131 = ~n9129 & ~n9130;
  assign n9132 = ~n9125 & ~n9126;
  assign n9133 = ~n9120 & ~n32923;
  assign n9134 = ~n9118 & ~n9133;
  assign n9135 = ~n2833 & ~n9134;
  assign n9136 = ~n8596 & ~n8598;
  assign n9137 = ~n8896 & n9136;
  assign n9138 = ~n32857 & ~n9137;
  assign n9139 = ~n8596 & n32857;
  assign n9140 = ~n8598 & n9139;
  assign n9141 = n32857 & n9137;
  assign n9142 = ~n8896 & n9140;
  assign n9143 = ~n9138 & ~n32924;
  assign n9144 = n2833 & ~n9118;
  assign n9145 = ~n9133 & n9144;
  assign n9146 = n2833 & n9134;
  assign n9147 = ~n9143 & ~n32925;
  assign n9148 = ~n9135 & ~n9147;
  assign n9149 = ~n2536 & ~n9148;
  assign n9150 = n2536 & ~n9135;
  assign n9151 = ~n9147 & n9150;
  assign n9152 = ~n8614 & ~n32859;
  assign n9153 = ~n8614 & ~n8896;
  assign n9154 = ~n32859 & n9153;
  assign n9155 = ~n8896 & n9152;
  assign n9156 = n8622 & ~n32926;
  assign n9157 = n8626 & n9153;
  assign n9158 = n8622 & ~n32859;
  assign n9159 = ~n8614 & n9158;
  assign n9160 = ~n8896 & n9159;
  assign n9161 = ~n8622 & ~n32926;
  assign n9162 = ~n9160 & ~n9161;
  assign n9163 = ~n9156 & ~n9157;
  assign n9164 = ~n9151 & ~n32927;
  assign n9165 = ~n9149 & ~n9164;
  assign n9166 = ~n2283 & ~n9165;
  assign n9167 = n2283 & ~n9149;
  assign n9168 = ~n9164 & n9167;
  assign n9169 = n2283 & n9165;
  assign n9170 = ~n8628 & ~n8638;
  assign n9171 = ~n8628 & ~n8896;
  assign n9172 = ~n8638 & n9171;
  assign n9173 = ~n8896 & n9170;
  assign n9174 = n8636 & ~n32929;
  assign n9175 = n8639 & n9171;
  assign n9176 = ~n8628 & n8636;
  assign n9177 = ~n8638 & n9176;
  assign n9178 = ~n8896 & n9177;
  assign n9179 = ~n8636 & ~n32929;
  assign n9180 = ~n9178 & ~n9179;
  assign n9181 = ~n9174 & ~n9175;
  assign n9182 = ~n32928 & ~n32930;
  assign n9183 = ~n9166 & ~n9182;
  assign n9184 = ~n2021 & ~n9183;
  assign n9185 = n2021 & ~n9166;
  assign n9186 = ~n9182 & n9185;
  assign n9187 = ~n8641 & ~n32862;
  assign n9188 = ~n8641 & ~n8896;
  assign n9189 = ~n32862 & n9188;
  assign n9190 = ~n8896 & n9187;
  assign n9191 = n8649 & ~n32931;
  assign n9192 = n8653 & n9188;
  assign n9193 = n8649 & ~n32862;
  assign n9194 = ~n8641 & n9193;
  assign n9195 = ~n8896 & n9194;
  assign n9196 = ~n8649 & ~n32931;
  assign n9197 = ~n9195 & ~n9196;
  assign n9198 = ~n9191 & ~n9192;
  assign n9199 = ~n9186 & ~n32932;
  assign n9200 = ~n9184 & ~n9199;
  assign n9201 = ~n1796 & ~n9200;
  assign n9202 = ~n8655 & ~n8657;
  assign n9203 = ~n8896 & n9202;
  assign n9204 = ~n32864 & ~n9203;
  assign n9205 = ~n8655 & n32864;
  assign n9206 = ~n8657 & n9205;
  assign n9207 = n32864 & n9203;
  assign n9208 = ~n8896 & n9206;
  assign n9209 = ~n9204 & ~n32933;
  assign n9210 = n1796 & ~n9184;
  assign n9211 = ~n9199 & n9210;
  assign n9212 = n1796 & n9200;
  assign n9213 = ~n9209 & ~n32934;
  assign n9214 = ~n9201 & ~n9213;
  assign n9215 = ~n1567 & ~n9214;
  assign n9216 = n1567 & ~n9201;
  assign n9217 = ~n9213 & n9216;
  assign n9218 = ~n8672 & ~n32866;
  assign n9219 = ~n8672 & ~n8896;
  assign n9220 = ~n32866 & n9219;
  assign n9221 = ~n8896 & n9218;
  assign n9222 = n8680 & ~n32935;
  assign n9223 = n8684 & n9219;
  assign n9224 = n8680 & ~n32866;
  assign n9225 = ~n8672 & n9224;
  assign n9226 = ~n8896 & n9225;
  assign n9227 = ~n8680 & ~n32935;
  assign n9228 = ~n9226 & ~n9227;
  assign n9229 = ~n9222 & ~n9223;
  assign n9230 = ~n9217 & ~n32936;
  assign n9231 = ~n9215 & ~n9230;
  assign n9232 = ~n1374 & ~n9231;
  assign n9233 = n1374 & ~n9215;
  assign n9234 = ~n9230 & n9233;
  assign n9235 = n1374 & n9231;
  assign n9236 = ~n8686 & ~n8696;
  assign n9237 = ~n8686 & ~n8896;
  assign n9238 = ~n8696 & n9237;
  assign n9239 = ~n8896 & n9236;
  assign n9240 = n8694 & ~n32938;
  assign n9241 = n8697 & n9237;
  assign n9242 = ~n8686 & n8694;
  assign n9243 = ~n8696 & n9242;
  assign n9244 = ~n8896 & n9243;
  assign n9245 = ~n8694 & ~n32938;
  assign n9246 = ~n9244 & ~n9245;
  assign n9247 = ~n9240 & ~n9241;
  assign n9248 = ~n32937 & ~n32939;
  assign n9249 = ~n9232 & ~n9248;
  assign n9250 = ~n1179 & ~n9249;
  assign n9251 = n1179 & ~n9232;
  assign n9252 = ~n9248 & n9251;
  assign n9253 = ~n8699 & ~n32869;
  assign n9254 = ~n8699 & ~n8896;
  assign n9255 = ~n32869 & n9254;
  assign n9256 = ~n8896 & n9253;
  assign n9257 = n8707 & ~n32940;
  assign n9258 = n8711 & n9254;
  assign n9259 = n8707 & ~n32869;
  assign n9260 = ~n8699 & n9259;
  assign n9261 = ~n8896 & n9260;
  assign n9262 = ~n8707 & ~n32940;
  assign n9263 = ~n9261 & ~n9262;
  assign n9264 = ~n9257 & ~n9258;
  assign n9265 = ~n9252 & ~n32941;
  assign n9266 = ~n9250 & ~n9265;
  assign n9267 = ~n1016 & ~n9266;
  assign n9268 = ~n8713 & ~n8715;
  assign n9269 = ~n8896 & n9268;
  assign n9270 = ~n32871 & ~n9269;
  assign n9271 = ~n8713 & n32871;
  assign n9272 = ~n8715 & n9271;
  assign n9273 = n32871 & n9269;
  assign n9274 = ~n8896 & n9272;
  assign n9275 = ~n9270 & ~n32942;
  assign n9276 = n1016 & ~n9250;
  assign n9277 = ~n9265 & n9276;
  assign n9278 = n1016 & n9266;
  assign n9279 = ~n9275 & ~n32943;
  assign n9280 = ~n9267 & ~n9279;
  assign n9281 = ~n855 & ~n9280;
  assign n9282 = n855 & ~n9267;
  assign n9283 = ~n9279 & n9282;
  assign n9284 = ~n8730 & ~n32873;
  assign n9285 = ~n8730 & ~n8896;
  assign n9286 = ~n32873 & n9285;
  assign n9287 = ~n8896 & n9284;
  assign n9288 = n8738 & ~n32944;
  assign n9289 = n8742 & n9285;
  assign n9290 = n8738 & ~n32873;
  assign n9291 = ~n8730 & n9290;
  assign n9292 = ~n8896 & n9291;
  assign n9293 = ~n8738 & ~n32944;
  assign n9294 = ~n9292 & ~n9293;
  assign n9295 = ~n9288 & ~n9289;
  assign n9296 = ~n9283 & ~n32945;
  assign n9297 = ~n9281 & ~n9296;
  assign n9298 = ~n720 & ~n9297;
  assign n9299 = n720 & ~n9281;
  assign n9300 = ~n9296 & n9299;
  assign n9301 = n720 & n9297;
  assign n9302 = ~n8744 & ~n8754;
  assign n9303 = ~n8744 & ~n8896;
  assign n9304 = ~n8754 & n9303;
  assign n9305 = ~n8896 & n9302;
  assign n9306 = n8752 & ~n32947;
  assign n9307 = n8755 & n9303;
  assign n9308 = ~n8744 & n8752;
  assign n9309 = ~n8754 & n9308;
  assign n9310 = ~n8896 & n9309;
  assign n9311 = ~n8752 & ~n32947;
  assign n9312 = ~n9310 & ~n9311;
  assign n9313 = ~n9306 & ~n9307;
  assign n9314 = ~n32946 & ~n32948;
  assign n9315 = ~n9298 & ~n9314;
  assign n9316 = ~n592 & ~n9315;
  assign n9317 = n592 & ~n9298;
  assign n9318 = ~n9314 & n9317;
  assign n9319 = ~n8757 & ~n32876;
  assign n9320 = ~n8757 & ~n8896;
  assign n9321 = ~n32876 & n9320;
  assign n9322 = ~n8896 & n9319;
  assign n9323 = n8765 & ~n32949;
  assign n9324 = n8769 & n9320;
  assign n9325 = n8765 & ~n32876;
  assign n9326 = ~n8757 & n9325;
  assign n9327 = ~n8896 & n9326;
  assign n9328 = ~n8765 & ~n32949;
  assign n9329 = ~n9327 & ~n9328;
  assign n9330 = ~n9323 & ~n9324;
  assign n9331 = ~n9318 & ~n32950;
  assign n9332 = ~n9316 & ~n9331;
  assign n9333 = ~n487 & ~n9332;
  assign n9334 = ~n8771 & ~n8773;
  assign n9335 = ~n8896 & n9334;
  assign n9336 = ~n32878 & ~n9335;
  assign n9337 = ~n8771 & n32878;
  assign n9338 = ~n8773 & n9337;
  assign n9339 = n32878 & n9335;
  assign n9340 = ~n8896 & n9338;
  assign n9341 = ~n9336 & ~n32951;
  assign n9342 = n487 & ~n9316;
  assign n9343 = ~n9331 & n9342;
  assign n9344 = n487 & n9332;
  assign n9345 = ~n9341 & ~n32952;
  assign n9346 = ~n9333 & ~n9345;
  assign n9347 = ~n393 & ~n9346;
  assign n9348 = n393 & ~n9333;
  assign n9349 = ~n9345 & n9348;
  assign n9350 = ~n8788 & ~n32880;
  assign n9351 = ~n8788 & ~n8896;
  assign n9352 = ~n32880 & n9351;
  assign n9353 = ~n8896 & n9350;
  assign n9354 = n8796 & ~n32953;
  assign n9355 = n8800 & n9351;
  assign n9356 = n8796 & ~n32880;
  assign n9357 = ~n8788 & n9356;
  assign n9358 = ~n8896 & n9357;
  assign n9359 = ~n8796 & ~n32953;
  assign n9360 = ~n9358 & ~n9359;
  assign n9361 = ~n9354 & ~n9355;
  assign n9362 = ~n9349 & ~n32954;
  assign n9363 = ~n9347 & ~n9362;
  assign n9364 = ~n321 & ~n9363;
  assign n9365 = n321 & ~n9347;
  assign n9366 = ~n9362 & n9365;
  assign n9367 = n321 & n9363;
  assign n9368 = ~n8802 & ~n8812;
  assign n9369 = ~n8802 & ~n8896;
  assign n9370 = ~n8812 & n9369;
  assign n9371 = ~n8896 & n9368;
  assign n9372 = n8810 & ~n32956;
  assign n9373 = n8813 & n9369;
  assign n9374 = ~n8802 & n8810;
  assign n9375 = ~n8812 & n9374;
  assign n9376 = ~n8896 & n9375;
  assign n9377 = ~n8810 & ~n32956;
  assign n9378 = ~n9376 & ~n9377;
  assign n9379 = ~n9372 & ~n9373;
  assign n9380 = ~n32955 & ~n32957;
  assign n9381 = ~n9364 & ~n9380;
  assign n9382 = ~n263 & ~n9381;
  assign n9383 = n263 & ~n9364;
  assign n9384 = ~n9380 & n9383;
  assign n9385 = ~n8815 & ~n32883;
  assign n9386 = ~n8815 & ~n8896;
  assign n9387 = ~n32883 & n9386;
  assign n9388 = ~n8896 & n9385;
  assign n9389 = n8823 & ~n32958;
  assign n9390 = n8827 & n9386;
  assign n9391 = n8823 & ~n32883;
  assign n9392 = ~n8815 & n9391;
  assign n9393 = ~n8896 & n9392;
  assign n9394 = ~n8823 & ~n32958;
  assign n9395 = ~n9393 & ~n9394;
  assign n9396 = ~n9389 & ~n9390;
  assign n9397 = ~n9384 & ~n32959;
  assign n9398 = ~n9382 & ~n9397;
  assign n9399 = ~n214 & ~n9398;
  assign n9400 = ~n8829 & ~n8831;
  assign n9401 = ~n8896 & n9400;
  assign n9402 = ~n32885 & ~n9401;
  assign n9403 = ~n8829 & n32885;
  assign n9404 = ~n8831 & n9403;
  assign n9405 = n32885 & n9401;
  assign n9406 = ~n8896 & n9404;
  assign n9407 = ~n9402 & ~n32960;
  assign n9408 = n214 & ~n9382;
  assign n9409 = ~n9397 & n9408;
  assign n9410 = n214 & n9398;
  assign n9411 = ~n9407 & ~n32961;
  assign n9412 = ~n9399 & ~n9411;
  assign n9413 = ~n197 & ~n9412;
  assign n9414 = n197 & ~n9399;
  assign n9415 = ~n9411 & n9414;
  assign n9416 = ~n8846 & ~n32887;
  assign n9417 = ~n8846 & ~n8896;
  assign n9418 = ~n32887 & n9417;
  assign n9419 = ~n8896 & n9416;
  assign n9420 = n8854 & ~n32962;
  assign n9421 = n8858 & n9417;
  assign n9422 = n8854 & ~n32887;
  assign n9423 = ~n8846 & n9422;
  assign n9424 = ~n8896 & n9423;
  assign n9425 = ~n8854 & ~n32962;
  assign n9426 = ~n9424 & ~n9425;
  assign n9427 = ~n9420 & ~n9421;
  assign n9428 = ~n9415 & ~n32963;
  assign n9429 = ~n9413 & ~n9428;
  assign n9430 = ~n8860 & ~n8870;
  assign n9431 = ~n8860 & ~n8896;
  assign n9432 = ~n8870 & n9431;
  assign n9433 = ~n8896 & n9430;
  assign n9434 = n8868 & ~n32964;
  assign n9435 = n8871 & n9431;
  assign n9436 = ~n8860 & n8868;
  assign n9437 = ~n8870 & n9436;
  assign n9438 = ~n8896 & n9437;
  assign n9439 = ~n8868 & ~n32964;
  assign n9440 = ~n9438 & ~n9439;
  assign n9441 = ~n9434 & ~n9435;
  assign n9442 = ~n8872 & ~n8880;
  assign n9443 = ~n8880 & ~n8896;
  assign n9444 = ~n8872 & n9443;
  assign n9445 = ~n8896 & n9442;
  assign n9446 = ~n32891 & ~n32966;
  assign n9447 = ~n32965 & n9446;
  assign n9448 = ~n9429 & n9447;
  assign n9449 = n193 & ~n9448;
  assign n9450 = ~n9413 & n32965;
  assign n9451 = ~n9428 & n9450;
  assign n9452 = n9429 & n32965;
  assign n9453 = n8872 & ~n9443;
  assign n9454 = ~n193 & ~n9442;
  assign n9455 = ~n9453 & n9454;
  assign n9456 = ~n32967 & ~n9455;
  assign n9457 = ~n9449 & n9456;
  assign n9458 = ~n8921 & ~n8923;
  assign n9459 = ~n9457 & n9458;
  assign n9460 = ~n8932 & ~n9459;
  assign n9461 = ~n8923 & n8932;
  assign n9462 = ~n8921 & n9461;
  assign n9463 = n8932 & n9459;
  assign n9464 = ~n9457 & n9462;
  assign n9465 = ~n9460 & ~n32968;
  assign n9466 = ~pi58  & ~n9457;
  assign n9467 = ~pi59  & n9466;
  assign n9468 = n8898 & ~n9457;
  assign n9469 = ~n8896 & ~n9455;
  assign n9470 = ~n32967 & n9469;
  assign n9471 = ~n9449 & n9470;
  assign n9472 = ~n32969 & ~n9471;
  assign n9473 = pi60  & ~n9472;
  assign n9474 = ~pi60  & ~n9471;
  assign n9475 = ~pi60  & n9472;
  assign n9476 = ~n32969 & n9474;
  assign n9477 = ~n9473 & ~n32970;
  assign n9478 = pi58  & ~n9457;
  assign n9479 = ~pi56  & ~pi57 ;
  assign n9480 = ~pi58  & n9479;
  assign n9481 = ~n32830 & ~n32893;
  assign n9482 = ~n8390 & n9481;
  assign n9483 = ~n8409 & n9482;
  assign n9484 = ~n32832 & n9483;
  assign n9485 = n8395 & n8411;
  assign n9486 = ~n8403 & n9484;
  assign n9487 = ~n9480 & ~n32971;
  assign n9488 = ~n8894 & n9487;
  assign n9489 = ~n32891 & n9488;
  assign n9490 = ~n8888 & n9489;
  assign n9491 = ~n9478 & ~n9480;
  assign n9492 = n8896 & n9491;
  assign n9493 = ~n9478 & n9490;
  assign n9494 = pi59  & ~n9466;
  assign n9495 = ~n32969 & ~n9494;
  assign n9496 = ~n32972 & n9495;
  assign n9497 = ~n8896 & ~n9491;
  assign n9498 = n8411 & ~n9497;
  assign n9499 = ~n9496 & ~n9497;
  assign n9500 = n8411 & n9499;
  assign n9501 = ~n9496 & n9498;
  assign n9502 = ~n9477 & ~n32973;
  assign n9503 = ~n8411 & ~n9499;
  assign n9504 = n7885 & ~n9503;
  assign n9505 = ~n9502 & n9504;
  assign n9506 = ~n8901 & ~n32894;
  assign n9507 = ~n9457 & n9506;
  assign n9508 = n8906 & ~n9507;
  assign n9509 = ~n8906 & n9506;
  assign n9510 = ~n8906 & n9507;
  assign n9511 = ~n9457 & n9509;
  assign n9512 = ~n9508 & ~n32974;
  assign n9513 = ~n9505 & ~n9512;
  assign n9514 = ~n9502 & ~n9503;
  assign n9515 = ~n7885 & ~n9514;
  assign n9516 = n7428 & ~n9515;
  assign n9517 = ~n9513 & ~n9515;
  assign n9518 = n7428 & n9517;
  assign n9519 = ~n9513 & n9516;
  assign n9520 = ~n9465 & ~n32975;
  assign n9521 = ~n7428 & ~n9517;
  assign n9522 = ~n9520 & ~n9521;
  assign n9523 = ~n6937 & ~n9522;
  assign n9524 = ~n8935 & n8942;
  assign n9525 = ~n32897 & n9524;
  assign n9526 = ~n8935 & ~n32897;
  assign n9527 = ~n9457 & n9526;
  assign n9528 = n8942 & n9527;
  assign n9529 = ~n9457 & n9525;
  assign n9530 = ~n8942 & ~n9527;
  assign n9531 = ~n32976 & ~n9530;
  assign n9532 = n6937 & ~n9521;
  assign n9533 = ~n9520 & n9532;
  assign n9534 = ~n9531 & ~n9533;
  assign n9535 = ~n9523 & ~n9534;
  assign n9536 = ~n6507 & ~n9535;
  assign n9537 = ~n8948 & ~n8950;
  assign n9538 = ~n9457 & n9537;
  assign n9539 = ~n32899 & ~n9538;
  assign n9540 = ~n8950 & n32899;
  assign n9541 = ~n8948 & n9540;
  assign n9542 = n32899 & n9538;
  assign n9543 = ~n9457 & n9541;
  assign n9544 = ~n9539 & ~n32977;
  assign n9545 = n6507 & ~n9523;
  assign n9546 = n6507 & n9535;
  assign n9547 = ~n9534 & n9545;
  assign n9548 = ~n9544 & ~n32978;
  assign n9549 = ~n9536 & ~n9548;
  assign n9550 = ~n6051 & ~n9549;
  assign n9551 = n6051 & ~n9536;
  assign n9552 = ~n9548 & n9551;
  assign n9553 = ~n8965 & ~n32900;
  assign n9554 = ~n9457 & n9553;
  assign n9555 = ~n32902 & ~n9554;
  assign n9556 = n32902 & n9554;
  assign n9557 = ~n8965 & ~n32902;
  assign n9558 = ~n32900 & n9557;
  assign n9559 = ~n9457 & n9558;
  assign n9560 = n32902 & ~n9554;
  assign n9561 = ~n9559 & ~n9560;
  assign n9562 = ~n9555 & ~n9556;
  assign n9563 = ~n9552 & ~n32979;
  assign n9564 = ~n9550 & ~n9563;
  assign n9565 = ~n5648 & ~n9564;
  assign n9566 = ~n8982 & ~n8984;
  assign n9567 = ~n9457 & n9566;
  assign n9568 = ~n32904 & ~n9567;
  assign n9569 = ~n8984 & n32904;
  assign n9570 = ~n8982 & n9569;
  assign n9571 = n32904 & n9567;
  assign n9572 = ~n9457 & n9570;
  assign n9573 = ~n9568 & ~n32980;
  assign n9574 = n5648 & ~n9550;
  assign n9575 = n5648 & n9564;
  assign n9576 = ~n9563 & n9574;
  assign n9577 = ~n9573 & ~n32981;
  assign n9578 = ~n9565 & ~n9577;
  assign n9579 = ~n5223 & ~n9578;
  assign n9580 = n5223 & ~n9565;
  assign n9581 = ~n9577 & n9580;
  assign n9582 = ~n8999 & ~n32905;
  assign n9583 = ~n9457 & n9582;
  assign n9584 = ~n32906 & n9583;
  assign n9585 = n32906 & ~n9583;
  assign n9586 = ~n8999 & n32906;
  assign n9587 = ~n32905 & n9586;
  assign n9588 = ~n9457 & n9587;
  assign n9589 = ~n32906 & ~n9583;
  assign n9590 = ~n9588 & ~n9589;
  assign n9591 = ~n9584 & ~n9585;
  assign n9592 = ~n9581 & ~n32982;
  assign n9593 = ~n9579 & ~n9592;
  assign n9594 = ~n4851 & ~n9593;
  assign n9595 = ~n9015 & ~n9017;
  assign n9596 = ~n9457 & n9595;
  assign n9597 = ~n32908 & ~n9596;
  assign n9598 = ~n9017 & n32908;
  assign n9599 = ~n9015 & n9598;
  assign n9600 = n32908 & n9596;
  assign n9601 = ~n9457 & n9599;
  assign n9602 = ~n9597 & ~n32983;
  assign n9603 = n4851 & ~n9579;
  assign n9604 = n4851 & n9593;
  assign n9605 = ~n9592 & n9603;
  assign n9606 = ~n9602 & ~n32984;
  assign n9607 = ~n9594 & ~n9606;
  assign n9608 = ~n4461 & ~n9607;
  assign n9609 = n4461 & ~n9594;
  assign n9610 = ~n9606 & n9609;
  assign n9611 = ~n9032 & ~n32909;
  assign n9612 = ~n9457 & n9611;
  assign n9613 = ~n32910 & n9612;
  assign n9614 = n32910 & ~n9612;
  assign n9615 = ~n32910 & ~n9612;
  assign n9616 = ~n9032 & n32910;
  assign n9617 = ~n32909 & n9616;
  assign n9618 = n32910 & n9612;
  assign n9619 = ~n9457 & n9617;
  assign n9620 = ~n9615 & ~n32985;
  assign n9621 = ~n9613 & ~n9614;
  assign n9622 = ~n9610 & ~n32986;
  assign n9623 = ~n9608 & ~n9622;
  assign n9624 = ~n4115 & ~n9623;
  assign n9625 = ~n9048 & ~n9050;
  assign n9626 = ~n9457 & n9625;
  assign n9627 = ~n32912 & ~n9626;
  assign n9628 = ~n9050 & n32912;
  assign n9629 = ~n9048 & n9628;
  assign n9630 = n32912 & n9626;
  assign n9631 = ~n9457 & n9629;
  assign n9632 = ~n9627 & ~n32987;
  assign n9633 = n4115 & ~n9608;
  assign n9634 = n4115 & n9623;
  assign n9635 = ~n9622 & n9633;
  assign n9636 = ~n9632 & ~n32988;
  assign n9637 = ~n9624 & ~n9636;
  assign n9638 = ~n3754 & ~n9637;
  assign n9639 = n3754 & ~n9624;
  assign n9640 = ~n9636 & n9639;
  assign n9641 = ~n9065 & ~n32913;
  assign n9642 = ~n9065 & ~n9457;
  assign n9643 = ~n32913 & n9642;
  assign n9644 = ~n9457 & n9641;
  assign n9645 = n32915 & ~n32989;
  assign n9646 = n9080 & n9642;
  assign n9647 = ~n32915 & n32989;
  assign n9648 = ~n9065 & n32915;
  assign n9649 = ~n32913 & n9648;
  assign n9650 = ~n9457 & n9649;
  assign n9651 = ~n32915 & ~n32989;
  assign n9652 = ~n9650 & ~n9651;
  assign n9653 = ~n9645 & ~n32990;
  assign n9654 = ~n9640 & ~n32991;
  assign n9655 = ~n9638 & ~n9654;
  assign n9656 = ~n3444 & ~n9655;
  assign n9657 = ~n9082 & ~n9084;
  assign n9658 = ~n9457 & n9657;
  assign n9659 = ~n32917 & ~n9658;
  assign n9660 = ~n9084 & n32917;
  assign n9661 = ~n9082 & n9660;
  assign n9662 = n32917 & n9658;
  assign n9663 = ~n9457 & n9661;
  assign n9664 = ~n9659 & ~n32992;
  assign n9665 = n3444 & ~n9638;
  assign n9666 = n3444 & n9655;
  assign n9667 = ~n9654 & n9665;
  assign n9668 = ~n9664 & ~n32993;
  assign n9669 = ~n9656 & ~n9668;
  assign n9670 = ~n3116 & ~n9669;
  assign n9671 = ~n9099 & ~n32918;
  assign n9672 = ~n9457 & n9671;
  assign n9673 = ~n32921 & ~n9672;
  assign n9674 = ~n9099 & n32921;
  assign n9675 = ~n32918 & n9674;
  assign n9676 = n32921 & n9672;
  assign n9677 = ~n9457 & n9675;
  assign n9678 = ~n9673 & ~n32994;
  assign n9679 = n3116 & ~n9656;
  assign n9680 = ~n9668 & n9679;
  assign n9681 = ~n9678 & ~n9680;
  assign n9682 = ~n9670 & ~n9681;
  assign n9683 = ~n2833 & ~n9682;
  assign n9684 = ~n9118 & ~n9120;
  assign n9685 = ~n9457 & n9684;
  assign n9686 = ~n32923 & ~n9685;
  assign n9687 = ~n9120 & n32923;
  assign n9688 = ~n9118 & n9687;
  assign n9689 = n32923 & n9685;
  assign n9690 = ~n9457 & n9688;
  assign n9691 = ~n9686 & ~n32995;
  assign n9692 = n2833 & ~n9670;
  assign n9693 = n2833 & n9682;
  assign n9694 = ~n9681 & n9692;
  assign n9695 = ~n9691 & ~n32996;
  assign n9696 = ~n9683 & ~n9695;
  assign n9697 = ~n2536 & ~n9696;
  assign n9698 = n2536 & ~n9683;
  assign n9699 = ~n9695 & n9698;
  assign n9700 = ~n9135 & ~n32925;
  assign n9701 = ~n9135 & ~n9457;
  assign n9702 = ~n32925 & n9701;
  assign n9703 = ~n9457 & n9700;
  assign n9704 = n9143 & ~n32997;
  assign n9705 = n9147 & n9701;
  assign n9706 = ~n9135 & n9143;
  assign n9707 = ~n32925 & n9706;
  assign n9708 = ~n9457 & n9707;
  assign n9709 = ~n9143 & ~n32997;
  assign n9710 = ~n9708 & ~n9709;
  assign n9711 = ~n9704 & ~n9705;
  assign n9712 = ~n9699 & ~n32998;
  assign n9713 = ~n9697 & ~n9712;
  assign n9714 = ~n2283 & ~n9713;
  assign n9715 = ~n9149 & ~n9151;
  assign n9716 = ~n9457 & n9715;
  assign n9717 = ~n32927 & ~n9716;
  assign n9718 = ~n9151 & n32927;
  assign n9719 = ~n9149 & n9718;
  assign n9720 = n32927 & n9716;
  assign n9721 = ~n9457 & n9719;
  assign n9722 = ~n9717 & ~n32999;
  assign n9723 = n2283 & ~n9697;
  assign n9724 = n2283 & n9713;
  assign n9725 = ~n9712 & n9723;
  assign n9726 = ~n9722 & ~n33000;
  assign n9727 = ~n9714 & ~n9726;
  assign n9728 = ~n2021 & ~n9727;
  assign n9729 = ~n9166 & ~n32928;
  assign n9730 = ~n9457 & n9729;
  assign n9731 = ~n32930 & ~n9730;
  assign n9732 = ~n9166 & n32930;
  assign n9733 = ~n32928 & n9732;
  assign n9734 = n32930 & n9730;
  assign n9735 = ~n9457 & n9733;
  assign n9736 = ~n9731 & ~n33001;
  assign n9737 = n2021 & ~n9714;
  assign n9738 = ~n9726 & n9737;
  assign n9739 = ~n9736 & ~n9738;
  assign n9740 = ~n9728 & ~n9739;
  assign n9741 = ~n1796 & ~n9740;
  assign n9742 = ~n9184 & ~n9186;
  assign n9743 = ~n9457 & n9742;
  assign n9744 = ~n32932 & ~n9743;
  assign n9745 = ~n9186 & n32932;
  assign n9746 = ~n9184 & n9745;
  assign n9747 = n32932 & n9743;
  assign n9748 = ~n9457 & n9746;
  assign n9749 = ~n9744 & ~n33002;
  assign n9750 = n1796 & ~n9728;
  assign n9751 = n1796 & n9740;
  assign n9752 = ~n9739 & n9750;
  assign n9753 = ~n9749 & ~n33003;
  assign n9754 = ~n9741 & ~n9753;
  assign n9755 = ~n1567 & ~n9754;
  assign n9756 = n1567 & ~n9741;
  assign n9757 = ~n9753 & n9756;
  assign n9758 = ~n9201 & ~n32934;
  assign n9759 = ~n9201 & ~n9457;
  assign n9760 = ~n32934 & n9759;
  assign n9761 = ~n9457 & n9758;
  assign n9762 = n9209 & ~n33004;
  assign n9763 = n9213 & n9759;
  assign n9764 = ~n9201 & n9209;
  assign n9765 = ~n32934 & n9764;
  assign n9766 = ~n9457 & n9765;
  assign n9767 = ~n9209 & ~n33004;
  assign n9768 = ~n9766 & ~n9767;
  assign n9769 = ~n9762 & ~n9763;
  assign n9770 = ~n9757 & ~n33005;
  assign n9771 = ~n9755 & ~n9770;
  assign n9772 = ~n1374 & ~n9771;
  assign n9773 = ~n9215 & ~n9217;
  assign n9774 = ~n9457 & n9773;
  assign n9775 = ~n32936 & ~n9774;
  assign n9776 = ~n9217 & n32936;
  assign n9777 = ~n9215 & n9776;
  assign n9778 = n32936 & n9774;
  assign n9779 = ~n9457 & n9777;
  assign n9780 = ~n9775 & ~n33006;
  assign n9781 = n1374 & ~n9755;
  assign n9782 = n1374 & n9771;
  assign n9783 = ~n9770 & n9781;
  assign n9784 = ~n9780 & ~n33007;
  assign n9785 = ~n9772 & ~n9784;
  assign n9786 = ~n1179 & ~n9785;
  assign n9787 = ~n9232 & ~n32937;
  assign n9788 = ~n9457 & n9787;
  assign n9789 = ~n32939 & ~n9788;
  assign n9790 = ~n9232 & n32939;
  assign n9791 = ~n32937 & n9790;
  assign n9792 = n32939 & n9788;
  assign n9793 = ~n9457 & n9791;
  assign n9794 = ~n9789 & ~n33008;
  assign n9795 = n1179 & ~n9772;
  assign n9796 = ~n9784 & n9795;
  assign n9797 = ~n9794 & ~n9796;
  assign n9798 = ~n9786 & ~n9797;
  assign n9799 = ~n1016 & ~n9798;
  assign n9800 = ~n9250 & ~n9252;
  assign n9801 = ~n9457 & n9800;
  assign n9802 = ~n32941 & ~n9801;
  assign n9803 = ~n9252 & n32941;
  assign n9804 = ~n9250 & n9803;
  assign n9805 = n32941 & n9801;
  assign n9806 = ~n9457 & n9804;
  assign n9807 = ~n9802 & ~n33009;
  assign n9808 = n1016 & ~n9786;
  assign n9809 = n1016 & n9798;
  assign n9810 = ~n9797 & n9808;
  assign n9811 = ~n9807 & ~n33010;
  assign n9812 = ~n9799 & ~n9811;
  assign n9813 = ~n855 & ~n9812;
  assign n9814 = n855 & ~n9799;
  assign n9815 = ~n9811 & n9814;
  assign n9816 = ~n9267 & ~n32943;
  assign n9817 = ~n9267 & ~n9457;
  assign n9818 = ~n32943 & n9817;
  assign n9819 = ~n9457 & n9816;
  assign n9820 = n9275 & ~n33011;
  assign n9821 = n9279 & n9817;
  assign n9822 = ~n9267 & n9275;
  assign n9823 = ~n32943 & n9822;
  assign n9824 = ~n9457 & n9823;
  assign n9825 = ~n9275 & ~n33011;
  assign n9826 = ~n9824 & ~n9825;
  assign n9827 = ~n9820 & ~n9821;
  assign n9828 = ~n9815 & ~n33012;
  assign n9829 = ~n9813 & ~n9828;
  assign n9830 = ~n720 & ~n9829;
  assign n9831 = ~n9281 & ~n9283;
  assign n9832 = ~n9457 & n9831;
  assign n9833 = ~n32945 & ~n9832;
  assign n9834 = ~n9283 & n32945;
  assign n9835 = ~n9281 & n9834;
  assign n9836 = n32945 & n9832;
  assign n9837 = ~n9457 & n9835;
  assign n9838 = ~n9833 & ~n33013;
  assign n9839 = n720 & ~n9813;
  assign n9840 = n720 & n9829;
  assign n9841 = ~n9828 & n9839;
  assign n9842 = ~n9838 & ~n33014;
  assign n9843 = ~n9830 & ~n9842;
  assign n9844 = ~n592 & ~n9843;
  assign n9845 = ~n9298 & ~n32946;
  assign n9846 = ~n9457 & n9845;
  assign n9847 = ~n32948 & ~n9846;
  assign n9848 = ~n9298 & n32948;
  assign n9849 = ~n32946 & n9848;
  assign n9850 = n32948 & n9846;
  assign n9851 = ~n9457 & n9849;
  assign n9852 = ~n9847 & ~n33015;
  assign n9853 = n592 & ~n9830;
  assign n9854 = ~n9842 & n9853;
  assign n9855 = ~n9852 & ~n9854;
  assign n9856 = ~n9844 & ~n9855;
  assign n9857 = ~n487 & ~n9856;
  assign n9858 = ~n9316 & ~n9318;
  assign n9859 = ~n9457 & n9858;
  assign n9860 = ~n32950 & ~n9859;
  assign n9861 = ~n9318 & n32950;
  assign n9862 = ~n9316 & n9861;
  assign n9863 = n32950 & n9859;
  assign n9864 = ~n9457 & n9862;
  assign n9865 = ~n9860 & ~n33016;
  assign n9866 = n487 & ~n9844;
  assign n9867 = n487 & n9856;
  assign n9868 = ~n9855 & n9866;
  assign n9869 = ~n9865 & ~n33017;
  assign n9870 = ~n9857 & ~n9869;
  assign n9871 = ~n393 & ~n9870;
  assign n9872 = n393 & ~n9857;
  assign n9873 = ~n9869 & n9872;
  assign n9874 = ~n9333 & ~n32952;
  assign n9875 = ~n9333 & ~n9457;
  assign n9876 = ~n32952 & n9875;
  assign n9877 = ~n9457 & n9874;
  assign n9878 = n9341 & ~n33018;
  assign n9879 = n9345 & n9875;
  assign n9880 = ~n9333 & n9341;
  assign n9881 = ~n32952 & n9880;
  assign n9882 = ~n9457 & n9881;
  assign n9883 = ~n9341 & ~n33018;
  assign n9884 = ~n9882 & ~n9883;
  assign n9885 = ~n9878 & ~n9879;
  assign n9886 = ~n9873 & ~n33019;
  assign n9887 = ~n9871 & ~n9886;
  assign n9888 = ~n321 & ~n9887;
  assign n9889 = ~n9347 & ~n9349;
  assign n9890 = ~n9457 & n9889;
  assign n9891 = ~n32954 & ~n9890;
  assign n9892 = ~n9349 & n32954;
  assign n9893 = ~n9347 & n9892;
  assign n9894 = n32954 & n9890;
  assign n9895 = ~n9457 & n9893;
  assign n9896 = ~n9891 & ~n33020;
  assign n9897 = n321 & ~n9871;
  assign n9898 = n321 & n9887;
  assign n9899 = ~n9886 & n9897;
  assign n9900 = ~n9896 & ~n33021;
  assign n9901 = ~n9888 & ~n9900;
  assign n9902 = ~n263 & ~n9901;
  assign n9903 = ~n9364 & ~n32955;
  assign n9904 = ~n9457 & n9903;
  assign n9905 = ~n32957 & ~n9904;
  assign n9906 = ~n9364 & n32957;
  assign n9907 = ~n32955 & n9906;
  assign n9908 = n32957 & n9904;
  assign n9909 = ~n9457 & n9907;
  assign n9910 = ~n9905 & ~n33022;
  assign n9911 = n263 & ~n9888;
  assign n9912 = ~n9900 & n9911;
  assign n9913 = ~n9910 & ~n9912;
  assign n9914 = ~n9902 & ~n9913;
  assign n9915 = ~n214 & ~n9914;
  assign n9916 = ~n9382 & ~n9384;
  assign n9917 = ~n9457 & n9916;
  assign n9918 = ~n32959 & ~n9917;
  assign n9919 = ~n9384 & n32959;
  assign n9920 = ~n9382 & n9919;
  assign n9921 = n32959 & n9917;
  assign n9922 = ~n9457 & n9920;
  assign n9923 = ~n9918 & ~n33023;
  assign n9924 = n214 & ~n9902;
  assign n9925 = n214 & n9914;
  assign n9926 = ~n9913 & n9924;
  assign n9927 = ~n9923 & ~n33024;
  assign n9928 = ~n9915 & ~n9927;
  assign n9929 = ~n197 & ~n9928;
  assign n9930 = n197 & ~n9915;
  assign n9931 = ~n9927 & n9930;
  assign n9932 = ~n9399 & ~n32961;
  assign n9933 = ~n9399 & ~n9457;
  assign n9934 = ~n32961 & n9933;
  assign n9935 = ~n9457 & n9932;
  assign n9936 = n9407 & ~n33025;
  assign n9937 = n9411 & n9933;
  assign n9938 = ~n9399 & n9407;
  assign n9939 = ~n32961 & n9938;
  assign n9940 = ~n9457 & n9939;
  assign n9941 = ~n9407 & ~n33025;
  assign n9942 = ~n9940 & ~n9941;
  assign n9943 = ~n9936 & ~n9937;
  assign n9944 = ~n9931 & ~n33026;
  assign n9945 = ~n9929 & ~n9944;
  assign n9946 = ~n9413 & ~n9415;
  assign n9947 = ~n9457 & n9946;
  assign n9948 = ~n32963 & ~n9947;
  assign n9949 = ~n9415 & n32963;
  assign n9950 = ~n9413 & n9949;
  assign n9951 = n32963 & n9947;
  assign n9952 = ~n9457 & n9950;
  assign n9953 = ~n9948 & ~n33027;
  assign n9954 = ~n9429 & ~n32965;
  assign n9955 = ~n32965 & ~n9457;
  assign n9956 = ~n9429 & n9955;
  assign n9957 = ~n9457 & n9954;
  assign n9958 = ~n32967 & ~n33028;
  assign n9959 = ~n9953 & n9958;
  assign n9960 = ~n9945 & n9959;
  assign n9961 = n193 & ~n9960;
  assign n9962 = ~n9929 & n9953;
  assign n9963 = n9945 & n9953;
  assign n9964 = ~n9944 & n9962;
  assign n9965 = n9429 & ~n9955;
  assign n9966 = ~n193 & ~n9954;
  assign n9967 = ~n9965 & n9966;
  assign n9968 = ~n33029 & ~n9967;
  assign n9969 = ~n9961 & n9968;
  assign n9970 = pi56  & ~n9969;
  assign n9971 = ~pi54  & ~pi55 ;
  assign n9972 = ~pi56  & n9971;
  assign n9973 = ~n9970 & ~n9972;
  assign n9974 = ~n9457 & ~n9973;
  assign n9975 = ~pi56  & ~n9969;
  assign n9976 = pi57  & ~n9975;
  assign n9977 = ~pi57  & n9975;
  assign n9978 = n9479 & ~n9969;
  assign n9979 = ~n9976 & ~n33030;
  assign n9980 = ~n32889 & ~n32971;
  assign n9981 = ~n8875 & n9980;
  assign n9982 = ~n8894 & n9981;
  assign n9983 = ~n32891 & n9982;
  assign n9984 = n8880 & n8896;
  assign n9985 = ~n8888 & n9983;
  assign n9986 = ~n9972 & ~n33031;
  assign n9987 = ~n9455 & n9986;
  assign n9988 = ~n32967 & n9987;
  assign n9989 = ~n9449 & n9988;
  assign n9990 = n9457 & n9973;
  assign n9991 = ~n9970 & n9989;
  assign n9992 = n9979 & ~n33032;
  assign n9993 = ~n9974 & ~n9992;
  assign n9994 = ~n8896 & ~n9993;
  assign n9995 = n8896 & ~n9974;
  assign n9996 = ~n9992 & n9995;
  assign n9997 = ~n9457 & ~n9967;
  assign n9998 = ~n33029 & n9997;
  assign n9999 = ~n9961 & n9998;
  assign n10000 = ~n33030 & ~n9999;
  assign n10001 = pi58  & ~n10000;
  assign n10002 = ~pi58  & ~n9999;
  assign n10003 = ~pi58  & n10000;
  assign n10004 = ~n33030 & n10002;
  assign n10005 = ~n10001 & ~n33033;
  assign n10006 = ~n9996 & ~n10005;
  assign n10007 = ~n9994 & ~n10006;
  assign n10008 = ~n8411 & ~n10007;
  assign n10009 = n8411 & ~n9994;
  assign n10010 = ~n10006 & n10009;
  assign n10011 = n8411 & n10007;
  assign n10012 = ~n32972 & ~n9497;
  assign n10013 = ~n9969 & n10012;
  assign n10014 = n9495 & ~n10013;
  assign n10015 = ~n9495 & n10012;
  assign n10016 = ~n9495 & n10013;
  assign n10017 = ~n9969 & n10015;
  assign n10018 = ~n10014 & ~n33035;
  assign n10019 = ~n33034 & ~n10018;
  assign n10020 = ~n10008 & ~n10019;
  assign n10021 = ~n7885 & ~n10020;
  assign n10022 = n7885 & ~n10008;
  assign n10023 = ~n10019 & n10022;
  assign n10024 = ~n32973 & ~n9503;
  assign n10025 = ~n9503 & ~n9969;
  assign n10026 = ~n32973 & n10025;
  assign n10027 = ~n9969 & n10024;
  assign n10028 = n9477 & ~n33036;
  assign n10029 = n9502 & n10025;
  assign n10030 = n9477 & ~n32973;
  assign n10031 = ~n9503 & n10030;
  assign n10032 = ~n9969 & n10031;
  assign n10033 = ~n9477 & ~n33036;
  assign n10034 = ~n10032 & ~n10033;
  assign n10035 = ~n10028 & ~n10029;
  assign n10036 = ~n10023 & ~n33037;
  assign n10037 = ~n10021 & ~n10036;
  assign n10038 = ~n7428 & ~n10037;
  assign n10039 = n7428 & ~n10021;
  assign n10040 = ~n10036 & n10039;
  assign n10041 = n7428 & n10037;
  assign n10042 = ~n9505 & ~n9515;
  assign n10043 = ~n9969 & n10042;
  assign n10044 = ~n9512 & ~n10043;
  assign n10045 = n9512 & ~n9515;
  assign n10046 = ~n9505 & n10045;
  assign n10047 = n9512 & n10043;
  assign n10048 = ~n9969 & n10046;
  assign n10049 = n9512 & ~n10043;
  assign n10050 = ~n9512 & n10043;
  assign n10051 = ~n10049 & ~n10050;
  assign n10052 = ~n10044 & ~n33039;
  assign n10053 = ~n33038 & n33040;
  assign n10054 = ~n10038 & ~n10053;
  assign n10055 = ~n6937 & ~n10054;
  assign n10056 = n6937 & ~n10038;
  assign n10057 = ~n10053 & n10056;
  assign n10058 = n9465 & ~n32975;
  assign n10059 = ~n9521 & n10058;
  assign n10060 = ~n32975 & ~n9521;
  assign n10061 = ~n9969 & n10060;
  assign n10062 = n9465 & n10061;
  assign n10063 = ~n9969 & n10059;
  assign n10064 = ~n9465 & ~n10061;
  assign n10065 = ~n33041 & ~n10064;
  assign n10066 = ~n10057 & ~n10065;
  assign n10067 = ~n10055 & ~n10066;
  assign n10068 = ~n6507 & ~n10067;
  assign n10069 = ~n9523 & ~n9533;
  assign n10070 = ~n9969 & n10069;
  assign n10071 = ~n9531 & ~n10070;
  assign n10072 = ~n9523 & n9531;
  assign n10073 = ~n9533 & n10072;
  assign n10074 = n9531 & n10070;
  assign n10075 = ~n9969 & n10073;
  assign n10076 = ~n10071 & ~n33042;
  assign n10077 = n6507 & ~n10055;
  assign n10078 = ~n10066 & n10077;
  assign n10079 = n6507 & n10067;
  assign n10080 = ~n10076 & ~n33043;
  assign n10081 = ~n10068 & ~n10080;
  assign n10082 = ~n6051 & ~n10081;
  assign n10083 = n6051 & ~n10068;
  assign n10084 = ~n10080 & n10083;
  assign n10085 = ~n9536 & ~n32978;
  assign n10086 = ~n9536 & ~n9969;
  assign n10087 = ~n32978 & n10086;
  assign n10088 = ~n9969 & n10085;
  assign n10089 = n9544 & ~n33044;
  assign n10090 = n9548 & n10086;
  assign n10091 = n9544 & ~n32978;
  assign n10092 = ~n9536 & n10091;
  assign n10093 = ~n9969 & n10092;
  assign n10094 = ~n9544 & ~n33044;
  assign n10095 = ~n10093 & ~n10094;
  assign n10096 = ~n10089 & ~n10090;
  assign n10097 = ~n10084 & ~n33045;
  assign n10098 = ~n10082 & ~n10097;
  assign n10099 = ~n5648 & ~n10098;
  assign n10100 = n5648 & ~n10082;
  assign n10101 = ~n10097 & n10100;
  assign n10102 = n5648 & n10098;
  assign n10103 = ~n9550 & ~n9552;
  assign n10104 = ~n9969 & n10103;
  assign n10105 = ~n32979 & n10104;
  assign n10106 = n32979 & ~n10104;
  assign n10107 = ~n9550 & n32979;
  assign n10108 = ~n9552 & n10107;
  assign n10109 = ~n9969 & n10108;
  assign n10110 = ~n32979 & ~n10104;
  assign n10111 = ~n10109 & ~n10110;
  assign n10112 = ~n10105 & ~n10106;
  assign n10113 = ~n33046 & ~n33047;
  assign n10114 = ~n10099 & ~n10113;
  assign n10115 = ~n5223 & ~n10114;
  assign n10116 = n5223 & ~n10099;
  assign n10117 = ~n10113 & n10116;
  assign n10118 = ~n9565 & ~n32981;
  assign n10119 = ~n9565 & ~n9969;
  assign n10120 = ~n32981 & n10119;
  assign n10121 = ~n9969 & n10118;
  assign n10122 = n9573 & ~n33048;
  assign n10123 = n9577 & n10119;
  assign n10124 = n9573 & ~n32981;
  assign n10125 = ~n9565 & n10124;
  assign n10126 = ~n9969 & n10125;
  assign n10127 = ~n9573 & ~n33048;
  assign n10128 = ~n10126 & ~n10127;
  assign n10129 = ~n10122 & ~n10123;
  assign n10130 = ~n10117 & ~n33049;
  assign n10131 = ~n10115 & ~n10130;
  assign n10132 = ~n4851 & ~n10131;
  assign n10133 = n4851 & ~n10115;
  assign n10134 = ~n10130 & n10133;
  assign n10135 = n4851 & n10131;
  assign n10136 = ~n9579 & ~n9581;
  assign n10137 = ~n9969 & n10136;
  assign n10138 = ~n32982 & n10137;
  assign n10139 = n32982 & ~n10137;
  assign n10140 = ~n32982 & ~n10137;
  assign n10141 = ~n9579 & n32982;
  assign n10142 = ~n9581 & n10141;
  assign n10143 = n32982 & n10137;
  assign n10144 = ~n9969 & n10142;
  assign n10145 = ~n10140 & ~n33051;
  assign n10146 = ~n10138 & ~n10139;
  assign n10147 = ~n33050 & ~n33052;
  assign n10148 = ~n10132 & ~n10147;
  assign n10149 = ~n4461 & ~n10148;
  assign n10150 = n4461 & ~n10132;
  assign n10151 = ~n10147 & n10150;
  assign n10152 = ~n9594 & ~n32984;
  assign n10153 = ~n9594 & ~n9969;
  assign n10154 = ~n32984 & n10153;
  assign n10155 = ~n9969 & n10152;
  assign n10156 = n9602 & ~n33053;
  assign n10157 = n9606 & n10153;
  assign n10158 = n9602 & ~n32984;
  assign n10159 = ~n9594 & n10158;
  assign n10160 = ~n9969 & n10159;
  assign n10161 = ~n9602 & ~n33053;
  assign n10162 = ~n10160 & ~n10161;
  assign n10163 = ~n10156 & ~n10157;
  assign n10164 = ~n10151 & ~n33054;
  assign n10165 = ~n10149 & ~n10164;
  assign n10166 = ~n4115 & ~n10165;
  assign n10167 = n4115 & ~n10149;
  assign n10168 = ~n10164 & n10167;
  assign n10169 = n4115 & n10165;
  assign n10170 = ~n9608 & ~n9610;
  assign n10171 = ~n9608 & ~n9969;
  assign n10172 = ~n9610 & n10171;
  assign n10173 = ~n9969 & n10170;
  assign n10174 = n32986 & ~n33056;
  assign n10175 = n9622 & n10171;
  assign n10176 = ~n32986 & n33056;
  assign n10177 = ~n9608 & n32986;
  assign n10178 = ~n9610 & n10177;
  assign n10179 = ~n9969 & n10178;
  assign n10180 = ~n32986 & ~n33056;
  assign n10181 = ~n10179 & ~n10180;
  assign n10182 = ~n10174 & ~n33057;
  assign n10183 = ~n33055 & ~n33058;
  assign n10184 = ~n10166 & ~n10183;
  assign n10185 = ~n3754 & ~n10184;
  assign n10186 = n3754 & ~n10166;
  assign n10187 = ~n10183 & n10186;
  assign n10188 = ~n9624 & ~n32988;
  assign n10189 = ~n9624 & ~n9969;
  assign n10190 = ~n32988 & n10189;
  assign n10191 = ~n9969 & n10188;
  assign n10192 = n9632 & ~n33059;
  assign n10193 = n9636 & n10189;
  assign n10194 = n9632 & ~n32988;
  assign n10195 = ~n9624 & n10194;
  assign n10196 = ~n9969 & n10195;
  assign n10197 = ~n9632 & ~n33059;
  assign n10198 = ~n10196 & ~n10197;
  assign n10199 = ~n10192 & ~n10193;
  assign n10200 = ~n10187 & ~n33060;
  assign n10201 = ~n10185 & ~n10200;
  assign n10202 = ~n3444 & ~n10201;
  assign n10203 = ~n9638 & ~n9640;
  assign n10204 = ~n9969 & n10203;
  assign n10205 = ~n32991 & ~n10204;
  assign n10206 = ~n9638 & n32991;
  assign n10207 = ~n9640 & n10206;
  assign n10208 = n32991 & n10204;
  assign n10209 = ~n9969 & n10207;
  assign n10210 = ~n10205 & ~n33061;
  assign n10211 = n3444 & ~n10185;
  assign n10212 = ~n10200 & n10211;
  assign n10213 = n3444 & n10201;
  assign n10214 = ~n10210 & ~n33062;
  assign n10215 = ~n10202 & ~n10214;
  assign n10216 = ~n3116 & ~n10215;
  assign n10217 = n3116 & ~n10202;
  assign n10218 = ~n10214 & n10217;
  assign n10219 = ~n9656 & ~n32993;
  assign n10220 = ~n9656 & ~n9969;
  assign n10221 = ~n32993 & n10220;
  assign n10222 = ~n9969 & n10219;
  assign n10223 = n9664 & ~n33063;
  assign n10224 = n9668 & n10220;
  assign n10225 = n9664 & ~n32993;
  assign n10226 = ~n9656 & n10225;
  assign n10227 = ~n9969 & n10226;
  assign n10228 = ~n9664 & ~n33063;
  assign n10229 = ~n10227 & ~n10228;
  assign n10230 = ~n10223 & ~n10224;
  assign n10231 = ~n10218 & ~n33064;
  assign n10232 = ~n10216 & ~n10231;
  assign n10233 = ~n2833 & ~n10232;
  assign n10234 = n2833 & ~n10216;
  assign n10235 = ~n10231 & n10234;
  assign n10236 = n2833 & n10232;
  assign n10237 = ~n9670 & ~n9680;
  assign n10238 = ~n9670 & ~n9969;
  assign n10239 = ~n9680 & n10238;
  assign n10240 = ~n9969 & n10237;
  assign n10241 = n9678 & ~n33066;
  assign n10242 = n9681 & n10238;
  assign n10243 = ~n9670 & n9678;
  assign n10244 = ~n9680 & n10243;
  assign n10245 = ~n9969 & n10244;
  assign n10246 = ~n9678 & ~n33066;
  assign n10247 = ~n10245 & ~n10246;
  assign n10248 = ~n10241 & ~n10242;
  assign n10249 = ~n33065 & ~n33067;
  assign n10250 = ~n10233 & ~n10249;
  assign n10251 = ~n2536 & ~n10250;
  assign n10252 = n2536 & ~n10233;
  assign n10253 = ~n10249 & n10252;
  assign n10254 = ~n9683 & ~n32996;
  assign n10255 = ~n9683 & ~n9969;
  assign n10256 = ~n32996 & n10255;
  assign n10257 = ~n9969 & n10254;
  assign n10258 = n9691 & ~n33068;
  assign n10259 = n9695 & n10255;
  assign n10260 = n9691 & ~n32996;
  assign n10261 = ~n9683 & n10260;
  assign n10262 = ~n9969 & n10261;
  assign n10263 = ~n9691 & ~n33068;
  assign n10264 = ~n10262 & ~n10263;
  assign n10265 = ~n10258 & ~n10259;
  assign n10266 = ~n10253 & ~n33069;
  assign n10267 = ~n10251 & ~n10266;
  assign n10268 = ~n2283 & ~n10267;
  assign n10269 = ~n9697 & ~n9699;
  assign n10270 = ~n9969 & n10269;
  assign n10271 = ~n32998 & ~n10270;
  assign n10272 = ~n9697 & n32998;
  assign n10273 = ~n9699 & n10272;
  assign n10274 = n32998 & n10270;
  assign n10275 = ~n9969 & n10273;
  assign n10276 = ~n10271 & ~n33070;
  assign n10277 = n2283 & ~n10251;
  assign n10278 = ~n10266 & n10277;
  assign n10279 = n2283 & n10267;
  assign n10280 = ~n10276 & ~n33071;
  assign n10281 = ~n10268 & ~n10280;
  assign n10282 = ~n2021 & ~n10281;
  assign n10283 = n2021 & ~n10268;
  assign n10284 = ~n10280 & n10283;
  assign n10285 = ~n9714 & ~n33000;
  assign n10286 = ~n9714 & ~n9969;
  assign n10287 = ~n33000 & n10286;
  assign n10288 = ~n9969 & n10285;
  assign n10289 = n9722 & ~n33072;
  assign n10290 = n9726 & n10286;
  assign n10291 = n9722 & ~n33000;
  assign n10292 = ~n9714 & n10291;
  assign n10293 = ~n9969 & n10292;
  assign n10294 = ~n9722 & ~n33072;
  assign n10295 = ~n10293 & ~n10294;
  assign n10296 = ~n10289 & ~n10290;
  assign n10297 = ~n10284 & ~n33073;
  assign n10298 = ~n10282 & ~n10297;
  assign n10299 = ~n1796 & ~n10298;
  assign n10300 = n1796 & ~n10282;
  assign n10301 = ~n10297 & n10300;
  assign n10302 = n1796 & n10298;
  assign n10303 = ~n9728 & ~n9738;
  assign n10304 = ~n9728 & ~n9969;
  assign n10305 = ~n9738 & n10304;
  assign n10306 = ~n9969 & n10303;
  assign n10307 = n9736 & ~n33075;
  assign n10308 = n9739 & n10304;
  assign n10309 = ~n9728 & n9736;
  assign n10310 = ~n9738 & n10309;
  assign n10311 = ~n9969 & n10310;
  assign n10312 = ~n9736 & ~n33075;
  assign n10313 = ~n10311 & ~n10312;
  assign n10314 = ~n10307 & ~n10308;
  assign n10315 = ~n33074 & ~n33076;
  assign n10316 = ~n10299 & ~n10315;
  assign n10317 = ~n1567 & ~n10316;
  assign n10318 = n1567 & ~n10299;
  assign n10319 = ~n10315 & n10318;
  assign n10320 = ~n9741 & ~n33003;
  assign n10321 = ~n9741 & ~n9969;
  assign n10322 = ~n33003 & n10321;
  assign n10323 = ~n9969 & n10320;
  assign n10324 = n9749 & ~n33077;
  assign n10325 = n9753 & n10321;
  assign n10326 = n9749 & ~n33003;
  assign n10327 = ~n9741 & n10326;
  assign n10328 = ~n9969 & n10327;
  assign n10329 = ~n9749 & ~n33077;
  assign n10330 = ~n10328 & ~n10329;
  assign n10331 = ~n10324 & ~n10325;
  assign n10332 = ~n10319 & ~n33078;
  assign n10333 = ~n10317 & ~n10332;
  assign n10334 = ~n1374 & ~n10333;
  assign n10335 = ~n9755 & ~n9757;
  assign n10336 = ~n9969 & n10335;
  assign n10337 = ~n33005 & ~n10336;
  assign n10338 = ~n9755 & n33005;
  assign n10339 = ~n9757 & n10338;
  assign n10340 = n33005 & n10336;
  assign n10341 = ~n9969 & n10339;
  assign n10342 = ~n10337 & ~n33079;
  assign n10343 = n1374 & ~n10317;
  assign n10344 = ~n10332 & n10343;
  assign n10345 = n1374 & n10333;
  assign n10346 = ~n10342 & ~n33080;
  assign n10347 = ~n10334 & ~n10346;
  assign n10348 = ~n1179 & ~n10347;
  assign n10349 = n1179 & ~n10334;
  assign n10350 = ~n10346 & n10349;
  assign n10351 = ~n9772 & ~n33007;
  assign n10352 = ~n9772 & ~n9969;
  assign n10353 = ~n33007 & n10352;
  assign n10354 = ~n9969 & n10351;
  assign n10355 = n9780 & ~n33081;
  assign n10356 = n9784 & n10352;
  assign n10357 = n9780 & ~n33007;
  assign n10358 = ~n9772 & n10357;
  assign n10359 = ~n9969 & n10358;
  assign n10360 = ~n9780 & ~n33081;
  assign n10361 = ~n10359 & ~n10360;
  assign n10362 = ~n10355 & ~n10356;
  assign n10363 = ~n10350 & ~n33082;
  assign n10364 = ~n10348 & ~n10363;
  assign n10365 = ~n1016 & ~n10364;
  assign n10366 = n1016 & ~n10348;
  assign n10367 = ~n10363 & n10366;
  assign n10368 = n1016 & n10364;
  assign n10369 = ~n9786 & ~n9796;
  assign n10370 = ~n9786 & ~n9969;
  assign n10371 = ~n9796 & n10370;
  assign n10372 = ~n9969 & n10369;
  assign n10373 = n9794 & ~n33084;
  assign n10374 = n9797 & n10370;
  assign n10375 = ~n9786 & n9794;
  assign n10376 = ~n9796 & n10375;
  assign n10377 = ~n9969 & n10376;
  assign n10378 = ~n9794 & ~n33084;
  assign n10379 = ~n10377 & ~n10378;
  assign n10380 = ~n10373 & ~n10374;
  assign n10381 = ~n33083 & ~n33085;
  assign n10382 = ~n10365 & ~n10381;
  assign n10383 = ~n855 & ~n10382;
  assign n10384 = n855 & ~n10365;
  assign n10385 = ~n10381 & n10384;
  assign n10386 = ~n9799 & ~n33010;
  assign n10387 = ~n9799 & ~n9969;
  assign n10388 = ~n33010 & n10387;
  assign n10389 = ~n9969 & n10386;
  assign n10390 = n9807 & ~n33086;
  assign n10391 = n9811 & n10387;
  assign n10392 = n9807 & ~n33010;
  assign n10393 = ~n9799 & n10392;
  assign n10394 = ~n9969 & n10393;
  assign n10395 = ~n9807 & ~n33086;
  assign n10396 = ~n10394 & ~n10395;
  assign n10397 = ~n10390 & ~n10391;
  assign n10398 = ~n10385 & ~n33087;
  assign n10399 = ~n10383 & ~n10398;
  assign n10400 = ~n720 & ~n10399;
  assign n10401 = ~n9813 & ~n9815;
  assign n10402 = ~n9969 & n10401;
  assign n10403 = ~n33012 & ~n10402;
  assign n10404 = ~n9813 & n33012;
  assign n10405 = ~n9815 & n10404;
  assign n10406 = n33012 & n10402;
  assign n10407 = ~n9969 & n10405;
  assign n10408 = ~n10403 & ~n33088;
  assign n10409 = n720 & ~n10383;
  assign n10410 = ~n10398 & n10409;
  assign n10411 = n720 & n10399;
  assign n10412 = ~n10408 & ~n33089;
  assign n10413 = ~n10400 & ~n10412;
  assign n10414 = ~n592 & ~n10413;
  assign n10415 = n592 & ~n10400;
  assign n10416 = ~n10412 & n10415;
  assign n10417 = ~n9830 & ~n33014;
  assign n10418 = ~n9830 & ~n9969;
  assign n10419 = ~n33014 & n10418;
  assign n10420 = ~n9969 & n10417;
  assign n10421 = n9838 & ~n33090;
  assign n10422 = n9842 & n10418;
  assign n10423 = n9838 & ~n33014;
  assign n10424 = ~n9830 & n10423;
  assign n10425 = ~n9969 & n10424;
  assign n10426 = ~n9838 & ~n33090;
  assign n10427 = ~n10425 & ~n10426;
  assign n10428 = ~n10421 & ~n10422;
  assign n10429 = ~n10416 & ~n33091;
  assign n10430 = ~n10414 & ~n10429;
  assign n10431 = ~n487 & ~n10430;
  assign n10432 = n487 & ~n10414;
  assign n10433 = ~n10429 & n10432;
  assign n10434 = n487 & n10430;
  assign n10435 = ~n9844 & ~n9854;
  assign n10436 = ~n9844 & ~n9969;
  assign n10437 = ~n9854 & n10436;
  assign n10438 = ~n9969 & n10435;
  assign n10439 = n9852 & ~n33093;
  assign n10440 = n9855 & n10436;
  assign n10441 = ~n9844 & n9852;
  assign n10442 = ~n9854 & n10441;
  assign n10443 = ~n9969 & n10442;
  assign n10444 = ~n9852 & ~n33093;
  assign n10445 = ~n10443 & ~n10444;
  assign n10446 = ~n10439 & ~n10440;
  assign n10447 = ~n33092 & ~n33094;
  assign n10448 = ~n10431 & ~n10447;
  assign n10449 = ~n393 & ~n10448;
  assign n10450 = n393 & ~n10431;
  assign n10451 = ~n10447 & n10450;
  assign n10452 = ~n9857 & ~n33017;
  assign n10453 = ~n9857 & ~n9969;
  assign n10454 = ~n33017 & n10453;
  assign n10455 = ~n9969 & n10452;
  assign n10456 = n9865 & ~n33095;
  assign n10457 = n9869 & n10453;
  assign n10458 = n9865 & ~n33017;
  assign n10459 = ~n9857 & n10458;
  assign n10460 = ~n9969 & n10459;
  assign n10461 = ~n9865 & ~n33095;
  assign n10462 = ~n10460 & ~n10461;
  assign n10463 = ~n10456 & ~n10457;
  assign n10464 = ~n10451 & ~n33096;
  assign n10465 = ~n10449 & ~n10464;
  assign n10466 = ~n321 & ~n10465;
  assign n10467 = ~n9871 & ~n9873;
  assign n10468 = ~n9969 & n10467;
  assign n10469 = ~n33019 & ~n10468;
  assign n10470 = ~n9871 & n33019;
  assign n10471 = ~n9873 & n10470;
  assign n10472 = n33019 & n10468;
  assign n10473 = ~n9969 & n10471;
  assign n10474 = ~n10469 & ~n33097;
  assign n10475 = n321 & ~n10449;
  assign n10476 = ~n10464 & n10475;
  assign n10477 = n321 & n10465;
  assign n10478 = ~n10474 & ~n33098;
  assign n10479 = ~n10466 & ~n10478;
  assign n10480 = ~n263 & ~n10479;
  assign n10481 = n263 & ~n10466;
  assign n10482 = ~n10478 & n10481;
  assign n10483 = ~n9888 & ~n33021;
  assign n10484 = ~n9888 & ~n9969;
  assign n10485 = ~n33021 & n10484;
  assign n10486 = ~n9969 & n10483;
  assign n10487 = n9896 & ~n33099;
  assign n10488 = n9900 & n10484;
  assign n10489 = n9896 & ~n33021;
  assign n10490 = ~n9888 & n10489;
  assign n10491 = ~n9969 & n10490;
  assign n10492 = ~n9896 & ~n33099;
  assign n10493 = ~n10491 & ~n10492;
  assign n10494 = ~n10487 & ~n10488;
  assign n10495 = ~n10482 & ~n33100;
  assign n10496 = ~n10480 & ~n10495;
  assign n10497 = ~n214 & ~n10496;
  assign n10498 = n214 & ~n10480;
  assign n10499 = ~n10495 & n10498;
  assign n10500 = n214 & n10496;
  assign n10501 = ~n9902 & ~n9912;
  assign n10502 = ~n9902 & ~n9969;
  assign n10503 = ~n9912 & n10502;
  assign n10504 = ~n9969 & n10501;
  assign n10505 = n9910 & ~n33102;
  assign n10506 = n9913 & n10502;
  assign n10507 = ~n9902 & n9910;
  assign n10508 = ~n9912 & n10507;
  assign n10509 = ~n9969 & n10508;
  assign n10510 = ~n9910 & ~n33102;
  assign n10511 = ~n10509 & ~n10510;
  assign n10512 = ~n10505 & ~n10506;
  assign n10513 = ~n33101 & ~n33103;
  assign n10514 = ~n10497 & ~n10513;
  assign n10515 = ~n197 & ~n10514;
  assign n10516 = n197 & ~n10497;
  assign n10517 = ~n10513 & n10516;
  assign n10518 = ~n9915 & ~n33024;
  assign n10519 = ~n9915 & ~n9969;
  assign n10520 = ~n33024 & n10519;
  assign n10521 = ~n9969 & n10518;
  assign n10522 = n9923 & ~n33104;
  assign n10523 = n9927 & n10519;
  assign n10524 = n9923 & ~n33024;
  assign n10525 = ~n9915 & n10524;
  assign n10526 = ~n9969 & n10525;
  assign n10527 = ~n9923 & ~n33104;
  assign n10528 = ~n10526 & ~n10527;
  assign n10529 = ~n10522 & ~n10523;
  assign n10530 = ~n10517 & ~n33105;
  assign n10531 = ~n10515 & ~n10530;
  assign n10532 = ~n9929 & ~n9931;
  assign n10533 = ~n9969 & n10532;
  assign n10534 = ~n33026 & ~n10533;
  assign n10535 = ~n9929 & n33026;
  assign n10536 = ~n9931 & n10535;
  assign n10537 = n33026 & n10533;
  assign n10538 = ~n9969 & n10536;
  assign n10539 = ~n10534 & ~n33106;
  assign n10540 = ~n9945 & ~n9953;
  assign n10541 = ~n9953 & ~n9969;
  assign n10542 = ~n9945 & n10541;
  assign n10543 = ~n9969 & n10540;
  assign n10544 = ~n33029 & ~n33107;
  assign n10545 = ~n10539 & n10544;
  assign n10546 = ~n10531 & n10545;
  assign n10547 = n193 & ~n10546;
  assign n10548 = ~n10515 & n10539;
  assign n10549 = ~n10530 & n10548;
  assign n10550 = n10531 & n10539;
  assign n10551 = n9945 & ~n10541;
  assign n10552 = ~n193 & ~n10540;
  assign n10553 = ~n10551 & n10552;
  assign n10554 = ~n33108 & ~n10553;
  assign n10555 = ~n10547 & n10554;
  assign n10556 = ~n10055 & ~n10057;
  assign n10557 = ~n10555 & n10556;
  assign n10558 = ~n10065 & ~n10557;
  assign n10559 = ~n10057 & n10065;
  assign n10560 = ~n10055 & n10559;
  assign n10561 = n10065 & n10557;
  assign n10562 = ~n10555 & n10560;
  assign n10563 = ~n10558 & ~n33109;
  assign n10564 = ~n10021 & ~n10023;
  assign n10565 = ~n10555 & n10564;
  assign n10566 = ~n33037 & ~n10565;
  assign n10567 = ~n10023 & n33037;
  assign n10568 = ~n10021 & n10567;
  assign n10569 = n33037 & n10565;
  assign n10570 = ~n10555 & n10568;
  assign n10571 = ~n10566 & ~n33110;
  assign n10572 = ~n9994 & ~n9996;
  assign n10573 = ~n10555 & n10572;
  assign n10574 = ~n10005 & ~n10573;
  assign n10575 = ~n9996 & n10005;
  assign n10576 = ~n9994 & n10575;
  assign n10577 = n10005 & n10573;
  assign n10578 = ~n10555 & n10576;
  assign n10579 = ~n10574 & ~n33111;
  assign n10580 = ~pi54  & ~n10555;
  assign n10581 = ~pi55  & n10580;
  assign n10582 = n9971 & ~n10555;
  assign n10583 = ~n9969 & ~n10553;
  assign n10584 = ~n33108 & n10583;
  assign n10585 = ~n10547 & n10584;
  assign n10586 = ~n33112 & ~n10585;
  assign n10587 = pi56  & ~n10586;
  assign n10588 = ~pi56  & ~n10585;
  assign n10589 = ~pi56  & n10586;
  assign n10590 = ~n33112 & n10588;
  assign n10591 = ~n10587 & ~n33113;
  assign n10592 = pi54  & ~n10555;
  assign n10593 = ~pi52  & ~pi53 ;
  assign n10594 = ~pi54  & n10593;
  assign n10595 = ~n9438 & ~n33031;
  assign n10596 = ~n9439 & n10595;
  assign n10597 = ~n9455 & n10596;
  assign n10598 = ~n32967 & n10597;
  assign n10599 = n32965 & n9457;
  assign n10600 = ~n9449 & n10598;
  assign n10601 = ~n10594 & ~n33114;
  assign n10602 = ~n9967 & n10601;
  assign n10603 = ~n33029 & n10602;
  assign n10604 = ~n9961 & n10603;
  assign n10605 = ~n10592 & ~n10594;
  assign n10606 = n9969 & n10605;
  assign n10607 = ~n10592 & n10604;
  assign n10608 = pi55  & ~n10580;
  assign n10609 = ~n33112 & ~n10608;
  assign n10610 = ~n33115 & n10609;
  assign n10611 = ~n9969 & ~n10605;
  assign n10612 = n9457 & ~n10611;
  assign n10613 = ~n10610 & ~n10611;
  assign n10614 = n9457 & n10613;
  assign n10615 = ~n10610 & n10612;
  assign n10616 = ~n10591 & ~n33116;
  assign n10617 = ~n9457 & ~n10613;
  assign n10618 = n8896 & ~n10617;
  assign n10619 = ~n10616 & n10618;
  assign n10620 = ~n9974 & ~n33032;
  assign n10621 = ~n10555 & n10620;
  assign n10622 = n9979 & ~n10621;
  assign n10623 = ~n9979 & n10620;
  assign n10624 = ~n9979 & n10621;
  assign n10625 = ~n10555 & n10623;
  assign n10626 = ~n10622 & ~n33117;
  assign n10627 = ~n10619 & ~n10626;
  assign n10628 = ~n10616 & ~n10617;
  assign n10629 = ~n8896 & ~n10628;
  assign n10630 = n8411 & ~n10629;
  assign n10631 = ~n10627 & ~n10629;
  assign n10632 = n8411 & n10631;
  assign n10633 = ~n10627 & n10630;
  assign n10634 = ~n10579 & ~n33118;
  assign n10635 = ~n8411 & ~n10631;
  assign n10636 = n7885 & ~n10635;
  assign n10637 = ~n10634 & n10636;
  assign n10638 = ~n10008 & ~n33034;
  assign n10639 = ~n10555 & n10638;
  assign n10640 = ~n10018 & ~n10639;
  assign n10641 = ~n10008 & n10018;
  assign n10642 = ~n33034 & n10641;
  assign n10643 = n10018 & n10639;
  assign n10644 = ~n10555 & n10642;
  assign n10645 = n10018 & ~n10639;
  assign n10646 = ~n10018 & n10639;
  assign n10647 = ~n10645 & ~n10646;
  assign n10648 = ~n10640 & ~n33119;
  assign n10649 = ~n10637 & n33120;
  assign n10650 = ~n10634 & ~n10635;
  assign n10651 = ~n7885 & ~n10650;
  assign n10652 = n7428 & ~n10651;
  assign n10653 = ~n10649 & ~n10651;
  assign n10654 = n7428 & n10653;
  assign n10655 = ~n10649 & n10652;
  assign n10656 = ~n10571 & ~n33121;
  assign n10657 = ~n7428 & ~n10653;
  assign n10658 = n6937 & ~n10657;
  assign n10659 = ~n10656 & n10658;
  assign n10660 = ~n10038 & ~n33038;
  assign n10661 = ~n10555 & n10660;
  assign n10662 = ~n33040 & ~n10661;
  assign n10663 = n33040 & n10661;
  assign n10664 = ~n10038 & ~n33040;
  assign n10665 = ~n33038 & n10664;
  assign n10666 = ~n10555 & n10665;
  assign n10667 = n33040 & ~n10661;
  assign n10668 = ~n10666 & ~n10667;
  assign n10669 = ~n10662 & ~n10663;
  assign n10670 = ~n10659 & ~n33122;
  assign n10671 = ~n10656 & ~n10657;
  assign n10672 = ~n6937 & ~n10671;
  assign n10673 = n6507 & ~n10672;
  assign n10674 = ~n10670 & ~n10672;
  assign n10675 = n6507 & n10674;
  assign n10676 = ~n10670 & n10673;
  assign n10677 = ~n10563 & ~n33123;
  assign n10678 = ~n6507 & ~n10674;
  assign n10679 = ~n10677 & ~n10678;
  assign n10680 = ~n6051 & ~n10679;
  assign n10681 = ~n10068 & ~n33043;
  assign n10682 = ~n10555 & n10681;
  assign n10683 = n10076 & ~n10682;
  assign n10684 = ~n10076 & n10682;
  assign n10685 = ~n10068 & n10076;
  assign n10686 = ~n33043 & n10685;
  assign n10687 = ~n10555 & n10686;
  assign n10688 = ~n10076 & ~n10682;
  assign n10689 = ~n10687 & ~n10688;
  assign n10690 = ~n10683 & ~n10684;
  assign n10691 = n6051 & ~n10678;
  assign n10692 = ~n10677 & n10691;
  assign n10693 = ~n33124 & ~n10692;
  assign n10694 = ~n10680 & ~n10693;
  assign n10695 = ~n5648 & ~n10694;
  assign n10696 = ~n10082 & ~n10084;
  assign n10697 = ~n10555 & n10696;
  assign n10698 = ~n33045 & ~n10697;
  assign n10699 = ~n10084 & n33045;
  assign n10700 = ~n10082 & n10699;
  assign n10701 = n33045 & n10697;
  assign n10702 = ~n10555 & n10700;
  assign n10703 = ~n10698 & ~n33125;
  assign n10704 = n5648 & ~n10680;
  assign n10705 = n5648 & n10694;
  assign n10706 = ~n10693 & n10704;
  assign n10707 = ~n10703 & ~n33126;
  assign n10708 = ~n10695 & ~n10707;
  assign n10709 = ~n5223 & ~n10708;
  assign n10710 = n5223 & ~n10695;
  assign n10711 = ~n10707 & n10710;
  assign n10712 = ~n10099 & ~n33046;
  assign n10713 = ~n10555 & n10712;
  assign n10714 = ~n33047 & ~n10713;
  assign n10715 = ~n10099 & n33047;
  assign n10716 = ~n33046 & n10715;
  assign n10717 = n33047 & n10713;
  assign n10718 = ~n10555 & n10716;
  assign n10719 = n33047 & ~n10713;
  assign n10720 = ~n33047 & n10713;
  assign n10721 = ~n10719 & ~n10720;
  assign n10722 = ~n10714 & ~n33127;
  assign n10723 = ~n10711 & n33128;
  assign n10724 = ~n10709 & ~n10723;
  assign n10725 = ~n4851 & ~n10724;
  assign n10726 = ~n10115 & ~n10117;
  assign n10727 = ~n10555 & n10726;
  assign n10728 = ~n33049 & ~n10727;
  assign n10729 = ~n10117 & n33049;
  assign n10730 = ~n10115 & n10729;
  assign n10731 = n33049 & n10727;
  assign n10732 = ~n10555 & n10730;
  assign n10733 = ~n10728 & ~n33129;
  assign n10734 = n4851 & ~n10709;
  assign n10735 = n4851 & n10724;
  assign n10736 = ~n10723 & n10734;
  assign n10737 = ~n10733 & ~n33130;
  assign n10738 = ~n10725 & ~n10737;
  assign n10739 = ~n4461 & ~n10738;
  assign n10740 = n4461 & ~n10725;
  assign n10741 = ~n10737 & n10740;
  assign n10742 = ~n10132 & ~n33050;
  assign n10743 = ~n10132 & ~n10555;
  assign n10744 = ~n33050 & n10743;
  assign n10745 = ~n10555 & n10742;
  assign n10746 = n33052 & ~n33131;
  assign n10747 = n10147 & n10743;
  assign n10748 = ~n33052 & n33131;
  assign n10749 = ~n10132 & n33052;
  assign n10750 = ~n33050 & n10749;
  assign n10751 = ~n10555 & n10750;
  assign n10752 = ~n33052 & ~n33131;
  assign n10753 = ~n10751 & ~n10752;
  assign n10754 = ~n10746 & ~n33132;
  assign n10755 = ~n10741 & ~n33133;
  assign n10756 = ~n10739 & ~n10755;
  assign n10757 = ~n4115 & ~n10756;
  assign n10758 = ~n10149 & ~n10151;
  assign n10759 = ~n10555 & n10758;
  assign n10760 = ~n33054 & ~n10759;
  assign n10761 = ~n10151 & n33054;
  assign n10762 = ~n10149 & n10761;
  assign n10763 = n33054 & n10759;
  assign n10764 = ~n10555 & n10762;
  assign n10765 = ~n10760 & ~n33134;
  assign n10766 = n4115 & ~n10739;
  assign n10767 = n4115 & n10756;
  assign n10768 = ~n10755 & n10766;
  assign n10769 = ~n10765 & ~n33135;
  assign n10770 = ~n10757 & ~n10769;
  assign n10771 = ~n3754 & ~n10770;
  assign n10772 = ~n10166 & ~n33055;
  assign n10773 = ~n10555 & n10772;
  assign n10774 = ~n33058 & ~n10773;
  assign n10775 = ~n10166 & n33058;
  assign n10776 = ~n33055 & n10775;
  assign n10777 = n33058 & n10773;
  assign n10778 = ~n10555 & n10776;
  assign n10779 = ~n10774 & ~n33136;
  assign n10780 = n3754 & ~n10757;
  assign n10781 = ~n10769 & n10780;
  assign n10782 = ~n10779 & ~n10781;
  assign n10783 = ~n10771 & ~n10782;
  assign n10784 = ~n3444 & ~n10783;
  assign n10785 = ~n10185 & ~n10187;
  assign n10786 = ~n10555 & n10785;
  assign n10787 = ~n33060 & ~n10786;
  assign n10788 = ~n10187 & n33060;
  assign n10789 = ~n10185 & n10788;
  assign n10790 = n33060 & n10786;
  assign n10791 = ~n10555 & n10789;
  assign n10792 = ~n10787 & ~n33137;
  assign n10793 = n3444 & ~n10771;
  assign n10794 = n3444 & n10783;
  assign n10795 = ~n10782 & n10793;
  assign n10796 = ~n10792 & ~n33138;
  assign n10797 = ~n10784 & ~n10796;
  assign n10798 = ~n3116 & ~n10797;
  assign n10799 = n3116 & ~n10784;
  assign n10800 = ~n10796 & n10799;
  assign n10801 = ~n10202 & ~n33062;
  assign n10802 = ~n10202 & ~n10555;
  assign n10803 = ~n33062 & n10802;
  assign n10804 = ~n10555 & n10801;
  assign n10805 = n10210 & ~n33139;
  assign n10806 = n10214 & n10802;
  assign n10807 = ~n10202 & n10210;
  assign n10808 = ~n33062 & n10807;
  assign n10809 = ~n10555 & n10808;
  assign n10810 = ~n10210 & ~n33139;
  assign n10811 = ~n10809 & ~n10810;
  assign n10812 = ~n10805 & ~n10806;
  assign n10813 = ~n10800 & ~n33140;
  assign n10814 = ~n10798 & ~n10813;
  assign n10815 = ~n2833 & ~n10814;
  assign n10816 = ~n10216 & ~n10218;
  assign n10817 = ~n10555 & n10816;
  assign n10818 = ~n33064 & ~n10817;
  assign n10819 = ~n10218 & n33064;
  assign n10820 = ~n10216 & n10819;
  assign n10821 = n33064 & n10817;
  assign n10822 = ~n10555 & n10820;
  assign n10823 = ~n10818 & ~n33141;
  assign n10824 = n2833 & ~n10798;
  assign n10825 = n2833 & n10814;
  assign n10826 = ~n10813 & n10824;
  assign n10827 = ~n10823 & ~n33142;
  assign n10828 = ~n10815 & ~n10827;
  assign n10829 = ~n2536 & ~n10828;
  assign n10830 = ~n10233 & ~n33065;
  assign n10831 = ~n10555 & n10830;
  assign n10832 = ~n33067 & ~n10831;
  assign n10833 = ~n10233 & n33067;
  assign n10834 = ~n33065 & n10833;
  assign n10835 = n33067 & n10831;
  assign n10836 = ~n10555 & n10834;
  assign n10837 = ~n10832 & ~n33143;
  assign n10838 = n2536 & ~n10815;
  assign n10839 = ~n10827 & n10838;
  assign n10840 = ~n10837 & ~n10839;
  assign n10841 = ~n10829 & ~n10840;
  assign n10842 = ~n2283 & ~n10841;
  assign n10843 = ~n10251 & ~n10253;
  assign n10844 = ~n10555 & n10843;
  assign n10845 = ~n33069 & ~n10844;
  assign n10846 = ~n10253 & n33069;
  assign n10847 = ~n10251 & n10846;
  assign n10848 = n33069 & n10844;
  assign n10849 = ~n10555 & n10847;
  assign n10850 = ~n10845 & ~n33144;
  assign n10851 = n2283 & ~n10829;
  assign n10852 = n2283 & n10841;
  assign n10853 = ~n10840 & n10851;
  assign n10854 = ~n10850 & ~n33145;
  assign n10855 = ~n10842 & ~n10854;
  assign n10856 = ~n2021 & ~n10855;
  assign n10857 = n2021 & ~n10842;
  assign n10858 = ~n10854 & n10857;
  assign n10859 = ~n10268 & ~n33071;
  assign n10860 = ~n10268 & ~n10555;
  assign n10861 = ~n33071 & n10860;
  assign n10862 = ~n10555 & n10859;
  assign n10863 = n10276 & ~n33146;
  assign n10864 = n10280 & n10860;
  assign n10865 = ~n10268 & n10276;
  assign n10866 = ~n33071 & n10865;
  assign n10867 = ~n10555 & n10866;
  assign n10868 = ~n10276 & ~n33146;
  assign n10869 = ~n10867 & ~n10868;
  assign n10870 = ~n10863 & ~n10864;
  assign n10871 = ~n10858 & ~n33147;
  assign n10872 = ~n10856 & ~n10871;
  assign n10873 = ~n1796 & ~n10872;
  assign n10874 = ~n10282 & ~n10284;
  assign n10875 = ~n10555 & n10874;
  assign n10876 = ~n33073 & ~n10875;
  assign n10877 = ~n10284 & n33073;
  assign n10878 = ~n10282 & n10877;
  assign n10879 = n33073 & n10875;
  assign n10880 = ~n10555 & n10878;
  assign n10881 = ~n10876 & ~n33148;
  assign n10882 = n1796 & ~n10856;
  assign n10883 = n1796 & n10872;
  assign n10884 = ~n10871 & n10882;
  assign n10885 = ~n10881 & ~n33149;
  assign n10886 = ~n10873 & ~n10885;
  assign n10887 = ~n1567 & ~n10886;
  assign n10888 = ~n10299 & ~n33074;
  assign n10889 = ~n10555 & n10888;
  assign n10890 = ~n33076 & ~n10889;
  assign n10891 = ~n10299 & n33076;
  assign n10892 = ~n33074 & n10891;
  assign n10893 = n33076 & n10889;
  assign n10894 = ~n10555 & n10892;
  assign n10895 = ~n10890 & ~n33150;
  assign n10896 = n1567 & ~n10873;
  assign n10897 = ~n10885 & n10896;
  assign n10898 = ~n10895 & ~n10897;
  assign n10899 = ~n10887 & ~n10898;
  assign n10900 = ~n1374 & ~n10899;
  assign n10901 = ~n10317 & ~n10319;
  assign n10902 = ~n10555 & n10901;
  assign n10903 = ~n33078 & ~n10902;
  assign n10904 = ~n10319 & n33078;
  assign n10905 = ~n10317 & n10904;
  assign n10906 = n33078 & n10902;
  assign n10907 = ~n10555 & n10905;
  assign n10908 = ~n10903 & ~n33151;
  assign n10909 = n1374 & ~n10887;
  assign n10910 = n1374 & n10899;
  assign n10911 = ~n10898 & n10909;
  assign n10912 = ~n10908 & ~n33152;
  assign n10913 = ~n10900 & ~n10912;
  assign n10914 = ~n1179 & ~n10913;
  assign n10915 = n1179 & ~n10900;
  assign n10916 = ~n10912 & n10915;
  assign n10917 = ~n10334 & ~n33080;
  assign n10918 = ~n10334 & ~n10555;
  assign n10919 = ~n33080 & n10918;
  assign n10920 = ~n10555 & n10917;
  assign n10921 = n10342 & ~n33153;
  assign n10922 = n10346 & n10918;
  assign n10923 = ~n10334 & n10342;
  assign n10924 = ~n33080 & n10923;
  assign n10925 = ~n10555 & n10924;
  assign n10926 = ~n10342 & ~n33153;
  assign n10927 = ~n10925 & ~n10926;
  assign n10928 = ~n10921 & ~n10922;
  assign n10929 = ~n10916 & ~n33154;
  assign n10930 = ~n10914 & ~n10929;
  assign n10931 = ~n1016 & ~n10930;
  assign n10932 = ~n10348 & ~n10350;
  assign n10933 = ~n10555 & n10932;
  assign n10934 = ~n33082 & ~n10933;
  assign n10935 = ~n10350 & n33082;
  assign n10936 = ~n10348 & n10935;
  assign n10937 = n33082 & n10933;
  assign n10938 = ~n10555 & n10936;
  assign n10939 = ~n10934 & ~n33155;
  assign n10940 = n1016 & ~n10914;
  assign n10941 = n1016 & n10930;
  assign n10942 = ~n10929 & n10940;
  assign n10943 = ~n10939 & ~n33156;
  assign n10944 = ~n10931 & ~n10943;
  assign n10945 = ~n855 & ~n10944;
  assign n10946 = ~n10365 & ~n33083;
  assign n10947 = ~n10555 & n10946;
  assign n10948 = ~n33085 & ~n10947;
  assign n10949 = ~n10365 & n33085;
  assign n10950 = ~n33083 & n10949;
  assign n10951 = n33085 & n10947;
  assign n10952 = ~n10555 & n10950;
  assign n10953 = ~n10948 & ~n33157;
  assign n10954 = n855 & ~n10931;
  assign n10955 = ~n10943 & n10954;
  assign n10956 = ~n10953 & ~n10955;
  assign n10957 = ~n10945 & ~n10956;
  assign n10958 = ~n720 & ~n10957;
  assign n10959 = ~n10383 & ~n10385;
  assign n10960 = ~n10555 & n10959;
  assign n10961 = ~n33087 & ~n10960;
  assign n10962 = ~n10385 & n33087;
  assign n10963 = ~n10383 & n10962;
  assign n10964 = n33087 & n10960;
  assign n10965 = ~n10555 & n10963;
  assign n10966 = ~n10961 & ~n33158;
  assign n10967 = n720 & ~n10945;
  assign n10968 = n720 & n10957;
  assign n10969 = ~n10956 & n10967;
  assign n10970 = ~n10966 & ~n33159;
  assign n10971 = ~n10958 & ~n10970;
  assign n10972 = ~n592 & ~n10971;
  assign n10973 = n592 & ~n10958;
  assign n10974 = ~n10970 & n10973;
  assign n10975 = ~n10400 & ~n33089;
  assign n10976 = ~n10400 & ~n10555;
  assign n10977 = ~n33089 & n10976;
  assign n10978 = ~n10555 & n10975;
  assign n10979 = n10408 & ~n33160;
  assign n10980 = n10412 & n10976;
  assign n10981 = ~n10400 & n10408;
  assign n10982 = ~n33089 & n10981;
  assign n10983 = ~n10555 & n10982;
  assign n10984 = ~n10408 & ~n33160;
  assign n10985 = ~n10983 & ~n10984;
  assign n10986 = ~n10979 & ~n10980;
  assign n10987 = ~n10974 & ~n33161;
  assign n10988 = ~n10972 & ~n10987;
  assign n10989 = ~n487 & ~n10988;
  assign n10990 = ~n10414 & ~n10416;
  assign n10991 = ~n10555 & n10990;
  assign n10992 = ~n33091 & ~n10991;
  assign n10993 = ~n10416 & n33091;
  assign n10994 = ~n10414 & n10993;
  assign n10995 = n33091 & n10991;
  assign n10996 = ~n10555 & n10994;
  assign n10997 = ~n10992 & ~n33162;
  assign n10998 = n487 & ~n10972;
  assign n10999 = n487 & n10988;
  assign n11000 = ~n10987 & n10998;
  assign n11001 = ~n10997 & ~n33163;
  assign n11002 = ~n10989 & ~n11001;
  assign n11003 = ~n393 & ~n11002;
  assign n11004 = ~n10431 & ~n33092;
  assign n11005 = ~n10555 & n11004;
  assign n11006 = ~n33094 & ~n11005;
  assign n11007 = ~n10431 & n33094;
  assign n11008 = ~n33092 & n11007;
  assign n11009 = n33094 & n11005;
  assign n11010 = ~n10555 & n11008;
  assign n11011 = ~n11006 & ~n33164;
  assign n11012 = n393 & ~n10989;
  assign n11013 = ~n11001 & n11012;
  assign n11014 = ~n11011 & ~n11013;
  assign n11015 = ~n11003 & ~n11014;
  assign n11016 = ~n321 & ~n11015;
  assign n11017 = ~n10449 & ~n10451;
  assign n11018 = ~n10555 & n11017;
  assign n11019 = ~n33096 & ~n11018;
  assign n11020 = ~n10451 & n33096;
  assign n11021 = ~n10449 & n11020;
  assign n11022 = n33096 & n11018;
  assign n11023 = ~n10555 & n11021;
  assign n11024 = ~n11019 & ~n33165;
  assign n11025 = n321 & ~n11003;
  assign n11026 = n321 & n11015;
  assign n11027 = ~n11014 & n11025;
  assign n11028 = ~n11024 & ~n33166;
  assign n11029 = ~n11016 & ~n11028;
  assign n11030 = ~n263 & ~n11029;
  assign n11031 = n263 & ~n11016;
  assign n11032 = ~n11028 & n11031;
  assign n11033 = ~n10466 & ~n33098;
  assign n11034 = ~n10466 & ~n10555;
  assign n11035 = ~n33098 & n11034;
  assign n11036 = ~n10555 & n11033;
  assign n11037 = n10474 & ~n33167;
  assign n11038 = n10478 & n11034;
  assign n11039 = ~n10466 & n10474;
  assign n11040 = ~n33098 & n11039;
  assign n11041 = ~n10555 & n11040;
  assign n11042 = ~n10474 & ~n33167;
  assign n11043 = ~n11041 & ~n11042;
  assign n11044 = ~n11037 & ~n11038;
  assign n11045 = ~n11032 & ~n33168;
  assign n11046 = ~n11030 & ~n11045;
  assign n11047 = ~n214 & ~n11046;
  assign n11048 = ~n10480 & ~n10482;
  assign n11049 = ~n10555 & n11048;
  assign n11050 = ~n33100 & ~n11049;
  assign n11051 = ~n10482 & n33100;
  assign n11052 = ~n10480 & n11051;
  assign n11053 = n33100 & n11049;
  assign n11054 = ~n10555 & n11052;
  assign n11055 = ~n11050 & ~n33169;
  assign n11056 = n214 & ~n11030;
  assign n11057 = n214 & n11046;
  assign n11058 = ~n11045 & n11056;
  assign n11059 = ~n11055 & ~n33170;
  assign n11060 = ~n11047 & ~n11059;
  assign n11061 = ~n197 & ~n11060;
  assign n11062 = ~n10497 & ~n33101;
  assign n11063 = ~n10555 & n11062;
  assign n11064 = ~n33103 & ~n11063;
  assign n11065 = ~n10497 & n33103;
  assign n11066 = ~n33101 & n11065;
  assign n11067 = n33103 & n11063;
  assign n11068 = ~n10555 & n11066;
  assign n11069 = ~n11064 & ~n33171;
  assign n11070 = n197 & ~n11047;
  assign n11071 = ~n11059 & n11070;
  assign n11072 = ~n11069 & ~n11071;
  assign n11073 = ~n11061 & ~n11072;
  assign n11074 = ~n10515 & ~n10517;
  assign n11075 = ~n10555 & n11074;
  assign n11076 = ~n33105 & ~n11075;
  assign n11077 = ~n10517 & n33105;
  assign n11078 = ~n10515 & n11077;
  assign n11079 = n33105 & n11075;
  assign n11080 = ~n10555 & n11078;
  assign n11081 = ~n11076 & ~n33172;
  assign n11082 = ~n10531 & ~n10539;
  assign n11083 = ~n10539 & ~n10555;
  assign n11084 = ~n10531 & n11083;
  assign n11085 = ~n10555 & n11082;
  assign n11086 = ~n33108 & ~n33173;
  assign n11087 = ~n11081 & n11086;
  assign n11088 = ~n11073 & n11087;
  assign n11089 = n193 & ~n11088;
  assign n11090 = ~n11061 & n11081;
  assign n11091 = n11073 & n11081;
  assign n11092 = ~n11072 & n11090;
  assign n11093 = n10531 & ~n11083;
  assign n11094 = ~n193 & ~n11082;
  assign n11095 = ~n11093 & n11094;
  assign n11096 = ~n33174 & ~n11095;
  assign n11097 = ~n11089 & n11096;
  assign n11098 = pi52  & ~n11097;
  assign n11099 = ~pi50  & ~pi51 ;
  assign n11100 = ~pi52  & n11099;
  assign n11101 = ~n11098 & ~n11100;
  assign n11102 = ~n10555 & ~n11101;
  assign n11103 = ~pi52  & ~n11097;
  assign n11104 = pi53  & ~n11103;
  assign n11105 = ~pi53  & n11103;
  assign n11106 = n10593 & ~n11097;
  assign n11107 = ~n11104 & ~n33175;
  assign n11108 = ~n33027 & ~n33114;
  assign n11109 = ~n9948 & n11108;
  assign n11110 = ~n9967 & n11109;
  assign n11111 = ~n33029 & n11110;
  assign n11112 = n9953 & n9969;
  assign n11113 = ~n9961 & n11111;
  assign n11114 = ~n11100 & ~n33176;
  assign n11115 = ~n10553 & n11114;
  assign n11116 = ~n33108 & n11115;
  assign n11117 = ~n10547 & n11116;
  assign n11118 = n10555 & n11101;
  assign n11119 = ~n11098 & n11117;
  assign n11120 = n11107 & ~n33177;
  assign n11121 = ~n11102 & ~n11120;
  assign n11122 = ~n9969 & ~n11121;
  assign n11123 = n9969 & ~n11102;
  assign n11124 = ~n11120 & n11123;
  assign n11125 = ~n10555 & ~n11095;
  assign n11126 = ~n33174 & n11125;
  assign n11127 = ~n11089 & n11126;
  assign n11128 = ~n33175 & ~n11127;
  assign n11129 = pi54  & ~n11128;
  assign n11130 = ~pi54  & ~n11127;
  assign n11131 = ~pi54  & n11128;
  assign n11132 = ~n33175 & n11130;
  assign n11133 = ~n11129 & ~n33178;
  assign n11134 = ~n11124 & ~n11133;
  assign n11135 = ~n11122 & ~n11134;
  assign n11136 = ~n9457 & ~n11135;
  assign n11137 = n9457 & ~n11122;
  assign n11138 = ~n11134 & n11137;
  assign n11139 = n9457 & n11135;
  assign n11140 = ~n33115 & ~n10611;
  assign n11141 = ~n11097 & n11140;
  assign n11142 = n10609 & ~n11141;
  assign n11143 = ~n10609 & n11140;
  assign n11144 = ~n10609 & n11141;
  assign n11145 = ~n11097 & n11143;
  assign n11146 = ~n11142 & ~n33180;
  assign n11147 = ~n33179 & ~n11146;
  assign n11148 = ~n11136 & ~n11147;
  assign n11149 = ~n8896 & ~n11148;
  assign n11150 = n8896 & ~n11136;
  assign n11151 = ~n11147 & n11150;
  assign n11152 = ~n33116 & ~n10617;
  assign n11153 = ~n10617 & ~n11097;
  assign n11154 = ~n33116 & n11153;
  assign n11155 = ~n11097 & n11152;
  assign n11156 = n10591 & ~n33181;
  assign n11157 = n10616 & n11153;
  assign n11158 = n10591 & ~n33116;
  assign n11159 = ~n10617 & n11158;
  assign n11160 = ~n11097 & n11159;
  assign n11161 = ~n10591 & ~n33181;
  assign n11162 = ~n11160 & ~n11161;
  assign n11163 = ~n11156 & ~n11157;
  assign n11164 = ~n11151 & ~n33182;
  assign n11165 = ~n11149 & ~n11164;
  assign n11166 = ~n8411 & ~n11165;
  assign n11167 = n8411 & ~n11149;
  assign n11168 = ~n11164 & n11167;
  assign n11169 = n8411 & n11165;
  assign n11170 = ~n10619 & ~n10629;
  assign n11171 = ~n11097 & n11170;
  assign n11172 = ~n10626 & ~n11171;
  assign n11173 = n10626 & ~n10629;
  assign n11174 = ~n10619 & n11173;
  assign n11175 = n10626 & n11171;
  assign n11176 = ~n11097 & n11174;
  assign n11177 = n10626 & ~n11171;
  assign n11178 = ~n10626 & n11171;
  assign n11179 = ~n11177 & ~n11178;
  assign n11180 = ~n11172 & ~n33184;
  assign n11181 = ~n33183 & n33185;
  assign n11182 = ~n11166 & ~n11181;
  assign n11183 = ~n7885 & ~n11182;
  assign n11184 = n7885 & ~n11166;
  assign n11185 = ~n11181 & n11184;
  assign n11186 = ~n33118 & ~n10635;
  assign n11187 = ~n10635 & ~n11097;
  assign n11188 = ~n33118 & n11187;
  assign n11189 = ~n11097 & n11186;
  assign n11190 = n10579 & ~n33186;
  assign n11191 = n10634 & n11187;
  assign n11192 = n10579 & ~n33118;
  assign n11193 = ~n10635 & n11192;
  assign n11194 = ~n11097 & n11193;
  assign n11195 = ~n10579 & ~n33186;
  assign n11196 = ~n11194 & ~n11195;
  assign n11197 = ~n11190 & ~n11191;
  assign n11198 = ~n11185 & ~n33187;
  assign n11199 = ~n11183 & ~n11198;
  assign n11200 = ~n7428 & ~n11199;
  assign n11201 = n7428 & ~n11183;
  assign n11202 = ~n11198 & n11201;
  assign n11203 = n7428 & n11199;
  assign n11204 = ~n10637 & ~n10651;
  assign n11205 = ~n11097 & n11204;
  assign n11206 = ~n33120 & ~n11205;
  assign n11207 = n33120 & n11205;
  assign n11208 = ~n33120 & ~n10651;
  assign n11209 = ~n10637 & n11208;
  assign n11210 = ~n11097 & n11209;
  assign n11211 = n33120 & ~n11205;
  assign n11212 = ~n11210 & ~n11211;
  assign n11213 = ~n11206 & ~n11207;
  assign n11214 = ~n33188 & ~n33189;
  assign n11215 = ~n11200 & ~n11214;
  assign n11216 = ~n6937 & ~n11215;
  assign n11217 = n6937 & ~n11200;
  assign n11218 = ~n11214 & n11217;
  assign n11219 = ~n33121 & ~n10657;
  assign n11220 = ~n10657 & ~n11097;
  assign n11221 = ~n33121 & n11220;
  assign n11222 = ~n11097 & n11219;
  assign n11223 = n10571 & ~n33190;
  assign n11224 = n10656 & n11220;
  assign n11225 = n10571 & ~n33121;
  assign n11226 = ~n10657 & n11225;
  assign n11227 = ~n11097 & n11226;
  assign n11228 = ~n10571 & ~n33190;
  assign n11229 = ~n11227 & ~n11228;
  assign n11230 = ~n11223 & ~n11224;
  assign n11231 = ~n11218 & ~n33191;
  assign n11232 = ~n11216 & ~n11231;
  assign n11233 = ~n6507 & ~n11232;
  assign n11234 = n6507 & ~n11216;
  assign n11235 = ~n11231 & n11234;
  assign n11236 = n6507 & n11232;
  assign n11237 = ~n10659 & ~n10672;
  assign n11238 = ~n11097 & n11237;
  assign n11239 = ~n33122 & n11238;
  assign n11240 = n33122 & ~n11238;
  assign n11241 = n33122 & ~n10672;
  assign n11242 = ~n10659 & n11241;
  assign n11243 = ~n11097 & n11242;
  assign n11244 = ~n33122 & ~n11238;
  assign n11245 = ~n11243 & ~n11244;
  assign n11246 = ~n11239 & ~n11240;
  assign n11247 = ~n33192 & ~n33193;
  assign n11248 = ~n11233 & ~n11247;
  assign n11249 = ~n6051 & ~n11248;
  assign n11250 = n6051 & ~n11233;
  assign n11251 = ~n11247 & n11250;
  assign n11252 = ~n33123 & ~n10678;
  assign n11253 = ~n11097 & n11252;
  assign n11254 = n10563 & ~n11253;
  assign n11255 = ~n10563 & n11253;
  assign n11256 = n10563 & ~n33123;
  assign n11257 = ~n10678 & n11256;
  assign n11258 = ~n11097 & n11257;
  assign n11259 = ~n10563 & ~n11253;
  assign n11260 = ~n11258 & ~n11259;
  assign n11261 = ~n11254 & ~n11255;
  assign n11262 = ~n11251 & ~n33194;
  assign n11263 = ~n11249 & ~n11262;
  assign n11264 = ~n5648 & ~n11263;
  assign n11265 = ~n10680 & ~n10692;
  assign n11266 = ~n11097 & n11265;
  assign n11267 = ~n33124 & n11266;
  assign n11268 = n33124 & ~n11266;
  assign n11269 = ~n10680 & n33124;
  assign n11270 = ~n10692 & n11269;
  assign n11271 = ~n11097 & n11270;
  assign n11272 = ~n33124 & ~n11266;
  assign n11273 = ~n11271 & ~n11272;
  assign n11274 = ~n11267 & ~n11268;
  assign n11275 = n5648 & ~n11249;
  assign n11276 = ~n11262 & n11275;
  assign n11277 = n5648 & n11263;
  assign n11278 = ~n33195 & ~n33196;
  assign n11279 = ~n11264 & ~n11278;
  assign n11280 = ~n5223 & ~n11279;
  assign n11281 = n5223 & ~n11264;
  assign n11282 = ~n11278 & n11281;
  assign n11283 = ~n10695 & ~n33126;
  assign n11284 = ~n10695 & ~n11097;
  assign n11285 = ~n33126 & n11284;
  assign n11286 = ~n11097 & n11283;
  assign n11287 = n10703 & ~n33197;
  assign n11288 = n10707 & n11284;
  assign n11289 = n10703 & ~n33126;
  assign n11290 = ~n10695 & n11289;
  assign n11291 = ~n11097 & n11290;
  assign n11292 = ~n10703 & ~n33197;
  assign n11293 = ~n11291 & ~n11292;
  assign n11294 = ~n11287 & ~n11288;
  assign n11295 = ~n11282 & ~n33198;
  assign n11296 = ~n11280 & ~n11295;
  assign n11297 = ~n4851 & ~n11296;
  assign n11298 = n4851 & ~n11280;
  assign n11299 = ~n11295 & n11298;
  assign n11300 = n4851 & n11296;
  assign n11301 = ~n10709 & ~n10711;
  assign n11302 = ~n11097 & n11301;
  assign n11303 = ~n33128 & ~n11302;
  assign n11304 = n33128 & n11302;
  assign n11305 = n33128 & ~n11302;
  assign n11306 = ~n10709 & ~n33128;
  assign n11307 = ~n10711 & n11306;
  assign n11308 = ~n33128 & n11302;
  assign n11309 = ~n11097 & n11307;
  assign n11310 = ~n11305 & ~n33200;
  assign n11311 = ~n11303 & ~n11304;
  assign n11312 = ~n33199 & ~n33201;
  assign n11313 = ~n11297 & ~n11312;
  assign n11314 = ~n4461 & ~n11313;
  assign n11315 = n4461 & ~n11297;
  assign n11316 = ~n11312 & n11315;
  assign n11317 = ~n10725 & ~n33130;
  assign n11318 = ~n10725 & ~n11097;
  assign n11319 = ~n33130 & n11318;
  assign n11320 = ~n11097 & n11317;
  assign n11321 = n10733 & ~n33202;
  assign n11322 = n10737 & n11318;
  assign n11323 = n10733 & ~n33130;
  assign n11324 = ~n10725 & n11323;
  assign n11325 = ~n11097 & n11324;
  assign n11326 = ~n10733 & ~n33202;
  assign n11327 = ~n11325 & ~n11326;
  assign n11328 = ~n11321 & ~n11322;
  assign n11329 = ~n11316 & ~n33203;
  assign n11330 = ~n11314 & ~n11329;
  assign n11331 = ~n4115 & ~n11330;
  assign n11332 = ~n10739 & ~n10741;
  assign n11333 = ~n11097 & n11332;
  assign n11334 = ~n33133 & ~n11333;
  assign n11335 = ~n10739 & n33133;
  assign n11336 = ~n10741 & n11335;
  assign n11337 = n33133 & n11333;
  assign n11338 = ~n11097 & n11336;
  assign n11339 = ~n11334 & ~n33204;
  assign n11340 = n4115 & ~n11314;
  assign n11341 = ~n11329 & n11340;
  assign n11342 = n4115 & n11330;
  assign n11343 = ~n11339 & ~n33205;
  assign n11344 = ~n11331 & ~n11343;
  assign n11345 = ~n3754 & ~n11344;
  assign n11346 = n3754 & ~n11331;
  assign n11347 = ~n11343 & n11346;
  assign n11348 = ~n10757 & ~n33135;
  assign n11349 = ~n10757 & ~n11097;
  assign n11350 = ~n33135 & n11349;
  assign n11351 = ~n11097 & n11348;
  assign n11352 = n10765 & ~n33206;
  assign n11353 = n10769 & n11349;
  assign n11354 = n10765 & ~n33135;
  assign n11355 = ~n10757 & n11354;
  assign n11356 = ~n11097 & n11355;
  assign n11357 = ~n10765 & ~n33206;
  assign n11358 = ~n11356 & ~n11357;
  assign n11359 = ~n11352 & ~n11353;
  assign n11360 = ~n11347 & ~n33207;
  assign n11361 = ~n11345 & ~n11360;
  assign n11362 = ~n3444 & ~n11361;
  assign n11363 = n3444 & ~n11345;
  assign n11364 = ~n11360 & n11363;
  assign n11365 = n3444 & n11361;
  assign n11366 = ~n10771 & ~n10781;
  assign n11367 = ~n10771 & ~n11097;
  assign n11368 = ~n10781 & n11367;
  assign n11369 = ~n11097 & n11366;
  assign n11370 = n10779 & ~n33209;
  assign n11371 = n10782 & n11367;
  assign n11372 = ~n10771 & n10779;
  assign n11373 = ~n10781 & n11372;
  assign n11374 = ~n11097 & n11373;
  assign n11375 = ~n10779 & ~n33209;
  assign n11376 = ~n11374 & ~n11375;
  assign n11377 = ~n11370 & ~n11371;
  assign n11378 = ~n33208 & ~n33210;
  assign n11379 = ~n11362 & ~n11378;
  assign n11380 = ~n3116 & ~n11379;
  assign n11381 = n3116 & ~n11362;
  assign n11382 = ~n11378 & n11381;
  assign n11383 = ~n10784 & ~n33138;
  assign n11384 = ~n10784 & ~n11097;
  assign n11385 = ~n33138 & n11384;
  assign n11386 = ~n11097 & n11383;
  assign n11387 = n10792 & ~n33211;
  assign n11388 = n10796 & n11384;
  assign n11389 = n10792 & ~n33138;
  assign n11390 = ~n10784 & n11389;
  assign n11391 = ~n11097 & n11390;
  assign n11392 = ~n10792 & ~n33211;
  assign n11393 = ~n11391 & ~n11392;
  assign n11394 = ~n11387 & ~n11388;
  assign n11395 = ~n11382 & ~n33212;
  assign n11396 = ~n11380 & ~n11395;
  assign n11397 = ~n2833 & ~n11396;
  assign n11398 = ~n10798 & ~n10800;
  assign n11399 = ~n11097 & n11398;
  assign n11400 = ~n33140 & ~n11399;
  assign n11401 = ~n10798 & n33140;
  assign n11402 = ~n10800 & n11401;
  assign n11403 = n33140 & n11399;
  assign n11404 = ~n11097 & n11402;
  assign n11405 = ~n11400 & ~n33213;
  assign n11406 = n2833 & ~n11380;
  assign n11407 = ~n11395 & n11406;
  assign n11408 = n2833 & n11396;
  assign n11409 = ~n11405 & ~n33214;
  assign n11410 = ~n11397 & ~n11409;
  assign n11411 = ~n2536 & ~n11410;
  assign n11412 = n2536 & ~n11397;
  assign n11413 = ~n11409 & n11412;
  assign n11414 = ~n10815 & ~n33142;
  assign n11415 = ~n10815 & ~n11097;
  assign n11416 = ~n33142 & n11415;
  assign n11417 = ~n11097 & n11414;
  assign n11418 = n10823 & ~n33215;
  assign n11419 = n10827 & n11415;
  assign n11420 = n10823 & ~n33142;
  assign n11421 = ~n10815 & n11420;
  assign n11422 = ~n11097 & n11421;
  assign n11423 = ~n10823 & ~n33215;
  assign n11424 = ~n11422 & ~n11423;
  assign n11425 = ~n11418 & ~n11419;
  assign n11426 = ~n11413 & ~n33216;
  assign n11427 = ~n11411 & ~n11426;
  assign n11428 = ~n2283 & ~n11427;
  assign n11429 = n2283 & ~n11411;
  assign n11430 = ~n11426 & n11429;
  assign n11431 = n2283 & n11427;
  assign n11432 = ~n10829 & ~n10839;
  assign n11433 = ~n10829 & ~n11097;
  assign n11434 = ~n10839 & n11433;
  assign n11435 = ~n11097 & n11432;
  assign n11436 = n10837 & ~n33218;
  assign n11437 = n10840 & n11433;
  assign n11438 = ~n10829 & n10837;
  assign n11439 = ~n10839 & n11438;
  assign n11440 = ~n11097 & n11439;
  assign n11441 = ~n10837 & ~n33218;
  assign n11442 = ~n11440 & ~n11441;
  assign n11443 = ~n11436 & ~n11437;
  assign n11444 = ~n33217 & ~n33219;
  assign n11445 = ~n11428 & ~n11444;
  assign n11446 = ~n2021 & ~n11445;
  assign n11447 = n2021 & ~n11428;
  assign n11448 = ~n11444 & n11447;
  assign n11449 = ~n10842 & ~n33145;
  assign n11450 = ~n10842 & ~n11097;
  assign n11451 = ~n33145 & n11450;
  assign n11452 = ~n11097 & n11449;
  assign n11453 = n10850 & ~n33220;
  assign n11454 = n10854 & n11450;
  assign n11455 = n10850 & ~n33145;
  assign n11456 = ~n10842 & n11455;
  assign n11457 = ~n11097 & n11456;
  assign n11458 = ~n10850 & ~n33220;
  assign n11459 = ~n11457 & ~n11458;
  assign n11460 = ~n11453 & ~n11454;
  assign n11461 = ~n11448 & ~n33221;
  assign n11462 = ~n11446 & ~n11461;
  assign n11463 = ~n1796 & ~n11462;
  assign n11464 = ~n10856 & ~n10858;
  assign n11465 = ~n11097 & n11464;
  assign n11466 = ~n33147 & ~n11465;
  assign n11467 = ~n10856 & n33147;
  assign n11468 = ~n10858 & n11467;
  assign n11469 = n33147 & n11465;
  assign n11470 = ~n11097 & n11468;
  assign n11471 = ~n11466 & ~n33222;
  assign n11472 = n1796 & ~n11446;
  assign n11473 = ~n11461 & n11472;
  assign n11474 = n1796 & n11462;
  assign n11475 = ~n11471 & ~n33223;
  assign n11476 = ~n11463 & ~n11475;
  assign n11477 = ~n1567 & ~n11476;
  assign n11478 = n1567 & ~n11463;
  assign n11479 = ~n11475 & n11478;
  assign n11480 = ~n10873 & ~n33149;
  assign n11481 = ~n10873 & ~n11097;
  assign n11482 = ~n33149 & n11481;
  assign n11483 = ~n11097 & n11480;
  assign n11484 = n10881 & ~n33224;
  assign n11485 = n10885 & n11481;
  assign n11486 = n10881 & ~n33149;
  assign n11487 = ~n10873 & n11486;
  assign n11488 = ~n11097 & n11487;
  assign n11489 = ~n10881 & ~n33224;
  assign n11490 = ~n11488 & ~n11489;
  assign n11491 = ~n11484 & ~n11485;
  assign n11492 = ~n11479 & ~n33225;
  assign n11493 = ~n11477 & ~n11492;
  assign n11494 = ~n1374 & ~n11493;
  assign n11495 = n1374 & ~n11477;
  assign n11496 = ~n11492 & n11495;
  assign n11497 = n1374 & n11493;
  assign n11498 = ~n10887 & ~n10897;
  assign n11499 = ~n10887 & ~n11097;
  assign n11500 = ~n10897 & n11499;
  assign n11501 = ~n11097 & n11498;
  assign n11502 = n10895 & ~n33227;
  assign n11503 = n10898 & n11499;
  assign n11504 = ~n10887 & n10895;
  assign n11505 = ~n10897 & n11504;
  assign n11506 = ~n11097 & n11505;
  assign n11507 = ~n10895 & ~n33227;
  assign n11508 = ~n11506 & ~n11507;
  assign n11509 = ~n11502 & ~n11503;
  assign n11510 = ~n33226 & ~n33228;
  assign n11511 = ~n11494 & ~n11510;
  assign n11512 = ~n1179 & ~n11511;
  assign n11513 = n1179 & ~n11494;
  assign n11514 = ~n11510 & n11513;
  assign n11515 = ~n10900 & ~n33152;
  assign n11516 = ~n10900 & ~n11097;
  assign n11517 = ~n33152 & n11516;
  assign n11518 = ~n11097 & n11515;
  assign n11519 = n10908 & ~n33229;
  assign n11520 = n10912 & n11516;
  assign n11521 = n10908 & ~n33152;
  assign n11522 = ~n10900 & n11521;
  assign n11523 = ~n11097 & n11522;
  assign n11524 = ~n10908 & ~n33229;
  assign n11525 = ~n11523 & ~n11524;
  assign n11526 = ~n11519 & ~n11520;
  assign n11527 = ~n11514 & ~n33230;
  assign n11528 = ~n11512 & ~n11527;
  assign n11529 = ~n1016 & ~n11528;
  assign n11530 = ~n10914 & ~n10916;
  assign n11531 = ~n11097 & n11530;
  assign n11532 = ~n33154 & ~n11531;
  assign n11533 = ~n10914 & n33154;
  assign n11534 = ~n10916 & n11533;
  assign n11535 = n33154 & n11531;
  assign n11536 = ~n11097 & n11534;
  assign n11537 = ~n11532 & ~n33231;
  assign n11538 = n1016 & ~n11512;
  assign n11539 = ~n11527 & n11538;
  assign n11540 = n1016 & n11528;
  assign n11541 = ~n11537 & ~n33232;
  assign n11542 = ~n11529 & ~n11541;
  assign n11543 = ~n855 & ~n11542;
  assign n11544 = n855 & ~n11529;
  assign n11545 = ~n11541 & n11544;
  assign n11546 = ~n10931 & ~n33156;
  assign n11547 = ~n10931 & ~n11097;
  assign n11548 = ~n33156 & n11547;
  assign n11549 = ~n11097 & n11546;
  assign n11550 = n10939 & ~n33233;
  assign n11551 = n10943 & n11547;
  assign n11552 = n10939 & ~n33156;
  assign n11553 = ~n10931 & n11552;
  assign n11554 = ~n11097 & n11553;
  assign n11555 = ~n10939 & ~n33233;
  assign n11556 = ~n11554 & ~n11555;
  assign n11557 = ~n11550 & ~n11551;
  assign n11558 = ~n11545 & ~n33234;
  assign n11559 = ~n11543 & ~n11558;
  assign n11560 = ~n720 & ~n11559;
  assign n11561 = n720 & ~n11543;
  assign n11562 = ~n11558 & n11561;
  assign n11563 = n720 & n11559;
  assign n11564 = ~n10945 & ~n10955;
  assign n11565 = ~n10945 & ~n11097;
  assign n11566 = ~n10955 & n11565;
  assign n11567 = ~n11097 & n11564;
  assign n11568 = n10953 & ~n33236;
  assign n11569 = n10956 & n11565;
  assign n11570 = ~n10945 & n10953;
  assign n11571 = ~n10955 & n11570;
  assign n11572 = ~n11097 & n11571;
  assign n11573 = ~n10953 & ~n33236;
  assign n11574 = ~n11572 & ~n11573;
  assign n11575 = ~n11568 & ~n11569;
  assign n11576 = ~n33235 & ~n33237;
  assign n11577 = ~n11560 & ~n11576;
  assign n11578 = ~n592 & ~n11577;
  assign n11579 = n592 & ~n11560;
  assign n11580 = ~n11576 & n11579;
  assign n11581 = ~n10958 & ~n33159;
  assign n11582 = ~n10958 & ~n11097;
  assign n11583 = ~n33159 & n11582;
  assign n11584 = ~n11097 & n11581;
  assign n11585 = n10966 & ~n33238;
  assign n11586 = n10970 & n11582;
  assign n11587 = n10966 & ~n33159;
  assign n11588 = ~n10958 & n11587;
  assign n11589 = ~n11097 & n11588;
  assign n11590 = ~n10966 & ~n33238;
  assign n11591 = ~n11589 & ~n11590;
  assign n11592 = ~n11585 & ~n11586;
  assign n11593 = ~n11580 & ~n33239;
  assign n11594 = ~n11578 & ~n11593;
  assign n11595 = ~n487 & ~n11594;
  assign n11596 = ~n10972 & ~n10974;
  assign n11597 = ~n11097 & n11596;
  assign n11598 = ~n33161 & ~n11597;
  assign n11599 = ~n10972 & n33161;
  assign n11600 = ~n10974 & n11599;
  assign n11601 = n33161 & n11597;
  assign n11602 = ~n11097 & n11600;
  assign n11603 = ~n11598 & ~n33240;
  assign n11604 = n487 & ~n11578;
  assign n11605 = ~n11593 & n11604;
  assign n11606 = n487 & n11594;
  assign n11607 = ~n11603 & ~n33241;
  assign n11608 = ~n11595 & ~n11607;
  assign n11609 = ~n393 & ~n11608;
  assign n11610 = n393 & ~n11595;
  assign n11611 = ~n11607 & n11610;
  assign n11612 = ~n10989 & ~n33163;
  assign n11613 = ~n10989 & ~n11097;
  assign n11614 = ~n33163 & n11613;
  assign n11615 = ~n11097 & n11612;
  assign n11616 = n10997 & ~n33242;
  assign n11617 = n11001 & n11613;
  assign n11618 = n10997 & ~n33163;
  assign n11619 = ~n10989 & n11618;
  assign n11620 = ~n11097 & n11619;
  assign n11621 = ~n10997 & ~n33242;
  assign n11622 = ~n11620 & ~n11621;
  assign n11623 = ~n11616 & ~n11617;
  assign n11624 = ~n11611 & ~n33243;
  assign n11625 = ~n11609 & ~n11624;
  assign n11626 = ~n321 & ~n11625;
  assign n11627 = n321 & ~n11609;
  assign n11628 = ~n11624 & n11627;
  assign n11629 = n321 & n11625;
  assign n11630 = ~n11003 & ~n11013;
  assign n11631 = ~n11003 & ~n11097;
  assign n11632 = ~n11013 & n11631;
  assign n11633 = ~n11097 & n11630;
  assign n11634 = n11011 & ~n33245;
  assign n11635 = n11014 & n11631;
  assign n11636 = ~n11003 & n11011;
  assign n11637 = ~n11013 & n11636;
  assign n11638 = ~n11097 & n11637;
  assign n11639 = ~n11011 & ~n33245;
  assign n11640 = ~n11638 & ~n11639;
  assign n11641 = ~n11634 & ~n11635;
  assign n11642 = ~n33244 & ~n33246;
  assign n11643 = ~n11626 & ~n11642;
  assign n11644 = ~n263 & ~n11643;
  assign n11645 = n263 & ~n11626;
  assign n11646 = ~n11642 & n11645;
  assign n11647 = ~n11016 & ~n33166;
  assign n11648 = ~n11016 & ~n11097;
  assign n11649 = ~n33166 & n11648;
  assign n11650 = ~n11097 & n11647;
  assign n11651 = n11024 & ~n33247;
  assign n11652 = n11028 & n11648;
  assign n11653 = n11024 & ~n33166;
  assign n11654 = ~n11016 & n11653;
  assign n11655 = ~n11097 & n11654;
  assign n11656 = ~n11024 & ~n33247;
  assign n11657 = ~n11655 & ~n11656;
  assign n11658 = ~n11651 & ~n11652;
  assign n11659 = ~n11646 & ~n33248;
  assign n11660 = ~n11644 & ~n11659;
  assign n11661 = ~n214 & ~n11660;
  assign n11662 = ~n11030 & ~n11032;
  assign n11663 = ~n11097 & n11662;
  assign n11664 = ~n33168 & ~n11663;
  assign n11665 = ~n11030 & n33168;
  assign n11666 = ~n11032 & n11665;
  assign n11667 = n33168 & n11663;
  assign n11668 = ~n11097 & n11666;
  assign n11669 = ~n11664 & ~n33249;
  assign n11670 = n214 & ~n11644;
  assign n11671 = ~n11659 & n11670;
  assign n11672 = n214 & n11660;
  assign n11673 = ~n11669 & ~n33250;
  assign n11674 = ~n11661 & ~n11673;
  assign n11675 = ~n197 & ~n11674;
  assign n11676 = n197 & ~n11661;
  assign n11677 = ~n11673 & n11676;
  assign n11678 = ~n11047 & ~n33170;
  assign n11679 = ~n11047 & ~n11097;
  assign n11680 = ~n33170 & n11679;
  assign n11681 = ~n11097 & n11678;
  assign n11682 = n11055 & ~n33251;
  assign n11683 = n11059 & n11679;
  assign n11684 = n11055 & ~n33170;
  assign n11685 = ~n11047 & n11684;
  assign n11686 = ~n11097 & n11685;
  assign n11687 = ~n11055 & ~n33251;
  assign n11688 = ~n11686 & ~n11687;
  assign n11689 = ~n11682 & ~n11683;
  assign n11690 = ~n11677 & ~n33252;
  assign n11691 = ~n11675 & ~n11690;
  assign n11692 = ~n11061 & ~n11071;
  assign n11693 = ~n11061 & ~n11097;
  assign n11694 = ~n11071 & n11693;
  assign n11695 = ~n11097 & n11692;
  assign n11696 = n11069 & ~n33253;
  assign n11697 = n11072 & n11693;
  assign n11698 = ~n11061 & n11069;
  assign n11699 = ~n11071 & n11698;
  assign n11700 = ~n11097 & n11699;
  assign n11701 = ~n11069 & ~n33253;
  assign n11702 = ~n11700 & ~n11701;
  assign n11703 = ~n11696 & ~n11697;
  assign n11704 = ~n11073 & ~n11081;
  assign n11705 = ~n11081 & ~n11097;
  assign n11706 = ~n11073 & n11705;
  assign n11707 = ~n11097 & n11704;
  assign n11708 = ~n33174 & ~n33255;
  assign n11709 = ~n33254 & n11708;
  assign n11710 = ~n11691 & n11709;
  assign n11711 = n193 & ~n11710;
  assign n11712 = ~n11675 & n33254;
  assign n11713 = ~n11690 & n11712;
  assign n11714 = n11691 & n33254;
  assign n11715 = n11073 & ~n11705;
  assign n11716 = ~n193 & ~n11704;
  assign n11717 = ~n11715 & n11716;
  assign n11718 = ~n33256 & ~n11717;
  assign n11719 = ~n11711 & n11718;
  assign n11720 = ~n11216 & ~n11218;
  assign n11721 = ~n11719 & n11720;
  assign n11722 = ~n33191 & ~n11721;
  assign n11723 = ~n11218 & n33191;
  assign n11724 = ~n11216 & n11723;
  assign n11725 = n33191 & n11721;
  assign n11726 = ~n11719 & n11724;
  assign n11727 = ~n11722 & ~n33257;
  assign n11728 = ~n11183 & ~n11185;
  assign n11729 = ~n11719 & n11728;
  assign n11730 = ~n33187 & ~n11729;
  assign n11731 = ~n11185 & n33187;
  assign n11732 = ~n11183 & n11731;
  assign n11733 = n33187 & n11729;
  assign n11734 = ~n11719 & n11732;
  assign n11735 = ~n11730 & ~n33258;
  assign n11736 = ~n11149 & ~n11151;
  assign n11737 = ~n11719 & n11736;
  assign n11738 = ~n33182 & ~n11737;
  assign n11739 = ~n11151 & n33182;
  assign n11740 = ~n11149 & n11739;
  assign n11741 = n33182 & n11737;
  assign n11742 = ~n11719 & n11740;
  assign n11743 = ~n11738 & ~n33259;
  assign n11744 = ~n11122 & ~n11124;
  assign n11745 = ~n11719 & n11744;
  assign n11746 = ~n11133 & ~n11745;
  assign n11747 = ~n11124 & n11133;
  assign n11748 = ~n11122 & n11747;
  assign n11749 = n11133 & n11745;
  assign n11750 = ~n11719 & n11748;
  assign n11751 = ~n11746 & ~n33260;
  assign n11752 = ~pi50  & ~n11719;
  assign n11753 = ~pi51  & n11752;
  assign n11754 = n11099 & ~n11719;
  assign n11755 = ~n11097 & ~n11717;
  assign n11756 = ~n33256 & n11755;
  assign n11757 = ~n11711 & n11756;
  assign n11758 = ~n33261 & ~n11757;
  assign n11759 = pi52  & ~n11758;
  assign n11760 = ~pi52  & ~n11757;
  assign n11761 = ~pi52  & n11758;
  assign n11762 = ~n33261 & n11760;
  assign n11763 = ~n11759 & ~n33262;
  assign n11764 = pi50  & ~n11719;
  assign n11765 = ~pi48  & ~pi49 ;
  assign n11766 = ~pi50  & n11765;
  assign n11767 = ~n33106 & ~n33176;
  assign n11768 = ~n10534 & n11767;
  assign n11769 = ~n10553 & n11768;
  assign n11770 = ~n33108 & n11769;
  assign n11771 = n10539 & n10555;
  assign n11772 = ~n10547 & n11770;
  assign n11773 = ~n11766 & ~n33263;
  assign n11774 = ~n11095 & n11773;
  assign n11775 = ~n33174 & n11774;
  assign n11776 = ~n11089 & n11775;
  assign n11777 = ~n11764 & ~n11766;
  assign n11778 = n11097 & n11777;
  assign n11779 = ~n11764 & n11776;
  assign n11780 = pi51  & ~n11752;
  assign n11781 = ~n33261 & ~n11780;
  assign n11782 = ~n33264 & n11781;
  assign n11783 = ~n11097 & ~n11777;
  assign n11784 = n10555 & ~n11783;
  assign n11785 = ~n11782 & ~n11783;
  assign n11786 = n10555 & n11785;
  assign n11787 = ~n11782 & n11784;
  assign n11788 = ~n11763 & ~n33265;
  assign n11789 = ~n10555 & ~n11785;
  assign n11790 = n9969 & ~n11789;
  assign n11791 = ~n11788 & n11790;
  assign n11792 = ~n11102 & ~n33177;
  assign n11793 = ~n11719 & n11792;
  assign n11794 = n11107 & ~n11793;
  assign n11795 = ~n11107 & n11792;
  assign n11796 = ~n11107 & n11793;
  assign n11797 = ~n11719 & n11795;
  assign n11798 = ~n11794 & ~n33266;
  assign n11799 = ~n11791 & ~n11798;
  assign n11800 = ~n11788 & ~n11789;
  assign n11801 = ~n9969 & ~n11800;
  assign n11802 = n9457 & ~n11801;
  assign n11803 = ~n11799 & ~n11801;
  assign n11804 = n9457 & n11803;
  assign n11805 = ~n11799 & n11802;
  assign n11806 = ~n11751 & ~n33267;
  assign n11807 = ~n9457 & ~n11803;
  assign n11808 = n8896 & ~n11807;
  assign n11809 = ~n11806 & n11808;
  assign n11810 = ~n11136 & ~n33179;
  assign n11811 = ~n11719 & n11810;
  assign n11812 = ~n11146 & ~n11811;
  assign n11813 = ~n11136 & n11146;
  assign n11814 = ~n33179 & n11813;
  assign n11815 = n11146 & n11811;
  assign n11816 = ~n11719 & n11814;
  assign n11817 = n11146 & ~n11811;
  assign n11818 = ~n11146 & n11811;
  assign n11819 = ~n11817 & ~n11818;
  assign n11820 = ~n11812 & ~n33268;
  assign n11821 = ~n11809 & n33269;
  assign n11822 = ~n11806 & ~n11807;
  assign n11823 = ~n8896 & ~n11822;
  assign n11824 = n8411 & ~n11823;
  assign n11825 = ~n11821 & ~n11823;
  assign n11826 = n8411 & n11825;
  assign n11827 = ~n11821 & n11824;
  assign n11828 = ~n11743 & ~n33270;
  assign n11829 = ~n8411 & ~n11825;
  assign n11830 = n7885 & ~n11829;
  assign n11831 = ~n11828 & n11830;
  assign n11832 = ~n11166 & ~n33183;
  assign n11833 = ~n11719 & n11832;
  assign n11834 = ~n33185 & ~n11833;
  assign n11835 = n33185 & n11833;
  assign n11836 = ~n11166 & ~n33185;
  assign n11837 = ~n33183 & n11836;
  assign n11838 = ~n11719 & n11837;
  assign n11839 = n33185 & ~n11833;
  assign n11840 = ~n11838 & ~n11839;
  assign n11841 = ~n11834 & ~n11835;
  assign n11842 = ~n11831 & ~n33271;
  assign n11843 = ~n11828 & ~n11829;
  assign n11844 = ~n7885 & ~n11843;
  assign n11845 = n7428 & ~n11844;
  assign n11846 = ~n11842 & ~n11844;
  assign n11847 = n7428 & n11846;
  assign n11848 = ~n11842 & n11845;
  assign n11849 = ~n11735 & ~n33272;
  assign n11850 = ~n7428 & ~n11846;
  assign n11851 = n6937 & ~n11850;
  assign n11852 = ~n11849 & n11851;
  assign n11853 = ~n11200 & ~n33188;
  assign n11854 = ~n11719 & n11853;
  assign n11855 = ~n33189 & n11854;
  assign n11856 = n33189 & ~n11854;
  assign n11857 = ~n11200 & n33189;
  assign n11858 = ~n33188 & n11857;
  assign n11859 = ~n11719 & n11858;
  assign n11860 = ~n33189 & ~n11854;
  assign n11861 = ~n11859 & ~n11860;
  assign n11862 = ~n11855 & ~n11856;
  assign n11863 = ~n11852 & ~n33273;
  assign n11864 = ~n11849 & ~n11850;
  assign n11865 = ~n6937 & ~n11864;
  assign n11866 = n6507 & ~n11865;
  assign n11867 = ~n11863 & ~n11865;
  assign n11868 = n6507 & n11867;
  assign n11869 = ~n11863 & n11866;
  assign n11870 = ~n11727 & ~n33274;
  assign n11871 = ~n6507 & ~n11867;
  assign n11872 = n6051 & ~n11871;
  assign n11873 = ~n11870 & n11872;
  assign n11874 = ~n11233 & ~n33192;
  assign n11875 = ~n11719 & n11874;
  assign n11876 = ~n33193 & n11875;
  assign n11877 = n33193 & ~n11875;
  assign n11878 = ~n33193 & ~n11875;
  assign n11879 = ~n11233 & n33193;
  assign n11880 = ~n33192 & n11879;
  assign n11881 = n33193 & n11875;
  assign n11882 = ~n11719 & n11880;
  assign n11883 = ~n11878 & ~n33275;
  assign n11884 = ~n11876 & ~n11877;
  assign n11885 = ~n11873 & ~n33276;
  assign n11886 = ~n11870 & ~n11871;
  assign n11887 = ~n6051 & ~n11886;
  assign n11888 = n5648 & ~n11887;
  assign n11889 = ~n11885 & ~n11887;
  assign n11890 = n5648 & n11889;
  assign n11891 = ~n11885 & n11888;
  assign n11892 = ~n11249 & ~n11251;
  assign n11893 = ~n11719 & n11892;
  assign n11894 = ~n33194 & n11893;
  assign n11895 = n33194 & ~n11893;
  assign n11896 = ~n11251 & n33194;
  assign n11897 = ~n11249 & n11896;
  assign n11898 = ~n11719 & n11897;
  assign n11899 = ~n33194 & ~n11893;
  assign n11900 = ~n11898 & ~n11899;
  assign n11901 = ~n11894 & ~n11895;
  assign n11902 = ~n33277 & ~n33278;
  assign n11903 = ~n5648 & ~n11889;
  assign n11904 = ~n11902 & ~n11903;
  assign n11905 = ~n5223 & ~n11904;
  assign n11906 = ~n11264 & ~n33196;
  assign n11907 = ~n11719 & n11906;
  assign n11908 = n33195 & ~n11907;
  assign n11909 = ~n33195 & n11907;
  assign n11910 = ~n11264 & n33195;
  assign n11911 = ~n33196 & n11910;
  assign n11912 = ~n11719 & n11911;
  assign n11913 = ~n33195 & ~n11907;
  assign n11914 = ~n11912 & ~n11913;
  assign n11915 = ~n11908 & ~n11909;
  assign n11916 = n5223 & ~n11903;
  assign n11917 = ~n11902 & n11916;
  assign n11918 = ~n33279 & ~n11917;
  assign n11919 = ~n11905 & ~n11918;
  assign n11920 = ~n4851 & ~n11919;
  assign n11921 = ~n11280 & ~n11282;
  assign n11922 = ~n11719 & n11921;
  assign n11923 = ~n33198 & ~n11922;
  assign n11924 = ~n11282 & n33198;
  assign n11925 = ~n11280 & n11924;
  assign n11926 = n33198 & n11922;
  assign n11927 = ~n11719 & n11925;
  assign n11928 = ~n11923 & ~n33280;
  assign n11929 = n4851 & ~n11905;
  assign n11930 = n4851 & n11919;
  assign n11931 = ~n11918 & n11929;
  assign n11932 = ~n11928 & ~n33281;
  assign n11933 = ~n11920 & ~n11932;
  assign n11934 = ~n4461 & ~n11933;
  assign n11935 = n4461 & ~n11920;
  assign n11936 = ~n11932 & n11935;
  assign n11937 = ~n11297 & ~n33199;
  assign n11938 = ~n11297 & ~n11719;
  assign n11939 = ~n33199 & n11938;
  assign n11940 = ~n11719 & n11937;
  assign n11941 = ~n33201 & ~n33282;
  assign n11942 = ~n11297 & n33201;
  assign n11943 = ~n33199 & n11942;
  assign n11944 = n33201 & n33282;
  assign n11945 = ~n11719 & n11943;
  assign n11946 = n33201 & ~n33282;
  assign n11947 = n11312 & n11938;
  assign n11948 = ~n11946 & ~n11947;
  assign n11949 = ~n11941 & ~n33283;
  assign n11950 = ~n11936 & n33284;
  assign n11951 = ~n11934 & ~n11950;
  assign n11952 = ~n4115 & ~n11951;
  assign n11953 = ~n11314 & ~n11316;
  assign n11954 = ~n11719 & n11953;
  assign n11955 = ~n33203 & ~n11954;
  assign n11956 = ~n11316 & n33203;
  assign n11957 = ~n11314 & n11956;
  assign n11958 = n33203 & n11954;
  assign n11959 = ~n11719 & n11957;
  assign n11960 = ~n11955 & ~n33285;
  assign n11961 = n4115 & ~n11934;
  assign n11962 = n4115 & n11951;
  assign n11963 = ~n11950 & n11961;
  assign n11964 = ~n11960 & ~n33286;
  assign n11965 = ~n11952 & ~n11964;
  assign n11966 = ~n3754 & ~n11965;
  assign n11967 = n3754 & ~n11952;
  assign n11968 = ~n11964 & n11967;
  assign n11969 = ~n11331 & ~n33205;
  assign n11970 = ~n11331 & ~n11719;
  assign n11971 = ~n33205 & n11970;
  assign n11972 = ~n11719 & n11969;
  assign n11973 = n11339 & ~n33287;
  assign n11974 = n11343 & n11970;
  assign n11975 = ~n11331 & n11339;
  assign n11976 = ~n33205 & n11975;
  assign n11977 = ~n11719 & n11976;
  assign n11978 = ~n11339 & ~n33287;
  assign n11979 = ~n11977 & ~n11978;
  assign n11980 = ~n11973 & ~n11974;
  assign n11981 = ~n11968 & ~n33288;
  assign n11982 = ~n11966 & ~n11981;
  assign n11983 = ~n3444 & ~n11982;
  assign n11984 = ~n11345 & ~n11347;
  assign n11985 = ~n11719 & n11984;
  assign n11986 = ~n33207 & ~n11985;
  assign n11987 = ~n11347 & n33207;
  assign n11988 = ~n11345 & n11987;
  assign n11989 = n33207 & n11985;
  assign n11990 = ~n11719 & n11988;
  assign n11991 = ~n11986 & ~n33289;
  assign n11992 = n3444 & ~n11966;
  assign n11993 = n3444 & n11982;
  assign n11994 = ~n11981 & n11992;
  assign n11995 = ~n11991 & ~n33290;
  assign n11996 = ~n11983 & ~n11995;
  assign n11997 = ~n3116 & ~n11996;
  assign n11998 = ~n11362 & ~n33208;
  assign n11999 = ~n11719 & n11998;
  assign n12000 = ~n33210 & ~n11999;
  assign n12001 = ~n11362 & n33210;
  assign n12002 = ~n33208 & n12001;
  assign n12003 = n33210 & n11999;
  assign n12004 = ~n11719 & n12002;
  assign n12005 = ~n12000 & ~n33291;
  assign n12006 = n3116 & ~n11983;
  assign n12007 = ~n11995 & n12006;
  assign n12008 = ~n12005 & ~n12007;
  assign n12009 = ~n11997 & ~n12008;
  assign n12010 = ~n2833 & ~n12009;
  assign n12011 = ~n11380 & ~n11382;
  assign n12012 = ~n11719 & n12011;
  assign n12013 = ~n33212 & ~n12012;
  assign n12014 = ~n11382 & n33212;
  assign n12015 = ~n11380 & n12014;
  assign n12016 = n33212 & n12012;
  assign n12017 = ~n11719 & n12015;
  assign n12018 = ~n12013 & ~n33292;
  assign n12019 = n2833 & ~n11997;
  assign n12020 = n2833 & n12009;
  assign n12021 = ~n12008 & n12019;
  assign n12022 = ~n12018 & ~n33293;
  assign n12023 = ~n12010 & ~n12022;
  assign n12024 = ~n2536 & ~n12023;
  assign n12025 = n2536 & ~n12010;
  assign n12026 = ~n12022 & n12025;
  assign n12027 = ~n11397 & ~n33214;
  assign n12028 = ~n11397 & ~n11719;
  assign n12029 = ~n33214 & n12028;
  assign n12030 = ~n11719 & n12027;
  assign n12031 = n11405 & ~n33294;
  assign n12032 = n11409 & n12028;
  assign n12033 = ~n11397 & n11405;
  assign n12034 = ~n33214 & n12033;
  assign n12035 = ~n11719 & n12034;
  assign n12036 = ~n11405 & ~n33294;
  assign n12037 = ~n12035 & ~n12036;
  assign n12038 = ~n12031 & ~n12032;
  assign n12039 = ~n12026 & ~n33295;
  assign n12040 = ~n12024 & ~n12039;
  assign n12041 = ~n2283 & ~n12040;
  assign n12042 = ~n11411 & ~n11413;
  assign n12043 = ~n11719 & n12042;
  assign n12044 = ~n33216 & ~n12043;
  assign n12045 = ~n11413 & n33216;
  assign n12046 = ~n11411 & n12045;
  assign n12047 = n33216 & n12043;
  assign n12048 = ~n11719 & n12046;
  assign n12049 = ~n12044 & ~n33296;
  assign n12050 = n2283 & ~n12024;
  assign n12051 = n2283 & n12040;
  assign n12052 = ~n12039 & n12050;
  assign n12053 = ~n12049 & ~n33297;
  assign n12054 = ~n12041 & ~n12053;
  assign n12055 = ~n2021 & ~n12054;
  assign n12056 = ~n11428 & ~n33217;
  assign n12057 = ~n11719 & n12056;
  assign n12058 = ~n33219 & ~n12057;
  assign n12059 = ~n11428 & n33219;
  assign n12060 = ~n33217 & n12059;
  assign n12061 = n33219 & n12057;
  assign n12062 = ~n11719 & n12060;
  assign n12063 = ~n12058 & ~n33298;
  assign n12064 = n2021 & ~n12041;
  assign n12065 = ~n12053 & n12064;
  assign n12066 = ~n12063 & ~n12065;
  assign n12067 = ~n12055 & ~n12066;
  assign n12068 = ~n1796 & ~n12067;
  assign n12069 = ~n11446 & ~n11448;
  assign n12070 = ~n11719 & n12069;
  assign n12071 = ~n33221 & ~n12070;
  assign n12072 = ~n11448 & n33221;
  assign n12073 = ~n11446 & n12072;
  assign n12074 = n33221 & n12070;
  assign n12075 = ~n11719 & n12073;
  assign n12076 = ~n12071 & ~n33299;
  assign n12077 = n1796 & ~n12055;
  assign n12078 = n1796 & n12067;
  assign n12079 = ~n12066 & n12077;
  assign n12080 = ~n12076 & ~n33300;
  assign n12081 = ~n12068 & ~n12080;
  assign n12082 = ~n1567 & ~n12081;
  assign n12083 = n1567 & ~n12068;
  assign n12084 = ~n12080 & n12083;
  assign n12085 = ~n11463 & ~n33223;
  assign n12086 = ~n11463 & ~n11719;
  assign n12087 = ~n33223 & n12086;
  assign n12088 = ~n11719 & n12085;
  assign n12089 = n11471 & ~n33301;
  assign n12090 = n11475 & n12086;
  assign n12091 = ~n11463 & n11471;
  assign n12092 = ~n33223 & n12091;
  assign n12093 = ~n11719 & n12092;
  assign n12094 = ~n11471 & ~n33301;
  assign n12095 = ~n12093 & ~n12094;
  assign n12096 = ~n12089 & ~n12090;
  assign n12097 = ~n12084 & ~n33302;
  assign n12098 = ~n12082 & ~n12097;
  assign n12099 = ~n1374 & ~n12098;
  assign n12100 = ~n11477 & ~n11479;
  assign n12101 = ~n11719 & n12100;
  assign n12102 = ~n33225 & ~n12101;
  assign n12103 = ~n11479 & n33225;
  assign n12104 = ~n11477 & n12103;
  assign n12105 = n33225 & n12101;
  assign n12106 = ~n11719 & n12104;
  assign n12107 = ~n12102 & ~n33303;
  assign n12108 = n1374 & ~n12082;
  assign n12109 = n1374 & n12098;
  assign n12110 = ~n12097 & n12108;
  assign n12111 = ~n12107 & ~n33304;
  assign n12112 = ~n12099 & ~n12111;
  assign n12113 = ~n1179 & ~n12112;
  assign n12114 = ~n11494 & ~n33226;
  assign n12115 = ~n11719 & n12114;
  assign n12116 = ~n33228 & ~n12115;
  assign n12117 = ~n11494 & n33228;
  assign n12118 = ~n33226 & n12117;
  assign n12119 = n33228 & n12115;
  assign n12120 = ~n11719 & n12118;
  assign n12121 = ~n12116 & ~n33305;
  assign n12122 = n1179 & ~n12099;
  assign n12123 = ~n12111 & n12122;
  assign n12124 = ~n12121 & ~n12123;
  assign n12125 = ~n12113 & ~n12124;
  assign n12126 = ~n1016 & ~n12125;
  assign n12127 = ~n11512 & ~n11514;
  assign n12128 = ~n11719 & n12127;
  assign n12129 = ~n33230 & ~n12128;
  assign n12130 = ~n11514 & n33230;
  assign n12131 = ~n11512 & n12130;
  assign n12132 = n33230 & n12128;
  assign n12133 = ~n11719 & n12131;
  assign n12134 = ~n12129 & ~n33306;
  assign n12135 = n1016 & ~n12113;
  assign n12136 = n1016 & n12125;
  assign n12137 = ~n12124 & n12135;
  assign n12138 = ~n12134 & ~n33307;
  assign n12139 = ~n12126 & ~n12138;
  assign n12140 = ~n855 & ~n12139;
  assign n12141 = n855 & ~n12126;
  assign n12142 = ~n12138 & n12141;
  assign n12143 = ~n11529 & ~n33232;
  assign n12144 = ~n11529 & ~n11719;
  assign n12145 = ~n33232 & n12144;
  assign n12146 = ~n11719 & n12143;
  assign n12147 = n11537 & ~n33308;
  assign n12148 = n11541 & n12144;
  assign n12149 = ~n11529 & n11537;
  assign n12150 = ~n33232 & n12149;
  assign n12151 = ~n11719 & n12150;
  assign n12152 = ~n11537 & ~n33308;
  assign n12153 = ~n12151 & ~n12152;
  assign n12154 = ~n12147 & ~n12148;
  assign n12155 = ~n12142 & ~n33309;
  assign n12156 = ~n12140 & ~n12155;
  assign n12157 = ~n720 & ~n12156;
  assign n12158 = ~n11543 & ~n11545;
  assign n12159 = ~n11719 & n12158;
  assign n12160 = ~n33234 & ~n12159;
  assign n12161 = ~n11545 & n33234;
  assign n12162 = ~n11543 & n12161;
  assign n12163 = n33234 & n12159;
  assign n12164 = ~n11719 & n12162;
  assign n12165 = ~n12160 & ~n33310;
  assign n12166 = n720 & ~n12140;
  assign n12167 = n720 & n12156;
  assign n12168 = ~n12155 & n12166;
  assign n12169 = ~n12165 & ~n33311;
  assign n12170 = ~n12157 & ~n12169;
  assign n12171 = ~n592 & ~n12170;
  assign n12172 = ~n11560 & ~n33235;
  assign n12173 = ~n11719 & n12172;
  assign n12174 = ~n33237 & ~n12173;
  assign n12175 = ~n11560 & n33237;
  assign n12176 = ~n33235 & n12175;
  assign n12177 = n33237 & n12173;
  assign n12178 = ~n11719 & n12176;
  assign n12179 = ~n12174 & ~n33312;
  assign n12180 = n592 & ~n12157;
  assign n12181 = ~n12169 & n12180;
  assign n12182 = ~n12179 & ~n12181;
  assign n12183 = ~n12171 & ~n12182;
  assign n12184 = ~n487 & ~n12183;
  assign n12185 = ~n11578 & ~n11580;
  assign n12186 = ~n11719 & n12185;
  assign n12187 = ~n33239 & ~n12186;
  assign n12188 = ~n11580 & n33239;
  assign n12189 = ~n11578 & n12188;
  assign n12190 = n33239 & n12186;
  assign n12191 = ~n11719 & n12189;
  assign n12192 = ~n12187 & ~n33313;
  assign n12193 = n487 & ~n12171;
  assign n12194 = n487 & n12183;
  assign n12195 = ~n12182 & n12193;
  assign n12196 = ~n12192 & ~n33314;
  assign n12197 = ~n12184 & ~n12196;
  assign n12198 = ~n393 & ~n12197;
  assign n12199 = n393 & ~n12184;
  assign n12200 = ~n12196 & n12199;
  assign n12201 = ~n11595 & ~n33241;
  assign n12202 = ~n11595 & ~n11719;
  assign n12203 = ~n33241 & n12202;
  assign n12204 = ~n11719 & n12201;
  assign n12205 = n11603 & ~n33315;
  assign n12206 = n11607 & n12202;
  assign n12207 = ~n11595 & n11603;
  assign n12208 = ~n33241 & n12207;
  assign n12209 = ~n11719 & n12208;
  assign n12210 = ~n11603 & ~n33315;
  assign n12211 = ~n12209 & ~n12210;
  assign n12212 = ~n12205 & ~n12206;
  assign n12213 = ~n12200 & ~n33316;
  assign n12214 = ~n12198 & ~n12213;
  assign n12215 = ~n321 & ~n12214;
  assign n12216 = ~n11609 & ~n11611;
  assign n12217 = ~n11719 & n12216;
  assign n12218 = ~n33243 & ~n12217;
  assign n12219 = ~n11611 & n33243;
  assign n12220 = ~n11609 & n12219;
  assign n12221 = n33243 & n12217;
  assign n12222 = ~n11719 & n12220;
  assign n12223 = ~n12218 & ~n33317;
  assign n12224 = n321 & ~n12198;
  assign n12225 = n321 & n12214;
  assign n12226 = ~n12213 & n12224;
  assign n12227 = ~n12223 & ~n33318;
  assign n12228 = ~n12215 & ~n12227;
  assign n12229 = ~n263 & ~n12228;
  assign n12230 = ~n11626 & ~n33244;
  assign n12231 = ~n11719 & n12230;
  assign n12232 = ~n33246 & ~n12231;
  assign n12233 = ~n11626 & n33246;
  assign n12234 = ~n33244 & n12233;
  assign n12235 = n33246 & n12231;
  assign n12236 = ~n11719 & n12234;
  assign n12237 = ~n12232 & ~n33319;
  assign n12238 = n263 & ~n12215;
  assign n12239 = ~n12227 & n12238;
  assign n12240 = ~n12237 & ~n12239;
  assign n12241 = ~n12229 & ~n12240;
  assign n12242 = ~n214 & ~n12241;
  assign n12243 = ~n11644 & ~n11646;
  assign n12244 = ~n11719 & n12243;
  assign n12245 = ~n33248 & ~n12244;
  assign n12246 = ~n11646 & n33248;
  assign n12247 = ~n11644 & n12246;
  assign n12248 = n33248 & n12244;
  assign n12249 = ~n11719 & n12247;
  assign n12250 = ~n12245 & ~n33320;
  assign n12251 = n214 & ~n12229;
  assign n12252 = n214 & n12241;
  assign n12253 = ~n12240 & n12251;
  assign n12254 = ~n12250 & ~n33321;
  assign n12255 = ~n12242 & ~n12254;
  assign n12256 = ~n197 & ~n12255;
  assign n12257 = n197 & ~n12242;
  assign n12258 = ~n12254 & n12257;
  assign n12259 = ~n11661 & ~n33250;
  assign n12260 = ~n11661 & ~n11719;
  assign n12261 = ~n33250 & n12260;
  assign n12262 = ~n11719 & n12259;
  assign n12263 = n11669 & ~n33322;
  assign n12264 = n11673 & n12260;
  assign n12265 = ~n11661 & n11669;
  assign n12266 = ~n33250 & n12265;
  assign n12267 = ~n11719 & n12266;
  assign n12268 = ~n11669 & ~n33322;
  assign n12269 = ~n12267 & ~n12268;
  assign n12270 = ~n12263 & ~n12264;
  assign n12271 = ~n12258 & ~n33323;
  assign n12272 = ~n12256 & ~n12271;
  assign n12273 = ~n11675 & ~n11677;
  assign n12274 = ~n11719 & n12273;
  assign n12275 = ~n33252 & ~n12274;
  assign n12276 = ~n11677 & n33252;
  assign n12277 = ~n11675 & n12276;
  assign n12278 = n33252 & n12274;
  assign n12279 = ~n11719 & n12277;
  assign n12280 = ~n12275 & ~n33324;
  assign n12281 = ~n11691 & ~n33254;
  assign n12282 = ~n33254 & ~n11719;
  assign n12283 = ~n11691 & n12282;
  assign n12284 = ~n11719 & n12281;
  assign n12285 = ~n33256 & ~n33325;
  assign n12286 = ~n12280 & n12285;
  assign n12287 = ~n12272 & n12286;
  assign n12288 = n193 & ~n12287;
  assign n12289 = ~n12256 & n12280;
  assign n12290 = n12272 & n12280;
  assign n12291 = ~n12271 & n12289;
  assign n12292 = n11691 & ~n12282;
  assign n12293 = ~n193 & ~n12281;
  assign n12294 = ~n12292 & n12293;
  assign n12295 = ~n33326 & ~n12294;
  assign n12296 = ~n12288 & n12295;
  assign n12297 = pi48  & ~n12296;
  assign n12298 = ~pi46  & ~pi47 ;
  assign n12299 = ~pi48  & n12298;
  assign n12300 = ~n12297 & ~n12299;
  assign n12301 = ~n11719 & ~n12300;
  assign n12302 = ~pi48  & ~n12296;
  assign n12303 = pi49  & ~n12302;
  assign n12304 = ~pi49  & n12302;
  assign n12305 = n11765 & ~n12296;
  assign n12306 = ~n12303 & ~n33327;
  assign n12307 = ~n33172 & ~n33263;
  assign n12308 = ~n11076 & n12307;
  assign n12309 = ~n11095 & n12308;
  assign n12310 = ~n33174 & n12309;
  assign n12311 = n11081 & n11097;
  assign n12312 = ~n11089 & n12310;
  assign n12313 = ~n12299 & ~n33328;
  assign n12314 = ~n11717 & n12313;
  assign n12315 = ~n33256 & n12314;
  assign n12316 = ~n11711 & n12315;
  assign n12317 = n11719 & n12300;
  assign n12318 = ~n12297 & n12316;
  assign n12319 = n12306 & ~n33329;
  assign n12320 = ~n12301 & ~n12319;
  assign n12321 = ~n11097 & ~n12320;
  assign n12322 = n11097 & ~n12301;
  assign n12323 = ~n12319 & n12322;
  assign n12324 = ~n11719 & ~n12294;
  assign n12325 = ~n33326 & n12324;
  assign n12326 = ~n12288 & n12325;
  assign n12327 = ~n33327 & ~n12326;
  assign n12328 = pi50  & ~n12327;
  assign n12329 = ~pi50  & ~n12326;
  assign n12330 = ~pi50  & n12327;
  assign n12331 = ~n33327 & n12329;
  assign n12332 = ~n12328 & ~n33330;
  assign n12333 = ~n12323 & ~n12332;
  assign n12334 = ~n12321 & ~n12333;
  assign n12335 = ~n10555 & ~n12334;
  assign n12336 = n10555 & ~n12321;
  assign n12337 = ~n12333 & n12336;
  assign n12338 = n10555 & n12334;
  assign n12339 = ~n33264 & ~n11783;
  assign n12340 = ~n12296 & n12339;
  assign n12341 = n11781 & ~n12340;
  assign n12342 = ~n11781 & n12339;
  assign n12343 = ~n11781 & n12340;
  assign n12344 = ~n12296 & n12342;
  assign n12345 = ~n12341 & ~n33332;
  assign n12346 = ~n33331 & ~n12345;
  assign n12347 = ~n12335 & ~n12346;
  assign n12348 = ~n9969 & ~n12347;
  assign n12349 = n9969 & ~n12335;
  assign n12350 = ~n12346 & n12349;
  assign n12351 = ~n33265 & ~n11789;
  assign n12352 = ~n11789 & ~n12296;
  assign n12353 = ~n33265 & n12352;
  assign n12354 = ~n12296 & n12351;
  assign n12355 = n11763 & ~n33333;
  assign n12356 = n11788 & n12352;
  assign n12357 = n11763 & ~n33265;
  assign n12358 = ~n11789 & n12357;
  assign n12359 = ~n12296 & n12358;
  assign n12360 = ~n11763 & ~n33333;
  assign n12361 = ~n12359 & ~n12360;
  assign n12362 = ~n12355 & ~n12356;
  assign n12363 = ~n12350 & ~n33334;
  assign n12364 = ~n12348 & ~n12363;
  assign n12365 = ~n9457 & ~n12364;
  assign n12366 = n9457 & ~n12348;
  assign n12367 = ~n12363 & n12366;
  assign n12368 = n9457 & n12364;
  assign n12369 = ~n11791 & ~n11801;
  assign n12370 = ~n12296 & n12369;
  assign n12371 = ~n11798 & ~n12370;
  assign n12372 = n11798 & ~n11801;
  assign n12373 = ~n11791 & n12372;
  assign n12374 = n11798 & n12370;
  assign n12375 = ~n12296 & n12373;
  assign n12376 = n11798 & ~n12370;
  assign n12377 = ~n11798 & n12370;
  assign n12378 = ~n12376 & ~n12377;
  assign n12379 = ~n12371 & ~n33336;
  assign n12380 = ~n33335 & n33337;
  assign n12381 = ~n12365 & ~n12380;
  assign n12382 = ~n8896 & ~n12381;
  assign n12383 = n8896 & ~n12365;
  assign n12384 = ~n12380 & n12383;
  assign n12385 = ~n33267 & ~n11807;
  assign n12386 = ~n11807 & ~n12296;
  assign n12387 = ~n33267 & n12386;
  assign n12388 = ~n12296 & n12385;
  assign n12389 = n11751 & ~n33338;
  assign n12390 = n11806 & n12386;
  assign n12391 = n11751 & ~n33267;
  assign n12392 = ~n11807 & n12391;
  assign n12393 = ~n12296 & n12392;
  assign n12394 = ~n11751 & ~n33338;
  assign n12395 = ~n12393 & ~n12394;
  assign n12396 = ~n12389 & ~n12390;
  assign n12397 = ~n12384 & ~n33339;
  assign n12398 = ~n12382 & ~n12397;
  assign n12399 = ~n8411 & ~n12398;
  assign n12400 = n8411 & ~n12382;
  assign n12401 = ~n12397 & n12400;
  assign n12402 = n8411 & n12398;
  assign n12403 = ~n11809 & ~n11823;
  assign n12404 = ~n12296 & n12403;
  assign n12405 = ~n33269 & ~n12404;
  assign n12406 = n33269 & n12404;
  assign n12407 = ~n33269 & ~n11823;
  assign n12408 = ~n11809 & n12407;
  assign n12409 = ~n12296 & n12408;
  assign n12410 = n33269 & ~n12404;
  assign n12411 = ~n12409 & ~n12410;
  assign n12412 = ~n12405 & ~n12406;
  assign n12413 = ~n33340 & ~n33341;
  assign n12414 = ~n12399 & ~n12413;
  assign n12415 = ~n7885 & ~n12414;
  assign n12416 = n7885 & ~n12399;
  assign n12417 = ~n12413 & n12416;
  assign n12418 = ~n33270 & ~n11829;
  assign n12419 = ~n11829 & ~n12296;
  assign n12420 = ~n33270 & n12419;
  assign n12421 = ~n12296 & n12418;
  assign n12422 = n11743 & ~n33342;
  assign n12423 = n11828 & n12419;
  assign n12424 = n11743 & ~n33270;
  assign n12425 = ~n11829 & n12424;
  assign n12426 = ~n12296 & n12425;
  assign n12427 = ~n11743 & ~n33342;
  assign n12428 = ~n12426 & ~n12427;
  assign n12429 = ~n12422 & ~n12423;
  assign n12430 = ~n12417 & ~n33343;
  assign n12431 = ~n12415 & ~n12430;
  assign n12432 = ~n7428 & ~n12431;
  assign n12433 = n7428 & ~n12415;
  assign n12434 = ~n12430 & n12433;
  assign n12435 = n7428 & n12431;
  assign n12436 = ~n11831 & ~n11844;
  assign n12437 = ~n12296 & n12436;
  assign n12438 = ~n33271 & n12437;
  assign n12439 = n33271 & ~n12437;
  assign n12440 = n33271 & ~n11844;
  assign n12441 = ~n11831 & n12440;
  assign n12442 = ~n12296 & n12441;
  assign n12443 = ~n33271 & ~n12437;
  assign n12444 = ~n12442 & ~n12443;
  assign n12445 = ~n12438 & ~n12439;
  assign n12446 = ~n33344 & ~n33345;
  assign n12447 = ~n12432 & ~n12446;
  assign n12448 = ~n6937 & ~n12447;
  assign n12449 = n6937 & ~n12432;
  assign n12450 = ~n12446 & n12449;
  assign n12451 = ~n33272 & ~n11850;
  assign n12452 = ~n11850 & ~n12296;
  assign n12453 = ~n33272 & n12452;
  assign n12454 = ~n12296 & n12451;
  assign n12455 = n11735 & ~n33346;
  assign n12456 = n11849 & n12452;
  assign n12457 = n11735 & ~n33272;
  assign n12458 = ~n11850 & n12457;
  assign n12459 = ~n12296 & n12458;
  assign n12460 = ~n11735 & ~n33346;
  assign n12461 = ~n12459 & ~n12460;
  assign n12462 = ~n12455 & ~n12456;
  assign n12463 = ~n12450 & ~n33347;
  assign n12464 = ~n12448 & ~n12463;
  assign n12465 = ~n6507 & ~n12464;
  assign n12466 = n6507 & ~n12448;
  assign n12467 = ~n12463 & n12466;
  assign n12468 = n6507 & n12464;
  assign n12469 = ~n11852 & ~n11865;
  assign n12470 = ~n12296 & n12469;
  assign n12471 = ~n33273 & n12470;
  assign n12472 = n33273 & ~n12470;
  assign n12473 = ~n33273 & ~n12470;
  assign n12474 = n33273 & ~n11865;
  assign n12475 = ~n11852 & n12474;
  assign n12476 = n33273 & n12470;
  assign n12477 = ~n12296 & n12475;
  assign n12478 = ~n12473 & ~n33349;
  assign n12479 = ~n12471 & ~n12472;
  assign n12480 = ~n33348 & ~n33350;
  assign n12481 = ~n12465 & ~n12480;
  assign n12482 = ~n6051 & ~n12481;
  assign n12483 = n6051 & ~n12465;
  assign n12484 = ~n12480 & n12483;
  assign n12485 = ~n33274 & ~n11871;
  assign n12486 = ~n11871 & ~n12296;
  assign n12487 = ~n33274 & n12486;
  assign n12488 = ~n12296 & n12485;
  assign n12489 = n11727 & ~n33351;
  assign n12490 = n11870 & n12486;
  assign n12491 = n11727 & ~n33274;
  assign n12492 = ~n11871 & n12491;
  assign n12493 = ~n12296 & n12492;
  assign n12494 = ~n11727 & ~n33351;
  assign n12495 = ~n12493 & ~n12494;
  assign n12496 = ~n12489 & ~n12490;
  assign n12497 = ~n12484 & ~n33352;
  assign n12498 = ~n12482 & ~n12497;
  assign n12499 = ~n5648 & ~n12498;
  assign n12500 = n5648 & ~n12482;
  assign n12501 = ~n12497 & n12500;
  assign n12502 = n5648 & n12498;
  assign n12503 = ~n11873 & ~n11887;
  assign n12504 = ~n11887 & ~n12296;
  assign n12505 = ~n11873 & n12504;
  assign n12506 = ~n12296 & n12503;
  assign n12507 = n33276 & ~n33354;
  assign n12508 = n11885 & n12504;
  assign n12509 = ~n33276 & n33354;
  assign n12510 = n33276 & ~n11887;
  assign n12511 = ~n11873 & n12510;
  assign n12512 = ~n12296 & n12511;
  assign n12513 = ~n33276 & ~n33354;
  assign n12514 = ~n12512 & ~n12513;
  assign n12515 = ~n12507 & ~n33355;
  assign n12516 = ~n33353 & ~n33356;
  assign n12517 = ~n12499 & ~n12516;
  assign n12518 = ~n5223 & ~n12517;
  assign n12519 = n5223 & ~n12499;
  assign n12520 = ~n12516 & n12519;
  assign n12521 = ~n33277 & ~n11903;
  assign n12522 = ~n12296 & n12521;
  assign n12523 = ~n33278 & n12522;
  assign n12524 = n33278 & ~n12522;
  assign n12525 = ~n33277 & n33278;
  assign n12526 = ~n11903 & n12525;
  assign n12527 = ~n12296 & n12526;
  assign n12528 = ~n33278 & ~n12522;
  assign n12529 = ~n12527 & ~n12528;
  assign n12530 = ~n12523 & ~n12524;
  assign n12531 = ~n12520 & ~n33357;
  assign n12532 = ~n12518 & ~n12531;
  assign n12533 = ~n4851 & ~n12532;
  assign n12534 = ~n11905 & ~n11917;
  assign n12535 = ~n12296 & n12534;
  assign n12536 = ~n33279 & ~n12535;
  assign n12537 = ~n11905 & n33279;
  assign n12538 = ~n11917 & n12537;
  assign n12539 = n33279 & n12535;
  assign n12540 = ~n12296 & n12538;
  assign n12541 = ~n12536 & ~n33358;
  assign n12542 = n4851 & ~n12518;
  assign n12543 = ~n12531 & n12542;
  assign n12544 = n4851 & n12532;
  assign n12545 = ~n12541 & ~n33359;
  assign n12546 = ~n12533 & ~n12545;
  assign n12547 = ~n4461 & ~n12546;
  assign n12548 = n4461 & ~n12533;
  assign n12549 = ~n12545 & n12548;
  assign n12550 = ~n11920 & ~n33281;
  assign n12551 = ~n11920 & ~n12296;
  assign n12552 = ~n33281 & n12551;
  assign n12553 = ~n12296 & n12550;
  assign n12554 = n11928 & ~n33360;
  assign n12555 = n11932 & n12551;
  assign n12556 = n11928 & ~n33281;
  assign n12557 = ~n11920 & n12556;
  assign n12558 = ~n12296 & n12557;
  assign n12559 = ~n11928 & ~n33360;
  assign n12560 = ~n12558 & ~n12559;
  assign n12561 = ~n12554 & ~n12555;
  assign n12562 = ~n12549 & ~n33361;
  assign n12563 = ~n12547 & ~n12562;
  assign n12564 = ~n4115 & ~n12563;
  assign n12565 = ~n11934 & ~n11936;
  assign n12566 = ~n12296 & n12565;
  assign n12567 = n33284 & ~n12566;
  assign n12568 = ~n11934 & ~n33284;
  assign n12569 = ~n11936 & n12568;
  assign n12570 = ~n33284 & n12566;
  assign n12571 = ~n12296 & n12569;
  assign n12572 = ~n12567 & ~n33362;
  assign n12573 = n4115 & ~n12547;
  assign n12574 = ~n12562 & n12573;
  assign n12575 = n4115 & n12563;
  assign n12576 = ~n12572 & ~n33363;
  assign n12577 = ~n12564 & ~n12576;
  assign n12578 = ~n3754 & ~n12577;
  assign n12579 = n3754 & ~n12564;
  assign n12580 = ~n12576 & n12579;
  assign n12581 = ~n11952 & ~n33286;
  assign n12582 = ~n11952 & ~n12296;
  assign n12583 = ~n33286 & n12582;
  assign n12584 = ~n12296 & n12581;
  assign n12585 = n11960 & ~n33364;
  assign n12586 = n11964 & n12582;
  assign n12587 = n11960 & ~n33286;
  assign n12588 = ~n11952 & n12587;
  assign n12589 = ~n12296 & n12588;
  assign n12590 = ~n11960 & ~n33364;
  assign n12591 = ~n12589 & ~n12590;
  assign n12592 = ~n12585 & ~n12586;
  assign n12593 = ~n12580 & ~n33365;
  assign n12594 = ~n12578 & ~n12593;
  assign n12595 = ~n3444 & ~n12594;
  assign n12596 = ~n11966 & ~n11968;
  assign n12597 = ~n12296 & n12596;
  assign n12598 = ~n33288 & ~n12597;
  assign n12599 = ~n11966 & n33288;
  assign n12600 = ~n11968 & n12599;
  assign n12601 = n33288 & n12597;
  assign n12602 = ~n12296 & n12600;
  assign n12603 = ~n12598 & ~n33366;
  assign n12604 = n3444 & ~n12578;
  assign n12605 = ~n12593 & n12604;
  assign n12606 = n3444 & n12594;
  assign n12607 = ~n12603 & ~n33367;
  assign n12608 = ~n12595 & ~n12607;
  assign n12609 = ~n3116 & ~n12608;
  assign n12610 = n3116 & ~n12595;
  assign n12611 = ~n12607 & n12610;
  assign n12612 = ~n11983 & ~n33290;
  assign n12613 = ~n11983 & ~n12296;
  assign n12614 = ~n33290 & n12613;
  assign n12615 = ~n12296 & n12612;
  assign n12616 = n11991 & ~n33368;
  assign n12617 = n11995 & n12613;
  assign n12618 = n11991 & ~n33290;
  assign n12619 = ~n11983 & n12618;
  assign n12620 = ~n12296 & n12619;
  assign n12621 = ~n11991 & ~n33368;
  assign n12622 = ~n12620 & ~n12621;
  assign n12623 = ~n12616 & ~n12617;
  assign n12624 = ~n12611 & ~n33369;
  assign n12625 = ~n12609 & ~n12624;
  assign n12626 = ~n2833 & ~n12625;
  assign n12627 = n2833 & ~n12609;
  assign n12628 = ~n12624 & n12627;
  assign n12629 = n2833 & n12625;
  assign n12630 = ~n11997 & ~n12007;
  assign n12631 = ~n11997 & ~n12296;
  assign n12632 = ~n12007 & n12631;
  assign n12633 = ~n12296 & n12630;
  assign n12634 = n12005 & ~n33371;
  assign n12635 = n12008 & n12631;
  assign n12636 = ~n11997 & n12005;
  assign n12637 = ~n12007 & n12636;
  assign n12638 = ~n12296 & n12637;
  assign n12639 = ~n12005 & ~n33371;
  assign n12640 = ~n12638 & ~n12639;
  assign n12641 = ~n12634 & ~n12635;
  assign n12642 = ~n33370 & ~n33372;
  assign n12643 = ~n12626 & ~n12642;
  assign n12644 = ~n2536 & ~n12643;
  assign n12645 = n2536 & ~n12626;
  assign n12646 = ~n12642 & n12645;
  assign n12647 = ~n12010 & ~n33293;
  assign n12648 = ~n12010 & ~n12296;
  assign n12649 = ~n33293 & n12648;
  assign n12650 = ~n12296 & n12647;
  assign n12651 = n12018 & ~n33373;
  assign n12652 = n12022 & n12648;
  assign n12653 = n12018 & ~n33293;
  assign n12654 = ~n12010 & n12653;
  assign n12655 = ~n12296 & n12654;
  assign n12656 = ~n12018 & ~n33373;
  assign n12657 = ~n12655 & ~n12656;
  assign n12658 = ~n12651 & ~n12652;
  assign n12659 = ~n12646 & ~n33374;
  assign n12660 = ~n12644 & ~n12659;
  assign n12661 = ~n2283 & ~n12660;
  assign n12662 = ~n12024 & ~n12026;
  assign n12663 = ~n12296 & n12662;
  assign n12664 = ~n33295 & ~n12663;
  assign n12665 = ~n12024 & n33295;
  assign n12666 = ~n12026 & n12665;
  assign n12667 = n33295 & n12663;
  assign n12668 = ~n12296 & n12666;
  assign n12669 = ~n12664 & ~n33375;
  assign n12670 = n2283 & ~n12644;
  assign n12671 = ~n12659 & n12670;
  assign n12672 = n2283 & n12660;
  assign n12673 = ~n12669 & ~n33376;
  assign n12674 = ~n12661 & ~n12673;
  assign n12675 = ~n2021 & ~n12674;
  assign n12676 = n2021 & ~n12661;
  assign n12677 = ~n12673 & n12676;
  assign n12678 = ~n12041 & ~n33297;
  assign n12679 = ~n12041 & ~n12296;
  assign n12680 = ~n33297 & n12679;
  assign n12681 = ~n12296 & n12678;
  assign n12682 = n12049 & ~n33377;
  assign n12683 = n12053 & n12679;
  assign n12684 = n12049 & ~n33297;
  assign n12685 = ~n12041 & n12684;
  assign n12686 = ~n12296 & n12685;
  assign n12687 = ~n12049 & ~n33377;
  assign n12688 = ~n12686 & ~n12687;
  assign n12689 = ~n12682 & ~n12683;
  assign n12690 = ~n12677 & ~n33378;
  assign n12691 = ~n12675 & ~n12690;
  assign n12692 = ~n1796 & ~n12691;
  assign n12693 = n1796 & ~n12675;
  assign n12694 = ~n12690 & n12693;
  assign n12695 = n1796 & n12691;
  assign n12696 = ~n12055 & ~n12065;
  assign n12697 = ~n12055 & ~n12296;
  assign n12698 = ~n12065 & n12697;
  assign n12699 = ~n12296 & n12696;
  assign n12700 = n12063 & ~n33380;
  assign n12701 = n12066 & n12697;
  assign n12702 = ~n12055 & n12063;
  assign n12703 = ~n12065 & n12702;
  assign n12704 = ~n12296 & n12703;
  assign n12705 = ~n12063 & ~n33380;
  assign n12706 = ~n12704 & ~n12705;
  assign n12707 = ~n12700 & ~n12701;
  assign n12708 = ~n33379 & ~n33381;
  assign n12709 = ~n12692 & ~n12708;
  assign n12710 = ~n1567 & ~n12709;
  assign n12711 = n1567 & ~n12692;
  assign n12712 = ~n12708 & n12711;
  assign n12713 = ~n12068 & ~n33300;
  assign n12714 = ~n12068 & ~n12296;
  assign n12715 = ~n33300 & n12714;
  assign n12716 = ~n12296 & n12713;
  assign n12717 = n12076 & ~n33382;
  assign n12718 = n12080 & n12714;
  assign n12719 = n12076 & ~n33300;
  assign n12720 = ~n12068 & n12719;
  assign n12721 = ~n12296 & n12720;
  assign n12722 = ~n12076 & ~n33382;
  assign n12723 = ~n12721 & ~n12722;
  assign n12724 = ~n12717 & ~n12718;
  assign n12725 = ~n12712 & ~n33383;
  assign n12726 = ~n12710 & ~n12725;
  assign n12727 = ~n1374 & ~n12726;
  assign n12728 = ~n12082 & ~n12084;
  assign n12729 = ~n12296 & n12728;
  assign n12730 = ~n33302 & ~n12729;
  assign n12731 = ~n12082 & n33302;
  assign n12732 = ~n12084 & n12731;
  assign n12733 = n33302 & n12729;
  assign n12734 = ~n12296 & n12732;
  assign n12735 = ~n12730 & ~n33384;
  assign n12736 = n1374 & ~n12710;
  assign n12737 = ~n12725 & n12736;
  assign n12738 = n1374 & n12726;
  assign n12739 = ~n12735 & ~n33385;
  assign n12740 = ~n12727 & ~n12739;
  assign n12741 = ~n1179 & ~n12740;
  assign n12742 = n1179 & ~n12727;
  assign n12743 = ~n12739 & n12742;
  assign n12744 = ~n12099 & ~n33304;
  assign n12745 = ~n12099 & ~n12296;
  assign n12746 = ~n33304 & n12745;
  assign n12747 = ~n12296 & n12744;
  assign n12748 = n12107 & ~n33386;
  assign n12749 = n12111 & n12745;
  assign n12750 = n12107 & ~n33304;
  assign n12751 = ~n12099 & n12750;
  assign n12752 = ~n12296 & n12751;
  assign n12753 = ~n12107 & ~n33386;
  assign n12754 = ~n12752 & ~n12753;
  assign n12755 = ~n12748 & ~n12749;
  assign n12756 = ~n12743 & ~n33387;
  assign n12757 = ~n12741 & ~n12756;
  assign n12758 = ~n1016 & ~n12757;
  assign n12759 = n1016 & ~n12741;
  assign n12760 = ~n12756 & n12759;
  assign n12761 = n1016 & n12757;
  assign n12762 = ~n12113 & ~n12123;
  assign n12763 = ~n12113 & ~n12296;
  assign n12764 = ~n12123 & n12763;
  assign n12765 = ~n12296 & n12762;
  assign n12766 = n12121 & ~n33389;
  assign n12767 = n12124 & n12763;
  assign n12768 = ~n12113 & n12121;
  assign n12769 = ~n12123 & n12768;
  assign n12770 = ~n12296 & n12769;
  assign n12771 = ~n12121 & ~n33389;
  assign n12772 = ~n12770 & ~n12771;
  assign n12773 = ~n12766 & ~n12767;
  assign n12774 = ~n33388 & ~n33390;
  assign n12775 = ~n12758 & ~n12774;
  assign n12776 = ~n855 & ~n12775;
  assign n12777 = n855 & ~n12758;
  assign n12778 = ~n12774 & n12777;
  assign n12779 = ~n12126 & ~n33307;
  assign n12780 = ~n12126 & ~n12296;
  assign n12781 = ~n33307 & n12780;
  assign n12782 = ~n12296 & n12779;
  assign n12783 = n12134 & ~n33391;
  assign n12784 = n12138 & n12780;
  assign n12785 = n12134 & ~n33307;
  assign n12786 = ~n12126 & n12785;
  assign n12787 = ~n12296 & n12786;
  assign n12788 = ~n12134 & ~n33391;
  assign n12789 = ~n12787 & ~n12788;
  assign n12790 = ~n12783 & ~n12784;
  assign n12791 = ~n12778 & ~n33392;
  assign n12792 = ~n12776 & ~n12791;
  assign n12793 = ~n720 & ~n12792;
  assign n12794 = ~n12140 & ~n12142;
  assign n12795 = ~n12296 & n12794;
  assign n12796 = ~n33309 & ~n12795;
  assign n12797 = ~n12140 & n33309;
  assign n12798 = ~n12142 & n12797;
  assign n12799 = n33309 & n12795;
  assign n12800 = ~n12296 & n12798;
  assign n12801 = ~n12796 & ~n33393;
  assign n12802 = n720 & ~n12776;
  assign n12803 = ~n12791 & n12802;
  assign n12804 = n720 & n12792;
  assign n12805 = ~n12801 & ~n33394;
  assign n12806 = ~n12793 & ~n12805;
  assign n12807 = ~n592 & ~n12806;
  assign n12808 = n592 & ~n12793;
  assign n12809 = ~n12805 & n12808;
  assign n12810 = ~n12157 & ~n33311;
  assign n12811 = ~n12157 & ~n12296;
  assign n12812 = ~n33311 & n12811;
  assign n12813 = ~n12296 & n12810;
  assign n12814 = n12165 & ~n33395;
  assign n12815 = n12169 & n12811;
  assign n12816 = n12165 & ~n33311;
  assign n12817 = ~n12157 & n12816;
  assign n12818 = ~n12296 & n12817;
  assign n12819 = ~n12165 & ~n33395;
  assign n12820 = ~n12818 & ~n12819;
  assign n12821 = ~n12814 & ~n12815;
  assign n12822 = ~n12809 & ~n33396;
  assign n12823 = ~n12807 & ~n12822;
  assign n12824 = ~n487 & ~n12823;
  assign n12825 = n487 & ~n12807;
  assign n12826 = ~n12822 & n12825;
  assign n12827 = n487 & n12823;
  assign n12828 = ~n12171 & ~n12181;
  assign n12829 = ~n12171 & ~n12296;
  assign n12830 = ~n12181 & n12829;
  assign n12831 = ~n12296 & n12828;
  assign n12832 = n12179 & ~n33398;
  assign n12833 = n12182 & n12829;
  assign n12834 = ~n12171 & n12179;
  assign n12835 = ~n12181 & n12834;
  assign n12836 = ~n12296 & n12835;
  assign n12837 = ~n12179 & ~n33398;
  assign n12838 = ~n12836 & ~n12837;
  assign n12839 = ~n12832 & ~n12833;
  assign n12840 = ~n33397 & ~n33399;
  assign n12841 = ~n12824 & ~n12840;
  assign n12842 = ~n393 & ~n12841;
  assign n12843 = n393 & ~n12824;
  assign n12844 = ~n12840 & n12843;
  assign n12845 = ~n12184 & ~n33314;
  assign n12846 = ~n12184 & ~n12296;
  assign n12847 = ~n33314 & n12846;
  assign n12848 = ~n12296 & n12845;
  assign n12849 = n12192 & ~n33400;
  assign n12850 = n12196 & n12846;
  assign n12851 = n12192 & ~n33314;
  assign n12852 = ~n12184 & n12851;
  assign n12853 = ~n12296 & n12852;
  assign n12854 = ~n12192 & ~n33400;
  assign n12855 = ~n12853 & ~n12854;
  assign n12856 = ~n12849 & ~n12850;
  assign n12857 = ~n12844 & ~n33401;
  assign n12858 = ~n12842 & ~n12857;
  assign n12859 = ~n321 & ~n12858;
  assign n12860 = ~n12198 & ~n12200;
  assign n12861 = ~n12296 & n12860;
  assign n12862 = ~n33316 & ~n12861;
  assign n12863 = ~n12198 & n33316;
  assign n12864 = ~n12200 & n12863;
  assign n12865 = n33316 & n12861;
  assign n12866 = ~n12296 & n12864;
  assign n12867 = ~n12862 & ~n33402;
  assign n12868 = n321 & ~n12842;
  assign n12869 = ~n12857 & n12868;
  assign n12870 = n321 & n12858;
  assign n12871 = ~n12867 & ~n33403;
  assign n12872 = ~n12859 & ~n12871;
  assign n12873 = ~n263 & ~n12872;
  assign n12874 = n263 & ~n12859;
  assign n12875 = ~n12871 & n12874;
  assign n12876 = ~n12215 & ~n33318;
  assign n12877 = ~n12215 & ~n12296;
  assign n12878 = ~n33318 & n12877;
  assign n12879 = ~n12296 & n12876;
  assign n12880 = n12223 & ~n33404;
  assign n12881 = n12227 & n12877;
  assign n12882 = n12223 & ~n33318;
  assign n12883 = ~n12215 & n12882;
  assign n12884 = ~n12296 & n12883;
  assign n12885 = ~n12223 & ~n33404;
  assign n12886 = ~n12884 & ~n12885;
  assign n12887 = ~n12880 & ~n12881;
  assign n12888 = ~n12875 & ~n33405;
  assign n12889 = ~n12873 & ~n12888;
  assign n12890 = ~n214 & ~n12889;
  assign n12891 = n214 & ~n12873;
  assign n12892 = ~n12888 & n12891;
  assign n12893 = n214 & n12889;
  assign n12894 = ~n12229 & ~n12239;
  assign n12895 = ~n12229 & ~n12296;
  assign n12896 = ~n12239 & n12895;
  assign n12897 = ~n12296 & n12894;
  assign n12898 = n12237 & ~n33407;
  assign n12899 = n12240 & n12895;
  assign n12900 = ~n12229 & n12237;
  assign n12901 = ~n12239 & n12900;
  assign n12902 = ~n12296 & n12901;
  assign n12903 = ~n12237 & ~n33407;
  assign n12904 = ~n12902 & ~n12903;
  assign n12905 = ~n12898 & ~n12899;
  assign n12906 = ~n33406 & ~n33408;
  assign n12907 = ~n12890 & ~n12906;
  assign n12908 = ~n197 & ~n12907;
  assign n12909 = n197 & ~n12890;
  assign n12910 = ~n12906 & n12909;
  assign n12911 = ~n12242 & ~n33321;
  assign n12912 = ~n12242 & ~n12296;
  assign n12913 = ~n33321 & n12912;
  assign n12914 = ~n12296 & n12911;
  assign n12915 = n12250 & ~n33409;
  assign n12916 = n12254 & n12912;
  assign n12917 = n12250 & ~n33321;
  assign n12918 = ~n12242 & n12917;
  assign n12919 = ~n12296 & n12918;
  assign n12920 = ~n12250 & ~n33409;
  assign n12921 = ~n12919 & ~n12920;
  assign n12922 = ~n12915 & ~n12916;
  assign n12923 = ~n12910 & ~n33410;
  assign n12924 = ~n12908 & ~n12923;
  assign n12925 = ~n12256 & ~n12258;
  assign n12926 = ~n12296 & n12925;
  assign n12927 = ~n33323 & ~n12926;
  assign n12928 = ~n12256 & n33323;
  assign n12929 = ~n12258 & n12928;
  assign n12930 = n33323 & n12926;
  assign n12931 = ~n12296 & n12929;
  assign n12932 = ~n12927 & ~n33411;
  assign n12933 = ~n12272 & ~n12280;
  assign n12934 = ~n12280 & ~n12296;
  assign n12935 = ~n12272 & n12934;
  assign n12936 = ~n12296 & n12933;
  assign n12937 = ~n33326 & ~n33412;
  assign n12938 = ~n12932 & n12937;
  assign n12939 = ~n12924 & n12938;
  assign n12940 = n193 & ~n12939;
  assign n12941 = ~n12908 & n12932;
  assign n12942 = ~n12923 & n12941;
  assign n12943 = n12924 & n12932;
  assign n12944 = n12272 & ~n12934;
  assign n12945 = ~n193 & ~n12933;
  assign n12946 = ~n12944 & n12945;
  assign n12947 = ~n33413 & ~n12946;
  assign n12948 = ~n12940 & n12947;
  assign n12949 = ~n12518 & ~n12520;
  assign n12950 = ~n12948 & n12949;
  assign n12951 = ~n33357 & ~n12950;
  assign n12952 = ~n12520 & n33357;
  assign n12953 = ~n12518 & n12952;
  assign n12954 = n33357 & n12950;
  assign n12955 = ~n12948 & n12953;
  assign n12956 = ~n12951 & ~n33414;
  assign n12957 = ~n12499 & ~n33353;
  assign n12958 = ~n12948 & n12957;
  assign n12959 = ~n33356 & ~n12958;
  assign n12960 = ~n12499 & n33356;
  assign n12961 = ~n33353 & n12960;
  assign n12962 = n33356 & n12958;
  assign n12963 = ~n12948 & n12961;
  assign n12964 = ~n12959 & ~n33415;
  assign n12965 = ~n12482 & ~n12484;
  assign n12966 = ~n12948 & n12965;
  assign n12967 = ~n33352 & ~n12966;
  assign n12968 = ~n12484 & n33352;
  assign n12969 = ~n12482 & n12968;
  assign n12970 = n33352 & n12966;
  assign n12971 = ~n12948 & n12969;
  assign n12972 = ~n12967 & ~n33416;
  assign n12973 = ~n12448 & ~n12450;
  assign n12974 = ~n12948 & n12973;
  assign n12975 = ~n33347 & ~n12974;
  assign n12976 = ~n12450 & n33347;
  assign n12977 = ~n12448 & n12976;
  assign n12978 = n33347 & n12974;
  assign n12979 = ~n12948 & n12977;
  assign n12980 = ~n12975 & ~n33417;
  assign n12981 = ~n12415 & ~n12417;
  assign n12982 = ~n12948 & n12981;
  assign n12983 = ~n33343 & ~n12982;
  assign n12984 = ~n12417 & n33343;
  assign n12985 = ~n12415 & n12984;
  assign n12986 = n33343 & n12982;
  assign n12987 = ~n12948 & n12985;
  assign n12988 = ~n12983 & ~n33418;
  assign n12989 = ~n12382 & ~n12384;
  assign n12990 = ~n12948 & n12989;
  assign n12991 = ~n33339 & ~n12990;
  assign n12992 = ~n12384 & n33339;
  assign n12993 = ~n12382 & n12992;
  assign n12994 = n33339 & n12990;
  assign n12995 = ~n12948 & n12993;
  assign n12996 = ~n12991 & ~n33419;
  assign n12997 = ~n12348 & ~n12350;
  assign n12998 = ~n12948 & n12997;
  assign n12999 = ~n33334 & ~n12998;
  assign n13000 = ~n12350 & n33334;
  assign n13001 = ~n12348 & n13000;
  assign n13002 = n33334 & n12998;
  assign n13003 = ~n12948 & n13001;
  assign n13004 = ~n12999 & ~n33420;
  assign n13005 = ~n12321 & ~n12323;
  assign n13006 = ~n12948 & n13005;
  assign n13007 = ~n12332 & ~n13006;
  assign n13008 = ~n12323 & n12332;
  assign n13009 = ~n12321 & n13008;
  assign n13010 = n12332 & n13006;
  assign n13011 = ~n12948 & n13009;
  assign n13012 = ~n13007 & ~n33421;
  assign n13013 = ~pi46  & ~n12948;
  assign n13014 = ~pi47  & n13013;
  assign n13015 = n12298 & ~n12948;
  assign n13016 = ~n12296 & ~n12946;
  assign n13017 = ~n33413 & n13016;
  assign n13018 = ~n12940 & n13017;
  assign n13019 = ~n33422 & ~n13018;
  assign n13020 = pi48  & ~n13019;
  assign n13021 = ~pi48  & ~n13018;
  assign n13022 = ~pi48  & n13019;
  assign n13023 = ~n33422 & n13021;
  assign n13024 = ~n13020 & ~n33423;
  assign n13025 = pi46  & ~n12948;
  assign n13026 = ~pi44  & ~pi45 ;
  assign n13027 = ~pi46  & n13026;
  assign n13028 = ~n11700 & ~n33328;
  assign n13029 = ~n11701 & n13028;
  assign n13030 = ~n11717 & n13029;
  assign n13031 = ~n33256 & n13030;
  assign n13032 = n33254 & n11719;
  assign n13033 = ~n11711 & n13031;
  assign n13034 = ~n13027 & ~n33424;
  assign n13035 = ~n12294 & n13034;
  assign n13036 = ~n33326 & n13035;
  assign n13037 = ~n12288 & n13036;
  assign n13038 = ~n13025 & ~n13027;
  assign n13039 = n12296 & n13038;
  assign n13040 = ~n13025 & n13037;
  assign n13041 = pi47  & ~n13013;
  assign n13042 = ~n33422 & ~n13041;
  assign n13043 = ~n33425 & n13042;
  assign n13044 = ~n12296 & ~n13038;
  assign n13045 = n11719 & ~n13044;
  assign n13046 = ~n13043 & ~n13044;
  assign n13047 = n11719 & n13046;
  assign n13048 = ~n13043 & n13045;
  assign n13049 = ~n13024 & ~n33426;
  assign n13050 = ~n11719 & ~n13046;
  assign n13051 = n11097 & ~n13050;
  assign n13052 = ~n13049 & n13051;
  assign n13053 = ~n12301 & ~n33329;
  assign n13054 = ~n12948 & n13053;
  assign n13055 = n12306 & ~n13054;
  assign n13056 = ~n12306 & n13053;
  assign n13057 = ~n12306 & n13054;
  assign n13058 = ~n12948 & n13056;
  assign n13059 = ~n13055 & ~n33427;
  assign n13060 = ~n13052 & ~n13059;
  assign n13061 = ~n13049 & ~n13050;
  assign n13062 = ~n11097 & ~n13061;
  assign n13063 = n10555 & ~n13062;
  assign n13064 = ~n13060 & ~n13062;
  assign n13065 = n10555 & n13064;
  assign n13066 = ~n13060 & n13063;
  assign n13067 = ~n13012 & ~n33428;
  assign n13068 = ~n10555 & ~n13064;
  assign n13069 = n9969 & ~n13068;
  assign n13070 = ~n13067 & n13069;
  assign n13071 = ~n12335 & ~n33331;
  assign n13072 = ~n12948 & n13071;
  assign n13073 = ~n12345 & ~n13072;
  assign n13074 = ~n12335 & n12345;
  assign n13075 = ~n33331 & n13074;
  assign n13076 = n12345 & n13072;
  assign n13077 = ~n12948 & n13075;
  assign n13078 = n12345 & ~n13072;
  assign n13079 = ~n12345 & n13072;
  assign n13080 = ~n13078 & ~n13079;
  assign n13081 = ~n13073 & ~n33429;
  assign n13082 = ~n13070 & n33430;
  assign n13083 = ~n13067 & ~n13068;
  assign n13084 = ~n9969 & ~n13083;
  assign n13085 = n9457 & ~n13084;
  assign n13086 = ~n13082 & ~n13084;
  assign n13087 = n9457 & n13086;
  assign n13088 = ~n13082 & n13085;
  assign n13089 = ~n13004 & ~n33431;
  assign n13090 = ~n9457 & ~n13086;
  assign n13091 = n8896 & ~n13090;
  assign n13092 = ~n13089 & n13091;
  assign n13093 = ~n12365 & ~n33335;
  assign n13094 = ~n12948 & n13093;
  assign n13095 = ~n33337 & ~n13094;
  assign n13096 = n33337 & n13094;
  assign n13097 = ~n12365 & ~n33337;
  assign n13098 = ~n33335 & n13097;
  assign n13099 = ~n12948 & n13098;
  assign n13100 = n33337 & ~n13094;
  assign n13101 = ~n13099 & ~n13100;
  assign n13102 = ~n13095 & ~n13096;
  assign n13103 = ~n13092 & ~n33432;
  assign n13104 = ~n13089 & ~n13090;
  assign n13105 = ~n8896 & ~n13104;
  assign n13106 = n8411 & ~n13105;
  assign n13107 = ~n13103 & ~n13105;
  assign n13108 = n8411 & n13107;
  assign n13109 = ~n13103 & n13106;
  assign n13110 = ~n12996 & ~n33433;
  assign n13111 = ~n8411 & ~n13107;
  assign n13112 = n7885 & ~n13111;
  assign n13113 = ~n13110 & n13112;
  assign n13114 = ~n12399 & ~n33340;
  assign n13115 = ~n12948 & n13114;
  assign n13116 = ~n33341 & n13115;
  assign n13117 = n33341 & ~n13115;
  assign n13118 = ~n12399 & n33341;
  assign n13119 = ~n33340 & n13118;
  assign n13120 = ~n12948 & n13119;
  assign n13121 = ~n33341 & ~n13115;
  assign n13122 = ~n13120 & ~n13121;
  assign n13123 = ~n13116 & ~n13117;
  assign n13124 = ~n13113 & ~n33434;
  assign n13125 = ~n13110 & ~n13111;
  assign n13126 = ~n7885 & ~n13125;
  assign n13127 = n7428 & ~n13126;
  assign n13128 = ~n13124 & ~n13126;
  assign n13129 = n7428 & n13128;
  assign n13130 = ~n13124 & n13127;
  assign n13131 = ~n12988 & ~n33435;
  assign n13132 = ~n7428 & ~n13128;
  assign n13133 = n6937 & ~n13132;
  assign n13134 = ~n13131 & n13133;
  assign n13135 = ~n12432 & ~n33344;
  assign n13136 = ~n12948 & n13135;
  assign n13137 = ~n33345 & n13136;
  assign n13138 = n33345 & ~n13136;
  assign n13139 = ~n33345 & ~n13136;
  assign n13140 = ~n12432 & n33345;
  assign n13141 = ~n33344 & n13140;
  assign n13142 = n33345 & n13136;
  assign n13143 = ~n12948 & n13141;
  assign n13144 = ~n13139 & ~n33436;
  assign n13145 = ~n13137 & ~n13138;
  assign n13146 = ~n13134 & ~n33437;
  assign n13147 = ~n13131 & ~n13132;
  assign n13148 = ~n6937 & ~n13147;
  assign n13149 = n6507 & ~n13148;
  assign n13150 = ~n13146 & ~n13148;
  assign n13151 = n6507 & n13150;
  assign n13152 = ~n13146 & n13149;
  assign n13153 = ~n12980 & ~n33438;
  assign n13154 = ~n6507 & ~n13150;
  assign n13155 = n6051 & ~n13154;
  assign n13156 = ~n13153 & n13155;
  assign n13157 = ~n12465 & ~n33348;
  assign n13158 = ~n12465 & ~n12948;
  assign n13159 = ~n33348 & n13158;
  assign n13160 = ~n12948 & n13157;
  assign n13161 = n33350 & ~n33439;
  assign n13162 = n12480 & n13158;
  assign n13163 = ~n33350 & n33439;
  assign n13164 = ~n12465 & n33350;
  assign n13165 = ~n33348 & n13164;
  assign n13166 = ~n12948 & n13165;
  assign n13167 = ~n33350 & ~n33439;
  assign n13168 = ~n13166 & ~n13167;
  assign n13169 = ~n13161 & ~n33440;
  assign n13170 = ~n13156 & ~n33441;
  assign n13171 = ~n13153 & ~n13154;
  assign n13172 = ~n6051 & ~n13171;
  assign n13173 = n5648 & ~n13172;
  assign n13174 = ~n13170 & ~n13172;
  assign n13175 = n5648 & n13174;
  assign n13176 = ~n13170 & n13173;
  assign n13177 = ~n12972 & ~n33442;
  assign n13178 = ~n5648 & ~n13174;
  assign n13179 = n5223 & ~n13178;
  assign n13180 = ~n13177 & n13179;
  assign n13181 = ~n12964 & ~n13180;
  assign n13182 = ~n13177 & ~n13178;
  assign n13183 = ~n5223 & ~n13182;
  assign n13184 = n4851 & ~n13183;
  assign n13185 = ~n13181 & ~n13183;
  assign n13186 = n4851 & n13185;
  assign n13187 = ~n13181 & n13184;
  assign n13188 = ~n12956 & ~n33443;
  assign n13189 = ~n4851 & ~n13185;
  assign n13190 = ~n13188 & ~n13189;
  assign n13191 = ~n4461 & ~n13190;
  assign n13192 = ~n12533 & n12541;
  assign n13193 = ~n33359 & n13192;
  assign n13194 = ~n12533 & ~n33359;
  assign n13195 = ~n12948 & n13194;
  assign n13196 = n12541 & n13195;
  assign n13197 = ~n12948 & n13193;
  assign n13198 = ~n12541 & ~n13195;
  assign n13199 = ~n33444 & ~n13198;
  assign n13200 = n4461 & ~n13189;
  assign n13201 = ~n13188 & n13200;
  assign n13202 = ~n13199 & ~n13201;
  assign n13203 = ~n13191 & ~n13202;
  assign n13204 = ~n4115 & ~n13203;
  assign n13205 = ~n12547 & ~n12549;
  assign n13206 = ~n12948 & n13205;
  assign n13207 = ~n33361 & ~n13206;
  assign n13208 = ~n12549 & n33361;
  assign n13209 = ~n12547 & n13208;
  assign n13210 = n33361 & n13206;
  assign n13211 = ~n12948 & n13209;
  assign n13212 = ~n13207 & ~n33445;
  assign n13213 = n4115 & ~n13191;
  assign n13214 = n4115 & n13203;
  assign n13215 = ~n13202 & n13213;
  assign n13216 = ~n13212 & ~n33446;
  assign n13217 = ~n13204 & ~n13216;
  assign n13218 = ~n3754 & ~n13217;
  assign n13219 = n3754 & ~n13204;
  assign n13220 = ~n13216 & n13219;
  assign n13221 = ~n12564 & ~n33363;
  assign n13222 = ~n12564 & ~n12948;
  assign n13223 = ~n33363 & n13222;
  assign n13224 = ~n12948 & n13221;
  assign n13225 = n12572 & ~n33447;
  assign n13226 = n12576 & n13222;
  assign n13227 = ~n12564 & n12572;
  assign n13228 = ~n33363 & n13227;
  assign n13229 = ~n12948 & n13228;
  assign n13230 = ~n12572 & ~n33447;
  assign n13231 = ~n13229 & ~n13230;
  assign n13232 = ~n13225 & ~n13226;
  assign n13233 = ~n13220 & ~n33448;
  assign n13234 = ~n13218 & ~n13233;
  assign n13235 = ~n3444 & ~n13234;
  assign n13236 = ~n12578 & ~n12580;
  assign n13237 = ~n12948 & n13236;
  assign n13238 = ~n33365 & ~n13237;
  assign n13239 = ~n12580 & n33365;
  assign n13240 = ~n12578 & n13239;
  assign n13241 = n33365 & n13237;
  assign n13242 = ~n12948 & n13240;
  assign n13243 = ~n13238 & ~n33449;
  assign n13244 = n3444 & ~n13218;
  assign n13245 = n3444 & n13234;
  assign n13246 = ~n13233 & n13244;
  assign n13247 = ~n13243 & ~n33450;
  assign n13248 = ~n13235 & ~n13247;
  assign n13249 = ~n3116 & ~n13248;
  assign n13250 = n3116 & ~n13235;
  assign n13251 = ~n13247 & n13250;
  assign n13252 = ~n12595 & ~n33367;
  assign n13253 = ~n12595 & ~n12948;
  assign n13254 = ~n33367 & n13253;
  assign n13255 = ~n12948 & n13252;
  assign n13256 = n12603 & ~n33451;
  assign n13257 = n12607 & n13253;
  assign n13258 = ~n12595 & n12603;
  assign n13259 = ~n33367 & n13258;
  assign n13260 = ~n12948 & n13259;
  assign n13261 = ~n12603 & ~n33451;
  assign n13262 = ~n13260 & ~n13261;
  assign n13263 = ~n13256 & ~n13257;
  assign n13264 = ~n13251 & ~n33452;
  assign n13265 = ~n13249 & ~n13264;
  assign n13266 = ~n2833 & ~n13265;
  assign n13267 = ~n12609 & ~n12611;
  assign n13268 = ~n12948 & n13267;
  assign n13269 = ~n33369 & ~n13268;
  assign n13270 = ~n12611 & n33369;
  assign n13271 = ~n12609 & n13270;
  assign n13272 = n33369 & n13268;
  assign n13273 = ~n12948 & n13271;
  assign n13274 = ~n13269 & ~n33453;
  assign n13275 = n2833 & ~n13249;
  assign n13276 = n2833 & n13265;
  assign n13277 = ~n13264 & n13275;
  assign n13278 = ~n13274 & ~n33454;
  assign n13279 = ~n13266 & ~n13278;
  assign n13280 = ~n2536 & ~n13279;
  assign n13281 = ~n12626 & ~n33370;
  assign n13282 = ~n12948 & n13281;
  assign n13283 = ~n33372 & ~n13282;
  assign n13284 = ~n12626 & n33372;
  assign n13285 = ~n33370 & n13284;
  assign n13286 = n33372 & n13282;
  assign n13287 = ~n12948 & n13285;
  assign n13288 = ~n13283 & ~n33455;
  assign n13289 = n2536 & ~n13266;
  assign n13290 = ~n13278 & n13289;
  assign n13291 = ~n13288 & ~n13290;
  assign n13292 = ~n13280 & ~n13291;
  assign n13293 = ~n2283 & ~n13292;
  assign n13294 = ~n12644 & ~n12646;
  assign n13295 = ~n12948 & n13294;
  assign n13296 = ~n33374 & ~n13295;
  assign n13297 = ~n12646 & n33374;
  assign n13298 = ~n12644 & n13297;
  assign n13299 = n33374 & n13295;
  assign n13300 = ~n12948 & n13298;
  assign n13301 = ~n13296 & ~n33456;
  assign n13302 = n2283 & ~n13280;
  assign n13303 = n2283 & n13292;
  assign n13304 = ~n13291 & n13302;
  assign n13305 = ~n13301 & ~n33457;
  assign n13306 = ~n13293 & ~n13305;
  assign n13307 = ~n2021 & ~n13306;
  assign n13308 = n2021 & ~n13293;
  assign n13309 = ~n13305 & n13308;
  assign n13310 = ~n12661 & ~n33376;
  assign n13311 = ~n12661 & ~n12948;
  assign n13312 = ~n33376 & n13311;
  assign n13313 = ~n12948 & n13310;
  assign n13314 = n12669 & ~n33458;
  assign n13315 = n12673 & n13311;
  assign n13316 = ~n12661 & n12669;
  assign n13317 = ~n33376 & n13316;
  assign n13318 = ~n12948 & n13317;
  assign n13319 = ~n12669 & ~n33458;
  assign n13320 = ~n13318 & ~n13319;
  assign n13321 = ~n13314 & ~n13315;
  assign n13322 = ~n13309 & ~n33459;
  assign n13323 = ~n13307 & ~n13322;
  assign n13324 = ~n1796 & ~n13323;
  assign n13325 = ~n12675 & ~n12677;
  assign n13326 = ~n12948 & n13325;
  assign n13327 = ~n33378 & ~n13326;
  assign n13328 = ~n12677 & n33378;
  assign n13329 = ~n12675 & n13328;
  assign n13330 = n33378 & n13326;
  assign n13331 = ~n12948 & n13329;
  assign n13332 = ~n13327 & ~n33460;
  assign n13333 = n1796 & ~n13307;
  assign n13334 = n1796 & n13323;
  assign n13335 = ~n13322 & n13333;
  assign n13336 = ~n13332 & ~n33461;
  assign n13337 = ~n13324 & ~n13336;
  assign n13338 = ~n1567 & ~n13337;
  assign n13339 = ~n12692 & ~n33379;
  assign n13340 = ~n12948 & n13339;
  assign n13341 = ~n33381 & ~n13340;
  assign n13342 = ~n12692 & n33381;
  assign n13343 = ~n33379 & n13342;
  assign n13344 = n33381 & n13340;
  assign n13345 = ~n12948 & n13343;
  assign n13346 = ~n13341 & ~n33462;
  assign n13347 = n1567 & ~n13324;
  assign n13348 = ~n13336 & n13347;
  assign n13349 = ~n13346 & ~n13348;
  assign n13350 = ~n13338 & ~n13349;
  assign n13351 = ~n1374 & ~n13350;
  assign n13352 = ~n12710 & ~n12712;
  assign n13353 = ~n12948 & n13352;
  assign n13354 = ~n33383 & ~n13353;
  assign n13355 = ~n12712 & n33383;
  assign n13356 = ~n12710 & n13355;
  assign n13357 = n33383 & n13353;
  assign n13358 = ~n12948 & n13356;
  assign n13359 = ~n13354 & ~n33463;
  assign n13360 = n1374 & ~n13338;
  assign n13361 = n1374 & n13350;
  assign n13362 = ~n13349 & n13360;
  assign n13363 = ~n13359 & ~n33464;
  assign n13364 = ~n13351 & ~n13363;
  assign n13365 = ~n1179 & ~n13364;
  assign n13366 = n1179 & ~n13351;
  assign n13367 = ~n13363 & n13366;
  assign n13368 = ~n12727 & ~n33385;
  assign n13369 = ~n12727 & ~n12948;
  assign n13370 = ~n33385 & n13369;
  assign n13371 = ~n12948 & n13368;
  assign n13372 = n12735 & ~n33465;
  assign n13373 = n12739 & n13369;
  assign n13374 = ~n12727 & n12735;
  assign n13375 = ~n33385 & n13374;
  assign n13376 = ~n12948 & n13375;
  assign n13377 = ~n12735 & ~n33465;
  assign n13378 = ~n13376 & ~n13377;
  assign n13379 = ~n13372 & ~n13373;
  assign n13380 = ~n13367 & ~n33466;
  assign n13381 = ~n13365 & ~n13380;
  assign n13382 = ~n1016 & ~n13381;
  assign n13383 = ~n12741 & ~n12743;
  assign n13384 = ~n12948 & n13383;
  assign n13385 = ~n33387 & ~n13384;
  assign n13386 = ~n12743 & n33387;
  assign n13387 = ~n12741 & n13386;
  assign n13388 = n33387 & n13384;
  assign n13389 = ~n12948 & n13387;
  assign n13390 = ~n13385 & ~n33467;
  assign n13391 = n1016 & ~n13365;
  assign n13392 = n1016 & n13381;
  assign n13393 = ~n13380 & n13391;
  assign n13394 = ~n13390 & ~n33468;
  assign n13395 = ~n13382 & ~n13394;
  assign n13396 = ~n855 & ~n13395;
  assign n13397 = ~n12758 & ~n33388;
  assign n13398 = ~n12948 & n13397;
  assign n13399 = ~n33390 & ~n13398;
  assign n13400 = ~n12758 & n33390;
  assign n13401 = ~n33388 & n13400;
  assign n13402 = n33390 & n13398;
  assign n13403 = ~n12948 & n13401;
  assign n13404 = ~n13399 & ~n33469;
  assign n13405 = n855 & ~n13382;
  assign n13406 = ~n13394 & n13405;
  assign n13407 = ~n13404 & ~n13406;
  assign n13408 = ~n13396 & ~n13407;
  assign n13409 = ~n720 & ~n13408;
  assign n13410 = ~n12776 & ~n12778;
  assign n13411 = ~n12948 & n13410;
  assign n13412 = ~n33392 & ~n13411;
  assign n13413 = ~n12778 & n33392;
  assign n13414 = ~n12776 & n13413;
  assign n13415 = n33392 & n13411;
  assign n13416 = ~n12948 & n13414;
  assign n13417 = ~n13412 & ~n33470;
  assign n13418 = n720 & ~n13396;
  assign n13419 = n720 & n13408;
  assign n13420 = ~n13407 & n13418;
  assign n13421 = ~n13417 & ~n33471;
  assign n13422 = ~n13409 & ~n13421;
  assign n13423 = ~n592 & ~n13422;
  assign n13424 = n592 & ~n13409;
  assign n13425 = ~n13421 & n13424;
  assign n13426 = ~n12793 & ~n33394;
  assign n13427 = ~n12793 & ~n12948;
  assign n13428 = ~n33394 & n13427;
  assign n13429 = ~n12948 & n13426;
  assign n13430 = n12801 & ~n33472;
  assign n13431 = n12805 & n13427;
  assign n13432 = ~n12793 & n12801;
  assign n13433 = ~n33394 & n13432;
  assign n13434 = ~n12948 & n13433;
  assign n13435 = ~n12801 & ~n33472;
  assign n13436 = ~n13434 & ~n13435;
  assign n13437 = ~n13430 & ~n13431;
  assign n13438 = ~n13425 & ~n33473;
  assign n13439 = ~n13423 & ~n13438;
  assign n13440 = ~n487 & ~n13439;
  assign n13441 = ~n12807 & ~n12809;
  assign n13442 = ~n12948 & n13441;
  assign n13443 = ~n33396 & ~n13442;
  assign n13444 = ~n12809 & n33396;
  assign n13445 = ~n12807 & n13444;
  assign n13446 = n33396 & n13442;
  assign n13447 = ~n12948 & n13445;
  assign n13448 = ~n13443 & ~n33474;
  assign n13449 = n487 & ~n13423;
  assign n13450 = n487 & n13439;
  assign n13451 = ~n13438 & n13449;
  assign n13452 = ~n13448 & ~n33475;
  assign n13453 = ~n13440 & ~n13452;
  assign n13454 = ~n393 & ~n13453;
  assign n13455 = ~n12824 & ~n33397;
  assign n13456 = ~n12948 & n13455;
  assign n13457 = ~n33399 & ~n13456;
  assign n13458 = ~n12824 & n33399;
  assign n13459 = ~n33397 & n13458;
  assign n13460 = n33399 & n13456;
  assign n13461 = ~n12948 & n13459;
  assign n13462 = ~n13457 & ~n33476;
  assign n13463 = n393 & ~n13440;
  assign n13464 = ~n13452 & n13463;
  assign n13465 = ~n13462 & ~n13464;
  assign n13466 = ~n13454 & ~n13465;
  assign n13467 = ~n321 & ~n13466;
  assign n13468 = ~n12842 & ~n12844;
  assign n13469 = ~n12948 & n13468;
  assign n13470 = ~n33401 & ~n13469;
  assign n13471 = ~n12844 & n33401;
  assign n13472 = ~n12842 & n13471;
  assign n13473 = n33401 & n13469;
  assign n13474 = ~n12948 & n13472;
  assign n13475 = ~n13470 & ~n33477;
  assign n13476 = n321 & ~n13454;
  assign n13477 = n321 & n13466;
  assign n13478 = ~n13465 & n13476;
  assign n13479 = ~n13475 & ~n33478;
  assign n13480 = ~n13467 & ~n13479;
  assign n13481 = ~n263 & ~n13480;
  assign n13482 = n263 & ~n13467;
  assign n13483 = ~n13479 & n13482;
  assign n13484 = ~n12859 & ~n33403;
  assign n13485 = ~n12859 & ~n12948;
  assign n13486 = ~n33403 & n13485;
  assign n13487 = ~n12948 & n13484;
  assign n13488 = n12867 & ~n33479;
  assign n13489 = n12871 & n13485;
  assign n13490 = ~n12859 & n12867;
  assign n13491 = ~n33403 & n13490;
  assign n13492 = ~n12948 & n13491;
  assign n13493 = ~n12867 & ~n33479;
  assign n13494 = ~n13492 & ~n13493;
  assign n13495 = ~n13488 & ~n13489;
  assign n13496 = ~n13483 & ~n33480;
  assign n13497 = ~n13481 & ~n13496;
  assign n13498 = ~n214 & ~n13497;
  assign n13499 = ~n12873 & ~n12875;
  assign n13500 = ~n12948 & n13499;
  assign n13501 = ~n33405 & ~n13500;
  assign n13502 = ~n12875 & n33405;
  assign n13503 = ~n12873 & n13502;
  assign n13504 = n33405 & n13500;
  assign n13505 = ~n12948 & n13503;
  assign n13506 = ~n13501 & ~n33481;
  assign n13507 = n214 & ~n13481;
  assign n13508 = n214 & n13497;
  assign n13509 = ~n13496 & n13507;
  assign n13510 = ~n13506 & ~n33482;
  assign n13511 = ~n13498 & ~n13510;
  assign n13512 = ~n197 & ~n13511;
  assign n13513 = ~n12890 & ~n33406;
  assign n13514 = ~n12948 & n13513;
  assign n13515 = ~n33408 & ~n13514;
  assign n13516 = ~n12890 & n33408;
  assign n13517 = ~n33406 & n13516;
  assign n13518 = n33408 & n13514;
  assign n13519 = ~n12948 & n13517;
  assign n13520 = ~n13515 & ~n33483;
  assign n13521 = n197 & ~n13498;
  assign n13522 = ~n13510 & n13521;
  assign n13523 = ~n13520 & ~n13522;
  assign n13524 = ~n13512 & ~n13523;
  assign n13525 = ~n12908 & ~n12910;
  assign n13526 = ~n12948 & n13525;
  assign n13527 = ~n33410 & ~n13526;
  assign n13528 = ~n12910 & n33410;
  assign n13529 = ~n12908 & n13528;
  assign n13530 = n33410 & n13526;
  assign n13531 = ~n12948 & n13529;
  assign n13532 = ~n13527 & ~n33484;
  assign n13533 = ~n12924 & ~n12932;
  assign n13534 = ~n12932 & ~n12948;
  assign n13535 = ~n12924 & n13534;
  assign n13536 = ~n12948 & n13533;
  assign n13537 = ~n33413 & ~n33485;
  assign n13538 = ~n13532 & n13537;
  assign n13539 = ~n13524 & n13538;
  assign n13540 = n193 & ~n13539;
  assign n13541 = ~n13512 & n13532;
  assign n13542 = n13524 & n13532;
  assign n13543 = ~n13523 & n13541;
  assign n13544 = n12924 & ~n13534;
  assign n13545 = ~n193 & ~n13533;
  assign n13546 = ~n13544 & n13545;
  assign n13547 = ~n33486 & ~n13546;
  assign n13548 = ~n13540 & n13547;
  assign n13549 = pi44  & ~n13548;
  assign n13550 = ~pi42  & ~pi43 ;
  assign n13551 = ~pi44  & n13550;
  assign n13552 = ~n13549 & ~n13551;
  assign n13553 = ~n12948 & ~n13552;
  assign n13554 = ~pi44  & ~n13548;
  assign n13555 = pi45  & ~n13554;
  assign n13556 = ~pi45  & n13554;
  assign n13557 = n13026 & ~n13548;
  assign n13558 = ~n13555 & ~n33487;
  assign n13559 = ~n33324 & ~n33424;
  assign n13560 = ~n12275 & n13559;
  assign n13561 = ~n12294 & n13560;
  assign n13562 = ~n33326 & n13561;
  assign n13563 = n12280 & n12296;
  assign n13564 = ~n12288 & n13562;
  assign n13565 = ~n13551 & ~n33488;
  assign n13566 = ~n12946 & n13565;
  assign n13567 = ~n33413 & n13566;
  assign n13568 = ~n12940 & n13567;
  assign n13569 = n12948 & n13552;
  assign n13570 = ~n13549 & n13568;
  assign n13571 = n13558 & ~n33489;
  assign n13572 = ~n13553 & ~n13571;
  assign n13573 = ~n12296 & ~n13572;
  assign n13574 = n12296 & ~n13553;
  assign n13575 = ~n13571 & n13574;
  assign n13576 = ~n12948 & ~n13546;
  assign n13577 = ~n33486 & n13576;
  assign n13578 = ~n13540 & n13577;
  assign n13579 = ~n33487 & ~n13578;
  assign n13580 = pi46  & ~n13579;
  assign n13581 = ~pi46  & ~n13578;
  assign n13582 = ~pi46  & n13579;
  assign n13583 = ~n33487 & n13581;
  assign n13584 = ~n13580 & ~n33490;
  assign n13585 = ~n13575 & ~n13584;
  assign n13586 = ~n13573 & ~n13585;
  assign n13587 = ~n11719 & ~n13586;
  assign n13588 = n11719 & ~n13573;
  assign n13589 = ~n13585 & n13588;
  assign n13590 = n11719 & n13586;
  assign n13591 = ~n33425 & ~n13044;
  assign n13592 = ~n13548 & n13591;
  assign n13593 = n13042 & ~n13592;
  assign n13594 = ~n13042 & n13591;
  assign n13595 = ~n13042 & n13592;
  assign n13596 = ~n13548 & n13594;
  assign n13597 = ~n13593 & ~n33492;
  assign n13598 = ~n33491 & ~n13597;
  assign n13599 = ~n13587 & ~n13598;
  assign n13600 = ~n11097 & ~n13599;
  assign n13601 = n11097 & ~n13587;
  assign n13602 = ~n13598 & n13601;
  assign n13603 = ~n33426 & ~n13050;
  assign n13604 = ~n13050 & ~n13548;
  assign n13605 = ~n33426 & n13604;
  assign n13606 = ~n13548 & n13603;
  assign n13607 = n13024 & ~n33493;
  assign n13608 = n13049 & n13604;
  assign n13609 = n13024 & ~n33426;
  assign n13610 = ~n13050 & n13609;
  assign n13611 = ~n13548 & n13610;
  assign n13612 = ~n13024 & ~n33493;
  assign n13613 = ~n13611 & ~n13612;
  assign n13614 = ~n13607 & ~n13608;
  assign n13615 = ~n13602 & ~n33494;
  assign n13616 = ~n13600 & ~n13615;
  assign n13617 = ~n10555 & ~n13616;
  assign n13618 = n10555 & ~n13600;
  assign n13619 = ~n13615 & n13618;
  assign n13620 = n10555 & n13616;
  assign n13621 = ~n13052 & ~n13062;
  assign n13622 = ~n13548 & n13621;
  assign n13623 = ~n13059 & ~n13622;
  assign n13624 = n13059 & ~n13062;
  assign n13625 = ~n13052 & n13624;
  assign n13626 = n13059 & n13622;
  assign n13627 = ~n13548 & n13625;
  assign n13628 = n13059 & ~n13622;
  assign n13629 = ~n13059 & n13622;
  assign n13630 = ~n13628 & ~n13629;
  assign n13631 = ~n13623 & ~n33496;
  assign n13632 = ~n33495 & n33497;
  assign n13633 = ~n13617 & ~n13632;
  assign n13634 = ~n9969 & ~n13633;
  assign n13635 = n9969 & ~n13617;
  assign n13636 = ~n13632 & n13635;
  assign n13637 = ~n33428 & ~n13068;
  assign n13638 = ~n13068 & ~n13548;
  assign n13639 = ~n33428 & n13638;
  assign n13640 = ~n13548 & n13637;
  assign n13641 = n13012 & ~n33498;
  assign n13642 = n13067 & n13638;
  assign n13643 = n13012 & ~n33428;
  assign n13644 = ~n13068 & n13643;
  assign n13645 = ~n13548 & n13644;
  assign n13646 = ~n13012 & ~n33498;
  assign n13647 = ~n13645 & ~n13646;
  assign n13648 = ~n13641 & ~n13642;
  assign n13649 = ~n13636 & ~n33499;
  assign n13650 = ~n13634 & ~n13649;
  assign n13651 = ~n9457 & ~n13650;
  assign n13652 = n9457 & ~n13634;
  assign n13653 = ~n13649 & n13652;
  assign n13654 = n9457 & n13650;
  assign n13655 = ~n13070 & ~n13084;
  assign n13656 = ~n13548 & n13655;
  assign n13657 = ~n33430 & ~n13656;
  assign n13658 = n33430 & n13656;
  assign n13659 = ~n33430 & ~n13084;
  assign n13660 = ~n13070 & n13659;
  assign n13661 = ~n13548 & n13660;
  assign n13662 = n33430 & ~n13656;
  assign n13663 = ~n13661 & ~n13662;
  assign n13664 = ~n13657 & ~n13658;
  assign n13665 = ~n33500 & ~n33501;
  assign n13666 = ~n13651 & ~n13665;
  assign n13667 = ~n8896 & ~n13666;
  assign n13668 = n8896 & ~n13651;
  assign n13669 = ~n13665 & n13668;
  assign n13670 = ~n33431 & ~n13090;
  assign n13671 = ~n13090 & ~n13548;
  assign n13672 = ~n33431 & n13671;
  assign n13673 = ~n13548 & n13670;
  assign n13674 = n13004 & ~n33502;
  assign n13675 = n13089 & n13671;
  assign n13676 = n13004 & ~n33431;
  assign n13677 = ~n13090 & n13676;
  assign n13678 = ~n13548 & n13677;
  assign n13679 = ~n13004 & ~n33502;
  assign n13680 = ~n13678 & ~n13679;
  assign n13681 = ~n13674 & ~n13675;
  assign n13682 = ~n13669 & ~n33503;
  assign n13683 = ~n13667 & ~n13682;
  assign n13684 = ~n8411 & ~n13683;
  assign n13685 = n8411 & ~n13667;
  assign n13686 = ~n13682 & n13685;
  assign n13687 = n8411 & n13683;
  assign n13688 = ~n13092 & ~n13105;
  assign n13689 = ~n13548 & n13688;
  assign n13690 = ~n33432 & n13689;
  assign n13691 = n33432 & ~n13689;
  assign n13692 = n33432 & ~n13105;
  assign n13693 = ~n13092 & n13692;
  assign n13694 = ~n13548 & n13693;
  assign n13695 = ~n33432 & ~n13689;
  assign n13696 = ~n13694 & ~n13695;
  assign n13697 = ~n13690 & ~n13691;
  assign n13698 = ~n33504 & ~n33505;
  assign n13699 = ~n13684 & ~n13698;
  assign n13700 = ~n7885 & ~n13699;
  assign n13701 = n7885 & ~n13684;
  assign n13702 = ~n13698 & n13701;
  assign n13703 = ~n33433 & ~n13111;
  assign n13704 = ~n13111 & ~n13548;
  assign n13705 = ~n33433 & n13704;
  assign n13706 = ~n13548 & n13703;
  assign n13707 = n12996 & ~n33506;
  assign n13708 = n13110 & n13704;
  assign n13709 = n12996 & ~n33433;
  assign n13710 = ~n13111 & n13709;
  assign n13711 = ~n13548 & n13710;
  assign n13712 = ~n12996 & ~n33506;
  assign n13713 = ~n13711 & ~n13712;
  assign n13714 = ~n13707 & ~n13708;
  assign n13715 = ~n13702 & ~n33507;
  assign n13716 = ~n13700 & ~n13715;
  assign n13717 = ~n7428 & ~n13716;
  assign n13718 = n7428 & ~n13700;
  assign n13719 = ~n13715 & n13718;
  assign n13720 = n7428 & n13716;
  assign n13721 = ~n13113 & ~n13126;
  assign n13722 = ~n13548 & n13721;
  assign n13723 = ~n33434 & n13722;
  assign n13724 = n33434 & ~n13722;
  assign n13725 = ~n33434 & ~n13722;
  assign n13726 = n33434 & ~n13126;
  assign n13727 = ~n13113 & n13726;
  assign n13728 = n33434 & n13722;
  assign n13729 = ~n13548 & n13727;
  assign n13730 = ~n13725 & ~n33509;
  assign n13731 = ~n13723 & ~n13724;
  assign n13732 = ~n33508 & ~n33510;
  assign n13733 = ~n13717 & ~n13732;
  assign n13734 = ~n6937 & ~n13733;
  assign n13735 = n6937 & ~n13717;
  assign n13736 = ~n13732 & n13735;
  assign n13737 = ~n33435 & ~n13132;
  assign n13738 = ~n13132 & ~n13548;
  assign n13739 = ~n33435 & n13738;
  assign n13740 = ~n13548 & n13737;
  assign n13741 = n12988 & ~n33511;
  assign n13742 = n13131 & n13738;
  assign n13743 = n12988 & ~n33435;
  assign n13744 = ~n13132 & n13743;
  assign n13745 = ~n13548 & n13744;
  assign n13746 = ~n12988 & ~n33511;
  assign n13747 = ~n13745 & ~n13746;
  assign n13748 = ~n13741 & ~n13742;
  assign n13749 = ~n13736 & ~n33512;
  assign n13750 = ~n13734 & ~n13749;
  assign n13751 = ~n6507 & ~n13750;
  assign n13752 = n6507 & ~n13734;
  assign n13753 = ~n13749 & n13752;
  assign n13754 = n6507 & n13750;
  assign n13755 = ~n13134 & ~n13148;
  assign n13756 = ~n13148 & ~n13548;
  assign n13757 = ~n13134 & n13756;
  assign n13758 = ~n13548 & n13755;
  assign n13759 = n33437 & ~n33514;
  assign n13760 = n13146 & n13756;
  assign n13761 = ~n33437 & n33514;
  assign n13762 = n33437 & ~n13148;
  assign n13763 = ~n13134 & n13762;
  assign n13764 = ~n13548 & n13763;
  assign n13765 = ~n33437 & ~n33514;
  assign n13766 = ~n13764 & ~n13765;
  assign n13767 = ~n13759 & ~n33515;
  assign n13768 = ~n33513 & ~n33516;
  assign n13769 = ~n13751 & ~n13768;
  assign n13770 = ~n6051 & ~n13769;
  assign n13771 = n6051 & ~n13751;
  assign n13772 = ~n13768 & n13771;
  assign n13773 = ~n33438 & ~n13154;
  assign n13774 = ~n13154 & ~n13548;
  assign n13775 = ~n33438 & n13774;
  assign n13776 = ~n13548 & n13773;
  assign n13777 = n12980 & ~n33517;
  assign n13778 = n13153 & n13774;
  assign n13779 = n12980 & ~n33438;
  assign n13780 = ~n13154 & n13779;
  assign n13781 = ~n13548 & n13780;
  assign n13782 = ~n12980 & ~n33517;
  assign n13783 = ~n13781 & ~n13782;
  assign n13784 = ~n13777 & ~n13778;
  assign n13785 = ~n13772 & ~n33518;
  assign n13786 = ~n13770 & ~n13785;
  assign n13787 = ~n5648 & ~n13786;
  assign n13788 = ~n13156 & ~n13172;
  assign n13789 = ~n13548 & n13788;
  assign n13790 = ~n33441 & ~n13789;
  assign n13791 = n33441 & ~n13172;
  assign n13792 = ~n13156 & n13791;
  assign n13793 = n33441 & n13789;
  assign n13794 = ~n13548 & n13792;
  assign n13795 = ~n13790 & ~n33519;
  assign n13796 = n5648 & ~n13770;
  assign n13797 = ~n13785 & n13796;
  assign n13798 = n5648 & n13786;
  assign n13799 = ~n13795 & ~n33520;
  assign n13800 = ~n13787 & ~n13799;
  assign n13801 = ~n5223 & ~n13800;
  assign n13802 = n5223 & ~n13787;
  assign n13803 = ~n13799 & n13802;
  assign n13804 = ~n33442 & ~n13178;
  assign n13805 = ~n13178 & ~n13548;
  assign n13806 = ~n33442 & n13805;
  assign n13807 = ~n13548 & n13804;
  assign n13808 = n12972 & ~n33521;
  assign n13809 = n13177 & n13805;
  assign n13810 = n12972 & ~n33442;
  assign n13811 = ~n13178 & n13810;
  assign n13812 = ~n13548 & n13811;
  assign n13813 = ~n12972 & ~n33521;
  assign n13814 = ~n13812 & ~n13813;
  assign n13815 = ~n13808 & ~n13809;
  assign n13816 = ~n13803 & ~n33522;
  assign n13817 = ~n13801 & ~n13816;
  assign n13818 = ~n4851 & ~n13817;
  assign n13819 = n4851 & ~n13801;
  assign n13820 = ~n13816 & n13819;
  assign n13821 = n4851 & n13817;
  assign n13822 = ~n13180 & ~n13183;
  assign n13823 = ~n13183 & ~n13548;
  assign n13824 = ~n13180 & n13823;
  assign n13825 = ~n13548 & n13822;
  assign n13826 = n12964 & ~n33524;
  assign n13827 = n13181 & n13823;
  assign n13828 = n12964 & ~n13183;
  assign n13829 = ~n13180 & n13828;
  assign n13830 = ~n13548 & n13829;
  assign n13831 = ~n12964 & ~n33524;
  assign n13832 = ~n13830 & ~n13831;
  assign n13833 = ~n13826 & ~n13827;
  assign n13834 = ~n33523 & ~n33525;
  assign n13835 = ~n13818 & ~n13834;
  assign n13836 = ~n4461 & ~n13835;
  assign n13837 = n4461 & ~n13818;
  assign n13838 = ~n13834 & n13837;
  assign n13839 = n12956 & ~n33443;
  assign n13840 = ~n13189 & n13839;
  assign n13841 = ~n33443 & ~n13189;
  assign n13842 = ~n13548 & n13841;
  assign n13843 = n12956 & n13842;
  assign n13844 = ~n13548 & n13840;
  assign n13845 = ~n12956 & ~n13842;
  assign n13846 = ~n33526 & ~n13845;
  assign n13847 = ~n13838 & ~n13846;
  assign n13848 = ~n13836 & ~n13847;
  assign n13849 = ~n4115 & ~n13848;
  assign n13850 = ~n13191 & ~n13201;
  assign n13851 = ~n13548 & n13850;
  assign n13852 = ~n13199 & ~n13851;
  assign n13853 = ~n13191 & n13199;
  assign n13854 = ~n13201 & n13853;
  assign n13855 = n13199 & n13851;
  assign n13856 = ~n13548 & n13854;
  assign n13857 = ~n13852 & ~n33527;
  assign n13858 = n4115 & ~n13836;
  assign n13859 = ~n13847 & n13858;
  assign n13860 = n4115 & n13848;
  assign n13861 = ~n13857 & ~n33528;
  assign n13862 = ~n13849 & ~n13861;
  assign n13863 = ~n3754 & ~n13862;
  assign n13864 = n3754 & ~n13849;
  assign n13865 = ~n13861 & n13864;
  assign n13866 = ~n13204 & ~n33446;
  assign n13867 = ~n13204 & ~n13548;
  assign n13868 = ~n33446 & n13867;
  assign n13869 = ~n13548 & n13866;
  assign n13870 = n13212 & ~n33529;
  assign n13871 = n13216 & n13867;
  assign n13872 = n13212 & ~n33446;
  assign n13873 = ~n13204 & n13872;
  assign n13874 = ~n13548 & n13873;
  assign n13875 = ~n13212 & ~n33529;
  assign n13876 = ~n13874 & ~n13875;
  assign n13877 = ~n13870 & ~n13871;
  assign n13878 = ~n13865 & ~n33530;
  assign n13879 = ~n13863 & ~n13878;
  assign n13880 = ~n3444 & ~n13879;
  assign n13881 = ~n13218 & ~n13220;
  assign n13882 = ~n13548 & n13881;
  assign n13883 = ~n33448 & ~n13882;
  assign n13884 = ~n13218 & n33448;
  assign n13885 = ~n13220 & n13884;
  assign n13886 = n33448 & n13882;
  assign n13887 = ~n13548 & n13885;
  assign n13888 = ~n13883 & ~n33531;
  assign n13889 = n3444 & ~n13863;
  assign n13890 = ~n13878 & n13889;
  assign n13891 = n3444 & n13879;
  assign n13892 = ~n13888 & ~n33532;
  assign n13893 = ~n13880 & ~n13892;
  assign n13894 = ~n3116 & ~n13893;
  assign n13895 = n3116 & ~n13880;
  assign n13896 = ~n13892 & n13895;
  assign n13897 = ~n13235 & ~n33450;
  assign n13898 = ~n13235 & ~n13548;
  assign n13899 = ~n33450 & n13898;
  assign n13900 = ~n13548 & n13897;
  assign n13901 = n13243 & ~n33533;
  assign n13902 = n13247 & n13898;
  assign n13903 = n13243 & ~n33450;
  assign n13904 = ~n13235 & n13903;
  assign n13905 = ~n13548 & n13904;
  assign n13906 = ~n13243 & ~n33533;
  assign n13907 = ~n13905 & ~n13906;
  assign n13908 = ~n13901 & ~n13902;
  assign n13909 = ~n13896 & ~n33534;
  assign n13910 = ~n13894 & ~n13909;
  assign n13911 = ~n2833 & ~n13910;
  assign n13912 = ~n13249 & ~n13251;
  assign n13913 = ~n13548 & n13912;
  assign n13914 = ~n33452 & ~n13913;
  assign n13915 = ~n13249 & n33452;
  assign n13916 = ~n13251 & n13915;
  assign n13917 = n33452 & n13913;
  assign n13918 = ~n13548 & n13916;
  assign n13919 = ~n13914 & ~n33535;
  assign n13920 = n2833 & ~n13894;
  assign n13921 = ~n13909 & n13920;
  assign n13922 = n2833 & n13910;
  assign n13923 = ~n13919 & ~n33536;
  assign n13924 = ~n13911 & ~n13923;
  assign n13925 = ~n2536 & ~n13924;
  assign n13926 = n2536 & ~n13911;
  assign n13927 = ~n13923 & n13926;
  assign n13928 = ~n13266 & ~n33454;
  assign n13929 = ~n13266 & ~n13548;
  assign n13930 = ~n33454 & n13929;
  assign n13931 = ~n13548 & n13928;
  assign n13932 = n13274 & ~n33537;
  assign n13933 = n13278 & n13929;
  assign n13934 = n13274 & ~n33454;
  assign n13935 = ~n13266 & n13934;
  assign n13936 = ~n13548 & n13935;
  assign n13937 = ~n13274 & ~n33537;
  assign n13938 = ~n13936 & ~n13937;
  assign n13939 = ~n13932 & ~n13933;
  assign n13940 = ~n13927 & ~n33538;
  assign n13941 = ~n13925 & ~n13940;
  assign n13942 = ~n2283 & ~n13941;
  assign n13943 = n2283 & ~n13925;
  assign n13944 = ~n13940 & n13943;
  assign n13945 = n2283 & n13941;
  assign n13946 = ~n13280 & ~n13290;
  assign n13947 = ~n13280 & ~n13548;
  assign n13948 = ~n13290 & n13947;
  assign n13949 = ~n13548 & n13946;
  assign n13950 = n13288 & ~n33540;
  assign n13951 = n13291 & n13947;
  assign n13952 = ~n13280 & n13288;
  assign n13953 = ~n13290 & n13952;
  assign n13954 = ~n13548 & n13953;
  assign n13955 = ~n13288 & ~n33540;
  assign n13956 = ~n13954 & ~n13955;
  assign n13957 = ~n13950 & ~n13951;
  assign n13958 = ~n33539 & ~n33541;
  assign n13959 = ~n13942 & ~n13958;
  assign n13960 = ~n2021 & ~n13959;
  assign n13961 = n2021 & ~n13942;
  assign n13962 = ~n13958 & n13961;
  assign n13963 = ~n13293 & ~n33457;
  assign n13964 = ~n13293 & ~n13548;
  assign n13965 = ~n33457 & n13964;
  assign n13966 = ~n13548 & n13963;
  assign n13967 = n13301 & ~n33542;
  assign n13968 = n13305 & n13964;
  assign n13969 = n13301 & ~n33457;
  assign n13970 = ~n13293 & n13969;
  assign n13971 = ~n13548 & n13970;
  assign n13972 = ~n13301 & ~n33542;
  assign n13973 = ~n13971 & ~n13972;
  assign n13974 = ~n13967 & ~n13968;
  assign n13975 = ~n13962 & ~n33543;
  assign n13976 = ~n13960 & ~n13975;
  assign n13977 = ~n1796 & ~n13976;
  assign n13978 = ~n13307 & ~n13309;
  assign n13979 = ~n13548 & n13978;
  assign n13980 = ~n33459 & ~n13979;
  assign n13981 = ~n13307 & n33459;
  assign n13982 = ~n13309 & n13981;
  assign n13983 = n33459 & n13979;
  assign n13984 = ~n13548 & n13982;
  assign n13985 = ~n13980 & ~n33544;
  assign n13986 = n1796 & ~n13960;
  assign n13987 = ~n13975 & n13986;
  assign n13988 = n1796 & n13976;
  assign n13989 = ~n13985 & ~n33545;
  assign n13990 = ~n13977 & ~n13989;
  assign n13991 = ~n1567 & ~n13990;
  assign n13992 = n1567 & ~n13977;
  assign n13993 = ~n13989 & n13992;
  assign n13994 = ~n13324 & ~n33461;
  assign n13995 = ~n13324 & ~n13548;
  assign n13996 = ~n33461 & n13995;
  assign n13997 = ~n13548 & n13994;
  assign n13998 = n13332 & ~n33546;
  assign n13999 = n13336 & n13995;
  assign n14000 = n13332 & ~n33461;
  assign n14001 = ~n13324 & n14000;
  assign n14002 = ~n13548 & n14001;
  assign n14003 = ~n13332 & ~n33546;
  assign n14004 = ~n14002 & ~n14003;
  assign n14005 = ~n13998 & ~n13999;
  assign n14006 = ~n13993 & ~n33547;
  assign n14007 = ~n13991 & ~n14006;
  assign n14008 = ~n1374 & ~n14007;
  assign n14009 = n1374 & ~n13991;
  assign n14010 = ~n14006 & n14009;
  assign n14011 = n1374 & n14007;
  assign n14012 = ~n13338 & ~n13348;
  assign n14013 = ~n13338 & ~n13548;
  assign n14014 = ~n13348 & n14013;
  assign n14015 = ~n13548 & n14012;
  assign n14016 = n13346 & ~n33549;
  assign n14017 = n13349 & n14013;
  assign n14018 = ~n13338 & n13346;
  assign n14019 = ~n13348 & n14018;
  assign n14020 = ~n13548 & n14019;
  assign n14021 = ~n13346 & ~n33549;
  assign n14022 = ~n14020 & ~n14021;
  assign n14023 = ~n14016 & ~n14017;
  assign n14024 = ~n33548 & ~n33550;
  assign n14025 = ~n14008 & ~n14024;
  assign n14026 = ~n1179 & ~n14025;
  assign n14027 = n1179 & ~n14008;
  assign n14028 = ~n14024 & n14027;
  assign n14029 = ~n13351 & ~n33464;
  assign n14030 = ~n13351 & ~n13548;
  assign n14031 = ~n33464 & n14030;
  assign n14032 = ~n13548 & n14029;
  assign n14033 = n13359 & ~n33551;
  assign n14034 = n13363 & n14030;
  assign n14035 = n13359 & ~n33464;
  assign n14036 = ~n13351 & n14035;
  assign n14037 = ~n13548 & n14036;
  assign n14038 = ~n13359 & ~n33551;
  assign n14039 = ~n14037 & ~n14038;
  assign n14040 = ~n14033 & ~n14034;
  assign n14041 = ~n14028 & ~n33552;
  assign n14042 = ~n14026 & ~n14041;
  assign n14043 = ~n1016 & ~n14042;
  assign n14044 = ~n13365 & ~n13367;
  assign n14045 = ~n13548 & n14044;
  assign n14046 = ~n33466 & ~n14045;
  assign n14047 = ~n13365 & n33466;
  assign n14048 = ~n13367 & n14047;
  assign n14049 = n33466 & n14045;
  assign n14050 = ~n13548 & n14048;
  assign n14051 = ~n14046 & ~n33553;
  assign n14052 = n1016 & ~n14026;
  assign n14053 = ~n14041 & n14052;
  assign n14054 = n1016 & n14042;
  assign n14055 = ~n14051 & ~n33554;
  assign n14056 = ~n14043 & ~n14055;
  assign n14057 = ~n855 & ~n14056;
  assign n14058 = n855 & ~n14043;
  assign n14059 = ~n14055 & n14058;
  assign n14060 = ~n13382 & ~n33468;
  assign n14061 = ~n13382 & ~n13548;
  assign n14062 = ~n33468 & n14061;
  assign n14063 = ~n13548 & n14060;
  assign n14064 = n13390 & ~n33555;
  assign n14065 = n13394 & n14061;
  assign n14066 = n13390 & ~n33468;
  assign n14067 = ~n13382 & n14066;
  assign n14068 = ~n13548 & n14067;
  assign n14069 = ~n13390 & ~n33555;
  assign n14070 = ~n14068 & ~n14069;
  assign n14071 = ~n14064 & ~n14065;
  assign n14072 = ~n14059 & ~n33556;
  assign n14073 = ~n14057 & ~n14072;
  assign n14074 = ~n720 & ~n14073;
  assign n14075 = n720 & ~n14057;
  assign n14076 = ~n14072 & n14075;
  assign n14077 = n720 & n14073;
  assign n14078 = ~n13396 & ~n13406;
  assign n14079 = ~n13396 & ~n13548;
  assign n14080 = ~n13406 & n14079;
  assign n14081 = ~n13548 & n14078;
  assign n14082 = n13404 & ~n33558;
  assign n14083 = n13407 & n14079;
  assign n14084 = ~n13396 & n13404;
  assign n14085 = ~n13406 & n14084;
  assign n14086 = ~n13548 & n14085;
  assign n14087 = ~n13404 & ~n33558;
  assign n14088 = ~n14086 & ~n14087;
  assign n14089 = ~n14082 & ~n14083;
  assign n14090 = ~n33557 & ~n33559;
  assign n14091 = ~n14074 & ~n14090;
  assign n14092 = ~n592 & ~n14091;
  assign n14093 = n592 & ~n14074;
  assign n14094 = ~n14090 & n14093;
  assign n14095 = ~n13409 & ~n33471;
  assign n14096 = ~n13409 & ~n13548;
  assign n14097 = ~n33471 & n14096;
  assign n14098 = ~n13548 & n14095;
  assign n14099 = n13417 & ~n33560;
  assign n14100 = n13421 & n14096;
  assign n14101 = n13417 & ~n33471;
  assign n14102 = ~n13409 & n14101;
  assign n14103 = ~n13548 & n14102;
  assign n14104 = ~n13417 & ~n33560;
  assign n14105 = ~n14103 & ~n14104;
  assign n14106 = ~n14099 & ~n14100;
  assign n14107 = ~n14094 & ~n33561;
  assign n14108 = ~n14092 & ~n14107;
  assign n14109 = ~n487 & ~n14108;
  assign n14110 = ~n13423 & ~n13425;
  assign n14111 = ~n13548 & n14110;
  assign n14112 = ~n33473 & ~n14111;
  assign n14113 = ~n13423 & n33473;
  assign n14114 = ~n13425 & n14113;
  assign n14115 = n33473 & n14111;
  assign n14116 = ~n13548 & n14114;
  assign n14117 = ~n14112 & ~n33562;
  assign n14118 = n487 & ~n14092;
  assign n14119 = ~n14107 & n14118;
  assign n14120 = n487 & n14108;
  assign n14121 = ~n14117 & ~n33563;
  assign n14122 = ~n14109 & ~n14121;
  assign n14123 = ~n393 & ~n14122;
  assign n14124 = n393 & ~n14109;
  assign n14125 = ~n14121 & n14124;
  assign n14126 = ~n13440 & ~n33475;
  assign n14127 = ~n13440 & ~n13548;
  assign n14128 = ~n33475 & n14127;
  assign n14129 = ~n13548 & n14126;
  assign n14130 = n13448 & ~n33564;
  assign n14131 = n13452 & n14127;
  assign n14132 = n13448 & ~n33475;
  assign n14133 = ~n13440 & n14132;
  assign n14134 = ~n13548 & n14133;
  assign n14135 = ~n13448 & ~n33564;
  assign n14136 = ~n14134 & ~n14135;
  assign n14137 = ~n14130 & ~n14131;
  assign n14138 = ~n14125 & ~n33565;
  assign n14139 = ~n14123 & ~n14138;
  assign n14140 = ~n321 & ~n14139;
  assign n14141 = n321 & ~n14123;
  assign n14142 = ~n14138 & n14141;
  assign n14143 = n321 & n14139;
  assign n14144 = ~n13454 & ~n13464;
  assign n14145 = ~n13454 & ~n13548;
  assign n14146 = ~n13464 & n14145;
  assign n14147 = ~n13548 & n14144;
  assign n14148 = n13462 & ~n33567;
  assign n14149 = n13465 & n14145;
  assign n14150 = ~n13454 & n13462;
  assign n14151 = ~n13464 & n14150;
  assign n14152 = ~n13548 & n14151;
  assign n14153 = ~n13462 & ~n33567;
  assign n14154 = ~n14152 & ~n14153;
  assign n14155 = ~n14148 & ~n14149;
  assign n14156 = ~n33566 & ~n33568;
  assign n14157 = ~n14140 & ~n14156;
  assign n14158 = ~n263 & ~n14157;
  assign n14159 = n263 & ~n14140;
  assign n14160 = ~n14156 & n14159;
  assign n14161 = ~n13467 & ~n33478;
  assign n14162 = ~n13467 & ~n13548;
  assign n14163 = ~n33478 & n14162;
  assign n14164 = ~n13548 & n14161;
  assign n14165 = n13475 & ~n33569;
  assign n14166 = n13479 & n14162;
  assign n14167 = n13475 & ~n33478;
  assign n14168 = ~n13467 & n14167;
  assign n14169 = ~n13548 & n14168;
  assign n14170 = ~n13475 & ~n33569;
  assign n14171 = ~n14169 & ~n14170;
  assign n14172 = ~n14165 & ~n14166;
  assign n14173 = ~n14160 & ~n33570;
  assign n14174 = ~n14158 & ~n14173;
  assign n14175 = ~n214 & ~n14174;
  assign n14176 = ~n13481 & ~n13483;
  assign n14177 = ~n13548 & n14176;
  assign n14178 = ~n33480 & ~n14177;
  assign n14179 = ~n13481 & n33480;
  assign n14180 = ~n13483 & n14179;
  assign n14181 = n33480 & n14177;
  assign n14182 = ~n13548 & n14180;
  assign n14183 = ~n14178 & ~n33571;
  assign n14184 = n214 & ~n14158;
  assign n14185 = ~n14173 & n14184;
  assign n14186 = n214 & n14174;
  assign n14187 = ~n14183 & ~n33572;
  assign n14188 = ~n14175 & ~n14187;
  assign n14189 = ~n197 & ~n14188;
  assign n14190 = n197 & ~n14175;
  assign n14191 = ~n14187 & n14190;
  assign n14192 = ~n13498 & ~n33482;
  assign n14193 = ~n13498 & ~n13548;
  assign n14194 = ~n33482 & n14193;
  assign n14195 = ~n13548 & n14192;
  assign n14196 = n13506 & ~n33573;
  assign n14197 = n13510 & n14193;
  assign n14198 = n13506 & ~n33482;
  assign n14199 = ~n13498 & n14198;
  assign n14200 = ~n13548 & n14199;
  assign n14201 = ~n13506 & ~n33573;
  assign n14202 = ~n14200 & ~n14201;
  assign n14203 = ~n14196 & ~n14197;
  assign n14204 = ~n14191 & ~n33574;
  assign n14205 = ~n14189 & ~n14204;
  assign n14206 = ~n13512 & ~n13522;
  assign n14207 = ~n13512 & ~n13548;
  assign n14208 = ~n13522 & n14207;
  assign n14209 = ~n13548 & n14206;
  assign n14210 = n13520 & ~n33575;
  assign n14211 = n13523 & n14207;
  assign n14212 = ~n13512 & n13520;
  assign n14213 = ~n13522 & n14212;
  assign n14214 = ~n13548 & n14213;
  assign n14215 = ~n13520 & ~n33575;
  assign n14216 = ~n14214 & ~n14215;
  assign n14217 = ~n14210 & ~n14211;
  assign n14218 = ~n13524 & ~n13532;
  assign n14219 = ~n13532 & ~n13548;
  assign n14220 = ~n13524 & n14219;
  assign n14221 = ~n13548 & n14218;
  assign n14222 = ~n33486 & ~n33577;
  assign n14223 = ~n33576 & n14222;
  assign n14224 = ~n14205 & n14223;
  assign n14225 = n193 & ~n14224;
  assign n14226 = ~n14189 & n33576;
  assign n14227 = ~n14204 & n14226;
  assign n14228 = n14205 & n33576;
  assign n14229 = n13524 & ~n14219;
  assign n14230 = ~n193 & ~n14218;
  assign n14231 = ~n14229 & n14230;
  assign n14232 = ~n33578 & ~n14231;
  assign n14233 = ~n14225 & n14232;
  assign n14234 = ~n13836 & ~n13838;
  assign n14235 = ~n14233 & n14234;
  assign n14236 = ~n13846 & ~n14235;
  assign n14237 = ~n13838 & n13846;
  assign n14238 = ~n13836 & n14237;
  assign n14239 = n13846 & n14235;
  assign n14240 = ~n14233 & n14238;
  assign n14241 = ~n14236 & ~n33579;
  assign n14242 = ~n13818 & ~n33523;
  assign n14243 = ~n14233 & n14242;
  assign n14244 = ~n33525 & ~n14243;
  assign n14245 = ~n13818 & n33525;
  assign n14246 = ~n33523 & n14245;
  assign n14247 = n33525 & n14243;
  assign n14248 = ~n14233 & n14246;
  assign n14249 = ~n14244 & ~n33580;
  assign n14250 = ~n13801 & ~n13803;
  assign n14251 = ~n14233 & n14250;
  assign n14252 = ~n33522 & ~n14251;
  assign n14253 = ~n13803 & n33522;
  assign n14254 = ~n13801 & n14253;
  assign n14255 = n33522 & n14251;
  assign n14256 = ~n14233 & n14254;
  assign n14257 = ~n14252 & ~n33581;
  assign n14258 = ~n13770 & ~n13772;
  assign n14259 = ~n14233 & n14258;
  assign n14260 = ~n33518 & ~n14259;
  assign n14261 = ~n13772 & n33518;
  assign n14262 = ~n13770 & n14261;
  assign n14263 = n33518 & n14259;
  assign n14264 = ~n14233 & n14262;
  assign n14265 = ~n14260 & ~n33582;
  assign n14266 = ~n13751 & ~n33513;
  assign n14267 = ~n14233 & n14266;
  assign n14268 = ~n33516 & ~n14267;
  assign n14269 = ~n13751 & n33516;
  assign n14270 = ~n33513 & n14269;
  assign n14271 = n33516 & n14267;
  assign n14272 = ~n14233 & n14270;
  assign n14273 = ~n14268 & ~n33583;
  assign n14274 = ~n13734 & ~n13736;
  assign n14275 = ~n14233 & n14274;
  assign n14276 = ~n33512 & ~n14275;
  assign n14277 = ~n13736 & n33512;
  assign n14278 = ~n13734 & n14277;
  assign n14279 = n33512 & n14275;
  assign n14280 = ~n14233 & n14278;
  assign n14281 = ~n14276 & ~n33584;
  assign n14282 = ~n13700 & ~n13702;
  assign n14283 = ~n14233 & n14282;
  assign n14284 = ~n33507 & ~n14283;
  assign n14285 = ~n13702 & n33507;
  assign n14286 = ~n13700 & n14285;
  assign n14287 = n33507 & n14283;
  assign n14288 = ~n14233 & n14286;
  assign n14289 = ~n14284 & ~n33585;
  assign n14290 = ~n13667 & ~n13669;
  assign n14291 = ~n14233 & n14290;
  assign n14292 = ~n33503 & ~n14291;
  assign n14293 = ~n13669 & n33503;
  assign n14294 = ~n13667 & n14293;
  assign n14295 = n33503 & n14291;
  assign n14296 = ~n14233 & n14294;
  assign n14297 = ~n14292 & ~n33586;
  assign n14298 = ~n13634 & ~n13636;
  assign n14299 = ~n14233 & n14298;
  assign n14300 = ~n33499 & ~n14299;
  assign n14301 = ~n13636 & n33499;
  assign n14302 = ~n13634 & n14301;
  assign n14303 = n33499 & n14299;
  assign n14304 = ~n14233 & n14302;
  assign n14305 = ~n14300 & ~n33587;
  assign n14306 = ~n13600 & ~n13602;
  assign n14307 = ~n14233 & n14306;
  assign n14308 = ~n33494 & ~n14307;
  assign n14309 = ~n13602 & n33494;
  assign n14310 = ~n13600 & n14309;
  assign n14311 = n33494 & n14307;
  assign n14312 = ~n14233 & n14310;
  assign n14313 = ~n14308 & ~n33588;
  assign n14314 = ~n13573 & ~n13575;
  assign n14315 = ~n14233 & n14314;
  assign n14316 = ~n13584 & ~n14315;
  assign n14317 = ~n13575 & n13584;
  assign n14318 = ~n13573 & n14317;
  assign n14319 = n13584 & n14315;
  assign n14320 = ~n14233 & n14318;
  assign n14321 = ~n14316 & ~n33589;
  assign n14322 = ~pi42  & ~n14233;
  assign n14323 = ~pi43  & n14322;
  assign n14324 = n13550 & ~n14233;
  assign n14325 = ~n13548 & ~n14231;
  assign n14326 = ~n33578 & n14325;
  assign n14327 = ~n14225 & n14326;
  assign n14328 = ~n33590 & ~n14327;
  assign n14329 = pi44  & ~n14328;
  assign n14330 = ~pi44  & ~n14327;
  assign n14331 = ~pi44  & n14328;
  assign n14332 = ~n33590 & n14330;
  assign n14333 = ~n14329 & ~n33591;
  assign n14334 = pi42  & ~n14233;
  assign n14335 = ~pi40  & ~pi41 ;
  assign n14336 = ~pi42  & n14335;
  assign n14337 = ~n33411 & ~n33488;
  assign n14338 = ~n12927 & n14337;
  assign n14339 = ~n12946 & n14338;
  assign n14340 = ~n33413 & n14339;
  assign n14341 = n12932 & n12948;
  assign n14342 = ~n12940 & n14340;
  assign n14343 = ~n14336 & ~n33592;
  assign n14344 = ~n13546 & n14343;
  assign n14345 = ~n33486 & n14344;
  assign n14346 = ~n13540 & n14345;
  assign n14347 = ~n14334 & ~n14336;
  assign n14348 = n13548 & n14347;
  assign n14349 = ~n14334 & n14346;
  assign n14350 = pi43  & ~n14322;
  assign n14351 = ~n33590 & ~n14350;
  assign n14352 = ~n33593 & n14351;
  assign n14353 = ~n13548 & ~n14347;
  assign n14354 = n12948 & ~n14353;
  assign n14355 = ~n14352 & ~n14353;
  assign n14356 = n12948 & n14355;
  assign n14357 = ~n14352 & n14354;
  assign n14358 = ~n14333 & ~n33594;
  assign n14359 = ~n12948 & ~n14355;
  assign n14360 = n12296 & ~n14359;
  assign n14361 = ~n14358 & n14360;
  assign n14362 = ~n13553 & ~n33489;
  assign n14363 = ~n14233 & n14362;
  assign n14364 = n13558 & ~n14363;
  assign n14365 = ~n13558 & n14362;
  assign n14366 = ~n13558 & n14363;
  assign n14367 = ~n14233 & n14365;
  assign n14368 = ~n14364 & ~n33595;
  assign n14369 = ~n14361 & ~n14368;
  assign n14370 = ~n14358 & ~n14359;
  assign n14371 = ~n12296 & ~n14370;
  assign n14372 = n11719 & ~n14371;
  assign n14373 = ~n14369 & ~n14371;
  assign n14374 = n11719 & n14373;
  assign n14375 = ~n14369 & n14372;
  assign n14376 = ~n14321 & ~n33596;
  assign n14377 = ~n11719 & ~n14373;
  assign n14378 = n11097 & ~n14377;
  assign n14379 = ~n14376 & n14378;
  assign n14380 = ~n13587 & ~n33491;
  assign n14381 = ~n14233 & n14380;
  assign n14382 = ~n13597 & ~n14381;
  assign n14383 = ~n13587 & n13597;
  assign n14384 = ~n33491 & n14383;
  assign n14385 = n13597 & n14381;
  assign n14386 = ~n14233 & n14384;
  assign n14387 = n13597 & ~n14381;
  assign n14388 = ~n13597 & n14381;
  assign n14389 = ~n14387 & ~n14388;
  assign n14390 = ~n14382 & ~n33597;
  assign n14391 = ~n14379 & n33598;
  assign n14392 = ~n14376 & ~n14377;
  assign n14393 = ~n11097 & ~n14392;
  assign n14394 = n10555 & ~n14393;
  assign n14395 = ~n14391 & ~n14393;
  assign n14396 = n10555 & n14395;
  assign n14397 = ~n14391 & n14394;
  assign n14398 = ~n14313 & ~n33599;
  assign n14399 = ~n10555 & ~n14395;
  assign n14400 = n9969 & ~n14399;
  assign n14401 = ~n14398 & n14400;
  assign n14402 = ~n13617 & ~n33495;
  assign n14403 = ~n14233 & n14402;
  assign n14404 = ~n33497 & ~n14403;
  assign n14405 = n33497 & n14403;
  assign n14406 = ~n13617 & ~n33497;
  assign n14407 = ~n33495 & n14406;
  assign n14408 = ~n14233 & n14407;
  assign n14409 = n33497 & ~n14403;
  assign n14410 = ~n14408 & ~n14409;
  assign n14411 = ~n14404 & ~n14405;
  assign n14412 = ~n14401 & ~n33600;
  assign n14413 = ~n14398 & ~n14399;
  assign n14414 = ~n9969 & ~n14413;
  assign n14415 = n9457 & ~n14414;
  assign n14416 = ~n14412 & ~n14414;
  assign n14417 = n9457 & n14416;
  assign n14418 = ~n14412 & n14415;
  assign n14419 = ~n14305 & ~n33601;
  assign n14420 = ~n9457 & ~n14416;
  assign n14421 = n8896 & ~n14420;
  assign n14422 = ~n14419 & n14421;
  assign n14423 = ~n13651 & ~n33500;
  assign n14424 = ~n14233 & n14423;
  assign n14425 = ~n33501 & n14424;
  assign n14426 = n33501 & ~n14424;
  assign n14427 = ~n13651 & n33501;
  assign n14428 = ~n33500 & n14427;
  assign n14429 = ~n14233 & n14428;
  assign n14430 = ~n33501 & ~n14424;
  assign n14431 = ~n14429 & ~n14430;
  assign n14432 = ~n14425 & ~n14426;
  assign n14433 = ~n14422 & ~n33602;
  assign n14434 = ~n14419 & ~n14420;
  assign n14435 = ~n8896 & ~n14434;
  assign n14436 = n8411 & ~n14435;
  assign n14437 = ~n14433 & ~n14435;
  assign n14438 = n8411 & n14437;
  assign n14439 = ~n14433 & n14436;
  assign n14440 = ~n14297 & ~n33603;
  assign n14441 = ~n8411 & ~n14437;
  assign n14442 = n7885 & ~n14441;
  assign n14443 = ~n14440 & n14442;
  assign n14444 = ~n13684 & ~n33504;
  assign n14445 = ~n14233 & n14444;
  assign n14446 = ~n33505 & n14445;
  assign n14447 = n33505 & ~n14445;
  assign n14448 = ~n33505 & ~n14445;
  assign n14449 = ~n13684 & n33505;
  assign n14450 = ~n33504 & n14449;
  assign n14451 = n33505 & n14445;
  assign n14452 = ~n14233 & n14450;
  assign n14453 = ~n14448 & ~n33604;
  assign n14454 = ~n14446 & ~n14447;
  assign n14455 = ~n14443 & ~n33605;
  assign n14456 = ~n14440 & ~n14441;
  assign n14457 = ~n7885 & ~n14456;
  assign n14458 = n7428 & ~n14457;
  assign n14459 = ~n14455 & ~n14457;
  assign n14460 = n7428 & n14459;
  assign n14461 = ~n14455 & n14458;
  assign n14462 = ~n14289 & ~n33606;
  assign n14463 = ~n7428 & ~n14459;
  assign n14464 = n6937 & ~n14463;
  assign n14465 = ~n14462 & n14464;
  assign n14466 = ~n13717 & ~n33508;
  assign n14467 = ~n13717 & ~n14233;
  assign n14468 = ~n33508 & n14467;
  assign n14469 = ~n14233 & n14466;
  assign n14470 = n33510 & ~n33607;
  assign n14471 = n13732 & n14467;
  assign n14472 = ~n33510 & n33607;
  assign n14473 = ~n13717 & n33510;
  assign n14474 = ~n33508 & n14473;
  assign n14475 = ~n14233 & n14474;
  assign n14476 = ~n33510 & ~n33607;
  assign n14477 = ~n14475 & ~n14476;
  assign n14478 = ~n14470 & ~n33608;
  assign n14479 = ~n14465 & ~n33609;
  assign n14480 = ~n14462 & ~n14463;
  assign n14481 = ~n6937 & ~n14480;
  assign n14482 = n6507 & ~n14481;
  assign n14483 = ~n14479 & ~n14481;
  assign n14484 = n6507 & n14483;
  assign n14485 = ~n14479 & n14482;
  assign n14486 = ~n14281 & ~n33610;
  assign n14487 = ~n6507 & ~n14483;
  assign n14488 = n6051 & ~n14487;
  assign n14489 = ~n14486 & n14488;
  assign n14490 = ~n14273 & ~n14489;
  assign n14491 = ~n14486 & ~n14487;
  assign n14492 = ~n6051 & ~n14491;
  assign n14493 = n5648 & ~n14492;
  assign n14494 = ~n14490 & ~n14492;
  assign n14495 = n5648 & n14494;
  assign n14496 = ~n14490 & n14493;
  assign n14497 = ~n14265 & ~n33611;
  assign n14498 = ~n5648 & ~n14494;
  assign n14499 = n5223 & ~n14498;
  assign n14500 = ~n14497 & n14499;
  assign n14501 = ~n13787 & ~n33520;
  assign n14502 = ~n13787 & ~n14233;
  assign n14503 = ~n33520 & n14502;
  assign n14504 = ~n14233 & n14501;
  assign n14505 = n13795 & ~n33612;
  assign n14506 = n13799 & n14502;
  assign n14507 = ~n13787 & n13795;
  assign n14508 = ~n33520 & n14507;
  assign n14509 = ~n14233 & n14508;
  assign n14510 = ~n13795 & ~n33612;
  assign n14511 = ~n14509 & ~n14510;
  assign n14512 = ~n14505 & ~n14506;
  assign n14513 = ~n14500 & ~n33613;
  assign n14514 = ~n14497 & ~n14498;
  assign n14515 = ~n5223 & ~n14514;
  assign n14516 = n4851 & ~n14515;
  assign n14517 = ~n14513 & ~n14515;
  assign n14518 = n4851 & n14517;
  assign n14519 = ~n14513 & n14516;
  assign n14520 = ~n14257 & ~n33614;
  assign n14521 = ~n4851 & ~n14517;
  assign n14522 = n4461 & ~n14521;
  assign n14523 = ~n14520 & n14522;
  assign n14524 = ~n14249 & ~n14523;
  assign n14525 = ~n14520 & ~n14521;
  assign n14526 = ~n4461 & ~n14525;
  assign n14527 = n4115 & ~n14526;
  assign n14528 = ~n14524 & ~n14526;
  assign n14529 = n4115 & n14528;
  assign n14530 = ~n14524 & n14527;
  assign n14531 = ~n14241 & ~n33615;
  assign n14532 = ~n4115 & ~n14528;
  assign n14533 = ~n14531 & ~n14532;
  assign n14534 = ~n3754 & ~n14533;
  assign n14535 = ~n13849 & ~n33528;
  assign n14536 = ~n14233 & n14535;
  assign n14537 = n13857 & ~n14536;
  assign n14538 = ~n13857 & n14536;
  assign n14539 = ~n13849 & n13857;
  assign n14540 = ~n33528 & n14539;
  assign n14541 = ~n14233 & n14540;
  assign n14542 = ~n13857 & ~n14536;
  assign n14543 = ~n14541 & ~n14542;
  assign n14544 = ~n14537 & ~n14538;
  assign n14545 = n3754 & ~n14532;
  assign n14546 = ~n14531 & n14545;
  assign n14547 = ~n33616 & ~n14546;
  assign n14548 = ~n14534 & ~n14547;
  assign n14549 = ~n3444 & ~n14548;
  assign n14550 = ~n13863 & ~n13865;
  assign n14551 = ~n14233 & n14550;
  assign n14552 = ~n33530 & ~n14551;
  assign n14553 = ~n13865 & n33530;
  assign n14554 = ~n13863 & n14553;
  assign n14555 = n33530 & n14551;
  assign n14556 = ~n14233 & n14554;
  assign n14557 = ~n14552 & ~n33617;
  assign n14558 = n3444 & ~n14534;
  assign n14559 = n3444 & n14548;
  assign n14560 = ~n14547 & n14558;
  assign n14561 = ~n14557 & ~n33618;
  assign n14562 = ~n14549 & ~n14561;
  assign n14563 = ~n3116 & ~n14562;
  assign n14564 = n3116 & ~n14549;
  assign n14565 = ~n14561 & n14564;
  assign n14566 = ~n13880 & ~n33532;
  assign n14567 = ~n13880 & ~n14233;
  assign n14568 = ~n33532 & n14567;
  assign n14569 = ~n14233 & n14566;
  assign n14570 = n13888 & ~n33619;
  assign n14571 = n13892 & n14567;
  assign n14572 = ~n13880 & n13888;
  assign n14573 = ~n33532 & n14572;
  assign n14574 = ~n14233 & n14573;
  assign n14575 = ~n13888 & ~n33619;
  assign n14576 = ~n14574 & ~n14575;
  assign n14577 = ~n14570 & ~n14571;
  assign n14578 = ~n14565 & ~n33620;
  assign n14579 = ~n14563 & ~n14578;
  assign n14580 = ~n2833 & ~n14579;
  assign n14581 = ~n13894 & ~n13896;
  assign n14582 = ~n14233 & n14581;
  assign n14583 = ~n33534 & ~n14582;
  assign n14584 = ~n13896 & n33534;
  assign n14585 = ~n13894 & n14584;
  assign n14586 = n33534 & n14582;
  assign n14587 = ~n14233 & n14585;
  assign n14588 = ~n14583 & ~n33621;
  assign n14589 = n2833 & ~n14563;
  assign n14590 = n2833 & n14579;
  assign n14591 = ~n14578 & n14589;
  assign n14592 = ~n14588 & ~n33622;
  assign n14593 = ~n14580 & ~n14592;
  assign n14594 = ~n2536 & ~n14593;
  assign n14595 = n2536 & ~n14580;
  assign n14596 = ~n14592 & n14595;
  assign n14597 = ~n13911 & ~n33536;
  assign n14598 = ~n13911 & ~n14233;
  assign n14599 = ~n33536 & n14598;
  assign n14600 = ~n14233 & n14597;
  assign n14601 = n13919 & ~n33623;
  assign n14602 = n13923 & n14598;
  assign n14603 = ~n13911 & n13919;
  assign n14604 = ~n33536 & n14603;
  assign n14605 = ~n14233 & n14604;
  assign n14606 = ~n13919 & ~n33623;
  assign n14607 = ~n14605 & ~n14606;
  assign n14608 = ~n14601 & ~n14602;
  assign n14609 = ~n14596 & ~n33624;
  assign n14610 = ~n14594 & ~n14609;
  assign n14611 = ~n2283 & ~n14610;
  assign n14612 = ~n13925 & ~n13927;
  assign n14613 = ~n14233 & n14612;
  assign n14614 = ~n33538 & ~n14613;
  assign n14615 = ~n13927 & n33538;
  assign n14616 = ~n13925 & n14615;
  assign n14617 = n33538 & n14613;
  assign n14618 = ~n14233 & n14616;
  assign n14619 = ~n14614 & ~n33625;
  assign n14620 = n2283 & ~n14594;
  assign n14621 = n2283 & n14610;
  assign n14622 = ~n14609 & n14620;
  assign n14623 = ~n14619 & ~n33626;
  assign n14624 = ~n14611 & ~n14623;
  assign n14625 = ~n2021 & ~n14624;
  assign n14626 = ~n13942 & ~n33539;
  assign n14627 = ~n14233 & n14626;
  assign n14628 = ~n33541 & ~n14627;
  assign n14629 = ~n13942 & n33541;
  assign n14630 = ~n33539 & n14629;
  assign n14631 = n33541 & n14627;
  assign n14632 = ~n14233 & n14630;
  assign n14633 = ~n14628 & ~n33627;
  assign n14634 = n2021 & ~n14611;
  assign n14635 = ~n14623 & n14634;
  assign n14636 = ~n14633 & ~n14635;
  assign n14637 = ~n14625 & ~n14636;
  assign n14638 = ~n1796 & ~n14637;
  assign n14639 = ~n13960 & ~n13962;
  assign n14640 = ~n14233 & n14639;
  assign n14641 = ~n33543 & ~n14640;
  assign n14642 = ~n13962 & n33543;
  assign n14643 = ~n13960 & n14642;
  assign n14644 = n33543 & n14640;
  assign n14645 = ~n14233 & n14643;
  assign n14646 = ~n14641 & ~n33628;
  assign n14647 = n1796 & ~n14625;
  assign n14648 = n1796 & n14637;
  assign n14649 = ~n14636 & n14647;
  assign n14650 = ~n14646 & ~n33629;
  assign n14651 = ~n14638 & ~n14650;
  assign n14652 = ~n1567 & ~n14651;
  assign n14653 = n1567 & ~n14638;
  assign n14654 = ~n14650 & n14653;
  assign n14655 = ~n13977 & ~n33545;
  assign n14656 = ~n13977 & ~n14233;
  assign n14657 = ~n33545 & n14656;
  assign n14658 = ~n14233 & n14655;
  assign n14659 = n13985 & ~n33630;
  assign n14660 = n13989 & n14656;
  assign n14661 = ~n13977 & n13985;
  assign n14662 = ~n33545 & n14661;
  assign n14663 = ~n14233 & n14662;
  assign n14664 = ~n13985 & ~n33630;
  assign n14665 = ~n14663 & ~n14664;
  assign n14666 = ~n14659 & ~n14660;
  assign n14667 = ~n14654 & ~n33631;
  assign n14668 = ~n14652 & ~n14667;
  assign n14669 = ~n1374 & ~n14668;
  assign n14670 = ~n13991 & ~n13993;
  assign n14671 = ~n14233 & n14670;
  assign n14672 = ~n33547 & ~n14671;
  assign n14673 = ~n13993 & n33547;
  assign n14674 = ~n13991 & n14673;
  assign n14675 = n33547 & n14671;
  assign n14676 = ~n14233 & n14674;
  assign n14677 = ~n14672 & ~n33632;
  assign n14678 = n1374 & ~n14652;
  assign n14679 = n1374 & n14668;
  assign n14680 = ~n14667 & n14678;
  assign n14681 = ~n14677 & ~n33633;
  assign n14682 = ~n14669 & ~n14681;
  assign n14683 = ~n1179 & ~n14682;
  assign n14684 = ~n14008 & ~n33548;
  assign n14685 = ~n14233 & n14684;
  assign n14686 = ~n33550 & ~n14685;
  assign n14687 = ~n14008 & n33550;
  assign n14688 = ~n33548 & n14687;
  assign n14689 = n33550 & n14685;
  assign n14690 = ~n14233 & n14688;
  assign n14691 = ~n14686 & ~n33634;
  assign n14692 = n1179 & ~n14669;
  assign n14693 = ~n14681 & n14692;
  assign n14694 = ~n14691 & ~n14693;
  assign n14695 = ~n14683 & ~n14694;
  assign n14696 = ~n1016 & ~n14695;
  assign n14697 = ~n14026 & ~n14028;
  assign n14698 = ~n14233 & n14697;
  assign n14699 = ~n33552 & ~n14698;
  assign n14700 = ~n14028 & n33552;
  assign n14701 = ~n14026 & n14700;
  assign n14702 = n33552 & n14698;
  assign n14703 = ~n14233 & n14701;
  assign n14704 = ~n14699 & ~n33635;
  assign n14705 = n1016 & ~n14683;
  assign n14706 = n1016 & n14695;
  assign n14707 = ~n14694 & n14705;
  assign n14708 = ~n14704 & ~n33636;
  assign n14709 = ~n14696 & ~n14708;
  assign n14710 = ~n855 & ~n14709;
  assign n14711 = n855 & ~n14696;
  assign n14712 = ~n14708 & n14711;
  assign n14713 = ~n14043 & ~n33554;
  assign n14714 = ~n14043 & ~n14233;
  assign n14715 = ~n33554 & n14714;
  assign n14716 = ~n14233 & n14713;
  assign n14717 = n14051 & ~n33637;
  assign n14718 = n14055 & n14714;
  assign n14719 = ~n14043 & n14051;
  assign n14720 = ~n33554 & n14719;
  assign n14721 = ~n14233 & n14720;
  assign n14722 = ~n14051 & ~n33637;
  assign n14723 = ~n14721 & ~n14722;
  assign n14724 = ~n14717 & ~n14718;
  assign n14725 = ~n14712 & ~n33638;
  assign n14726 = ~n14710 & ~n14725;
  assign n14727 = ~n720 & ~n14726;
  assign n14728 = ~n14057 & ~n14059;
  assign n14729 = ~n14233 & n14728;
  assign n14730 = ~n33556 & ~n14729;
  assign n14731 = ~n14059 & n33556;
  assign n14732 = ~n14057 & n14731;
  assign n14733 = n33556 & n14729;
  assign n14734 = ~n14233 & n14732;
  assign n14735 = ~n14730 & ~n33639;
  assign n14736 = n720 & ~n14710;
  assign n14737 = n720 & n14726;
  assign n14738 = ~n14725 & n14736;
  assign n14739 = ~n14735 & ~n33640;
  assign n14740 = ~n14727 & ~n14739;
  assign n14741 = ~n592 & ~n14740;
  assign n14742 = ~n14074 & ~n33557;
  assign n14743 = ~n14233 & n14742;
  assign n14744 = ~n33559 & ~n14743;
  assign n14745 = ~n14074 & n33559;
  assign n14746 = ~n33557 & n14745;
  assign n14747 = n33559 & n14743;
  assign n14748 = ~n14233 & n14746;
  assign n14749 = ~n14744 & ~n33641;
  assign n14750 = n592 & ~n14727;
  assign n14751 = ~n14739 & n14750;
  assign n14752 = ~n14749 & ~n14751;
  assign n14753 = ~n14741 & ~n14752;
  assign n14754 = ~n487 & ~n14753;
  assign n14755 = ~n14092 & ~n14094;
  assign n14756 = ~n14233 & n14755;
  assign n14757 = ~n33561 & ~n14756;
  assign n14758 = ~n14094 & n33561;
  assign n14759 = ~n14092 & n14758;
  assign n14760 = n33561 & n14756;
  assign n14761 = ~n14233 & n14759;
  assign n14762 = ~n14757 & ~n33642;
  assign n14763 = n487 & ~n14741;
  assign n14764 = n487 & n14753;
  assign n14765 = ~n14752 & n14763;
  assign n14766 = ~n14762 & ~n33643;
  assign n14767 = ~n14754 & ~n14766;
  assign n14768 = ~n393 & ~n14767;
  assign n14769 = n393 & ~n14754;
  assign n14770 = ~n14766 & n14769;
  assign n14771 = ~n14109 & ~n33563;
  assign n14772 = ~n14109 & ~n14233;
  assign n14773 = ~n33563 & n14772;
  assign n14774 = ~n14233 & n14771;
  assign n14775 = n14117 & ~n33644;
  assign n14776 = n14121 & n14772;
  assign n14777 = ~n14109 & n14117;
  assign n14778 = ~n33563 & n14777;
  assign n14779 = ~n14233 & n14778;
  assign n14780 = ~n14117 & ~n33644;
  assign n14781 = ~n14779 & ~n14780;
  assign n14782 = ~n14775 & ~n14776;
  assign n14783 = ~n14770 & ~n33645;
  assign n14784 = ~n14768 & ~n14783;
  assign n14785 = ~n321 & ~n14784;
  assign n14786 = ~n14123 & ~n14125;
  assign n14787 = ~n14233 & n14786;
  assign n14788 = ~n33565 & ~n14787;
  assign n14789 = ~n14125 & n33565;
  assign n14790 = ~n14123 & n14789;
  assign n14791 = n33565 & n14787;
  assign n14792 = ~n14233 & n14790;
  assign n14793 = ~n14788 & ~n33646;
  assign n14794 = n321 & ~n14768;
  assign n14795 = n321 & n14784;
  assign n14796 = ~n14783 & n14794;
  assign n14797 = ~n14793 & ~n33647;
  assign n14798 = ~n14785 & ~n14797;
  assign n14799 = ~n263 & ~n14798;
  assign n14800 = ~n14140 & ~n33566;
  assign n14801 = ~n14233 & n14800;
  assign n14802 = ~n33568 & ~n14801;
  assign n14803 = ~n14140 & n33568;
  assign n14804 = ~n33566 & n14803;
  assign n14805 = n33568 & n14801;
  assign n14806 = ~n14233 & n14804;
  assign n14807 = ~n14802 & ~n33648;
  assign n14808 = n263 & ~n14785;
  assign n14809 = ~n14797 & n14808;
  assign n14810 = ~n14807 & ~n14809;
  assign n14811 = ~n14799 & ~n14810;
  assign n14812 = ~n214 & ~n14811;
  assign n14813 = ~n14158 & ~n14160;
  assign n14814 = ~n14233 & n14813;
  assign n14815 = ~n33570 & ~n14814;
  assign n14816 = ~n14160 & n33570;
  assign n14817 = ~n14158 & n14816;
  assign n14818 = n33570 & n14814;
  assign n14819 = ~n14233 & n14817;
  assign n14820 = ~n14815 & ~n33649;
  assign n14821 = n214 & ~n14799;
  assign n14822 = n214 & n14811;
  assign n14823 = ~n14810 & n14821;
  assign n14824 = ~n14820 & ~n33650;
  assign n14825 = ~n14812 & ~n14824;
  assign n14826 = ~n197 & ~n14825;
  assign n14827 = n197 & ~n14812;
  assign n14828 = ~n14824 & n14827;
  assign n14829 = ~n14175 & ~n33572;
  assign n14830 = ~n14175 & ~n14233;
  assign n14831 = ~n33572 & n14830;
  assign n14832 = ~n14233 & n14829;
  assign n14833 = n14183 & ~n33651;
  assign n14834 = n14187 & n14830;
  assign n14835 = ~n14175 & n14183;
  assign n14836 = ~n33572 & n14835;
  assign n14837 = ~n14233 & n14836;
  assign n14838 = ~n14183 & ~n33651;
  assign n14839 = ~n14837 & ~n14838;
  assign n14840 = ~n14833 & ~n14834;
  assign n14841 = ~n14828 & ~n33652;
  assign n14842 = ~n14826 & ~n14841;
  assign n14843 = ~n14189 & ~n14191;
  assign n14844 = ~n14233 & n14843;
  assign n14845 = ~n33574 & ~n14844;
  assign n14846 = ~n14191 & n33574;
  assign n14847 = ~n14189 & n14846;
  assign n14848 = n33574 & n14844;
  assign n14849 = ~n14233 & n14847;
  assign n14850 = ~n14845 & ~n33653;
  assign n14851 = ~n14205 & ~n33576;
  assign n14852 = ~n33576 & ~n14233;
  assign n14853 = ~n14205 & n14852;
  assign n14854 = ~n14233 & n14851;
  assign n14855 = ~n33578 & ~n33654;
  assign n14856 = ~n14850 & n14855;
  assign n14857 = ~n14842 & n14856;
  assign n14858 = n193 & ~n14857;
  assign n14859 = ~n14826 & n14850;
  assign n14860 = n14842 & n14850;
  assign n14861 = ~n14841 & n14859;
  assign n14862 = n14205 & ~n14852;
  assign n14863 = ~n193 & ~n14851;
  assign n14864 = ~n14862 & n14863;
  assign n14865 = ~n33655 & ~n14864;
  assign n14866 = ~n14858 & n14865;
  assign n14867 = pi40  & ~n14866;
  assign n14868 = ~pi38  & ~pi39 ;
  assign n14869 = ~pi40  & n14868;
  assign n14870 = ~n14867 & ~n14869;
  assign n14871 = ~n14233 & ~n14870;
  assign n14872 = ~pi40  & ~n14866;
  assign n14873 = pi41  & ~n14872;
  assign n14874 = ~pi41  & n14872;
  assign n14875 = n14335 & ~n14866;
  assign n14876 = ~n14873 & ~n33656;
  assign n14877 = ~n33484 & ~n33592;
  assign n14878 = ~n13527 & n14877;
  assign n14879 = ~n13546 & n14878;
  assign n14880 = ~n33486 & n14879;
  assign n14881 = n13532 & n13548;
  assign n14882 = ~n13540 & n14880;
  assign n14883 = ~n14869 & ~n33657;
  assign n14884 = ~n14231 & n14883;
  assign n14885 = ~n33578 & n14884;
  assign n14886 = ~n14225 & n14885;
  assign n14887 = n14233 & n14870;
  assign n14888 = ~n14867 & n14886;
  assign n14889 = n14876 & ~n33658;
  assign n14890 = ~n14871 & ~n14889;
  assign n14891 = ~n13548 & ~n14890;
  assign n14892 = n13548 & ~n14871;
  assign n14893 = ~n14889 & n14892;
  assign n14894 = ~n14233 & ~n14864;
  assign n14895 = ~n33655 & n14894;
  assign n14896 = ~n14858 & n14895;
  assign n14897 = ~n33656 & ~n14896;
  assign n14898 = pi42  & ~n14897;
  assign n14899 = ~pi42  & ~n14896;
  assign n14900 = ~pi42  & n14897;
  assign n14901 = ~n33656 & n14899;
  assign n14902 = ~n14898 & ~n33659;
  assign n14903 = ~n14893 & ~n14902;
  assign n14904 = ~n14891 & ~n14903;
  assign n14905 = ~n12948 & ~n14904;
  assign n14906 = n12948 & ~n14891;
  assign n14907 = ~n14903 & n14906;
  assign n14908 = n12948 & n14904;
  assign n14909 = ~n33593 & ~n14353;
  assign n14910 = ~n14866 & n14909;
  assign n14911 = n14351 & ~n14910;
  assign n14912 = ~n14351 & n14909;
  assign n14913 = ~n14351 & n14910;
  assign n14914 = ~n14866 & n14912;
  assign n14915 = ~n14911 & ~n33661;
  assign n14916 = ~n33660 & ~n14915;
  assign n14917 = ~n14905 & ~n14916;
  assign n14918 = ~n12296 & ~n14917;
  assign n14919 = n12296 & ~n14905;
  assign n14920 = ~n14916 & n14919;
  assign n14921 = ~n33594 & ~n14359;
  assign n14922 = ~n14359 & ~n14866;
  assign n14923 = ~n33594 & n14922;
  assign n14924 = ~n14866 & n14921;
  assign n14925 = n14333 & ~n33662;
  assign n14926 = n14358 & n14922;
  assign n14927 = n14333 & ~n33594;
  assign n14928 = ~n14359 & n14927;
  assign n14929 = ~n14866 & n14928;
  assign n14930 = ~n14333 & ~n33662;
  assign n14931 = ~n14929 & ~n14930;
  assign n14932 = ~n14925 & ~n14926;
  assign n14933 = ~n14920 & ~n33663;
  assign n14934 = ~n14918 & ~n14933;
  assign n14935 = ~n11719 & ~n14934;
  assign n14936 = n11719 & ~n14918;
  assign n14937 = ~n14933 & n14936;
  assign n14938 = n11719 & n14934;
  assign n14939 = ~n14361 & ~n14371;
  assign n14940 = ~n14866 & n14939;
  assign n14941 = ~n14368 & ~n14940;
  assign n14942 = n14368 & ~n14371;
  assign n14943 = ~n14361 & n14942;
  assign n14944 = n14368 & n14940;
  assign n14945 = ~n14866 & n14943;
  assign n14946 = n14368 & ~n14940;
  assign n14947 = ~n14368 & n14940;
  assign n14948 = ~n14946 & ~n14947;
  assign n14949 = ~n14941 & ~n33665;
  assign n14950 = ~n33664 & n33666;
  assign n14951 = ~n14935 & ~n14950;
  assign n14952 = ~n11097 & ~n14951;
  assign n14953 = n11097 & ~n14935;
  assign n14954 = ~n14950 & n14953;
  assign n14955 = ~n33596 & ~n14377;
  assign n14956 = ~n14377 & ~n14866;
  assign n14957 = ~n33596 & n14956;
  assign n14958 = ~n14866 & n14955;
  assign n14959 = n14321 & ~n33667;
  assign n14960 = n14376 & n14956;
  assign n14961 = n14321 & ~n33596;
  assign n14962 = ~n14377 & n14961;
  assign n14963 = ~n14866 & n14962;
  assign n14964 = ~n14321 & ~n33667;
  assign n14965 = ~n14963 & ~n14964;
  assign n14966 = ~n14959 & ~n14960;
  assign n14967 = ~n14954 & ~n33668;
  assign n14968 = ~n14952 & ~n14967;
  assign n14969 = ~n10555 & ~n14968;
  assign n14970 = n10555 & ~n14952;
  assign n14971 = ~n14967 & n14970;
  assign n14972 = n10555 & n14968;
  assign n14973 = ~n14379 & ~n14393;
  assign n14974 = ~n14866 & n14973;
  assign n14975 = ~n33598 & ~n14974;
  assign n14976 = n33598 & n14974;
  assign n14977 = ~n33598 & ~n14393;
  assign n14978 = ~n14379 & n14977;
  assign n14979 = ~n14866 & n14978;
  assign n14980 = n33598 & ~n14974;
  assign n14981 = ~n14979 & ~n14980;
  assign n14982 = ~n14975 & ~n14976;
  assign n14983 = ~n33669 & ~n33670;
  assign n14984 = ~n14969 & ~n14983;
  assign n14985 = ~n9969 & ~n14984;
  assign n14986 = n9969 & ~n14969;
  assign n14987 = ~n14983 & n14986;
  assign n14988 = ~n33599 & ~n14399;
  assign n14989 = ~n14399 & ~n14866;
  assign n14990 = ~n33599 & n14989;
  assign n14991 = ~n14866 & n14988;
  assign n14992 = n14313 & ~n33671;
  assign n14993 = n14398 & n14989;
  assign n14994 = n14313 & ~n33599;
  assign n14995 = ~n14399 & n14994;
  assign n14996 = ~n14866 & n14995;
  assign n14997 = ~n14313 & ~n33671;
  assign n14998 = ~n14996 & ~n14997;
  assign n14999 = ~n14992 & ~n14993;
  assign n15000 = ~n14987 & ~n33672;
  assign n15001 = ~n14985 & ~n15000;
  assign n15002 = ~n9457 & ~n15001;
  assign n15003 = n9457 & ~n14985;
  assign n15004 = ~n15000 & n15003;
  assign n15005 = n9457 & n15001;
  assign n15006 = ~n14401 & ~n14414;
  assign n15007 = ~n14866 & n15006;
  assign n15008 = ~n33600 & n15007;
  assign n15009 = n33600 & ~n15007;
  assign n15010 = n33600 & ~n14414;
  assign n15011 = ~n14401 & n15010;
  assign n15012 = ~n14866 & n15011;
  assign n15013 = ~n33600 & ~n15007;
  assign n15014 = ~n15012 & ~n15013;
  assign n15015 = ~n15008 & ~n15009;
  assign n15016 = ~n33673 & ~n33674;
  assign n15017 = ~n15002 & ~n15016;
  assign n15018 = ~n8896 & ~n15017;
  assign n15019 = n8896 & ~n15002;
  assign n15020 = ~n15016 & n15019;
  assign n15021 = ~n33601 & ~n14420;
  assign n15022 = ~n14420 & ~n14866;
  assign n15023 = ~n33601 & n15022;
  assign n15024 = ~n14866 & n15021;
  assign n15025 = n14305 & ~n33675;
  assign n15026 = n14419 & n15022;
  assign n15027 = n14305 & ~n33601;
  assign n15028 = ~n14420 & n15027;
  assign n15029 = ~n14866 & n15028;
  assign n15030 = ~n14305 & ~n33675;
  assign n15031 = ~n15029 & ~n15030;
  assign n15032 = ~n15025 & ~n15026;
  assign n15033 = ~n15020 & ~n33676;
  assign n15034 = ~n15018 & ~n15033;
  assign n15035 = ~n8411 & ~n15034;
  assign n15036 = n8411 & ~n15018;
  assign n15037 = ~n15033 & n15036;
  assign n15038 = n8411 & n15034;
  assign n15039 = ~n14422 & ~n14435;
  assign n15040 = ~n14866 & n15039;
  assign n15041 = ~n33602 & n15040;
  assign n15042 = n33602 & ~n15040;
  assign n15043 = ~n33602 & ~n15040;
  assign n15044 = n33602 & ~n14435;
  assign n15045 = ~n14422 & n15044;
  assign n15046 = n33602 & n15040;
  assign n15047 = ~n14866 & n15045;
  assign n15048 = ~n15043 & ~n33678;
  assign n15049 = ~n15041 & ~n15042;
  assign n15050 = ~n33677 & ~n33679;
  assign n15051 = ~n15035 & ~n15050;
  assign n15052 = ~n7885 & ~n15051;
  assign n15053 = n7885 & ~n15035;
  assign n15054 = ~n15050 & n15053;
  assign n15055 = ~n33603 & ~n14441;
  assign n15056 = ~n14441 & ~n14866;
  assign n15057 = ~n33603 & n15056;
  assign n15058 = ~n14866 & n15055;
  assign n15059 = n14297 & ~n33680;
  assign n15060 = n14440 & n15056;
  assign n15061 = n14297 & ~n33603;
  assign n15062 = ~n14441 & n15061;
  assign n15063 = ~n14866 & n15062;
  assign n15064 = ~n14297 & ~n33680;
  assign n15065 = ~n15063 & ~n15064;
  assign n15066 = ~n15059 & ~n15060;
  assign n15067 = ~n15054 & ~n33681;
  assign n15068 = ~n15052 & ~n15067;
  assign n15069 = ~n7428 & ~n15068;
  assign n15070 = n7428 & ~n15052;
  assign n15071 = ~n15067 & n15070;
  assign n15072 = n7428 & n15068;
  assign n15073 = ~n14443 & ~n14457;
  assign n15074 = ~n14457 & ~n14866;
  assign n15075 = ~n14443 & n15074;
  assign n15076 = ~n14866 & n15073;
  assign n15077 = n33605 & ~n33683;
  assign n15078 = n14455 & n15074;
  assign n15079 = ~n33605 & n33683;
  assign n15080 = n33605 & ~n14457;
  assign n15081 = ~n14443 & n15080;
  assign n15082 = ~n14866 & n15081;
  assign n15083 = ~n33605 & ~n33683;
  assign n15084 = ~n15082 & ~n15083;
  assign n15085 = ~n15077 & ~n33684;
  assign n15086 = ~n33682 & ~n33685;
  assign n15087 = ~n15069 & ~n15086;
  assign n15088 = ~n6937 & ~n15087;
  assign n15089 = n6937 & ~n15069;
  assign n15090 = ~n15086 & n15089;
  assign n15091 = ~n33606 & ~n14463;
  assign n15092 = ~n14463 & ~n14866;
  assign n15093 = ~n33606 & n15092;
  assign n15094 = ~n14866 & n15091;
  assign n15095 = n14289 & ~n33686;
  assign n15096 = n14462 & n15092;
  assign n15097 = n14289 & ~n33606;
  assign n15098 = ~n14463 & n15097;
  assign n15099 = ~n14866 & n15098;
  assign n15100 = ~n14289 & ~n33686;
  assign n15101 = ~n15099 & ~n15100;
  assign n15102 = ~n15095 & ~n15096;
  assign n15103 = ~n15090 & ~n33687;
  assign n15104 = ~n15088 & ~n15103;
  assign n15105 = ~n6507 & ~n15104;
  assign n15106 = ~n14465 & ~n14481;
  assign n15107 = ~n14866 & n15106;
  assign n15108 = ~n33609 & ~n15107;
  assign n15109 = n33609 & ~n14481;
  assign n15110 = ~n14465 & n15109;
  assign n15111 = n33609 & n15107;
  assign n15112 = ~n14866 & n15110;
  assign n15113 = ~n15108 & ~n33688;
  assign n15114 = n6507 & ~n15088;
  assign n15115 = ~n15103 & n15114;
  assign n15116 = n6507 & n15104;
  assign n15117 = ~n15113 & ~n33689;
  assign n15118 = ~n15105 & ~n15117;
  assign n15119 = ~n6051 & ~n15118;
  assign n15120 = n6051 & ~n15105;
  assign n15121 = ~n15117 & n15120;
  assign n15122 = ~n33610 & ~n14487;
  assign n15123 = ~n14487 & ~n14866;
  assign n15124 = ~n33610 & n15123;
  assign n15125 = ~n14866 & n15122;
  assign n15126 = n14281 & ~n33690;
  assign n15127 = n14486 & n15123;
  assign n15128 = n14281 & ~n33610;
  assign n15129 = ~n14487 & n15128;
  assign n15130 = ~n14866 & n15129;
  assign n15131 = ~n14281 & ~n33690;
  assign n15132 = ~n15130 & ~n15131;
  assign n15133 = ~n15126 & ~n15127;
  assign n15134 = ~n15121 & ~n33691;
  assign n15135 = ~n15119 & ~n15134;
  assign n15136 = ~n5648 & ~n15135;
  assign n15137 = n5648 & ~n15119;
  assign n15138 = ~n15134 & n15137;
  assign n15139 = n5648 & n15135;
  assign n15140 = ~n14489 & ~n14492;
  assign n15141 = ~n14492 & ~n14866;
  assign n15142 = ~n14489 & n15141;
  assign n15143 = ~n14866 & n15140;
  assign n15144 = n14273 & ~n33693;
  assign n15145 = n14490 & n15141;
  assign n15146 = n14273 & ~n14492;
  assign n15147 = ~n14489 & n15146;
  assign n15148 = ~n14866 & n15147;
  assign n15149 = ~n14273 & ~n33693;
  assign n15150 = ~n15148 & ~n15149;
  assign n15151 = ~n15144 & ~n15145;
  assign n15152 = ~n33692 & ~n33694;
  assign n15153 = ~n15136 & ~n15152;
  assign n15154 = ~n5223 & ~n15153;
  assign n15155 = n5223 & ~n15136;
  assign n15156 = ~n15152 & n15155;
  assign n15157 = ~n33611 & ~n14498;
  assign n15158 = ~n14498 & ~n14866;
  assign n15159 = ~n33611 & n15158;
  assign n15160 = ~n14866 & n15157;
  assign n15161 = n14265 & ~n33695;
  assign n15162 = n14497 & n15158;
  assign n15163 = n14265 & ~n33611;
  assign n15164 = ~n14498 & n15163;
  assign n15165 = ~n14866 & n15164;
  assign n15166 = ~n14265 & ~n33695;
  assign n15167 = ~n15165 & ~n15166;
  assign n15168 = ~n15161 & ~n15162;
  assign n15169 = ~n15156 & ~n33696;
  assign n15170 = ~n15154 & ~n15169;
  assign n15171 = ~n4851 & ~n15170;
  assign n15172 = ~n14500 & ~n14515;
  assign n15173 = ~n14866 & n15172;
  assign n15174 = ~n33613 & ~n15173;
  assign n15175 = n33613 & ~n14515;
  assign n15176 = ~n14500 & n15175;
  assign n15177 = n33613 & n15173;
  assign n15178 = ~n14866 & n15176;
  assign n15179 = ~n15174 & ~n33697;
  assign n15180 = n4851 & ~n15154;
  assign n15181 = ~n15169 & n15180;
  assign n15182 = n4851 & n15170;
  assign n15183 = ~n15179 & ~n33698;
  assign n15184 = ~n15171 & ~n15183;
  assign n15185 = ~n4461 & ~n15184;
  assign n15186 = n4461 & ~n15171;
  assign n15187 = ~n15183 & n15186;
  assign n15188 = ~n33614 & ~n14521;
  assign n15189 = ~n14521 & ~n14866;
  assign n15190 = ~n33614 & n15189;
  assign n15191 = ~n14866 & n15188;
  assign n15192 = n14257 & ~n33699;
  assign n15193 = n14520 & n15189;
  assign n15194 = n14257 & ~n33614;
  assign n15195 = ~n14521 & n15194;
  assign n15196 = ~n14866 & n15195;
  assign n15197 = ~n14257 & ~n33699;
  assign n15198 = ~n15196 & ~n15197;
  assign n15199 = ~n15192 & ~n15193;
  assign n15200 = ~n15187 & ~n33700;
  assign n15201 = ~n15185 & ~n15200;
  assign n15202 = ~n4115 & ~n15201;
  assign n15203 = n4115 & ~n15185;
  assign n15204 = ~n15200 & n15203;
  assign n15205 = n4115 & n15201;
  assign n15206 = ~n14523 & ~n14526;
  assign n15207 = ~n14526 & ~n14866;
  assign n15208 = ~n14523 & n15207;
  assign n15209 = ~n14866 & n15206;
  assign n15210 = n14249 & ~n33702;
  assign n15211 = n14524 & n15207;
  assign n15212 = n14249 & ~n14526;
  assign n15213 = ~n14523 & n15212;
  assign n15214 = ~n14866 & n15213;
  assign n15215 = ~n14249 & ~n33702;
  assign n15216 = ~n15214 & ~n15215;
  assign n15217 = ~n15210 & ~n15211;
  assign n15218 = ~n33701 & ~n33703;
  assign n15219 = ~n15202 & ~n15218;
  assign n15220 = ~n3754 & ~n15219;
  assign n15221 = n3754 & ~n15202;
  assign n15222 = ~n15218 & n15221;
  assign n15223 = ~n33615 & ~n14532;
  assign n15224 = ~n14866 & n15223;
  assign n15225 = n14241 & ~n15224;
  assign n15226 = ~n14241 & n15224;
  assign n15227 = n14241 & ~n33615;
  assign n15228 = ~n14532 & n15227;
  assign n15229 = ~n14866 & n15228;
  assign n15230 = ~n14241 & ~n15224;
  assign n15231 = ~n15229 & ~n15230;
  assign n15232 = ~n15225 & ~n15226;
  assign n15233 = ~n15222 & ~n33704;
  assign n15234 = ~n15220 & ~n15233;
  assign n15235 = ~n3444 & ~n15234;
  assign n15236 = ~n14534 & ~n14546;
  assign n15237 = ~n14866 & n15236;
  assign n15238 = ~n33616 & n15237;
  assign n15239 = n33616 & ~n15237;
  assign n15240 = ~n14534 & n33616;
  assign n15241 = ~n14546 & n15240;
  assign n15242 = ~n14866 & n15241;
  assign n15243 = ~n33616 & ~n15237;
  assign n15244 = ~n15242 & ~n15243;
  assign n15245 = ~n15238 & ~n15239;
  assign n15246 = n3444 & ~n15220;
  assign n15247 = ~n15233 & n15246;
  assign n15248 = n3444 & n15234;
  assign n15249 = ~n33705 & ~n33706;
  assign n15250 = ~n15235 & ~n15249;
  assign n15251 = ~n3116 & ~n15250;
  assign n15252 = n3116 & ~n15235;
  assign n15253 = ~n15249 & n15252;
  assign n15254 = ~n14549 & ~n33618;
  assign n15255 = ~n14549 & ~n14866;
  assign n15256 = ~n33618 & n15255;
  assign n15257 = ~n14866 & n15254;
  assign n15258 = n14557 & ~n33707;
  assign n15259 = n14561 & n15255;
  assign n15260 = n14557 & ~n33618;
  assign n15261 = ~n14549 & n15260;
  assign n15262 = ~n14866 & n15261;
  assign n15263 = ~n14557 & ~n33707;
  assign n15264 = ~n15262 & ~n15263;
  assign n15265 = ~n15258 & ~n15259;
  assign n15266 = ~n15253 & ~n33708;
  assign n15267 = ~n15251 & ~n15266;
  assign n15268 = ~n2833 & ~n15267;
  assign n15269 = ~n14563 & ~n14565;
  assign n15270 = ~n14866 & n15269;
  assign n15271 = ~n33620 & ~n15270;
  assign n15272 = ~n14563 & n33620;
  assign n15273 = ~n14565 & n15272;
  assign n15274 = n33620 & n15270;
  assign n15275 = ~n14866 & n15273;
  assign n15276 = ~n15271 & ~n33709;
  assign n15277 = n2833 & ~n15251;
  assign n15278 = ~n15266 & n15277;
  assign n15279 = n2833 & n15267;
  assign n15280 = ~n15276 & ~n33710;
  assign n15281 = ~n15268 & ~n15280;
  assign n15282 = ~n2536 & ~n15281;
  assign n15283 = n2536 & ~n15268;
  assign n15284 = ~n15280 & n15283;
  assign n15285 = ~n14580 & ~n33622;
  assign n15286 = ~n14580 & ~n14866;
  assign n15287 = ~n33622 & n15286;
  assign n15288 = ~n14866 & n15285;
  assign n15289 = n14588 & ~n33711;
  assign n15290 = n14592 & n15286;
  assign n15291 = n14588 & ~n33622;
  assign n15292 = ~n14580 & n15291;
  assign n15293 = ~n14866 & n15292;
  assign n15294 = ~n14588 & ~n33711;
  assign n15295 = ~n15293 & ~n15294;
  assign n15296 = ~n15289 & ~n15290;
  assign n15297 = ~n15284 & ~n33712;
  assign n15298 = ~n15282 & ~n15297;
  assign n15299 = ~n2283 & ~n15298;
  assign n15300 = ~n14594 & ~n14596;
  assign n15301 = ~n14866 & n15300;
  assign n15302 = ~n33624 & ~n15301;
  assign n15303 = ~n14594 & n33624;
  assign n15304 = ~n14596 & n15303;
  assign n15305 = n33624 & n15301;
  assign n15306 = ~n14866 & n15304;
  assign n15307 = ~n15302 & ~n33713;
  assign n15308 = n2283 & ~n15282;
  assign n15309 = ~n15297 & n15308;
  assign n15310 = n2283 & n15298;
  assign n15311 = ~n15307 & ~n33714;
  assign n15312 = ~n15299 & ~n15311;
  assign n15313 = ~n2021 & ~n15312;
  assign n15314 = n2021 & ~n15299;
  assign n15315 = ~n15311 & n15314;
  assign n15316 = ~n14611 & ~n33626;
  assign n15317 = ~n14611 & ~n14866;
  assign n15318 = ~n33626 & n15317;
  assign n15319 = ~n14866 & n15316;
  assign n15320 = n14619 & ~n33715;
  assign n15321 = n14623 & n15317;
  assign n15322 = n14619 & ~n33626;
  assign n15323 = ~n14611 & n15322;
  assign n15324 = ~n14866 & n15323;
  assign n15325 = ~n14619 & ~n33715;
  assign n15326 = ~n15324 & ~n15325;
  assign n15327 = ~n15320 & ~n15321;
  assign n15328 = ~n15315 & ~n33716;
  assign n15329 = ~n15313 & ~n15328;
  assign n15330 = ~n1796 & ~n15329;
  assign n15331 = n1796 & ~n15313;
  assign n15332 = ~n15328 & n15331;
  assign n15333 = n1796 & n15329;
  assign n15334 = ~n14625 & ~n14635;
  assign n15335 = ~n14625 & ~n14866;
  assign n15336 = ~n14635 & n15335;
  assign n15337 = ~n14866 & n15334;
  assign n15338 = n14633 & ~n33718;
  assign n15339 = n14636 & n15335;
  assign n15340 = ~n14625 & n14633;
  assign n15341 = ~n14635 & n15340;
  assign n15342 = ~n14866 & n15341;
  assign n15343 = ~n14633 & ~n33718;
  assign n15344 = ~n15342 & ~n15343;
  assign n15345 = ~n15338 & ~n15339;
  assign n15346 = ~n33717 & ~n33719;
  assign n15347 = ~n15330 & ~n15346;
  assign n15348 = ~n1567 & ~n15347;
  assign n15349 = n1567 & ~n15330;
  assign n15350 = ~n15346 & n15349;
  assign n15351 = ~n14638 & ~n33629;
  assign n15352 = ~n14638 & ~n14866;
  assign n15353 = ~n33629 & n15352;
  assign n15354 = ~n14866 & n15351;
  assign n15355 = n14646 & ~n33720;
  assign n15356 = n14650 & n15352;
  assign n15357 = n14646 & ~n33629;
  assign n15358 = ~n14638 & n15357;
  assign n15359 = ~n14866 & n15358;
  assign n15360 = ~n14646 & ~n33720;
  assign n15361 = ~n15359 & ~n15360;
  assign n15362 = ~n15355 & ~n15356;
  assign n15363 = ~n15350 & ~n33721;
  assign n15364 = ~n15348 & ~n15363;
  assign n15365 = ~n1374 & ~n15364;
  assign n15366 = ~n14652 & ~n14654;
  assign n15367 = ~n14866 & n15366;
  assign n15368 = ~n33631 & ~n15367;
  assign n15369 = ~n14652 & n33631;
  assign n15370 = ~n14654 & n15369;
  assign n15371 = n33631 & n15367;
  assign n15372 = ~n14866 & n15370;
  assign n15373 = ~n15368 & ~n33722;
  assign n15374 = n1374 & ~n15348;
  assign n15375 = ~n15363 & n15374;
  assign n15376 = n1374 & n15364;
  assign n15377 = ~n15373 & ~n33723;
  assign n15378 = ~n15365 & ~n15377;
  assign n15379 = ~n1179 & ~n15378;
  assign n15380 = n1179 & ~n15365;
  assign n15381 = ~n15377 & n15380;
  assign n15382 = ~n14669 & ~n33633;
  assign n15383 = ~n14669 & ~n14866;
  assign n15384 = ~n33633 & n15383;
  assign n15385 = ~n14866 & n15382;
  assign n15386 = n14677 & ~n33724;
  assign n15387 = n14681 & n15383;
  assign n15388 = n14677 & ~n33633;
  assign n15389 = ~n14669 & n15388;
  assign n15390 = ~n14866 & n15389;
  assign n15391 = ~n14677 & ~n33724;
  assign n15392 = ~n15390 & ~n15391;
  assign n15393 = ~n15386 & ~n15387;
  assign n15394 = ~n15381 & ~n33725;
  assign n15395 = ~n15379 & ~n15394;
  assign n15396 = ~n1016 & ~n15395;
  assign n15397 = n1016 & ~n15379;
  assign n15398 = ~n15394 & n15397;
  assign n15399 = n1016 & n15395;
  assign n15400 = ~n14683 & ~n14693;
  assign n15401 = ~n14683 & ~n14866;
  assign n15402 = ~n14693 & n15401;
  assign n15403 = ~n14866 & n15400;
  assign n15404 = n14691 & ~n33727;
  assign n15405 = n14694 & n15401;
  assign n15406 = ~n14683 & n14691;
  assign n15407 = ~n14693 & n15406;
  assign n15408 = ~n14866 & n15407;
  assign n15409 = ~n14691 & ~n33727;
  assign n15410 = ~n15408 & ~n15409;
  assign n15411 = ~n15404 & ~n15405;
  assign n15412 = ~n33726 & ~n33728;
  assign n15413 = ~n15396 & ~n15412;
  assign n15414 = ~n855 & ~n15413;
  assign n15415 = n855 & ~n15396;
  assign n15416 = ~n15412 & n15415;
  assign n15417 = ~n14696 & ~n33636;
  assign n15418 = ~n14696 & ~n14866;
  assign n15419 = ~n33636 & n15418;
  assign n15420 = ~n14866 & n15417;
  assign n15421 = n14704 & ~n33729;
  assign n15422 = n14708 & n15418;
  assign n15423 = n14704 & ~n33636;
  assign n15424 = ~n14696 & n15423;
  assign n15425 = ~n14866 & n15424;
  assign n15426 = ~n14704 & ~n33729;
  assign n15427 = ~n15425 & ~n15426;
  assign n15428 = ~n15421 & ~n15422;
  assign n15429 = ~n15416 & ~n33730;
  assign n15430 = ~n15414 & ~n15429;
  assign n15431 = ~n720 & ~n15430;
  assign n15432 = ~n14710 & ~n14712;
  assign n15433 = ~n14866 & n15432;
  assign n15434 = ~n33638 & ~n15433;
  assign n15435 = ~n14710 & n33638;
  assign n15436 = ~n14712 & n15435;
  assign n15437 = n33638 & n15433;
  assign n15438 = ~n14866 & n15436;
  assign n15439 = ~n15434 & ~n33731;
  assign n15440 = n720 & ~n15414;
  assign n15441 = ~n15429 & n15440;
  assign n15442 = n720 & n15430;
  assign n15443 = ~n15439 & ~n33732;
  assign n15444 = ~n15431 & ~n15443;
  assign n15445 = ~n592 & ~n15444;
  assign n15446 = n592 & ~n15431;
  assign n15447 = ~n15443 & n15446;
  assign n15448 = ~n14727 & ~n33640;
  assign n15449 = ~n14727 & ~n14866;
  assign n15450 = ~n33640 & n15449;
  assign n15451 = ~n14866 & n15448;
  assign n15452 = n14735 & ~n33733;
  assign n15453 = n14739 & n15449;
  assign n15454 = n14735 & ~n33640;
  assign n15455 = ~n14727 & n15454;
  assign n15456 = ~n14866 & n15455;
  assign n15457 = ~n14735 & ~n33733;
  assign n15458 = ~n15456 & ~n15457;
  assign n15459 = ~n15452 & ~n15453;
  assign n15460 = ~n15447 & ~n33734;
  assign n15461 = ~n15445 & ~n15460;
  assign n15462 = ~n487 & ~n15461;
  assign n15463 = n487 & ~n15445;
  assign n15464 = ~n15460 & n15463;
  assign n15465 = n487 & n15461;
  assign n15466 = ~n14741 & ~n14751;
  assign n15467 = ~n14741 & ~n14866;
  assign n15468 = ~n14751 & n15467;
  assign n15469 = ~n14866 & n15466;
  assign n15470 = n14749 & ~n33736;
  assign n15471 = n14752 & n15467;
  assign n15472 = ~n14741 & n14749;
  assign n15473 = ~n14751 & n15472;
  assign n15474 = ~n14866 & n15473;
  assign n15475 = ~n14749 & ~n33736;
  assign n15476 = ~n15474 & ~n15475;
  assign n15477 = ~n15470 & ~n15471;
  assign n15478 = ~n33735 & ~n33737;
  assign n15479 = ~n15462 & ~n15478;
  assign n15480 = ~n393 & ~n15479;
  assign n15481 = n393 & ~n15462;
  assign n15482 = ~n15478 & n15481;
  assign n15483 = ~n14754 & ~n33643;
  assign n15484 = ~n14754 & ~n14866;
  assign n15485 = ~n33643 & n15484;
  assign n15486 = ~n14866 & n15483;
  assign n15487 = n14762 & ~n33738;
  assign n15488 = n14766 & n15484;
  assign n15489 = n14762 & ~n33643;
  assign n15490 = ~n14754 & n15489;
  assign n15491 = ~n14866 & n15490;
  assign n15492 = ~n14762 & ~n33738;
  assign n15493 = ~n15491 & ~n15492;
  assign n15494 = ~n15487 & ~n15488;
  assign n15495 = ~n15482 & ~n33739;
  assign n15496 = ~n15480 & ~n15495;
  assign n15497 = ~n321 & ~n15496;
  assign n15498 = ~n14768 & ~n14770;
  assign n15499 = ~n14866 & n15498;
  assign n15500 = ~n33645 & ~n15499;
  assign n15501 = ~n14768 & n33645;
  assign n15502 = ~n14770 & n15501;
  assign n15503 = n33645 & n15499;
  assign n15504 = ~n14866 & n15502;
  assign n15505 = ~n15500 & ~n33740;
  assign n15506 = n321 & ~n15480;
  assign n15507 = ~n15495 & n15506;
  assign n15508 = n321 & n15496;
  assign n15509 = ~n15505 & ~n33741;
  assign n15510 = ~n15497 & ~n15509;
  assign n15511 = ~n263 & ~n15510;
  assign n15512 = n263 & ~n15497;
  assign n15513 = ~n15509 & n15512;
  assign n15514 = ~n14785 & ~n33647;
  assign n15515 = ~n14785 & ~n14866;
  assign n15516 = ~n33647 & n15515;
  assign n15517 = ~n14866 & n15514;
  assign n15518 = n14793 & ~n33742;
  assign n15519 = n14797 & n15515;
  assign n15520 = n14793 & ~n33647;
  assign n15521 = ~n14785 & n15520;
  assign n15522 = ~n14866 & n15521;
  assign n15523 = ~n14793 & ~n33742;
  assign n15524 = ~n15522 & ~n15523;
  assign n15525 = ~n15518 & ~n15519;
  assign n15526 = ~n15513 & ~n33743;
  assign n15527 = ~n15511 & ~n15526;
  assign n15528 = ~n214 & ~n15527;
  assign n15529 = n214 & ~n15511;
  assign n15530 = ~n15526 & n15529;
  assign n15531 = n214 & n15527;
  assign n15532 = ~n14799 & ~n14809;
  assign n15533 = ~n14799 & ~n14866;
  assign n15534 = ~n14809 & n15533;
  assign n15535 = ~n14866 & n15532;
  assign n15536 = n14807 & ~n33745;
  assign n15537 = n14810 & n15533;
  assign n15538 = ~n14799 & n14807;
  assign n15539 = ~n14809 & n15538;
  assign n15540 = ~n14866 & n15539;
  assign n15541 = ~n14807 & ~n33745;
  assign n15542 = ~n15540 & ~n15541;
  assign n15543 = ~n15536 & ~n15537;
  assign n15544 = ~n33744 & ~n33746;
  assign n15545 = ~n15528 & ~n15544;
  assign n15546 = ~n197 & ~n15545;
  assign n15547 = n197 & ~n15528;
  assign n15548 = ~n15544 & n15547;
  assign n15549 = ~n14812 & ~n33650;
  assign n15550 = ~n14812 & ~n14866;
  assign n15551 = ~n33650 & n15550;
  assign n15552 = ~n14866 & n15549;
  assign n15553 = n14820 & ~n33747;
  assign n15554 = n14824 & n15550;
  assign n15555 = n14820 & ~n33650;
  assign n15556 = ~n14812 & n15555;
  assign n15557 = ~n14866 & n15556;
  assign n15558 = ~n14820 & ~n33747;
  assign n15559 = ~n15557 & ~n15558;
  assign n15560 = ~n15553 & ~n15554;
  assign n15561 = ~n15548 & ~n33748;
  assign n15562 = ~n15546 & ~n15561;
  assign n15563 = ~n14826 & ~n14828;
  assign n15564 = ~n14866 & n15563;
  assign n15565 = ~n33652 & ~n15564;
  assign n15566 = ~n14826 & n33652;
  assign n15567 = ~n14828 & n15566;
  assign n15568 = n33652 & n15564;
  assign n15569 = ~n14866 & n15567;
  assign n15570 = ~n15565 & ~n33749;
  assign n15571 = ~n14842 & ~n14850;
  assign n15572 = ~n14850 & ~n14866;
  assign n15573 = ~n14842 & n15572;
  assign n15574 = ~n14866 & n15571;
  assign n15575 = ~n33655 & ~n33750;
  assign n15576 = ~n15570 & n15575;
  assign n15577 = ~n15562 & n15576;
  assign n15578 = n193 & ~n15577;
  assign n15579 = ~n15546 & n15570;
  assign n15580 = ~n15561 & n15579;
  assign n15581 = n15562 & n15570;
  assign n15582 = n14842 & ~n15572;
  assign n15583 = ~n193 & ~n15571;
  assign n15584 = ~n15582 & n15583;
  assign n15585 = ~n33751 & ~n15584;
  assign n15586 = ~n15578 & n15585;
  assign n15587 = ~n15202 & ~n33701;
  assign n15588 = ~n15586 & n15587;
  assign n15589 = ~n33703 & ~n15588;
  assign n15590 = ~n15202 & n33703;
  assign n15591 = ~n33701 & n15590;
  assign n15592 = n33703 & n15588;
  assign n15593 = ~n15586 & n15591;
  assign n15594 = ~n15589 & ~n33752;
  assign n15595 = ~n15185 & ~n15187;
  assign n15596 = ~n15586 & n15595;
  assign n15597 = ~n33700 & ~n15596;
  assign n15598 = ~n15187 & n33700;
  assign n15599 = ~n15185 & n15598;
  assign n15600 = n33700 & n15596;
  assign n15601 = ~n15586 & n15599;
  assign n15602 = ~n15597 & ~n33753;
  assign n15603 = ~n15154 & ~n15156;
  assign n15604 = ~n15586 & n15603;
  assign n15605 = ~n33696 & ~n15604;
  assign n15606 = ~n15156 & n33696;
  assign n15607 = ~n15154 & n15606;
  assign n15608 = n33696 & n15604;
  assign n15609 = ~n15586 & n15607;
  assign n15610 = ~n15605 & ~n33754;
  assign n15611 = ~n15136 & ~n33692;
  assign n15612 = ~n15586 & n15611;
  assign n15613 = ~n33694 & ~n15612;
  assign n15614 = ~n15136 & n33694;
  assign n15615 = ~n33692 & n15614;
  assign n15616 = n33694 & n15612;
  assign n15617 = ~n15586 & n15615;
  assign n15618 = ~n15613 & ~n33755;
  assign n15619 = ~n15119 & ~n15121;
  assign n15620 = ~n15586 & n15619;
  assign n15621 = ~n33691 & ~n15620;
  assign n15622 = ~n15121 & n33691;
  assign n15623 = ~n15119 & n15622;
  assign n15624 = n33691 & n15620;
  assign n15625 = ~n15586 & n15623;
  assign n15626 = ~n15621 & ~n33756;
  assign n15627 = ~n15088 & ~n15090;
  assign n15628 = ~n15586 & n15627;
  assign n15629 = ~n33687 & ~n15628;
  assign n15630 = ~n15090 & n33687;
  assign n15631 = ~n15088 & n15630;
  assign n15632 = n33687 & n15628;
  assign n15633 = ~n15586 & n15631;
  assign n15634 = ~n15629 & ~n33757;
  assign n15635 = ~n15069 & ~n33682;
  assign n15636 = ~n15586 & n15635;
  assign n15637 = ~n33685 & ~n15636;
  assign n15638 = ~n15069 & n33685;
  assign n15639 = ~n33682 & n15638;
  assign n15640 = n33685 & n15636;
  assign n15641 = ~n15586 & n15639;
  assign n15642 = ~n15637 & ~n33758;
  assign n15643 = ~n15052 & ~n15054;
  assign n15644 = ~n15586 & n15643;
  assign n15645 = ~n33681 & ~n15644;
  assign n15646 = ~n15054 & n33681;
  assign n15647 = ~n15052 & n15646;
  assign n15648 = n33681 & n15644;
  assign n15649 = ~n15586 & n15647;
  assign n15650 = ~n15645 & ~n33759;
  assign n15651 = ~n15018 & ~n15020;
  assign n15652 = ~n15586 & n15651;
  assign n15653 = ~n33676 & ~n15652;
  assign n15654 = ~n15020 & n33676;
  assign n15655 = ~n15018 & n15654;
  assign n15656 = n33676 & n15652;
  assign n15657 = ~n15586 & n15655;
  assign n15658 = ~n15653 & ~n33760;
  assign n15659 = ~n14985 & ~n14987;
  assign n15660 = ~n15586 & n15659;
  assign n15661 = ~n33672 & ~n15660;
  assign n15662 = ~n14987 & n33672;
  assign n15663 = ~n14985 & n15662;
  assign n15664 = n33672 & n15660;
  assign n15665 = ~n15586 & n15663;
  assign n15666 = ~n15661 & ~n33761;
  assign n15667 = ~n14952 & ~n14954;
  assign n15668 = ~n15586 & n15667;
  assign n15669 = ~n33668 & ~n15668;
  assign n15670 = ~n14954 & n33668;
  assign n15671 = ~n14952 & n15670;
  assign n15672 = n33668 & n15668;
  assign n15673 = ~n15586 & n15671;
  assign n15674 = ~n15669 & ~n33762;
  assign n15675 = ~n14918 & ~n14920;
  assign n15676 = ~n15586 & n15675;
  assign n15677 = ~n33663 & ~n15676;
  assign n15678 = ~n14920 & n33663;
  assign n15679 = ~n14918 & n15678;
  assign n15680 = n33663 & n15676;
  assign n15681 = ~n15586 & n15679;
  assign n15682 = ~n15677 & ~n33763;
  assign n15683 = ~n14891 & ~n14893;
  assign n15684 = ~n15586 & n15683;
  assign n15685 = ~n14902 & ~n15684;
  assign n15686 = ~n14893 & n14902;
  assign n15687 = ~n14891 & n15686;
  assign n15688 = n14902 & n15684;
  assign n15689 = ~n15586 & n15687;
  assign n15690 = ~n15685 & ~n33764;
  assign n15691 = ~pi38  & ~n15586;
  assign n15692 = ~pi39  & n15691;
  assign n15693 = n14868 & ~n15586;
  assign n15694 = ~n14866 & ~n15584;
  assign n15695 = ~n33751 & n15694;
  assign n15696 = ~n15578 & n15695;
  assign n15697 = ~n33765 & ~n15696;
  assign n15698 = pi40  & ~n15697;
  assign n15699 = ~pi40  & ~n15696;
  assign n15700 = ~pi40  & n15697;
  assign n15701 = ~n33765 & n15699;
  assign n15702 = ~n15698 & ~n33766;
  assign n15703 = pi38  & ~n15586;
  assign n15704 = ~pi36  & ~pi37 ;
  assign n15705 = ~pi38  & n15704;
  assign n15706 = ~n14214 & ~n33657;
  assign n15707 = ~n14215 & n15706;
  assign n15708 = ~n14231 & n15707;
  assign n15709 = ~n33578 & n15708;
  assign n15710 = n33576 & n14233;
  assign n15711 = ~n14225 & n15709;
  assign n15712 = ~n15705 & ~n33767;
  assign n15713 = ~n14864 & n15712;
  assign n15714 = ~n33655 & n15713;
  assign n15715 = ~n14858 & n15714;
  assign n15716 = ~n15703 & ~n15705;
  assign n15717 = n14866 & n15716;
  assign n15718 = ~n15703 & n15715;
  assign n15719 = pi39  & ~n15691;
  assign n15720 = ~n33765 & ~n15719;
  assign n15721 = ~n33768 & n15720;
  assign n15722 = ~n14866 & ~n15716;
  assign n15723 = n14233 & ~n15722;
  assign n15724 = ~n15721 & ~n15722;
  assign n15725 = n14233 & n15724;
  assign n15726 = ~n15721 & n15723;
  assign n15727 = ~n15702 & ~n33769;
  assign n15728 = ~n14233 & ~n15724;
  assign n15729 = n13548 & ~n15728;
  assign n15730 = ~n15727 & n15729;
  assign n15731 = ~n14871 & ~n33658;
  assign n15732 = ~n15586 & n15731;
  assign n15733 = n14876 & ~n15732;
  assign n15734 = ~n14876 & n15731;
  assign n15735 = ~n14876 & n15732;
  assign n15736 = ~n15586 & n15734;
  assign n15737 = ~n15733 & ~n33770;
  assign n15738 = ~n15730 & ~n15737;
  assign n15739 = ~n15727 & ~n15728;
  assign n15740 = ~n13548 & ~n15739;
  assign n15741 = n12948 & ~n15740;
  assign n15742 = ~n15738 & ~n15740;
  assign n15743 = n12948 & n15742;
  assign n15744 = ~n15738 & n15741;
  assign n15745 = ~n15690 & ~n33771;
  assign n15746 = ~n12948 & ~n15742;
  assign n15747 = n12296 & ~n15746;
  assign n15748 = ~n15745 & n15747;
  assign n15749 = ~n14905 & ~n33660;
  assign n15750 = ~n15586 & n15749;
  assign n15751 = ~n14915 & ~n15750;
  assign n15752 = ~n14905 & n14915;
  assign n15753 = ~n33660 & n15752;
  assign n15754 = n14915 & n15750;
  assign n15755 = ~n15586 & n15753;
  assign n15756 = n14915 & ~n15750;
  assign n15757 = ~n14915 & n15750;
  assign n15758 = ~n15756 & ~n15757;
  assign n15759 = ~n15751 & ~n33772;
  assign n15760 = ~n15748 & n33773;
  assign n15761 = ~n15745 & ~n15746;
  assign n15762 = ~n12296 & ~n15761;
  assign n15763 = n11719 & ~n15762;
  assign n15764 = ~n15760 & ~n15762;
  assign n15765 = n11719 & n15764;
  assign n15766 = ~n15760 & n15763;
  assign n15767 = ~n15682 & ~n33774;
  assign n15768 = ~n11719 & ~n15764;
  assign n15769 = n11097 & ~n15768;
  assign n15770 = ~n15767 & n15769;
  assign n15771 = ~n14935 & ~n33664;
  assign n15772 = ~n15586 & n15771;
  assign n15773 = ~n33666 & ~n15772;
  assign n15774 = n33666 & n15772;
  assign n15775 = ~n14935 & ~n33666;
  assign n15776 = ~n33664 & n15775;
  assign n15777 = ~n15586 & n15776;
  assign n15778 = n33666 & ~n15772;
  assign n15779 = ~n15777 & ~n15778;
  assign n15780 = ~n15773 & ~n15774;
  assign n15781 = ~n15770 & ~n33775;
  assign n15782 = ~n15767 & ~n15768;
  assign n15783 = ~n11097 & ~n15782;
  assign n15784 = n10555 & ~n15783;
  assign n15785 = ~n15781 & ~n15783;
  assign n15786 = n10555 & n15785;
  assign n15787 = ~n15781 & n15784;
  assign n15788 = ~n15674 & ~n33776;
  assign n15789 = ~n10555 & ~n15785;
  assign n15790 = n9969 & ~n15789;
  assign n15791 = ~n15788 & n15790;
  assign n15792 = ~n14969 & ~n33669;
  assign n15793 = ~n15586 & n15792;
  assign n15794 = ~n33670 & n15793;
  assign n15795 = n33670 & ~n15793;
  assign n15796 = ~n14969 & n33670;
  assign n15797 = ~n33669 & n15796;
  assign n15798 = ~n15586 & n15797;
  assign n15799 = ~n33670 & ~n15793;
  assign n15800 = ~n15798 & ~n15799;
  assign n15801 = ~n15794 & ~n15795;
  assign n15802 = ~n15791 & ~n33777;
  assign n15803 = ~n15788 & ~n15789;
  assign n15804 = ~n9969 & ~n15803;
  assign n15805 = n9457 & ~n15804;
  assign n15806 = ~n15802 & ~n15804;
  assign n15807 = n9457 & n15806;
  assign n15808 = ~n15802 & n15805;
  assign n15809 = ~n15666 & ~n33778;
  assign n15810 = ~n9457 & ~n15806;
  assign n15811 = n8896 & ~n15810;
  assign n15812 = ~n15809 & n15811;
  assign n15813 = ~n15002 & ~n33673;
  assign n15814 = ~n15586 & n15813;
  assign n15815 = ~n33674 & n15814;
  assign n15816 = n33674 & ~n15814;
  assign n15817 = ~n33674 & ~n15814;
  assign n15818 = ~n15002 & n33674;
  assign n15819 = ~n33673 & n15818;
  assign n15820 = n33674 & n15814;
  assign n15821 = ~n15586 & n15819;
  assign n15822 = ~n15817 & ~n33779;
  assign n15823 = ~n15815 & ~n15816;
  assign n15824 = ~n15812 & ~n33780;
  assign n15825 = ~n15809 & ~n15810;
  assign n15826 = ~n8896 & ~n15825;
  assign n15827 = n8411 & ~n15826;
  assign n15828 = ~n15824 & ~n15826;
  assign n15829 = n8411 & n15828;
  assign n15830 = ~n15824 & n15827;
  assign n15831 = ~n15658 & ~n33781;
  assign n15832 = ~n8411 & ~n15828;
  assign n15833 = n7885 & ~n15832;
  assign n15834 = ~n15831 & n15833;
  assign n15835 = ~n15035 & ~n33677;
  assign n15836 = ~n15035 & ~n15586;
  assign n15837 = ~n33677 & n15836;
  assign n15838 = ~n15586 & n15835;
  assign n15839 = n33679 & ~n33782;
  assign n15840 = n15050 & n15836;
  assign n15841 = ~n33679 & n33782;
  assign n15842 = ~n15035 & n33679;
  assign n15843 = ~n33677 & n15842;
  assign n15844 = ~n15586 & n15843;
  assign n15845 = ~n33679 & ~n33782;
  assign n15846 = ~n15844 & ~n15845;
  assign n15847 = ~n15839 & ~n33783;
  assign n15848 = ~n15834 & ~n33784;
  assign n15849 = ~n15831 & ~n15832;
  assign n15850 = ~n7885 & ~n15849;
  assign n15851 = n7428 & ~n15850;
  assign n15852 = ~n15848 & ~n15850;
  assign n15853 = n7428 & n15852;
  assign n15854 = ~n15848 & n15851;
  assign n15855 = ~n15650 & ~n33785;
  assign n15856 = ~n7428 & ~n15852;
  assign n15857 = n6937 & ~n15856;
  assign n15858 = ~n15855 & n15857;
  assign n15859 = ~n15642 & ~n15858;
  assign n15860 = ~n15855 & ~n15856;
  assign n15861 = ~n6937 & ~n15860;
  assign n15862 = n6507 & ~n15861;
  assign n15863 = ~n15859 & ~n15861;
  assign n15864 = n6507 & n15863;
  assign n15865 = ~n15859 & n15862;
  assign n15866 = ~n15634 & ~n33786;
  assign n15867 = ~n6507 & ~n15863;
  assign n15868 = n6051 & ~n15867;
  assign n15869 = ~n15866 & n15868;
  assign n15870 = ~n15105 & ~n33689;
  assign n15871 = ~n15105 & ~n15586;
  assign n15872 = ~n33689 & n15871;
  assign n15873 = ~n15586 & n15870;
  assign n15874 = n15113 & ~n33787;
  assign n15875 = n15117 & n15871;
  assign n15876 = ~n15105 & n15113;
  assign n15877 = ~n33689 & n15876;
  assign n15878 = ~n15586 & n15877;
  assign n15879 = ~n15113 & ~n33787;
  assign n15880 = ~n15878 & ~n15879;
  assign n15881 = ~n15874 & ~n15875;
  assign n15882 = ~n15869 & ~n33788;
  assign n15883 = ~n15866 & ~n15867;
  assign n15884 = ~n6051 & ~n15883;
  assign n15885 = n5648 & ~n15884;
  assign n15886 = ~n15882 & ~n15884;
  assign n15887 = n5648 & n15886;
  assign n15888 = ~n15882 & n15885;
  assign n15889 = ~n15626 & ~n33789;
  assign n15890 = ~n5648 & ~n15886;
  assign n15891 = n5223 & ~n15890;
  assign n15892 = ~n15889 & n15891;
  assign n15893 = ~n15618 & ~n15892;
  assign n15894 = ~n15889 & ~n15890;
  assign n15895 = ~n5223 & ~n15894;
  assign n15896 = n4851 & ~n15895;
  assign n15897 = ~n15893 & ~n15895;
  assign n15898 = n4851 & n15897;
  assign n15899 = ~n15893 & n15896;
  assign n15900 = ~n15610 & ~n33790;
  assign n15901 = ~n4851 & ~n15897;
  assign n15902 = n4461 & ~n15901;
  assign n15903 = ~n15900 & n15902;
  assign n15904 = ~n15171 & ~n33698;
  assign n15905 = ~n15171 & ~n15586;
  assign n15906 = ~n33698 & n15905;
  assign n15907 = ~n15586 & n15904;
  assign n15908 = n15179 & ~n33791;
  assign n15909 = n15183 & n15905;
  assign n15910 = ~n15171 & n15179;
  assign n15911 = ~n33698 & n15910;
  assign n15912 = ~n15586 & n15911;
  assign n15913 = ~n15179 & ~n33791;
  assign n15914 = ~n15912 & ~n15913;
  assign n15915 = ~n15908 & ~n15909;
  assign n15916 = ~n15903 & ~n33792;
  assign n15917 = ~n15900 & ~n15901;
  assign n15918 = ~n4461 & ~n15917;
  assign n15919 = n4115 & ~n15918;
  assign n15920 = ~n15916 & ~n15918;
  assign n15921 = n4115 & n15920;
  assign n15922 = ~n15916 & n15919;
  assign n15923 = ~n15602 & ~n33793;
  assign n15924 = ~n4115 & ~n15920;
  assign n15925 = n3754 & ~n15924;
  assign n15926 = ~n15923 & n15925;
  assign n15927 = ~n15594 & ~n15926;
  assign n15928 = ~n15923 & ~n15924;
  assign n15929 = ~n3754 & ~n15928;
  assign n15930 = n3444 & ~n15929;
  assign n15931 = ~n15927 & ~n15929;
  assign n15932 = n3444 & n15931;
  assign n15933 = ~n15927 & n15930;
  assign n15934 = ~n15220 & ~n15222;
  assign n15935 = ~n15586 & n15934;
  assign n15936 = ~n33704 & n15935;
  assign n15937 = n33704 & ~n15935;
  assign n15938 = ~n15222 & n33704;
  assign n15939 = ~n15220 & n15938;
  assign n15940 = ~n15586 & n15939;
  assign n15941 = ~n33704 & ~n15935;
  assign n15942 = ~n15940 & ~n15941;
  assign n15943 = ~n15936 & ~n15937;
  assign n15944 = ~n33794 & ~n33795;
  assign n15945 = ~n3444 & ~n15931;
  assign n15946 = ~n15944 & ~n15945;
  assign n15947 = ~n3116 & ~n15946;
  assign n15948 = ~n15235 & ~n33706;
  assign n15949 = ~n15586 & n15948;
  assign n15950 = n33705 & ~n15949;
  assign n15951 = ~n33705 & n15949;
  assign n15952 = ~n15235 & n33705;
  assign n15953 = ~n33706 & n15952;
  assign n15954 = ~n15586 & n15953;
  assign n15955 = ~n33705 & ~n15949;
  assign n15956 = ~n15954 & ~n15955;
  assign n15957 = ~n15950 & ~n15951;
  assign n15958 = n3116 & ~n15945;
  assign n15959 = ~n15944 & n15958;
  assign n15960 = ~n33796 & ~n15959;
  assign n15961 = ~n15947 & ~n15960;
  assign n15962 = ~n2833 & ~n15961;
  assign n15963 = ~n15251 & ~n15253;
  assign n15964 = ~n15586 & n15963;
  assign n15965 = ~n33708 & ~n15964;
  assign n15966 = ~n15253 & n33708;
  assign n15967 = ~n15251 & n15966;
  assign n15968 = n33708 & n15964;
  assign n15969 = ~n15586 & n15967;
  assign n15970 = ~n15965 & ~n33797;
  assign n15971 = n2833 & ~n15947;
  assign n15972 = n2833 & n15961;
  assign n15973 = ~n15960 & n15971;
  assign n15974 = ~n15970 & ~n33798;
  assign n15975 = ~n15962 & ~n15974;
  assign n15976 = ~n2536 & ~n15975;
  assign n15977 = n2536 & ~n15962;
  assign n15978 = ~n15974 & n15977;
  assign n15979 = ~n15268 & ~n33710;
  assign n15980 = ~n15268 & ~n15586;
  assign n15981 = ~n33710 & n15980;
  assign n15982 = ~n15586 & n15979;
  assign n15983 = n15276 & ~n33799;
  assign n15984 = n15280 & n15980;
  assign n15985 = ~n15268 & n15276;
  assign n15986 = ~n33710 & n15985;
  assign n15987 = ~n15586 & n15986;
  assign n15988 = ~n15276 & ~n33799;
  assign n15989 = ~n15987 & ~n15988;
  assign n15990 = ~n15983 & ~n15984;
  assign n15991 = ~n15978 & ~n33800;
  assign n15992 = ~n15976 & ~n15991;
  assign n15993 = ~n2283 & ~n15992;
  assign n15994 = ~n15282 & ~n15284;
  assign n15995 = ~n15586 & n15994;
  assign n15996 = ~n33712 & ~n15995;
  assign n15997 = ~n15284 & n33712;
  assign n15998 = ~n15282 & n15997;
  assign n15999 = n33712 & n15995;
  assign n16000 = ~n15586 & n15998;
  assign n16001 = ~n15996 & ~n33801;
  assign n16002 = n2283 & ~n15976;
  assign n16003 = n2283 & n15992;
  assign n16004 = ~n15991 & n16002;
  assign n16005 = ~n16001 & ~n33802;
  assign n16006 = ~n15993 & ~n16005;
  assign n16007 = ~n2021 & ~n16006;
  assign n16008 = n2021 & ~n15993;
  assign n16009 = ~n16005 & n16008;
  assign n16010 = ~n15299 & ~n33714;
  assign n16011 = ~n15299 & ~n15586;
  assign n16012 = ~n33714 & n16011;
  assign n16013 = ~n15586 & n16010;
  assign n16014 = n15307 & ~n33803;
  assign n16015 = n15311 & n16011;
  assign n16016 = ~n15299 & n15307;
  assign n16017 = ~n33714 & n16016;
  assign n16018 = ~n15586 & n16017;
  assign n16019 = ~n15307 & ~n33803;
  assign n16020 = ~n16018 & ~n16019;
  assign n16021 = ~n16014 & ~n16015;
  assign n16022 = ~n16009 & ~n33804;
  assign n16023 = ~n16007 & ~n16022;
  assign n16024 = ~n1796 & ~n16023;
  assign n16025 = ~n15313 & ~n15315;
  assign n16026 = ~n15586 & n16025;
  assign n16027 = ~n33716 & ~n16026;
  assign n16028 = ~n15315 & n33716;
  assign n16029 = ~n15313 & n16028;
  assign n16030 = n33716 & n16026;
  assign n16031 = ~n15586 & n16029;
  assign n16032 = ~n16027 & ~n33805;
  assign n16033 = n1796 & ~n16007;
  assign n16034 = n1796 & n16023;
  assign n16035 = ~n16022 & n16033;
  assign n16036 = ~n16032 & ~n33806;
  assign n16037 = ~n16024 & ~n16036;
  assign n16038 = ~n1567 & ~n16037;
  assign n16039 = ~n15330 & ~n33717;
  assign n16040 = ~n15586 & n16039;
  assign n16041 = ~n33719 & ~n16040;
  assign n16042 = ~n15330 & n33719;
  assign n16043 = ~n33717 & n16042;
  assign n16044 = n33719 & n16040;
  assign n16045 = ~n15586 & n16043;
  assign n16046 = ~n16041 & ~n33807;
  assign n16047 = n1567 & ~n16024;
  assign n16048 = ~n16036 & n16047;
  assign n16049 = ~n16046 & ~n16048;
  assign n16050 = ~n16038 & ~n16049;
  assign n16051 = ~n1374 & ~n16050;
  assign n16052 = ~n15348 & ~n15350;
  assign n16053 = ~n15586 & n16052;
  assign n16054 = ~n33721 & ~n16053;
  assign n16055 = ~n15350 & n33721;
  assign n16056 = ~n15348 & n16055;
  assign n16057 = n33721 & n16053;
  assign n16058 = ~n15586 & n16056;
  assign n16059 = ~n16054 & ~n33808;
  assign n16060 = n1374 & ~n16038;
  assign n16061 = n1374 & n16050;
  assign n16062 = ~n16049 & n16060;
  assign n16063 = ~n16059 & ~n33809;
  assign n16064 = ~n16051 & ~n16063;
  assign n16065 = ~n1179 & ~n16064;
  assign n16066 = n1179 & ~n16051;
  assign n16067 = ~n16063 & n16066;
  assign n16068 = ~n15365 & ~n33723;
  assign n16069 = ~n15365 & ~n15586;
  assign n16070 = ~n33723 & n16069;
  assign n16071 = ~n15586 & n16068;
  assign n16072 = n15373 & ~n33810;
  assign n16073 = n15377 & n16069;
  assign n16074 = ~n15365 & n15373;
  assign n16075 = ~n33723 & n16074;
  assign n16076 = ~n15586 & n16075;
  assign n16077 = ~n15373 & ~n33810;
  assign n16078 = ~n16076 & ~n16077;
  assign n16079 = ~n16072 & ~n16073;
  assign n16080 = ~n16067 & ~n33811;
  assign n16081 = ~n16065 & ~n16080;
  assign n16082 = ~n1016 & ~n16081;
  assign n16083 = ~n15379 & ~n15381;
  assign n16084 = ~n15586 & n16083;
  assign n16085 = ~n33725 & ~n16084;
  assign n16086 = ~n15381 & n33725;
  assign n16087 = ~n15379 & n16086;
  assign n16088 = n33725 & n16084;
  assign n16089 = ~n15586 & n16087;
  assign n16090 = ~n16085 & ~n33812;
  assign n16091 = n1016 & ~n16065;
  assign n16092 = n1016 & n16081;
  assign n16093 = ~n16080 & n16091;
  assign n16094 = ~n16090 & ~n33813;
  assign n16095 = ~n16082 & ~n16094;
  assign n16096 = ~n855 & ~n16095;
  assign n16097 = ~n15396 & ~n33726;
  assign n16098 = ~n15586 & n16097;
  assign n16099 = ~n33728 & ~n16098;
  assign n16100 = ~n15396 & n33728;
  assign n16101 = ~n33726 & n16100;
  assign n16102 = n33728 & n16098;
  assign n16103 = ~n15586 & n16101;
  assign n16104 = ~n16099 & ~n33814;
  assign n16105 = n855 & ~n16082;
  assign n16106 = ~n16094 & n16105;
  assign n16107 = ~n16104 & ~n16106;
  assign n16108 = ~n16096 & ~n16107;
  assign n16109 = ~n720 & ~n16108;
  assign n16110 = ~n15414 & ~n15416;
  assign n16111 = ~n15586 & n16110;
  assign n16112 = ~n33730 & ~n16111;
  assign n16113 = ~n15416 & n33730;
  assign n16114 = ~n15414 & n16113;
  assign n16115 = n33730 & n16111;
  assign n16116 = ~n15586 & n16114;
  assign n16117 = ~n16112 & ~n33815;
  assign n16118 = n720 & ~n16096;
  assign n16119 = n720 & n16108;
  assign n16120 = ~n16107 & n16118;
  assign n16121 = ~n16117 & ~n33816;
  assign n16122 = ~n16109 & ~n16121;
  assign n16123 = ~n592 & ~n16122;
  assign n16124 = n592 & ~n16109;
  assign n16125 = ~n16121 & n16124;
  assign n16126 = ~n15431 & ~n33732;
  assign n16127 = ~n15431 & ~n15586;
  assign n16128 = ~n33732 & n16127;
  assign n16129 = ~n15586 & n16126;
  assign n16130 = n15439 & ~n33817;
  assign n16131 = n15443 & n16127;
  assign n16132 = ~n15431 & n15439;
  assign n16133 = ~n33732 & n16132;
  assign n16134 = ~n15586 & n16133;
  assign n16135 = ~n15439 & ~n33817;
  assign n16136 = ~n16134 & ~n16135;
  assign n16137 = ~n16130 & ~n16131;
  assign n16138 = ~n16125 & ~n33818;
  assign n16139 = ~n16123 & ~n16138;
  assign n16140 = ~n487 & ~n16139;
  assign n16141 = ~n15445 & ~n15447;
  assign n16142 = ~n15586 & n16141;
  assign n16143 = ~n33734 & ~n16142;
  assign n16144 = ~n15447 & n33734;
  assign n16145 = ~n15445 & n16144;
  assign n16146 = n33734 & n16142;
  assign n16147 = ~n15586 & n16145;
  assign n16148 = ~n16143 & ~n33819;
  assign n16149 = n487 & ~n16123;
  assign n16150 = n487 & n16139;
  assign n16151 = ~n16138 & n16149;
  assign n16152 = ~n16148 & ~n33820;
  assign n16153 = ~n16140 & ~n16152;
  assign n16154 = ~n393 & ~n16153;
  assign n16155 = ~n15462 & ~n33735;
  assign n16156 = ~n15586 & n16155;
  assign n16157 = ~n33737 & ~n16156;
  assign n16158 = ~n15462 & n33737;
  assign n16159 = ~n33735 & n16158;
  assign n16160 = n33737 & n16156;
  assign n16161 = ~n15586 & n16159;
  assign n16162 = ~n16157 & ~n33821;
  assign n16163 = n393 & ~n16140;
  assign n16164 = ~n16152 & n16163;
  assign n16165 = ~n16162 & ~n16164;
  assign n16166 = ~n16154 & ~n16165;
  assign n16167 = ~n321 & ~n16166;
  assign n16168 = ~n15480 & ~n15482;
  assign n16169 = ~n15586 & n16168;
  assign n16170 = ~n33739 & ~n16169;
  assign n16171 = ~n15482 & n33739;
  assign n16172 = ~n15480 & n16171;
  assign n16173 = n33739 & n16169;
  assign n16174 = ~n15586 & n16172;
  assign n16175 = ~n16170 & ~n33822;
  assign n16176 = n321 & ~n16154;
  assign n16177 = n321 & n16166;
  assign n16178 = ~n16165 & n16176;
  assign n16179 = ~n16175 & ~n33823;
  assign n16180 = ~n16167 & ~n16179;
  assign n16181 = ~n263 & ~n16180;
  assign n16182 = n263 & ~n16167;
  assign n16183 = ~n16179 & n16182;
  assign n16184 = ~n15497 & ~n33741;
  assign n16185 = ~n15497 & ~n15586;
  assign n16186 = ~n33741 & n16185;
  assign n16187 = ~n15586 & n16184;
  assign n16188 = n15505 & ~n33824;
  assign n16189 = n15509 & n16185;
  assign n16190 = ~n15497 & n15505;
  assign n16191 = ~n33741 & n16190;
  assign n16192 = ~n15586 & n16191;
  assign n16193 = ~n15505 & ~n33824;
  assign n16194 = ~n16192 & ~n16193;
  assign n16195 = ~n16188 & ~n16189;
  assign n16196 = ~n16183 & ~n33825;
  assign n16197 = ~n16181 & ~n16196;
  assign n16198 = ~n214 & ~n16197;
  assign n16199 = ~n15511 & ~n15513;
  assign n16200 = ~n15586 & n16199;
  assign n16201 = ~n33743 & ~n16200;
  assign n16202 = ~n15513 & n33743;
  assign n16203 = ~n15511 & n16202;
  assign n16204 = n33743 & n16200;
  assign n16205 = ~n15586 & n16203;
  assign n16206 = ~n16201 & ~n33826;
  assign n16207 = n214 & ~n16181;
  assign n16208 = n214 & n16197;
  assign n16209 = ~n16196 & n16207;
  assign n16210 = ~n16206 & ~n33827;
  assign n16211 = ~n16198 & ~n16210;
  assign n16212 = ~n197 & ~n16211;
  assign n16213 = ~n15528 & ~n33744;
  assign n16214 = ~n15586 & n16213;
  assign n16215 = ~n33746 & ~n16214;
  assign n16216 = ~n15528 & n33746;
  assign n16217 = ~n33744 & n16216;
  assign n16218 = n33746 & n16214;
  assign n16219 = ~n15586 & n16217;
  assign n16220 = ~n16215 & ~n33828;
  assign n16221 = n197 & ~n16198;
  assign n16222 = ~n16210 & n16221;
  assign n16223 = ~n16220 & ~n16222;
  assign n16224 = ~n16212 & ~n16223;
  assign n16225 = ~n15546 & ~n15548;
  assign n16226 = ~n15586 & n16225;
  assign n16227 = ~n33748 & ~n16226;
  assign n16228 = ~n15548 & n33748;
  assign n16229 = ~n15546 & n16228;
  assign n16230 = n33748 & n16226;
  assign n16231 = ~n15586 & n16229;
  assign n16232 = ~n16227 & ~n33829;
  assign n16233 = ~n15562 & ~n15570;
  assign n16234 = ~n15570 & ~n15586;
  assign n16235 = ~n15562 & n16234;
  assign n16236 = ~n15586 & n16233;
  assign n16237 = ~n33751 & ~n33830;
  assign n16238 = ~n16232 & n16237;
  assign n16239 = ~n16224 & n16238;
  assign n16240 = n193 & ~n16239;
  assign n16241 = ~n16212 & n16232;
  assign n16242 = n16224 & n16232;
  assign n16243 = ~n16223 & n16241;
  assign n16244 = n15562 & ~n16234;
  assign n16245 = ~n193 & ~n16233;
  assign n16246 = ~n16244 & n16245;
  assign n16247 = ~n33831 & ~n16246;
  assign n16248 = ~n16240 & n16247;
  assign n16249 = pi36  & ~n16248;
  assign n16250 = ~pi34  & ~pi35 ;
  assign n16251 = ~pi36  & n16250;
  assign n16252 = ~n16249 & ~n16251;
  assign n16253 = ~n15586 & ~n16252;
  assign n16254 = ~pi36  & ~n16248;
  assign n16255 = pi37  & ~n16254;
  assign n16256 = ~pi37  & n16254;
  assign n16257 = n15704 & ~n16248;
  assign n16258 = ~n16255 & ~n33832;
  assign n16259 = ~n33653 & ~n33767;
  assign n16260 = ~n14845 & n16259;
  assign n16261 = ~n14864 & n16260;
  assign n16262 = ~n33655 & n16261;
  assign n16263 = n14850 & n14866;
  assign n16264 = ~n14858 & n16262;
  assign n16265 = ~n16251 & ~n33833;
  assign n16266 = ~n15584 & n16265;
  assign n16267 = ~n33751 & n16266;
  assign n16268 = ~n15578 & n16267;
  assign n16269 = n15586 & n16252;
  assign n16270 = ~n16249 & n16268;
  assign n16271 = n16258 & ~n33834;
  assign n16272 = ~n16253 & ~n16271;
  assign n16273 = ~n14866 & ~n16272;
  assign n16274 = n14866 & ~n16253;
  assign n16275 = ~n16271 & n16274;
  assign n16276 = ~n15586 & ~n16246;
  assign n16277 = ~n33831 & n16276;
  assign n16278 = ~n16240 & n16277;
  assign n16279 = ~n33832 & ~n16278;
  assign n16280 = pi38  & ~n16279;
  assign n16281 = ~pi38  & ~n16278;
  assign n16282 = ~pi38  & n16279;
  assign n16283 = ~n33832 & n16281;
  assign n16284 = ~n16280 & ~n33835;
  assign n16285 = ~n16275 & ~n16284;
  assign n16286 = ~n16273 & ~n16285;
  assign n16287 = ~n14233 & ~n16286;
  assign n16288 = n14233 & ~n16273;
  assign n16289 = ~n16285 & n16288;
  assign n16290 = n14233 & n16286;
  assign n16291 = ~n33768 & ~n15722;
  assign n16292 = ~n16248 & n16291;
  assign n16293 = n15720 & ~n16292;
  assign n16294 = ~n15720 & n16291;
  assign n16295 = ~n15720 & n16292;
  assign n16296 = ~n16248 & n16294;
  assign n16297 = ~n16293 & ~n33837;
  assign n16298 = ~n33836 & ~n16297;
  assign n16299 = ~n16287 & ~n16298;
  assign n16300 = ~n13548 & ~n16299;
  assign n16301 = n13548 & ~n16287;
  assign n16302 = ~n16298 & n16301;
  assign n16303 = ~n33769 & ~n15728;
  assign n16304 = ~n15728 & ~n16248;
  assign n16305 = ~n33769 & n16304;
  assign n16306 = ~n16248 & n16303;
  assign n16307 = n15702 & ~n33838;
  assign n16308 = n15727 & n16304;
  assign n16309 = n15702 & ~n33769;
  assign n16310 = ~n15728 & n16309;
  assign n16311 = ~n16248 & n16310;
  assign n16312 = ~n15702 & ~n33838;
  assign n16313 = ~n16311 & ~n16312;
  assign n16314 = ~n16307 & ~n16308;
  assign n16315 = ~n16302 & ~n33839;
  assign n16316 = ~n16300 & ~n16315;
  assign n16317 = ~n12948 & ~n16316;
  assign n16318 = n12948 & ~n16300;
  assign n16319 = ~n16315 & n16318;
  assign n16320 = n12948 & n16316;
  assign n16321 = ~n15730 & ~n15740;
  assign n16322 = ~n16248 & n16321;
  assign n16323 = ~n15737 & ~n16322;
  assign n16324 = n15737 & ~n15740;
  assign n16325 = ~n15730 & n16324;
  assign n16326 = n15737 & n16322;
  assign n16327 = ~n16248 & n16325;
  assign n16328 = n15737 & ~n16322;
  assign n16329 = ~n15737 & n16322;
  assign n16330 = ~n16328 & ~n16329;
  assign n16331 = ~n16323 & ~n33841;
  assign n16332 = ~n33840 & n33842;
  assign n16333 = ~n16317 & ~n16332;
  assign n16334 = ~n12296 & ~n16333;
  assign n16335 = n12296 & ~n16317;
  assign n16336 = ~n16332 & n16335;
  assign n16337 = ~n33771 & ~n15746;
  assign n16338 = ~n15746 & ~n16248;
  assign n16339 = ~n33771 & n16338;
  assign n16340 = ~n16248 & n16337;
  assign n16341 = n15690 & ~n33843;
  assign n16342 = n15745 & n16338;
  assign n16343 = n15690 & ~n33771;
  assign n16344 = ~n15746 & n16343;
  assign n16345 = ~n16248 & n16344;
  assign n16346 = ~n15690 & ~n33843;
  assign n16347 = ~n16345 & ~n16346;
  assign n16348 = ~n16341 & ~n16342;
  assign n16349 = ~n16336 & ~n33844;
  assign n16350 = ~n16334 & ~n16349;
  assign n16351 = ~n11719 & ~n16350;
  assign n16352 = n11719 & ~n16334;
  assign n16353 = ~n16349 & n16352;
  assign n16354 = n11719 & n16350;
  assign n16355 = ~n15748 & ~n15762;
  assign n16356 = ~n16248 & n16355;
  assign n16357 = ~n33773 & ~n16356;
  assign n16358 = n33773 & n16356;
  assign n16359 = ~n33773 & ~n15762;
  assign n16360 = ~n15748 & n16359;
  assign n16361 = ~n16248 & n16360;
  assign n16362 = n33773 & ~n16356;
  assign n16363 = ~n16361 & ~n16362;
  assign n16364 = ~n16357 & ~n16358;
  assign n16365 = ~n33845 & ~n33846;
  assign n16366 = ~n16351 & ~n16365;
  assign n16367 = ~n11097 & ~n16366;
  assign n16368 = n11097 & ~n16351;
  assign n16369 = ~n16365 & n16368;
  assign n16370 = ~n33774 & ~n15768;
  assign n16371 = ~n15768 & ~n16248;
  assign n16372 = ~n33774 & n16371;
  assign n16373 = ~n16248 & n16370;
  assign n16374 = n15682 & ~n33847;
  assign n16375 = n15767 & n16371;
  assign n16376 = n15682 & ~n33774;
  assign n16377 = ~n15768 & n16376;
  assign n16378 = ~n16248 & n16377;
  assign n16379 = ~n15682 & ~n33847;
  assign n16380 = ~n16378 & ~n16379;
  assign n16381 = ~n16374 & ~n16375;
  assign n16382 = ~n16369 & ~n33848;
  assign n16383 = ~n16367 & ~n16382;
  assign n16384 = ~n10555 & ~n16383;
  assign n16385 = n10555 & ~n16367;
  assign n16386 = ~n16382 & n16385;
  assign n16387 = n10555 & n16383;
  assign n16388 = ~n15770 & ~n15783;
  assign n16389 = ~n16248 & n16388;
  assign n16390 = ~n33775 & n16389;
  assign n16391 = n33775 & ~n16389;
  assign n16392 = n33775 & ~n15783;
  assign n16393 = ~n15770 & n16392;
  assign n16394 = ~n16248 & n16393;
  assign n16395 = ~n33775 & ~n16389;
  assign n16396 = ~n16394 & ~n16395;
  assign n16397 = ~n16390 & ~n16391;
  assign n16398 = ~n33849 & ~n33850;
  assign n16399 = ~n16384 & ~n16398;
  assign n16400 = ~n9969 & ~n16399;
  assign n16401 = n9969 & ~n16384;
  assign n16402 = ~n16398 & n16401;
  assign n16403 = ~n33776 & ~n15789;
  assign n16404 = ~n15789 & ~n16248;
  assign n16405 = ~n33776 & n16404;
  assign n16406 = ~n16248 & n16403;
  assign n16407 = n15674 & ~n33851;
  assign n16408 = n15788 & n16404;
  assign n16409 = n15674 & ~n33776;
  assign n16410 = ~n15789 & n16409;
  assign n16411 = ~n16248 & n16410;
  assign n16412 = ~n15674 & ~n33851;
  assign n16413 = ~n16411 & ~n16412;
  assign n16414 = ~n16407 & ~n16408;
  assign n16415 = ~n16402 & ~n33852;
  assign n16416 = ~n16400 & ~n16415;
  assign n16417 = ~n9457 & ~n16416;
  assign n16418 = n9457 & ~n16400;
  assign n16419 = ~n16415 & n16418;
  assign n16420 = n9457 & n16416;
  assign n16421 = ~n15791 & ~n15804;
  assign n16422 = ~n16248 & n16421;
  assign n16423 = ~n33777 & n16422;
  assign n16424 = n33777 & ~n16422;
  assign n16425 = ~n33777 & ~n16422;
  assign n16426 = n33777 & ~n15804;
  assign n16427 = ~n15791 & n16426;
  assign n16428 = n33777 & n16422;
  assign n16429 = ~n16248 & n16427;
  assign n16430 = ~n16425 & ~n33854;
  assign n16431 = ~n16423 & ~n16424;
  assign n16432 = ~n33853 & ~n33855;
  assign n16433 = ~n16417 & ~n16432;
  assign n16434 = ~n8896 & ~n16433;
  assign n16435 = n8896 & ~n16417;
  assign n16436 = ~n16432 & n16435;
  assign n16437 = ~n33778 & ~n15810;
  assign n16438 = ~n15810 & ~n16248;
  assign n16439 = ~n33778 & n16438;
  assign n16440 = ~n16248 & n16437;
  assign n16441 = n15666 & ~n33856;
  assign n16442 = n15809 & n16438;
  assign n16443 = n15666 & ~n33778;
  assign n16444 = ~n15810 & n16443;
  assign n16445 = ~n16248 & n16444;
  assign n16446 = ~n15666 & ~n33856;
  assign n16447 = ~n16445 & ~n16446;
  assign n16448 = ~n16441 & ~n16442;
  assign n16449 = ~n16436 & ~n33857;
  assign n16450 = ~n16434 & ~n16449;
  assign n16451 = ~n8411 & ~n16450;
  assign n16452 = n8411 & ~n16434;
  assign n16453 = ~n16449 & n16452;
  assign n16454 = n8411 & n16450;
  assign n16455 = ~n15812 & ~n15826;
  assign n16456 = ~n15826 & ~n16248;
  assign n16457 = ~n15812 & n16456;
  assign n16458 = ~n16248 & n16455;
  assign n16459 = n33780 & ~n33859;
  assign n16460 = n15824 & n16456;
  assign n16461 = ~n33780 & n33859;
  assign n16462 = n33780 & ~n15826;
  assign n16463 = ~n15812 & n16462;
  assign n16464 = ~n16248 & n16463;
  assign n16465 = ~n33780 & ~n33859;
  assign n16466 = ~n16464 & ~n16465;
  assign n16467 = ~n16459 & ~n33860;
  assign n16468 = ~n33858 & ~n33861;
  assign n16469 = ~n16451 & ~n16468;
  assign n16470 = ~n7885 & ~n16469;
  assign n16471 = n7885 & ~n16451;
  assign n16472 = ~n16468 & n16471;
  assign n16473 = ~n33781 & ~n15832;
  assign n16474 = ~n15832 & ~n16248;
  assign n16475 = ~n33781 & n16474;
  assign n16476 = ~n16248 & n16473;
  assign n16477 = n15658 & ~n33862;
  assign n16478 = n15831 & n16474;
  assign n16479 = n15658 & ~n33781;
  assign n16480 = ~n15832 & n16479;
  assign n16481 = ~n16248 & n16480;
  assign n16482 = ~n15658 & ~n33862;
  assign n16483 = ~n16481 & ~n16482;
  assign n16484 = ~n16477 & ~n16478;
  assign n16485 = ~n16472 & ~n33863;
  assign n16486 = ~n16470 & ~n16485;
  assign n16487 = ~n7428 & ~n16486;
  assign n16488 = ~n15834 & ~n15850;
  assign n16489 = ~n16248 & n16488;
  assign n16490 = ~n33784 & ~n16489;
  assign n16491 = n33784 & ~n15850;
  assign n16492 = ~n15834 & n16491;
  assign n16493 = n33784 & n16489;
  assign n16494 = ~n16248 & n16492;
  assign n16495 = ~n16490 & ~n33864;
  assign n16496 = n7428 & ~n16470;
  assign n16497 = ~n16485 & n16496;
  assign n16498 = n7428 & n16486;
  assign n16499 = ~n16495 & ~n33865;
  assign n16500 = ~n16487 & ~n16499;
  assign n16501 = ~n6937 & ~n16500;
  assign n16502 = n6937 & ~n16487;
  assign n16503 = ~n16499 & n16502;
  assign n16504 = ~n33785 & ~n15856;
  assign n16505 = ~n15856 & ~n16248;
  assign n16506 = ~n33785 & n16505;
  assign n16507 = ~n16248 & n16504;
  assign n16508 = n15650 & ~n33866;
  assign n16509 = n15855 & n16505;
  assign n16510 = n15650 & ~n33785;
  assign n16511 = ~n15856 & n16510;
  assign n16512 = ~n16248 & n16511;
  assign n16513 = ~n15650 & ~n33866;
  assign n16514 = ~n16512 & ~n16513;
  assign n16515 = ~n16508 & ~n16509;
  assign n16516 = ~n16503 & ~n33867;
  assign n16517 = ~n16501 & ~n16516;
  assign n16518 = ~n6507 & ~n16517;
  assign n16519 = n6507 & ~n16501;
  assign n16520 = ~n16516 & n16519;
  assign n16521 = n6507 & n16517;
  assign n16522 = ~n15858 & ~n15861;
  assign n16523 = ~n15861 & ~n16248;
  assign n16524 = ~n15858 & n16523;
  assign n16525 = ~n16248 & n16522;
  assign n16526 = n15642 & ~n33869;
  assign n16527 = n15859 & n16523;
  assign n16528 = n15642 & ~n15861;
  assign n16529 = ~n15858 & n16528;
  assign n16530 = ~n16248 & n16529;
  assign n16531 = ~n15642 & ~n33869;
  assign n16532 = ~n16530 & ~n16531;
  assign n16533 = ~n16526 & ~n16527;
  assign n16534 = ~n33868 & ~n33870;
  assign n16535 = ~n16518 & ~n16534;
  assign n16536 = ~n6051 & ~n16535;
  assign n16537 = n6051 & ~n16518;
  assign n16538 = ~n16534 & n16537;
  assign n16539 = ~n33786 & ~n15867;
  assign n16540 = ~n15867 & ~n16248;
  assign n16541 = ~n33786 & n16540;
  assign n16542 = ~n16248 & n16539;
  assign n16543 = n15634 & ~n33871;
  assign n16544 = n15866 & n16540;
  assign n16545 = n15634 & ~n33786;
  assign n16546 = ~n15867 & n16545;
  assign n16547 = ~n16248 & n16546;
  assign n16548 = ~n15634 & ~n33871;
  assign n16549 = ~n16547 & ~n16548;
  assign n16550 = ~n16543 & ~n16544;
  assign n16551 = ~n16538 & ~n33872;
  assign n16552 = ~n16536 & ~n16551;
  assign n16553 = ~n5648 & ~n16552;
  assign n16554 = ~n15869 & ~n15884;
  assign n16555 = ~n16248 & n16554;
  assign n16556 = ~n33788 & ~n16555;
  assign n16557 = n33788 & ~n15884;
  assign n16558 = ~n15869 & n16557;
  assign n16559 = n33788 & n16555;
  assign n16560 = ~n16248 & n16558;
  assign n16561 = ~n16556 & ~n33873;
  assign n16562 = n5648 & ~n16536;
  assign n16563 = ~n16551 & n16562;
  assign n16564 = n5648 & n16552;
  assign n16565 = ~n16561 & ~n33874;
  assign n16566 = ~n16553 & ~n16565;
  assign n16567 = ~n5223 & ~n16566;
  assign n16568 = n5223 & ~n16553;
  assign n16569 = ~n16565 & n16568;
  assign n16570 = ~n33789 & ~n15890;
  assign n16571 = ~n15890 & ~n16248;
  assign n16572 = ~n33789 & n16571;
  assign n16573 = ~n16248 & n16570;
  assign n16574 = n15626 & ~n33875;
  assign n16575 = n15889 & n16571;
  assign n16576 = n15626 & ~n33789;
  assign n16577 = ~n15890 & n16576;
  assign n16578 = ~n16248 & n16577;
  assign n16579 = ~n15626 & ~n33875;
  assign n16580 = ~n16578 & ~n16579;
  assign n16581 = ~n16574 & ~n16575;
  assign n16582 = ~n16569 & ~n33876;
  assign n16583 = ~n16567 & ~n16582;
  assign n16584 = ~n4851 & ~n16583;
  assign n16585 = n4851 & ~n16567;
  assign n16586 = ~n16582 & n16585;
  assign n16587 = n4851 & n16583;
  assign n16588 = ~n15892 & ~n15895;
  assign n16589 = ~n15895 & ~n16248;
  assign n16590 = ~n15892 & n16589;
  assign n16591 = ~n16248 & n16588;
  assign n16592 = n15618 & ~n33878;
  assign n16593 = n15893 & n16589;
  assign n16594 = n15618 & ~n15895;
  assign n16595 = ~n15892 & n16594;
  assign n16596 = ~n16248 & n16595;
  assign n16597 = ~n15618 & ~n33878;
  assign n16598 = ~n16596 & ~n16597;
  assign n16599 = ~n16592 & ~n16593;
  assign n16600 = ~n33877 & ~n33879;
  assign n16601 = ~n16584 & ~n16600;
  assign n16602 = ~n4461 & ~n16601;
  assign n16603 = n4461 & ~n16584;
  assign n16604 = ~n16600 & n16603;
  assign n16605 = ~n33790 & ~n15901;
  assign n16606 = ~n15901 & ~n16248;
  assign n16607 = ~n33790 & n16606;
  assign n16608 = ~n16248 & n16605;
  assign n16609 = n15610 & ~n33880;
  assign n16610 = n15900 & n16606;
  assign n16611 = n15610 & ~n33790;
  assign n16612 = ~n15901 & n16611;
  assign n16613 = ~n16248 & n16612;
  assign n16614 = ~n15610 & ~n33880;
  assign n16615 = ~n16613 & ~n16614;
  assign n16616 = ~n16609 & ~n16610;
  assign n16617 = ~n16604 & ~n33881;
  assign n16618 = ~n16602 & ~n16617;
  assign n16619 = ~n4115 & ~n16618;
  assign n16620 = ~n15903 & ~n15918;
  assign n16621 = ~n16248 & n16620;
  assign n16622 = ~n33792 & ~n16621;
  assign n16623 = n33792 & ~n15918;
  assign n16624 = ~n15903 & n16623;
  assign n16625 = n33792 & n16621;
  assign n16626 = ~n16248 & n16624;
  assign n16627 = ~n16622 & ~n33882;
  assign n16628 = n4115 & ~n16602;
  assign n16629 = ~n16617 & n16628;
  assign n16630 = n4115 & n16618;
  assign n16631 = ~n16627 & ~n33883;
  assign n16632 = ~n16619 & ~n16631;
  assign n16633 = ~n3754 & ~n16632;
  assign n16634 = n3754 & ~n16619;
  assign n16635 = ~n16631 & n16634;
  assign n16636 = ~n33793 & ~n15924;
  assign n16637 = ~n15924 & ~n16248;
  assign n16638 = ~n33793 & n16637;
  assign n16639 = ~n16248 & n16636;
  assign n16640 = n15602 & ~n33884;
  assign n16641 = n15923 & n16637;
  assign n16642 = n15602 & ~n33793;
  assign n16643 = ~n15924 & n16642;
  assign n16644 = ~n16248 & n16643;
  assign n16645 = ~n15602 & ~n33884;
  assign n16646 = ~n16644 & ~n16645;
  assign n16647 = ~n16640 & ~n16641;
  assign n16648 = ~n16635 & ~n33885;
  assign n16649 = ~n16633 & ~n16648;
  assign n16650 = ~n3444 & ~n16649;
  assign n16651 = n3444 & ~n16633;
  assign n16652 = ~n16648 & n16651;
  assign n16653 = n3444 & n16649;
  assign n16654 = ~n15926 & ~n15929;
  assign n16655 = ~n15929 & ~n16248;
  assign n16656 = ~n15926 & n16655;
  assign n16657 = ~n16248 & n16654;
  assign n16658 = n15594 & ~n33887;
  assign n16659 = n15927 & n16655;
  assign n16660 = n15594 & ~n15929;
  assign n16661 = ~n15926 & n16660;
  assign n16662 = ~n16248 & n16661;
  assign n16663 = ~n15594 & ~n33887;
  assign n16664 = ~n16662 & ~n16663;
  assign n16665 = ~n16658 & ~n16659;
  assign n16666 = ~n33886 & ~n33888;
  assign n16667 = ~n16650 & ~n16666;
  assign n16668 = ~n3116 & ~n16667;
  assign n16669 = n3116 & ~n16650;
  assign n16670 = ~n16666 & n16669;
  assign n16671 = ~n33794 & ~n15945;
  assign n16672 = ~n16248 & n16671;
  assign n16673 = ~n33795 & n16672;
  assign n16674 = n33795 & ~n16672;
  assign n16675 = ~n33794 & n33795;
  assign n16676 = ~n15945 & n16675;
  assign n16677 = ~n16248 & n16676;
  assign n16678 = ~n33795 & ~n16672;
  assign n16679 = ~n16677 & ~n16678;
  assign n16680 = ~n16673 & ~n16674;
  assign n16681 = ~n16670 & ~n33889;
  assign n16682 = ~n16668 & ~n16681;
  assign n16683 = ~n2833 & ~n16682;
  assign n16684 = ~n15947 & ~n15959;
  assign n16685 = ~n16248 & n16684;
  assign n16686 = ~n33796 & ~n16685;
  assign n16687 = ~n15947 & n33796;
  assign n16688 = ~n15959 & n16687;
  assign n16689 = n33796 & n16685;
  assign n16690 = ~n16248 & n16688;
  assign n16691 = ~n16686 & ~n33890;
  assign n16692 = n2833 & ~n16668;
  assign n16693 = ~n16681 & n16692;
  assign n16694 = n2833 & n16682;
  assign n16695 = ~n16691 & ~n33891;
  assign n16696 = ~n16683 & ~n16695;
  assign n16697 = ~n2536 & ~n16696;
  assign n16698 = n2536 & ~n16683;
  assign n16699 = ~n16695 & n16698;
  assign n16700 = ~n15962 & ~n33798;
  assign n16701 = ~n15962 & ~n16248;
  assign n16702 = ~n33798 & n16701;
  assign n16703 = ~n16248 & n16700;
  assign n16704 = n15970 & ~n33892;
  assign n16705 = n15974 & n16701;
  assign n16706 = n15970 & ~n33798;
  assign n16707 = ~n15962 & n16706;
  assign n16708 = ~n16248 & n16707;
  assign n16709 = ~n15970 & ~n33892;
  assign n16710 = ~n16708 & ~n16709;
  assign n16711 = ~n16704 & ~n16705;
  assign n16712 = ~n16699 & ~n33893;
  assign n16713 = ~n16697 & ~n16712;
  assign n16714 = ~n2283 & ~n16713;
  assign n16715 = ~n15976 & ~n15978;
  assign n16716 = ~n16248 & n16715;
  assign n16717 = ~n33800 & ~n16716;
  assign n16718 = ~n15976 & n33800;
  assign n16719 = ~n15978 & n16718;
  assign n16720 = n33800 & n16716;
  assign n16721 = ~n16248 & n16719;
  assign n16722 = ~n16717 & ~n33894;
  assign n16723 = n2283 & ~n16697;
  assign n16724 = ~n16712 & n16723;
  assign n16725 = n2283 & n16713;
  assign n16726 = ~n16722 & ~n33895;
  assign n16727 = ~n16714 & ~n16726;
  assign n16728 = ~n2021 & ~n16727;
  assign n16729 = n2021 & ~n16714;
  assign n16730 = ~n16726 & n16729;
  assign n16731 = ~n15993 & ~n33802;
  assign n16732 = ~n15993 & ~n16248;
  assign n16733 = ~n33802 & n16732;
  assign n16734 = ~n16248 & n16731;
  assign n16735 = n16001 & ~n33896;
  assign n16736 = n16005 & n16732;
  assign n16737 = n16001 & ~n33802;
  assign n16738 = ~n15993 & n16737;
  assign n16739 = ~n16248 & n16738;
  assign n16740 = ~n16001 & ~n33896;
  assign n16741 = ~n16739 & ~n16740;
  assign n16742 = ~n16735 & ~n16736;
  assign n16743 = ~n16730 & ~n33897;
  assign n16744 = ~n16728 & ~n16743;
  assign n16745 = ~n1796 & ~n16744;
  assign n16746 = ~n16007 & ~n16009;
  assign n16747 = ~n16248 & n16746;
  assign n16748 = ~n33804 & ~n16747;
  assign n16749 = ~n16007 & n33804;
  assign n16750 = ~n16009 & n16749;
  assign n16751 = n33804 & n16747;
  assign n16752 = ~n16248 & n16750;
  assign n16753 = ~n16748 & ~n33898;
  assign n16754 = n1796 & ~n16728;
  assign n16755 = ~n16743 & n16754;
  assign n16756 = n1796 & n16744;
  assign n16757 = ~n16753 & ~n33899;
  assign n16758 = ~n16745 & ~n16757;
  assign n16759 = ~n1567 & ~n16758;
  assign n16760 = n1567 & ~n16745;
  assign n16761 = ~n16757 & n16760;
  assign n16762 = ~n16024 & ~n33806;
  assign n16763 = ~n16024 & ~n16248;
  assign n16764 = ~n33806 & n16763;
  assign n16765 = ~n16248 & n16762;
  assign n16766 = n16032 & ~n33900;
  assign n16767 = n16036 & n16763;
  assign n16768 = n16032 & ~n33806;
  assign n16769 = ~n16024 & n16768;
  assign n16770 = ~n16248 & n16769;
  assign n16771 = ~n16032 & ~n33900;
  assign n16772 = ~n16770 & ~n16771;
  assign n16773 = ~n16766 & ~n16767;
  assign n16774 = ~n16761 & ~n33901;
  assign n16775 = ~n16759 & ~n16774;
  assign n16776 = ~n1374 & ~n16775;
  assign n16777 = n1374 & ~n16759;
  assign n16778 = ~n16774 & n16777;
  assign n16779 = n1374 & n16775;
  assign n16780 = ~n16038 & ~n16048;
  assign n16781 = ~n16038 & ~n16248;
  assign n16782 = ~n16048 & n16781;
  assign n16783 = ~n16248 & n16780;
  assign n16784 = n16046 & ~n33903;
  assign n16785 = n16049 & n16781;
  assign n16786 = ~n16038 & n16046;
  assign n16787 = ~n16048 & n16786;
  assign n16788 = ~n16248 & n16787;
  assign n16789 = ~n16046 & ~n33903;
  assign n16790 = ~n16788 & ~n16789;
  assign n16791 = ~n16784 & ~n16785;
  assign n16792 = ~n33902 & ~n33904;
  assign n16793 = ~n16776 & ~n16792;
  assign n16794 = ~n1179 & ~n16793;
  assign n16795 = n1179 & ~n16776;
  assign n16796 = ~n16792 & n16795;
  assign n16797 = ~n16051 & ~n33809;
  assign n16798 = ~n16051 & ~n16248;
  assign n16799 = ~n33809 & n16798;
  assign n16800 = ~n16248 & n16797;
  assign n16801 = n16059 & ~n33905;
  assign n16802 = n16063 & n16798;
  assign n16803 = n16059 & ~n33809;
  assign n16804 = ~n16051 & n16803;
  assign n16805 = ~n16248 & n16804;
  assign n16806 = ~n16059 & ~n33905;
  assign n16807 = ~n16805 & ~n16806;
  assign n16808 = ~n16801 & ~n16802;
  assign n16809 = ~n16796 & ~n33906;
  assign n16810 = ~n16794 & ~n16809;
  assign n16811 = ~n1016 & ~n16810;
  assign n16812 = ~n16065 & ~n16067;
  assign n16813 = ~n16248 & n16812;
  assign n16814 = ~n33811 & ~n16813;
  assign n16815 = ~n16065 & n33811;
  assign n16816 = ~n16067 & n16815;
  assign n16817 = n33811 & n16813;
  assign n16818 = ~n16248 & n16816;
  assign n16819 = ~n16814 & ~n33907;
  assign n16820 = n1016 & ~n16794;
  assign n16821 = ~n16809 & n16820;
  assign n16822 = n1016 & n16810;
  assign n16823 = ~n16819 & ~n33908;
  assign n16824 = ~n16811 & ~n16823;
  assign n16825 = ~n855 & ~n16824;
  assign n16826 = n855 & ~n16811;
  assign n16827 = ~n16823 & n16826;
  assign n16828 = ~n16082 & ~n33813;
  assign n16829 = ~n16082 & ~n16248;
  assign n16830 = ~n33813 & n16829;
  assign n16831 = ~n16248 & n16828;
  assign n16832 = n16090 & ~n33909;
  assign n16833 = n16094 & n16829;
  assign n16834 = n16090 & ~n33813;
  assign n16835 = ~n16082 & n16834;
  assign n16836 = ~n16248 & n16835;
  assign n16837 = ~n16090 & ~n33909;
  assign n16838 = ~n16836 & ~n16837;
  assign n16839 = ~n16832 & ~n16833;
  assign n16840 = ~n16827 & ~n33910;
  assign n16841 = ~n16825 & ~n16840;
  assign n16842 = ~n720 & ~n16841;
  assign n16843 = n720 & ~n16825;
  assign n16844 = ~n16840 & n16843;
  assign n16845 = n720 & n16841;
  assign n16846 = ~n16096 & ~n16106;
  assign n16847 = ~n16096 & ~n16248;
  assign n16848 = ~n16106 & n16847;
  assign n16849 = ~n16248 & n16846;
  assign n16850 = n16104 & ~n33912;
  assign n16851 = n16107 & n16847;
  assign n16852 = ~n16096 & n16104;
  assign n16853 = ~n16106 & n16852;
  assign n16854 = ~n16248 & n16853;
  assign n16855 = ~n16104 & ~n33912;
  assign n16856 = ~n16854 & ~n16855;
  assign n16857 = ~n16850 & ~n16851;
  assign n16858 = ~n33911 & ~n33913;
  assign n16859 = ~n16842 & ~n16858;
  assign n16860 = ~n592 & ~n16859;
  assign n16861 = n592 & ~n16842;
  assign n16862 = ~n16858 & n16861;
  assign n16863 = ~n16109 & ~n33816;
  assign n16864 = ~n16109 & ~n16248;
  assign n16865 = ~n33816 & n16864;
  assign n16866 = ~n16248 & n16863;
  assign n16867 = n16117 & ~n33914;
  assign n16868 = n16121 & n16864;
  assign n16869 = n16117 & ~n33816;
  assign n16870 = ~n16109 & n16869;
  assign n16871 = ~n16248 & n16870;
  assign n16872 = ~n16117 & ~n33914;
  assign n16873 = ~n16871 & ~n16872;
  assign n16874 = ~n16867 & ~n16868;
  assign n16875 = ~n16862 & ~n33915;
  assign n16876 = ~n16860 & ~n16875;
  assign n16877 = ~n487 & ~n16876;
  assign n16878 = ~n16123 & ~n16125;
  assign n16879 = ~n16248 & n16878;
  assign n16880 = ~n33818 & ~n16879;
  assign n16881 = ~n16123 & n33818;
  assign n16882 = ~n16125 & n16881;
  assign n16883 = n33818 & n16879;
  assign n16884 = ~n16248 & n16882;
  assign n16885 = ~n16880 & ~n33916;
  assign n16886 = n487 & ~n16860;
  assign n16887 = ~n16875 & n16886;
  assign n16888 = n487 & n16876;
  assign n16889 = ~n16885 & ~n33917;
  assign n16890 = ~n16877 & ~n16889;
  assign n16891 = ~n393 & ~n16890;
  assign n16892 = n393 & ~n16877;
  assign n16893 = ~n16889 & n16892;
  assign n16894 = ~n16140 & ~n33820;
  assign n16895 = ~n16140 & ~n16248;
  assign n16896 = ~n33820 & n16895;
  assign n16897 = ~n16248 & n16894;
  assign n16898 = n16148 & ~n33918;
  assign n16899 = n16152 & n16895;
  assign n16900 = n16148 & ~n33820;
  assign n16901 = ~n16140 & n16900;
  assign n16902 = ~n16248 & n16901;
  assign n16903 = ~n16148 & ~n33918;
  assign n16904 = ~n16902 & ~n16903;
  assign n16905 = ~n16898 & ~n16899;
  assign n16906 = ~n16893 & ~n33919;
  assign n16907 = ~n16891 & ~n16906;
  assign n16908 = ~n321 & ~n16907;
  assign n16909 = n321 & ~n16891;
  assign n16910 = ~n16906 & n16909;
  assign n16911 = n321 & n16907;
  assign n16912 = ~n16154 & ~n16164;
  assign n16913 = ~n16154 & ~n16248;
  assign n16914 = ~n16164 & n16913;
  assign n16915 = ~n16248 & n16912;
  assign n16916 = n16162 & ~n33921;
  assign n16917 = n16165 & n16913;
  assign n16918 = ~n16154 & n16162;
  assign n16919 = ~n16164 & n16918;
  assign n16920 = ~n16248 & n16919;
  assign n16921 = ~n16162 & ~n33921;
  assign n16922 = ~n16920 & ~n16921;
  assign n16923 = ~n16916 & ~n16917;
  assign n16924 = ~n33920 & ~n33922;
  assign n16925 = ~n16908 & ~n16924;
  assign n16926 = ~n263 & ~n16925;
  assign n16927 = n263 & ~n16908;
  assign n16928 = ~n16924 & n16927;
  assign n16929 = ~n16167 & ~n33823;
  assign n16930 = ~n16167 & ~n16248;
  assign n16931 = ~n33823 & n16930;
  assign n16932 = ~n16248 & n16929;
  assign n16933 = n16175 & ~n33923;
  assign n16934 = n16179 & n16930;
  assign n16935 = n16175 & ~n33823;
  assign n16936 = ~n16167 & n16935;
  assign n16937 = ~n16248 & n16936;
  assign n16938 = ~n16175 & ~n33923;
  assign n16939 = ~n16937 & ~n16938;
  assign n16940 = ~n16933 & ~n16934;
  assign n16941 = ~n16928 & ~n33924;
  assign n16942 = ~n16926 & ~n16941;
  assign n16943 = ~n214 & ~n16942;
  assign n16944 = ~n16181 & ~n16183;
  assign n16945 = ~n16248 & n16944;
  assign n16946 = ~n33825 & ~n16945;
  assign n16947 = ~n16181 & n33825;
  assign n16948 = ~n16183 & n16947;
  assign n16949 = n33825 & n16945;
  assign n16950 = ~n16248 & n16948;
  assign n16951 = ~n16946 & ~n33925;
  assign n16952 = n214 & ~n16926;
  assign n16953 = ~n16941 & n16952;
  assign n16954 = n214 & n16942;
  assign n16955 = ~n16951 & ~n33926;
  assign n16956 = ~n16943 & ~n16955;
  assign n16957 = ~n197 & ~n16956;
  assign n16958 = n197 & ~n16943;
  assign n16959 = ~n16955 & n16958;
  assign n16960 = ~n16198 & ~n33827;
  assign n16961 = ~n16198 & ~n16248;
  assign n16962 = ~n33827 & n16961;
  assign n16963 = ~n16248 & n16960;
  assign n16964 = n16206 & ~n33927;
  assign n16965 = n16210 & n16961;
  assign n16966 = n16206 & ~n33827;
  assign n16967 = ~n16198 & n16966;
  assign n16968 = ~n16248 & n16967;
  assign n16969 = ~n16206 & ~n33927;
  assign n16970 = ~n16968 & ~n16969;
  assign n16971 = ~n16964 & ~n16965;
  assign n16972 = ~n16959 & ~n33928;
  assign n16973 = ~n16957 & ~n16972;
  assign n16974 = ~n16212 & ~n16222;
  assign n16975 = ~n16212 & ~n16248;
  assign n16976 = ~n16222 & n16975;
  assign n16977 = ~n16248 & n16974;
  assign n16978 = n16220 & ~n33929;
  assign n16979 = n16223 & n16975;
  assign n16980 = ~n16212 & n16220;
  assign n16981 = ~n16222 & n16980;
  assign n16982 = ~n16248 & n16981;
  assign n16983 = ~n16220 & ~n33929;
  assign n16984 = ~n16982 & ~n16983;
  assign n16985 = ~n16978 & ~n16979;
  assign n16986 = ~n16224 & ~n16232;
  assign n16987 = ~n16232 & ~n16248;
  assign n16988 = ~n16224 & n16987;
  assign n16989 = ~n16248 & n16986;
  assign n16990 = ~n33831 & ~n33931;
  assign n16991 = ~n33930 & n16990;
  assign n16992 = ~n16973 & n16991;
  assign n16993 = n193 & ~n16992;
  assign n16994 = ~n16957 & n33930;
  assign n16995 = ~n16972 & n16994;
  assign n16996 = n16973 & n33930;
  assign n16997 = n16224 & ~n16987;
  assign n16998 = ~n193 & ~n16986;
  assign n16999 = ~n16997 & n16998;
  assign n17000 = ~n33932 & ~n16999;
  assign n17001 = ~n16993 & n17000;
  assign n17002 = ~n16668 & ~n16670;
  assign n17003 = ~n17001 & n17002;
  assign n17004 = ~n33889 & ~n17003;
  assign n17005 = ~n16670 & n33889;
  assign n17006 = ~n16668 & n17005;
  assign n17007 = n33889 & n17003;
  assign n17008 = ~n17001 & n17006;
  assign n17009 = ~n17004 & ~n33933;
  assign n17010 = ~n16650 & ~n33886;
  assign n17011 = ~n17001 & n17010;
  assign n17012 = ~n33888 & ~n17011;
  assign n17013 = ~n16650 & n33888;
  assign n17014 = ~n33886 & n17013;
  assign n17015 = n33888 & n17011;
  assign n17016 = ~n17001 & n17014;
  assign n17017 = ~n17012 & ~n33934;
  assign n17018 = ~n16633 & ~n16635;
  assign n17019 = ~n17001 & n17018;
  assign n17020 = ~n33885 & ~n17019;
  assign n17021 = ~n16635 & n33885;
  assign n17022 = ~n16633 & n17021;
  assign n17023 = n33885 & n17019;
  assign n17024 = ~n17001 & n17022;
  assign n17025 = ~n17020 & ~n33935;
  assign n17026 = ~n16602 & ~n16604;
  assign n17027 = ~n17001 & n17026;
  assign n17028 = ~n33881 & ~n17027;
  assign n17029 = ~n16604 & n33881;
  assign n17030 = ~n16602 & n17029;
  assign n17031 = n33881 & n17027;
  assign n17032 = ~n17001 & n17030;
  assign n17033 = ~n17028 & ~n33936;
  assign n17034 = ~n16584 & ~n33877;
  assign n17035 = ~n17001 & n17034;
  assign n17036 = ~n33879 & ~n17035;
  assign n17037 = ~n16584 & n33879;
  assign n17038 = ~n33877 & n17037;
  assign n17039 = n33879 & n17035;
  assign n17040 = ~n17001 & n17038;
  assign n17041 = ~n17036 & ~n33937;
  assign n17042 = ~n16567 & ~n16569;
  assign n17043 = ~n17001 & n17042;
  assign n17044 = ~n33876 & ~n17043;
  assign n17045 = ~n16569 & n33876;
  assign n17046 = ~n16567 & n17045;
  assign n17047 = n33876 & n17043;
  assign n17048 = ~n17001 & n17046;
  assign n17049 = ~n17044 & ~n33938;
  assign n17050 = ~n16536 & ~n16538;
  assign n17051 = ~n17001 & n17050;
  assign n17052 = ~n33872 & ~n17051;
  assign n17053 = ~n16538 & n33872;
  assign n17054 = ~n16536 & n17053;
  assign n17055 = n33872 & n17051;
  assign n17056 = ~n17001 & n17054;
  assign n17057 = ~n17052 & ~n33939;
  assign n17058 = ~n16518 & ~n33868;
  assign n17059 = ~n17001 & n17058;
  assign n17060 = ~n33870 & ~n17059;
  assign n17061 = ~n16518 & n33870;
  assign n17062 = ~n33868 & n17061;
  assign n17063 = n33870 & n17059;
  assign n17064 = ~n17001 & n17062;
  assign n17065 = ~n17060 & ~n33940;
  assign n17066 = ~n16501 & ~n16503;
  assign n17067 = ~n17001 & n17066;
  assign n17068 = ~n33867 & ~n17067;
  assign n17069 = ~n16503 & n33867;
  assign n17070 = ~n16501 & n17069;
  assign n17071 = n33867 & n17067;
  assign n17072 = ~n17001 & n17070;
  assign n17073 = ~n17068 & ~n33941;
  assign n17074 = ~n16470 & ~n16472;
  assign n17075 = ~n17001 & n17074;
  assign n17076 = ~n33863 & ~n17075;
  assign n17077 = ~n16472 & n33863;
  assign n17078 = ~n16470 & n17077;
  assign n17079 = n33863 & n17075;
  assign n17080 = ~n17001 & n17078;
  assign n17081 = ~n17076 & ~n33942;
  assign n17082 = ~n16451 & ~n33858;
  assign n17083 = ~n17001 & n17082;
  assign n17084 = ~n33861 & ~n17083;
  assign n17085 = ~n16451 & n33861;
  assign n17086 = ~n33858 & n17085;
  assign n17087 = n33861 & n17083;
  assign n17088 = ~n17001 & n17086;
  assign n17089 = ~n17084 & ~n33943;
  assign n17090 = ~n16434 & ~n16436;
  assign n17091 = ~n17001 & n17090;
  assign n17092 = ~n33857 & ~n17091;
  assign n17093 = ~n16436 & n33857;
  assign n17094 = ~n16434 & n17093;
  assign n17095 = n33857 & n17091;
  assign n17096 = ~n17001 & n17094;
  assign n17097 = ~n17092 & ~n33944;
  assign n17098 = ~n16400 & ~n16402;
  assign n17099 = ~n17001 & n17098;
  assign n17100 = ~n33852 & ~n17099;
  assign n17101 = ~n16402 & n33852;
  assign n17102 = ~n16400 & n17101;
  assign n17103 = n33852 & n17099;
  assign n17104 = ~n17001 & n17102;
  assign n17105 = ~n17100 & ~n33945;
  assign n17106 = ~n16367 & ~n16369;
  assign n17107 = ~n17001 & n17106;
  assign n17108 = ~n33848 & ~n17107;
  assign n17109 = ~n16369 & n33848;
  assign n17110 = ~n16367 & n17109;
  assign n17111 = n33848 & n17107;
  assign n17112 = ~n17001 & n17110;
  assign n17113 = ~n17108 & ~n33946;
  assign n17114 = ~n16334 & ~n16336;
  assign n17115 = ~n17001 & n17114;
  assign n17116 = ~n33844 & ~n17115;
  assign n17117 = ~n16336 & n33844;
  assign n17118 = ~n16334 & n17117;
  assign n17119 = n33844 & n17115;
  assign n17120 = ~n17001 & n17118;
  assign n17121 = ~n17116 & ~n33947;
  assign n17122 = ~n16300 & ~n16302;
  assign n17123 = ~n17001 & n17122;
  assign n17124 = ~n33839 & ~n17123;
  assign n17125 = ~n16302 & n33839;
  assign n17126 = ~n16300 & n17125;
  assign n17127 = n33839 & n17123;
  assign n17128 = ~n17001 & n17126;
  assign n17129 = ~n17124 & ~n33948;
  assign n17130 = ~n16273 & ~n16275;
  assign n17131 = ~n17001 & n17130;
  assign n17132 = ~n16284 & ~n17131;
  assign n17133 = ~n16275 & n16284;
  assign n17134 = ~n16273 & n17133;
  assign n17135 = n16284 & n17131;
  assign n17136 = ~n17001 & n17134;
  assign n17137 = ~n17132 & ~n33949;
  assign n17138 = ~pi34  & ~n17001;
  assign n17139 = ~pi35  & n17138;
  assign n17140 = n16250 & ~n17001;
  assign n17141 = ~n16248 & ~n16999;
  assign n17142 = ~n33932 & n17141;
  assign n17143 = ~n16993 & n17142;
  assign n17144 = ~n33950 & ~n17143;
  assign n17145 = pi36  & ~n17144;
  assign n17146 = ~pi36  & ~n17143;
  assign n17147 = ~pi36  & n17144;
  assign n17148 = ~n33950 & n17146;
  assign n17149 = ~n17145 & ~n33951;
  assign n17150 = pi34  & ~n17001;
  assign n17151 = ~pi32  & ~pi33 ;
  assign n17152 = ~pi34  & n17151;
  assign n17153 = ~n33749 & ~n33833;
  assign n17154 = ~n15565 & n17153;
  assign n17155 = ~n15584 & n17154;
  assign n17156 = ~n33751 & n17155;
  assign n17157 = n15570 & n15586;
  assign n17158 = ~n15578 & n17156;
  assign n17159 = ~n17152 & ~n33952;
  assign n17160 = ~n16246 & n17159;
  assign n17161 = ~n33831 & n17160;
  assign n17162 = ~n16240 & n17161;
  assign n17163 = ~n17150 & ~n17152;
  assign n17164 = n16248 & n17163;
  assign n17165 = ~n17150 & n17162;
  assign n17166 = pi35  & ~n17138;
  assign n17167 = ~n33950 & ~n17166;
  assign n17168 = ~n33953 & n17167;
  assign n17169 = ~n16248 & ~n17163;
  assign n17170 = n15586 & ~n17169;
  assign n17171 = ~n17168 & ~n17169;
  assign n17172 = n15586 & n17171;
  assign n17173 = ~n17168 & n17170;
  assign n17174 = ~n17149 & ~n33954;
  assign n17175 = ~n15586 & ~n17171;
  assign n17176 = n14866 & ~n17175;
  assign n17177 = ~n17174 & n17176;
  assign n17178 = ~n16253 & ~n33834;
  assign n17179 = ~n17001 & n17178;
  assign n17180 = n16258 & ~n17179;
  assign n17181 = ~n16258 & n17178;
  assign n17182 = ~n16258 & n17179;
  assign n17183 = ~n17001 & n17181;
  assign n17184 = ~n17180 & ~n33955;
  assign n17185 = ~n17177 & ~n17184;
  assign n17186 = ~n17174 & ~n17175;
  assign n17187 = ~n14866 & ~n17186;
  assign n17188 = n14233 & ~n17187;
  assign n17189 = ~n17185 & ~n17187;
  assign n17190 = n14233 & n17189;
  assign n17191 = ~n17185 & n17188;
  assign n17192 = ~n17137 & ~n33956;
  assign n17193 = ~n14233 & ~n17189;
  assign n17194 = n13548 & ~n17193;
  assign n17195 = ~n17192 & n17194;
  assign n17196 = ~n16287 & ~n33836;
  assign n17197 = ~n17001 & n17196;
  assign n17198 = ~n16297 & ~n17197;
  assign n17199 = ~n16287 & n16297;
  assign n17200 = ~n33836 & n17199;
  assign n17201 = n16297 & n17197;
  assign n17202 = ~n17001 & n17200;
  assign n17203 = n16297 & ~n17197;
  assign n17204 = ~n16297 & n17197;
  assign n17205 = ~n17203 & ~n17204;
  assign n17206 = ~n17198 & ~n33957;
  assign n17207 = ~n17195 & n33958;
  assign n17208 = ~n17192 & ~n17193;
  assign n17209 = ~n13548 & ~n17208;
  assign n17210 = n12948 & ~n17209;
  assign n17211 = ~n17207 & ~n17209;
  assign n17212 = n12948 & n17211;
  assign n17213 = ~n17207 & n17210;
  assign n17214 = ~n17129 & ~n33959;
  assign n17215 = ~n12948 & ~n17211;
  assign n17216 = n12296 & ~n17215;
  assign n17217 = ~n17214 & n17216;
  assign n17218 = ~n16317 & ~n33840;
  assign n17219 = ~n17001 & n17218;
  assign n17220 = ~n33842 & ~n17219;
  assign n17221 = n33842 & n17219;
  assign n17222 = ~n16317 & ~n33842;
  assign n17223 = ~n33840 & n17222;
  assign n17224 = ~n17001 & n17223;
  assign n17225 = n33842 & ~n17219;
  assign n17226 = ~n17224 & ~n17225;
  assign n17227 = ~n17220 & ~n17221;
  assign n17228 = ~n17217 & ~n33960;
  assign n17229 = ~n17214 & ~n17215;
  assign n17230 = ~n12296 & ~n17229;
  assign n17231 = n11719 & ~n17230;
  assign n17232 = ~n17228 & ~n17230;
  assign n17233 = n11719 & n17232;
  assign n17234 = ~n17228 & n17231;
  assign n17235 = ~n17121 & ~n33961;
  assign n17236 = ~n11719 & ~n17232;
  assign n17237 = n11097 & ~n17236;
  assign n17238 = ~n17235 & n17237;
  assign n17239 = ~n16351 & ~n33845;
  assign n17240 = ~n17001 & n17239;
  assign n17241 = ~n33846 & n17240;
  assign n17242 = n33846 & ~n17240;
  assign n17243 = ~n16351 & n33846;
  assign n17244 = ~n33845 & n17243;
  assign n17245 = ~n17001 & n17244;
  assign n17246 = ~n33846 & ~n17240;
  assign n17247 = ~n17245 & ~n17246;
  assign n17248 = ~n17241 & ~n17242;
  assign n17249 = ~n17238 & ~n33962;
  assign n17250 = ~n17235 & ~n17236;
  assign n17251 = ~n11097 & ~n17250;
  assign n17252 = n10555 & ~n17251;
  assign n17253 = ~n17249 & ~n17251;
  assign n17254 = n10555 & n17253;
  assign n17255 = ~n17249 & n17252;
  assign n17256 = ~n17113 & ~n33963;
  assign n17257 = ~n10555 & ~n17253;
  assign n17258 = n9969 & ~n17257;
  assign n17259 = ~n17256 & n17258;
  assign n17260 = ~n16384 & ~n33849;
  assign n17261 = ~n17001 & n17260;
  assign n17262 = ~n33850 & n17261;
  assign n17263 = n33850 & ~n17261;
  assign n17264 = ~n33850 & ~n17261;
  assign n17265 = ~n16384 & n33850;
  assign n17266 = ~n33849 & n17265;
  assign n17267 = n33850 & n17261;
  assign n17268 = ~n17001 & n17266;
  assign n17269 = ~n17264 & ~n33964;
  assign n17270 = ~n17262 & ~n17263;
  assign n17271 = ~n17259 & ~n33965;
  assign n17272 = ~n17256 & ~n17257;
  assign n17273 = ~n9969 & ~n17272;
  assign n17274 = n9457 & ~n17273;
  assign n17275 = ~n17271 & ~n17273;
  assign n17276 = n9457 & n17275;
  assign n17277 = ~n17271 & n17274;
  assign n17278 = ~n17105 & ~n33966;
  assign n17279 = ~n9457 & ~n17275;
  assign n17280 = n8896 & ~n17279;
  assign n17281 = ~n17278 & n17280;
  assign n17282 = ~n16417 & ~n33853;
  assign n17283 = ~n16417 & ~n17001;
  assign n17284 = ~n33853 & n17283;
  assign n17285 = ~n17001 & n17282;
  assign n17286 = n33855 & ~n33967;
  assign n17287 = n16432 & n17283;
  assign n17288 = ~n33855 & n33967;
  assign n17289 = ~n16417 & n33855;
  assign n17290 = ~n33853 & n17289;
  assign n17291 = ~n17001 & n17290;
  assign n17292 = ~n33855 & ~n33967;
  assign n17293 = ~n17291 & ~n17292;
  assign n17294 = ~n17286 & ~n33968;
  assign n17295 = ~n17281 & ~n33969;
  assign n17296 = ~n17278 & ~n17279;
  assign n17297 = ~n8896 & ~n17296;
  assign n17298 = n8411 & ~n17297;
  assign n17299 = ~n17295 & ~n17297;
  assign n17300 = n8411 & n17299;
  assign n17301 = ~n17295 & n17298;
  assign n17302 = ~n17097 & ~n33970;
  assign n17303 = ~n8411 & ~n17299;
  assign n17304 = n7885 & ~n17303;
  assign n17305 = ~n17302 & n17304;
  assign n17306 = ~n17089 & ~n17305;
  assign n17307 = ~n17302 & ~n17303;
  assign n17308 = ~n7885 & ~n17307;
  assign n17309 = n7428 & ~n17308;
  assign n17310 = ~n17306 & ~n17308;
  assign n17311 = n7428 & n17310;
  assign n17312 = ~n17306 & n17309;
  assign n17313 = ~n17081 & ~n33971;
  assign n17314 = ~n7428 & ~n17310;
  assign n17315 = n6937 & ~n17314;
  assign n17316 = ~n17313 & n17315;
  assign n17317 = ~n16487 & ~n33865;
  assign n17318 = ~n16487 & ~n17001;
  assign n17319 = ~n33865 & n17318;
  assign n17320 = ~n17001 & n17317;
  assign n17321 = n16495 & ~n33972;
  assign n17322 = n16499 & n17318;
  assign n17323 = ~n16487 & n16495;
  assign n17324 = ~n33865 & n17323;
  assign n17325 = ~n17001 & n17324;
  assign n17326 = ~n16495 & ~n33972;
  assign n17327 = ~n17325 & ~n17326;
  assign n17328 = ~n17321 & ~n17322;
  assign n17329 = ~n17316 & ~n33973;
  assign n17330 = ~n17313 & ~n17314;
  assign n17331 = ~n6937 & ~n17330;
  assign n17332 = n6507 & ~n17331;
  assign n17333 = ~n17329 & ~n17331;
  assign n17334 = n6507 & n17333;
  assign n17335 = ~n17329 & n17332;
  assign n17336 = ~n17073 & ~n33974;
  assign n17337 = ~n6507 & ~n17333;
  assign n17338 = n6051 & ~n17337;
  assign n17339 = ~n17336 & n17338;
  assign n17340 = ~n17065 & ~n17339;
  assign n17341 = ~n17336 & ~n17337;
  assign n17342 = ~n6051 & ~n17341;
  assign n17343 = n5648 & ~n17342;
  assign n17344 = ~n17340 & ~n17342;
  assign n17345 = n5648 & n17344;
  assign n17346 = ~n17340 & n17343;
  assign n17347 = ~n17057 & ~n33975;
  assign n17348 = ~n5648 & ~n17344;
  assign n17349 = n5223 & ~n17348;
  assign n17350 = ~n17347 & n17349;
  assign n17351 = ~n16553 & ~n33874;
  assign n17352 = ~n16553 & ~n17001;
  assign n17353 = ~n33874 & n17352;
  assign n17354 = ~n17001 & n17351;
  assign n17355 = n16561 & ~n33976;
  assign n17356 = n16565 & n17352;
  assign n17357 = ~n16553 & n16561;
  assign n17358 = ~n33874 & n17357;
  assign n17359 = ~n17001 & n17358;
  assign n17360 = ~n16561 & ~n33976;
  assign n17361 = ~n17359 & ~n17360;
  assign n17362 = ~n17355 & ~n17356;
  assign n17363 = ~n17350 & ~n33977;
  assign n17364 = ~n17347 & ~n17348;
  assign n17365 = ~n5223 & ~n17364;
  assign n17366 = n4851 & ~n17365;
  assign n17367 = ~n17363 & ~n17365;
  assign n17368 = n4851 & n17367;
  assign n17369 = ~n17363 & n17366;
  assign n17370 = ~n17049 & ~n33978;
  assign n17371 = ~n4851 & ~n17367;
  assign n17372 = n4461 & ~n17371;
  assign n17373 = ~n17370 & n17372;
  assign n17374 = ~n17041 & ~n17373;
  assign n17375 = ~n17370 & ~n17371;
  assign n17376 = ~n4461 & ~n17375;
  assign n17377 = n4115 & ~n17376;
  assign n17378 = ~n17374 & ~n17376;
  assign n17379 = n4115 & n17378;
  assign n17380 = ~n17374 & n17377;
  assign n17381 = ~n17033 & ~n33979;
  assign n17382 = ~n4115 & ~n17378;
  assign n17383 = n3754 & ~n17382;
  assign n17384 = ~n17381 & n17383;
  assign n17385 = ~n16619 & ~n33883;
  assign n17386 = ~n16619 & ~n17001;
  assign n17387 = ~n33883 & n17386;
  assign n17388 = ~n17001 & n17385;
  assign n17389 = n16627 & ~n33980;
  assign n17390 = n16631 & n17386;
  assign n17391 = ~n16619 & n16627;
  assign n17392 = ~n33883 & n17391;
  assign n17393 = ~n17001 & n17392;
  assign n17394 = ~n16627 & ~n33980;
  assign n17395 = ~n17393 & ~n17394;
  assign n17396 = ~n17389 & ~n17390;
  assign n17397 = ~n17384 & ~n33981;
  assign n17398 = ~n17381 & ~n17382;
  assign n17399 = ~n3754 & ~n17398;
  assign n17400 = n3444 & ~n17399;
  assign n17401 = ~n17397 & ~n17399;
  assign n17402 = n3444 & n17401;
  assign n17403 = ~n17397 & n17400;
  assign n17404 = ~n17025 & ~n33982;
  assign n17405 = ~n3444 & ~n17401;
  assign n17406 = n3116 & ~n17405;
  assign n17407 = ~n17404 & n17406;
  assign n17408 = ~n17017 & ~n17407;
  assign n17409 = ~n17404 & ~n17405;
  assign n17410 = ~n3116 & ~n17409;
  assign n17411 = n2833 & ~n17410;
  assign n17412 = ~n17408 & ~n17410;
  assign n17413 = n2833 & n17412;
  assign n17414 = ~n17408 & n17411;
  assign n17415 = ~n17009 & ~n33983;
  assign n17416 = ~n2833 & ~n17412;
  assign n17417 = ~n17415 & ~n17416;
  assign n17418 = ~n2536 & ~n17417;
  assign n17419 = ~n16683 & n16691;
  assign n17420 = ~n33891 & n17419;
  assign n17421 = ~n16683 & ~n33891;
  assign n17422 = ~n17001 & n17421;
  assign n17423 = n16691 & n17422;
  assign n17424 = ~n17001 & n17420;
  assign n17425 = ~n16691 & ~n17422;
  assign n17426 = ~n33984 & ~n17425;
  assign n17427 = n2536 & ~n17416;
  assign n17428 = ~n17415 & n17427;
  assign n17429 = ~n17426 & ~n17428;
  assign n17430 = ~n17418 & ~n17429;
  assign n17431 = ~n2283 & ~n17430;
  assign n17432 = ~n16697 & ~n16699;
  assign n17433 = ~n17001 & n17432;
  assign n17434 = ~n33893 & ~n17433;
  assign n17435 = ~n16699 & n33893;
  assign n17436 = ~n16697 & n17435;
  assign n17437 = n33893 & n17433;
  assign n17438 = ~n17001 & n17436;
  assign n17439 = ~n17434 & ~n33985;
  assign n17440 = n2283 & ~n17418;
  assign n17441 = n2283 & n17430;
  assign n17442 = ~n17429 & n17440;
  assign n17443 = ~n17439 & ~n33986;
  assign n17444 = ~n17431 & ~n17443;
  assign n17445 = ~n2021 & ~n17444;
  assign n17446 = n2021 & ~n17431;
  assign n17447 = ~n17443 & n17446;
  assign n17448 = ~n16714 & ~n33895;
  assign n17449 = ~n16714 & ~n17001;
  assign n17450 = ~n33895 & n17449;
  assign n17451 = ~n17001 & n17448;
  assign n17452 = n16722 & ~n33987;
  assign n17453 = n16726 & n17449;
  assign n17454 = ~n16714 & n16722;
  assign n17455 = ~n33895 & n17454;
  assign n17456 = ~n17001 & n17455;
  assign n17457 = ~n16722 & ~n33987;
  assign n17458 = ~n17456 & ~n17457;
  assign n17459 = ~n17452 & ~n17453;
  assign n17460 = ~n17447 & ~n33988;
  assign n17461 = ~n17445 & ~n17460;
  assign n17462 = ~n1796 & ~n17461;
  assign n17463 = ~n16728 & ~n16730;
  assign n17464 = ~n17001 & n17463;
  assign n17465 = ~n33897 & ~n17464;
  assign n17466 = ~n16730 & n33897;
  assign n17467 = ~n16728 & n17466;
  assign n17468 = n33897 & n17464;
  assign n17469 = ~n17001 & n17467;
  assign n17470 = ~n17465 & ~n33989;
  assign n17471 = n1796 & ~n17445;
  assign n17472 = n1796 & n17461;
  assign n17473 = ~n17460 & n17471;
  assign n17474 = ~n17470 & ~n33990;
  assign n17475 = ~n17462 & ~n17474;
  assign n17476 = ~n1567 & ~n17475;
  assign n17477 = n1567 & ~n17462;
  assign n17478 = ~n17474 & n17477;
  assign n17479 = ~n16745 & ~n33899;
  assign n17480 = ~n16745 & ~n17001;
  assign n17481 = ~n33899 & n17480;
  assign n17482 = ~n17001 & n17479;
  assign n17483 = n16753 & ~n33991;
  assign n17484 = n16757 & n17480;
  assign n17485 = ~n16745 & n16753;
  assign n17486 = ~n33899 & n17485;
  assign n17487 = ~n17001 & n17486;
  assign n17488 = ~n16753 & ~n33991;
  assign n17489 = ~n17487 & ~n17488;
  assign n17490 = ~n17483 & ~n17484;
  assign n17491 = ~n17478 & ~n33992;
  assign n17492 = ~n17476 & ~n17491;
  assign n17493 = ~n1374 & ~n17492;
  assign n17494 = ~n16759 & ~n16761;
  assign n17495 = ~n17001 & n17494;
  assign n17496 = ~n33901 & ~n17495;
  assign n17497 = ~n16761 & n33901;
  assign n17498 = ~n16759 & n17497;
  assign n17499 = n33901 & n17495;
  assign n17500 = ~n17001 & n17498;
  assign n17501 = ~n17496 & ~n33993;
  assign n17502 = n1374 & ~n17476;
  assign n17503 = n1374 & n17492;
  assign n17504 = ~n17491 & n17502;
  assign n17505 = ~n17501 & ~n33994;
  assign n17506 = ~n17493 & ~n17505;
  assign n17507 = ~n1179 & ~n17506;
  assign n17508 = ~n16776 & ~n33902;
  assign n17509 = ~n17001 & n17508;
  assign n17510 = ~n33904 & ~n17509;
  assign n17511 = ~n16776 & n33904;
  assign n17512 = ~n33902 & n17511;
  assign n17513 = n33904 & n17509;
  assign n17514 = ~n17001 & n17512;
  assign n17515 = ~n17510 & ~n33995;
  assign n17516 = n1179 & ~n17493;
  assign n17517 = ~n17505 & n17516;
  assign n17518 = ~n17515 & ~n17517;
  assign n17519 = ~n17507 & ~n17518;
  assign n17520 = ~n1016 & ~n17519;
  assign n17521 = ~n16794 & ~n16796;
  assign n17522 = ~n17001 & n17521;
  assign n17523 = ~n33906 & ~n17522;
  assign n17524 = ~n16796 & n33906;
  assign n17525 = ~n16794 & n17524;
  assign n17526 = n33906 & n17522;
  assign n17527 = ~n17001 & n17525;
  assign n17528 = ~n17523 & ~n33996;
  assign n17529 = n1016 & ~n17507;
  assign n17530 = n1016 & n17519;
  assign n17531 = ~n17518 & n17529;
  assign n17532 = ~n17528 & ~n33997;
  assign n17533 = ~n17520 & ~n17532;
  assign n17534 = ~n855 & ~n17533;
  assign n17535 = n855 & ~n17520;
  assign n17536 = ~n17532 & n17535;
  assign n17537 = ~n16811 & ~n33908;
  assign n17538 = ~n16811 & ~n17001;
  assign n17539 = ~n33908 & n17538;
  assign n17540 = ~n17001 & n17537;
  assign n17541 = n16819 & ~n33998;
  assign n17542 = n16823 & n17538;
  assign n17543 = ~n16811 & n16819;
  assign n17544 = ~n33908 & n17543;
  assign n17545 = ~n17001 & n17544;
  assign n17546 = ~n16819 & ~n33998;
  assign n17547 = ~n17545 & ~n17546;
  assign n17548 = ~n17541 & ~n17542;
  assign n17549 = ~n17536 & ~n33999;
  assign n17550 = ~n17534 & ~n17549;
  assign n17551 = ~n720 & ~n17550;
  assign n17552 = ~n16825 & ~n16827;
  assign n17553 = ~n17001 & n17552;
  assign n17554 = ~n33910 & ~n17553;
  assign n17555 = ~n16827 & n33910;
  assign n17556 = ~n16825 & n17555;
  assign n17557 = n33910 & n17553;
  assign n17558 = ~n17001 & n17556;
  assign n17559 = ~n17554 & ~n34000;
  assign n17560 = n720 & ~n17534;
  assign n17561 = n720 & n17550;
  assign n17562 = ~n17549 & n17560;
  assign n17563 = ~n17559 & ~n34001;
  assign n17564 = ~n17551 & ~n17563;
  assign n17565 = ~n592 & ~n17564;
  assign n17566 = ~n16842 & ~n33911;
  assign n17567 = ~n17001 & n17566;
  assign n17568 = ~n33913 & ~n17567;
  assign n17569 = ~n16842 & n33913;
  assign n17570 = ~n33911 & n17569;
  assign n17571 = n33913 & n17567;
  assign n17572 = ~n17001 & n17570;
  assign n17573 = ~n17568 & ~n34002;
  assign n17574 = n592 & ~n17551;
  assign n17575 = ~n17563 & n17574;
  assign n17576 = ~n17573 & ~n17575;
  assign n17577 = ~n17565 & ~n17576;
  assign n17578 = ~n487 & ~n17577;
  assign n17579 = ~n16860 & ~n16862;
  assign n17580 = ~n17001 & n17579;
  assign n17581 = ~n33915 & ~n17580;
  assign n17582 = ~n16862 & n33915;
  assign n17583 = ~n16860 & n17582;
  assign n17584 = n33915 & n17580;
  assign n17585 = ~n17001 & n17583;
  assign n17586 = ~n17581 & ~n34003;
  assign n17587 = n487 & ~n17565;
  assign n17588 = n487 & n17577;
  assign n17589 = ~n17576 & n17587;
  assign n17590 = ~n17586 & ~n34004;
  assign n17591 = ~n17578 & ~n17590;
  assign n17592 = ~n393 & ~n17591;
  assign n17593 = n393 & ~n17578;
  assign n17594 = ~n17590 & n17593;
  assign n17595 = ~n16877 & ~n33917;
  assign n17596 = ~n16877 & ~n17001;
  assign n17597 = ~n33917 & n17596;
  assign n17598 = ~n17001 & n17595;
  assign n17599 = n16885 & ~n34005;
  assign n17600 = n16889 & n17596;
  assign n17601 = ~n16877 & n16885;
  assign n17602 = ~n33917 & n17601;
  assign n17603 = ~n17001 & n17602;
  assign n17604 = ~n16885 & ~n34005;
  assign n17605 = ~n17603 & ~n17604;
  assign n17606 = ~n17599 & ~n17600;
  assign n17607 = ~n17594 & ~n34006;
  assign n17608 = ~n17592 & ~n17607;
  assign n17609 = ~n321 & ~n17608;
  assign n17610 = ~n16891 & ~n16893;
  assign n17611 = ~n17001 & n17610;
  assign n17612 = ~n33919 & ~n17611;
  assign n17613 = ~n16893 & n33919;
  assign n17614 = ~n16891 & n17613;
  assign n17615 = n33919 & n17611;
  assign n17616 = ~n17001 & n17614;
  assign n17617 = ~n17612 & ~n34007;
  assign n17618 = n321 & ~n17592;
  assign n17619 = n321 & n17608;
  assign n17620 = ~n17607 & n17618;
  assign n17621 = ~n17617 & ~n34008;
  assign n17622 = ~n17609 & ~n17621;
  assign n17623 = ~n263 & ~n17622;
  assign n17624 = ~n16908 & ~n33920;
  assign n17625 = ~n17001 & n17624;
  assign n17626 = ~n33922 & ~n17625;
  assign n17627 = ~n16908 & n33922;
  assign n17628 = ~n33920 & n17627;
  assign n17629 = n33922 & n17625;
  assign n17630 = ~n17001 & n17628;
  assign n17631 = ~n17626 & ~n34009;
  assign n17632 = n263 & ~n17609;
  assign n17633 = ~n17621 & n17632;
  assign n17634 = ~n17631 & ~n17633;
  assign n17635 = ~n17623 & ~n17634;
  assign n17636 = ~n214 & ~n17635;
  assign n17637 = ~n16926 & ~n16928;
  assign n17638 = ~n17001 & n17637;
  assign n17639 = ~n33924 & ~n17638;
  assign n17640 = ~n16928 & n33924;
  assign n17641 = ~n16926 & n17640;
  assign n17642 = n33924 & n17638;
  assign n17643 = ~n17001 & n17641;
  assign n17644 = ~n17639 & ~n34010;
  assign n17645 = n214 & ~n17623;
  assign n17646 = n214 & n17635;
  assign n17647 = ~n17634 & n17645;
  assign n17648 = ~n17644 & ~n34011;
  assign n17649 = ~n17636 & ~n17648;
  assign n17650 = ~n197 & ~n17649;
  assign n17651 = n197 & ~n17636;
  assign n17652 = ~n17648 & n17651;
  assign n17653 = ~n16943 & ~n33926;
  assign n17654 = ~n16943 & ~n17001;
  assign n17655 = ~n33926 & n17654;
  assign n17656 = ~n17001 & n17653;
  assign n17657 = n16951 & ~n34012;
  assign n17658 = n16955 & n17654;
  assign n17659 = ~n16943 & n16951;
  assign n17660 = ~n33926 & n17659;
  assign n17661 = ~n17001 & n17660;
  assign n17662 = ~n16951 & ~n34012;
  assign n17663 = ~n17661 & ~n17662;
  assign n17664 = ~n17657 & ~n17658;
  assign n17665 = ~n17652 & ~n34013;
  assign n17666 = ~n17650 & ~n17665;
  assign n17667 = ~n16957 & ~n16959;
  assign n17668 = ~n17001 & n17667;
  assign n17669 = ~n33928 & ~n17668;
  assign n17670 = ~n16959 & n33928;
  assign n17671 = ~n16957 & n17670;
  assign n17672 = n33928 & n17668;
  assign n17673 = ~n17001 & n17671;
  assign n17674 = ~n17669 & ~n34014;
  assign n17675 = ~n16973 & ~n33930;
  assign n17676 = ~n33930 & ~n17001;
  assign n17677 = ~n16973 & n17676;
  assign n17678 = ~n17001 & n17675;
  assign n17679 = ~n33932 & ~n34015;
  assign n17680 = ~n17674 & n17679;
  assign n17681 = ~n17666 & n17680;
  assign n17682 = n193 & ~n17681;
  assign n17683 = ~n17650 & n17674;
  assign n17684 = n17666 & n17674;
  assign n17685 = ~n17665 & n17683;
  assign n17686 = n16973 & ~n17676;
  assign n17687 = ~n193 & ~n17675;
  assign n17688 = ~n17686 & n17687;
  assign n17689 = ~n34016 & ~n17688;
  assign n17690 = ~n17682 & n17689;
  assign n17691 = pi32  & ~n17690;
  assign n17692 = ~pi30  & ~pi31 ;
  assign n17693 = ~pi32  & n17692;
  assign n17694 = ~n17691 & ~n17693;
  assign n17695 = ~n17001 & ~n17694;
  assign n17696 = ~pi32  & ~n17690;
  assign n17697 = pi33  & ~n17696;
  assign n17698 = ~pi33  & n17696;
  assign n17699 = n17151 & ~n17690;
  assign n17700 = ~n17697 & ~n34017;
  assign n17701 = ~n33829 & ~n33952;
  assign n17702 = ~n16227 & n17701;
  assign n17703 = ~n16246 & n17702;
  assign n17704 = ~n33831 & n17703;
  assign n17705 = n16232 & n16248;
  assign n17706 = ~n16240 & n17704;
  assign n17707 = ~n17693 & ~n34018;
  assign n17708 = ~n16999 & n17707;
  assign n17709 = ~n33932 & n17708;
  assign n17710 = ~n16993 & n17709;
  assign n17711 = n17001 & n17694;
  assign n17712 = ~n17691 & n17710;
  assign n17713 = n17700 & ~n34019;
  assign n17714 = ~n17695 & ~n17713;
  assign n17715 = ~n16248 & ~n17714;
  assign n17716 = n16248 & ~n17695;
  assign n17717 = ~n17713 & n17716;
  assign n17718 = ~n17001 & ~n17688;
  assign n17719 = ~n34016 & n17718;
  assign n17720 = ~n17682 & n17719;
  assign n17721 = ~n34017 & ~n17720;
  assign n17722 = pi34  & ~n17721;
  assign n17723 = ~pi34  & ~n17720;
  assign n17724 = ~pi34  & n17721;
  assign n17725 = ~n34017 & n17723;
  assign n17726 = ~n17722 & ~n34020;
  assign n17727 = ~n17717 & ~n17726;
  assign n17728 = ~n17715 & ~n17727;
  assign n17729 = ~n15586 & ~n17728;
  assign n17730 = n15586 & ~n17715;
  assign n17731 = ~n17727 & n17730;
  assign n17732 = n15586 & n17728;
  assign n17733 = ~n33953 & ~n17169;
  assign n17734 = ~n17690 & n17733;
  assign n17735 = n17167 & ~n17734;
  assign n17736 = ~n17167 & n17733;
  assign n17737 = ~n17167 & n17734;
  assign n17738 = ~n17690 & n17736;
  assign n17739 = ~n17735 & ~n34022;
  assign n17740 = ~n34021 & ~n17739;
  assign n17741 = ~n17729 & ~n17740;
  assign n17742 = ~n14866 & ~n17741;
  assign n17743 = n14866 & ~n17729;
  assign n17744 = ~n17740 & n17743;
  assign n17745 = ~n33954 & ~n17175;
  assign n17746 = ~n17175 & ~n17690;
  assign n17747 = ~n33954 & n17746;
  assign n17748 = ~n17690 & n17745;
  assign n17749 = n17149 & ~n34023;
  assign n17750 = n17174 & n17746;
  assign n17751 = n17149 & ~n33954;
  assign n17752 = ~n17175 & n17751;
  assign n17753 = ~n17690 & n17752;
  assign n17754 = ~n17149 & ~n34023;
  assign n17755 = ~n17753 & ~n17754;
  assign n17756 = ~n17749 & ~n17750;
  assign n17757 = ~n17744 & ~n34024;
  assign n17758 = ~n17742 & ~n17757;
  assign n17759 = ~n14233 & ~n17758;
  assign n17760 = n14233 & ~n17742;
  assign n17761 = ~n17757 & n17760;
  assign n17762 = n14233 & n17758;
  assign n17763 = ~n17177 & ~n17187;
  assign n17764 = ~n17690 & n17763;
  assign n17765 = ~n17184 & ~n17764;
  assign n17766 = n17184 & ~n17187;
  assign n17767 = ~n17177 & n17766;
  assign n17768 = n17184 & n17764;
  assign n17769 = ~n17690 & n17767;
  assign n17770 = n17184 & ~n17764;
  assign n17771 = ~n17184 & n17764;
  assign n17772 = ~n17770 & ~n17771;
  assign n17773 = ~n17765 & ~n34026;
  assign n17774 = ~n34025 & n34027;
  assign n17775 = ~n17759 & ~n17774;
  assign n17776 = ~n13548 & ~n17775;
  assign n17777 = n13548 & ~n17759;
  assign n17778 = ~n17774 & n17777;
  assign n17779 = ~n33956 & ~n17193;
  assign n17780 = ~n17193 & ~n17690;
  assign n17781 = ~n33956 & n17780;
  assign n17782 = ~n17690 & n17779;
  assign n17783 = n17137 & ~n34028;
  assign n17784 = n17192 & n17780;
  assign n17785 = n17137 & ~n33956;
  assign n17786 = ~n17193 & n17785;
  assign n17787 = ~n17690 & n17786;
  assign n17788 = ~n17137 & ~n34028;
  assign n17789 = ~n17787 & ~n17788;
  assign n17790 = ~n17783 & ~n17784;
  assign n17791 = ~n17778 & ~n34029;
  assign n17792 = ~n17776 & ~n17791;
  assign n17793 = ~n12948 & ~n17792;
  assign n17794 = n12948 & ~n17776;
  assign n17795 = ~n17791 & n17794;
  assign n17796 = n12948 & n17792;
  assign n17797 = ~n17195 & ~n17209;
  assign n17798 = ~n17690 & n17797;
  assign n17799 = ~n33958 & ~n17798;
  assign n17800 = n33958 & n17798;
  assign n17801 = ~n33958 & ~n17209;
  assign n17802 = ~n17195 & n17801;
  assign n17803 = ~n17690 & n17802;
  assign n17804 = n33958 & ~n17798;
  assign n17805 = ~n17803 & ~n17804;
  assign n17806 = ~n17799 & ~n17800;
  assign n17807 = ~n34030 & ~n34031;
  assign n17808 = ~n17793 & ~n17807;
  assign n17809 = ~n12296 & ~n17808;
  assign n17810 = n12296 & ~n17793;
  assign n17811 = ~n17807 & n17810;
  assign n17812 = ~n33959 & ~n17215;
  assign n17813 = ~n17215 & ~n17690;
  assign n17814 = ~n33959 & n17813;
  assign n17815 = ~n17690 & n17812;
  assign n17816 = n17129 & ~n34032;
  assign n17817 = n17214 & n17813;
  assign n17818 = n17129 & ~n33959;
  assign n17819 = ~n17215 & n17818;
  assign n17820 = ~n17690 & n17819;
  assign n17821 = ~n17129 & ~n34032;
  assign n17822 = ~n17820 & ~n17821;
  assign n17823 = ~n17816 & ~n17817;
  assign n17824 = ~n17811 & ~n34033;
  assign n17825 = ~n17809 & ~n17824;
  assign n17826 = ~n11719 & ~n17825;
  assign n17827 = n11719 & ~n17809;
  assign n17828 = ~n17824 & n17827;
  assign n17829 = n11719 & n17825;
  assign n17830 = ~n17217 & ~n17230;
  assign n17831 = ~n17690 & n17830;
  assign n17832 = ~n33960 & n17831;
  assign n17833 = n33960 & ~n17831;
  assign n17834 = n33960 & ~n17230;
  assign n17835 = ~n17217 & n17834;
  assign n17836 = ~n17690 & n17835;
  assign n17837 = ~n33960 & ~n17831;
  assign n17838 = ~n17836 & ~n17837;
  assign n17839 = ~n17832 & ~n17833;
  assign n17840 = ~n34034 & ~n34035;
  assign n17841 = ~n17826 & ~n17840;
  assign n17842 = ~n11097 & ~n17841;
  assign n17843 = n11097 & ~n17826;
  assign n17844 = ~n17840 & n17843;
  assign n17845 = ~n33961 & ~n17236;
  assign n17846 = ~n17236 & ~n17690;
  assign n17847 = ~n33961 & n17846;
  assign n17848 = ~n17690 & n17845;
  assign n17849 = n17121 & ~n34036;
  assign n17850 = n17235 & n17846;
  assign n17851 = n17121 & ~n33961;
  assign n17852 = ~n17236 & n17851;
  assign n17853 = ~n17690 & n17852;
  assign n17854 = ~n17121 & ~n34036;
  assign n17855 = ~n17853 & ~n17854;
  assign n17856 = ~n17849 & ~n17850;
  assign n17857 = ~n17844 & ~n34037;
  assign n17858 = ~n17842 & ~n17857;
  assign n17859 = ~n10555 & ~n17858;
  assign n17860 = n10555 & ~n17842;
  assign n17861 = ~n17857 & n17860;
  assign n17862 = n10555 & n17858;
  assign n17863 = ~n17238 & ~n17251;
  assign n17864 = ~n17690 & n17863;
  assign n17865 = ~n33962 & n17864;
  assign n17866 = n33962 & ~n17864;
  assign n17867 = ~n33962 & ~n17864;
  assign n17868 = n33962 & ~n17251;
  assign n17869 = ~n17238 & n17868;
  assign n17870 = n33962 & n17864;
  assign n17871 = ~n17690 & n17869;
  assign n17872 = ~n17867 & ~n34039;
  assign n17873 = ~n17865 & ~n17866;
  assign n17874 = ~n34038 & ~n34040;
  assign n17875 = ~n17859 & ~n17874;
  assign n17876 = ~n9969 & ~n17875;
  assign n17877 = n9969 & ~n17859;
  assign n17878 = ~n17874 & n17877;
  assign n17879 = ~n33963 & ~n17257;
  assign n17880 = ~n17257 & ~n17690;
  assign n17881 = ~n33963 & n17880;
  assign n17882 = ~n17690 & n17879;
  assign n17883 = n17113 & ~n34041;
  assign n17884 = n17256 & n17880;
  assign n17885 = n17113 & ~n33963;
  assign n17886 = ~n17257 & n17885;
  assign n17887 = ~n17690 & n17886;
  assign n17888 = ~n17113 & ~n34041;
  assign n17889 = ~n17887 & ~n17888;
  assign n17890 = ~n17883 & ~n17884;
  assign n17891 = ~n17878 & ~n34042;
  assign n17892 = ~n17876 & ~n17891;
  assign n17893 = ~n9457 & ~n17892;
  assign n17894 = n9457 & ~n17876;
  assign n17895 = ~n17891 & n17894;
  assign n17896 = n9457 & n17892;
  assign n17897 = ~n17259 & ~n17273;
  assign n17898 = ~n17273 & ~n17690;
  assign n17899 = ~n17259 & n17898;
  assign n17900 = ~n17690 & n17897;
  assign n17901 = n33965 & ~n34044;
  assign n17902 = n17271 & n17898;
  assign n17903 = ~n33965 & n34044;
  assign n17904 = n33965 & ~n17273;
  assign n17905 = ~n17259 & n17904;
  assign n17906 = ~n17690 & n17905;
  assign n17907 = ~n33965 & ~n34044;
  assign n17908 = ~n17906 & ~n17907;
  assign n17909 = ~n17901 & ~n34045;
  assign n17910 = ~n34043 & ~n34046;
  assign n17911 = ~n17893 & ~n17910;
  assign n17912 = ~n8896 & ~n17911;
  assign n17913 = n8896 & ~n17893;
  assign n17914 = ~n17910 & n17913;
  assign n17915 = ~n33966 & ~n17279;
  assign n17916 = ~n17279 & ~n17690;
  assign n17917 = ~n33966 & n17916;
  assign n17918 = ~n17690 & n17915;
  assign n17919 = n17105 & ~n34047;
  assign n17920 = n17278 & n17916;
  assign n17921 = n17105 & ~n33966;
  assign n17922 = ~n17279 & n17921;
  assign n17923 = ~n17690 & n17922;
  assign n17924 = ~n17105 & ~n34047;
  assign n17925 = ~n17923 & ~n17924;
  assign n17926 = ~n17919 & ~n17920;
  assign n17927 = ~n17914 & ~n34048;
  assign n17928 = ~n17912 & ~n17927;
  assign n17929 = ~n8411 & ~n17928;
  assign n17930 = ~n17281 & ~n17297;
  assign n17931 = ~n17690 & n17930;
  assign n17932 = ~n33969 & ~n17931;
  assign n17933 = n33969 & ~n17297;
  assign n17934 = ~n17281 & n17933;
  assign n17935 = n33969 & n17931;
  assign n17936 = ~n17690 & n17934;
  assign n17937 = ~n17932 & ~n34049;
  assign n17938 = n8411 & ~n17912;
  assign n17939 = ~n17927 & n17938;
  assign n17940 = n8411 & n17928;
  assign n17941 = ~n17937 & ~n34050;
  assign n17942 = ~n17929 & ~n17941;
  assign n17943 = ~n7885 & ~n17942;
  assign n17944 = n7885 & ~n17929;
  assign n17945 = ~n17941 & n17944;
  assign n17946 = ~n33970 & ~n17303;
  assign n17947 = ~n17303 & ~n17690;
  assign n17948 = ~n33970 & n17947;
  assign n17949 = ~n17690 & n17946;
  assign n17950 = n17097 & ~n34051;
  assign n17951 = n17302 & n17947;
  assign n17952 = n17097 & ~n33970;
  assign n17953 = ~n17303 & n17952;
  assign n17954 = ~n17690 & n17953;
  assign n17955 = ~n17097 & ~n34051;
  assign n17956 = ~n17954 & ~n17955;
  assign n17957 = ~n17950 & ~n17951;
  assign n17958 = ~n17945 & ~n34052;
  assign n17959 = ~n17943 & ~n17958;
  assign n17960 = ~n7428 & ~n17959;
  assign n17961 = n7428 & ~n17943;
  assign n17962 = ~n17958 & n17961;
  assign n17963 = n7428 & n17959;
  assign n17964 = ~n17305 & ~n17308;
  assign n17965 = ~n17308 & ~n17690;
  assign n17966 = ~n17305 & n17965;
  assign n17967 = ~n17690 & n17964;
  assign n17968 = n17089 & ~n34054;
  assign n17969 = n17306 & n17965;
  assign n17970 = n17089 & ~n17308;
  assign n17971 = ~n17305 & n17970;
  assign n17972 = ~n17690 & n17971;
  assign n17973 = ~n17089 & ~n34054;
  assign n17974 = ~n17972 & ~n17973;
  assign n17975 = ~n17968 & ~n17969;
  assign n17976 = ~n34053 & ~n34055;
  assign n17977 = ~n17960 & ~n17976;
  assign n17978 = ~n6937 & ~n17977;
  assign n17979 = n6937 & ~n17960;
  assign n17980 = ~n17976 & n17979;
  assign n17981 = ~n33971 & ~n17314;
  assign n17982 = ~n17314 & ~n17690;
  assign n17983 = ~n33971 & n17982;
  assign n17984 = ~n17690 & n17981;
  assign n17985 = n17081 & ~n34056;
  assign n17986 = n17313 & n17982;
  assign n17987 = n17081 & ~n33971;
  assign n17988 = ~n17314 & n17987;
  assign n17989 = ~n17690 & n17988;
  assign n17990 = ~n17081 & ~n34056;
  assign n17991 = ~n17989 & ~n17990;
  assign n17992 = ~n17985 & ~n17986;
  assign n17993 = ~n17980 & ~n34057;
  assign n17994 = ~n17978 & ~n17993;
  assign n17995 = ~n6507 & ~n17994;
  assign n17996 = ~n17316 & ~n17331;
  assign n17997 = ~n17690 & n17996;
  assign n17998 = ~n33973 & ~n17997;
  assign n17999 = n33973 & ~n17331;
  assign n18000 = ~n17316 & n17999;
  assign n18001 = n33973 & n17997;
  assign n18002 = ~n17690 & n18000;
  assign n18003 = ~n17998 & ~n34058;
  assign n18004 = n6507 & ~n17978;
  assign n18005 = ~n17993 & n18004;
  assign n18006 = n6507 & n17994;
  assign n18007 = ~n18003 & ~n34059;
  assign n18008 = ~n17995 & ~n18007;
  assign n18009 = ~n6051 & ~n18008;
  assign n18010 = n6051 & ~n17995;
  assign n18011 = ~n18007 & n18010;
  assign n18012 = ~n33974 & ~n17337;
  assign n18013 = ~n17337 & ~n17690;
  assign n18014 = ~n33974 & n18013;
  assign n18015 = ~n17690 & n18012;
  assign n18016 = n17073 & ~n34060;
  assign n18017 = n17336 & n18013;
  assign n18018 = n17073 & ~n33974;
  assign n18019 = ~n17337 & n18018;
  assign n18020 = ~n17690 & n18019;
  assign n18021 = ~n17073 & ~n34060;
  assign n18022 = ~n18020 & ~n18021;
  assign n18023 = ~n18016 & ~n18017;
  assign n18024 = ~n18011 & ~n34061;
  assign n18025 = ~n18009 & ~n18024;
  assign n18026 = ~n5648 & ~n18025;
  assign n18027 = n5648 & ~n18009;
  assign n18028 = ~n18024 & n18027;
  assign n18029 = n5648 & n18025;
  assign n18030 = ~n17339 & ~n17342;
  assign n18031 = ~n17342 & ~n17690;
  assign n18032 = ~n17339 & n18031;
  assign n18033 = ~n17690 & n18030;
  assign n18034 = n17065 & ~n34063;
  assign n18035 = n17340 & n18031;
  assign n18036 = n17065 & ~n17342;
  assign n18037 = ~n17339 & n18036;
  assign n18038 = ~n17690 & n18037;
  assign n18039 = ~n17065 & ~n34063;
  assign n18040 = ~n18038 & ~n18039;
  assign n18041 = ~n18034 & ~n18035;
  assign n18042 = ~n34062 & ~n34064;
  assign n18043 = ~n18026 & ~n18042;
  assign n18044 = ~n5223 & ~n18043;
  assign n18045 = n5223 & ~n18026;
  assign n18046 = ~n18042 & n18045;
  assign n18047 = ~n33975 & ~n17348;
  assign n18048 = ~n17348 & ~n17690;
  assign n18049 = ~n33975 & n18048;
  assign n18050 = ~n17690 & n18047;
  assign n18051 = n17057 & ~n34065;
  assign n18052 = n17347 & n18048;
  assign n18053 = n17057 & ~n33975;
  assign n18054 = ~n17348 & n18053;
  assign n18055 = ~n17690 & n18054;
  assign n18056 = ~n17057 & ~n34065;
  assign n18057 = ~n18055 & ~n18056;
  assign n18058 = ~n18051 & ~n18052;
  assign n18059 = ~n18046 & ~n34066;
  assign n18060 = ~n18044 & ~n18059;
  assign n18061 = ~n4851 & ~n18060;
  assign n18062 = ~n17350 & ~n17365;
  assign n18063 = ~n17690 & n18062;
  assign n18064 = ~n33977 & ~n18063;
  assign n18065 = n33977 & ~n17365;
  assign n18066 = ~n17350 & n18065;
  assign n18067 = n33977 & n18063;
  assign n18068 = ~n17690 & n18066;
  assign n18069 = ~n18064 & ~n34067;
  assign n18070 = n4851 & ~n18044;
  assign n18071 = ~n18059 & n18070;
  assign n18072 = n4851 & n18060;
  assign n18073 = ~n18069 & ~n34068;
  assign n18074 = ~n18061 & ~n18073;
  assign n18075 = ~n4461 & ~n18074;
  assign n18076 = n4461 & ~n18061;
  assign n18077 = ~n18073 & n18076;
  assign n18078 = ~n33978 & ~n17371;
  assign n18079 = ~n17371 & ~n17690;
  assign n18080 = ~n33978 & n18079;
  assign n18081 = ~n17690 & n18078;
  assign n18082 = n17049 & ~n34069;
  assign n18083 = n17370 & n18079;
  assign n18084 = n17049 & ~n33978;
  assign n18085 = ~n17371 & n18084;
  assign n18086 = ~n17690 & n18085;
  assign n18087 = ~n17049 & ~n34069;
  assign n18088 = ~n18086 & ~n18087;
  assign n18089 = ~n18082 & ~n18083;
  assign n18090 = ~n18077 & ~n34070;
  assign n18091 = ~n18075 & ~n18090;
  assign n18092 = ~n4115 & ~n18091;
  assign n18093 = n4115 & ~n18075;
  assign n18094 = ~n18090 & n18093;
  assign n18095 = n4115 & n18091;
  assign n18096 = ~n17373 & ~n17376;
  assign n18097 = ~n17376 & ~n17690;
  assign n18098 = ~n17373 & n18097;
  assign n18099 = ~n17690 & n18096;
  assign n18100 = n17041 & ~n34072;
  assign n18101 = n17374 & n18097;
  assign n18102 = n17041 & ~n17376;
  assign n18103 = ~n17373 & n18102;
  assign n18104 = ~n17690 & n18103;
  assign n18105 = ~n17041 & ~n34072;
  assign n18106 = ~n18104 & ~n18105;
  assign n18107 = ~n18100 & ~n18101;
  assign n18108 = ~n34071 & ~n34073;
  assign n18109 = ~n18092 & ~n18108;
  assign n18110 = ~n3754 & ~n18109;
  assign n18111 = n3754 & ~n18092;
  assign n18112 = ~n18108 & n18111;
  assign n18113 = ~n33979 & ~n17382;
  assign n18114 = ~n17382 & ~n17690;
  assign n18115 = ~n33979 & n18114;
  assign n18116 = ~n17690 & n18113;
  assign n18117 = n17033 & ~n34074;
  assign n18118 = n17381 & n18114;
  assign n18119 = n17033 & ~n33979;
  assign n18120 = ~n17382 & n18119;
  assign n18121 = ~n17690 & n18120;
  assign n18122 = ~n17033 & ~n34074;
  assign n18123 = ~n18121 & ~n18122;
  assign n18124 = ~n18117 & ~n18118;
  assign n18125 = ~n18112 & ~n34075;
  assign n18126 = ~n18110 & ~n18125;
  assign n18127 = ~n3444 & ~n18126;
  assign n18128 = ~n17384 & ~n17399;
  assign n18129 = ~n17690 & n18128;
  assign n18130 = ~n33981 & ~n18129;
  assign n18131 = n33981 & ~n17399;
  assign n18132 = ~n17384 & n18131;
  assign n18133 = n33981 & n18129;
  assign n18134 = ~n17690 & n18132;
  assign n18135 = ~n18130 & ~n34076;
  assign n18136 = n3444 & ~n18110;
  assign n18137 = ~n18125 & n18136;
  assign n18138 = n3444 & n18126;
  assign n18139 = ~n18135 & ~n34077;
  assign n18140 = ~n18127 & ~n18139;
  assign n18141 = ~n3116 & ~n18140;
  assign n18142 = n3116 & ~n18127;
  assign n18143 = ~n18139 & n18142;
  assign n18144 = ~n33982 & ~n17405;
  assign n18145 = ~n17405 & ~n17690;
  assign n18146 = ~n33982 & n18145;
  assign n18147 = ~n17690 & n18144;
  assign n18148 = n17025 & ~n34078;
  assign n18149 = n17404 & n18145;
  assign n18150 = n17025 & ~n33982;
  assign n18151 = ~n17405 & n18150;
  assign n18152 = ~n17690 & n18151;
  assign n18153 = ~n17025 & ~n34078;
  assign n18154 = ~n18152 & ~n18153;
  assign n18155 = ~n18148 & ~n18149;
  assign n18156 = ~n18143 & ~n34079;
  assign n18157 = ~n18141 & ~n18156;
  assign n18158 = ~n2833 & ~n18157;
  assign n18159 = n2833 & ~n18141;
  assign n18160 = ~n18156 & n18159;
  assign n18161 = n2833 & n18157;
  assign n18162 = ~n17407 & ~n17410;
  assign n18163 = ~n17410 & ~n17690;
  assign n18164 = ~n17407 & n18163;
  assign n18165 = ~n17690 & n18162;
  assign n18166 = n17017 & ~n34081;
  assign n18167 = n17408 & n18163;
  assign n18168 = n17017 & ~n17410;
  assign n18169 = ~n17407 & n18168;
  assign n18170 = ~n17690 & n18169;
  assign n18171 = ~n17017 & ~n34081;
  assign n18172 = ~n18170 & ~n18171;
  assign n18173 = ~n18166 & ~n18167;
  assign n18174 = ~n34080 & ~n34082;
  assign n18175 = ~n18158 & ~n18174;
  assign n18176 = ~n2536 & ~n18175;
  assign n18177 = n2536 & ~n18158;
  assign n18178 = ~n18174 & n18177;
  assign n18179 = n17009 & ~n33983;
  assign n18180 = ~n17416 & n18179;
  assign n18181 = ~n33983 & ~n17416;
  assign n18182 = ~n17690 & n18181;
  assign n18183 = n17009 & n18182;
  assign n18184 = ~n17690 & n18180;
  assign n18185 = ~n17009 & ~n18182;
  assign n18186 = ~n34083 & ~n18185;
  assign n18187 = ~n18178 & ~n18186;
  assign n18188 = ~n18176 & ~n18187;
  assign n18189 = ~n2283 & ~n18188;
  assign n18190 = ~n17418 & ~n17428;
  assign n18191 = ~n17690 & n18190;
  assign n18192 = ~n17426 & ~n18191;
  assign n18193 = ~n17418 & n17426;
  assign n18194 = ~n17428 & n18193;
  assign n18195 = n17426 & n18191;
  assign n18196 = ~n17690 & n18194;
  assign n18197 = ~n18192 & ~n34084;
  assign n18198 = n2283 & ~n18176;
  assign n18199 = ~n18187 & n18198;
  assign n18200 = n2283 & n18188;
  assign n18201 = ~n18197 & ~n34085;
  assign n18202 = ~n18189 & ~n18201;
  assign n18203 = ~n2021 & ~n18202;
  assign n18204 = n2021 & ~n18189;
  assign n18205 = ~n18201 & n18204;
  assign n18206 = ~n17431 & ~n33986;
  assign n18207 = ~n17431 & ~n17690;
  assign n18208 = ~n33986 & n18207;
  assign n18209 = ~n17690 & n18206;
  assign n18210 = n17439 & ~n34086;
  assign n18211 = n17443 & n18207;
  assign n18212 = n17439 & ~n33986;
  assign n18213 = ~n17431 & n18212;
  assign n18214 = ~n17690 & n18213;
  assign n18215 = ~n17439 & ~n34086;
  assign n18216 = ~n18214 & ~n18215;
  assign n18217 = ~n18210 & ~n18211;
  assign n18218 = ~n18205 & ~n34087;
  assign n18219 = ~n18203 & ~n18218;
  assign n18220 = ~n1796 & ~n18219;
  assign n18221 = ~n17445 & ~n17447;
  assign n18222 = ~n17690 & n18221;
  assign n18223 = ~n33988 & ~n18222;
  assign n18224 = ~n17445 & n33988;
  assign n18225 = ~n17447 & n18224;
  assign n18226 = n33988 & n18222;
  assign n18227 = ~n17690 & n18225;
  assign n18228 = ~n18223 & ~n34088;
  assign n18229 = n1796 & ~n18203;
  assign n18230 = ~n18218 & n18229;
  assign n18231 = n1796 & n18219;
  assign n18232 = ~n18228 & ~n34089;
  assign n18233 = ~n18220 & ~n18232;
  assign n18234 = ~n1567 & ~n18233;
  assign n18235 = n1567 & ~n18220;
  assign n18236 = ~n18232 & n18235;
  assign n18237 = ~n17462 & ~n33990;
  assign n18238 = ~n17462 & ~n17690;
  assign n18239 = ~n33990 & n18238;
  assign n18240 = ~n17690 & n18237;
  assign n18241 = n17470 & ~n34090;
  assign n18242 = n17474 & n18238;
  assign n18243 = n17470 & ~n33990;
  assign n18244 = ~n17462 & n18243;
  assign n18245 = ~n17690 & n18244;
  assign n18246 = ~n17470 & ~n34090;
  assign n18247 = ~n18245 & ~n18246;
  assign n18248 = ~n18241 & ~n18242;
  assign n18249 = ~n18236 & ~n34091;
  assign n18250 = ~n18234 & ~n18249;
  assign n18251 = ~n1374 & ~n18250;
  assign n18252 = ~n17476 & ~n17478;
  assign n18253 = ~n17690 & n18252;
  assign n18254 = ~n33992 & ~n18253;
  assign n18255 = ~n17476 & n33992;
  assign n18256 = ~n17478 & n18255;
  assign n18257 = n33992 & n18253;
  assign n18258 = ~n17690 & n18256;
  assign n18259 = ~n18254 & ~n34092;
  assign n18260 = n1374 & ~n18234;
  assign n18261 = ~n18249 & n18260;
  assign n18262 = n1374 & n18250;
  assign n18263 = ~n18259 & ~n34093;
  assign n18264 = ~n18251 & ~n18263;
  assign n18265 = ~n1179 & ~n18264;
  assign n18266 = n1179 & ~n18251;
  assign n18267 = ~n18263 & n18266;
  assign n18268 = ~n17493 & ~n33994;
  assign n18269 = ~n17493 & ~n17690;
  assign n18270 = ~n33994 & n18269;
  assign n18271 = ~n17690 & n18268;
  assign n18272 = n17501 & ~n34094;
  assign n18273 = n17505 & n18269;
  assign n18274 = n17501 & ~n33994;
  assign n18275 = ~n17493 & n18274;
  assign n18276 = ~n17690 & n18275;
  assign n18277 = ~n17501 & ~n34094;
  assign n18278 = ~n18276 & ~n18277;
  assign n18279 = ~n18272 & ~n18273;
  assign n18280 = ~n18267 & ~n34095;
  assign n18281 = ~n18265 & ~n18280;
  assign n18282 = ~n1016 & ~n18281;
  assign n18283 = n1016 & ~n18265;
  assign n18284 = ~n18280 & n18283;
  assign n18285 = n1016 & n18281;
  assign n18286 = ~n17507 & ~n17517;
  assign n18287 = ~n17507 & ~n17690;
  assign n18288 = ~n17517 & n18287;
  assign n18289 = ~n17690 & n18286;
  assign n18290 = n17515 & ~n34097;
  assign n18291 = n17518 & n18287;
  assign n18292 = ~n17507 & n17515;
  assign n18293 = ~n17517 & n18292;
  assign n18294 = ~n17690 & n18293;
  assign n18295 = ~n17515 & ~n34097;
  assign n18296 = ~n18294 & ~n18295;
  assign n18297 = ~n18290 & ~n18291;
  assign n18298 = ~n34096 & ~n34098;
  assign n18299 = ~n18282 & ~n18298;
  assign n18300 = ~n855 & ~n18299;
  assign n18301 = n855 & ~n18282;
  assign n18302 = ~n18298 & n18301;
  assign n18303 = ~n17520 & ~n33997;
  assign n18304 = ~n17520 & ~n17690;
  assign n18305 = ~n33997 & n18304;
  assign n18306 = ~n17690 & n18303;
  assign n18307 = n17528 & ~n34099;
  assign n18308 = n17532 & n18304;
  assign n18309 = n17528 & ~n33997;
  assign n18310 = ~n17520 & n18309;
  assign n18311 = ~n17690 & n18310;
  assign n18312 = ~n17528 & ~n34099;
  assign n18313 = ~n18311 & ~n18312;
  assign n18314 = ~n18307 & ~n18308;
  assign n18315 = ~n18302 & ~n34100;
  assign n18316 = ~n18300 & ~n18315;
  assign n18317 = ~n720 & ~n18316;
  assign n18318 = ~n17534 & ~n17536;
  assign n18319 = ~n17690 & n18318;
  assign n18320 = ~n33999 & ~n18319;
  assign n18321 = ~n17534 & n33999;
  assign n18322 = ~n17536 & n18321;
  assign n18323 = n33999 & n18319;
  assign n18324 = ~n17690 & n18322;
  assign n18325 = ~n18320 & ~n34101;
  assign n18326 = n720 & ~n18300;
  assign n18327 = ~n18315 & n18326;
  assign n18328 = n720 & n18316;
  assign n18329 = ~n18325 & ~n34102;
  assign n18330 = ~n18317 & ~n18329;
  assign n18331 = ~n592 & ~n18330;
  assign n18332 = n592 & ~n18317;
  assign n18333 = ~n18329 & n18332;
  assign n18334 = ~n17551 & ~n34001;
  assign n18335 = ~n17551 & ~n17690;
  assign n18336 = ~n34001 & n18335;
  assign n18337 = ~n17690 & n18334;
  assign n18338 = n17559 & ~n34103;
  assign n18339 = n17563 & n18335;
  assign n18340 = n17559 & ~n34001;
  assign n18341 = ~n17551 & n18340;
  assign n18342 = ~n17690 & n18341;
  assign n18343 = ~n17559 & ~n34103;
  assign n18344 = ~n18342 & ~n18343;
  assign n18345 = ~n18338 & ~n18339;
  assign n18346 = ~n18333 & ~n34104;
  assign n18347 = ~n18331 & ~n18346;
  assign n18348 = ~n487 & ~n18347;
  assign n18349 = n487 & ~n18331;
  assign n18350 = ~n18346 & n18349;
  assign n18351 = n487 & n18347;
  assign n18352 = ~n17565 & ~n17575;
  assign n18353 = ~n17565 & ~n17690;
  assign n18354 = ~n17575 & n18353;
  assign n18355 = ~n17690 & n18352;
  assign n18356 = n17573 & ~n34106;
  assign n18357 = n17576 & n18353;
  assign n18358 = ~n17565 & n17573;
  assign n18359 = ~n17575 & n18358;
  assign n18360 = ~n17690 & n18359;
  assign n18361 = ~n17573 & ~n34106;
  assign n18362 = ~n18360 & ~n18361;
  assign n18363 = ~n18356 & ~n18357;
  assign n18364 = ~n34105 & ~n34107;
  assign n18365 = ~n18348 & ~n18364;
  assign n18366 = ~n393 & ~n18365;
  assign n18367 = n393 & ~n18348;
  assign n18368 = ~n18364 & n18367;
  assign n18369 = ~n17578 & ~n34004;
  assign n18370 = ~n17578 & ~n17690;
  assign n18371 = ~n34004 & n18370;
  assign n18372 = ~n17690 & n18369;
  assign n18373 = n17586 & ~n34108;
  assign n18374 = n17590 & n18370;
  assign n18375 = n17586 & ~n34004;
  assign n18376 = ~n17578 & n18375;
  assign n18377 = ~n17690 & n18376;
  assign n18378 = ~n17586 & ~n34108;
  assign n18379 = ~n18377 & ~n18378;
  assign n18380 = ~n18373 & ~n18374;
  assign n18381 = ~n18368 & ~n34109;
  assign n18382 = ~n18366 & ~n18381;
  assign n18383 = ~n321 & ~n18382;
  assign n18384 = ~n17592 & ~n17594;
  assign n18385 = ~n17690 & n18384;
  assign n18386 = ~n34006 & ~n18385;
  assign n18387 = ~n17592 & n34006;
  assign n18388 = ~n17594 & n18387;
  assign n18389 = n34006 & n18385;
  assign n18390 = ~n17690 & n18388;
  assign n18391 = ~n18386 & ~n34110;
  assign n18392 = n321 & ~n18366;
  assign n18393 = ~n18381 & n18392;
  assign n18394 = n321 & n18382;
  assign n18395 = ~n18391 & ~n34111;
  assign n18396 = ~n18383 & ~n18395;
  assign n18397 = ~n263 & ~n18396;
  assign n18398 = n263 & ~n18383;
  assign n18399 = ~n18395 & n18398;
  assign n18400 = ~n17609 & ~n34008;
  assign n18401 = ~n17609 & ~n17690;
  assign n18402 = ~n34008 & n18401;
  assign n18403 = ~n17690 & n18400;
  assign n18404 = n17617 & ~n34112;
  assign n18405 = n17621 & n18401;
  assign n18406 = n17617 & ~n34008;
  assign n18407 = ~n17609 & n18406;
  assign n18408 = ~n17690 & n18407;
  assign n18409 = ~n17617 & ~n34112;
  assign n18410 = ~n18408 & ~n18409;
  assign n18411 = ~n18404 & ~n18405;
  assign n18412 = ~n18399 & ~n34113;
  assign n18413 = ~n18397 & ~n18412;
  assign n18414 = ~n214 & ~n18413;
  assign n18415 = n214 & ~n18397;
  assign n18416 = ~n18412 & n18415;
  assign n18417 = n214 & n18413;
  assign n18418 = ~n17623 & ~n17633;
  assign n18419 = ~n17623 & ~n17690;
  assign n18420 = ~n17633 & n18419;
  assign n18421 = ~n17690 & n18418;
  assign n18422 = n17631 & ~n34115;
  assign n18423 = n17634 & n18419;
  assign n18424 = ~n17623 & n17631;
  assign n18425 = ~n17633 & n18424;
  assign n18426 = ~n17690 & n18425;
  assign n18427 = ~n17631 & ~n34115;
  assign n18428 = ~n18426 & ~n18427;
  assign n18429 = ~n18422 & ~n18423;
  assign n18430 = ~n34114 & ~n34116;
  assign n18431 = ~n18414 & ~n18430;
  assign n18432 = ~n197 & ~n18431;
  assign n18433 = n197 & ~n18414;
  assign n18434 = ~n18430 & n18433;
  assign n18435 = ~n17636 & ~n34011;
  assign n18436 = ~n17636 & ~n17690;
  assign n18437 = ~n34011 & n18436;
  assign n18438 = ~n17690 & n18435;
  assign n18439 = n17644 & ~n34117;
  assign n18440 = n17648 & n18436;
  assign n18441 = n17644 & ~n34011;
  assign n18442 = ~n17636 & n18441;
  assign n18443 = ~n17690 & n18442;
  assign n18444 = ~n17644 & ~n34117;
  assign n18445 = ~n18443 & ~n18444;
  assign n18446 = ~n18439 & ~n18440;
  assign n18447 = ~n18434 & ~n34118;
  assign n18448 = ~n18432 & ~n18447;
  assign n18449 = ~n17650 & ~n17652;
  assign n18450 = ~n17690 & n18449;
  assign n18451 = ~n34013 & ~n18450;
  assign n18452 = ~n17650 & n34013;
  assign n18453 = ~n17652 & n18452;
  assign n18454 = n34013 & n18450;
  assign n18455 = ~n17690 & n18453;
  assign n18456 = ~n18451 & ~n34119;
  assign n18457 = ~n17666 & ~n17674;
  assign n18458 = ~n17674 & ~n17690;
  assign n18459 = ~n17666 & n18458;
  assign n18460 = ~n17690 & n18457;
  assign n18461 = ~n34016 & ~n34120;
  assign n18462 = ~n18456 & n18461;
  assign n18463 = ~n18448 & n18462;
  assign n18464 = n193 & ~n18463;
  assign n18465 = ~n18432 & n18456;
  assign n18466 = ~n18447 & n18465;
  assign n18467 = n18448 & n18456;
  assign n18468 = n17666 & ~n18458;
  assign n18469 = ~n193 & ~n18457;
  assign n18470 = ~n18468 & n18469;
  assign n18471 = ~n34121 & ~n18470;
  assign n18472 = ~n18464 & n18471;
  assign n18473 = ~n18176 & ~n18178;
  assign n18474 = ~n18472 & n18473;
  assign n18475 = ~n18186 & ~n18474;
  assign n18476 = ~n18178 & n18186;
  assign n18477 = ~n18176 & n18476;
  assign n18478 = n18186 & n18474;
  assign n18479 = ~n18472 & n18477;
  assign n18480 = ~n18475 & ~n34122;
  assign n18481 = ~n18158 & ~n34080;
  assign n18482 = ~n18472 & n18481;
  assign n18483 = ~n34082 & ~n18482;
  assign n18484 = ~n18158 & n34082;
  assign n18485 = ~n34080 & n18484;
  assign n18486 = n34082 & n18482;
  assign n18487 = ~n18472 & n18485;
  assign n18488 = ~n18483 & ~n34123;
  assign n18489 = ~n18141 & ~n18143;
  assign n18490 = ~n18472 & n18489;
  assign n18491 = ~n34079 & ~n18490;
  assign n18492 = ~n18143 & n34079;
  assign n18493 = ~n18141 & n18492;
  assign n18494 = n34079 & n18490;
  assign n18495 = ~n18472 & n18493;
  assign n18496 = ~n18491 & ~n34124;
  assign n18497 = ~n18110 & ~n18112;
  assign n18498 = ~n18472 & n18497;
  assign n18499 = ~n34075 & ~n18498;
  assign n18500 = ~n18112 & n34075;
  assign n18501 = ~n18110 & n18500;
  assign n18502 = n34075 & n18498;
  assign n18503 = ~n18472 & n18501;
  assign n18504 = ~n18499 & ~n34125;
  assign n18505 = ~n18092 & ~n34071;
  assign n18506 = ~n18472 & n18505;
  assign n18507 = ~n34073 & ~n18506;
  assign n18508 = ~n18092 & n34073;
  assign n18509 = ~n34071 & n18508;
  assign n18510 = n34073 & n18506;
  assign n18511 = ~n18472 & n18509;
  assign n18512 = ~n18507 & ~n34126;
  assign n18513 = ~n18075 & ~n18077;
  assign n18514 = ~n18472 & n18513;
  assign n18515 = ~n34070 & ~n18514;
  assign n18516 = ~n18077 & n34070;
  assign n18517 = ~n18075 & n18516;
  assign n18518 = n34070 & n18514;
  assign n18519 = ~n18472 & n18517;
  assign n18520 = ~n18515 & ~n34127;
  assign n18521 = ~n18044 & ~n18046;
  assign n18522 = ~n18472 & n18521;
  assign n18523 = ~n34066 & ~n18522;
  assign n18524 = ~n18046 & n34066;
  assign n18525 = ~n18044 & n18524;
  assign n18526 = n34066 & n18522;
  assign n18527 = ~n18472 & n18525;
  assign n18528 = ~n18523 & ~n34128;
  assign n18529 = ~n18026 & ~n34062;
  assign n18530 = ~n18472 & n18529;
  assign n18531 = ~n34064 & ~n18530;
  assign n18532 = ~n18026 & n34064;
  assign n18533 = ~n34062 & n18532;
  assign n18534 = n34064 & n18530;
  assign n18535 = ~n18472 & n18533;
  assign n18536 = ~n18531 & ~n34129;
  assign n18537 = ~n18009 & ~n18011;
  assign n18538 = ~n18472 & n18537;
  assign n18539 = ~n34061 & ~n18538;
  assign n18540 = ~n18011 & n34061;
  assign n18541 = ~n18009 & n18540;
  assign n18542 = n34061 & n18538;
  assign n18543 = ~n18472 & n18541;
  assign n18544 = ~n18539 & ~n34130;
  assign n18545 = ~n17978 & ~n17980;
  assign n18546 = ~n18472 & n18545;
  assign n18547 = ~n34057 & ~n18546;
  assign n18548 = ~n17980 & n34057;
  assign n18549 = ~n17978 & n18548;
  assign n18550 = n34057 & n18546;
  assign n18551 = ~n18472 & n18549;
  assign n18552 = ~n18547 & ~n34131;
  assign n18553 = ~n17960 & ~n34053;
  assign n18554 = ~n18472 & n18553;
  assign n18555 = ~n34055 & ~n18554;
  assign n18556 = ~n17960 & n34055;
  assign n18557 = ~n34053 & n18556;
  assign n18558 = n34055 & n18554;
  assign n18559 = ~n18472 & n18557;
  assign n18560 = ~n18555 & ~n34132;
  assign n18561 = ~n17943 & ~n17945;
  assign n18562 = ~n18472 & n18561;
  assign n18563 = ~n34052 & ~n18562;
  assign n18564 = ~n17945 & n34052;
  assign n18565 = ~n17943 & n18564;
  assign n18566 = n34052 & n18562;
  assign n18567 = ~n18472 & n18565;
  assign n18568 = ~n18563 & ~n34133;
  assign n18569 = ~n17912 & ~n17914;
  assign n18570 = ~n18472 & n18569;
  assign n18571 = ~n34048 & ~n18570;
  assign n18572 = ~n17914 & n34048;
  assign n18573 = ~n17912 & n18572;
  assign n18574 = n34048 & n18570;
  assign n18575 = ~n18472 & n18573;
  assign n18576 = ~n18571 & ~n34134;
  assign n18577 = ~n17893 & ~n34043;
  assign n18578 = ~n18472 & n18577;
  assign n18579 = ~n34046 & ~n18578;
  assign n18580 = ~n17893 & n34046;
  assign n18581 = ~n34043 & n18580;
  assign n18582 = n34046 & n18578;
  assign n18583 = ~n18472 & n18581;
  assign n18584 = ~n18579 & ~n34135;
  assign n18585 = ~n17876 & ~n17878;
  assign n18586 = ~n18472 & n18585;
  assign n18587 = ~n34042 & ~n18586;
  assign n18588 = ~n17878 & n34042;
  assign n18589 = ~n17876 & n18588;
  assign n18590 = n34042 & n18586;
  assign n18591 = ~n18472 & n18589;
  assign n18592 = ~n18587 & ~n34136;
  assign n18593 = ~n17842 & ~n17844;
  assign n18594 = ~n18472 & n18593;
  assign n18595 = ~n34037 & ~n18594;
  assign n18596 = ~n17844 & n34037;
  assign n18597 = ~n17842 & n18596;
  assign n18598 = n34037 & n18594;
  assign n18599 = ~n18472 & n18597;
  assign n18600 = ~n18595 & ~n34137;
  assign n18601 = ~n17809 & ~n17811;
  assign n18602 = ~n18472 & n18601;
  assign n18603 = ~n34033 & ~n18602;
  assign n18604 = ~n17811 & n34033;
  assign n18605 = ~n17809 & n18604;
  assign n18606 = n34033 & n18602;
  assign n18607 = ~n18472 & n18605;
  assign n18608 = ~n18603 & ~n34138;
  assign n18609 = ~n17776 & ~n17778;
  assign n18610 = ~n18472 & n18609;
  assign n18611 = ~n34029 & ~n18610;
  assign n18612 = ~n17778 & n34029;
  assign n18613 = ~n17776 & n18612;
  assign n18614 = n34029 & n18610;
  assign n18615 = ~n18472 & n18613;
  assign n18616 = ~n18611 & ~n34139;
  assign n18617 = ~n17742 & ~n17744;
  assign n18618 = ~n18472 & n18617;
  assign n18619 = ~n34024 & ~n18618;
  assign n18620 = ~n17744 & n34024;
  assign n18621 = ~n17742 & n18620;
  assign n18622 = n34024 & n18618;
  assign n18623 = ~n18472 & n18621;
  assign n18624 = ~n18619 & ~n34140;
  assign n18625 = ~n17715 & ~n17717;
  assign n18626 = ~n18472 & n18625;
  assign n18627 = ~n17726 & ~n18626;
  assign n18628 = ~n17717 & n17726;
  assign n18629 = ~n17715 & n18628;
  assign n18630 = n17726 & n18626;
  assign n18631 = ~n18472 & n18629;
  assign n18632 = ~n18627 & ~n34141;
  assign n18633 = ~pi30  & ~n18472;
  assign n18634 = ~pi31  & n18633;
  assign n18635 = n17692 & ~n18472;
  assign n18636 = ~n17690 & ~n18470;
  assign n18637 = ~n34121 & n18636;
  assign n18638 = ~n18464 & n18637;
  assign n18639 = ~n34142 & ~n18638;
  assign n18640 = pi32  & ~n18639;
  assign n18641 = ~pi32  & ~n18638;
  assign n18642 = ~pi32  & n18639;
  assign n18643 = ~n34142 & n18641;
  assign n18644 = ~n18640 & ~n34143;
  assign n18645 = pi30  & ~n18472;
  assign n18646 = ~pi28  & ~pi29 ;
  assign n18647 = ~pi30  & n18646;
  assign n18648 = ~n16982 & ~n34018;
  assign n18649 = ~n16983 & n18648;
  assign n18650 = ~n16999 & n18649;
  assign n18651 = ~n33932 & n18650;
  assign n18652 = n33930 & n17001;
  assign n18653 = ~n16993 & n18651;
  assign n18654 = ~n18647 & ~n34144;
  assign n18655 = ~n17688 & n18654;
  assign n18656 = ~n34016 & n18655;
  assign n18657 = ~n17682 & n18656;
  assign n18658 = ~n18645 & ~n18647;
  assign n18659 = n17690 & n18658;
  assign n18660 = ~n18645 & n18657;
  assign n18661 = pi31  & ~n18633;
  assign n18662 = ~n34142 & ~n18661;
  assign n18663 = ~n34145 & n18662;
  assign n18664 = ~n17690 & ~n18658;
  assign n18665 = n17001 & ~n18664;
  assign n18666 = ~n18663 & ~n18664;
  assign n18667 = n17001 & n18666;
  assign n18668 = ~n18663 & n18665;
  assign n18669 = ~n18644 & ~n34146;
  assign n18670 = ~n17001 & ~n18666;
  assign n18671 = n16248 & ~n18670;
  assign n18672 = ~n18669 & n18671;
  assign n18673 = ~n17695 & ~n34019;
  assign n18674 = ~n18472 & n18673;
  assign n18675 = n17700 & ~n18674;
  assign n18676 = ~n17700 & n18673;
  assign n18677 = ~n17700 & n18674;
  assign n18678 = ~n18472 & n18676;
  assign n18679 = ~n18675 & ~n34147;
  assign n18680 = ~n18672 & ~n18679;
  assign n18681 = ~n18669 & ~n18670;
  assign n18682 = ~n16248 & ~n18681;
  assign n18683 = n15586 & ~n18682;
  assign n18684 = ~n18680 & ~n18682;
  assign n18685 = n15586 & n18684;
  assign n18686 = ~n18680 & n18683;
  assign n18687 = ~n18632 & ~n34148;
  assign n18688 = ~n15586 & ~n18684;
  assign n18689 = n14866 & ~n18688;
  assign n18690 = ~n18687 & n18689;
  assign n18691 = ~n17729 & ~n34021;
  assign n18692 = ~n18472 & n18691;
  assign n18693 = ~n17739 & ~n18692;
  assign n18694 = ~n17729 & n17739;
  assign n18695 = ~n34021 & n18694;
  assign n18696 = n17739 & n18692;
  assign n18697 = ~n18472 & n18695;
  assign n18698 = n17739 & ~n18692;
  assign n18699 = ~n17739 & n18692;
  assign n18700 = ~n18698 & ~n18699;
  assign n18701 = ~n18693 & ~n34149;
  assign n18702 = ~n18690 & n34150;
  assign n18703 = ~n18687 & ~n18688;
  assign n18704 = ~n14866 & ~n18703;
  assign n18705 = n14233 & ~n18704;
  assign n18706 = ~n18702 & ~n18704;
  assign n18707 = n14233 & n18706;
  assign n18708 = ~n18702 & n18705;
  assign n18709 = ~n18624 & ~n34151;
  assign n18710 = ~n14233 & ~n18706;
  assign n18711 = n13548 & ~n18710;
  assign n18712 = ~n18709 & n18711;
  assign n18713 = ~n17759 & ~n34025;
  assign n18714 = ~n18472 & n18713;
  assign n18715 = ~n34027 & ~n18714;
  assign n18716 = n34027 & n18714;
  assign n18717 = ~n17759 & ~n34027;
  assign n18718 = ~n34025 & n18717;
  assign n18719 = ~n18472 & n18718;
  assign n18720 = n34027 & ~n18714;
  assign n18721 = ~n18719 & ~n18720;
  assign n18722 = ~n18715 & ~n18716;
  assign n18723 = ~n18712 & ~n34152;
  assign n18724 = ~n18709 & ~n18710;
  assign n18725 = ~n13548 & ~n18724;
  assign n18726 = n12948 & ~n18725;
  assign n18727 = ~n18723 & ~n18725;
  assign n18728 = n12948 & n18727;
  assign n18729 = ~n18723 & n18726;
  assign n18730 = ~n18616 & ~n34153;
  assign n18731 = ~n12948 & ~n18727;
  assign n18732 = n12296 & ~n18731;
  assign n18733 = ~n18730 & n18732;
  assign n18734 = ~n17793 & ~n34030;
  assign n18735 = ~n18472 & n18734;
  assign n18736 = ~n34031 & n18735;
  assign n18737 = n34031 & ~n18735;
  assign n18738 = ~n17793 & n34031;
  assign n18739 = ~n34030 & n18738;
  assign n18740 = ~n18472 & n18739;
  assign n18741 = ~n34031 & ~n18735;
  assign n18742 = ~n18740 & ~n18741;
  assign n18743 = ~n18736 & ~n18737;
  assign n18744 = ~n18733 & ~n34154;
  assign n18745 = ~n18730 & ~n18731;
  assign n18746 = ~n12296 & ~n18745;
  assign n18747 = n11719 & ~n18746;
  assign n18748 = ~n18744 & ~n18746;
  assign n18749 = n11719 & n18748;
  assign n18750 = ~n18744 & n18747;
  assign n18751 = ~n18608 & ~n34155;
  assign n18752 = ~n11719 & ~n18748;
  assign n18753 = n11097 & ~n18752;
  assign n18754 = ~n18751 & n18753;
  assign n18755 = ~n17826 & ~n34034;
  assign n18756 = ~n18472 & n18755;
  assign n18757 = ~n34035 & n18756;
  assign n18758 = n34035 & ~n18756;
  assign n18759 = ~n34035 & ~n18756;
  assign n18760 = ~n17826 & n34035;
  assign n18761 = ~n34034 & n18760;
  assign n18762 = n34035 & n18756;
  assign n18763 = ~n18472 & n18761;
  assign n18764 = ~n18759 & ~n34156;
  assign n18765 = ~n18757 & ~n18758;
  assign n18766 = ~n18754 & ~n34157;
  assign n18767 = ~n18751 & ~n18752;
  assign n18768 = ~n11097 & ~n18767;
  assign n18769 = n10555 & ~n18768;
  assign n18770 = ~n18766 & ~n18768;
  assign n18771 = n10555 & n18770;
  assign n18772 = ~n18766 & n18769;
  assign n18773 = ~n18600 & ~n34158;
  assign n18774 = ~n10555 & ~n18770;
  assign n18775 = n9969 & ~n18774;
  assign n18776 = ~n18773 & n18775;
  assign n18777 = ~n17859 & ~n34038;
  assign n18778 = ~n17859 & ~n18472;
  assign n18779 = ~n34038 & n18778;
  assign n18780 = ~n18472 & n18777;
  assign n18781 = n34040 & ~n34159;
  assign n18782 = n17874 & n18778;
  assign n18783 = ~n34040 & n34159;
  assign n18784 = ~n17859 & n34040;
  assign n18785 = ~n34038 & n18784;
  assign n18786 = ~n18472 & n18785;
  assign n18787 = ~n34040 & ~n34159;
  assign n18788 = ~n18786 & ~n18787;
  assign n18789 = ~n18781 & ~n34160;
  assign n18790 = ~n18776 & ~n34161;
  assign n18791 = ~n18773 & ~n18774;
  assign n18792 = ~n9969 & ~n18791;
  assign n18793 = n9457 & ~n18792;
  assign n18794 = ~n18790 & ~n18792;
  assign n18795 = n9457 & n18794;
  assign n18796 = ~n18790 & n18793;
  assign n18797 = ~n18592 & ~n34162;
  assign n18798 = ~n9457 & ~n18794;
  assign n18799 = n8896 & ~n18798;
  assign n18800 = ~n18797 & n18799;
  assign n18801 = ~n18584 & ~n18800;
  assign n18802 = ~n18797 & ~n18798;
  assign n18803 = ~n8896 & ~n18802;
  assign n18804 = n8411 & ~n18803;
  assign n18805 = ~n18801 & ~n18803;
  assign n18806 = n8411 & n18805;
  assign n18807 = ~n18801 & n18804;
  assign n18808 = ~n18576 & ~n34163;
  assign n18809 = ~n8411 & ~n18805;
  assign n18810 = n7885 & ~n18809;
  assign n18811 = ~n18808 & n18810;
  assign n18812 = ~n17929 & ~n34050;
  assign n18813 = ~n17929 & ~n18472;
  assign n18814 = ~n34050 & n18813;
  assign n18815 = ~n18472 & n18812;
  assign n18816 = n17937 & ~n34164;
  assign n18817 = n17941 & n18813;
  assign n18818 = ~n17929 & n17937;
  assign n18819 = ~n34050 & n18818;
  assign n18820 = ~n18472 & n18819;
  assign n18821 = ~n17937 & ~n34164;
  assign n18822 = ~n18820 & ~n18821;
  assign n18823 = ~n18816 & ~n18817;
  assign n18824 = ~n18811 & ~n34165;
  assign n18825 = ~n18808 & ~n18809;
  assign n18826 = ~n7885 & ~n18825;
  assign n18827 = n7428 & ~n18826;
  assign n18828 = ~n18824 & ~n18826;
  assign n18829 = n7428 & n18828;
  assign n18830 = ~n18824 & n18827;
  assign n18831 = ~n18568 & ~n34166;
  assign n18832 = ~n7428 & ~n18828;
  assign n18833 = n6937 & ~n18832;
  assign n18834 = ~n18831 & n18833;
  assign n18835 = ~n18560 & ~n18834;
  assign n18836 = ~n18831 & ~n18832;
  assign n18837 = ~n6937 & ~n18836;
  assign n18838 = n6507 & ~n18837;
  assign n18839 = ~n18835 & ~n18837;
  assign n18840 = n6507 & n18839;
  assign n18841 = ~n18835 & n18838;
  assign n18842 = ~n18552 & ~n34167;
  assign n18843 = ~n6507 & ~n18839;
  assign n18844 = n6051 & ~n18843;
  assign n18845 = ~n18842 & n18844;
  assign n18846 = ~n17995 & ~n34059;
  assign n18847 = ~n17995 & ~n18472;
  assign n18848 = ~n34059 & n18847;
  assign n18849 = ~n18472 & n18846;
  assign n18850 = n18003 & ~n34168;
  assign n18851 = n18007 & n18847;
  assign n18852 = ~n17995 & n18003;
  assign n18853 = ~n34059 & n18852;
  assign n18854 = ~n18472 & n18853;
  assign n18855 = ~n18003 & ~n34168;
  assign n18856 = ~n18854 & ~n18855;
  assign n18857 = ~n18850 & ~n18851;
  assign n18858 = ~n18845 & ~n34169;
  assign n18859 = ~n18842 & ~n18843;
  assign n18860 = ~n6051 & ~n18859;
  assign n18861 = n5648 & ~n18860;
  assign n18862 = ~n18858 & ~n18860;
  assign n18863 = n5648 & n18862;
  assign n18864 = ~n18858 & n18861;
  assign n18865 = ~n18544 & ~n34170;
  assign n18866 = ~n5648 & ~n18862;
  assign n18867 = n5223 & ~n18866;
  assign n18868 = ~n18865 & n18867;
  assign n18869 = ~n18536 & ~n18868;
  assign n18870 = ~n18865 & ~n18866;
  assign n18871 = ~n5223 & ~n18870;
  assign n18872 = n4851 & ~n18871;
  assign n18873 = ~n18869 & ~n18871;
  assign n18874 = n4851 & n18873;
  assign n18875 = ~n18869 & n18872;
  assign n18876 = ~n18528 & ~n34171;
  assign n18877 = ~n4851 & ~n18873;
  assign n18878 = n4461 & ~n18877;
  assign n18879 = ~n18876 & n18878;
  assign n18880 = ~n18061 & ~n34068;
  assign n18881 = ~n18061 & ~n18472;
  assign n18882 = ~n34068 & n18881;
  assign n18883 = ~n18472 & n18880;
  assign n18884 = n18069 & ~n34172;
  assign n18885 = n18073 & n18881;
  assign n18886 = ~n18061 & n18069;
  assign n18887 = ~n34068 & n18886;
  assign n18888 = ~n18472 & n18887;
  assign n18889 = ~n18069 & ~n34172;
  assign n18890 = ~n18888 & ~n18889;
  assign n18891 = ~n18884 & ~n18885;
  assign n18892 = ~n18879 & ~n34173;
  assign n18893 = ~n18876 & ~n18877;
  assign n18894 = ~n4461 & ~n18893;
  assign n18895 = n4115 & ~n18894;
  assign n18896 = ~n18892 & ~n18894;
  assign n18897 = n4115 & n18896;
  assign n18898 = ~n18892 & n18895;
  assign n18899 = ~n18520 & ~n34174;
  assign n18900 = ~n4115 & ~n18896;
  assign n18901 = n3754 & ~n18900;
  assign n18902 = ~n18899 & n18901;
  assign n18903 = ~n18512 & ~n18902;
  assign n18904 = ~n18899 & ~n18900;
  assign n18905 = ~n3754 & ~n18904;
  assign n18906 = n3444 & ~n18905;
  assign n18907 = ~n18903 & ~n18905;
  assign n18908 = n3444 & n18907;
  assign n18909 = ~n18903 & n18906;
  assign n18910 = ~n18504 & ~n34175;
  assign n18911 = ~n3444 & ~n18907;
  assign n18912 = n3116 & ~n18911;
  assign n18913 = ~n18910 & n18912;
  assign n18914 = ~n18127 & ~n34077;
  assign n18915 = ~n18127 & ~n18472;
  assign n18916 = ~n34077 & n18915;
  assign n18917 = ~n18472 & n18914;
  assign n18918 = n18135 & ~n34176;
  assign n18919 = n18139 & n18915;
  assign n18920 = ~n18127 & n18135;
  assign n18921 = ~n34077 & n18920;
  assign n18922 = ~n18472 & n18921;
  assign n18923 = ~n18135 & ~n34176;
  assign n18924 = ~n18922 & ~n18923;
  assign n18925 = ~n18918 & ~n18919;
  assign n18926 = ~n18913 & ~n34177;
  assign n18927 = ~n18910 & ~n18911;
  assign n18928 = ~n3116 & ~n18927;
  assign n18929 = n2833 & ~n18928;
  assign n18930 = ~n18926 & ~n18928;
  assign n18931 = n2833 & n18930;
  assign n18932 = ~n18926 & n18929;
  assign n18933 = ~n18496 & ~n34178;
  assign n18934 = ~n2833 & ~n18930;
  assign n18935 = n2536 & ~n18934;
  assign n18936 = ~n18933 & n18935;
  assign n18937 = ~n18488 & ~n18936;
  assign n18938 = ~n18933 & ~n18934;
  assign n18939 = ~n2536 & ~n18938;
  assign n18940 = n2283 & ~n18939;
  assign n18941 = ~n18937 & ~n18939;
  assign n18942 = n2283 & n18941;
  assign n18943 = ~n18937 & n18940;
  assign n18944 = ~n18480 & ~n34179;
  assign n18945 = ~n2283 & ~n18941;
  assign n18946 = ~n18944 & ~n18945;
  assign n18947 = ~n2021 & ~n18946;
  assign n18948 = ~n18189 & ~n34085;
  assign n18949 = ~n18472 & n18948;
  assign n18950 = n18197 & ~n18949;
  assign n18951 = ~n18197 & n18949;
  assign n18952 = ~n18189 & n18197;
  assign n18953 = ~n34085 & n18952;
  assign n18954 = ~n18472 & n18953;
  assign n18955 = ~n18197 & ~n18949;
  assign n18956 = ~n18954 & ~n18955;
  assign n18957 = ~n18950 & ~n18951;
  assign n18958 = n2021 & ~n18945;
  assign n18959 = ~n18944 & n18958;
  assign n18960 = ~n34180 & ~n18959;
  assign n18961 = ~n18947 & ~n18960;
  assign n18962 = ~n1796 & ~n18961;
  assign n18963 = ~n18203 & ~n18205;
  assign n18964 = ~n18472 & n18963;
  assign n18965 = ~n34087 & ~n18964;
  assign n18966 = ~n18205 & n34087;
  assign n18967 = ~n18203 & n18966;
  assign n18968 = n34087 & n18964;
  assign n18969 = ~n18472 & n18967;
  assign n18970 = ~n18965 & ~n34181;
  assign n18971 = n1796 & ~n18947;
  assign n18972 = n1796 & n18961;
  assign n18973 = ~n18960 & n18971;
  assign n18974 = ~n18970 & ~n34182;
  assign n18975 = ~n18962 & ~n18974;
  assign n18976 = ~n1567 & ~n18975;
  assign n18977 = n1567 & ~n18962;
  assign n18978 = ~n18974 & n18977;
  assign n18979 = ~n18220 & ~n34089;
  assign n18980 = ~n18220 & ~n18472;
  assign n18981 = ~n34089 & n18980;
  assign n18982 = ~n18472 & n18979;
  assign n18983 = n18228 & ~n34183;
  assign n18984 = n18232 & n18980;
  assign n18985 = ~n18220 & n18228;
  assign n18986 = ~n34089 & n18985;
  assign n18987 = ~n18472 & n18986;
  assign n18988 = ~n18228 & ~n34183;
  assign n18989 = ~n18987 & ~n18988;
  assign n18990 = ~n18983 & ~n18984;
  assign n18991 = ~n18978 & ~n34184;
  assign n18992 = ~n18976 & ~n18991;
  assign n18993 = ~n1374 & ~n18992;
  assign n18994 = ~n18234 & ~n18236;
  assign n18995 = ~n18472 & n18994;
  assign n18996 = ~n34091 & ~n18995;
  assign n18997 = ~n18236 & n34091;
  assign n18998 = ~n18234 & n18997;
  assign n18999 = n34091 & n18995;
  assign n19000 = ~n18472 & n18998;
  assign n19001 = ~n18996 & ~n34185;
  assign n19002 = n1374 & ~n18976;
  assign n19003 = n1374 & n18992;
  assign n19004 = ~n18991 & n19002;
  assign n19005 = ~n19001 & ~n34186;
  assign n19006 = ~n18993 & ~n19005;
  assign n19007 = ~n1179 & ~n19006;
  assign n19008 = n1179 & ~n18993;
  assign n19009 = ~n19005 & n19008;
  assign n19010 = ~n18251 & ~n34093;
  assign n19011 = ~n18251 & ~n18472;
  assign n19012 = ~n34093 & n19011;
  assign n19013 = ~n18472 & n19010;
  assign n19014 = n18259 & ~n34187;
  assign n19015 = n18263 & n19011;
  assign n19016 = ~n18251 & n18259;
  assign n19017 = ~n34093 & n19016;
  assign n19018 = ~n18472 & n19017;
  assign n19019 = ~n18259 & ~n34187;
  assign n19020 = ~n19018 & ~n19019;
  assign n19021 = ~n19014 & ~n19015;
  assign n19022 = ~n19009 & ~n34188;
  assign n19023 = ~n19007 & ~n19022;
  assign n19024 = ~n1016 & ~n19023;
  assign n19025 = ~n18265 & ~n18267;
  assign n19026 = ~n18472 & n19025;
  assign n19027 = ~n34095 & ~n19026;
  assign n19028 = ~n18267 & n34095;
  assign n19029 = ~n18265 & n19028;
  assign n19030 = n34095 & n19026;
  assign n19031 = ~n18472 & n19029;
  assign n19032 = ~n19027 & ~n34189;
  assign n19033 = n1016 & ~n19007;
  assign n19034 = n1016 & n19023;
  assign n19035 = ~n19022 & n19033;
  assign n19036 = ~n19032 & ~n34190;
  assign n19037 = ~n19024 & ~n19036;
  assign n19038 = ~n855 & ~n19037;
  assign n19039 = ~n18282 & ~n34096;
  assign n19040 = ~n18472 & n19039;
  assign n19041 = ~n34098 & ~n19040;
  assign n19042 = ~n18282 & n34098;
  assign n19043 = ~n34096 & n19042;
  assign n19044 = n34098 & n19040;
  assign n19045 = ~n18472 & n19043;
  assign n19046 = ~n19041 & ~n34191;
  assign n19047 = n855 & ~n19024;
  assign n19048 = ~n19036 & n19047;
  assign n19049 = ~n19046 & ~n19048;
  assign n19050 = ~n19038 & ~n19049;
  assign n19051 = ~n720 & ~n19050;
  assign n19052 = ~n18300 & ~n18302;
  assign n19053 = ~n18472 & n19052;
  assign n19054 = ~n34100 & ~n19053;
  assign n19055 = ~n18302 & n34100;
  assign n19056 = ~n18300 & n19055;
  assign n19057 = n34100 & n19053;
  assign n19058 = ~n18472 & n19056;
  assign n19059 = ~n19054 & ~n34192;
  assign n19060 = n720 & ~n19038;
  assign n19061 = n720 & n19050;
  assign n19062 = ~n19049 & n19060;
  assign n19063 = ~n19059 & ~n34193;
  assign n19064 = ~n19051 & ~n19063;
  assign n19065 = ~n592 & ~n19064;
  assign n19066 = n592 & ~n19051;
  assign n19067 = ~n19063 & n19066;
  assign n19068 = ~n18317 & ~n34102;
  assign n19069 = ~n18317 & ~n18472;
  assign n19070 = ~n34102 & n19069;
  assign n19071 = ~n18472 & n19068;
  assign n19072 = n18325 & ~n34194;
  assign n19073 = n18329 & n19069;
  assign n19074 = ~n18317 & n18325;
  assign n19075 = ~n34102 & n19074;
  assign n19076 = ~n18472 & n19075;
  assign n19077 = ~n18325 & ~n34194;
  assign n19078 = ~n19076 & ~n19077;
  assign n19079 = ~n19072 & ~n19073;
  assign n19080 = ~n19067 & ~n34195;
  assign n19081 = ~n19065 & ~n19080;
  assign n19082 = ~n487 & ~n19081;
  assign n19083 = ~n18331 & ~n18333;
  assign n19084 = ~n18472 & n19083;
  assign n19085 = ~n34104 & ~n19084;
  assign n19086 = ~n18333 & n34104;
  assign n19087 = ~n18331 & n19086;
  assign n19088 = n34104 & n19084;
  assign n19089 = ~n18472 & n19087;
  assign n19090 = ~n19085 & ~n34196;
  assign n19091 = n487 & ~n19065;
  assign n19092 = n487 & n19081;
  assign n19093 = ~n19080 & n19091;
  assign n19094 = ~n19090 & ~n34197;
  assign n19095 = ~n19082 & ~n19094;
  assign n19096 = ~n393 & ~n19095;
  assign n19097 = ~n18348 & ~n34105;
  assign n19098 = ~n18472 & n19097;
  assign n19099 = ~n34107 & ~n19098;
  assign n19100 = ~n18348 & n34107;
  assign n19101 = ~n34105 & n19100;
  assign n19102 = n34107 & n19098;
  assign n19103 = ~n18472 & n19101;
  assign n19104 = ~n19099 & ~n34198;
  assign n19105 = n393 & ~n19082;
  assign n19106 = ~n19094 & n19105;
  assign n19107 = ~n19104 & ~n19106;
  assign n19108 = ~n19096 & ~n19107;
  assign n19109 = ~n321 & ~n19108;
  assign n19110 = ~n18366 & ~n18368;
  assign n19111 = ~n18472 & n19110;
  assign n19112 = ~n34109 & ~n19111;
  assign n19113 = ~n18368 & n34109;
  assign n19114 = ~n18366 & n19113;
  assign n19115 = n34109 & n19111;
  assign n19116 = ~n18472 & n19114;
  assign n19117 = ~n19112 & ~n34199;
  assign n19118 = n321 & ~n19096;
  assign n19119 = n321 & n19108;
  assign n19120 = ~n19107 & n19118;
  assign n19121 = ~n19117 & ~n34200;
  assign n19122 = ~n19109 & ~n19121;
  assign n19123 = ~n263 & ~n19122;
  assign n19124 = n263 & ~n19109;
  assign n19125 = ~n19121 & n19124;
  assign n19126 = ~n18383 & ~n34111;
  assign n19127 = ~n18383 & ~n18472;
  assign n19128 = ~n34111 & n19127;
  assign n19129 = ~n18472 & n19126;
  assign n19130 = n18391 & ~n34201;
  assign n19131 = n18395 & n19127;
  assign n19132 = ~n18383 & n18391;
  assign n19133 = ~n34111 & n19132;
  assign n19134 = ~n18472 & n19133;
  assign n19135 = ~n18391 & ~n34201;
  assign n19136 = ~n19134 & ~n19135;
  assign n19137 = ~n19130 & ~n19131;
  assign n19138 = ~n19125 & ~n34202;
  assign n19139 = ~n19123 & ~n19138;
  assign n19140 = ~n214 & ~n19139;
  assign n19141 = ~n18397 & ~n18399;
  assign n19142 = ~n18472 & n19141;
  assign n19143 = ~n34113 & ~n19142;
  assign n19144 = ~n18399 & n34113;
  assign n19145 = ~n18397 & n19144;
  assign n19146 = n34113 & n19142;
  assign n19147 = ~n18472 & n19145;
  assign n19148 = ~n19143 & ~n34203;
  assign n19149 = n214 & ~n19123;
  assign n19150 = n214 & n19139;
  assign n19151 = ~n19138 & n19149;
  assign n19152 = ~n19148 & ~n34204;
  assign n19153 = ~n19140 & ~n19152;
  assign n19154 = ~n197 & ~n19153;
  assign n19155 = ~n18414 & ~n34114;
  assign n19156 = ~n18472 & n19155;
  assign n19157 = ~n34116 & ~n19156;
  assign n19158 = ~n18414 & n34116;
  assign n19159 = ~n34114 & n19158;
  assign n19160 = n34116 & n19156;
  assign n19161 = ~n18472 & n19159;
  assign n19162 = ~n19157 & ~n34205;
  assign n19163 = n197 & ~n19140;
  assign n19164 = ~n19152 & n19163;
  assign n19165 = ~n19162 & ~n19164;
  assign n19166 = ~n19154 & ~n19165;
  assign n19167 = ~n18432 & ~n18434;
  assign n19168 = ~n18472 & n19167;
  assign n19169 = ~n34118 & ~n19168;
  assign n19170 = ~n18434 & n34118;
  assign n19171 = ~n18432 & n19170;
  assign n19172 = n34118 & n19168;
  assign n19173 = ~n18472 & n19171;
  assign n19174 = ~n19169 & ~n34206;
  assign n19175 = ~n18448 & ~n18456;
  assign n19176 = ~n18456 & ~n18472;
  assign n19177 = ~n18448 & n19176;
  assign n19178 = ~n18472 & n19175;
  assign n19179 = ~n34121 & ~n34207;
  assign n19180 = ~n19174 & n19179;
  assign n19181 = ~n19166 & n19180;
  assign n19182 = n193 & ~n19181;
  assign n19183 = ~n19154 & n19174;
  assign n19184 = n19166 & n19174;
  assign n19185 = ~n19165 & n19183;
  assign n19186 = n18448 & ~n19176;
  assign n19187 = ~n193 & ~n19175;
  assign n19188 = ~n19186 & n19187;
  assign n19189 = ~n34208 & ~n19188;
  assign n19190 = ~n19182 & n19189;
  assign n19191 = pi28  & ~n19190;
  assign n19192 = ~pi26  & ~pi27 ;
  assign n19193 = ~pi28  & n19192;
  assign n19194 = ~n19191 & ~n19193;
  assign n19195 = ~n18472 & ~n19194;
  assign n19196 = ~pi28  & ~n19190;
  assign n19197 = pi29  & ~n19196;
  assign n19198 = ~pi29  & n19196;
  assign n19199 = n18646 & ~n19190;
  assign n19200 = ~n19197 & ~n34209;
  assign n19201 = ~n34014 & ~n34144;
  assign n19202 = ~n17669 & n19201;
  assign n19203 = ~n17688 & n19202;
  assign n19204 = ~n34016 & n19203;
  assign n19205 = n17674 & n17690;
  assign n19206 = ~n17682 & n19204;
  assign n19207 = ~n19193 & ~n34210;
  assign n19208 = ~n18470 & n19207;
  assign n19209 = ~n34121 & n19208;
  assign n19210 = ~n18464 & n19209;
  assign n19211 = n18472 & n19194;
  assign n19212 = ~n19191 & n19210;
  assign n19213 = n19200 & ~n34211;
  assign n19214 = ~n19195 & ~n19213;
  assign n19215 = ~n17690 & ~n19214;
  assign n19216 = n17690 & ~n19195;
  assign n19217 = ~n19213 & n19216;
  assign n19218 = ~n18472 & ~n19188;
  assign n19219 = ~n34208 & n19218;
  assign n19220 = ~n19182 & n19219;
  assign n19221 = ~n34209 & ~n19220;
  assign n19222 = pi30  & ~n19221;
  assign n19223 = ~pi30  & ~n19220;
  assign n19224 = ~pi30  & n19221;
  assign n19225 = ~n34209 & n19223;
  assign n19226 = ~n19222 & ~n34212;
  assign n19227 = ~n19217 & ~n19226;
  assign n19228 = ~n19215 & ~n19227;
  assign n19229 = ~n17001 & ~n19228;
  assign n19230 = n17001 & ~n19215;
  assign n19231 = ~n19227 & n19230;
  assign n19232 = n17001 & n19228;
  assign n19233 = ~n34145 & ~n18664;
  assign n19234 = ~n19190 & n19233;
  assign n19235 = n18662 & ~n19234;
  assign n19236 = ~n18662 & n19233;
  assign n19237 = ~n18662 & n19234;
  assign n19238 = ~n19190 & n19236;
  assign n19239 = ~n19235 & ~n34214;
  assign n19240 = ~n34213 & ~n19239;
  assign n19241 = ~n19229 & ~n19240;
  assign n19242 = ~n16248 & ~n19241;
  assign n19243 = n16248 & ~n19229;
  assign n19244 = ~n19240 & n19243;
  assign n19245 = ~n34146 & ~n18670;
  assign n19246 = ~n18670 & ~n19190;
  assign n19247 = ~n34146 & n19246;
  assign n19248 = ~n19190 & n19245;
  assign n19249 = n18644 & ~n34215;
  assign n19250 = n18669 & n19246;
  assign n19251 = n18644 & ~n34146;
  assign n19252 = ~n18670 & n19251;
  assign n19253 = ~n19190 & n19252;
  assign n19254 = ~n18644 & ~n34215;
  assign n19255 = ~n19253 & ~n19254;
  assign n19256 = ~n19249 & ~n19250;
  assign n19257 = ~n19244 & ~n34216;
  assign n19258 = ~n19242 & ~n19257;
  assign n19259 = ~n15586 & ~n19258;
  assign n19260 = n15586 & ~n19242;
  assign n19261 = ~n19257 & n19260;
  assign n19262 = n15586 & n19258;
  assign n19263 = ~n18672 & ~n18682;
  assign n19264 = ~n19190 & n19263;
  assign n19265 = ~n18679 & ~n19264;
  assign n19266 = n18679 & ~n18682;
  assign n19267 = ~n18672 & n19266;
  assign n19268 = n18679 & n19264;
  assign n19269 = ~n19190 & n19267;
  assign n19270 = n18679 & ~n19264;
  assign n19271 = ~n18679 & n19264;
  assign n19272 = ~n19270 & ~n19271;
  assign n19273 = ~n19265 & ~n34218;
  assign n19274 = ~n34217 & n34219;
  assign n19275 = ~n19259 & ~n19274;
  assign n19276 = ~n14866 & ~n19275;
  assign n19277 = n14866 & ~n19259;
  assign n19278 = ~n19274 & n19277;
  assign n19279 = ~n34148 & ~n18688;
  assign n19280 = ~n18688 & ~n19190;
  assign n19281 = ~n34148 & n19280;
  assign n19282 = ~n19190 & n19279;
  assign n19283 = n18632 & ~n34220;
  assign n19284 = n18687 & n19280;
  assign n19285 = n18632 & ~n34148;
  assign n19286 = ~n18688 & n19285;
  assign n19287 = ~n19190 & n19286;
  assign n19288 = ~n18632 & ~n34220;
  assign n19289 = ~n19287 & ~n19288;
  assign n19290 = ~n19283 & ~n19284;
  assign n19291 = ~n19278 & ~n34221;
  assign n19292 = ~n19276 & ~n19291;
  assign n19293 = ~n14233 & ~n19292;
  assign n19294 = n14233 & ~n19276;
  assign n19295 = ~n19291 & n19294;
  assign n19296 = n14233 & n19292;
  assign n19297 = ~n18690 & ~n18704;
  assign n19298 = ~n19190 & n19297;
  assign n19299 = ~n34150 & ~n19298;
  assign n19300 = n34150 & n19298;
  assign n19301 = ~n34150 & ~n18704;
  assign n19302 = ~n18690 & n19301;
  assign n19303 = ~n19190 & n19302;
  assign n19304 = n34150 & ~n19298;
  assign n19305 = ~n19303 & ~n19304;
  assign n19306 = ~n19299 & ~n19300;
  assign n19307 = ~n34222 & ~n34223;
  assign n19308 = ~n19293 & ~n19307;
  assign n19309 = ~n13548 & ~n19308;
  assign n19310 = n13548 & ~n19293;
  assign n19311 = ~n19307 & n19310;
  assign n19312 = ~n34151 & ~n18710;
  assign n19313 = ~n18710 & ~n19190;
  assign n19314 = ~n34151 & n19313;
  assign n19315 = ~n19190 & n19312;
  assign n19316 = n18624 & ~n34224;
  assign n19317 = n18709 & n19313;
  assign n19318 = n18624 & ~n34151;
  assign n19319 = ~n18710 & n19318;
  assign n19320 = ~n19190 & n19319;
  assign n19321 = ~n18624 & ~n34224;
  assign n19322 = ~n19320 & ~n19321;
  assign n19323 = ~n19316 & ~n19317;
  assign n19324 = ~n19311 & ~n34225;
  assign n19325 = ~n19309 & ~n19324;
  assign n19326 = ~n12948 & ~n19325;
  assign n19327 = n12948 & ~n19309;
  assign n19328 = ~n19324 & n19327;
  assign n19329 = n12948 & n19325;
  assign n19330 = ~n18712 & ~n18725;
  assign n19331 = ~n19190 & n19330;
  assign n19332 = ~n34152 & n19331;
  assign n19333 = n34152 & ~n19331;
  assign n19334 = n34152 & ~n18725;
  assign n19335 = ~n18712 & n19334;
  assign n19336 = ~n19190 & n19335;
  assign n19337 = ~n34152 & ~n19331;
  assign n19338 = ~n19336 & ~n19337;
  assign n19339 = ~n19332 & ~n19333;
  assign n19340 = ~n34226 & ~n34227;
  assign n19341 = ~n19326 & ~n19340;
  assign n19342 = ~n12296 & ~n19341;
  assign n19343 = n12296 & ~n19326;
  assign n19344 = ~n19340 & n19343;
  assign n19345 = ~n34153 & ~n18731;
  assign n19346 = ~n18731 & ~n19190;
  assign n19347 = ~n34153 & n19346;
  assign n19348 = ~n19190 & n19345;
  assign n19349 = n18616 & ~n34228;
  assign n19350 = n18730 & n19346;
  assign n19351 = n18616 & ~n34153;
  assign n19352 = ~n18731 & n19351;
  assign n19353 = ~n19190 & n19352;
  assign n19354 = ~n18616 & ~n34228;
  assign n19355 = ~n19353 & ~n19354;
  assign n19356 = ~n19349 & ~n19350;
  assign n19357 = ~n19344 & ~n34229;
  assign n19358 = ~n19342 & ~n19357;
  assign n19359 = ~n11719 & ~n19358;
  assign n19360 = n11719 & ~n19342;
  assign n19361 = ~n19357 & n19360;
  assign n19362 = n11719 & n19358;
  assign n19363 = ~n18733 & ~n18746;
  assign n19364 = ~n19190 & n19363;
  assign n19365 = ~n34154 & n19364;
  assign n19366 = n34154 & ~n19364;
  assign n19367 = ~n34154 & ~n19364;
  assign n19368 = n34154 & ~n18746;
  assign n19369 = ~n18733 & n19368;
  assign n19370 = n34154 & n19364;
  assign n19371 = ~n19190 & n19369;
  assign n19372 = ~n19367 & ~n34231;
  assign n19373 = ~n19365 & ~n19366;
  assign n19374 = ~n34230 & ~n34232;
  assign n19375 = ~n19359 & ~n19374;
  assign n19376 = ~n11097 & ~n19375;
  assign n19377 = n11097 & ~n19359;
  assign n19378 = ~n19374 & n19377;
  assign n19379 = ~n34155 & ~n18752;
  assign n19380 = ~n18752 & ~n19190;
  assign n19381 = ~n34155 & n19380;
  assign n19382 = ~n19190 & n19379;
  assign n19383 = n18608 & ~n34233;
  assign n19384 = n18751 & n19380;
  assign n19385 = n18608 & ~n34155;
  assign n19386 = ~n18752 & n19385;
  assign n19387 = ~n19190 & n19386;
  assign n19388 = ~n18608 & ~n34233;
  assign n19389 = ~n19387 & ~n19388;
  assign n19390 = ~n19383 & ~n19384;
  assign n19391 = ~n19378 & ~n34234;
  assign n19392 = ~n19376 & ~n19391;
  assign n19393 = ~n10555 & ~n19392;
  assign n19394 = n10555 & ~n19376;
  assign n19395 = ~n19391 & n19394;
  assign n19396 = n10555 & n19392;
  assign n19397 = ~n18754 & ~n18768;
  assign n19398 = ~n18768 & ~n19190;
  assign n19399 = ~n18754 & n19398;
  assign n19400 = ~n19190 & n19397;
  assign n19401 = n34157 & ~n34236;
  assign n19402 = n18766 & n19398;
  assign n19403 = ~n34157 & n34236;
  assign n19404 = n34157 & ~n18768;
  assign n19405 = ~n18754 & n19404;
  assign n19406 = ~n19190 & n19405;
  assign n19407 = ~n34157 & ~n34236;
  assign n19408 = ~n19406 & ~n19407;
  assign n19409 = ~n19401 & ~n34237;
  assign n19410 = ~n34235 & ~n34238;
  assign n19411 = ~n19393 & ~n19410;
  assign n19412 = ~n9969 & ~n19411;
  assign n19413 = n9969 & ~n19393;
  assign n19414 = ~n19410 & n19413;
  assign n19415 = ~n34158 & ~n18774;
  assign n19416 = ~n18774 & ~n19190;
  assign n19417 = ~n34158 & n19416;
  assign n19418 = ~n19190 & n19415;
  assign n19419 = n18600 & ~n34239;
  assign n19420 = n18773 & n19416;
  assign n19421 = n18600 & ~n34158;
  assign n19422 = ~n18774 & n19421;
  assign n19423 = ~n19190 & n19422;
  assign n19424 = ~n18600 & ~n34239;
  assign n19425 = ~n19423 & ~n19424;
  assign n19426 = ~n19419 & ~n19420;
  assign n19427 = ~n19414 & ~n34240;
  assign n19428 = ~n19412 & ~n19427;
  assign n19429 = ~n9457 & ~n19428;
  assign n19430 = ~n18776 & ~n18792;
  assign n19431 = ~n19190 & n19430;
  assign n19432 = ~n34161 & ~n19431;
  assign n19433 = n34161 & ~n18792;
  assign n19434 = ~n18776 & n19433;
  assign n19435 = n34161 & n19431;
  assign n19436 = ~n19190 & n19434;
  assign n19437 = ~n19432 & ~n34241;
  assign n19438 = n9457 & ~n19412;
  assign n19439 = ~n19427 & n19438;
  assign n19440 = n9457 & n19428;
  assign n19441 = ~n19437 & ~n34242;
  assign n19442 = ~n19429 & ~n19441;
  assign n19443 = ~n8896 & ~n19442;
  assign n19444 = n8896 & ~n19429;
  assign n19445 = ~n19441 & n19444;
  assign n19446 = ~n34162 & ~n18798;
  assign n19447 = ~n18798 & ~n19190;
  assign n19448 = ~n34162 & n19447;
  assign n19449 = ~n19190 & n19446;
  assign n19450 = n18592 & ~n34243;
  assign n19451 = n18797 & n19447;
  assign n19452 = n18592 & ~n34162;
  assign n19453 = ~n18798 & n19452;
  assign n19454 = ~n19190 & n19453;
  assign n19455 = ~n18592 & ~n34243;
  assign n19456 = ~n19454 & ~n19455;
  assign n19457 = ~n19450 & ~n19451;
  assign n19458 = ~n19445 & ~n34244;
  assign n19459 = ~n19443 & ~n19458;
  assign n19460 = ~n8411 & ~n19459;
  assign n19461 = n8411 & ~n19443;
  assign n19462 = ~n19458 & n19461;
  assign n19463 = n8411 & n19459;
  assign n19464 = ~n18800 & ~n18803;
  assign n19465 = ~n18803 & ~n19190;
  assign n19466 = ~n18800 & n19465;
  assign n19467 = ~n19190 & n19464;
  assign n19468 = n18584 & ~n34246;
  assign n19469 = n18801 & n19465;
  assign n19470 = n18584 & ~n18803;
  assign n19471 = ~n18800 & n19470;
  assign n19472 = ~n19190 & n19471;
  assign n19473 = ~n18584 & ~n34246;
  assign n19474 = ~n19472 & ~n19473;
  assign n19475 = ~n19468 & ~n19469;
  assign n19476 = ~n34245 & ~n34247;
  assign n19477 = ~n19460 & ~n19476;
  assign n19478 = ~n7885 & ~n19477;
  assign n19479 = n7885 & ~n19460;
  assign n19480 = ~n19476 & n19479;
  assign n19481 = ~n34163 & ~n18809;
  assign n19482 = ~n18809 & ~n19190;
  assign n19483 = ~n34163 & n19482;
  assign n19484 = ~n19190 & n19481;
  assign n19485 = n18576 & ~n34248;
  assign n19486 = n18808 & n19482;
  assign n19487 = n18576 & ~n34163;
  assign n19488 = ~n18809 & n19487;
  assign n19489 = ~n19190 & n19488;
  assign n19490 = ~n18576 & ~n34248;
  assign n19491 = ~n19489 & ~n19490;
  assign n19492 = ~n19485 & ~n19486;
  assign n19493 = ~n19480 & ~n34249;
  assign n19494 = ~n19478 & ~n19493;
  assign n19495 = ~n7428 & ~n19494;
  assign n19496 = ~n18811 & ~n18826;
  assign n19497 = ~n19190 & n19496;
  assign n19498 = ~n34165 & ~n19497;
  assign n19499 = n34165 & ~n18826;
  assign n19500 = ~n18811 & n19499;
  assign n19501 = n34165 & n19497;
  assign n19502 = ~n19190 & n19500;
  assign n19503 = ~n19498 & ~n34250;
  assign n19504 = n7428 & ~n19478;
  assign n19505 = ~n19493 & n19504;
  assign n19506 = n7428 & n19494;
  assign n19507 = ~n19503 & ~n34251;
  assign n19508 = ~n19495 & ~n19507;
  assign n19509 = ~n6937 & ~n19508;
  assign n19510 = n6937 & ~n19495;
  assign n19511 = ~n19507 & n19510;
  assign n19512 = ~n34166 & ~n18832;
  assign n19513 = ~n18832 & ~n19190;
  assign n19514 = ~n34166 & n19513;
  assign n19515 = ~n19190 & n19512;
  assign n19516 = n18568 & ~n34252;
  assign n19517 = n18831 & n19513;
  assign n19518 = n18568 & ~n34166;
  assign n19519 = ~n18832 & n19518;
  assign n19520 = ~n19190 & n19519;
  assign n19521 = ~n18568 & ~n34252;
  assign n19522 = ~n19520 & ~n19521;
  assign n19523 = ~n19516 & ~n19517;
  assign n19524 = ~n19511 & ~n34253;
  assign n19525 = ~n19509 & ~n19524;
  assign n19526 = ~n6507 & ~n19525;
  assign n19527 = n6507 & ~n19509;
  assign n19528 = ~n19524 & n19527;
  assign n19529 = n6507 & n19525;
  assign n19530 = ~n18834 & ~n18837;
  assign n19531 = ~n18837 & ~n19190;
  assign n19532 = ~n18834 & n19531;
  assign n19533 = ~n19190 & n19530;
  assign n19534 = n18560 & ~n34255;
  assign n19535 = n18835 & n19531;
  assign n19536 = n18560 & ~n18837;
  assign n19537 = ~n18834 & n19536;
  assign n19538 = ~n19190 & n19537;
  assign n19539 = ~n18560 & ~n34255;
  assign n19540 = ~n19538 & ~n19539;
  assign n19541 = ~n19534 & ~n19535;
  assign n19542 = ~n34254 & ~n34256;
  assign n19543 = ~n19526 & ~n19542;
  assign n19544 = ~n6051 & ~n19543;
  assign n19545 = n6051 & ~n19526;
  assign n19546 = ~n19542 & n19545;
  assign n19547 = ~n34167 & ~n18843;
  assign n19548 = ~n18843 & ~n19190;
  assign n19549 = ~n34167 & n19548;
  assign n19550 = ~n19190 & n19547;
  assign n19551 = n18552 & ~n34257;
  assign n19552 = n18842 & n19548;
  assign n19553 = n18552 & ~n34167;
  assign n19554 = ~n18843 & n19553;
  assign n19555 = ~n19190 & n19554;
  assign n19556 = ~n18552 & ~n34257;
  assign n19557 = ~n19555 & ~n19556;
  assign n19558 = ~n19551 & ~n19552;
  assign n19559 = ~n19546 & ~n34258;
  assign n19560 = ~n19544 & ~n19559;
  assign n19561 = ~n5648 & ~n19560;
  assign n19562 = ~n18845 & ~n18860;
  assign n19563 = ~n19190 & n19562;
  assign n19564 = ~n34169 & ~n19563;
  assign n19565 = n34169 & ~n18860;
  assign n19566 = ~n18845 & n19565;
  assign n19567 = n34169 & n19563;
  assign n19568 = ~n19190 & n19566;
  assign n19569 = ~n19564 & ~n34259;
  assign n19570 = n5648 & ~n19544;
  assign n19571 = ~n19559 & n19570;
  assign n19572 = n5648 & n19560;
  assign n19573 = ~n19569 & ~n34260;
  assign n19574 = ~n19561 & ~n19573;
  assign n19575 = ~n5223 & ~n19574;
  assign n19576 = n5223 & ~n19561;
  assign n19577 = ~n19573 & n19576;
  assign n19578 = ~n34170 & ~n18866;
  assign n19579 = ~n18866 & ~n19190;
  assign n19580 = ~n34170 & n19579;
  assign n19581 = ~n19190 & n19578;
  assign n19582 = n18544 & ~n34261;
  assign n19583 = n18865 & n19579;
  assign n19584 = n18544 & ~n34170;
  assign n19585 = ~n18866 & n19584;
  assign n19586 = ~n19190 & n19585;
  assign n19587 = ~n18544 & ~n34261;
  assign n19588 = ~n19586 & ~n19587;
  assign n19589 = ~n19582 & ~n19583;
  assign n19590 = ~n19577 & ~n34262;
  assign n19591 = ~n19575 & ~n19590;
  assign n19592 = ~n4851 & ~n19591;
  assign n19593 = n4851 & ~n19575;
  assign n19594 = ~n19590 & n19593;
  assign n19595 = n4851 & n19591;
  assign n19596 = ~n18868 & ~n18871;
  assign n19597 = ~n18871 & ~n19190;
  assign n19598 = ~n18868 & n19597;
  assign n19599 = ~n19190 & n19596;
  assign n19600 = n18536 & ~n34264;
  assign n19601 = n18869 & n19597;
  assign n19602 = n18536 & ~n18871;
  assign n19603 = ~n18868 & n19602;
  assign n19604 = ~n19190 & n19603;
  assign n19605 = ~n18536 & ~n34264;
  assign n19606 = ~n19604 & ~n19605;
  assign n19607 = ~n19600 & ~n19601;
  assign n19608 = ~n34263 & ~n34265;
  assign n19609 = ~n19592 & ~n19608;
  assign n19610 = ~n4461 & ~n19609;
  assign n19611 = n4461 & ~n19592;
  assign n19612 = ~n19608 & n19611;
  assign n19613 = ~n34171 & ~n18877;
  assign n19614 = ~n18877 & ~n19190;
  assign n19615 = ~n34171 & n19614;
  assign n19616 = ~n19190 & n19613;
  assign n19617 = n18528 & ~n34266;
  assign n19618 = n18876 & n19614;
  assign n19619 = n18528 & ~n34171;
  assign n19620 = ~n18877 & n19619;
  assign n19621 = ~n19190 & n19620;
  assign n19622 = ~n18528 & ~n34266;
  assign n19623 = ~n19621 & ~n19622;
  assign n19624 = ~n19617 & ~n19618;
  assign n19625 = ~n19612 & ~n34267;
  assign n19626 = ~n19610 & ~n19625;
  assign n19627 = ~n4115 & ~n19626;
  assign n19628 = ~n18879 & ~n18894;
  assign n19629 = ~n19190 & n19628;
  assign n19630 = ~n34173 & ~n19629;
  assign n19631 = n34173 & ~n18894;
  assign n19632 = ~n18879 & n19631;
  assign n19633 = n34173 & n19629;
  assign n19634 = ~n19190 & n19632;
  assign n19635 = ~n19630 & ~n34268;
  assign n19636 = n4115 & ~n19610;
  assign n19637 = ~n19625 & n19636;
  assign n19638 = n4115 & n19626;
  assign n19639 = ~n19635 & ~n34269;
  assign n19640 = ~n19627 & ~n19639;
  assign n19641 = ~n3754 & ~n19640;
  assign n19642 = n3754 & ~n19627;
  assign n19643 = ~n19639 & n19642;
  assign n19644 = ~n34174 & ~n18900;
  assign n19645 = ~n18900 & ~n19190;
  assign n19646 = ~n34174 & n19645;
  assign n19647 = ~n19190 & n19644;
  assign n19648 = n18520 & ~n34270;
  assign n19649 = n18899 & n19645;
  assign n19650 = n18520 & ~n34174;
  assign n19651 = ~n18900 & n19650;
  assign n19652 = ~n19190 & n19651;
  assign n19653 = ~n18520 & ~n34270;
  assign n19654 = ~n19652 & ~n19653;
  assign n19655 = ~n19648 & ~n19649;
  assign n19656 = ~n19643 & ~n34271;
  assign n19657 = ~n19641 & ~n19656;
  assign n19658 = ~n3444 & ~n19657;
  assign n19659 = n3444 & ~n19641;
  assign n19660 = ~n19656 & n19659;
  assign n19661 = n3444 & n19657;
  assign n19662 = ~n18902 & ~n18905;
  assign n19663 = ~n18905 & ~n19190;
  assign n19664 = ~n18902 & n19663;
  assign n19665 = ~n19190 & n19662;
  assign n19666 = n18512 & ~n34273;
  assign n19667 = n18903 & n19663;
  assign n19668 = n18512 & ~n18905;
  assign n19669 = ~n18902 & n19668;
  assign n19670 = ~n19190 & n19669;
  assign n19671 = ~n18512 & ~n34273;
  assign n19672 = ~n19670 & ~n19671;
  assign n19673 = ~n19666 & ~n19667;
  assign n19674 = ~n34272 & ~n34274;
  assign n19675 = ~n19658 & ~n19674;
  assign n19676 = ~n3116 & ~n19675;
  assign n19677 = n3116 & ~n19658;
  assign n19678 = ~n19674 & n19677;
  assign n19679 = ~n34175 & ~n18911;
  assign n19680 = ~n18911 & ~n19190;
  assign n19681 = ~n34175 & n19680;
  assign n19682 = ~n19190 & n19679;
  assign n19683 = n18504 & ~n34275;
  assign n19684 = n18910 & n19680;
  assign n19685 = n18504 & ~n34175;
  assign n19686 = ~n18911 & n19685;
  assign n19687 = ~n19190 & n19686;
  assign n19688 = ~n18504 & ~n34275;
  assign n19689 = ~n19687 & ~n19688;
  assign n19690 = ~n19683 & ~n19684;
  assign n19691 = ~n19678 & ~n34276;
  assign n19692 = ~n19676 & ~n19691;
  assign n19693 = ~n2833 & ~n19692;
  assign n19694 = ~n18913 & ~n18928;
  assign n19695 = ~n19190 & n19694;
  assign n19696 = ~n34177 & ~n19695;
  assign n19697 = n34177 & ~n18928;
  assign n19698 = ~n18913 & n19697;
  assign n19699 = n34177 & n19695;
  assign n19700 = ~n19190 & n19698;
  assign n19701 = ~n19696 & ~n34277;
  assign n19702 = n2833 & ~n19676;
  assign n19703 = ~n19691 & n19702;
  assign n19704 = n2833 & n19692;
  assign n19705 = ~n19701 & ~n34278;
  assign n19706 = ~n19693 & ~n19705;
  assign n19707 = ~n2536 & ~n19706;
  assign n19708 = n2536 & ~n19693;
  assign n19709 = ~n19705 & n19708;
  assign n19710 = ~n34178 & ~n18934;
  assign n19711 = ~n18934 & ~n19190;
  assign n19712 = ~n34178 & n19711;
  assign n19713 = ~n19190 & n19710;
  assign n19714 = n18496 & ~n34279;
  assign n19715 = n18933 & n19711;
  assign n19716 = n18496 & ~n34178;
  assign n19717 = ~n18934 & n19716;
  assign n19718 = ~n19190 & n19717;
  assign n19719 = ~n18496 & ~n34279;
  assign n19720 = ~n19718 & ~n19719;
  assign n19721 = ~n19714 & ~n19715;
  assign n19722 = ~n19709 & ~n34280;
  assign n19723 = ~n19707 & ~n19722;
  assign n19724 = ~n2283 & ~n19723;
  assign n19725 = n2283 & ~n19707;
  assign n19726 = ~n19722 & n19725;
  assign n19727 = n2283 & n19723;
  assign n19728 = ~n18936 & ~n18939;
  assign n19729 = ~n18939 & ~n19190;
  assign n19730 = ~n18936 & n19729;
  assign n19731 = ~n19190 & n19728;
  assign n19732 = n18488 & ~n34282;
  assign n19733 = n18937 & n19729;
  assign n19734 = n18488 & ~n18939;
  assign n19735 = ~n18936 & n19734;
  assign n19736 = ~n19190 & n19735;
  assign n19737 = ~n18488 & ~n34282;
  assign n19738 = ~n19736 & ~n19737;
  assign n19739 = ~n19732 & ~n19733;
  assign n19740 = ~n34281 & ~n34283;
  assign n19741 = ~n19724 & ~n19740;
  assign n19742 = ~n2021 & ~n19741;
  assign n19743 = n2021 & ~n19724;
  assign n19744 = ~n19740 & n19743;
  assign n19745 = ~n34179 & ~n18945;
  assign n19746 = ~n19190 & n19745;
  assign n19747 = n18480 & ~n19746;
  assign n19748 = ~n18480 & n19746;
  assign n19749 = n18480 & ~n34179;
  assign n19750 = ~n18945 & n19749;
  assign n19751 = ~n19190 & n19750;
  assign n19752 = ~n18480 & ~n19746;
  assign n19753 = ~n19751 & ~n19752;
  assign n19754 = ~n19747 & ~n19748;
  assign n19755 = ~n19744 & ~n34284;
  assign n19756 = ~n19742 & ~n19755;
  assign n19757 = ~n1796 & ~n19756;
  assign n19758 = ~n18947 & ~n18959;
  assign n19759 = ~n19190 & n19758;
  assign n19760 = ~n34180 & n19759;
  assign n19761 = n34180 & ~n19759;
  assign n19762 = ~n18947 & n34180;
  assign n19763 = ~n18959 & n19762;
  assign n19764 = ~n19190 & n19763;
  assign n19765 = ~n34180 & ~n19759;
  assign n19766 = ~n19764 & ~n19765;
  assign n19767 = ~n19760 & ~n19761;
  assign n19768 = n1796 & ~n19742;
  assign n19769 = ~n19755 & n19768;
  assign n19770 = n1796 & n19756;
  assign n19771 = ~n34285 & ~n34286;
  assign n19772 = ~n19757 & ~n19771;
  assign n19773 = ~n1567 & ~n19772;
  assign n19774 = n1567 & ~n19757;
  assign n19775 = ~n19771 & n19774;
  assign n19776 = ~n18962 & ~n34182;
  assign n19777 = ~n18962 & ~n19190;
  assign n19778 = ~n34182 & n19777;
  assign n19779 = ~n19190 & n19776;
  assign n19780 = n18970 & ~n34287;
  assign n19781 = n18974 & n19777;
  assign n19782 = n18970 & ~n34182;
  assign n19783 = ~n18962 & n19782;
  assign n19784 = ~n19190 & n19783;
  assign n19785 = ~n18970 & ~n34287;
  assign n19786 = ~n19784 & ~n19785;
  assign n19787 = ~n19780 & ~n19781;
  assign n19788 = ~n19775 & ~n34288;
  assign n19789 = ~n19773 & ~n19788;
  assign n19790 = ~n1374 & ~n19789;
  assign n19791 = ~n18976 & ~n18978;
  assign n19792 = ~n19190 & n19791;
  assign n19793 = ~n34184 & ~n19792;
  assign n19794 = ~n18976 & n34184;
  assign n19795 = ~n18978 & n19794;
  assign n19796 = n34184 & n19792;
  assign n19797 = ~n19190 & n19795;
  assign n19798 = ~n19793 & ~n34289;
  assign n19799 = n1374 & ~n19773;
  assign n19800 = ~n19788 & n19799;
  assign n19801 = n1374 & n19789;
  assign n19802 = ~n19798 & ~n34290;
  assign n19803 = ~n19790 & ~n19802;
  assign n19804 = ~n1179 & ~n19803;
  assign n19805 = n1179 & ~n19790;
  assign n19806 = ~n19802 & n19805;
  assign n19807 = ~n18993 & ~n34186;
  assign n19808 = ~n18993 & ~n19190;
  assign n19809 = ~n34186 & n19808;
  assign n19810 = ~n19190 & n19807;
  assign n19811 = n19001 & ~n34291;
  assign n19812 = n19005 & n19808;
  assign n19813 = n19001 & ~n34186;
  assign n19814 = ~n18993 & n19813;
  assign n19815 = ~n19190 & n19814;
  assign n19816 = ~n19001 & ~n34291;
  assign n19817 = ~n19815 & ~n19816;
  assign n19818 = ~n19811 & ~n19812;
  assign n19819 = ~n19806 & ~n34292;
  assign n19820 = ~n19804 & ~n19819;
  assign n19821 = ~n1016 & ~n19820;
  assign n19822 = ~n19007 & ~n19009;
  assign n19823 = ~n19190 & n19822;
  assign n19824 = ~n34188 & ~n19823;
  assign n19825 = ~n19007 & n34188;
  assign n19826 = ~n19009 & n19825;
  assign n19827 = n34188 & n19823;
  assign n19828 = ~n19190 & n19826;
  assign n19829 = ~n19824 & ~n34293;
  assign n19830 = n1016 & ~n19804;
  assign n19831 = ~n19819 & n19830;
  assign n19832 = n1016 & n19820;
  assign n19833 = ~n19829 & ~n34294;
  assign n19834 = ~n19821 & ~n19833;
  assign n19835 = ~n855 & ~n19834;
  assign n19836 = n855 & ~n19821;
  assign n19837 = ~n19833 & n19836;
  assign n19838 = ~n19024 & ~n34190;
  assign n19839 = ~n19024 & ~n19190;
  assign n19840 = ~n34190 & n19839;
  assign n19841 = ~n19190 & n19838;
  assign n19842 = n19032 & ~n34295;
  assign n19843 = n19036 & n19839;
  assign n19844 = n19032 & ~n34190;
  assign n19845 = ~n19024 & n19844;
  assign n19846 = ~n19190 & n19845;
  assign n19847 = ~n19032 & ~n34295;
  assign n19848 = ~n19846 & ~n19847;
  assign n19849 = ~n19842 & ~n19843;
  assign n19850 = ~n19837 & ~n34296;
  assign n19851 = ~n19835 & ~n19850;
  assign n19852 = ~n720 & ~n19851;
  assign n19853 = n720 & ~n19835;
  assign n19854 = ~n19850 & n19853;
  assign n19855 = n720 & n19851;
  assign n19856 = ~n19038 & ~n19048;
  assign n19857 = ~n19038 & ~n19190;
  assign n19858 = ~n19048 & n19857;
  assign n19859 = ~n19190 & n19856;
  assign n19860 = n19046 & ~n34298;
  assign n19861 = n19049 & n19857;
  assign n19862 = ~n19038 & n19046;
  assign n19863 = ~n19048 & n19862;
  assign n19864 = ~n19190 & n19863;
  assign n19865 = ~n19046 & ~n34298;
  assign n19866 = ~n19864 & ~n19865;
  assign n19867 = ~n19860 & ~n19861;
  assign n19868 = ~n34297 & ~n34299;
  assign n19869 = ~n19852 & ~n19868;
  assign n19870 = ~n592 & ~n19869;
  assign n19871 = n592 & ~n19852;
  assign n19872 = ~n19868 & n19871;
  assign n19873 = ~n19051 & ~n34193;
  assign n19874 = ~n19051 & ~n19190;
  assign n19875 = ~n34193 & n19874;
  assign n19876 = ~n19190 & n19873;
  assign n19877 = n19059 & ~n34300;
  assign n19878 = n19063 & n19874;
  assign n19879 = n19059 & ~n34193;
  assign n19880 = ~n19051 & n19879;
  assign n19881 = ~n19190 & n19880;
  assign n19882 = ~n19059 & ~n34300;
  assign n19883 = ~n19881 & ~n19882;
  assign n19884 = ~n19877 & ~n19878;
  assign n19885 = ~n19872 & ~n34301;
  assign n19886 = ~n19870 & ~n19885;
  assign n19887 = ~n487 & ~n19886;
  assign n19888 = ~n19065 & ~n19067;
  assign n19889 = ~n19190 & n19888;
  assign n19890 = ~n34195 & ~n19889;
  assign n19891 = ~n19065 & n34195;
  assign n19892 = ~n19067 & n19891;
  assign n19893 = n34195 & n19889;
  assign n19894 = ~n19190 & n19892;
  assign n19895 = ~n19890 & ~n34302;
  assign n19896 = n487 & ~n19870;
  assign n19897 = ~n19885 & n19896;
  assign n19898 = n487 & n19886;
  assign n19899 = ~n19895 & ~n34303;
  assign n19900 = ~n19887 & ~n19899;
  assign n19901 = ~n393 & ~n19900;
  assign n19902 = n393 & ~n19887;
  assign n19903 = ~n19899 & n19902;
  assign n19904 = ~n19082 & ~n34197;
  assign n19905 = ~n19082 & ~n19190;
  assign n19906 = ~n34197 & n19905;
  assign n19907 = ~n19190 & n19904;
  assign n19908 = n19090 & ~n34304;
  assign n19909 = n19094 & n19905;
  assign n19910 = n19090 & ~n34197;
  assign n19911 = ~n19082 & n19910;
  assign n19912 = ~n19190 & n19911;
  assign n19913 = ~n19090 & ~n34304;
  assign n19914 = ~n19912 & ~n19913;
  assign n19915 = ~n19908 & ~n19909;
  assign n19916 = ~n19903 & ~n34305;
  assign n19917 = ~n19901 & ~n19916;
  assign n19918 = ~n321 & ~n19917;
  assign n19919 = n321 & ~n19901;
  assign n19920 = ~n19916 & n19919;
  assign n19921 = n321 & n19917;
  assign n19922 = ~n19096 & ~n19106;
  assign n19923 = ~n19096 & ~n19190;
  assign n19924 = ~n19106 & n19923;
  assign n19925 = ~n19190 & n19922;
  assign n19926 = n19104 & ~n34307;
  assign n19927 = n19107 & n19923;
  assign n19928 = ~n19096 & n19104;
  assign n19929 = ~n19106 & n19928;
  assign n19930 = ~n19190 & n19929;
  assign n19931 = ~n19104 & ~n34307;
  assign n19932 = ~n19930 & ~n19931;
  assign n19933 = ~n19926 & ~n19927;
  assign n19934 = ~n34306 & ~n34308;
  assign n19935 = ~n19918 & ~n19934;
  assign n19936 = ~n263 & ~n19935;
  assign n19937 = n263 & ~n19918;
  assign n19938 = ~n19934 & n19937;
  assign n19939 = ~n19109 & ~n34200;
  assign n19940 = ~n19109 & ~n19190;
  assign n19941 = ~n34200 & n19940;
  assign n19942 = ~n19190 & n19939;
  assign n19943 = n19117 & ~n34309;
  assign n19944 = n19121 & n19940;
  assign n19945 = n19117 & ~n34200;
  assign n19946 = ~n19109 & n19945;
  assign n19947 = ~n19190 & n19946;
  assign n19948 = ~n19117 & ~n34309;
  assign n19949 = ~n19947 & ~n19948;
  assign n19950 = ~n19943 & ~n19944;
  assign n19951 = ~n19938 & ~n34310;
  assign n19952 = ~n19936 & ~n19951;
  assign n19953 = ~n214 & ~n19952;
  assign n19954 = ~n19123 & ~n19125;
  assign n19955 = ~n19190 & n19954;
  assign n19956 = ~n34202 & ~n19955;
  assign n19957 = ~n19123 & n34202;
  assign n19958 = ~n19125 & n19957;
  assign n19959 = n34202 & n19955;
  assign n19960 = ~n19190 & n19958;
  assign n19961 = ~n19956 & ~n34311;
  assign n19962 = n214 & ~n19936;
  assign n19963 = ~n19951 & n19962;
  assign n19964 = n214 & n19952;
  assign n19965 = ~n19961 & ~n34312;
  assign n19966 = ~n19953 & ~n19965;
  assign n19967 = ~n197 & ~n19966;
  assign n19968 = n197 & ~n19953;
  assign n19969 = ~n19965 & n19968;
  assign n19970 = ~n19140 & ~n34204;
  assign n19971 = ~n19140 & ~n19190;
  assign n19972 = ~n34204 & n19971;
  assign n19973 = ~n19190 & n19970;
  assign n19974 = n19148 & ~n34313;
  assign n19975 = n19152 & n19971;
  assign n19976 = n19148 & ~n34204;
  assign n19977 = ~n19140 & n19976;
  assign n19978 = ~n19190 & n19977;
  assign n19979 = ~n19148 & ~n34313;
  assign n19980 = ~n19978 & ~n19979;
  assign n19981 = ~n19974 & ~n19975;
  assign n19982 = ~n19969 & ~n34314;
  assign n19983 = ~n19967 & ~n19982;
  assign n19984 = ~n19154 & ~n19164;
  assign n19985 = ~n19154 & ~n19190;
  assign n19986 = ~n19164 & n19985;
  assign n19987 = ~n19190 & n19984;
  assign n19988 = n19162 & ~n34315;
  assign n19989 = n19165 & n19985;
  assign n19990 = ~n19154 & n19162;
  assign n19991 = ~n19164 & n19990;
  assign n19992 = ~n19190 & n19991;
  assign n19993 = ~n19162 & ~n34315;
  assign n19994 = ~n19992 & ~n19993;
  assign n19995 = ~n19988 & ~n19989;
  assign n19996 = ~n19166 & ~n19174;
  assign n19997 = ~n19174 & ~n19190;
  assign n19998 = ~n19166 & n19997;
  assign n19999 = ~n19190 & n19996;
  assign n20000 = ~n34208 & ~n34317;
  assign n20001 = ~n34316 & n20000;
  assign n20002 = ~n19983 & n20001;
  assign n20003 = n193 & ~n20002;
  assign n20004 = ~n19967 & n34316;
  assign n20005 = ~n19982 & n20004;
  assign n20006 = n19983 & n34316;
  assign n20007 = n19166 & ~n19997;
  assign n20008 = ~n193 & ~n19996;
  assign n20009 = ~n20007 & n20008;
  assign n20010 = ~n34318 & ~n20009;
  assign n20011 = ~n20003 & n20010;
  assign n20012 = ~n19724 & ~n34281;
  assign n20013 = ~n20011 & n20012;
  assign n20014 = ~n34283 & ~n20013;
  assign n20015 = ~n19724 & n34283;
  assign n20016 = ~n34281 & n20015;
  assign n20017 = n34283 & n20013;
  assign n20018 = ~n20011 & n20016;
  assign n20019 = ~n20014 & ~n34319;
  assign n20020 = ~n19707 & ~n19709;
  assign n20021 = ~n20011 & n20020;
  assign n20022 = ~n34280 & ~n20021;
  assign n20023 = ~n19709 & n34280;
  assign n20024 = ~n19707 & n20023;
  assign n20025 = n34280 & n20021;
  assign n20026 = ~n20011 & n20024;
  assign n20027 = ~n20022 & ~n34320;
  assign n20028 = ~n19676 & ~n19678;
  assign n20029 = ~n20011 & n20028;
  assign n20030 = ~n34276 & ~n20029;
  assign n20031 = ~n19678 & n34276;
  assign n20032 = ~n19676 & n20031;
  assign n20033 = n34276 & n20029;
  assign n20034 = ~n20011 & n20032;
  assign n20035 = ~n20030 & ~n34321;
  assign n20036 = ~n19658 & ~n34272;
  assign n20037 = ~n20011 & n20036;
  assign n20038 = ~n34274 & ~n20037;
  assign n20039 = ~n19658 & n34274;
  assign n20040 = ~n34272 & n20039;
  assign n20041 = n34274 & n20037;
  assign n20042 = ~n20011 & n20040;
  assign n20043 = ~n20038 & ~n34322;
  assign n20044 = ~n19641 & ~n19643;
  assign n20045 = ~n20011 & n20044;
  assign n20046 = ~n34271 & ~n20045;
  assign n20047 = ~n19643 & n34271;
  assign n20048 = ~n19641 & n20047;
  assign n20049 = n34271 & n20045;
  assign n20050 = ~n20011 & n20048;
  assign n20051 = ~n20046 & ~n34323;
  assign n20052 = ~n19610 & ~n19612;
  assign n20053 = ~n20011 & n20052;
  assign n20054 = ~n34267 & ~n20053;
  assign n20055 = ~n19612 & n34267;
  assign n20056 = ~n19610 & n20055;
  assign n20057 = n34267 & n20053;
  assign n20058 = ~n20011 & n20056;
  assign n20059 = ~n20054 & ~n34324;
  assign n20060 = ~n19592 & ~n34263;
  assign n20061 = ~n20011 & n20060;
  assign n20062 = ~n34265 & ~n20061;
  assign n20063 = ~n19592 & n34265;
  assign n20064 = ~n34263 & n20063;
  assign n20065 = n34265 & n20061;
  assign n20066 = ~n20011 & n20064;
  assign n20067 = ~n20062 & ~n34325;
  assign n20068 = ~n19575 & ~n19577;
  assign n20069 = ~n20011 & n20068;
  assign n20070 = ~n34262 & ~n20069;
  assign n20071 = ~n19577 & n34262;
  assign n20072 = ~n19575 & n20071;
  assign n20073 = n34262 & n20069;
  assign n20074 = ~n20011 & n20072;
  assign n20075 = ~n20070 & ~n34326;
  assign n20076 = ~n19544 & ~n19546;
  assign n20077 = ~n20011 & n20076;
  assign n20078 = ~n34258 & ~n20077;
  assign n20079 = ~n19546 & n34258;
  assign n20080 = ~n19544 & n20079;
  assign n20081 = n34258 & n20077;
  assign n20082 = ~n20011 & n20080;
  assign n20083 = ~n20078 & ~n34327;
  assign n20084 = ~n19526 & ~n34254;
  assign n20085 = ~n20011 & n20084;
  assign n20086 = ~n34256 & ~n20085;
  assign n20087 = ~n19526 & n34256;
  assign n20088 = ~n34254 & n20087;
  assign n20089 = n34256 & n20085;
  assign n20090 = ~n20011 & n20088;
  assign n20091 = ~n20086 & ~n34328;
  assign n20092 = ~n19509 & ~n19511;
  assign n20093 = ~n20011 & n20092;
  assign n20094 = ~n34253 & ~n20093;
  assign n20095 = ~n19511 & n34253;
  assign n20096 = ~n19509 & n20095;
  assign n20097 = n34253 & n20093;
  assign n20098 = ~n20011 & n20096;
  assign n20099 = ~n20094 & ~n34329;
  assign n20100 = ~n19478 & ~n19480;
  assign n20101 = ~n20011 & n20100;
  assign n20102 = ~n34249 & ~n20101;
  assign n20103 = ~n19480 & n34249;
  assign n20104 = ~n19478 & n20103;
  assign n20105 = n34249 & n20101;
  assign n20106 = ~n20011 & n20104;
  assign n20107 = ~n20102 & ~n34330;
  assign n20108 = ~n19460 & ~n34245;
  assign n20109 = ~n20011 & n20108;
  assign n20110 = ~n34247 & ~n20109;
  assign n20111 = ~n19460 & n34247;
  assign n20112 = ~n34245 & n20111;
  assign n20113 = n34247 & n20109;
  assign n20114 = ~n20011 & n20112;
  assign n20115 = ~n20110 & ~n34331;
  assign n20116 = ~n19443 & ~n19445;
  assign n20117 = ~n20011 & n20116;
  assign n20118 = ~n34244 & ~n20117;
  assign n20119 = ~n19445 & n34244;
  assign n20120 = ~n19443 & n20119;
  assign n20121 = n34244 & n20117;
  assign n20122 = ~n20011 & n20120;
  assign n20123 = ~n20118 & ~n34332;
  assign n20124 = ~n19412 & ~n19414;
  assign n20125 = ~n20011 & n20124;
  assign n20126 = ~n34240 & ~n20125;
  assign n20127 = ~n19414 & n34240;
  assign n20128 = ~n19412 & n20127;
  assign n20129 = n34240 & n20125;
  assign n20130 = ~n20011 & n20128;
  assign n20131 = ~n20126 & ~n34333;
  assign n20132 = ~n19393 & ~n34235;
  assign n20133 = ~n20011 & n20132;
  assign n20134 = ~n34238 & ~n20133;
  assign n20135 = ~n19393 & n34238;
  assign n20136 = ~n34235 & n20135;
  assign n20137 = n34238 & n20133;
  assign n20138 = ~n20011 & n20136;
  assign n20139 = ~n20134 & ~n34334;
  assign n20140 = ~n19376 & ~n19378;
  assign n20141 = ~n20011 & n20140;
  assign n20142 = ~n34234 & ~n20141;
  assign n20143 = ~n19378 & n34234;
  assign n20144 = ~n19376 & n20143;
  assign n20145 = n34234 & n20141;
  assign n20146 = ~n20011 & n20144;
  assign n20147 = ~n20142 & ~n34335;
  assign n20148 = ~n19342 & ~n19344;
  assign n20149 = ~n20011 & n20148;
  assign n20150 = ~n34229 & ~n20149;
  assign n20151 = ~n19344 & n34229;
  assign n20152 = ~n19342 & n20151;
  assign n20153 = n34229 & n20149;
  assign n20154 = ~n20011 & n20152;
  assign n20155 = ~n20150 & ~n34336;
  assign n20156 = ~n19309 & ~n19311;
  assign n20157 = ~n20011 & n20156;
  assign n20158 = ~n34225 & ~n20157;
  assign n20159 = ~n19311 & n34225;
  assign n20160 = ~n19309 & n20159;
  assign n20161 = n34225 & n20157;
  assign n20162 = ~n20011 & n20160;
  assign n20163 = ~n20158 & ~n34337;
  assign n20164 = ~n19276 & ~n19278;
  assign n20165 = ~n20011 & n20164;
  assign n20166 = ~n34221 & ~n20165;
  assign n20167 = ~n19278 & n34221;
  assign n20168 = ~n19276 & n20167;
  assign n20169 = n34221 & n20165;
  assign n20170 = ~n20011 & n20168;
  assign n20171 = ~n20166 & ~n34338;
  assign n20172 = ~n19242 & ~n19244;
  assign n20173 = ~n20011 & n20172;
  assign n20174 = ~n34216 & ~n20173;
  assign n20175 = ~n19244 & n34216;
  assign n20176 = ~n19242 & n20175;
  assign n20177 = n34216 & n20173;
  assign n20178 = ~n20011 & n20176;
  assign n20179 = ~n20174 & ~n34339;
  assign n20180 = ~n19215 & ~n19217;
  assign n20181 = ~n20011 & n20180;
  assign n20182 = ~n19226 & ~n20181;
  assign n20183 = ~n19217 & n19226;
  assign n20184 = ~n19215 & n20183;
  assign n20185 = n19226 & n20181;
  assign n20186 = ~n20011 & n20184;
  assign n20187 = ~n20182 & ~n34340;
  assign n20188 = ~pi26  & ~n20011;
  assign n20189 = ~pi27  & n20188;
  assign n20190 = n19192 & ~n20011;
  assign n20191 = ~n19190 & ~n20009;
  assign n20192 = ~n34318 & n20191;
  assign n20193 = ~n20003 & n20192;
  assign n20194 = ~n34341 & ~n20193;
  assign n20195 = pi28  & ~n20194;
  assign n20196 = ~pi28  & ~n20193;
  assign n20197 = ~pi28  & n20194;
  assign n20198 = ~n34341 & n20196;
  assign n20199 = ~n20195 & ~n34342;
  assign n20200 = pi26  & ~n20011;
  assign n20201 = ~pi24  & ~pi25 ;
  assign n20202 = ~pi26  & n20201;
  assign n20203 = ~n34119 & ~n34210;
  assign n20204 = ~n18451 & n20203;
  assign n20205 = ~n18470 & n20204;
  assign n20206 = ~n34121 & n20205;
  assign n20207 = n18456 & n18472;
  assign n20208 = ~n18464 & n20206;
  assign n20209 = ~n20202 & ~n34343;
  assign n20210 = ~n19188 & n20209;
  assign n20211 = ~n34208 & n20210;
  assign n20212 = ~n19182 & n20211;
  assign n20213 = ~n20200 & ~n20202;
  assign n20214 = n19190 & n20213;
  assign n20215 = ~n20200 & n20212;
  assign n20216 = pi27  & ~n20188;
  assign n20217 = ~n34341 & ~n20216;
  assign n20218 = ~n34344 & n20217;
  assign n20219 = ~n19190 & ~n20213;
  assign n20220 = n18472 & ~n20219;
  assign n20221 = ~n20218 & ~n20219;
  assign n20222 = n18472 & n20221;
  assign n20223 = ~n20218 & n20220;
  assign n20224 = ~n20199 & ~n34345;
  assign n20225 = ~n18472 & ~n20221;
  assign n20226 = n17690 & ~n20225;
  assign n20227 = ~n20224 & n20226;
  assign n20228 = ~n19195 & ~n34211;
  assign n20229 = ~n20011 & n20228;
  assign n20230 = n19200 & ~n20229;
  assign n20231 = ~n19200 & n20228;
  assign n20232 = ~n19200 & n20229;
  assign n20233 = ~n20011 & n20231;
  assign n20234 = ~n20230 & ~n34346;
  assign n20235 = ~n20227 & ~n20234;
  assign n20236 = ~n20224 & ~n20225;
  assign n20237 = ~n17690 & ~n20236;
  assign n20238 = n17001 & ~n20237;
  assign n20239 = ~n20235 & ~n20237;
  assign n20240 = n17001 & n20239;
  assign n20241 = ~n20235 & n20238;
  assign n20242 = ~n20187 & ~n34347;
  assign n20243 = ~n17001 & ~n20239;
  assign n20244 = n16248 & ~n20243;
  assign n20245 = ~n20242 & n20244;
  assign n20246 = ~n19229 & ~n34213;
  assign n20247 = ~n20011 & n20246;
  assign n20248 = ~n19239 & ~n20247;
  assign n20249 = ~n19229 & n19239;
  assign n20250 = ~n34213 & n20249;
  assign n20251 = n19239 & n20247;
  assign n20252 = ~n20011 & n20250;
  assign n20253 = n19239 & ~n20247;
  assign n20254 = ~n19239 & n20247;
  assign n20255 = ~n20253 & ~n20254;
  assign n20256 = ~n20248 & ~n34348;
  assign n20257 = ~n20245 & n34349;
  assign n20258 = ~n20242 & ~n20243;
  assign n20259 = ~n16248 & ~n20258;
  assign n20260 = n15586 & ~n20259;
  assign n20261 = ~n20257 & ~n20259;
  assign n20262 = n15586 & n20261;
  assign n20263 = ~n20257 & n20260;
  assign n20264 = ~n20179 & ~n34350;
  assign n20265 = ~n15586 & ~n20261;
  assign n20266 = n14866 & ~n20265;
  assign n20267 = ~n20264 & n20266;
  assign n20268 = ~n19259 & ~n34217;
  assign n20269 = ~n20011 & n20268;
  assign n20270 = ~n34219 & ~n20269;
  assign n20271 = n34219 & n20269;
  assign n20272 = ~n19259 & ~n34219;
  assign n20273 = ~n34217 & n20272;
  assign n20274 = ~n20011 & n20273;
  assign n20275 = n34219 & ~n20269;
  assign n20276 = ~n20274 & ~n20275;
  assign n20277 = ~n20270 & ~n20271;
  assign n20278 = ~n20267 & ~n34351;
  assign n20279 = ~n20264 & ~n20265;
  assign n20280 = ~n14866 & ~n20279;
  assign n20281 = n14233 & ~n20280;
  assign n20282 = ~n20278 & ~n20280;
  assign n20283 = n14233 & n20282;
  assign n20284 = ~n20278 & n20281;
  assign n20285 = ~n20171 & ~n34352;
  assign n20286 = ~n14233 & ~n20282;
  assign n20287 = n13548 & ~n20286;
  assign n20288 = ~n20285 & n20287;
  assign n20289 = ~n19293 & ~n34222;
  assign n20290 = ~n20011 & n20289;
  assign n20291 = ~n34223 & n20290;
  assign n20292 = n34223 & ~n20290;
  assign n20293 = ~n19293 & n34223;
  assign n20294 = ~n34222 & n20293;
  assign n20295 = ~n20011 & n20294;
  assign n20296 = ~n34223 & ~n20290;
  assign n20297 = ~n20295 & ~n20296;
  assign n20298 = ~n20291 & ~n20292;
  assign n20299 = ~n20288 & ~n34353;
  assign n20300 = ~n20285 & ~n20286;
  assign n20301 = ~n13548 & ~n20300;
  assign n20302 = n12948 & ~n20301;
  assign n20303 = ~n20299 & ~n20301;
  assign n20304 = n12948 & n20303;
  assign n20305 = ~n20299 & n20302;
  assign n20306 = ~n20163 & ~n34354;
  assign n20307 = ~n12948 & ~n20303;
  assign n20308 = n12296 & ~n20307;
  assign n20309 = ~n20306 & n20308;
  assign n20310 = ~n19326 & ~n34226;
  assign n20311 = ~n20011 & n20310;
  assign n20312 = ~n34227 & n20311;
  assign n20313 = n34227 & ~n20311;
  assign n20314 = ~n34227 & ~n20311;
  assign n20315 = ~n19326 & n34227;
  assign n20316 = ~n34226 & n20315;
  assign n20317 = n34227 & n20311;
  assign n20318 = ~n20011 & n20316;
  assign n20319 = ~n20314 & ~n34355;
  assign n20320 = ~n20312 & ~n20313;
  assign n20321 = ~n20309 & ~n34356;
  assign n20322 = ~n20306 & ~n20307;
  assign n20323 = ~n12296 & ~n20322;
  assign n20324 = n11719 & ~n20323;
  assign n20325 = ~n20321 & ~n20323;
  assign n20326 = n11719 & n20325;
  assign n20327 = ~n20321 & n20324;
  assign n20328 = ~n20155 & ~n34357;
  assign n20329 = ~n11719 & ~n20325;
  assign n20330 = n11097 & ~n20329;
  assign n20331 = ~n20328 & n20330;
  assign n20332 = ~n19359 & ~n34230;
  assign n20333 = ~n19359 & ~n20011;
  assign n20334 = ~n34230 & n20333;
  assign n20335 = ~n20011 & n20332;
  assign n20336 = n34232 & ~n34358;
  assign n20337 = n19374 & n20333;
  assign n20338 = ~n34232 & n34358;
  assign n20339 = ~n19359 & n34232;
  assign n20340 = ~n34230 & n20339;
  assign n20341 = ~n20011 & n20340;
  assign n20342 = ~n34232 & ~n34358;
  assign n20343 = ~n20341 & ~n20342;
  assign n20344 = ~n20336 & ~n34359;
  assign n20345 = ~n20331 & ~n34360;
  assign n20346 = ~n20328 & ~n20329;
  assign n20347 = ~n11097 & ~n20346;
  assign n20348 = n10555 & ~n20347;
  assign n20349 = ~n20345 & ~n20347;
  assign n20350 = n10555 & n20349;
  assign n20351 = ~n20345 & n20348;
  assign n20352 = ~n20147 & ~n34361;
  assign n20353 = ~n10555 & ~n20349;
  assign n20354 = n9969 & ~n20353;
  assign n20355 = ~n20352 & n20354;
  assign n20356 = ~n20139 & ~n20355;
  assign n20357 = ~n20352 & ~n20353;
  assign n20358 = ~n9969 & ~n20357;
  assign n20359 = n9457 & ~n20358;
  assign n20360 = ~n20356 & ~n20358;
  assign n20361 = n9457 & n20360;
  assign n20362 = ~n20356 & n20359;
  assign n20363 = ~n20131 & ~n34362;
  assign n20364 = ~n9457 & ~n20360;
  assign n20365 = n8896 & ~n20364;
  assign n20366 = ~n20363 & n20365;
  assign n20367 = ~n19429 & ~n34242;
  assign n20368 = ~n19429 & ~n20011;
  assign n20369 = ~n34242 & n20368;
  assign n20370 = ~n20011 & n20367;
  assign n20371 = n19437 & ~n34363;
  assign n20372 = n19441 & n20368;
  assign n20373 = ~n19429 & n19437;
  assign n20374 = ~n34242 & n20373;
  assign n20375 = ~n20011 & n20374;
  assign n20376 = ~n19437 & ~n34363;
  assign n20377 = ~n20375 & ~n20376;
  assign n20378 = ~n20371 & ~n20372;
  assign n20379 = ~n20366 & ~n34364;
  assign n20380 = ~n20363 & ~n20364;
  assign n20381 = ~n8896 & ~n20380;
  assign n20382 = n8411 & ~n20381;
  assign n20383 = ~n20379 & ~n20381;
  assign n20384 = n8411 & n20383;
  assign n20385 = ~n20379 & n20382;
  assign n20386 = ~n20123 & ~n34365;
  assign n20387 = ~n8411 & ~n20383;
  assign n20388 = n7885 & ~n20387;
  assign n20389 = ~n20386 & n20388;
  assign n20390 = ~n20115 & ~n20389;
  assign n20391 = ~n20386 & ~n20387;
  assign n20392 = ~n7885 & ~n20391;
  assign n20393 = n7428 & ~n20392;
  assign n20394 = ~n20390 & ~n20392;
  assign n20395 = n7428 & n20394;
  assign n20396 = ~n20390 & n20393;
  assign n20397 = ~n20107 & ~n34366;
  assign n20398 = ~n7428 & ~n20394;
  assign n20399 = n6937 & ~n20398;
  assign n20400 = ~n20397 & n20399;
  assign n20401 = ~n19495 & ~n34251;
  assign n20402 = ~n19495 & ~n20011;
  assign n20403 = ~n34251 & n20402;
  assign n20404 = ~n20011 & n20401;
  assign n20405 = n19503 & ~n34367;
  assign n20406 = n19507 & n20402;
  assign n20407 = ~n19495 & n19503;
  assign n20408 = ~n34251 & n20407;
  assign n20409 = ~n20011 & n20408;
  assign n20410 = ~n19503 & ~n34367;
  assign n20411 = ~n20409 & ~n20410;
  assign n20412 = ~n20405 & ~n20406;
  assign n20413 = ~n20400 & ~n34368;
  assign n20414 = ~n20397 & ~n20398;
  assign n20415 = ~n6937 & ~n20414;
  assign n20416 = n6507 & ~n20415;
  assign n20417 = ~n20413 & ~n20415;
  assign n20418 = n6507 & n20417;
  assign n20419 = ~n20413 & n20416;
  assign n20420 = ~n20099 & ~n34369;
  assign n20421 = ~n6507 & ~n20417;
  assign n20422 = n6051 & ~n20421;
  assign n20423 = ~n20420 & n20422;
  assign n20424 = ~n20091 & ~n20423;
  assign n20425 = ~n20420 & ~n20421;
  assign n20426 = ~n6051 & ~n20425;
  assign n20427 = n5648 & ~n20426;
  assign n20428 = ~n20424 & ~n20426;
  assign n20429 = n5648 & n20428;
  assign n20430 = ~n20424 & n20427;
  assign n20431 = ~n20083 & ~n34370;
  assign n20432 = ~n5648 & ~n20428;
  assign n20433 = n5223 & ~n20432;
  assign n20434 = ~n20431 & n20433;
  assign n20435 = ~n19561 & ~n34260;
  assign n20436 = ~n19561 & ~n20011;
  assign n20437 = ~n34260 & n20436;
  assign n20438 = ~n20011 & n20435;
  assign n20439 = n19569 & ~n34371;
  assign n20440 = n19573 & n20436;
  assign n20441 = ~n19561 & n19569;
  assign n20442 = ~n34260 & n20441;
  assign n20443 = ~n20011 & n20442;
  assign n20444 = ~n19569 & ~n34371;
  assign n20445 = ~n20443 & ~n20444;
  assign n20446 = ~n20439 & ~n20440;
  assign n20447 = ~n20434 & ~n34372;
  assign n20448 = ~n20431 & ~n20432;
  assign n20449 = ~n5223 & ~n20448;
  assign n20450 = n4851 & ~n20449;
  assign n20451 = ~n20447 & ~n20449;
  assign n20452 = n4851 & n20451;
  assign n20453 = ~n20447 & n20450;
  assign n20454 = ~n20075 & ~n34373;
  assign n20455 = ~n4851 & ~n20451;
  assign n20456 = n4461 & ~n20455;
  assign n20457 = ~n20454 & n20456;
  assign n20458 = ~n20067 & ~n20457;
  assign n20459 = ~n20454 & ~n20455;
  assign n20460 = ~n4461 & ~n20459;
  assign n20461 = n4115 & ~n20460;
  assign n20462 = ~n20458 & ~n20460;
  assign n20463 = n4115 & n20462;
  assign n20464 = ~n20458 & n20461;
  assign n20465 = ~n20059 & ~n34374;
  assign n20466 = ~n4115 & ~n20462;
  assign n20467 = n3754 & ~n20466;
  assign n20468 = ~n20465 & n20467;
  assign n20469 = ~n19627 & ~n34269;
  assign n20470 = ~n19627 & ~n20011;
  assign n20471 = ~n34269 & n20470;
  assign n20472 = ~n20011 & n20469;
  assign n20473 = n19635 & ~n34375;
  assign n20474 = n19639 & n20470;
  assign n20475 = ~n19627 & n19635;
  assign n20476 = ~n34269 & n20475;
  assign n20477 = ~n20011 & n20476;
  assign n20478 = ~n19635 & ~n34375;
  assign n20479 = ~n20477 & ~n20478;
  assign n20480 = ~n20473 & ~n20474;
  assign n20481 = ~n20468 & ~n34376;
  assign n20482 = ~n20465 & ~n20466;
  assign n20483 = ~n3754 & ~n20482;
  assign n20484 = n3444 & ~n20483;
  assign n20485 = ~n20481 & ~n20483;
  assign n20486 = n3444 & n20485;
  assign n20487 = ~n20481 & n20484;
  assign n20488 = ~n20051 & ~n34377;
  assign n20489 = ~n3444 & ~n20485;
  assign n20490 = n3116 & ~n20489;
  assign n20491 = ~n20488 & n20490;
  assign n20492 = ~n20043 & ~n20491;
  assign n20493 = ~n20488 & ~n20489;
  assign n20494 = ~n3116 & ~n20493;
  assign n20495 = n2833 & ~n20494;
  assign n20496 = ~n20492 & ~n20494;
  assign n20497 = n2833 & n20496;
  assign n20498 = ~n20492 & n20495;
  assign n20499 = ~n20035 & ~n34378;
  assign n20500 = ~n2833 & ~n20496;
  assign n20501 = n2536 & ~n20500;
  assign n20502 = ~n20499 & n20501;
  assign n20503 = ~n19693 & ~n34278;
  assign n20504 = ~n19693 & ~n20011;
  assign n20505 = ~n34278 & n20504;
  assign n20506 = ~n20011 & n20503;
  assign n20507 = n19701 & ~n34379;
  assign n20508 = n19705 & n20504;
  assign n20509 = ~n19693 & n19701;
  assign n20510 = ~n34278 & n20509;
  assign n20511 = ~n20011 & n20510;
  assign n20512 = ~n19701 & ~n34379;
  assign n20513 = ~n20511 & ~n20512;
  assign n20514 = ~n20507 & ~n20508;
  assign n20515 = ~n20502 & ~n34380;
  assign n20516 = ~n20499 & ~n20500;
  assign n20517 = ~n2536 & ~n20516;
  assign n20518 = n2283 & ~n20517;
  assign n20519 = ~n20515 & ~n20517;
  assign n20520 = n2283 & n20519;
  assign n20521 = ~n20515 & n20518;
  assign n20522 = ~n20027 & ~n34381;
  assign n20523 = ~n2283 & ~n20519;
  assign n20524 = n2021 & ~n20523;
  assign n20525 = ~n20522 & n20524;
  assign n20526 = ~n20019 & ~n20525;
  assign n20527 = ~n20522 & ~n20523;
  assign n20528 = ~n2021 & ~n20527;
  assign n20529 = n1796 & ~n20528;
  assign n20530 = ~n20526 & ~n20528;
  assign n20531 = n1796 & n20530;
  assign n20532 = ~n20526 & n20529;
  assign n20533 = ~n19742 & ~n19744;
  assign n20534 = ~n20011 & n20533;
  assign n20535 = ~n34284 & n20534;
  assign n20536 = n34284 & ~n20534;
  assign n20537 = ~n19744 & n34284;
  assign n20538 = ~n19742 & n20537;
  assign n20539 = ~n20011 & n20538;
  assign n20540 = ~n34284 & ~n20534;
  assign n20541 = ~n20539 & ~n20540;
  assign n20542 = ~n20535 & ~n20536;
  assign n20543 = ~n34382 & ~n34383;
  assign n20544 = ~n1796 & ~n20530;
  assign n20545 = ~n20543 & ~n20544;
  assign n20546 = ~n1567 & ~n20545;
  assign n20547 = ~n19757 & ~n34286;
  assign n20548 = ~n20011 & n20547;
  assign n20549 = n34285 & ~n20548;
  assign n20550 = ~n34285 & n20548;
  assign n20551 = ~n19757 & n34285;
  assign n20552 = ~n34286 & n20551;
  assign n20553 = ~n20011 & n20552;
  assign n20554 = ~n34285 & ~n20548;
  assign n20555 = ~n20553 & ~n20554;
  assign n20556 = ~n20549 & ~n20550;
  assign n20557 = n1567 & ~n20544;
  assign n20558 = ~n20543 & n20557;
  assign n20559 = ~n34384 & ~n20558;
  assign n20560 = ~n20546 & ~n20559;
  assign n20561 = ~n1374 & ~n20560;
  assign n20562 = ~n19773 & ~n19775;
  assign n20563 = ~n20011 & n20562;
  assign n20564 = ~n34288 & ~n20563;
  assign n20565 = ~n19775 & n34288;
  assign n20566 = ~n19773 & n20565;
  assign n20567 = n34288 & n20563;
  assign n20568 = ~n20011 & n20566;
  assign n20569 = ~n20564 & ~n34385;
  assign n20570 = n1374 & ~n20546;
  assign n20571 = n1374 & n20560;
  assign n20572 = ~n20559 & n20570;
  assign n20573 = ~n20569 & ~n34386;
  assign n20574 = ~n20561 & ~n20573;
  assign n20575 = ~n1179 & ~n20574;
  assign n20576 = n1179 & ~n20561;
  assign n20577 = ~n20573 & n20576;
  assign n20578 = ~n19790 & ~n34290;
  assign n20579 = ~n19790 & ~n20011;
  assign n20580 = ~n34290 & n20579;
  assign n20581 = ~n20011 & n20578;
  assign n20582 = n19798 & ~n34387;
  assign n20583 = n19802 & n20579;
  assign n20584 = ~n19790 & n19798;
  assign n20585 = ~n34290 & n20584;
  assign n20586 = ~n20011 & n20585;
  assign n20587 = ~n19798 & ~n34387;
  assign n20588 = ~n20586 & ~n20587;
  assign n20589 = ~n20582 & ~n20583;
  assign n20590 = ~n20577 & ~n34388;
  assign n20591 = ~n20575 & ~n20590;
  assign n20592 = ~n1016 & ~n20591;
  assign n20593 = ~n19804 & ~n19806;
  assign n20594 = ~n20011 & n20593;
  assign n20595 = ~n34292 & ~n20594;
  assign n20596 = ~n19806 & n34292;
  assign n20597 = ~n19804 & n20596;
  assign n20598 = n34292 & n20594;
  assign n20599 = ~n20011 & n20597;
  assign n20600 = ~n20595 & ~n34389;
  assign n20601 = n1016 & ~n20575;
  assign n20602 = n1016 & n20591;
  assign n20603 = ~n20590 & n20601;
  assign n20604 = ~n20600 & ~n34390;
  assign n20605 = ~n20592 & ~n20604;
  assign n20606 = ~n855 & ~n20605;
  assign n20607 = n855 & ~n20592;
  assign n20608 = ~n20604 & n20607;
  assign n20609 = ~n19821 & ~n34294;
  assign n20610 = ~n19821 & ~n20011;
  assign n20611 = ~n34294 & n20610;
  assign n20612 = ~n20011 & n20609;
  assign n20613 = n19829 & ~n34391;
  assign n20614 = n19833 & n20610;
  assign n20615 = ~n19821 & n19829;
  assign n20616 = ~n34294 & n20615;
  assign n20617 = ~n20011 & n20616;
  assign n20618 = ~n19829 & ~n34391;
  assign n20619 = ~n20617 & ~n20618;
  assign n20620 = ~n20613 & ~n20614;
  assign n20621 = ~n20608 & ~n34392;
  assign n20622 = ~n20606 & ~n20621;
  assign n20623 = ~n720 & ~n20622;
  assign n20624 = ~n19835 & ~n19837;
  assign n20625 = ~n20011 & n20624;
  assign n20626 = ~n34296 & ~n20625;
  assign n20627 = ~n19837 & n34296;
  assign n20628 = ~n19835 & n20627;
  assign n20629 = n34296 & n20625;
  assign n20630 = ~n20011 & n20628;
  assign n20631 = ~n20626 & ~n34393;
  assign n20632 = n720 & ~n20606;
  assign n20633 = n720 & n20622;
  assign n20634 = ~n20621 & n20632;
  assign n20635 = ~n20631 & ~n34394;
  assign n20636 = ~n20623 & ~n20635;
  assign n20637 = ~n592 & ~n20636;
  assign n20638 = ~n19852 & ~n34297;
  assign n20639 = ~n20011 & n20638;
  assign n20640 = ~n34299 & ~n20639;
  assign n20641 = ~n19852 & n34299;
  assign n20642 = ~n34297 & n20641;
  assign n20643 = n34299 & n20639;
  assign n20644 = ~n20011 & n20642;
  assign n20645 = ~n20640 & ~n34395;
  assign n20646 = n592 & ~n20623;
  assign n20647 = ~n20635 & n20646;
  assign n20648 = ~n20645 & ~n20647;
  assign n20649 = ~n20637 & ~n20648;
  assign n20650 = ~n487 & ~n20649;
  assign n20651 = ~n19870 & ~n19872;
  assign n20652 = ~n20011 & n20651;
  assign n20653 = ~n34301 & ~n20652;
  assign n20654 = ~n19872 & n34301;
  assign n20655 = ~n19870 & n20654;
  assign n20656 = n34301 & n20652;
  assign n20657 = ~n20011 & n20655;
  assign n20658 = ~n20653 & ~n34396;
  assign n20659 = n487 & ~n20637;
  assign n20660 = n487 & n20649;
  assign n20661 = ~n20648 & n20659;
  assign n20662 = ~n20658 & ~n34397;
  assign n20663 = ~n20650 & ~n20662;
  assign n20664 = ~n393 & ~n20663;
  assign n20665 = n393 & ~n20650;
  assign n20666 = ~n20662 & n20665;
  assign n20667 = ~n19887 & ~n34303;
  assign n20668 = ~n19887 & ~n20011;
  assign n20669 = ~n34303 & n20668;
  assign n20670 = ~n20011 & n20667;
  assign n20671 = n19895 & ~n34398;
  assign n20672 = n19899 & n20668;
  assign n20673 = ~n19887 & n19895;
  assign n20674 = ~n34303 & n20673;
  assign n20675 = ~n20011 & n20674;
  assign n20676 = ~n19895 & ~n34398;
  assign n20677 = ~n20675 & ~n20676;
  assign n20678 = ~n20671 & ~n20672;
  assign n20679 = ~n20666 & ~n34399;
  assign n20680 = ~n20664 & ~n20679;
  assign n20681 = ~n321 & ~n20680;
  assign n20682 = ~n19901 & ~n19903;
  assign n20683 = ~n20011 & n20682;
  assign n20684 = ~n34305 & ~n20683;
  assign n20685 = ~n19903 & n34305;
  assign n20686 = ~n19901 & n20685;
  assign n20687 = n34305 & n20683;
  assign n20688 = ~n20011 & n20686;
  assign n20689 = ~n20684 & ~n34400;
  assign n20690 = n321 & ~n20664;
  assign n20691 = n321 & n20680;
  assign n20692 = ~n20679 & n20690;
  assign n20693 = ~n20689 & ~n34401;
  assign n20694 = ~n20681 & ~n20693;
  assign n20695 = ~n263 & ~n20694;
  assign n20696 = ~n19918 & ~n34306;
  assign n20697 = ~n20011 & n20696;
  assign n20698 = ~n34308 & ~n20697;
  assign n20699 = ~n19918 & n34308;
  assign n20700 = ~n34306 & n20699;
  assign n20701 = n34308 & n20697;
  assign n20702 = ~n20011 & n20700;
  assign n20703 = ~n20698 & ~n34402;
  assign n20704 = n263 & ~n20681;
  assign n20705 = ~n20693 & n20704;
  assign n20706 = ~n20703 & ~n20705;
  assign n20707 = ~n20695 & ~n20706;
  assign n20708 = ~n214 & ~n20707;
  assign n20709 = ~n19936 & ~n19938;
  assign n20710 = ~n20011 & n20709;
  assign n20711 = ~n34310 & ~n20710;
  assign n20712 = ~n19938 & n34310;
  assign n20713 = ~n19936 & n20712;
  assign n20714 = n34310 & n20710;
  assign n20715 = ~n20011 & n20713;
  assign n20716 = ~n20711 & ~n34403;
  assign n20717 = n214 & ~n20695;
  assign n20718 = n214 & n20707;
  assign n20719 = ~n20706 & n20717;
  assign n20720 = ~n20716 & ~n34404;
  assign n20721 = ~n20708 & ~n20720;
  assign n20722 = ~n197 & ~n20721;
  assign n20723 = n197 & ~n20708;
  assign n20724 = ~n20720 & n20723;
  assign n20725 = ~n19953 & ~n34312;
  assign n20726 = ~n19953 & ~n20011;
  assign n20727 = ~n34312 & n20726;
  assign n20728 = ~n20011 & n20725;
  assign n20729 = n19961 & ~n34405;
  assign n20730 = n19965 & n20726;
  assign n20731 = ~n19953 & n19961;
  assign n20732 = ~n34312 & n20731;
  assign n20733 = ~n20011 & n20732;
  assign n20734 = ~n19961 & ~n34405;
  assign n20735 = ~n20733 & ~n20734;
  assign n20736 = ~n20729 & ~n20730;
  assign n20737 = ~n20724 & ~n34406;
  assign n20738 = ~n20722 & ~n20737;
  assign n20739 = ~n19967 & ~n19969;
  assign n20740 = ~n20011 & n20739;
  assign n20741 = ~n34314 & ~n20740;
  assign n20742 = ~n19969 & n34314;
  assign n20743 = ~n19967 & n20742;
  assign n20744 = n34314 & n20740;
  assign n20745 = ~n20011 & n20743;
  assign n20746 = ~n20741 & ~n34407;
  assign n20747 = ~n19983 & ~n34316;
  assign n20748 = ~n34316 & ~n20011;
  assign n20749 = ~n19983 & n20748;
  assign n20750 = ~n20011 & n20747;
  assign n20751 = ~n34318 & ~n34408;
  assign n20752 = ~n20746 & n20751;
  assign n20753 = ~n20738 & n20752;
  assign n20754 = n193 & ~n20753;
  assign n20755 = ~n20722 & n20746;
  assign n20756 = n20738 & n20746;
  assign n20757 = ~n20737 & n20755;
  assign n20758 = n19983 & ~n20748;
  assign n20759 = ~n193 & ~n20747;
  assign n20760 = ~n20758 & n20759;
  assign n20761 = ~n34409 & ~n20760;
  assign n20762 = ~n20754 & n20761;
  assign n20763 = pi24  & ~n20762;
  assign n20764 = ~pi22  & ~pi23 ;
  assign n20765 = ~pi24  & n20764;
  assign n20766 = ~n20763 & ~n20765;
  assign n20767 = ~n20011 & ~n20766;
  assign n20768 = ~pi24  & ~n20762;
  assign n20769 = pi25  & ~n20768;
  assign n20770 = ~pi25  & n20768;
  assign n20771 = n20201 & ~n20762;
  assign n20772 = ~n20769 & ~n34410;
  assign n20773 = ~n34206 & ~n34343;
  assign n20774 = ~n19169 & n20773;
  assign n20775 = ~n19188 & n20774;
  assign n20776 = ~n34208 & n20775;
  assign n20777 = n19174 & n19190;
  assign n20778 = ~n19182 & n20776;
  assign n20779 = ~n20765 & ~n34411;
  assign n20780 = ~n20009 & n20779;
  assign n20781 = ~n34318 & n20780;
  assign n20782 = ~n20003 & n20781;
  assign n20783 = n20011 & n20766;
  assign n20784 = ~n20763 & n20782;
  assign n20785 = n20772 & ~n34412;
  assign n20786 = ~n20767 & ~n20785;
  assign n20787 = ~n19190 & ~n20786;
  assign n20788 = n19190 & ~n20767;
  assign n20789 = ~n20785 & n20788;
  assign n20790 = ~n20011 & ~n20760;
  assign n20791 = ~n34409 & n20790;
  assign n20792 = ~n20754 & n20791;
  assign n20793 = ~n34410 & ~n20792;
  assign n20794 = pi26  & ~n20793;
  assign n20795 = ~pi26  & ~n20792;
  assign n20796 = ~pi26  & n20793;
  assign n20797 = ~n34410 & n20795;
  assign n20798 = ~n20794 & ~n34413;
  assign n20799 = ~n20789 & ~n20798;
  assign n20800 = ~n20787 & ~n20799;
  assign n20801 = ~n18472 & ~n20800;
  assign n20802 = n18472 & ~n20787;
  assign n20803 = ~n20799 & n20802;
  assign n20804 = n18472 & n20800;
  assign n20805 = ~n34344 & ~n20219;
  assign n20806 = ~n20762 & n20805;
  assign n20807 = n20217 & ~n20806;
  assign n20808 = ~n20217 & n20805;
  assign n20809 = ~n20217 & n20806;
  assign n20810 = ~n20762 & n20808;
  assign n20811 = ~n20807 & ~n34415;
  assign n20812 = ~n34414 & ~n20811;
  assign n20813 = ~n20801 & ~n20812;
  assign n20814 = ~n17690 & ~n20813;
  assign n20815 = n17690 & ~n20801;
  assign n20816 = ~n20812 & n20815;
  assign n20817 = ~n34345 & ~n20225;
  assign n20818 = ~n20225 & ~n20762;
  assign n20819 = ~n34345 & n20818;
  assign n20820 = ~n20762 & n20817;
  assign n20821 = n20199 & ~n34416;
  assign n20822 = n20224 & n20818;
  assign n20823 = n20199 & ~n34345;
  assign n20824 = ~n20225 & n20823;
  assign n20825 = ~n20762 & n20824;
  assign n20826 = ~n20199 & ~n34416;
  assign n20827 = ~n20825 & ~n20826;
  assign n20828 = ~n20821 & ~n20822;
  assign n20829 = ~n20816 & ~n34417;
  assign n20830 = ~n20814 & ~n20829;
  assign n20831 = ~n17001 & ~n20830;
  assign n20832 = n17001 & ~n20814;
  assign n20833 = ~n20829 & n20832;
  assign n20834 = n17001 & n20830;
  assign n20835 = ~n20227 & ~n20237;
  assign n20836 = ~n20762 & n20835;
  assign n20837 = ~n20234 & ~n20836;
  assign n20838 = n20234 & ~n20237;
  assign n20839 = ~n20227 & n20838;
  assign n20840 = n20234 & n20836;
  assign n20841 = ~n20762 & n20839;
  assign n20842 = n20234 & ~n20836;
  assign n20843 = ~n20234 & n20836;
  assign n20844 = ~n20842 & ~n20843;
  assign n20845 = ~n20837 & ~n34419;
  assign n20846 = ~n34418 & n34420;
  assign n20847 = ~n20831 & ~n20846;
  assign n20848 = ~n16248 & ~n20847;
  assign n20849 = n16248 & ~n20831;
  assign n20850 = ~n20846 & n20849;
  assign n20851 = ~n34347 & ~n20243;
  assign n20852 = ~n20243 & ~n20762;
  assign n20853 = ~n34347 & n20852;
  assign n20854 = ~n20762 & n20851;
  assign n20855 = n20187 & ~n34421;
  assign n20856 = n20242 & n20852;
  assign n20857 = n20187 & ~n34347;
  assign n20858 = ~n20243 & n20857;
  assign n20859 = ~n20762 & n20858;
  assign n20860 = ~n20187 & ~n34421;
  assign n20861 = ~n20859 & ~n20860;
  assign n20862 = ~n20855 & ~n20856;
  assign n20863 = ~n20850 & ~n34422;
  assign n20864 = ~n20848 & ~n20863;
  assign n20865 = ~n15586 & ~n20864;
  assign n20866 = n15586 & ~n20848;
  assign n20867 = ~n20863 & n20866;
  assign n20868 = n15586 & n20864;
  assign n20869 = ~n20245 & ~n20259;
  assign n20870 = ~n20762 & n20869;
  assign n20871 = ~n34349 & ~n20870;
  assign n20872 = n34349 & n20870;
  assign n20873 = ~n34349 & ~n20259;
  assign n20874 = ~n20245 & n20873;
  assign n20875 = ~n20762 & n20874;
  assign n20876 = n34349 & ~n20870;
  assign n20877 = ~n20875 & ~n20876;
  assign n20878 = ~n20871 & ~n20872;
  assign n20879 = ~n34423 & ~n34424;
  assign n20880 = ~n20865 & ~n20879;
  assign n20881 = ~n14866 & ~n20880;
  assign n20882 = n14866 & ~n20865;
  assign n20883 = ~n20879 & n20882;
  assign n20884 = ~n34350 & ~n20265;
  assign n20885 = ~n20265 & ~n20762;
  assign n20886 = ~n34350 & n20885;
  assign n20887 = ~n20762 & n20884;
  assign n20888 = n20179 & ~n34425;
  assign n20889 = n20264 & n20885;
  assign n20890 = n20179 & ~n34350;
  assign n20891 = ~n20265 & n20890;
  assign n20892 = ~n20762 & n20891;
  assign n20893 = ~n20179 & ~n34425;
  assign n20894 = ~n20892 & ~n20893;
  assign n20895 = ~n20888 & ~n20889;
  assign n20896 = ~n20883 & ~n34426;
  assign n20897 = ~n20881 & ~n20896;
  assign n20898 = ~n14233 & ~n20897;
  assign n20899 = n14233 & ~n20881;
  assign n20900 = ~n20896 & n20899;
  assign n20901 = n14233 & n20897;
  assign n20902 = ~n20267 & ~n20280;
  assign n20903 = ~n20762 & n20902;
  assign n20904 = ~n34351 & n20903;
  assign n20905 = n34351 & ~n20903;
  assign n20906 = n34351 & ~n20280;
  assign n20907 = ~n20267 & n20906;
  assign n20908 = ~n20762 & n20907;
  assign n20909 = ~n34351 & ~n20903;
  assign n20910 = ~n20908 & ~n20909;
  assign n20911 = ~n20904 & ~n20905;
  assign n20912 = ~n34427 & ~n34428;
  assign n20913 = ~n20898 & ~n20912;
  assign n20914 = ~n13548 & ~n20913;
  assign n20915 = n13548 & ~n20898;
  assign n20916 = ~n20912 & n20915;
  assign n20917 = ~n34352 & ~n20286;
  assign n20918 = ~n20286 & ~n20762;
  assign n20919 = ~n34352 & n20918;
  assign n20920 = ~n20762 & n20917;
  assign n20921 = n20171 & ~n34429;
  assign n20922 = n20285 & n20918;
  assign n20923 = n20171 & ~n34352;
  assign n20924 = ~n20286 & n20923;
  assign n20925 = ~n20762 & n20924;
  assign n20926 = ~n20171 & ~n34429;
  assign n20927 = ~n20925 & ~n20926;
  assign n20928 = ~n20921 & ~n20922;
  assign n20929 = ~n20916 & ~n34430;
  assign n20930 = ~n20914 & ~n20929;
  assign n20931 = ~n12948 & ~n20930;
  assign n20932 = n12948 & ~n20914;
  assign n20933 = ~n20929 & n20932;
  assign n20934 = n12948 & n20930;
  assign n20935 = ~n20288 & ~n20301;
  assign n20936 = ~n20762 & n20935;
  assign n20937 = ~n34353 & n20936;
  assign n20938 = n34353 & ~n20936;
  assign n20939 = ~n34353 & ~n20936;
  assign n20940 = n34353 & ~n20301;
  assign n20941 = ~n20288 & n20940;
  assign n20942 = n34353 & n20936;
  assign n20943 = ~n20762 & n20941;
  assign n20944 = ~n20939 & ~n34432;
  assign n20945 = ~n20937 & ~n20938;
  assign n20946 = ~n34431 & ~n34433;
  assign n20947 = ~n20931 & ~n20946;
  assign n20948 = ~n12296 & ~n20947;
  assign n20949 = n12296 & ~n20931;
  assign n20950 = ~n20946 & n20949;
  assign n20951 = ~n34354 & ~n20307;
  assign n20952 = ~n20307 & ~n20762;
  assign n20953 = ~n34354 & n20952;
  assign n20954 = ~n20762 & n20951;
  assign n20955 = n20163 & ~n34434;
  assign n20956 = n20306 & n20952;
  assign n20957 = n20163 & ~n34354;
  assign n20958 = ~n20307 & n20957;
  assign n20959 = ~n20762 & n20958;
  assign n20960 = ~n20163 & ~n34434;
  assign n20961 = ~n20959 & ~n20960;
  assign n20962 = ~n20955 & ~n20956;
  assign n20963 = ~n20950 & ~n34435;
  assign n20964 = ~n20948 & ~n20963;
  assign n20965 = ~n11719 & ~n20964;
  assign n20966 = n11719 & ~n20948;
  assign n20967 = ~n20963 & n20966;
  assign n20968 = n11719 & n20964;
  assign n20969 = ~n20309 & ~n20323;
  assign n20970 = ~n20323 & ~n20762;
  assign n20971 = ~n20309 & n20970;
  assign n20972 = ~n20762 & n20969;
  assign n20973 = n34356 & ~n34437;
  assign n20974 = n20321 & n20970;
  assign n20975 = ~n34356 & n34437;
  assign n20976 = n34356 & ~n20323;
  assign n20977 = ~n20309 & n20976;
  assign n20978 = ~n20762 & n20977;
  assign n20979 = ~n34356 & ~n34437;
  assign n20980 = ~n20978 & ~n20979;
  assign n20981 = ~n20973 & ~n34438;
  assign n20982 = ~n34436 & ~n34439;
  assign n20983 = ~n20965 & ~n20982;
  assign n20984 = ~n11097 & ~n20983;
  assign n20985 = n11097 & ~n20965;
  assign n20986 = ~n20982 & n20985;
  assign n20987 = ~n34357 & ~n20329;
  assign n20988 = ~n20329 & ~n20762;
  assign n20989 = ~n34357 & n20988;
  assign n20990 = ~n20762 & n20987;
  assign n20991 = n20155 & ~n34440;
  assign n20992 = n20328 & n20988;
  assign n20993 = n20155 & ~n34357;
  assign n20994 = ~n20329 & n20993;
  assign n20995 = ~n20762 & n20994;
  assign n20996 = ~n20155 & ~n34440;
  assign n20997 = ~n20995 & ~n20996;
  assign n20998 = ~n20991 & ~n20992;
  assign n20999 = ~n20986 & ~n34441;
  assign n21000 = ~n20984 & ~n20999;
  assign n21001 = ~n10555 & ~n21000;
  assign n21002 = ~n20331 & ~n20347;
  assign n21003 = ~n20762 & n21002;
  assign n21004 = ~n34360 & ~n21003;
  assign n21005 = n34360 & ~n20347;
  assign n21006 = ~n20331 & n21005;
  assign n21007 = n34360 & n21003;
  assign n21008 = ~n20762 & n21006;
  assign n21009 = ~n21004 & ~n34442;
  assign n21010 = n10555 & ~n20984;
  assign n21011 = ~n20999 & n21010;
  assign n21012 = n10555 & n21000;
  assign n21013 = ~n21009 & ~n34443;
  assign n21014 = ~n21001 & ~n21013;
  assign n21015 = ~n9969 & ~n21014;
  assign n21016 = n9969 & ~n21001;
  assign n21017 = ~n21013 & n21016;
  assign n21018 = ~n34361 & ~n20353;
  assign n21019 = ~n20353 & ~n20762;
  assign n21020 = ~n34361 & n21019;
  assign n21021 = ~n20762 & n21018;
  assign n21022 = n20147 & ~n34444;
  assign n21023 = n20352 & n21019;
  assign n21024 = n20147 & ~n34361;
  assign n21025 = ~n20353 & n21024;
  assign n21026 = ~n20762 & n21025;
  assign n21027 = ~n20147 & ~n34444;
  assign n21028 = ~n21026 & ~n21027;
  assign n21029 = ~n21022 & ~n21023;
  assign n21030 = ~n21017 & ~n34445;
  assign n21031 = ~n21015 & ~n21030;
  assign n21032 = ~n9457 & ~n21031;
  assign n21033 = n9457 & ~n21015;
  assign n21034 = ~n21030 & n21033;
  assign n21035 = n9457 & n21031;
  assign n21036 = ~n20355 & ~n20358;
  assign n21037 = ~n20358 & ~n20762;
  assign n21038 = ~n20355 & n21037;
  assign n21039 = ~n20762 & n21036;
  assign n21040 = n20139 & ~n34447;
  assign n21041 = n20356 & n21037;
  assign n21042 = n20139 & ~n20358;
  assign n21043 = ~n20355 & n21042;
  assign n21044 = ~n20762 & n21043;
  assign n21045 = ~n20139 & ~n34447;
  assign n21046 = ~n21044 & ~n21045;
  assign n21047 = ~n21040 & ~n21041;
  assign n21048 = ~n34446 & ~n34448;
  assign n21049 = ~n21032 & ~n21048;
  assign n21050 = ~n8896 & ~n21049;
  assign n21051 = n8896 & ~n21032;
  assign n21052 = ~n21048 & n21051;
  assign n21053 = ~n34362 & ~n20364;
  assign n21054 = ~n20364 & ~n20762;
  assign n21055 = ~n34362 & n21054;
  assign n21056 = ~n20762 & n21053;
  assign n21057 = n20131 & ~n34449;
  assign n21058 = n20363 & n21054;
  assign n21059 = n20131 & ~n34362;
  assign n21060 = ~n20364 & n21059;
  assign n21061 = ~n20762 & n21060;
  assign n21062 = ~n20131 & ~n34449;
  assign n21063 = ~n21061 & ~n21062;
  assign n21064 = ~n21057 & ~n21058;
  assign n21065 = ~n21052 & ~n34450;
  assign n21066 = ~n21050 & ~n21065;
  assign n21067 = ~n8411 & ~n21066;
  assign n21068 = ~n20366 & ~n20381;
  assign n21069 = ~n20762 & n21068;
  assign n21070 = ~n34364 & ~n21069;
  assign n21071 = n34364 & ~n20381;
  assign n21072 = ~n20366 & n21071;
  assign n21073 = n34364 & n21069;
  assign n21074 = ~n20762 & n21072;
  assign n21075 = ~n21070 & ~n34451;
  assign n21076 = n8411 & ~n21050;
  assign n21077 = ~n21065 & n21076;
  assign n21078 = n8411 & n21066;
  assign n21079 = ~n21075 & ~n34452;
  assign n21080 = ~n21067 & ~n21079;
  assign n21081 = ~n7885 & ~n21080;
  assign n21082 = n7885 & ~n21067;
  assign n21083 = ~n21079 & n21082;
  assign n21084 = ~n34365 & ~n20387;
  assign n21085 = ~n20387 & ~n20762;
  assign n21086 = ~n34365 & n21085;
  assign n21087 = ~n20762 & n21084;
  assign n21088 = n20123 & ~n34453;
  assign n21089 = n20386 & n21085;
  assign n21090 = n20123 & ~n34365;
  assign n21091 = ~n20387 & n21090;
  assign n21092 = ~n20762 & n21091;
  assign n21093 = ~n20123 & ~n34453;
  assign n21094 = ~n21092 & ~n21093;
  assign n21095 = ~n21088 & ~n21089;
  assign n21096 = ~n21083 & ~n34454;
  assign n21097 = ~n21081 & ~n21096;
  assign n21098 = ~n7428 & ~n21097;
  assign n21099 = n7428 & ~n21081;
  assign n21100 = ~n21096 & n21099;
  assign n21101 = n7428 & n21097;
  assign n21102 = ~n20389 & ~n20392;
  assign n21103 = ~n20392 & ~n20762;
  assign n21104 = ~n20389 & n21103;
  assign n21105 = ~n20762 & n21102;
  assign n21106 = n20115 & ~n34456;
  assign n21107 = n20390 & n21103;
  assign n21108 = n20115 & ~n20392;
  assign n21109 = ~n20389 & n21108;
  assign n21110 = ~n20762 & n21109;
  assign n21111 = ~n20115 & ~n34456;
  assign n21112 = ~n21110 & ~n21111;
  assign n21113 = ~n21106 & ~n21107;
  assign n21114 = ~n34455 & ~n34457;
  assign n21115 = ~n21098 & ~n21114;
  assign n21116 = ~n6937 & ~n21115;
  assign n21117 = n6937 & ~n21098;
  assign n21118 = ~n21114 & n21117;
  assign n21119 = ~n34366 & ~n20398;
  assign n21120 = ~n20398 & ~n20762;
  assign n21121 = ~n34366 & n21120;
  assign n21122 = ~n20762 & n21119;
  assign n21123 = n20107 & ~n34458;
  assign n21124 = n20397 & n21120;
  assign n21125 = n20107 & ~n34366;
  assign n21126 = ~n20398 & n21125;
  assign n21127 = ~n20762 & n21126;
  assign n21128 = ~n20107 & ~n34458;
  assign n21129 = ~n21127 & ~n21128;
  assign n21130 = ~n21123 & ~n21124;
  assign n21131 = ~n21118 & ~n34459;
  assign n21132 = ~n21116 & ~n21131;
  assign n21133 = ~n6507 & ~n21132;
  assign n21134 = ~n20400 & ~n20415;
  assign n21135 = ~n20762 & n21134;
  assign n21136 = ~n34368 & ~n21135;
  assign n21137 = n34368 & ~n20415;
  assign n21138 = ~n20400 & n21137;
  assign n21139 = n34368 & n21135;
  assign n21140 = ~n20762 & n21138;
  assign n21141 = ~n21136 & ~n34460;
  assign n21142 = n6507 & ~n21116;
  assign n21143 = ~n21131 & n21142;
  assign n21144 = n6507 & n21132;
  assign n21145 = ~n21141 & ~n34461;
  assign n21146 = ~n21133 & ~n21145;
  assign n21147 = ~n6051 & ~n21146;
  assign n21148 = n6051 & ~n21133;
  assign n21149 = ~n21145 & n21148;
  assign n21150 = ~n34369 & ~n20421;
  assign n21151 = ~n20421 & ~n20762;
  assign n21152 = ~n34369 & n21151;
  assign n21153 = ~n20762 & n21150;
  assign n21154 = n20099 & ~n34462;
  assign n21155 = n20420 & n21151;
  assign n21156 = n20099 & ~n34369;
  assign n21157 = ~n20421 & n21156;
  assign n21158 = ~n20762 & n21157;
  assign n21159 = ~n20099 & ~n34462;
  assign n21160 = ~n21158 & ~n21159;
  assign n21161 = ~n21154 & ~n21155;
  assign n21162 = ~n21149 & ~n34463;
  assign n21163 = ~n21147 & ~n21162;
  assign n21164 = ~n5648 & ~n21163;
  assign n21165 = n5648 & ~n21147;
  assign n21166 = ~n21162 & n21165;
  assign n21167 = n5648 & n21163;
  assign n21168 = ~n20423 & ~n20426;
  assign n21169 = ~n20426 & ~n20762;
  assign n21170 = ~n20423 & n21169;
  assign n21171 = ~n20762 & n21168;
  assign n21172 = n20091 & ~n34465;
  assign n21173 = n20424 & n21169;
  assign n21174 = n20091 & ~n20426;
  assign n21175 = ~n20423 & n21174;
  assign n21176 = ~n20762 & n21175;
  assign n21177 = ~n20091 & ~n34465;
  assign n21178 = ~n21176 & ~n21177;
  assign n21179 = ~n21172 & ~n21173;
  assign n21180 = ~n34464 & ~n34466;
  assign n21181 = ~n21164 & ~n21180;
  assign n21182 = ~n5223 & ~n21181;
  assign n21183 = n5223 & ~n21164;
  assign n21184 = ~n21180 & n21183;
  assign n21185 = ~n34370 & ~n20432;
  assign n21186 = ~n20432 & ~n20762;
  assign n21187 = ~n34370 & n21186;
  assign n21188 = ~n20762 & n21185;
  assign n21189 = n20083 & ~n34467;
  assign n21190 = n20431 & n21186;
  assign n21191 = n20083 & ~n34370;
  assign n21192 = ~n20432 & n21191;
  assign n21193 = ~n20762 & n21192;
  assign n21194 = ~n20083 & ~n34467;
  assign n21195 = ~n21193 & ~n21194;
  assign n21196 = ~n21189 & ~n21190;
  assign n21197 = ~n21184 & ~n34468;
  assign n21198 = ~n21182 & ~n21197;
  assign n21199 = ~n4851 & ~n21198;
  assign n21200 = ~n20434 & ~n20449;
  assign n21201 = ~n20762 & n21200;
  assign n21202 = ~n34372 & ~n21201;
  assign n21203 = n34372 & ~n20449;
  assign n21204 = ~n20434 & n21203;
  assign n21205 = n34372 & n21201;
  assign n21206 = ~n20762 & n21204;
  assign n21207 = ~n21202 & ~n34469;
  assign n21208 = n4851 & ~n21182;
  assign n21209 = ~n21197 & n21208;
  assign n21210 = n4851 & n21198;
  assign n21211 = ~n21207 & ~n34470;
  assign n21212 = ~n21199 & ~n21211;
  assign n21213 = ~n4461 & ~n21212;
  assign n21214 = n4461 & ~n21199;
  assign n21215 = ~n21211 & n21214;
  assign n21216 = ~n34373 & ~n20455;
  assign n21217 = ~n20455 & ~n20762;
  assign n21218 = ~n34373 & n21217;
  assign n21219 = ~n20762 & n21216;
  assign n21220 = n20075 & ~n34471;
  assign n21221 = n20454 & n21217;
  assign n21222 = n20075 & ~n34373;
  assign n21223 = ~n20455 & n21222;
  assign n21224 = ~n20762 & n21223;
  assign n21225 = ~n20075 & ~n34471;
  assign n21226 = ~n21224 & ~n21225;
  assign n21227 = ~n21220 & ~n21221;
  assign n21228 = ~n21215 & ~n34472;
  assign n21229 = ~n21213 & ~n21228;
  assign n21230 = ~n4115 & ~n21229;
  assign n21231 = n4115 & ~n21213;
  assign n21232 = ~n21228 & n21231;
  assign n21233 = n4115 & n21229;
  assign n21234 = ~n20457 & ~n20460;
  assign n21235 = ~n20460 & ~n20762;
  assign n21236 = ~n20457 & n21235;
  assign n21237 = ~n20762 & n21234;
  assign n21238 = n20067 & ~n34474;
  assign n21239 = n20458 & n21235;
  assign n21240 = n20067 & ~n20460;
  assign n21241 = ~n20457 & n21240;
  assign n21242 = ~n20762 & n21241;
  assign n21243 = ~n20067 & ~n34474;
  assign n21244 = ~n21242 & ~n21243;
  assign n21245 = ~n21238 & ~n21239;
  assign n21246 = ~n34473 & ~n34475;
  assign n21247 = ~n21230 & ~n21246;
  assign n21248 = ~n3754 & ~n21247;
  assign n21249 = n3754 & ~n21230;
  assign n21250 = ~n21246 & n21249;
  assign n21251 = ~n34374 & ~n20466;
  assign n21252 = ~n20466 & ~n20762;
  assign n21253 = ~n34374 & n21252;
  assign n21254 = ~n20762 & n21251;
  assign n21255 = n20059 & ~n34476;
  assign n21256 = n20465 & n21252;
  assign n21257 = n20059 & ~n34374;
  assign n21258 = ~n20466 & n21257;
  assign n21259 = ~n20762 & n21258;
  assign n21260 = ~n20059 & ~n34476;
  assign n21261 = ~n21259 & ~n21260;
  assign n21262 = ~n21255 & ~n21256;
  assign n21263 = ~n21250 & ~n34477;
  assign n21264 = ~n21248 & ~n21263;
  assign n21265 = ~n3444 & ~n21264;
  assign n21266 = ~n20468 & ~n20483;
  assign n21267 = ~n20762 & n21266;
  assign n21268 = ~n34376 & ~n21267;
  assign n21269 = n34376 & ~n20483;
  assign n21270 = ~n20468 & n21269;
  assign n21271 = n34376 & n21267;
  assign n21272 = ~n20762 & n21270;
  assign n21273 = ~n21268 & ~n34478;
  assign n21274 = n3444 & ~n21248;
  assign n21275 = ~n21263 & n21274;
  assign n21276 = n3444 & n21264;
  assign n21277 = ~n21273 & ~n34479;
  assign n21278 = ~n21265 & ~n21277;
  assign n21279 = ~n3116 & ~n21278;
  assign n21280 = n3116 & ~n21265;
  assign n21281 = ~n21277 & n21280;
  assign n21282 = ~n34377 & ~n20489;
  assign n21283 = ~n20489 & ~n20762;
  assign n21284 = ~n34377 & n21283;
  assign n21285 = ~n20762 & n21282;
  assign n21286 = n20051 & ~n34480;
  assign n21287 = n20488 & n21283;
  assign n21288 = n20051 & ~n34377;
  assign n21289 = ~n20489 & n21288;
  assign n21290 = ~n20762 & n21289;
  assign n21291 = ~n20051 & ~n34480;
  assign n21292 = ~n21290 & ~n21291;
  assign n21293 = ~n21286 & ~n21287;
  assign n21294 = ~n21281 & ~n34481;
  assign n21295 = ~n21279 & ~n21294;
  assign n21296 = ~n2833 & ~n21295;
  assign n21297 = n2833 & ~n21279;
  assign n21298 = ~n21294 & n21297;
  assign n21299 = n2833 & n21295;
  assign n21300 = ~n20491 & ~n20494;
  assign n21301 = ~n20494 & ~n20762;
  assign n21302 = ~n20491 & n21301;
  assign n21303 = ~n20762 & n21300;
  assign n21304 = n20043 & ~n34483;
  assign n21305 = n20492 & n21301;
  assign n21306 = n20043 & ~n20494;
  assign n21307 = ~n20491 & n21306;
  assign n21308 = ~n20762 & n21307;
  assign n21309 = ~n20043 & ~n34483;
  assign n21310 = ~n21308 & ~n21309;
  assign n21311 = ~n21304 & ~n21305;
  assign n21312 = ~n34482 & ~n34484;
  assign n21313 = ~n21296 & ~n21312;
  assign n21314 = ~n2536 & ~n21313;
  assign n21315 = n2536 & ~n21296;
  assign n21316 = ~n21312 & n21315;
  assign n21317 = ~n34378 & ~n20500;
  assign n21318 = ~n20500 & ~n20762;
  assign n21319 = ~n34378 & n21318;
  assign n21320 = ~n20762 & n21317;
  assign n21321 = n20035 & ~n34485;
  assign n21322 = n20499 & n21318;
  assign n21323 = n20035 & ~n34378;
  assign n21324 = ~n20500 & n21323;
  assign n21325 = ~n20762 & n21324;
  assign n21326 = ~n20035 & ~n34485;
  assign n21327 = ~n21325 & ~n21326;
  assign n21328 = ~n21321 & ~n21322;
  assign n21329 = ~n21316 & ~n34486;
  assign n21330 = ~n21314 & ~n21329;
  assign n21331 = ~n2283 & ~n21330;
  assign n21332 = ~n20502 & ~n20517;
  assign n21333 = ~n20762 & n21332;
  assign n21334 = ~n34380 & ~n21333;
  assign n21335 = n34380 & ~n20517;
  assign n21336 = ~n20502 & n21335;
  assign n21337 = n34380 & n21333;
  assign n21338 = ~n20762 & n21336;
  assign n21339 = ~n21334 & ~n34487;
  assign n21340 = n2283 & ~n21314;
  assign n21341 = ~n21329 & n21340;
  assign n21342 = n2283 & n21330;
  assign n21343 = ~n21339 & ~n34488;
  assign n21344 = ~n21331 & ~n21343;
  assign n21345 = ~n2021 & ~n21344;
  assign n21346 = n2021 & ~n21331;
  assign n21347 = ~n21343 & n21346;
  assign n21348 = ~n34381 & ~n20523;
  assign n21349 = ~n20523 & ~n20762;
  assign n21350 = ~n34381 & n21349;
  assign n21351 = ~n20762 & n21348;
  assign n21352 = n20027 & ~n34489;
  assign n21353 = n20522 & n21349;
  assign n21354 = n20027 & ~n34381;
  assign n21355 = ~n20523 & n21354;
  assign n21356 = ~n20762 & n21355;
  assign n21357 = ~n20027 & ~n34489;
  assign n21358 = ~n21356 & ~n21357;
  assign n21359 = ~n21352 & ~n21353;
  assign n21360 = ~n21347 & ~n34490;
  assign n21361 = ~n21345 & ~n21360;
  assign n21362 = ~n1796 & ~n21361;
  assign n21363 = n1796 & ~n21345;
  assign n21364 = ~n21360 & n21363;
  assign n21365 = n1796 & n21361;
  assign n21366 = ~n20525 & ~n20528;
  assign n21367 = ~n20528 & ~n20762;
  assign n21368 = ~n20525 & n21367;
  assign n21369 = ~n20762 & n21366;
  assign n21370 = n20019 & ~n34492;
  assign n21371 = n20526 & n21367;
  assign n21372 = n20019 & ~n20528;
  assign n21373 = ~n20525 & n21372;
  assign n21374 = ~n20762 & n21373;
  assign n21375 = ~n20019 & ~n34492;
  assign n21376 = ~n21374 & ~n21375;
  assign n21377 = ~n21370 & ~n21371;
  assign n21378 = ~n34491 & ~n34493;
  assign n21379 = ~n21362 & ~n21378;
  assign n21380 = ~n1567 & ~n21379;
  assign n21381 = n1567 & ~n21362;
  assign n21382 = ~n21378 & n21381;
  assign n21383 = ~n34382 & ~n20544;
  assign n21384 = ~n20762 & n21383;
  assign n21385 = ~n34383 & n21384;
  assign n21386 = n34383 & ~n21384;
  assign n21387 = ~n34382 & n34383;
  assign n21388 = ~n20544 & n21387;
  assign n21389 = ~n20762 & n21388;
  assign n21390 = ~n34383 & ~n21384;
  assign n21391 = ~n21389 & ~n21390;
  assign n21392 = ~n21385 & ~n21386;
  assign n21393 = ~n21382 & ~n34494;
  assign n21394 = ~n21380 & ~n21393;
  assign n21395 = ~n1374 & ~n21394;
  assign n21396 = ~n20546 & ~n20558;
  assign n21397 = ~n20762 & n21396;
  assign n21398 = ~n34384 & ~n21397;
  assign n21399 = ~n20546 & n34384;
  assign n21400 = ~n20558 & n21399;
  assign n21401 = n34384 & n21397;
  assign n21402 = ~n20762 & n21400;
  assign n21403 = ~n21398 & ~n34495;
  assign n21404 = n1374 & ~n21380;
  assign n21405 = ~n21393 & n21404;
  assign n21406 = n1374 & n21394;
  assign n21407 = ~n21403 & ~n34496;
  assign n21408 = ~n21395 & ~n21407;
  assign n21409 = ~n1179 & ~n21408;
  assign n21410 = n1179 & ~n21395;
  assign n21411 = ~n21407 & n21410;
  assign n21412 = ~n20561 & ~n34386;
  assign n21413 = ~n20561 & ~n20762;
  assign n21414 = ~n34386 & n21413;
  assign n21415 = ~n20762 & n21412;
  assign n21416 = n20569 & ~n34497;
  assign n21417 = n20573 & n21413;
  assign n21418 = n20569 & ~n34386;
  assign n21419 = ~n20561 & n21418;
  assign n21420 = ~n20762 & n21419;
  assign n21421 = ~n20569 & ~n34497;
  assign n21422 = ~n21420 & ~n21421;
  assign n21423 = ~n21416 & ~n21417;
  assign n21424 = ~n21411 & ~n34498;
  assign n21425 = ~n21409 & ~n21424;
  assign n21426 = ~n1016 & ~n21425;
  assign n21427 = ~n20575 & ~n20577;
  assign n21428 = ~n20762 & n21427;
  assign n21429 = ~n34388 & ~n21428;
  assign n21430 = ~n20575 & n34388;
  assign n21431 = ~n20577 & n21430;
  assign n21432 = n34388 & n21428;
  assign n21433 = ~n20762 & n21431;
  assign n21434 = ~n21429 & ~n34499;
  assign n21435 = n1016 & ~n21409;
  assign n21436 = ~n21424 & n21435;
  assign n21437 = n1016 & n21425;
  assign n21438 = ~n21434 & ~n34500;
  assign n21439 = ~n21426 & ~n21438;
  assign n21440 = ~n855 & ~n21439;
  assign n21441 = n855 & ~n21426;
  assign n21442 = ~n21438 & n21441;
  assign n21443 = ~n20592 & ~n34390;
  assign n21444 = ~n20592 & ~n20762;
  assign n21445 = ~n34390 & n21444;
  assign n21446 = ~n20762 & n21443;
  assign n21447 = n20600 & ~n34501;
  assign n21448 = n20604 & n21444;
  assign n21449 = n20600 & ~n34390;
  assign n21450 = ~n20592 & n21449;
  assign n21451 = ~n20762 & n21450;
  assign n21452 = ~n20600 & ~n34501;
  assign n21453 = ~n21451 & ~n21452;
  assign n21454 = ~n21447 & ~n21448;
  assign n21455 = ~n21442 & ~n34502;
  assign n21456 = ~n21440 & ~n21455;
  assign n21457 = ~n720 & ~n21456;
  assign n21458 = ~n20606 & ~n20608;
  assign n21459 = ~n20762 & n21458;
  assign n21460 = ~n34392 & ~n21459;
  assign n21461 = ~n20606 & n34392;
  assign n21462 = ~n20608 & n21461;
  assign n21463 = n34392 & n21459;
  assign n21464 = ~n20762 & n21462;
  assign n21465 = ~n21460 & ~n34503;
  assign n21466 = n720 & ~n21440;
  assign n21467 = ~n21455 & n21466;
  assign n21468 = n720 & n21456;
  assign n21469 = ~n21465 & ~n34504;
  assign n21470 = ~n21457 & ~n21469;
  assign n21471 = ~n592 & ~n21470;
  assign n21472 = n592 & ~n21457;
  assign n21473 = ~n21469 & n21472;
  assign n21474 = ~n20623 & ~n34394;
  assign n21475 = ~n20623 & ~n20762;
  assign n21476 = ~n34394 & n21475;
  assign n21477 = ~n20762 & n21474;
  assign n21478 = n20631 & ~n34505;
  assign n21479 = n20635 & n21475;
  assign n21480 = n20631 & ~n34394;
  assign n21481 = ~n20623 & n21480;
  assign n21482 = ~n20762 & n21481;
  assign n21483 = ~n20631 & ~n34505;
  assign n21484 = ~n21482 & ~n21483;
  assign n21485 = ~n21478 & ~n21479;
  assign n21486 = ~n21473 & ~n34506;
  assign n21487 = ~n21471 & ~n21486;
  assign n21488 = ~n487 & ~n21487;
  assign n21489 = n487 & ~n21471;
  assign n21490 = ~n21486 & n21489;
  assign n21491 = n487 & n21487;
  assign n21492 = ~n20637 & ~n20647;
  assign n21493 = ~n20637 & ~n20762;
  assign n21494 = ~n20647 & n21493;
  assign n21495 = ~n20762 & n21492;
  assign n21496 = n20645 & ~n34508;
  assign n21497 = n20648 & n21493;
  assign n21498 = ~n20637 & n20645;
  assign n21499 = ~n20647 & n21498;
  assign n21500 = ~n20762 & n21499;
  assign n21501 = ~n20645 & ~n34508;
  assign n21502 = ~n21500 & ~n21501;
  assign n21503 = ~n21496 & ~n21497;
  assign n21504 = ~n34507 & ~n34509;
  assign n21505 = ~n21488 & ~n21504;
  assign n21506 = ~n393 & ~n21505;
  assign n21507 = n393 & ~n21488;
  assign n21508 = ~n21504 & n21507;
  assign n21509 = ~n20650 & ~n34397;
  assign n21510 = ~n20650 & ~n20762;
  assign n21511 = ~n34397 & n21510;
  assign n21512 = ~n20762 & n21509;
  assign n21513 = n20658 & ~n34510;
  assign n21514 = n20662 & n21510;
  assign n21515 = n20658 & ~n34397;
  assign n21516 = ~n20650 & n21515;
  assign n21517 = ~n20762 & n21516;
  assign n21518 = ~n20658 & ~n34510;
  assign n21519 = ~n21517 & ~n21518;
  assign n21520 = ~n21513 & ~n21514;
  assign n21521 = ~n21508 & ~n34511;
  assign n21522 = ~n21506 & ~n21521;
  assign n21523 = ~n321 & ~n21522;
  assign n21524 = ~n20664 & ~n20666;
  assign n21525 = ~n20762 & n21524;
  assign n21526 = ~n34399 & ~n21525;
  assign n21527 = ~n20664 & n34399;
  assign n21528 = ~n20666 & n21527;
  assign n21529 = n34399 & n21525;
  assign n21530 = ~n20762 & n21528;
  assign n21531 = ~n21526 & ~n34512;
  assign n21532 = n321 & ~n21506;
  assign n21533 = ~n21521 & n21532;
  assign n21534 = n321 & n21522;
  assign n21535 = ~n21531 & ~n34513;
  assign n21536 = ~n21523 & ~n21535;
  assign n21537 = ~n263 & ~n21536;
  assign n21538 = n263 & ~n21523;
  assign n21539 = ~n21535 & n21538;
  assign n21540 = ~n20681 & ~n34401;
  assign n21541 = ~n20681 & ~n20762;
  assign n21542 = ~n34401 & n21541;
  assign n21543 = ~n20762 & n21540;
  assign n21544 = n20689 & ~n34514;
  assign n21545 = n20693 & n21541;
  assign n21546 = n20689 & ~n34401;
  assign n21547 = ~n20681 & n21546;
  assign n21548 = ~n20762 & n21547;
  assign n21549 = ~n20689 & ~n34514;
  assign n21550 = ~n21548 & ~n21549;
  assign n21551 = ~n21544 & ~n21545;
  assign n21552 = ~n21539 & ~n34515;
  assign n21553 = ~n21537 & ~n21552;
  assign n21554 = ~n214 & ~n21553;
  assign n21555 = n214 & ~n21537;
  assign n21556 = ~n21552 & n21555;
  assign n21557 = n214 & n21553;
  assign n21558 = ~n20695 & ~n20705;
  assign n21559 = ~n20695 & ~n20762;
  assign n21560 = ~n20705 & n21559;
  assign n21561 = ~n20762 & n21558;
  assign n21562 = n20703 & ~n34517;
  assign n21563 = n20706 & n21559;
  assign n21564 = ~n20695 & n20703;
  assign n21565 = ~n20705 & n21564;
  assign n21566 = ~n20762 & n21565;
  assign n21567 = ~n20703 & ~n34517;
  assign n21568 = ~n21566 & ~n21567;
  assign n21569 = ~n21562 & ~n21563;
  assign n21570 = ~n34516 & ~n34518;
  assign n21571 = ~n21554 & ~n21570;
  assign n21572 = ~n197 & ~n21571;
  assign n21573 = n197 & ~n21554;
  assign n21574 = ~n21570 & n21573;
  assign n21575 = ~n20708 & ~n34404;
  assign n21576 = ~n20708 & ~n20762;
  assign n21577 = ~n34404 & n21576;
  assign n21578 = ~n20762 & n21575;
  assign n21579 = n20716 & ~n34519;
  assign n21580 = n20720 & n21576;
  assign n21581 = n20716 & ~n34404;
  assign n21582 = ~n20708 & n21581;
  assign n21583 = ~n20762 & n21582;
  assign n21584 = ~n20716 & ~n34519;
  assign n21585 = ~n21583 & ~n21584;
  assign n21586 = ~n21579 & ~n21580;
  assign n21587 = ~n21574 & ~n34520;
  assign n21588 = ~n21572 & ~n21587;
  assign n21589 = ~n20722 & ~n20724;
  assign n21590 = ~n20762 & n21589;
  assign n21591 = ~n34406 & ~n21590;
  assign n21592 = ~n20722 & n34406;
  assign n21593 = ~n20724 & n21592;
  assign n21594 = n34406 & n21590;
  assign n21595 = ~n20762 & n21593;
  assign n21596 = ~n21591 & ~n34521;
  assign n21597 = ~n20738 & ~n20746;
  assign n21598 = ~n20746 & ~n20762;
  assign n21599 = ~n20738 & n21598;
  assign n21600 = ~n20762 & n21597;
  assign n21601 = ~n34409 & ~n34522;
  assign n21602 = ~n21596 & n21601;
  assign n21603 = ~n21588 & n21602;
  assign n21604 = n193 & ~n21603;
  assign n21605 = ~n21572 & n21596;
  assign n21606 = ~n21587 & n21605;
  assign n21607 = n21588 & n21596;
  assign n21608 = n20738 & ~n21598;
  assign n21609 = ~n193 & ~n21597;
  assign n21610 = ~n21608 & n21609;
  assign n21611 = ~n34523 & ~n21610;
  assign n21612 = ~n21604 & n21611;
  assign n21613 = ~n21380 & ~n21382;
  assign n21614 = ~n21612 & n21613;
  assign n21615 = ~n34494 & ~n21614;
  assign n21616 = ~n21382 & n34494;
  assign n21617 = ~n21380 & n21616;
  assign n21618 = n34494 & n21614;
  assign n21619 = ~n21612 & n21617;
  assign n21620 = ~n21615 & ~n34524;
  assign n21621 = ~n21362 & ~n34491;
  assign n21622 = ~n21612 & n21621;
  assign n21623 = ~n34493 & ~n21622;
  assign n21624 = ~n21362 & n34493;
  assign n21625 = ~n34491 & n21624;
  assign n21626 = n34493 & n21622;
  assign n21627 = ~n21612 & n21625;
  assign n21628 = ~n21623 & ~n34525;
  assign n21629 = ~n21345 & ~n21347;
  assign n21630 = ~n21612 & n21629;
  assign n21631 = ~n34490 & ~n21630;
  assign n21632 = ~n21347 & n34490;
  assign n21633 = ~n21345 & n21632;
  assign n21634 = n34490 & n21630;
  assign n21635 = ~n21612 & n21633;
  assign n21636 = ~n21631 & ~n34526;
  assign n21637 = ~n21314 & ~n21316;
  assign n21638 = ~n21612 & n21637;
  assign n21639 = ~n34486 & ~n21638;
  assign n21640 = ~n21316 & n34486;
  assign n21641 = ~n21314 & n21640;
  assign n21642 = n34486 & n21638;
  assign n21643 = ~n21612 & n21641;
  assign n21644 = ~n21639 & ~n34527;
  assign n21645 = ~n21296 & ~n34482;
  assign n21646 = ~n21612 & n21645;
  assign n21647 = ~n34484 & ~n21646;
  assign n21648 = ~n21296 & n34484;
  assign n21649 = ~n34482 & n21648;
  assign n21650 = n34484 & n21646;
  assign n21651 = ~n21612 & n21649;
  assign n21652 = ~n21647 & ~n34528;
  assign n21653 = ~n21279 & ~n21281;
  assign n21654 = ~n21612 & n21653;
  assign n21655 = ~n34481 & ~n21654;
  assign n21656 = ~n21281 & n34481;
  assign n21657 = ~n21279 & n21656;
  assign n21658 = n34481 & n21654;
  assign n21659 = ~n21612 & n21657;
  assign n21660 = ~n21655 & ~n34529;
  assign n21661 = ~n21248 & ~n21250;
  assign n21662 = ~n21612 & n21661;
  assign n21663 = ~n34477 & ~n21662;
  assign n21664 = ~n21250 & n34477;
  assign n21665 = ~n21248 & n21664;
  assign n21666 = n34477 & n21662;
  assign n21667 = ~n21612 & n21665;
  assign n21668 = ~n21663 & ~n34530;
  assign n21669 = ~n21230 & ~n34473;
  assign n21670 = ~n21612 & n21669;
  assign n21671 = ~n34475 & ~n21670;
  assign n21672 = ~n21230 & n34475;
  assign n21673 = ~n34473 & n21672;
  assign n21674 = n34475 & n21670;
  assign n21675 = ~n21612 & n21673;
  assign n21676 = ~n21671 & ~n34531;
  assign n21677 = ~n21213 & ~n21215;
  assign n21678 = ~n21612 & n21677;
  assign n21679 = ~n34472 & ~n21678;
  assign n21680 = ~n21215 & n34472;
  assign n21681 = ~n21213 & n21680;
  assign n21682 = n34472 & n21678;
  assign n21683 = ~n21612 & n21681;
  assign n21684 = ~n21679 & ~n34532;
  assign n21685 = ~n21182 & ~n21184;
  assign n21686 = ~n21612 & n21685;
  assign n21687 = ~n34468 & ~n21686;
  assign n21688 = ~n21184 & n34468;
  assign n21689 = ~n21182 & n21688;
  assign n21690 = n34468 & n21686;
  assign n21691 = ~n21612 & n21689;
  assign n21692 = ~n21687 & ~n34533;
  assign n21693 = ~n21164 & ~n34464;
  assign n21694 = ~n21612 & n21693;
  assign n21695 = ~n34466 & ~n21694;
  assign n21696 = ~n21164 & n34466;
  assign n21697 = ~n34464 & n21696;
  assign n21698 = n34466 & n21694;
  assign n21699 = ~n21612 & n21697;
  assign n21700 = ~n21695 & ~n34534;
  assign n21701 = ~n21147 & ~n21149;
  assign n21702 = ~n21612 & n21701;
  assign n21703 = ~n34463 & ~n21702;
  assign n21704 = ~n21149 & n34463;
  assign n21705 = ~n21147 & n21704;
  assign n21706 = n34463 & n21702;
  assign n21707 = ~n21612 & n21705;
  assign n21708 = ~n21703 & ~n34535;
  assign n21709 = ~n21116 & ~n21118;
  assign n21710 = ~n21612 & n21709;
  assign n21711 = ~n34459 & ~n21710;
  assign n21712 = ~n21118 & n34459;
  assign n21713 = ~n21116 & n21712;
  assign n21714 = n34459 & n21710;
  assign n21715 = ~n21612 & n21713;
  assign n21716 = ~n21711 & ~n34536;
  assign n21717 = ~n21098 & ~n34455;
  assign n21718 = ~n21612 & n21717;
  assign n21719 = ~n34457 & ~n21718;
  assign n21720 = ~n21098 & n34457;
  assign n21721 = ~n34455 & n21720;
  assign n21722 = n34457 & n21718;
  assign n21723 = ~n21612 & n21721;
  assign n21724 = ~n21719 & ~n34537;
  assign n21725 = ~n21081 & ~n21083;
  assign n21726 = ~n21612 & n21725;
  assign n21727 = ~n34454 & ~n21726;
  assign n21728 = ~n21083 & n34454;
  assign n21729 = ~n21081 & n21728;
  assign n21730 = n34454 & n21726;
  assign n21731 = ~n21612 & n21729;
  assign n21732 = ~n21727 & ~n34538;
  assign n21733 = ~n21050 & ~n21052;
  assign n21734 = ~n21612 & n21733;
  assign n21735 = ~n34450 & ~n21734;
  assign n21736 = ~n21052 & n34450;
  assign n21737 = ~n21050 & n21736;
  assign n21738 = n34450 & n21734;
  assign n21739 = ~n21612 & n21737;
  assign n21740 = ~n21735 & ~n34539;
  assign n21741 = ~n21032 & ~n34446;
  assign n21742 = ~n21612 & n21741;
  assign n21743 = ~n34448 & ~n21742;
  assign n21744 = ~n21032 & n34448;
  assign n21745 = ~n34446 & n21744;
  assign n21746 = n34448 & n21742;
  assign n21747 = ~n21612 & n21745;
  assign n21748 = ~n21743 & ~n34540;
  assign n21749 = ~n21015 & ~n21017;
  assign n21750 = ~n21612 & n21749;
  assign n21751 = ~n34445 & ~n21750;
  assign n21752 = ~n21017 & n34445;
  assign n21753 = ~n21015 & n21752;
  assign n21754 = n34445 & n21750;
  assign n21755 = ~n21612 & n21753;
  assign n21756 = ~n21751 & ~n34541;
  assign n21757 = ~n20984 & ~n20986;
  assign n21758 = ~n21612 & n21757;
  assign n21759 = ~n34441 & ~n21758;
  assign n21760 = ~n20986 & n34441;
  assign n21761 = ~n20984 & n21760;
  assign n21762 = n34441 & n21758;
  assign n21763 = ~n21612 & n21761;
  assign n21764 = ~n21759 & ~n34542;
  assign n21765 = ~n20965 & ~n34436;
  assign n21766 = ~n21612 & n21765;
  assign n21767 = ~n34439 & ~n21766;
  assign n21768 = ~n20965 & n34439;
  assign n21769 = ~n34436 & n21768;
  assign n21770 = n34439 & n21766;
  assign n21771 = ~n21612 & n21769;
  assign n21772 = ~n21767 & ~n34543;
  assign n21773 = ~n20948 & ~n20950;
  assign n21774 = ~n21612 & n21773;
  assign n21775 = ~n34435 & ~n21774;
  assign n21776 = ~n20950 & n34435;
  assign n21777 = ~n20948 & n21776;
  assign n21778 = n34435 & n21774;
  assign n21779 = ~n21612 & n21777;
  assign n21780 = ~n21775 & ~n34544;
  assign n21781 = ~n20914 & ~n20916;
  assign n21782 = ~n21612 & n21781;
  assign n21783 = ~n34430 & ~n21782;
  assign n21784 = ~n20916 & n34430;
  assign n21785 = ~n20914 & n21784;
  assign n21786 = n34430 & n21782;
  assign n21787 = ~n21612 & n21785;
  assign n21788 = ~n21783 & ~n34545;
  assign n21789 = ~n20881 & ~n20883;
  assign n21790 = ~n21612 & n21789;
  assign n21791 = ~n34426 & ~n21790;
  assign n21792 = ~n20883 & n34426;
  assign n21793 = ~n20881 & n21792;
  assign n21794 = n34426 & n21790;
  assign n21795 = ~n21612 & n21793;
  assign n21796 = ~n21791 & ~n34546;
  assign n21797 = ~n20848 & ~n20850;
  assign n21798 = ~n21612 & n21797;
  assign n21799 = ~n34422 & ~n21798;
  assign n21800 = ~n20850 & n34422;
  assign n21801 = ~n20848 & n21800;
  assign n21802 = n34422 & n21798;
  assign n21803 = ~n21612 & n21801;
  assign n21804 = ~n21799 & ~n34547;
  assign n21805 = ~n20814 & ~n20816;
  assign n21806 = ~n21612 & n21805;
  assign n21807 = ~n34417 & ~n21806;
  assign n21808 = ~n20816 & n34417;
  assign n21809 = ~n20814 & n21808;
  assign n21810 = n34417 & n21806;
  assign n21811 = ~n21612 & n21809;
  assign n21812 = ~n21807 & ~n34548;
  assign n21813 = ~n20787 & ~n20789;
  assign n21814 = ~n21612 & n21813;
  assign n21815 = ~n20798 & ~n21814;
  assign n21816 = ~n20789 & n20798;
  assign n21817 = ~n20787 & n21816;
  assign n21818 = n20798 & n21814;
  assign n21819 = ~n21612 & n21817;
  assign n21820 = ~n21815 & ~n34549;
  assign n21821 = ~pi22  & ~n21612;
  assign n21822 = ~pi23  & n21821;
  assign n21823 = n20764 & ~n21612;
  assign n21824 = ~n20762 & ~n21610;
  assign n21825 = ~n34523 & n21824;
  assign n21826 = ~n21604 & n21825;
  assign n21827 = ~n34550 & ~n21826;
  assign n21828 = pi24  & ~n21827;
  assign n21829 = ~pi24  & ~n21826;
  assign n21830 = ~pi24  & n21827;
  assign n21831 = ~n34550 & n21829;
  assign n21832 = ~n21828 & ~n34551;
  assign n21833 = pi22  & ~n21612;
  assign n21834 = ~pi20  & ~pi21 ;
  assign n21835 = ~pi22  & n21834;
  assign n21836 = ~n19992 & ~n34411;
  assign n21837 = ~n19993 & n21836;
  assign n21838 = ~n20009 & n21837;
  assign n21839 = ~n34318 & n21838;
  assign n21840 = n34316 & n20011;
  assign n21841 = ~n20003 & n21839;
  assign n21842 = ~n21835 & ~n34552;
  assign n21843 = ~n20760 & n21842;
  assign n21844 = ~n34409 & n21843;
  assign n21845 = ~n20754 & n21844;
  assign n21846 = ~n21833 & ~n21835;
  assign n21847 = n20762 & n21846;
  assign n21848 = ~n21833 & n21845;
  assign n21849 = pi23  & ~n21821;
  assign n21850 = ~n34550 & ~n21849;
  assign n21851 = ~n34553 & n21850;
  assign n21852 = ~n20762 & ~n21846;
  assign n21853 = n20011 & ~n21852;
  assign n21854 = ~n21851 & ~n21852;
  assign n21855 = n20011 & n21854;
  assign n21856 = ~n21851 & n21853;
  assign n21857 = ~n21832 & ~n34554;
  assign n21858 = ~n20011 & ~n21854;
  assign n21859 = n19190 & ~n21858;
  assign n21860 = ~n21857 & n21859;
  assign n21861 = ~n20767 & ~n34412;
  assign n21862 = ~n21612 & n21861;
  assign n21863 = n20772 & ~n21862;
  assign n21864 = ~n20772 & n21861;
  assign n21865 = ~n20772 & n21862;
  assign n21866 = ~n21612 & n21864;
  assign n21867 = ~n21863 & ~n34555;
  assign n21868 = ~n21860 & ~n21867;
  assign n21869 = ~n21857 & ~n21858;
  assign n21870 = ~n19190 & ~n21869;
  assign n21871 = n18472 & ~n21870;
  assign n21872 = ~n21868 & ~n21870;
  assign n21873 = n18472 & n21872;
  assign n21874 = ~n21868 & n21871;
  assign n21875 = ~n21820 & ~n34556;
  assign n21876 = ~n18472 & ~n21872;
  assign n21877 = n17690 & ~n21876;
  assign n21878 = ~n21875 & n21877;
  assign n21879 = ~n20801 & ~n34414;
  assign n21880 = ~n21612 & n21879;
  assign n21881 = ~n20811 & ~n21880;
  assign n21882 = ~n20801 & n20811;
  assign n21883 = ~n34414 & n21882;
  assign n21884 = n20811 & n21880;
  assign n21885 = ~n21612 & n21883;
  assign n21886 = n20811 & ~n21880;
  assign n21887 = ~n20811 & n21880;
  assign n21888 = ~n21886 & ~n21887;
  assign n21889 = ~n21881 & ~n34557;
  assign n21890 = ~n21878 & n34558;
  assign n21891 = ~n21875 & ~n21876;
  assign n21892 = ~n17690 & ~n21891;
  assign n21893 = n17001 & ~n21892;
  assign n21894 = ~n21890 & ~n21892;
  assign n21895 = n17001 & n21894;
  assign n21896 = ~n21890 & n21893;
  assign n21897 = ~n21812 & ~n34559;
  assign n21898 = ~n17001 & ~n21894;
  assign n21899 = n16248 & ~n21898;
  assign n21900 = ~n21897 & n21899;
  assign n21901 = ~n20831 & ~n34418;
  assign n21902 = ~n21612 & n21901;
  assign n21903 = ~n34420 & ~n21902;
  assign n21904 = n34420 & n21902;
  assign n21905 = ~n20831 & ~n34420;
  assign n21906 = ~n34418 & n21905;
  assign n21907 = ~n21612 & n21906;
  assign n21908 = n34420 & ~n21902;
  assign n21909 = ~n21907 & ~n21908;
  assign n21910 = ~n21903 & ~n21904;
  assign n21911 = ~n21900 & ~n34560;
  assign n21912 = ~n21897 & ~n21898;
  assign n21913 = ~n16248 & ~n21912;
  assign n21914 = n15586 & ~n21913;
  assign n21915 = ~n21911 & ~n21913;
  assign n21916 = n15586 & n21915;
  assign n21917 = ~n21911 & n21914;
  assign n21918 = ~n21804 & ~n34561;
  assign n21919 = ~n15586 & ~n21915;
  assign n21920 = n14866 & ~n21919;
  assign n21921 = ~n21918 & n21920;
  assign n21922 = ~n20865 & ~n34423;
  assign n21923 = ~n21612 & n21922;
  assign n21924 = ~n34424 & n21923;
  assign n21925 = n34424 & ~n21923;
  assign n21926 = ~n20865 & n34424;
  assign n21927 = ~n34423 & n21926;
  assign n21928 = ~n21612 & n21927;
  assign n21929 = ~n34424 & ~n21923;
  assign n21930 = ~n21928 & ~n21929;
  assign n21931 = ~n21924 & ~n21925;
  assign n21932 = ~n21921 & ~n34562;
  assign n21933 = ~n21918 & ~n21919;
  assign n21934 = ~n14866 & ~n21933;
  assign n21935 = n14233 & ~n21934;
  assign n21936 = ~n21932 & ~n21934;
  assign n21937 = n14233 & n21936;
  assign n21938 = ~n21932 & n21935;
  assign n21939 = ~n21796 & ~n34563;
  assign n21940 = ~n14233 & ~n21936;
  assign n21941 = n13548 & ~n21940;
  assign n21942 = ~n21939 & n21941;
  assign n21943 = ~n20898 & ~n34427;
  assign n21944 = ~n21612 & n21943;
  assign n21945 = ~n34428 & n21944;
  assign n21946 = n34428 & ~n21944;
  assign n21947 = ~n34428 & ~n21944;
  assign n21948 = ~n20898 & n34428;
  assign n21949 = ~n34427 & n21948;
  assign n21950 = n34428 & n21944;
  assign n21951 = ~n21612 & n21949;
  assign n21952 = ~n21947 & ~n34564;
  assign n21953 = ~n21945 & ~n21946;
  assign n21954 = ~n21942 & ~n34565;
  assign n21955 = ~n21939 & ~n21940;
  assign n21956 = ~n13548 & ~n21955;
  assign n21957 = n12948 & ~n21956;
  assign n21958 = ~n21954 & ~n21956;
  assign n21959 = n12948 & n21958;
  assign n21960 = ~n21954 & n21957;
  assign n21961 = ~n21788 & ~n34566;
  assign n21962 = ~n12948 & ~n21958;
  assign n21963 = n12296 & ~n21962;
  assign n21964 = ~n21961 & n21963;
  assign n21965 = ~n20931 & ~n34431;
  assign n21966 = ~n20931 & ~n21612;
  assign n21967 = ~n34431 & n21966;
  assign n21968 = ~n21612 & n21965;
  assign n21969 = n34433 & ~n34567;
  assign n21970 = n20946 & n21966;
  assign n21971 = ~n34433 & n34567;
  assign n21972 = ~n20931 & n34433;
  assign n21973 = ~n34431 & n21972;
  assign n21974 = ~n21612 & n21973;
  assign n21975 = ~n34433 & ~n34567;
  assign n21976 = ~n21974 & ~n21975;
  assign n21977 = ~n21969 & ~n34568;
  assign n21978 = ~n21964 & ~n34569;
  assign n21979 = ~n21961 & ~n21962;
  assign n21980 = ~n12296 & ~n21979;
  assign n21981 = n11719 & ~n21980;
  assign n21982 = ~n21978 & ~n21980;
  assign n21983 = n11719 & n21982;
  assign n21984 = ~n21978 & n21981;
  assign n21985 = ~n21780 & ~n34570;
  assign n21986 = ~n11719 & ~n21982;
  assign n21987 = n11097 & ~n21986;
  assign n21988 = ~n21985 & n21987;
  assign n21989 = ~n21772 & ~n21988;
  assign n21990 = ~n21985 & ~n21986;
  assign n21991 = ~n11097 & ~n21990;
  assign n21992 = n10555 & ~n21991;
  assign n21993 = ~n21989 & ~n21991;
  assign n21994 = n10555 & n21993;
  assign n21995 = ~n21989 & n21992;
  assign n21996 = ~n21764 & ~n34571;
  assign n21997 = ~n10555 & ~n21993;
  assign n21998 = n9969 & ~n21997;
  assign n21999 = ~n21996 & n21998;
  assign n22000 = ~n21001 & ~n34443;
  assign n22001 = ~n21001 & ~n21612;
  assign n22002 = ~n34443 & n22001;
  assign n22003 = ~n21612 & n22000;
  assign n22004 = n21009 & ~n34572;
  assign n22005 = n21013 & n22001;
  assign n22006 = ~n21001 & n21009;
  assign n22007 = ~n34443 & n22006;
  assign n22008 = ~n21612 & n22007;
  assign n22009 = ~n21009 & ~n34572;
  assign n22010 = ~n22008 & ~n22009;
  assign n22011 = ~n22004 & ~n22005;
  assign n22012 = ~n21999 & ~n34573;
  assign n22013 = ~n21996 & ~n21997;
  assign n22014 = ~n9969 & ~n22013;
  assign n22015 = n9457 & ~n22014;
  assign n22016 = ~n22012 & ~n22014;
  assign n22017 = n9457 & n22016;
  assign n22018 = ~n22012 & n22015;
  assign n22019 = ~n21756 & ~n34574;
  assign n22020 = ~n9457 & ~n22016;
  assign n22021 = n8896 & ~n22020;
  assign n22022 = ~n22019 & n22021;
  assign n22023 = ~n21748 & ~n22022;
  assign n22024 = ~n22019 & ~n22020;
  assign n22025 = ~n8896 & ~n22024;
  assign n22026 = n8411 & ~n22025;
  assign n22027 = ~n22023 & ~n22025;
  assign n22028 = n8411 & n22027;
  assign n22029 = ~n22023 & n22026;
  assign n22030 = ~n21740 & ~n34575;
  assign n22031 = ~n8411 & ~n22027;
  assign n22032 = n7885 & ~n22031;
  assign n22033 = ~n22030 & n22032;
  assign n22034 = ~n21067 & ~n34452;
  assign n22035 = ~n21067 & ~n21612;
  assign n22036 = ~n34452 & n22035;
  assign n22037 = ~n21612 & n22034;
  assign n22038 = n21075 & ~n34576;
  assign n22039 = n21079 & n22035;
  assign n22040 = ~n21067 & n21075;
  assign n22041 = ~n34452 & n22040;
  assign n22042 = ~n21612 & n22041;
  assign n22043 = ~n21075 & ~n34576;
  assign n22044 = ~n22042 & ~n22043;
  assign n22045 = ~n22038 & ~n22039;
  assign n22046 = ~n22033 & ~n34577;
  assign n22047 = ~n22030 & ~n22031;
  assign n22048 = ~n7885 & ~n22047;
  assign n22049 = n7428 & ~n22048;
  assign n22050 = ~n22046 & ~n22048;
  assign n22051 = n7428 & n22050;
  assign n22052 = ~n22046 & n22049;
  assign n22053 = ~n21732 & ~n34578;
  assign n22054 = ~n7428 & ~n22050;
  assign n22055 = n6937 & ~n22054;
  assign n22056 = ~n22053 & n22055;
  assign n22057 = ~n21724 & ~n22056;
  assign n22058 = ~n22053 & ~n22054;
  assign n22059 = ~n6937 & ~n22058;
  assign n22060 = n6507 & ~n22059;
  assign n22061 = ~n22057 & ~n22059;
  assign n22062 = n6507 & n22061;
  assign n22063 = ~n22057 & n22060;
  assign n22064 = ~n21716 & ~n34579;
  assign n22065 = ~n6507 & ~n22061;
  assign n22066 = n6051 & ~n22065;
  assign n22067 = ~n22064 & n22066;
  assign n22068 = ~n21133 & ~n34461;
  assign n22069 = ~n21133 & ~n21612;
  assign n22070 = ~n34461 & n22069;
  assign n22071 = ~n21612 & n22068;
  assign n22072 = n21141 & ~n34580;
  assign n22073 = n21145 & n22069;
  assign n22074 = ~n21133 & n21141;
  assign n22075 = ~n34461 & n22074;
  assign n22076 = ~n21612 & n22075;
  assign n22077 = ~n21141 & ~n34580;
  assign n22078 = ~n22076 & ~n22077;
  assign n22079 = ~n22072 & ~n22073;
  assign n22080 = ~n22067 & ~n34581;
  assign n22081 = ~n22064 & ~n22065;
  assign n22082 = ~n6051 & ~n22081;
  assign n22083 = n5648 & ~n22082;
  assign n22084 = ~n22080 & ~n22082;
  assign n22085 = n5648 & n22084;
  assign n22086 = ~n22080 & n22083;
  assign n22087 = ~n21708 & ~n34582;
  assign n22088 = ~n5648 & ~n22084;
  assign n22089 = n5223 & ~n22088;
  assign n22090 = ~n22087 & n22089;
  assign n22091 = ~n21700 & ~n22090;
  assign n22092 = ~n22087 & ~n22088;
  assign n22093 = ~n5223 & ~n22092;
  assign n22094 = n4851 & ~n22093;
  assign n22095 = ~n22091 & ~n22093;
  assign n22096 = n4851 & n22095;
  assign n22097 = ~n22091 & n22094;
  assign n22098 = ~n21692 & ~n34583;
  assign n22099 = ~n4851 & ~n22095;
  assign n22100 = n4461 & ~n22099;
  assign n22101 = ~n22098 & n22100;
  assign n22102 = ~n21199 & ~n34470;
  assign n22103 = ~n21199 & ~n21612;
  assign n22104 = ~n34470 & n22103;
  assign n22105 = ~n21612 & n22102;
  assign n22106 = n21207 & ~n34584;
  assign n22107 = n21211 & n22103;
  assign n22108 = ~n21199 & n21207;
  assign n22109 = ~n34470 & n22108;
  assign n22110 = ~n21612 & n22109;
  assign n22111 = ~n21207 & ~n34584;
  assign n22112 = ~n22110 & ~n22111;
  assign n22113 = ~n22106 & ~n22107;
  assign n22114 = ~n22101 & ~n34585;
  assign n22115 = ~n22098 & ~n22099;
  assign n22116 = ~n4461 & ~n22115;
  assign n22117 = n4115 & ~n22116;
  assign n22118 = ~n22114 & ~n22116;
  assign n22119 = n4115 & n22118;
  assign n22120 = ~n22114 & n22117;
  assign n22121 = ~n21684 & ~n34586;
  assign n22122 = ~n4115 & ~n22118;
  assign n22123 = n3754 & ~n22122;
  assign n22124 = ~n22121 & n22123;
  assign n22125 = ~n21676 & ~n22124;
  assign n22126 = ~n22121 & ~n22122;
  assign n22127 = ~n3754 & ~n22126;
  assign n22128 = n3444 & ~n22127;
  assign n22129 = ~n22125 & ~n22127;
  assign n22130 = n3444 & n22129;
  assign n22131 = ~n22125 & n22128;
  assign n22132 = ~n21668 & ~n34587;
  assign n22133 = ~n3444 & ~n22129;
  assign n22134 = n3116 & ~n22133;
  assign n22135 = ~n22132 & n22134;
  assign n22136 = ~n21265 & ~n34479;
  assign n22137 = ~n21265 & ~n21612;
  assign n22138 = ~n34479 & n22137;
  assign n22139 = ~n21612 & n22136;
  assign n22140 = n21273 & ~n34588;
  assign n22141 = n21277 & n22137;
  assign n22142 = ~n21265 & n21273;
  assign n22143 = ~n34479 & n22142;
  assign n22144 = ~n21612 & n22143;
  assign n22145 = ~n21273 & ~n34588;
  assign n22146 = ~n22144 & ~n22145;
  assign n22147 = ~n22140 & ~n22141;
  assign n22148 = ~n22135 & ~n34589;
  assign n22149 = ~n22132 & ~n22133;
  assign n22150 = ~n3116 & ~n22149;
  assign n22151 = n2833 & ~n22150;
  assign n22152 = ~n22148 & ~n22150;
  assign n22153 = n2833 & n22152;
  assign n22154 = ~n22148 & n22151;
  assign n22155 = ~n21660 & ~n34590;
  assign n22156 = ~n2833 & ~n22152;
  assign n22157 = n2536 & ~n22156;
  assign n22158 = ~n22155 & n22157;
  assign n22159 = ~n21652 & ~n22158;
  assign n22160 = ~n22155 & ~n22156;
  assign n22161 = ~n2536 & ~n22160;
  assign n22162 = n2283 & ~n22161;
  assign n22163 = ~n22159 & ~n22161;
  assign n22164 = n2283 & n22163;
  assign n22165 = ~n22159 & n22162;
  assign n22166 = ~n21644 & ~n34591;
  assign n22167 = ~n2283 & ~n22163;
  assign n22168 = n2021 & ~n22167;
  assign n22169 = ~n22166 & n22168;
  assign n22170 = ~n21331 & ~n34488;
  assign n22171 = ~n21331 & ~n21612;
  assign n22172 = ~n34488 & n22171;
  assign n22173 = ~n21612 & n22170;
  assign n22174 = n21339 & ~n34592;
  assign n22175 = n21343 & n22171;
  assign n22176 = ~n21331 & n21339;
  assign n22177 = ~n34488 & n22176;
  assign n22178 = ~n21612 & n22177;
  assign n22179 = ~n21339 & ~n34592;
  assign n22180 = ~n22178 & ~n22179;
  assign n22181 = ~n22174 & ~n22175;
  assign n22182 = ~n22169 & ~n34593;
  assign n22183 = ~n22166 & ~n22167;
  assign n22184 = ~n2021 & ~n22183;
  assign n22185 = n1796 & ~n22184;
  assign n22186 = ~n22182 & ~n22184;
  assign n22187 = n1796 & n22186;
  assign n22188 = ~n22182 & n22185;
  assign n22189 = ~n21636 & ~n34594;
  assign n22190 = ~n1796 & ~n22186;
  assign n22191 = n1567 & ~n22190;
  assign n22192 = ~n22189 & n22191;
  assign n22193 = ~n21628 & ~n22192;
  assign n22194 = ~n22189 & ~n22190;
  assign n22195 = ~n1567 & ~n22194;
  assign n22196 = n1374 & ~n22195;
  assign n22197 = ~n22193 & ~n22195;
  assign n22198 = n1374 & n22197;
  assign n22199 = ~n22193 & n22196;
  assign n22200 = ~n21620 & ~n34595;
  assign n22201 = ~n1374 & ~n22197;
  assign n22202 = ~n22200 & ~n22201;
  assign n22203 = ~n1179 & ~n22202;
  assign n22204 = ~n21395 & n21403;
  assign n22205 = ~n34496 & n22204;
  assign n22206 = ~n21395 & ~n34496;
  assign n22207 = ~n21612 & n22206;
  assign n22208 = n21403 & n22207;
  assign n22209 = ~n21612 & n22205;
  assign n22210 = ~n21403 & ~n22207;
  assign n22211 = ~n34596 & ~n22210;
  assign n22212 = n1179 & ~n22201;
  assign n22213 = ~n22200 & n22212;
  assign n22214 = ~n22211 & ~n22213;
  assign n22215 = ~n22203 & ~n22214;
  assign n22216 = ~n1016 & ~n22215;
  assign n22217 = ~n21409 & ~n21411;
  assign n22218 = ~n21612 & n22217;
  assign n22219 = ~n34498 & ~n22218;
  assign n22220 = ~n21411 & n34498;
  assign n22221 = ~n21409 & n22220;
  assign n22222 = n34498 & n22218;
  assign n22223 = ~n21612 & n22221;
  assign n22224 = ~n22219 & ~n34597;
  assign n22225 = n1016 & ~n22203;
  assign n22226 = n1016 & n22215;
  assign n22227 = ~n22214 & n22225;
  assign n22228 = ~n22224 & ~n34598;
  assign n22229 = ~n22216 & ~n22228;
  assign n22230 = ~n855 & ~n22229;
  assign n22231 = n855 & ~n22216;
  assign n22232 = ~n22228 & n22231;
  assign n22233 = ~n21426 & ~n34500;
  assign n22234 = ~n21426 & ~n21612;
  assign n22235 = ~n34500 & n22234;
  assign n22236 = ~n21612 & n22233;
  assign n22237 = n21434 & ~n34599;
  assign n22238 = n21438 & n22234;
  assign n22239 = ~n21426 & n21434;
  assign n22240 = ~n34500 & n22239;
  assign n22241 = ~n21612 & n22240;
  assign n22242 = ~n21434 & ~n34599;
  assign n22243 = ~n22241 & ~n22242;
  assign n22244 = ~n22237 & ~n22238;
  assign n22245 = ~n22232 & ~n34600;
  assign n22246 = ~n22230 & ~n22245;
  assign n22247 = ~n720 & ~n22246;
  assign n22248 = ~n21440 & ~n21442;
  assign n22249 = ~n21612 & n22248;
  assign n22250 = ~n34502 & ~n22249;
  assign n22251 = ~n21442 & n34502;
  assign n22252 = ~n21440 & n22251;
  assign n22253 = n34502 & n22249;
  assign n22254 = ~n21612 & n22252;
  assign n22255 = ~n22250 & ~n34601;
  assign n22256 = n720 & ~n22230;
  assign n22257 = n720 & n22246;
  assign n22258 = ~n22245 & n22256;
  assign n22259 = ~n22255 & ~n34602;
  assign n22260 = ~n22247 & ~n22259;
  assign n22261 = ~n592 & ~n22260;
  assign n22262 = n592 & ~n22247;
  assign n22263 = ~n22259 & n22262;
  assign n22264 = ~n21457 & ~n34504;
  assign n22265 = ~n21457 & ~n21612;
  assign n22266 = ~n34504 & n22265;
  assign n22267 = ~n21612 & n22264;
  assign n22268 = n21465 & ~n34603;
  assign n22269 = n21469 & n22265;
  assign n22270 = ~n21457 & n21465;
  assign n22271 = ~n34504 & n22270;
  assign n22272 = ~n21612 & n22271;
  assign n22273 = ~n21465 & ~n34603;
  assign n22274 = ~n22272 & ~n22273;
  assign n22275 = ~n22268 & ~n22269;
  assign n22276 = ~n22263 & ~n34604;
  assign n22277 = ~n22261 & ~n22276;
  assign n22278 = ~n487 & ~n22277;
  assign n22279 = ~n21471 & ~n21473;
  assign n22280 = ~n21612 & n22279;
  assign n22281 = ~n34506 & ~n22280;
  assign n22282 = ~n21473 & n34506;
  assign n22283 = ~n21471 & n22282;
  assign n22284 = n34506 & n22280;
  assign n22285 = ~n21612 & n22283;
  assign n22286 = ~n22281 & ~n34605;
  assign n22287 = n487 & ~n22261;
  assign n22288 = n487 & n22277;
  assign n22289 = ~n22276 & n22287;
  assign n22290 = ~n22286 & ~n34606;
  assign n22291 = ~n22278 & ~n22290;
  assign n22292 = ~n393 & ~n22291;
  assign n22293 = ~n21488 & ~n34507;
  assign n22294 = ~n21612 & n22293;
  assign n22295 = ~n34509 & ~n22294;
  assign n22296 = ~n21488 & n34509;
  assign n22297 = ~n34507 & n22296;
  assign n22298 = n34509 & n22294;
  assign n22299 = ~n21612 & n22297;
  assign n22300 = ~n22295 & ~n34607;
  assign n22301 = n393 & ~n22278;
  assign n22302 = ~n22290 & n22301;
  assign n22303 = ~n22300 & ~n22302;
  assign n22304 = ~n22292 & ~n22303;
  assign n22305 = ~n321 & ~n22304;
  assign n22306 = ~n21506 & ~n21508;
  assign n22307 = ~n21612 & n22306;
  assign n22308 = ~n34511 & ~n22307;
  assign n22309 = ~n21508 & n34511;
  assign n22310 = ~n21506 & n22309;
  assign n22311 = n34511 & n22307;
  assign n22312 = ~n21612 & n22310;
  assign n22313 = ~n22308 & ~n34608;
  assign n22314 = n321 & ~n22292;
  assign n22315 = n321 & n22304;
  assign n22316 = ~n22303 & n22314;
  assign n22317 = ~n22313 & ~n34609;
  assign n22318 = ~n22305 & ~n22317;
  assign n22319 = ~n263 & ~n22318;
  assign n22320 = n263 & ~n22305;
  assign n22321 = ~n22317 & n22320;
  assign n22322 = ~n21523 & ~n34513;
  assign n22323 = ~n21523 & ~n21612;
  assign n22324 = ~n34513 & n22323;
  assign n22325 = ~n21612 & n22322;
  assign n22326 = n21531 & ~n34610;
  assign n22327 = n21535 & n22323;
  assign n22328 = ~n21523 & n21531;
  assign n22329 = ~n34513 & n22328;
  assign n22330 = ~n21612 & n22329;
  assign n22331 = ~n21531 & ~n34610;
  assign n22332 = ~n22330 & ~n22331;
  assign n22333 = ~n22326 & ~n22327;
  assign n22334 = ~n22321 & ~n34611;
  assign n22335 = ~n22319 & ~n22334;
  assign n22336 = ~n214 & ~n22335;
  assign n22337 = ~n21537 & ~n21539;
  assign n22338 = ~n21612 & n22337;
  assign n22339 = ~n34515 & ~n22338;
  assign n22340 = ~n21539 & n34515;
  assign n22341 = ~n21537 & n22340;
  assign n22342 = n34515 & n22338;
  assign n22343 = ~n21612 & n22341;
  assign n22344 = ~n22339 & ~n34612;
  assign n22345 = n214 & ~n22319;
  assign n22346 = n214 & n22335;
  assign n22347 = ~n22334 & n22345;
  assign n22348 = ~n22344 & ~n34613;
  assign n22349 = ~n22336 & ~n22348;
  assign n22350 = ~n197 & ~n22349;
  assign n22351 = ~n21554 & ~n34516;
  assign n22352 = ~n21612 & n22351;
  assign n22353 = ~n34518 & ~n22352;
  assign n22354 = ~n21554 & n34518;
  assign n22355 = ~n34516 & n22354;
  assign n22356 = n34518 & n22352;
  assign n22357 = ~n21612 & n22355;
  assign n22358 = ~n22353 & ~n34614;
  assign n22359 = n197 & ~n22336;
  assign n22360 = ~n22348 & n22359;
  assign n22361 = ~n22358 & ~n22360;
  assign n22362 = ~n22350 & ~n22361;
  assign n22363 = ~n21572 & ~n21574;
  assign n22364 = ~n21612 & n22363;
  assign n22365 = ~n34520 & ~n22364;
  assign n22366 = ~n21574 & n34520;
  assign n22367 = ~n21572 & n22366;
  assign n22368 = n34520 & n22364;
  assign n22369 = ~n21612 & n22367;
  assign n22370 = ~n22365 & ~n34615;
  assign n22371 = ~n21588 & ~n21596;
  assign n22372 = ~n21596 & ~n21612;
  assign n22373 = ~n21588 & n22372;
  assign n22374 = ~n21612 & n22371;
  assign n22375 = ~n34523 & ~n34616;
  assign n22376 = ~n22370 & n22375;
  assign n22377 = ~n22362 & n22376;
  assign n22378 = n193 & ~n22377;
  assign n22379 = ~n22350 & n22370;
  assign n22380 = n22362 & n22370;
  assign n22381 = ~n22361 & n22379;
  assign n22382 = n21588 & ~n22372;
  assign n22383 = ~n193 & ~n22371;
  assign n22384 = ~n22382 & n22383;
  assign n22385 = ~n34617 & ~n22384;
  assign n22386 = ~n22378 & n22385;
  assign n22387 = pi20  & ~n22386;
  assign n22388 = ~pi18  & ~pi19 ;
  assign n22389 = ~pi20  & n22388;
  assign n22390 = ~n22387 & ~n22389;
  assign n22391 = ~n21612 & ~n22390;
  assign n22392 = ~pi20  & ~n22386;
  assign n22393 = pi21  & ~n22392;
  assign n22394 = ~pi21  & n22392;
  assign n22395 = n21834 & ~n22386;
  assign n22396 = ~n22393 & ~n34618;
  assign n22397 = ~n34407 & ~n34552;
  assign n22398 = ~n20741 & n22397;
  assign n22399 = ~n20760 & n22398;
  assign n22400 = ~n34409 & n22399;
  assign n22401 = n20746 & n20762;
  assign n22402 = ~n20754 & n22400;
  assign n22403 = ~n22389 & ~n34619;
  assign n22404 = ~n21610 & n22403;
  assign n22405 = ~n34523 & n22404;
  assign n22406 = ~n21604 & n22405;
  assign n22407 = n21612 & n22390;
  assign n22408 = ~n22387 & n22406;
  assign n22409 = n22396 & ~n34620;
  assign n22410 = ~n22391 & ~n22409;
  assign n22411 = ~n20762 & ~n22410;
  assign n22412 = n20762 & ~n22391;
  assign n22413 = ~n22409 & n22412;
  assign n22414 = ~n21612 & ~n22384;
  assign n22415 = ~n34617 & n22414;
  assign n22416 = ~n22378 & n22415;
  assign n22417 = ~n34618 & ~n22416;
  assign n22418 = pi22  & ~n22417;
  assign n22419 = ~pi22  & ~n22416;
  assign n22420 = ~pi22  & n22417;
  assign n22421 = ~n34618 & n22419;
  assign n22422 = ~n22418 & ~n34621;
  assign n22423 = ~n22413 & ~n22422;
  assign n22424 = ~n22411 & ~n22423;
  assign n22425 = ~n20011 & ~n22424;
  assign n22426 = n20011 & ~n22411;
  assign n22427 = ~n22423 & n22426;
  assign n22428 = n20011 & n22424;
  assign n22429 = ~n34553 & ~n21852;
  assign n22430 = ~n22386 & n22429;
  assign n22431 = n21850 & ~n22430;
  assign n22432 = ~n21850 & n22429;
  assign n22433 = ~n21850 & n22430;
  assign n22434 = ~n22386 & n22432;
  assign n22435 = ~n22431 & ~n34623;
  assign n22436 = ~n34622 & ~n22435;
  assign n22437 = ~n22425 & ~n22436;
  assign n22438 = ~n19190 & ~n22437;
  assign n22439 = n19190 & ~n22425;
  assign n22440 = ~n22436 & n22439;
  assign n22441 = ~n34554 & ~n21858;
  assign n22442 = ~n21858 & ~n22386;
  assign n22443 = ~n34554 & n22442;
  assign n22444 = ~n22386 & n22441;
  assign n22445 = n21832 & ~n34624;
  assign n22446 = n21857 & n22442;
  assign n22447 = n21832 & ~n34554;
  assign n22448 = ~n21858 & n22447;
  assign n22449 = ~n22386 & n22448;
  assign n22450 = ~n21832 & ~n34624;
  assign n22451 = ~n22449 & ~n22450;
  assign n22452 = ~n22445 & ~n22446;
  assign n22453 = ~n22440 & ~n34625;
  assign n22454 = ~n22438 & ~n22453;
  assign n22455 = ~n18472 & ~n22454;
  assign n22456 = n18472 & ~n22438;
  assign n22457 = ~n22453 & n22456;
  assign n22458 = n18472 & n22454;
  assign n22459 = ~n21860 & ~n21870;
  assign n22460 = ~n22386 & n22459;
  assign n22461 = ~n21867 & ~n22460;
  assign n22462 = n21867 & ~n21870;
  assign n22463 = ~n21860 & n22462;
  assign n22464 = n21867 & n22460;
  assign n22465 = ~n22386 & n22463;
  assign n22466 = n21867 & ~n22460;
  assign n22467 = ~n21867 & n22460;
  assign n22468 = ~n22466 & ~n22467;
  assign n22469 = ~n22461 & ~n34627;
  assign n22470 = ~n34626 & n34628;
  assign n22471 = ~n22455 & ~n22470;
  assign n22472 = ~n17690 & ~n22471;
  assign n22473 = n17690 & ~n22455;
  assign n22474 = ~n22470 & n22473;
  assign n22475 = ~n34556 & ~n21876;
  assign n22476 = ~n21876 & ~n22386;
  assign n22477 = ~n34556 & n22476;
  assign n22478 = ~n22386 & n22475;
  assign n22479 = n21820 & ~n34629;
  assign n22480 = n21875 & n22476;
  assign n22481 = n21820 & ~n34556;
  assign n22482 = ~n21876 & n22481;
  assign n22483 = ~n22386 & n22482;
  assign n22484 = ~n21820 & ~n34629;
  assign n22485 = ~n22483 & ~n22484;
  assign n22486 = ~n22479 & ~n22480;
  assign n22487 = ~n22474 & ~n34630;
  assign n22488 = ~n22472 & ~n22487;
  assign n22489 = ~n17001 & ~n22488;
  assign n22490 = n17001 & ~n22472;
  assign n22491 = ~n22487 & n22490;
  assign n22492 = n17001 & n22488;
  assign n22493 = ~n21878 & ~n21892;
  assign n22494 = ~n22386 & n22493;
  assign n22495 = ~n34558 & ~n22494;
  assign n22496 = n34558 & n22494;
  assign n22497 = ~n34558 & ~n21892;
  assign n22498 = ~n21878 & n22497;
  assign n22499 = ~n22386 & n22498;
  assign n22500 = n34558 & ~n22494;
  assign n22501 = ~n22499 & ~n22500;
  assign n22502 = ~n22495 & ~n22496;
  assign n22503 = ~n34631 & ~n34632;
  assign n22504 = ~n22489 & ~n22503;
  assign n22505 = ~n16248 & ~n22504;
  assign n22506 = n16248 & ~n22489;
  assign n22507 = ~n22503 & n22506;
  assign n22508 = ~n34559 & ~n21898;
  assign n22509 = ~n21898 & ~n22386;
  assign n22510 = ~n34559 & n22509;
  assign n22511 = ~n22386 & n22508;
  assign n22512 = n21812 & ~n34633;
  assign n22513 = n21897 & n22509;
  assign n22514 = n21812 & ~n34559;
  assign n22515 = ~n21898 & n22514;
  assign n22516 = ~n22386 & n22515;
  assign n22517 = ~n21812 & ~n34633;
  assign n22518 = ~n22516 & ~n22517;
  assign n22519 = ~n22512 & ~n22513;
  assign n22520 = ~n22507 & ~n34634;
  assign n22521 = ~n22505 & ~n22520;
  assign n22522 = ~n15586 & ~n22521;
  assign n22523 = n15586 & ~n22505;
  assign n22524 = ~n22520 & n22523;
  assign n22525 = n15586 & n22521;
  assign n22526 = ~n21900 & ~n21913;
  assign n22527 = ~n22386 & n22526;
  assign n22528 = ~n34560 & n22527;
  assign n22529 = n34560 & ~n22527;
  assign n22530 = n34560 & ~n21913;
  assign n22531 = ~n21900 & n22530;
  assign n22532 = ~n22386 & n22531;
  assign n22533 = ~n34560 & ~n22527;
  assign n22534 = ~n22532 & ~n22533;
  assign n22535 = ~n22528 & ~n22529;
  assign n22536 = ~n34635 & ~n34636;
  assign n22537 = ~n22522 & ~n22536;
  assign n22538 = ~n14866 & ~n22537;
  assign n22539 = n14866 & ~n22522;
  assign n22540 = ~n22536 & n22539;
  assign n22541 = ~n34561 & ~n21919;
  assign n22542 = ~n21919 & ~n22386;
  assign n22543 = ~n34561 & n22542;
  assign n22544 = ~n22386 & n22541;
  assign n22545 = n21804 & ~n34637;
  assign n22546 = n21918 & n22542;
  assign n22547 = n21804 & ~n34561;
  assign n22548 = ~n21919 & n22547;
  assign n22549 = ~n22386 & n22548;
  assign n22550 = ~n21804 & ~n34637;
  assign n22551 = ~n22549 & ~n22550;
  assign n22552 = ~n22545 & ~n22546;
  assign n22553 = ~n22540 & ~n34638;
  assign n22554 = ~n22538 & ~n22553;
  assign n22555 = ~n14233 & ~n22554;
  assign n22556 = n14233 & ~n22538;
  assign n22557 = ~n22553 & n22556;
  assign n22558 = n14233 & n22554;
  assign n22559 = ~n21921 & ~n21934;
  assign n22560 = ~n22386 & n22559;
  assign n22561 = ~n34562 & n22560;
  assign n22562 = n34562 & ~n22560;
  assign n22563 = ~n34562 & ~n22560;
  assign n22564 = n34562 & ~n21934;
  assign n22565 = ~n21921 & n22564;
  assign n22566 = n34562 & n22560;
  assign n22567 = ~n22386 & n22565;
  assign n22568 = ~n22563 & ~n34640;
  assign n22569 = ~n22561 & ~n22562;
  assign n22570 = ~n34639 & ~n34641;
  assign n22571 = ~n22555 & ~n22570;
  assign n22572 = ~n13548 & ~n22571;
  assign n22573 = n13548 & ~n22555;
  assign n22574 = ~n22570 & n22573;
  assign n22575 = ~n34563 & ~n21940;
  assign n22576 = ~n21940 & ~n22386;
  assign n22577 = ~n34563 & n22576;
  assign n22578 = ~n22386 & n22575;
  assign n22579 = n21796 & ~n34642;
  assign n22580 = n21939 & n22576;
  assign n22581 = n21796 & ~n34563;
  assign n22582 = ~n21940 & n22581;
  assign n22583 = ~n22386 & n22582;
  assign n22584 = ~n21796 & ~n34642;
  assign n22585 = ~n22583 & ~n22584;
  assign n22586 = ~n22579 & ~n22580;
  assign n22587 = ~n22574 & ~n34643;
  assign n22588 = ~n22572 & ~n22587;
  assign n22589 = ~n12948 & ~n22588;
  assign n22590 = n12948 & ~n22572;
  assign n22591 = ~n22587 & n22590;
  assign n22592 = n12948 & n22588;
  assign n22593 = ~n21942 & ~n21956;
  assign n22594 = ~n21956 & ~n22386;
  assign n22595 = ~n21942 & n22594;
  assign n22596 = ~n22386 & n22593;
  assign n22597 = n34565 & ~n34645;
  assign n22598 = n21954 & n22594;
  assign n22599 = ~n34565 & n34645;
  assign n22600 = n34565 & ~n21956;
  assign n22601 = ~n21942 & n22600;
  assign n22602 = ~n22386 & n22601;
  assign n22603 = ~n34565 & ~n34645;
  assign n22604 = ~n22602 & ~n22603;
  assign n22605 = ~n22597 & ~n34646;
  assign n22606 = ~n34644 & ~n34647;
  assign n22607 = ~n22589 & ~n22606;
  assign n22608 = ~n12296 & ~n22607;
  assign n22609 = n12296 & ~n22589;
  assign n22610 = ~n22606 & n22609;
  assign n22611 = ~n34566 & ~n21962;
  assign n22612 = ~n21962 & ~n22386;
  assign n22613 = ~n34566 & n22612;
  assign n22614 = ~n22386 & n22611;
  assign n22615 = n21788 & ~n34648;
  assign n22616 = n21961 & n22612;
  assign n22617 = n21788 & ~n34566;
  assign n22618 = ~n21962 & n22617;
  assign n22619 = ~n22386 & n22618;
  assign n22620 = ~n21788 & ~n34648;
  assign n22621 = ~n22619 & ~n22620;
  assign n22622 = ~n22615 & ~n22616;
  assign n22623 = ~n22610 & ~n34649;
  assign n22624 = ~n22608 & ~n22623;
  assign n22625 = ~n11719 & ~n22624;
  assign n22626 = ~n21964 & ~n21980;
  assign n22627 = ~n22386 & n22626;
  assign n22628 = ~n34569 & ~n22627;
  assign n22629 = n34569 & ~n21980;
  assign n22630 = ~n21964 & n22629;
  assign n22631 = n34569 & n22627;
  assign n22632 = ~n22386 & n22630;
  assign n22633 = ~n22628 & ~n34650;
  assign n22634 = n11719 & ~n22608;
  assign n22635 = ~n22623 & n22634;
  assign n22636 = n11719 & n22624;
  assign n22637 = ~n22633 & ~n34651;
  assign n22638 = ~n22625 & ~n22637;
  assign n22639 = ~n11097 & ~n22638;
  assign n22640 = n11097 & ~n22625;
  assign n22641 = ~n22637 & n22640;
  assign n22642 = ~n34570 & ~n21986;
  assign n22643 = ~n21986 & ~n22386;
  assign n22644 = ~n34570 & n22643;
  assign n22645 = ~n22386 & n22642;
  assign n22646 = n21780 & ~n34652;
  assign n22647 = n21985 & n22643;
  assign n22648 = n21780 & ~n34570;
  assign n22649 = ~n21986 & n22648;
  assign n22650 = ~n22386 & n22649;
  assign n22651 = ~n21780 & ~n34652;
  assign n22652 = ~n22650 & ~n22651;
  assign n22653 = ~n22646 & ~n22647;
  assign n22654 = ~n22641 & ~n34653;
  assign n22655 = ~n22639 & ~n22654;
  assign n22656 = ~n10555 & ~n22655;
  assign n22657 = n10555 & ~n22639;
  assign n22658 = ~n22654 & n22657;
  assign n22659 = n10555 & n22655;
  assign n22660 = ~n21988 & ~n21991;
  assign n22661 = ~n21991 & ~n22386;
  assign n22662 = ~n21988 & n22661;
  assign n22663 = ~n22386 & n22660;
  assign n22664 = n21772 & ~n34655;
  assign n22665 = n21989 & n22661;
  assign n22666 = n21772 & ~n21991;
  assign n22667 = ~n21988 & n22666;
  assign n22668 = ~n22386 & n22667;
  assign n22669 = ~n21772 & ~n34655;
  assign n22670 = ~n22668 & ~n22669;
  assign n22671 = ~n22664 & ~n22665;
  assign n22672 = ~n34654 & ~n34656;
  assign n22673 = ~n22656 & ~n22672;
  assign n22674 = ~n9969 & ~n22673;
  assign n22675 = n9969 & ~n22656;
  assign n22676 = ~n22672 & n22675;
  assign n22677 = ~n34571 & ~n21997;
  assign n22678 = ~n21997 & ~n22386;
  assign n22679 = ~n34571 & n22678;
  assign n22680 = ~n22386 & n22677;
  assign n22681 = n21764 & ~n34657;
  assign n22682 = n21996 & n22678;
  assign n22683 = n21764 & ~n34571;
  assign n22684 = ~n21997 & n22683;
  assign n22685 = ~n22386 & n22684;
  assign n22686 = ~n21764 & ~n34657;
  assign n22687 = ~n22685 & ~n22686;
  assign n22688 = ~n22681 & ~n22682;
  assign n22689 = ~n22676 & ~n34658;
  assign n22690 = ~n22674 & ~n22689;
  assign n22691 = ~n9457 & ~n22690;
  assign n22692 = ~n21999 & ~n22014;
  assign n22693 = ~n22386 & n22692;
  assign n22694 = ~n34573 & ~n22693;
  assign n22695 = n34573 & ~n22014;
  assign n22696 = ~n21999 & n22695;
  assign n22697 = n34573 & n22693;
  assign n22698 = ~n22386 & n22696;
  assign n22699 = ~n22694 & ~n34659;
  assign n22700 = n9457 & ~n22674;
  assign n22701 = ~n22689 & n22700;
  assign n22702 = n9457 & n22690;
  assign n22703 = ~n22699 & ~n34660;
  assign n22704 = ~n22691 & ~n22703;
  assign n22705 = ~n8896 & ~n22704;
  assign n22706 = n8896 & ~n22691;
  assign n22707 = ~n22703 & n22706;
  assign n22708 = ~n34574 & ~n22020;
  assign n22709 = ~n22020 & ~n22386;
  assign n22710 = ~n34574 & n22709;
  assign n22711 = ~n22386 & n22708;
  assign n22712 = n21756 & ~n34661;
  assign n22713 = n22019 & n22709;
  assign n22714 = n21756 & ~n34574;
  assign n22715 = ~n22020 & n22714;
  assign n22716 = ~n22386 & n22715;
  assign n22717 = ~n21756 & ~n34661;
  assign n22718 = ~n22716 & ~n22717;
  assign n22719 = ~n22712 & ~n22713;
  assign n22720 = ~n22707 & ~n34662;
  assign n22721 = ~n22705 & ~n22720;
  assign n22722 = ~n8411 & ~n22721;
  assign n22723 = n8411 & ~n22705;
  assign n22724 = ~n22720 & n22723;
  assign n22725 = n8411 & n22721;
  assign n22726 = ~n22022 & ~n22025;
  assign n22727 = ~n22025 & ~n22386;
  assign n22728 = ~n22022 & n22727;
  assign n22729 = ~n22386 & n22726;
  assign n22730 = n21748 & ~n34664;
  assign n22731 = n22023 & n22727;
  assign n22732 = n21748 & ~n22025;
  assign n22733 = ~n22022 & n22732;
  assign n22734 = ~n22386 & n22733;
  assign n22735 = ~n21748 & ~n34664;
  assign n22736 = ~n22734 & ~n22735;
  assign n22737 = ~n22730 & ~n22731;
  assign n22738 = ~n34663 & ~n34665;
  assign n22739 = ~n22722 & ~n22738;
  assign n22740 = ~n7885 & ~n22739;
  assign n22741 = n7885 & ~n22722;
  assign n22742 = ~n22738 & n22741;
  assign n22743 = ~n34575 & ~n22031;
  assign n22744 = ~n22031 & ~n22386;
  assign n22745 = ~n34575 & n22744;
  assign n22746 = ~n22386 & n22743;
  assign n22747 = n21740 & ~n34666;
  assign n22748 = n22030 & n22744;
  assign n22749 = n21740 & ~n34575;
  assign n22750 = ~n22031 & n22749;
  assign n22751 = ~n22386 & n22750;
  assign n22752 = ~n21740 & ~n34666;
  assign n22753 = ~n22751 & ~n22752;
  assign n22754 = ~n22747 & ~n22748;
  assign n22755 = ~n22742 & ~n34667;
  assign n22756 = ~n22740 & ~n22755;
  assign n22757 = ~n7428 & ~n22756;
  assign n22758 = ~n22033 & ~n22048;
  assign n22759 = ~n22386 & n22758;
  assign n22760 = ~n34577 & ~n22759;
  assign n22761 = n34577 & ~n22048;
  assign n22762 = ~n22033 & n22761;
  assign n22763 = n34577 & n22759;
  assign n22764 = ~n22386 & n22762;
  assign n22765 = ~n22760 & ~n34668;
  assign n22766 = n7428 & ~n22740;
  assign n22767 = ~n22755 & n22766;
  assign n22768 = n7428 & n22756;
  assign n22769 = ~n22765 & ~n34669;
  assign n22770 = ~n22757 & ~n22769;
  assign n22771 = ~n6937 & ~n22770;
  assign n22772 = n6937 & ~n22757;
  assign n22773 = ~n22769 & n22772;
  assign n22774 = ~n34578 & ~n22054;
  assign n22775 = ~n22054 & ~n22386;
  assign n22776 = ~n34578 & n22775;
  assign n22777 = ~n22386 & n22774;
  assign n22778 = n21732 & ~n34670;
  assign n22779 = n22053 & n22775;
  assign n22780 = n21732 & ~n34578;
  assign n22781 = ~n22054 & n22780;
  assign n22782 = ~n22386 & n22781;
  assign n22783 = ~n21732 & ~n34670;
  assign n22784 = ~n22782 & ~n22783;
  assign n22785 = ~n22778 & ~n22779;
  assign n22786 = ~n22773 & ~n34671;
  assign n22787 = ~n22771 & ~n22786;
  assign n22788 = ~n6507 & ~n22787;
  assign n22789 = n6507 & ~n22771;
  assign n22790 = ~n22786 & n22789;
  assign n22791 = n6507 & n22787;
  assign n22792 = ~n22056 & ~n22059;
  assign n22793 = ~n22059 & ~n22386;
  assign n22794 = ~n22056 & n22793;
  assign n22795 = ~n22386 & n22792;
  assign n22796 = n21724 & ~n34673;
  assign n22797 = n22057 & n22793;
  assign n22798 = n21724 & ~n22059;
  assign n22799 = ~n22056 & n22798;
  assign n22800 = ~n22386 & n22799;
  assign n22801 = ~n21724 & ~n34673;
  assign n22802 = ~n22800 & ~n22801;
  assign n22803 = ~n22796 & ~n22797;
  assign n22804 = ~n34672 & ~n34674;
  assign n22805 = ~n22788 & ~n22804;
  assign n22806 = ~n6051 & ~n22805;
  assign n22807 = n6051 & ~n22788;
  assign n22808 = ~n22804 & n22807;
  assign n22809 = ~n34579 & ~n22065;
  assign n22810 = ~n22065 & ~n22386;
  assign n22811 = ~n34579 & n22810;
  assign n22812 = ~n22386 & n22809;
  assign n22813 = n21716 & ~n34675;
  assign n22814 = n22064 & n22810;
  assign n22815 = n21716 & ~n34579;
  assign n22816 = ~n22065 & n22815;
  assign n22817 = ~n22386 & n22816;
  assign n22818 = ~n21716 & ~n34675;
  assign n22819 = ~n22817 & ~n22818;
  assign n22820 = ~n22813 & ~n22814;
  assign n22821 = ~n22808 & ~n34676;
  assign n22822 = ~n22806 & ~n22821;
  assign n22823 = ~n5648 & ~n22822;
  assign n22824 = ~n22067 & ~n22082;
  assign n22825 = ~n22386 & n22824;
  assign n22826 = ~n34581 & ~n22825;
  assign n22827 = n34581 & ~n22082;
  assign n22828 = ~n22067 & n22827;
  assign n22829 = n34581 & n22825;
  assign n22830 = ~n22386 & n22828;
  assign n22831 = ~n22826 & ~n34677;
  assign n22832 = n5648 & ~n22806;
  assign n22833 = ~n22821 & n22832;
  assign n22834 = n5648 & n22822;
  assign n22835 = ~n22831 & ~n34678;
  assign n22836 = ~n22823 & ~n22835;
  assign n22837 = ~n5223 & ~n22836;
  assign n22838 = n5223 & ~n22823;
  assign n22839 = ~n22835 & n22838;
  assign n22840 = ~n34582 & ~n22088;
  assign n22841 = ~n22088 & ~n22386;
  assign n22842 = ~n34582 & n22841;
  assign n22843 = ~n22386 & n22840;
  assign n22844 = n21708 & ~n34679;
  assign n22845 = n22087 & n22841;
  assign n22846 = n21708 & ~n34582;
  assign n22847 = ~n22088 & n22846;
  assign n22848 = ~n22386 & n22847;
  assign n22849 = ~n21708 & ~n34679;
  assign n22850 = ~n22848 & ~n22849;
  assign n22851 = ~n22844 & ~n22845;
  assign n22852 = ~n22839 & ~n34680;
  assign n22853 = ~n22837 & ~n22852;
  assign n22854 = ~n4851 & ~n22853;
  assign n22855 = n4851 & ~n22837;
  assign n22856 = ~n22852 & n22855;
  assign n22857 = n4851 & n22853;
  assign n22858 = ~n22090 & ~n22093;
  assign n22859 = ~n22093 & ~n22386;
  assign n22860 = ~n22090 & n22859;
  assign n22861 = ~n22386 & n22858;
  assign n22862 = n21700 & ~n34682;
  assign n22863 = n22091 & n22859;
  assign n22864 = n21700 & ~n22093;
  assign n22865 = ~n22090 & n22864;
  assign n22866 = ~n22386 & n22865;
  assign n22867 = ~n21700 & ~n34682;
  assign n22868 = ~n22866 & ~n22867;
  assign n22869 = ~n22862 & ~n22863;
  assign n22870 = ~n34681 & ~n34683;
  assign n22871 = ~n22854 & ~n22870;
  assign n22872 = ~n4461 & ~n22871;
  assign n22873 = n4461 & ~n22854;
  assign n22874 = ~n22870 & n22873;
  assign n22875 = ~n34583 & ~n22099;
  assign n22876 = ~n22099 & ~n22386;
  assign n22877 = ~n34583 & n22876;
  assign n22878 = ~n22386 & n22875;
  assign n22879 = n21692 & ~n34684;
  assign n22880 = n22098 & n22876;
  assign n22881 = n21692 & ~n34583;
  assign n22882 = ~n22099 & n22881;
  assign n22883 = ~n22386 & n22882;
  assign n22884 = ~n21692 & ~n34684;
  assign n22885 = ~n22883 & ~n22884;
  assign n22886 = ~n22879 & ~n22880;
  assign n22887 = ~n22874 & ~n34685;
  assign n22888 = ~n22872 & ~n22887;
  assign n22889 = ~n4115 & ~n22888;
  assign n22890 = ~n22101 & ~n22116;
  assign n22891 = ~n22386 & n22890;
  assign n22892 = ~n34585 & ~n22891;
  assign n22893 = n34585 & ~n22116;
  assign n22894 = ~n22101 & n22893;
  assign n22895 = n34585 & n22891;
  assign n22896 = ~n22386 & n22894;
  assign n22897 = ~n22892 & ~n34686;
  assign n22898 = n4115 & ~n22872;
  assign n22899 = ~n22887 & n22898;
  assign n22900 = n4115 & n22888;
  assign n22901 = ~n22897 & ~n34687;
  assign n22902 = ~n22889 & ~n22901;
  assign n22903 = ~n3754 & ~n22902;
  assign n22904 = n3754 & ~n22889;
  assign n22905 = ~n22901 & n22904;
  assign n22906 = ~n34586 & ~n22122;
  assign n22907 = ~n22122 & ~n22386;
  assign n22908 = ~n34586 & n22907;
  assign n22909 = ~n22386 & n22906;
  assign n22910 = n21684 & ~n34688;
  assign n22911 = n22121 & n22907;
  assign n22912 = n21684 & ~n34586;
  assign n22913 = ~n22122 & n22912;
  assign n22914 = ~n22386 & n22913;
  assign n22915 = ~n21684 & ~n34688;
  assign n22916 = ~n22914 & ~n22915;
  assign n22917 = ~n22910 & ~n22911;
  assign n22918 = ~n22905 & ~n34689;
  assign n22919 = ~n22903 & ~n22918;
  assign n22920 = ~n3444 & ~n22919;
  assign n22921 = n3444 & ~n22903;
  assign n22922 = ~n22918 & n22921;
  assign n22923 = n3444 & n22919;
  assign n22924 = ~n22124 & ~n22127;
  assign n22925 = ~n22127 & ~n22386;
  assign n22926 = ~n22124 & n22925;
  assign n22927 = ~n22386 & n22924;
  assign n22928 = n21676 & ~n34691;
  assign n22929 = n22125 & n22925;
  assign n22930 = n21676 & ~n22127;
  assign n22931 = ~n22124 & n22930;
  assign n22932 = ~n22386 & n22931;
  assign n22933 = ~n21676 & ~n34691;
  assign n22934 = ~n22932 & ~n22933;
  assign n22935 = ~n22928 & ~n22929;
  assign n22936 = ~n34690 & ~n34692;
  assign n22937 = ~n22920 & ~n22936;
  assign n22938 = ~n3116 & ~n22937;
  assign n22939 = n3116 & ~n22920;
  assign n22940 = ~n22936 & n22939;
  assign n22941 = ~n34587 & ~n22133;
  assign n22942 = ~n22133 & ~n22386;
  assign n22943 = ~n34587 & n22942;
  assign n22944 = ~n22386 & n22941;
  assign n22945 = n21668 & ~n34693;
  assign n22946 = n22132 & n22942;
  assign n22947 = n21668 & ~n34587;
  assign n22948 = ~n22133 & n22947;
  assign n22949 = ~n22386 & n22948;
  assign n22950 = ~n21668 & ~n34693;
  assign n22951 = ~n22949 & ~n22950;
  assign n22952 = ~n22945 & ~n22946;
  assign n22953 = ~n22940 & ~n34694;
  assign n22954 = ~n22938 & ~n22953;
  assign n22955 = ~n2833 & ~n22954;
  assign n22956 = ~n22135 & ~n22150;
  assign n22957 = ~n22386 & n22956;
  assign n22958 = ~n34589 & ~n22957;
  assign n22959 = n34589 & ~n22150;
  assign n22960 = ~n22135 & n22959;
  assign n22961 = n34589 & n22957;
  assign n22962 = ~n22386 & n22960;
  assign n22963 = ~n22958 & ~n34695;
  assign n22964 = n2833 & ~n22938;
  assign n22965 = ~n22953 & n22964;
  assign n22966 = n2833 & n22954;
  assign n22967 = ~n22963 & ~n34696;
  assign n22968 = ~n22955 & ~n22967;
  assign n22969 = ~n2536 & ~n22968;
  assign n22970 = n2536 & ~n22955;
  assign n22971 = ~n22967 & n22970;
  assign n22972 = ~n34590 & ~n22156;
  assign n22973 = ~n22156 & ~n22386;
  assign n22974 = ~n34590 & n22973;
  assign n22975 = ~n22386 & n22972;
  assign n22976 = n21660 & ~n34697;
  assign n22977 = n22155 & n22973;
  assign n22978 = n21660 & ~n34590;
  assign n22979 = ~n22156 & n22978;
  assign n22980 = ~n22386 & n22979;
  assign n22981 = ~n21660 & ~n34697;
  assign n22982 = ~n22980 & ~n22981;
  assign n22983 = ~n22976 & ~n22977;
  assign n22984 = ~n22971 & ~n34698;
  assign n22985 = ~n22969 & ~n22984;
  assign n22986 = ~n2283 & ~n22985;
  assign n22987 = n2283 & ~n22969;
  assign n22988 = ~n22984 & n22987;
  assign n22989 = n2283 & n22985;
  assign n22990 = ~n22158 & ~n22161;
  assign n22991 = ~n22161 & ~n22386;
  assign n22992 = ~n22158 & n22991;
  assign n22993 = ~n22386 & n22990;
  assign n22994 = n21652 & ~n34700;
  assign n22995 = n22159 & n22991;
  assign n22996 = n21652 & ~n22161;
  assign n22997 = ~n22158 & n22996;
  assign n22998 = ~n22386 & n22997;
  assign n22999 = ~n21652 & ~n34700;
  assign n23000 = ~n22998 & ~n22999;
  assign n23001 = ~n22994 & ~n22995;
  assign n23002 = ~n34699 & ~n34701;
  assign n23003 = ~n22986 & ~n23002;
  assign n23004 = ~n2021 & ~n23003;
  assign n23005 = n2021 & ~n22986;
  assign n23006 = ~n23002 & n23005;
  assign n23007 = ~n34591 & ~n22167;
  assign n23008 = ~n22167 & ~n22386;
  assign n23009 = ~n34591 & n23008;
  assign n23010 = ~n22386 & n23007;
  assign n23011 = n21644 & ~n34702;
  assign n23012 = n22166 & n23008;
  assign n23013 = n21644 & ~n34591;
  assign n23014 = ~n22167 & n23013;
  assign n23015 = ~n22386 & n23014;
  assign n23016 = ~n21644 & ~n34702;
  assign n23017 = ~n23015 & ~n23016;
  assign n23018 = ~n23011 & ~n23012;
  assign n23019 = ~n23006 & ~n34703;
  assign n23020 = ~n23004 & ~n23019;
  assign n23021 = ~n1796 & ~n23020;
  assign n23022 = ~n22169 & ~n22184;
  assign n23023 = ~n22386 & n23022;
  assign n23024 = ~n34593 & ~n23023;
  assign n23025 = n34593 & ~n22184;
  assign n23026 = ~n22169 & n23025;
  assign n23027 = n34593 & n23023;
  assign n23028 = ~n22386 & n23026;
  assign n23029 = ~n23024 & ~n34704;
  assign n23030 = n1796 & ~n23004;
  assign n23031 = ~n23019 & n23030;
  assign n23032 = n1796 & n23020;
  assign n23033 = ~n23029 & ~n34705;
  assign n23034 = ~n23021 & ~n23033;
  assign n23035 = ~n1567 & ~n23034;
  assign n23036 = n1567 & ~n23021;
  assign n23037 = ~n23033 & n23036;
  assign n23038 = ~n34594 & ~n22190;
  assign n23039 = ~n22190 & ~n22386;
  assign n23040 = ~n34594 & n23039;
  assign n23041 = ~n22386 & n23038;
  assign n23042 = n21636 & ~n34706;
  assign n23043 = n22189 & n23039;
  assign n23044 = n21636 & ~n34594;
  assign n23045 = ~n22190 & n23044;
  assign n23046 = ~n22386 & n23045;
  assign n23047 = ~n21636 & ~n34706;
  assign n23048 = ~n23046 & ~n23047;
  assign n23049 = ~n23042 & ~n23043;
  assign n23050 = ~n23037 & ~n34707;
  assign n23051 = ~n23035 & ~n23050;
  assign n23052 = ~n1374 & ~n23051;
  assign n23053 = n1374 & ~n23035;
  assign n23054 = ~n23050 & n23053;
  assign n23055 = n1374 & n23051;
  assign n23056 = ~n22192 & ~n22195;
  assign n23057 = ~n22195 & ~n22386;
  assign n23058 = ~n22192 & n23057;
  assign n23059 = ~n22386 & n23056;
  assign n23060 = n21628 & ~n34709;
  assign n23061 = n22193 & n23057;
  assign n23062 = n21628 & ~n22195;
  assign n23063 = ~n22192 & n23062;
  assign n23064 = ~n22386 & n23063;
  assign n23065 = ~n21628 & ~n34709;
  assign n23066 = ~n23064 & ~n23065;
  assign n23067 = ~n23060 & ~n23061;
  assign n23068 = ~n34708 & ~n34710;
  assign n23069 = ~n23052 & ~n23068;
  assign n23070 = ~n1179 & ~n23069;
  assign n23071 = n1179 & ~n23052;
  assign n23072 = ~n23068 & n23071;
  assign n23073 = n21620 & ~n34595;
  assign n23074 = ~n22201 & n23073;
  assign n23075 = ~n34595 & ~n22201;
  assign n23076 = ~n22386 & n23075;
  assign n23077 = n21620 & n23076;
  assign n23078 = ~n22386 & n23074;
  assign n23079 = ~n21620 & ~n23076;
  assign n23080 = ~n34711 & ~n23079;
  assign n23081 = ~n23072 & ~n23080;
  assign n23082 = ~n23070 & ~n23081;
  assign n23083 = ~n1016 & ~n23082;
  assign n23084 = ~n22203 & ~n22213;
  assign n23085 = ~n22386 & n23084;
  assign n23086 = ~n22211 & ~n23085;
  assign n23087 = ~n22203 & n22211;
  assign n23088 = ~n22213 & n23087;
  assign n23089 = n22211 & n23085;
  assign n23090 = ~n22386 & n23088;
  assign n23091 = ~n23086 & ~n34712;
  assign n23092 = n1016 & ~n23070;
  assign n23093 = ~n23081 & n23092;
  assign n23094 = n1016 & n23082;
  assign n23095 = ~n23091 & ~n34713;
  assign n23096 = ~n23083 & ~n23095;
  assign n23097 = ~n855 & ~n23096;
  assign n23098 = n855 & ~n23083;
  assign n23099 = ~n23095 & n23098;
  assign n23100 = ~n22216 & ~n34598;
  assign n23101 = ~n22216 & ~n22386;
  assign n23102 = ~n34598 & n23101;
  assign n23103 = ~n22386 & n23100;
  assign n23104 = n22224 & ~n34714;
  assign n23105 = n22228 & n23101;
  assign n23106 = n22224 & ~n34598;
  assign n23107 = ~n22216 & n23106;
  assign n23108 = ~n22386 & n23107;
  assign n23109 = ~n22224 & ~n34714;
  assign n23110 = ~n23108 & ~n23109;
  assign n23111 = ~n23104 & ~n23105;
  assign n23112 = ~n23099 & ~n34715;
  assign n23113 = ~n23097 & ~n23112;
  assign n23114 = ~n720 & ~n23113;
  assign n23115 = ~n22230 & ~n22232;
  assign n23116 = ~n22386 & n23115;
  assign n23117 = ~n34600 & ~n23116;
  assign n23118 = ~n22230 & n34600;
  assign n23119 = ~n22232 & n23118;
  assign n23120 = n34600 & n23116;
  assign n23121 = ~n22386 & n23119;
  assign n23122 = ~n23117 & ~n34716;
  assign n23123 = n720 & ~n23097;
  assign n23124 = ~n23112 & n23123;
  assign n23125 = n720 & n23113;
  assign n23126 = ~n23122 & ~n34717;
  assign n23127 = ~n23114 & ~n23126;
  assign n23128 = ~n592 & ~n23127;
  assign n23129 = n592 & ~n23114;
  assign n23130 = ~n23126 & n23129;
  assign n23131 = ~n22247 & ~n34602;
  assign n23132 = ~n22247 & ~n22386;
  assign n23133 = ~n34602 & n23132;
  assign n23134 = ~n22386 & n23131;
  assign n23135 = n22255 & ~n34718;
  assign n23136 = n22259 & n23132;
  assign n23137 = n22255 & ~n34602;
  assign n23138 = ~n22247 & n23137;
  assign n23139 = ~n22386 & n23138;
  assign n23140 = ~n22255 & ~n34718;
  assign n23141 = ~n23139 & ~n23140;
  assign n23142 = ~n23135 & ~n23136;
  assign n23143 = ~n23130 & ~n34719;
  assign n23144 = ~n23128 & ~n23143;
  assign n23145 = ~n487 & ~n23144;
  assign n23146 = ~n22261 & ~n22263;
  assign n23147 = ~n22386 & n23146;
  assign n23148 = ~n34604 & ~n23147;
  assign n23149 = ~n22261 & n34604;
  assign n23150 = ~n22263 & n23149;
  assign n23151 = n34604 & n23147;
  assign n23152 = ~n22386 & n23150;
  assign n23153 = ~n23148 & ~n34720;
  assign n23154 = n487 & ~n23128;
  assign n23155 = ~n23143 & n23154;
  assign n23156 = n487 & n23144;
  assign n23157 = ~n23153 & ~n34721;
  assign n23158 = ~n23145 & ~n23157;
  assign n23159 = ~n393 & ~n23158;
  assign n23160 = n393 & ~n23145;
  assign n23161 = ~n23157 & n23160;
  assign n23162 = ~n22278 & ~n34606;
  assign n23163 = ~n22278 & ~n22386;
  assign n23164 = ~n34606 & n23163;
  assign n23165 = ~n22386 & n23162;
  assign n23166 = n22286 & ~n34722;
  assign n23167 = n22290 & n23163;
  assign n23168 = n22286 & ~n34606;
  assign n23169 = ~n22278 & n23168;
  assign n23170 = ~n22386 & n23169;
  assign n23171 = ~n22286 & ~n34722;
  assign n23172 = ~n23170 & ~n23171;
  assign n23173 = ~n23166 & ~n23167;
  assign n23174 = ~n23161 & ~n34723;
  assign n23175 = ~n23159 & ~n23174;
  assign n23176 = ~n321 & ~n23175;
  assign n23177 = n321 & ~n23159;
  assign n23178 = ~n23174 & n23177;
  assign n23179 = n321 & n23175;
  assign n23180 = ~n22292 & ~n22302;
  assign n23181 = ~n22292 & ~n22386;
  assign n23182 = ~n22302 & n23181;
  assign n23183 = ~n22386 & n23180;
  assign n23184 = n22300 & ~n34725;
  assign n23185 = n22303 & n23181;
  assign n23186 = ~n22292 & n22300;
  assign n23187 = ~n22302 & n23186;
  assign n23188 = ~n22386 & n23187;
  assign n23189 = ~n22300 & ~n34725;
  assign n23190 = ~n23188 & ~n23189;
  assign n23191 = ~n23184 & ~n23185;
  assign n23192 = ~n34724 & ~n34726;
  assign n23193 = ~n23176 & ~n23192;
  assign n23194 = ~n263 & ~n23193;
  assign n23195 = n263 & ~n23176;
  assign n23196 = ~n23192 & n23195;
  assign n23197 = ~n22305 & ~n34609;
  assign n23198 = ~n22305 & ~n22386;
  assign n23199 = ~n34609 & n23198;
  assign n23200 = ~n22386 & n23197;
  assign n23201 = n22313 & ~n34727;
  assign n23202 = n22317 & n23198;
  assign n23203 = n22313 & ~n34609;
  assign n23204 = ~n22305 & n23203;
  assign n23205 = ~n22386 & n23204;
  assign n23206 = ~n22313 & ~n34727;
  assign n23207 = ~n23205 & ~n23206;
  assign n23208 = ~n23201 & ~n23202;
  assign n23209 = ~n23196 & ~n34728;
  assign n23210 = ~n23194 & ~n23209;
  assign n23211 = ~n214 & ~n23210;
  assign n23212 = ~n22319 & ~n22321;
  assign n23213 = ~n22386 & n23212;
  assign n23214 = ~n34611 & ~n23213;
  assign n23215 = ~n22319 & n34611;
  assign n23216 = ~n22321 & n23215;
  assign n23217 = n34611 & n23213;
  assign n23218 = ~n22386 & n23216;
  assign n23219 = ~n23214 & ~n34729;
  assign n23220 = n214 & ~n23194;
  assign n23221 = ~n23209 & n23220;
  assign n23222 = n214 & n23210;
  assign n23223 = ~n23219 & ~n34730;
  assign n23224 = ~n23211 & ~n23223;
  assign n23225 = ~n197 & ~n23224;
  assign n23226 = n197 & ~n23211;
  assign n23227 = ~n23223 & n23226;
  assign n23228 = ~n22336 & ~n34613;
  assign n23229 = ~n22336 & ~n22386;
  assign n23230 = ~n34613 & n23229;
  assign n23231 = ~n22386 & n23228;
  assign n23232 = n22344 & ~n34731;
  assign n23233 = n22348 & n23229;
  assign n23234 = n22344 & ~n34613;
  assign n23235 = ~n22336 & n23234;
  assign n23236 = ~n22386 & n23235;
  assign n23237 = ~n22344 & ~n34731;
  assign n23238 = ~n23236 & ~n23237;
  assign n23239 = ~n23232 & ~n23233;
  assign n23240 = ~n23227 & ~n34732;
  assign n23241 = ~n23225 & ~n23240;
  assign n23242 = ~n22350 & ~n22360;
  assign n23243 = ~n22350 & ~n22386;
  assign n23244 = ~n22360 & n23243;
  assign n23245 = ~n22386 & n23242;
  assign n23246 = n22358 & ~n34733;
  assign n23247 = n22361 & n23243;
  assign n23248 = ~n22350 & n22358;
  assign n23249 = ~n22360 & n23248;
  assign n23250 = ~n22386 & n23249;
  assign n23251 = ~n22358 & ~n34733;
  assign n23252 = ~n23250 & ~n23251;
  assign n23253 = ~n23246 & ~n23247;
  assign n23254 = ~n22362 & ~n22370;
  assign n23255 = ~n22370 & ~n22386;
  assign n23256 = ~n22362 & n23255;
  assign n23257 = ~n22386 & n23254;
  assign n23258 = ~n34617 & ~n34735;
  assign n23259 = ~n34734 & n23258;
  assign n23260 = ~n23241 & n23259;
  assign n23261 = n193 & ~n23260;
  assign n23262 = ~n23225 & n34734;
  assign n23263 = ~n23240 & n23262;
  assign n23264 = n23241 & n34734;
  assign n23265 = n22362 & ~n23255;
  assign n23266 = ~n193 & ~n23254;
  assign n23267 = ~n23265 & n23266;
  assign n23268 = ~n34736 & ~n23267;
  assign n23269 = ~n23261 & n23268;
  assign n23270 = ~n23070 & ~n23072;
  assign n23271 = ~n23269 & n23270;
  assign n23272 = ~n23080 & ~n23271;
  assign n23273 = ~n23072 & n23080;
  assign n23274 = ~n23070 & n23273;
  assign n23275 = n23080 & n23271;
  assign n23276 = ~n23269 & n23274;
  assign n23277 = ~n23272 & ~n34737;
  assign n23278 = ~n23052 & ~n34708;
  assign n23279 = ~n23269 & n23278;
  assign n23280 = ~n34710 & ~n23279;
  assign n23281 = ~n23052 & n34710;
  assign n23282 = ~n34708 & n23281;
  assign n23283 = n34710 & n23279;
  assign n23284 = ~n23269 & n23282;
  assign n23285 = ~n23280 & ~n34738;
  assign n23286 = ~n23035 & ~n23037;
  assign n23287 = ~n23269 & n23286;
  assign n23288 = ~n34707 & ~n23287;
  assign n23289 = ~n23037 & n34707;
  assign n23290 = ~n23035 & n23289;
  assign n23291 = n34707 & n23287;
  assign n23292 = ~n23269 & n23290;
  assign n23293 = ~n23288 & ~n34739;
  assign n23294 = ~n23004 & ~n23006;
  assign n23295 = ~n23269 & n23294;
  assign n23296 = ~n34703 & ~n23295;
  assign n23297 = ~n23006 & n34703;
  assign n23298 = ~n23004 & n23297;
  assign n23299 = n34703 & n23295;
  assign n23300 = ~n23269 & n23298;
  assign n23301 = ~n23296 & ~n34740;
  assign n23302 = ~n22986 & ~n34699;
  assign n23303 = ~n23269 & n23302;
  assign n23304 = ~n34701 & ~n23303;
  assign n23305 = ~n22986 & n34701;
  assign n23306 = ~n34699 & n23305;
  assign n23307 = n34701 & n23303;
  assign n23308 = ~n23269 & n23306;
  assign n23309 = ~n23304 & ~n34741;
  assign n23310 = ~n22969 & ~n22971;
  assign n23311 = ~n23269 & n23310;
  assign n23312 = ~n34698 & ~n23311;
  assign n23313 = ~n22971 & n34698;
  assign n23314 = ~n22969 & n23313;
  assign n23315 = n34698 & n23311;
  assign n23316 = ~n23269 & n23314;
  assign n23317 = ~n23312 & ~n34742;
  assign n23318 = ~n22938 & ~n22940;
  assign n23319 = ~n23269 & n23318;
  assign n23320 = ~n34694 & ~n23319;
  assign n23321 = ~n22940 & n34694;
  assign n23322 = ~n22938 & n23321;
  assign n23323 = n34694 & n23319;
  assign n23324 = ~n23269 & n23322;
  assign n23325 = ~n23320 & ~n34743;
  assign n23326 = ~n22920 & ~n34690;
  assign n23327 = ~n23269 & n23326;
  assign n23328 = ~n34692 & ~n23327;
  assign n23329 = ~n22920 & n34692;
  assign n23330 = ~n34690 & n23329;
  assign n23331 = n34692 & n23327;
  assign n23332 = ~n23269 & n23330;
  assign n23333 = ~n23328 & ~n34744;
  assign n23334 = ~n22903 & ~n22905;
  assign n23335 = ~n23269 & n23334;
  assign n23336 = ~n34689 & ~n23335;
  assign n23337 = ~n22905 & n34689;
  assign n23338 = ~n22903 & n23337;
  assign n23339 = n34689 & n23335;
  assign n23340 = ~n23269 & n23338;
  assign n23341 = ~n23336 & ~n34745;
  assign n23342 = ~n22872 & ~n22874;
  assign n23343 = ~n23269 & n23342;
  assign n23344 = ~n34685 & ~n23343;
  assign n23345 = ~n22874 & n34685;
  assign n23346 = ~n22872 & n23345;
  assign n23347 = n34685 & n23343;
  assign n23348 = ~n23269 & n23346;
  assign n23349 = ~n23344 & ~n34746;
  assign n23350 = ~n22854 & ~n34681;
  assign n23351 = ~n23269 & n23350;
  assign n23352 = ~n34683 & ~n23351;
  assign n23353 = ~n22854 & n34683;
  assign n23354 = ~n34681 & n23353;
  assign n23355 = n34683 & n23351;
  assign n23356 = ~n23269 & n23354;
  assign n23357 = ~n23352 & ~n34747;
  assign n23358 = ~n22837 & ~n22839;
  assign n23359 = ~n23269 & n23358;
  assign n23360 = ~n34680 & ~n23359;
  assign n23361 = ~n22839 & n34680;
  assign n23362 = ~n22837 & n23361;
  assign n23363 = n34680 & n23359;
  assign n23364 = ~n23269 & n23362;
  assign n23365 = ~n23360 & ~n34748;
  assign n23366 = ~n22806 & ~n22808;
  assign n23367 = ~n23269 & n23366;
  assign n23368 = ~n34676 & ~n23367;
  assign n23369 = ~n22808 & n34676;
  assign n23370 = ~n22806 & n23369;
  assign n23371 = n34676 & n23367;
  assign n23372 = ~n23269 & n23370;
  assign n23373 = ~n23368 & ~n34749;
  assign n23374 = ~n22788 & ~n34672;
  assign n23375 = ~n23269 & n23374;
  assign n23376 = ~n34674 & ~n23375;
  assign n23377 = ~n22788 & n34674;
  assign n23378 = ~n34672 & n23377;
  assign n23379 = n34674 & n23375;
  assign n23380 = ~n23269 & n23378;
  assign n23381 = ~n23376 & ~n34750;
  assign n23382 = ~n22771 & ~n22773;
  assign n23383 = ~n23269 & n23382;
  assign n23384 = ~n34671 & ~n23383;
  assign n23385 = ~n22773 & n34671;
  assign n23386 = ~n22771 & n23385;
  assign n23387 = n34671 & n23383;
  assign n23388 = ~n23269 & n23386;
  assign n23389 = ~n23384 & ~n34751;
  assign n23390 = ~n22740 & ~n22742;
  assign n23391 = ~n23269 & n23390;
  assign n23392 = ~n34667 & ~n23391;
  assign n23393 = ~n22742 & n34667;
  assign n23394 = ~n22740 & n23393;
  assign n23395 = n34667 & n23391;
  assign n23396 = ~n23269 & n23394;
  assign n23397 = ~n23392 & ~n34752;
  assign n23398 = ~n22722 & ~n34663;
  assign n23399 = ~n23269 & n23398;
  assign n23400 = ~n34665 & ~n23399;
  assign n23401 = ~n22722 & n34665;
  assign n23402 = ~n34663 & n23401;
  assign n23403 = n34665 & n23399;
  assign n23404 = ~n23269 & n23402;
  assign n23405 = ~n23400 & ~n34753;
  assign n23406 = ~n22705 & ~n22707;
  assign n23407 = ~n23269 & n23406;
  assign n23408 = ~n34662 & ~n23407;
  assign n23409 = ~n22707 & n34662;
  assign n23410 = ~n22705 & n23409;
  assign n23411 = n34662 & n23407;
  assign n23412 = ~n23269 & n23410;
  assign n23413 = ~n23408 & ~n34754;
  assign n23414 = ~n22674 & ~n22676;
  assign n23415 = ~n23269 & n23414;
  assign n23416 = ~n34658 & ~n23415;
  assign n23417 = ~n22676 & n34658;
  assign n23418 = ~n22674 & n23417;
  assign n23419 = n34658 & n23415;
  assign n23420 = ~n23269 & n23418;
  assign n23421 = ~n23416 & ~n34755;
  assign n23422 = ~n22656 & ~n34654;
  assign n23423 = ~n23269 & n23422;
  assign n23424 = ~n34656 & ~n23423;
  assign n23425 = ~n22656 & n34656;
  assign n23426 = ~n34654 & n23425;
  assign n23427 = n34656 & n23423;
  assign n23428 = ~n23269 & n23426;
  assign n23429 = ~n23424 & ~n34756;
  assign n23430 = ~n22639 & ~n22641;
  assign n23431 = ~n23269 & n23430;
  assign n23432 = ~n34653 & ~n23431;
  assign n23433 = ~n22641 & n34653;
  assign n23434 = ~n22639 & n23433;
  assign n23435 = n34653 & n23431;
  assign n23436 = ~n23269 & n23434;
  assign n23437 = ~n23432 & ~n34757;
  assign n23438 = ~n22608 & ~n22610;
  assign n23439 = ~n23269 & n23438;
  assign n23440 = ~n34649 & ~n23439;
  assign n23441 = ~n22610 & n34649;
  assign n23442 = ~n22608 & n23441;
  assign n23443 = n34649 & n23439;
  assign n23444 = ~n23269 & n23442;
  assign n23445 = ~n23440 & ~n34758;
  assign n23446 = ~n22589 & ~n34644;
  assign n23447 = ~n23269 & n23446;
  assign n23448 = ~n34647 & ~n23447;
  assign n23449 = ~n22589 & n34647;
  assign n23450 = ~n34644 & n23449;
  assign n23451 = n34647 & n23447;
  assign n23452 = ~n23269 & n23450;
  assign n23453 = ~n23448 & ~n34759;
  assign n23454 = ~n22572 & ~n22574;
  assign n23455 = ~n23269 & n23454;
  assign n23456 = ~n34643 & ~n23455;
  assign n23457 = ~n22574 & n34643;
  assign n23458 = ~n22572 & n23457;
  assign n23459 = n34643 & n23455;
  assign n23460 = ~n23269 & n23458;
  assign n23461 = ~n23456 & ~n34760;
  assign n23462 = ~n22538 & ~n22540;
  assign n23463 = ~n23269 & n23462;
  assign n23464 = ~n34638 & ~n23463;
  assign n23465 = ~n22540 & n34638;
  assign n23466 = ~n22538 & n23465;
  assign n23467 = n34638 & n23463;
  assign n23468 = ~n23269 & n23466;
  assign n23469 = ~n23464 & ~n34761;
  assign n23470 = ~n22505 & ~n22507;
  assign n23471 = ~n23269 & n23470;
  assign n23472 = ~n34634 & ~n23471;
  assign n23473 = ~n22507 & n34634;
  assign n23474 = ~n22505 & n23473;
  assign n23475 = n34634 & n23471;
  assign n23476 = ~n23269 & n23474;
  assign n23477 = ~n23472 & ~n34762;
  assign n23478 = ~n22472 & ~n22474;
  assign n23479 = ~n23269 & n23478;
  assign n23480 = ~n34630 & ~n23479;
  assign n23481 = ~n22474 & n34630;
  assign n23482 = ~n22472 & n23481;
  assign n23483 = n34630 & n23479;
  assign n23484 = ~n23269 & n23482;
  assign n23485 = ~n23480 & ~n34763;
  assign n23486 = ~n22438 & ~n22440;
  assign n23487 = ~n23269 & n23486;
  assign n23488 = ~n34625 & ~n23487;
  assign n23489 = ~n22440 & n34625;
  assign n23490 = ~n22438 & n23489;
  assign n23491 = n34625 & n23487;
  assign n23492 = ~n23269 & n23490;
  assign n23493 = ~n23488 & ~n34764;
  assign n23494 = ~n22411 & ~n22413;
  assign n23495 = ~n23269 & n23494;
  assign n23496 = ~n22422 & ~n23495;
  assign n23497 = ~n22413 & n22422;
  assign n23498 = ~n22411 & n23497;
  assign n23499 = n22422 & n23495;
  assign n23500 = ~n23269 & n23498;
  assign n23501 = ~n23496 & ~n34765;
  assign n23502 = ~pi18  & ~n23269;
  assign n23503 = ~pi19  & n23502;
  assign n23504 = n22388 & ~n23269;
  assign n23505 = ~n22386 & ~n23267;
  assign n23506 = ~n34736 & n23505;
  assign n23507 = ~n23261 & n23506;
  assign n23508 = ~n34766 & ~n23507;
  assign n23509 = pi20  & ~n23508;
  assign n23510 = ~pi20  & ~n23507;
  assign n23511 = ~pi20  & n23508;
  assign n23512 = ~n34766 & n23510;
  assign n23513 = ~n23509 & ~n34767;
  assign n23514 = pi18  & ~n23269;
  assign n23515 = ~pi16  & ~pi17 ;
  assign n23516 = ~pi18  & n23515;
  assign n23517 = ~n34521 & ~n34619;
  assign n23518 = ~n21591 & n23517;
  assign n23519 = ~n21610 & n23518;
  assign n23520 = ~n34523 & n23519;
  assign n23521 = n21596 & n21612;
  assign n23522 = ~n21604 & n23520;
  assign n23523 = ~n23516 & ~n34768;
  assign n23524 = ~n22384 & n23523;
  assign n23525 = ~n34617 & n23524;
  assign n23526 = ~n22378 & n23525;
  assign n23527 = ~n23514 & ~n23516;
  assign n23528 = n22386 & n23527;
  assign n23529 = ~n23514 & n23526;
  assign n23530 = pi19  & ~n23502;
  assign n23531 = ~n34766 & ~n23530;
  assign n23532 = ~n34769 & n23531;
  assign n23533 = ~n22386 & ~n23527;
  assign n23534 = n21612 & ~n23533;
  assign n23535 = ~n23532 & ~n23533;
  assign n23536 = n21612 & n23535;
  assign n23537 = ~n23532 & n23534;
  assign n23538 = ~n23513 & ~n34770;
  assign n23539 = ~n21612 & ~n23535;
  assign n23540 = n20762 & ~n23539;
  assign n23541 = ~n23538 & n23540;
  assign n23542 = ~n22391 & ~n34620;
  assign n23543 = ~n23269 & n23542;
  assign n23544 = n22396 & ~n23543;
  assign n23545 = ~n22396 & n23542;
  assign n23546 = ~n22396 & n23543;
  assign n23547 = ~n23269 & n23545;
  assign n23548 = ~n23544 & ~n34771;
  assign n23549 = ~n23541 & ~n23548;
  assign n23550 = ~n23538 & ~n23539;
  assign n23551 = ~n20762 & ~n23550;
  assign n23552 = n20011 & ~n23551;
  assign n23553 = ~n23549 & ~n23551;
  assign n23554 = n20011 & n23553;
  assign n23555 = ~n23549 & n23552;
  assign n23556 = ~n23501 & ~n34772;
  assign n23557 = ~n20011 & ~n23553;
  assign n23558 = n19190 & ~n23557;
  assign n23559 = ~n23556 & n23558;
  assign n23560 = ~n22425 & ~n34622;
  assign n23561 = ~n23269 & n23560;
  assign n23562 = ~n22435 & ~n23561;
  assign n23563 = ~n22425 & n22435;
  assign n23564 = ~n34622 & n23563;
  assign n23565 = n22435 & n23561;
  assign n23566 = ~n23269 & n23564;
  assign n23567 = n22435 & ~n23561;
  assign n23568 = ~n22435 & n23561;
  assign n23569 = ~n23567 & ~n23568;
  assign n23570 = ~n23562 & ~n34773;
  assign n23571 = ~n23559 & n34774;
  assign n23572 = ~n23556 & ~n23557;
  assign n23573 = ~n19190 & ~n23572;
  assign n23574 = n18472 & ~n23573;
  assign n23575 = ~n23571 & ~n23573;
  assign n23576 = n18472 & n23575;
  assign n23577 = ~n23571 & n23574;
  assign n23578 = ~n23493 & ~n34775;
  assign n23579 = ~n18472 & ~n23575;
  assign n23580 = n17690 & ~n23579;
  assign n23581 = ~n23578 & n23580;
  assign n23582 = ~n22455 & ~n34626;
  assign n23583 = ~n23269 & n23582;
  assign n23584 = ~n34628 & ~n23583;
  assign n23585 = n34628 & n23583;
  assign n23586 = ~n22455 & ~n34628;
  assign n23587 = ~n34626 & n23586;
  assign n23588 = ~n23269 & n23587;
  assign n23589 = n34628 & ~n23583;
  assign n23590 = ~n23588 & ~n23589;
  assign n23591 = ~n23584 & ~n23585;
  assign n23592 = ~n23581 & ~n34776;
  assign n23593 = ~n23578 & ~n23579;
  assign n23594 = ~n17690 & ~n23593;
  assign n23595 = n17001 & ~n23594;
  assign n23596 = ~n23592 & ~n23594;
  assign n23597 = n17001 & n23596;
  assign n23598 = ~n23592 & n23595;
  assign n23599 = ~n23485 & ~n34777;
  assign n23600 = ~n17001 & ~n23596;
  assign n23601 = n16248 & ~n23600;
  assign n23602 = ~n23599 & n23601;
  assign n23603 = ~n22489 & ~n34631;
  assign n23604 = ~n23269 & n23603;
  assign n23605 = ~n34632 & n23604;
  assign n23606 = n34632 & ~n23604;
  assign n23607 = ~n22489 & n34632;
  assign n23608 = ~n34631 & n23607;
  assign n23609 = ~n23269 & n23608;
  assign n23610 = ~n34632 & ~n23604;
  assign n23611 = ~n23609 & ~n23610;
  assign n23612 = ~n23605 & ~n23606;
  assign n23613 = ~n23602 & ~n34778;
  assign n23614 = ~n23599 & ~n23600;
  assign n23615 = ~n16248 & ~n23614;
  assign n23616 = n15586 & ~n23615;
  assign n23617 = ~n23613 & ~n23615;
  assign n23618 = n15586 & n23617;
  assign n23619 = ~n23613 & n23616;
  assign n23620 = ~n23477 & ~n34779;
  assign n23621 = ~n15586 & ~n23617;
  assign n23622 = n14866 & ~n23621;
  assign n23623 = ~n23620 & n23622;
  assign n23624 = ~n22522 & ~n34635;
  assign n23625 = ~n23269 & n23624;
  assign n23626 = ~n34636 & n23625;
  assign n23627 = n34636 & ~n23625;
  assign n23628 = ~n34636 & ~n23625;
  assign n23629 = ~n22522 & n34636;
  assign n23630 = ~n34635 & n23629;
  assign n23631 = n34636 & n23625;
  assign n23632 = ~n23269 & n23630;
  assign n23633 = ~n23628 & ~n34780;
  assign n23634 = ~n23626 & ~n23627;
  assign n23635 = ~n23623 & ~n34781;
  assign n23636 = ~n23620 & ~n23621;
  assign n23637 = ~n14866 & ~n23636;
  assign n23638 = n14233 & ~n23637;
  assign n23639 = ~n23635 & ~n23637;
  assign n23640 = n14233 & n23639;
  assign n23641 = ~n23635 & n23638;
  assign n23642 = ~n23469 & ~n34782;
  assign n23643 = ~n14233 & ~n23639;
  assign n23644 = n13548 & ~n23643;
  assign n23645 = ~n23642 & n23644;
  assign n23646 = ~n22555 & ~n34639;
  assign n23647 = ~n22555 & ~n23269;
  assign n23648 = ~n34639 & n23647;
  assign n23649 = ~n23269 & n23646;
  assign n23650 = n34641 & ~n34783;
  assign n23651 = n22570 & n23647;
  assign n23652 = ~n34641 & n34783;
  assign n23653 = ~n22555 & n34641;
  assign n23654 = ~n34639 & n23653;
  assign n23655 = ~n23269 & n23654;
  assign n23656 = ~n34641 & ~n34783;
  assign n23657 = ~n23655 & ~n23656;
  assign n23658 = ~n23650 & ~n34784;
  assign n23659 = ~n23645 & ~n34785;
  assign n23660 = ~n23642 & ~n23643;
  assign n23661 = ~n13548 & ~n23660;
  assign n23662 = n12948 & ~n23661;
  assign n23663 = ~n23659 & ~n23661;
  assign n23664 = n12948 & n23663;
  assign n23665 = ~n23659 & n23662;
  assign n23666 = ~n23461 & ~n34786;
  assign n23667 = ~n12948 & ~n23663;
  assign n23668 = n12296 & ~n23667;
  assign n23669 = ~n23666 & n23668;
  assign n23670 = ~n23453 & ~n23669;
  assign n23671 = ~n23666 & ~n23667;
  assign n23672 = ~n12296 & ~n23671;
  assign n23673 = n11719 & ~n23672;
  assign n23674 = ~n23670 & ~n23672;
  assign n23675 = n11719 & n23674;
  assign n23676 = ~n23670 & n23673;
  assign n23677 = ~n23445 & ~n34787;
  assign n23678 = ~n11719 & ~n23674;
  assign n23679 = n11097 & ~n23678;
  assign n23680 = ~n23677 & n23679;
  assign n23681 = ~n22625 & ~n34651;
  assign n23682 = ~n22625 & ~n23269;
  assign n23683 = ~n34651 & n23682;
  assign n23684 = ~n23269 & n23681;
  assign n23685 = n22633 & ~n34788;
  assign n23686 = n22637 & n23682;
  assign n23687 = ~n22625 & n22633;
  assign n23688 = ~n34651 & n23687;
  assign n23689 = ~n23269 & n23688;
  assign n23690 = ~n22633 & ~n34788;
  assign n23691 = ~n23689 & ~n23690;
  assign n23692 = ~n23685 & ~n23686;
  assign n23693 = ~n23680 & ~n34789;
  assign n23694 = ~n23677 & ~n23678;
  assign n23695 = ~n11097 & ~n23694;
  assign n23696 = n10555 & ~n23695;
  assign n23697 = ~n23693 & ~n23695;
  assign n23698 = n10555 & n23697;
  assign n23699 = ~n23693 & n23696;
  assign n23700 = ~n23437 & ~n34790;
  assign n23701 = ~n10555 & ~n23697;
  assign n23702 = n9969 & ~n23701;
  assign n23703 = ~n23700 & n23702;
  assign n23704 = ~n23429 & ~n23703;
  assign n23705 = ~n23700 & ~n23701;
  assign n23706 = ~n9969 & ~n23705;
  assign n23707 = n9457 & ~n23706;
  assign n23708 = ~n23704 & ~n23706;
  assign n23709 = n9457 & n23708;
  assign n23710 = ~n23704 & n23707;
  assign n23711 = ~n23421 & ~n34791;
  assign n23712 = ~n9457 & ~n23708;
  assign n23713 = n8896 & ~n23712;
  assign n23714 = ~n23711 & n23713;
  assign n23715 = ~n22691 & ~n34660;
  assign n23716 = ~n22691 & ~n23269;
  assign n23717 = ~n34660 & n23716;
  assign n23718 = ~n23269 & n23715;
  assign n23719 = n22699 & ~n34792;
  assign n23720 = n22703 & n23716;
  assign n23721 = ~n22691 & n22699;
  assign n23722 = ~n34660 & n23721;
  assign n23723 = ~n23269 & n23722;
  assign n23724 = ~n22699 & ~n34792;
  assign n23725 = ~n23723 & ~n23724;
  assign n23726 = ~n23719 & ~n23720;
  assign n23727 = ~n23714 & ~n34793;
  assign n23728 = ~n23711 & ~n23712;
  assign n23729 = ~n8896 & ~n23728;
  assign n23730 = n8411 & ~n23729;
  assign n23731 = ~n23727 & ~n23729;
  assign n23732 = n8411 & n23731;
  assign n23733 = ~n23727 & n23730;
  assign n23734 = ~n23413 & ~n34794;
  assign n23735 = ~n8411 & ~n23731;
  assign n23736 = n7885 & ~n23735;
  assign n23737 = ~n23734 & n23736;
  assign n23738 = ~n23405 & ~n23737;
  assign n23739 = ~n23734 & ~n23735;
  assign n23740 = ~n7885 & ~n23739;
  assign n23741 = n7428 & ~n23740;
  assign n23742 = ~n23738 & ~n23740;
  assign n23743 = n7428 & n23742;
  assign n23744 = ~n23738 & n23741;
  assign n23745 = ~n23397 & ~n34795;
  assign n23746 = ~n7428 & ~n23742;
  assign n23747 = n6937 & ~n23746;
  assign n23748 = ~n23745 & n23747;
  assign n23749 = ~n22757 & ~n34669;
  assign n23750 = ~n22757 & ~n23269;
  assign n23751 = ~n34669 & n23750;
  assign n23752 = ~n23269 & n23749;
  assign n23753 = n22765 & ~n34796;
  assign n23754 = n22769 & n23750;
  assign n23755 = ~n22757 & n22765;
  assign n23756 = ~n34669 & n23755;
  assign n23757 = ~n23269 & n23756;
  assign n23758 = ~n22765 & ~n34796;
  assign n23759 = ~n23757 & ~n23758;
  assign n23760 = ~n23753 & ~n23754;
  assign n23761 = ~n23748 & ~n34797;
  assign n23762 = ~n23745 & ~n23746;
  assign n23763 = ~n6937 & ~n23762;
  assign n23764 = n6507 & ~n23763;
  assign n23765 = ~n23761 & ~n23763;
  assign n23766 = n6507 & n23765;
  assign n23767 = ~n23761 & n23764;
  assign n23768 = ~n23389 & ~n34798;
  assign n23769 = ~n6507 & ~n23765;
  assign n23770 = n6051 & ~n23769;
  assign n23771 = ~n23768 & n23770;
  assign n23772 = ~n23381 & ~n23771;
  assign n23773 = ~n23768 & ~n23769;
  assign n23774 = ~n6051 & ~n23773;
  assign n23775 = n5648 & ~n23774;
  assign n23776 = ~n23772 & ~n23774;
  assign n23777 = n5648 & n23776;
  assign n23778 = ~n23772 & n23775;
  assign n23779 = ~n23373 & ~n34799;
  assign n23780 = ~n5648 & ~n23776;
  assign n23781 = n5223 & ~n23780;
  assign n23782 = ~n23779 & n23781;
  assign n23783 = ~n22823 & ~n34678;
  assign n23784 = ~n22823 & ~n23269;
  assign n23785 = ~n34678 & n23784;
  assign n23786 = ~n23269 & n23783;
  assign n23787 = n22831 & ~n34800;
  assign n23788 = n22835 & n23784;
  assign n23789 = ~n22823 & n22831;
  assign n23790 = ~n34678 & n23789;
  assign n23791 = ~n23269 & n23790;
  assign n23792 = ~n22831 & ~n34800;
  assign n23793 = ~n23791 & ~n23792;
  assign n23794 = ~n23787 & ~n23788;
  assign n23795 = ~n23782 & ~n34801;
  assign n23796 = ~n23779 & ~n23780;
  assign n23797 = ~n5223 & ~n23796;
  assign n23798 = n4851 & ~n23797;
  assign n23799 = ~n23795 & ~n23797;
  assign n23800 = n4851 & n23799;
  assign n23801 = ~n23795 & n23798;
  assign n23802 = ~n23365 & ~n34802;
  assign n23803 = ~n4851 & ~n23799;
  assign n23804 = n4461 & ~n23803;
  assign n23805 = ~n23802 & n23804;
  assign n23806 = ~n23357 & ~n23805;
  assign n23807 = ~n23802 & ~n23803;
  assign n23808 = ~n4461 & ~n23807;
  assign n23809 = n4115 & ~n23808;
  assign n23810 = ~n23806 & ~n23808;
  assign n23811 = n4115 & n23810;
  assign n23812 = ~n23806 & n23809;
  assign n23813 = ~n23349 & ~n34803;
  assign n23814 = ~n4115 & ~n23810;
  assign n23815 = n3754 & ~n23814;
  assign n23816 = ~n23813 & n23815;
  assign n23817 = ~n22889 & ~n34687;
  assign n23818 = ~n22889 & ~n23269;
  assign n23819 = ~n34687 & n23818;
  assign n23820 = ~n23269 & n23817;
  assign n23821 = n22897 & ~n34804;
  assign n23822 = n22901 & n23818;
  assign n23823 = ~n22889 & n22897;
  assign n23824 = ~n34687 & n23823;
  assign n23825 = ~n23269 & n23824;
  assign n23826 = ~n22897 & ~n34804;
  assign n23827 = ~n23825 & ~n23826;
  assign n23828 = ~n23821 & ~n23822;
  assign n23829 = ~n23816 & ~n34805;
  assign n23830 = ~n23813 & ~n23814;
  assign n23831 = ~n3754 & ~n23830;
  assign n23832 = n3444 & ~n23831;
  assign n23833 = ~n23829 & ~n23831;
  assign n23834 = n3444 & n23833;
  assign n23835 = ~n23829 & n23832;
  assign n23836 = ~n23341 & ~n34806;
  assign n23837 = ~n3444 & ~n23833;
  assign n23838 = n3116 & ~n23837;
  assign n23839 = ~n23836 & n23838;
  assign n23840 = ~n23333 & ~n23839;
  assign n23841 = ~n23836 & ~n23837;
  assign n23842 = ~n3116 & ~n23841;
  assign n23843 = n2833 & ~n23842;
  assign n23844 = ~n23840 & ~n23842;
  assign n23845 = n2833 & n23844;
  assign n23846 = ~n23840 & n23843;
  assign n23847 = ~n23325 & ~n34807;
  assign n23848 = ~n2833 & ~n23844;
  assign n23849 = n2536 & ~n23848;
  assign n23850 = ~n23847 & n23849;
  assign n23851 = ~n22955 & ~n34696;
  assign n23852 = ~n22955 & ~n23269;
  assign n23853 = ~n34696 & n23852;
  assign n23854 = ~n23269 & n23851;
  assign n23855 = n22963 & ~n34808;
  assign n23856 = n22967 & n23852;
  assign n23857 = ~n22955 & n22963;
  assign n23858 = ~n34696 & n23857;
  assign n23859 = ~n23269 & n23858;
  assign n23860 = ~n22963 & ~n34808;
  assign n23861 = ~n23859 & ~n23860;
  assign n23862 = ~n23855 & ~n23856;
  assign n23863 = ~n23850 & ~n34809;
  assign n23864 = ~n23847 & ~n23848;
  assign n23865 = ~n2536 & ~n23864;
  assign n23866 = n2283 & ~n23865;
  assign n23867 = ~n23863 & ~n23865;
  assign n23868 = n2283 & n23867;
  assign n23869 = ~n23863 & n23866;
  assign n23870 = ~n23317 & ~n34810;
  assign n23871 = ~n2283 & ~n23867;
  assign n23872 = n2021 & ~n23871;
  assign n23873 = ~n23870 & n23872;
  assign n23874 = ~n23309 & ~n23873;
  assign n23875 = ~n23870 & ~n23871;
  assign n23876 = ~n2021 & ~n23875;
  assign n23877 = n1796 & ~n23876;
  assign n23878 = ~n23874 & ~n23876;
  assign n23879 = n1796 & n23878;
  assign n23880 = ~n23874 & n23877;
  assign n23881 = ~n23301 & ~n34811;
  assign n23882 = ~n1796 & ~n23878;
  assign n23883 = n1567 & ~n23882;
  assign n23884 = ~n23881 & n23883;
  assign n23885 = ~n23021 & ~n34705;
  assign n23886 = ~n23021 & ~n23269;
  assign n23887 = ~n34705 & n23886;
  assign n23888 = ~n23269 & n23885;
  assign n23889 = n23029 & ~n34812;
  assign n23890 = n23033 & n23886;
  assign n23891 = ~n23021 & n23029;
  assign n23892 = ~n34705 & n23891;
  assign n23893 = ~n23269 & n23892;
  assign n23894 = ~n23029 & ~n34812;
  assign n23895 = ~n23893 & ~n23894;
  assign n23896 = ~n23889 & ~n23890;
  assign n23897 = ~n23884 & ~n34813;
  assign n23898 = ~n23881 & ~n23882;
  assign n23899 = ~n1567 & ~n23898;
  assign n23900 = n1374 & ~n23899;
  assign n23901 = ~n23897 & ~n23899;
  assign n23902 = n1374 & n23901;
  assign n23903 = ~n23897 & n23900;
  assign n23904 = ~n23293 & ~n34814;
  assign n23905 = ~n1374 & ~n23901;
  assign n23906 = n1179 & ~n23905;
  assign n23907 = ~n23904 & n23906;
  assign n23908 = ~n23285 & ~n23907;
  assign n23909 = ~n23904 & ~n23905;
  assign n23910 = ~n1179 & ~n23909;
  assign n23911 = n1016 & ~n23910;
  assign n23912 = ~n23908 & ~n23910;
  assign n23913 = n1016 & n23912;
  assign n23914 = ~n23908 & n23911;
  assign n23915 = ~n23277 & ~n34815;
  assign n23916 = ~n1016 & ~n23912;
  assign n23917 = ~n23915 & ~n23916;
  assign n23918 = ~n855 & ~n23917;
  assign n23919 = ~n23083 & ~n34713;
  assign n23920 = ~n23269 & n23919;
  assign n23921 = n23091 & ~n23920;
  assign n23922 = ~n23091 & n23920;
  assign n23923 = ~n23083 & n23091;
  assign n23924 = ~n34713 & n23923;
  assign n23925 = ~n23269 & n23924;
  assign n23926 = ~n23091 & ~n23920;
  assign n23927 = ~n23925 & ~n23926;
  assign n23928 = ~n23921 & ~n23922;
  assign n23929 = n855 & ~n23916;
  assign n23930 = ~n23915 & n23929;
  assign n23931 = ~n34816 & ~n23930;
  assign n23932 = ~n23918 & ~n23931;
  assign n23933 = ~n720 & ~n23932;
  assign n23934 = ~n23097 & ~n23099;
  assign n23935 = ~n23269 & n23934;
  assign n23936 = ~n34715 & ~n23935;
  assign n23937 = ~n23099 & n34715;
  assign n23938 = ~n23097 & n23937;
  assign n23939 = n34715 & n23935;
  assign n23940 = ~n23269 & n23938;
  assign n23941 = ~n23936 & ~n34817;
  assign n23942 = n720 & ~n23918;
  assign n23943 = n720 & n23932;
  assign n23944 = ~n23931 & n23942;
  assign n23945 = ~n23941 & ~n34818;
  assign n23946 = ~n23933 & ~n23945;
  assign n23947 = ~n592 & ~n23946;
  assign n23948 = n592 & ~n23933;
  assign n23949 = ~n23945 & n23948;
  assign n23950 = ~n23114 & ~n34717;
  assign n23951 = ~n23114 & ~n23269;
  assign n23952 = ~n34717 & n23951;
  assign n23953 = ~n23269 & n23950;
  assign n23954 = n23122 & ~n34819;
  assign n23955 = n23126 & n23951;
  assign n23956 = ~n23114 & n23122;
  assign n23957 = ~n34717 & n23956;
  assign n23958 = ~n23269 & n23957;
  assign n23959 = ~n23122 & ~n34819;
  assign n23960 = ~n23958 & ~n23959;
  assign n23961 = ~n23954 & ~n23955;
  assign n23962 = ~n23949 & ~n34820;
  assign n23963 = ~n23947 & ~n23962;
  assign n23964 = ~n487 & ~n23963;
  assign n23965 = ~n23128 & ~n23130;
  assign n23966 = ~n23269 & n23965;
  assign n23967 = ~n34719 & ~n23966;
  assign n23968 = ~n23130 & n34719;
  assign n23969 = ~n23128 & n23968;
  assign n23970 = n34719 & n23966;
  assign n23971 = ~n23269 & n23969;
  assign n23972 = ~n23967 & ~n34821;
  assign n23973 = n487 & ~n23947;
  assign n23974 = n487 & n23963;
  assign n23975 = ~n23962 & n23973;
  assign n23976 = ~n23972 & ~n34822;
  assign n23977 = ~n23964 & ~n23976;
  assign n23978 = ~n393 & ~n23977;
  assign n23979 = n393 & ~n23964;
  assign n23980 = ~n23976 & n23979;
  assign n23981 = ~n23145 & ~n34721;
  assign n23982 = ~n23145 & ~n23269;
  assign n23983 = ~n34721 & n23982;
  assign n23984 = ~n23269 & n23981;
  assign n23985 = n23153 & ~n34823;
  assign n23986 = n23157 & n23982;
  assign n23987 = ~n23145 & n23153;
  assign n23988 = ~n34721 & n23987;
  assign n23989 = ~n23269 & n23988;
  assign n23990 = ~n23153 & ~n34823;
  assign n23991 = ~n23989 & ~n23990;
  assign n23992 = ~n23985 & ~n23986;
  assign n23993 = ~n23980 & ~n34824;
  assign n23994 = ~n23978 & ~n23993;
  assign n23995 = ~n321 & ~n23994;
  assign n23996 = ~n23159 & ~n23161;
  assign n23997 = ~n23269 & n23996;
  assign n23998 = ~n34723 & ~n23997;
  assign n23999 = ~n23161 & n34723;
  assign n24000 = ~n23159 & n23999;
  assign n24001 = n34723 & n23997;
  assign n24002 = ~n23269 & n24000;
  assign n24003 = ~n23998 & ~n34825;
  assign n24004 = n321 & ~n23978;
  assign n24005 = n321 & n23994;
  assign n24006 = ~n23993 & n24004;
  assign n24007 = ~n24003 & ~n34826;
  assign n24008 = ~n23995 & ~n24007;
  assign n24009 = ~n263 & ~n24008;
  assign n24010 = ~n23176 & ~n34724;
  assign n24011 = ~n23269 & n24010;
  assign n24012 = ~n34726 & ~n24011;
  assign n24013 = ~n23176 & n34726;
  assign n24014 = ~n34724 & n24013;
  assign n24015 = n34726 & n24011;
  assign n24016 = ~n23269 & n24014;
  assign n24017 = ~n24012 & ~n34827;
  assign n24018 = n263 & ~n23995;
  assign n24019 = ~n24007 & n24018;
  assign n24020 = ~n24017 & ~n24019;
  assign n24021 = ~n24009 & ~n24020;
  assign n24022 = ~n214 & ~n24021;
  assign n24023 = ~n23194 & ~n23196;
  assign n24024 = ~n23269 & n24023;
  assign n24025 = ~n34728 & ~n24024;
  assign n24026 = ~n23196 & n34728;
  assign n24027 = ~n23194 & n24026;
  assign n24028 = n34728 & n24024;
  assign n24029 = ~n23269 & n24027;
  assign n24030 = ~n24025 & ~n34828;
  assign n24031 = n214 & ~n24009;
  assign n24032 = n214 & n24021;
  assign n24033 = ~n24020 & n24031;
  assign n24034 = ~n24030 & ~n34829;
  assign n24035 = ~n24022 & ~n24034;
  assign n24036 = ~n197 & ~n24035;
  assign n24037 = n197 & ~n24022;
  assign n24038 = ~n24034 & n24037;
  assign n24039 = ~n23211 & ~n34730;
  assign n24040 = ~n23211 & ~n23269;
  assign n24041 = ~n34730 & n24040;
  assign n24042 = ~n23269 & n24039;
  assign n24043 = n23219 & ~n34830;
  assign n24044 = n23223 & n24040;
  assign n24045 = ~n23211 & n23219;
  assign n24046 = ~n34730 & n24045;
  assign n24047 = ~n23269 & n24046;
  assign n24048 = ~n23219 & ~n34830;
  assign n24049 = ~n24047 & ~n24048;
  assign n24050 = ~n24043 & ~n24044;
  assign n24051 = ~n24038 & ~n34831;
  assign n24052 = ~n24036 & ~n24051;
  assign n24053 = ~n23225 & ~n23227;
  assign n24054 = ~n23269 & n24053;
  assign n24055 = ~n34732 & ~n24054;
  assign n24056 = ~n23227 & n34732;
  assign n24057 = ~n23225 & n24056;
  assign n24058 = n34732 & n24054;
  assign n24059 = ~n23269 & n24057;
  assign n24060 = ~n24055 & ~n34832;
  assign n24061 = ~n23241 & ~n34734;
  assign n24062 = ~n34734 & ~n23269;
  assign n24063 = ~n23241 & n24062;
  assign n24064 = ~n23269 & n24061;
  assign n24065 = ~n34736 & ~n34833;
  assign n24066 = ~n24060 & n24065;
  assign n24067 = ~n24052 & n24066;
  assign n24068 = n193 & ~n24067;
  assign n24069 = ~n24036 & n24060;
  assign n24070 = n24052 & n24060;
  assign n24071 = ~n24051 & n24069;
  assign n24072 = n23241 & ~n24062;
  assign n24073 = ~n193 & ~n24061;
  assign n24074 = ~n24072 & n24073;
  assign n24075 = ~n34834 & ~n24074;
  assign n24076 = ~n24068 & n24075;
  assign n24077 = pi16  & ~n24076;
  assign n24078 = ~pi14  & ~pi15 ;
  assign n24079 = ~pi16  & n24078;
  assign n24080 = ~n24077 & ~n24079;
  assign n24081 = ~n23269 & ~n24080;
  assign n24082 = ~pi16  & ~n24076;
  assign n24083 = pi17  & ~n24082;
  assign n24084 = ~pi17  & n24082;
  assign n24085 = n23515 & ~n24076;
  assign n24086 = ~n24083 & ~n34835;
  assign n24087 = ~n34615 & ~n34768;
  assign n24088 = ~n22365 & n24087;
  assign n24089 = ~n22384 & n24088;
  assign n24090 = ~n34617 & n24089;
  assign n24091 = n22370 & n22386;
  assign n24092 = ~n22378 & n24090;
  assign n24093 = ~n24079 & ~n34836;
  assign n24094 = ~n23267 & n24093;
  assign n24095 = ~n34736 & n24094;
  assign n24096 = ~n23261 & n24095;
  assign n24097 = n23269 & n24080;
  assign n24098 = ~n24077 & n24096;
  assign n24099 = n24086 & ~n34837;
  assign n24100 = ~n24081 & ~n24099;
  assign n24101 = ~n22386 & ~n24100;
  assign n24102 = n22386 & ~n24081;
  assign n24103 = ~n24099 & n24102;
  assign n24104 = ~n23269 & ~n24074;
  assign n24105 = ~n34834 & n24104;
  assign n24106 = ~n24068 & n24105;
  assign n24107 = ~n34835 & ~n24106;
  assign n24108 = pi18  & ~n24107;
  assign n24109 = ~pi18  & ~n24106;
  assign n24110 = ~pi18  & n24107;
  assign n24111 = ~n34835 & n24109;
  assign n24112 = ~n24108 & ~n34838;
  assign n24113 = ~n24103 & ~n24112;
  assign n24114 = ~n24101 & ~n24113;
  assign n24115 = ~n21612 & ~n24114;
  assign n24116 = n21612 & ~n24101;
  assign n24117 = ~n24113 & n24116;
  assign n24118 = n21612 & n24114;
  assign n24119 = ~n34769 & ~n23533;
  assign n24120 = ~n24076 & n24119;
  assign n24121 = n23531 & ~n24120;
  assign n24122 = ~n23531 & n24119;
  assign n24123 = ~n23531 & n24120;
  assign n24124 = ~n24076 & n24122;
  assign n24125 = ~n24121 & ~n34840;
  assign n24126 = ~n34839 & ~n24125;
  assign n24127 = ~n24115 & ~n24126;
  assign n24128 = ~n20762 & ~n24127;
  assign n24129 = n20762 & ~n24115;
  assign n24130 = ~n24126 & n24129;
  assign n24131 = ~n34770 & ~n23539;
  assign n24132 = ~n23539 & ~n24076;
  assign n24133 = ~n34770 & n24132;
  assign n24134 = ~n24076 & n24131;
  assign n24135 = n23513 & ~n34841;
  assign n24136 = n23538 & n24132;
  assign n24137 = n23513 & ~n34770;
  assign n24138 = ~n23539 & n24137;
  assign n24139 = ~n24076 & n24138;
  assign n24140 = ~n23513 & ~n34841;
  assign n24141 = ~n24139 & ~n24140;
  assign n24142 = ~n24135 & ~n24136;
  assign n24143 = ~n24130 & ~n34842;
  assign n24144 = ~n24128 & ~n24143;
  assign n24145 = ~n20011 & ~n24144;
  assign n24146 = n20011 & ~n24128;
  assign n24147 = ~n24143 & n24146;
  assign n24148 = n20011 & n24144;
  assign n24149 = ~n23541 & ~n23551;
  assign n24150 = ~n24076 & n24149;
  assign n24151 = ~n23548 & ~n24150;
  assign n24152 = n23548 & ~n23551;
  assign n24153 = ~n23541 & n24152;
  assign n24154 = n23548 & n24150;
  assign n24155 = ~n24076 & n24153;
  assign n24156 = n23548 & ~n24150;
  assign n24157 = ~n23548 & n24150;
  assign n24158 = ~n24156 & ~n24157;
  assign n24159 = ~n24151 & ~n34844;
  assign n24160 = ~n34843 & n34845;
  assign n24161 = ~n24145 & ~n24160;
  assign n24162 = ~n19190 & ~n24161;
  assign n24163 = n19190 & ~n24145;
  assign n24164 = ~n24160 & n24163;
  assign n24165 = ~n34772 & ~n23557;
  assign n24166 = ~n23557 & ~n24076;
  assign n24167 = ~n34772 & n24166;
  assign n24168 = ~n24076 & n24165;
  assign n24169 = n23501 & ~n34846;
  assign n24170 = n23556 & n24166;
  assign n24171 = n23501 & ~n34772;
  assign n24172 = ~n23557 & n24171;
  assign n24173 = ~n24076 & n24172;
  assign n24174 = ~n23501 & ~n34846;
  assign n24175 = ~n24173 & ~n24174;
  assign n24176 = ~n24169 & ~n24170;
  assign n24177 = ~n24164 & ~n34847;
  assign n24178 = ~n24162 & ~n24177;
  assign n24179 = ~n18472 & ~n24178;
  assign n24180 = n18472 & ~n24162;
  assign n24181 = ~n24177 & n24180;
  assign n24182 = n18472 & n24178;
  assign n24183 = ~n23559 & ~n23573;
  assign n24184 = ~n24076 & n24183;
  assign n24185 = ~n34774 & ~n24184;
  assign n24186 = n34774 & n24184;
  assign n24187 = ~n34774 & ~n23573;
  assign n24188 = ~n23559 & n24187;
  assign n24189 = ~n24076 & n24188;
  assign n24190 = n34774 & ~n24184;
  assign n24191 = ~n24189 & ~n24190;
  assign n24192 = ~n24185 & ~n24186;
  assign n24193 = ~n34848 & ~n34849;
  assign n24194 = ~n24179 & ~n24193;
  assign n24195 = ~n17690 & ~n24194;
  assign n24196 = n17690 & ~n24179;
  assign n24197 = ~n24193 & n24196;
  assign n24198 = ~n34775 & ~n23579;
  assign n24199 = ~n23579 & ~n24076;
  assign n24200 = ~n34775 & n24199;
  assign n24201 = ~n24076 & n24198;
  assign n24202 = n23493 & ~n34850;
  assign n24203 = n23578 & n24199;
  assign n24204 = n23493 & ~n34775;
  assign n24205 = ~n23579 & n24204;
  assign n24206 = ~n24076 & n24205;
  assign n24207 = ~n23493 & ~n34850;
  assign n24208 = ~n24206 & ~n24207;
  assign n24209 = ~n24202 & ~n24203;
  assign n24210 = ~n24197 & ~n34851;
  assign n24211 = ~n24195 & ~n24210;
  assign n24212 = ~n17001 & ~n24211;
  assign n24213 = n17001 & ~n24195;
  assign n24214 = ~n24210 & n24213;
  assign n24215 = n17001 & n24211;
  assign n24216 = ~n23581 & ~n23594;
  assign n24217 = ~n24076 & n24216;
  assign n24218 = ~n34776 & n24217;
  assign n24219 = n34776 & ~n24217;
  assign n24220 = n34776 & ~n23594;
  assign n24221 = ~n23581 & n24220;
  assign n24222 = ~n24076 & n24221;
  assign n24223 = ~n34776 & ~n24217;
  assign n24224 = ~n24222 & ~n24223;
  assign n24225 = ~n24218 & ~n24219;
  assign n24226 = ~n34852 & ~n34853;
  assign n24227 = ~n24212 & ~n24226;
  assign n24228 = ~n16248 & ~n24227;
  assign n24229 = n16248 & ~n24212;
  assign n24230 = ~n24226 & n24229;
  assign n24231 = ~n34777 & ~n23600;
  assign n24232 = ~n23600 & ~n24076;
  assign n24233 = ~n34777 & n24232;
  assign n24234 = ~n24076 & n24231;
  assign n24235 = n23485 & ~n34854;
  assign n24236 = n23599 & n24232;
  assign n24237 = n23485 & ~n34777;
  assign n24238 = ~n23600 & n24237;
  assign n24239 = ~n24076 & n24238;
  assign n24240 = ~n23485 & ~n34854;
  assign n24241 = ~n24239 & ~n24240;
  assign n24242 = ~n24235 & ~n24236;
  assign n24243 = ~n24230 & ~n34855;
  assign n24244 = ~n24228 & ~n24243;
  assign n24245 = ~n15586 & ~n24244;
  assign n24246 = n15586 & ~n24228;
  assign n24247 = ~n24243 & n24246;
  assign n24248 = n15586 & n24244;
  assign n24249 = ~n23602 & ~n23615;
  assign n24250 = ~n24076 & n24249;
  assign n24251 = ~n34778 & n24250;
  assign n24252 = n34778 & ~n24250;
  assign n24253 = ~n34778 & ~n24250;
  assign n24254 = n34778 & ~n23615;
  assign n24255 = ~n23602 & n24254;
  assign n24256 = n34778 & n24250;
  assign n24257 = ~n24076 & n24255;
  assign n24258 = ~n24253 & ~n34857;
  assign n24259 = ~n24251 & ~n24252;
  assign n24260 = ~n34856 & ~n34858;
  assign n24261 = ~n24245 & ~n24260;
  assign n24262 = ~n14866 & ~n24261;
  assign n24263 = n14866 & ~n24245;
  assign n24264 = ~n24260 & n24263;
  assign n24265 = ~n34779 & ~n23621;
  assign n24266 = ~n23621 & ~n24076;
  assign n24267 = ~n34779 & n24266;
  assign n24268 = ~n24076 & n24265;
  assign n24269 = n23477 & ~n34859;
  assign n24270 = n23620 & n24266;
  assign n24271 = n23477 & ~n34779;
  assign n24272 = ~n23621 & n24271;
  assign n24273 = ~n24076 & n24272;
  assign n24274 = ~n23477 & ~n34859;
  assign n24275 = ~n24273 & ~n24274;
  assign n24276 = ~n24269 & ~n24270;
  assign n24277 = ~n24264 & ~n34860;
  assign n24278 = ~n24262 & ~n24277;
  assign n24279 = ~n14233 & ~n24278;
  assign n24280 = n14233 & ~n24262;
  assign n24281 = ~n24277 & n24280;
  assign n24282 = n14233 & n24278;
  assign n24283 = ~n23623 & ~n23637;
  assign n24284 = ~n23637 & ~n24076;
  assign n24285 = ~n23623 & n24284;
  assign n24286 = ~n24076 & n24283;
  assign n24287 = n34781 & ~n34862;
  assign n24288 = n23635 & n24284;
  assign n24289 = ~n34781 & n34862;
  assign n24290 = n34781 & ~n23637;
  assign n24291 = ~n23623 & n24290;
  assign n24292 = ~n24076 & n24291;
  assign n24293 = ~n34781 & ~n34862;
  assign n24294 = ~n24292 & ~n24293;
  assign n24295 = ~n24287 & ~n34863;
  assign n24296 = ~n34861 & ~n34864;
  assign n24297 = ~n24279 & ~n24296;
  assign n24298 = ~n13548 & ~n24297;
  assign n24299 = n13548 & ~n24279;
  assign n24300 = ~n24296 & n24299;
  assign n24301 = ~n34782 & ~n23643;
  assign n24302 = ~n23643 & ~n24076;
  assign n24303 = ~n34782 & n24302;
  assign n24304 = ~n24076 & n24301;
  assign n24305 = n23469 & ~n34865;
  assign n24306 = n23642 & n24302;
  assign n24307 = n23469 & ~n34782;
  assign n24308 = ~n23643 & n24307;
  assign n24309 = ~n24076 & n24308;
  assign n24310 = ~n23469 & ~n34865;
  assign n24311 = ~n24309 & ~n24310;
  assign n24312 = ~n24305 & ~n24306;
  assign n24313 = ~n24300 & ~n34866;
  assign n24314 = ~n24298 & ~n24313;
  assign n24315 = ~n12948 & ~n24314;
  assign n24316 = ~n23645 & ~n23661;
  assign n24317 = ~n24076 & n24316;
  assign n24318 = ~n34785 & ~n24317;
  assign n24319 = n34785 & ~n23661;
  assign n24320 = ~n23645 & n24319;
  assign n24321 = n34785 & n24317;
  assign n24322 = ~n24076 & n24320;
  assign n24323 = ~n24318 & ~n34867;
  assign n24324 = n12948 & ~n24298;
  assign n24325 = ~n24313 & n24324;
  assign n24326 = n12948 & n24314;
  assign n24327 = ~n24323 & ~n34868;
  assign n24328 = ~n24315 & ~n24327;
  assign n24329 = ~n12296 & ~n24328;
  assign n24330 = n12296 & ~n24315;
  assign n24331 = ~n24327 & n24330;
  assign n24332 = ~n34786 & ~n23667;
  assign n24333 = ~n23667 & ~n24076;
  assign n24334 = ~n34786 & n24333;
  assign n24335 = ~n24076 & n24332;
  assign n24336 = n23461 & ~n34869;
  assign n24337 = n23666 & n24333;
  assign n24338 = n23461 & ~n34786;
  assign n24339 = ~n23667 & n24338;
  assign n24340 = ~n24076 & n24339;
  assign n24341 = ~n23461 & ~n34869;
  assign n24342 = ~n24340 & ~n24341;
  assign n24343 = ~n24336 & ~n24337;
  assign n24344 = ~n24331 & ~n34870;
  assign n24345 = ~n24329 & ~n24344;
  assign n24346 = ~n11719 & ~n24345;
  assign n24347 = n11719 & ~n24329;
  assign n24348 = ~n24344 & n24347;
  assign n24349 = n11719 & n24345;
  assign n24350 = ~n23669 & ~n23672;
  assign n24351 = ~n23672 & ~n24076;
  assign n24352 = ~n23669 & n24351;
  assign n24353 = ~n24076 & n24350;
  assign n24354 = n23453 & ~n34872;
  assign n24355 = n23670 & n24351;
  assign n24356 = n23453 & ~n23672;
  assign n24357 = ~n23669 & n24356;
  assign n24358 = ~n24076 & n24357;
  assign n24359 = ~n23453 & ~n34872;
  assign n24360 = ~n24358 & ~n24359;
  assign n24361 = ~n24354 & ~n24355;
  assign n24362 = ~n34871 & ~n34873;
  assign n24363 = ~n24346 & ~n24362;
  assign n24364 = ~n11097 & ~n24363;
  assign n24365 = n11097 & ~n24346;
  assign n24366 = ~n24362 & n24365;
  assign n24367 = ~n34787 & ~n23678;
  assign n24368 = ~n23678 & ~n24076;
  assign n24369 = ~n34787 & n24368;
  assign n24370 = ~n24076 & n24367;
  assign n24371 = n23445 & ~n34874;
  assign n24372 = n23677 & n24368;
  assign n24373 = n23445 & ~n34787;
  assign n24374 = ~n23678 & n24373;
  assign n24375 = ~n24076 & n24374;
  assign n24376 = ~n23445 & ~n34874;
  assign n24377 = ~n24375 & ~n24376;
  assign n24378 = ~n24371 & ~n24372;
  assign n24379 = ~n24366 & ~n34875;
  assign n24380 = ~n24364 & ~n24379;
  assign n24381 = ~n10555 & ~n24380;
  assign n24382 = ~n23680 & ~n23695;
  assign n24383 = ~n24076 & n24382;
  assign n24384 = ~n34789 & ~n24383;
  assign n24385 = n34789 & ~n23695;
  assign n24386 = ~n23680 & n24385;
  assign n24387 = n34789 & n24383;
  assign n24388 = ~n24076 & n24386;
  assign n24389 = ~n24384 & ~n34876;
  assign n24390 = n10555 & ~n24364;
  assign n24391 = ~n24379 & n24390;
  assign n24392 = n10555 & n24380;
  assign n24393 = ~n24389 & ~n34877;
  assign n24394 = ~n24381 & ~n24393;
  assign n24395 = ~n9969 & ~n24394;
  assign n24396 = n9969 & ~n24381;
  assign n24397 = ~n24393 & n24396;
  assign n24398 = ~n34790 & ~n23701;
  assign n24399 = ~n23701 & ~n24076;
  assign n24400 = ~n34790 & n24399;
  assign n24401 = ~n24076 & n24398;
  assign n24402 = n23437 & ~n34878;
  assign n24403 = n23700 & n24399;
  assign n24404 = n23437 & ~n34790;
  assign n24405 = ~n23701 & n24404;
  assign n24406 = ~n24076 & n24405;
  assign n24407 = ~n23437 & ~n34878;
  assign n24408 = ~n24406 & ~n24407;
  assign n24409 = ~n24402 & ~n24403;
  assign n24410 = ~n24397 & ~n34879;
  assign n24411 = ~n24395 & ~n24410;
  assign n24412 = ~n9457 & ~n24411;
  assign n24413 = n9457 & ~n24395;
  assign n24414 = ~n24410 & n24413;
  assign n24415 = n9457 & n24411;
  assign n24416 = ~n23703 & ~n23706;
  assign n24417 = ~n23706 & ~n24076;
  assign n24418 = ~n23703 & n24417;
  assign n24419 = ~n24076 & n24416;
  assign n24420 = n23429 & ~n34881;
  assign n24421 = n23704 & n24417;
  assign n24422 = n23429 & ~n23706;
  assign n24423 = ~n23703 & n24422;
  assign n24424 = ~n24076 & n24423;
  assign n24425 = ~n23429 & ~n34881;
  assign n24426 = ~n24424 & ~n24425;
  assign n24427 = ~n24420 & ~n24421;
  assign n24428 = ~n34880 & ~n34882;
  assign n24429 = ~n24412 & ~n24428;
  assign n24430 = ~n8896 & ~n24429;
  assign n24431 = n8896 & ~n24412;
  assign n24432 = ~n24428 & n24431;
  assign n24433 = ~n34791 & ~n23712;
  assign n24434 = ~n23712 & ~n24076;
  assign n24435 = ~n34791 & n24434;
  assign n24436 = ~n24076 & n24433;
  assign n24437 = n23421 & ~n34883;
  assign n24438 = n23711 & n24434;
  assign n24439 = n23421 & ~n34791;
  assign n24440 = ~n23712 & n24439;
  assign n24441 = ~n24076 & n24440;
  assign n24442 = ~n23421 & ~n34883;
  assign n24443 = ~n24441 & ~n24442;
  assign n24444 = ~n24437 & ~n24438;
  assign n24445 = ~n24432 & ~n34884;
  assign n24446 = ~n24430 & ~n24445;
  assign n24447 = ~n8411 & ~n24446;
  assign n24448 = ~n23714 & ~n23729;
  assign n24449 = ~n24076 & n24448;
  assign n24450 = ~n34793 & ~n24449;
  assign n24451 = n34793 & ~n23729;
  assign n24452 = ~n23714 & n24451;
  assign n24453 = n34793 & n24449;
  assign n24454 = ~n24076 & n24452;
  assign n24455 = ~n24450 & ~n34885;
  assign n24456 = n8411 & ~n24430;
  assign n24457 = ~n24445 & n24456;
  assign n24458 = n8411 & n24446;
  assign n24459 = ~n24455 & ~n34886;
  assign n24460 = ~n24447 & ~n24459;
  assign n24461 = ~n7885 & ~n24460;
  assign n24462 = n7885 & ~n24447;
  assign n24463 = ~n24459 & n24462;
  assign n24464 = ~n34794 & ~n23735;
  assign n24465 = ~n23735 & ~n24076;
  assign n24466 = ~n34794 & n24465;
  assign n24467 = ~n24076 & n24464;
  assign n24468 = n23413 & ~n34887;
  assign n24469 = n23734 & n24465;
  assign n24470 = n23413 & ~n34794;
  assign n24471 = ~n23735 & n24470;
  assign n24472 = ~n24076 & n24471;
  assign n24473 = ~n23413 & ~n34887;
  assign n24474 = ~n24472 & ~n24473;
  assign n24475 = ~n24468 & ~n24469;
  assign n24476 = ~n24463 & ~n34888;
  assign n24477 = ~n24461 & ~n24476;
  assign n24478 = ~n7428 & ~n24477;
  assign n24479 = n7428 & ~n24461;
  assign n24480 = ~n24476 & n24479;
  assign n24481 = n7428 & n24477;
  assign n24482 = ~n23737 & ~n23740;
  assign n24483 = ~n23740 & ~n24076;
  assign n24484 = ~n23737 & n24483;
  assign n24485 = ~n24076 & n24482;
  assign n24486 = n23405 & ~n34890;
  assign n24487 = n23738 & n24483;
  assign n24488 = n23405 & ~n23740;
  assign n24489 = ~n23737 & n24488;
  assign n24490 = ~n24076 & n24489;
  assign n24491 = ~n23405 & ~n34890;
  assign n24492 = ~n24490 & ~n24491;
  assign n24493 = ~n24486 & ~n24487;
  assign n24494 = ~n34889 & ~n34891;
  assign n24495 = ~n24478 & ~n24494;
  assign n24496 = ~n6937 & ~n24495;
  assign n24497 = n6937 & ~n24478;
  assign n24498 = ~n24494 & n24497;
  assign n24499 = ~n34795 & ~n23746;
  assign n24500 = ~n23746 & ~n24076;
  assign n24501 = ~n34795 & n24500;
  assign n24502 = ~n24076 & n24499;
  assign n24503 = n23397 & ~n34892;
  assign n24504 = n23745 & n24500;
  assign n24505 = n23397 & ~n34795;
  assign n24506 = ~n23746 & n24505;
  assign n24507 = ~n24076 & n24506;
  assign n24508 = ~n23397 & ~n34892;
  assign n24509 = ~n24507 & ~n24508;
  assign n24510 = ~n24503 & ~n24504;
  assign n24511 = ~n24498 & ~n34893;
  assign n24512 = ~n24496 & ~n24511;
  assign n24513 = ~n6507 & ~n24512;
  assign n24514 = ~n23748 & ~n23763;
  assign n24515 = ~n24076 & n24514;
  assign n24516 = ~n34797 & ~n24515;
  assign n24517 = n34797 & ~n23763;
  assign n24518 = ~n23748 & n24517;
  assign n24519 = n34797 & n24515;
  assign n24520 = ~n24076 & n24518;
  assign n24521 = ~n24516 & ~n34894;
  assign n24522 = n6507 & ~n24496;
  assign n24523 = ~n24511 & n24522;
  assign n24524 = n6507 & n24512;
  assign n24525 = ~n24521 & ~n34895;
  assign n24526 = ~n24513 & ~n24525;
  assign n24527 = ~n6051 & ~n24526;
  assign n24528 = n6051 & ~n24513;
  assign n24529 = ~n24525 & n24528;
  assign n24530 = ~n34798 & ~n23769;
  assign n24531 = ~n23769 & ~n24076;
  assign n24532 = ~n34798 & n24531;
  assign n24533 = ~n24076 & n24530;
  assign n24534 = n23389 & ~n34896;
  assign n24535 = n23768 & n24531;
  assign n24536 = n23389 & ~n34798;
  assign n24537 = ~n23769 & n24536;
  assign n24538 = ~n24076 & n24537;
  assign n24539 = ~n23389 & ~n34896;
  assign n24540 = ~n24538 & ~n24539;
  assign n24541 = ~n24534 & ~n24535;
  assign n24542 = ~n24529 & ~n34897;
  assign n24543 = ~n24527 & ~n24542;
  assign n24544 = ~n5648 & ~n24543;
  assign n24545 = n5648 & ~n24527;
  assign n24546 = ~n24542 & n24545;
  assign n24547 = n5648 & n24543;
  assign n24548 = ~n23771 & ~n23774;
  assign n24549 = ~n23774 & ~n24076;
  assign n24550 = ~n23771 & n24549;
  assign n24551 = ~n24076 & n24548;
  assign n24552 = n23381 & ~n34899;
  assign n24553 = n23772 & n24549;
  assign n24554 = n23381 & ~n23774;
  assign n24555 = ~n23771 & n24554;
  assign n24556 = ~n24076 & n24555;
  assign n24557 = ~n23381 & ~n34899;
  assign n24558 = ~n24556 & ~n24557;
  assign n24559 = ~n24552 & ~n24553;
  assign n24560 = ~n34898 & ~n34900;
  assign n24561 = ~n24544 & ~n24560;
  assign n24562 = ~n5223 & ~n24561;
  assign n24563 = n5223 & ~n24544;
  assign n24564 = ~n24560 & n24563;
  assign n24565 = ~n34799 & ~n23780;
  assign n24566 = ~n23780 & ~n24076;
  assign n24567 = ~n34799 & n24566;
  assign n24568 = ~n24076 & n24565;
  assign n24569 = n23373 & ~n34901;
  assign n24570 = n23779 & n24566;
  assign n24571 = n23373 & ~n34799;
  assign n24572 = ~n23780 & n24571;
  assign n24573 = ~n24076 & n24572;
  assign n24574 = ~n23373 & ~n34901;
  assign n24575 = ~n24573 & ~n24574;
  assign n24576 = ~n24569 & ~n24570;
  assign n24577 = ~n24564 & ~n34902;
  assign n24578 = ~n24562 & ~n24577;
  assign n24579 = ~n4851 & ~n24578;
  assign n24580 = ~n23782 & ~n23797;
  assign n24581 = ~n24076 & n24580;
  assign n24582 = ~n34801 & ~n24581;
  assign n24583 = n34801 & ~n23797;
  assign n24584 = ~n23782 & n24583;
  assign n24585 = n34801 & n24581;
  assign n24586 = ~n24076 & n24584;
  assign n24587 = ~n24582 & ~n34903;
  assign n24588 = n4851 & ~n24562;
  assign n24589 = ~n24577 & n24588;
  assign n24590 = n4851 & n24578;
  assign n24591 = ~n24587 & ~n34904;
  assign n24592 = ~n24579 & ~n24591;
  assign n24593 = ~n4461 & ~n24592;
  assign n24594 = n4461 & ~n24579;
  assign n24595 = ~n24591 & n24594;
  assign n24596 = ~n34802 & ~n23803;
  assign n24597 = ~n23803 & ~n24076;
  assign n24598 = ~n34802 & n24597;
  assign n24599 = ~n24076 & n24596;
  assign n24600 = n23365 & ~n34905;
  assign n24601 = n23802 & n24597;
  assign n24602 = n23365 & ~n34802;
  assign n24603 = ~n23803 & n24602;
  assign n24604 = ~n24076 & n24603;
  assign n24605 = ~n23365 & ~n34905;
  assign n24606 = ~n24604 & ~n24605;
  assign n24607 = ~n24600 & ~n24601;
  assign n24608 = ~n24595 & ~n34906;
  assign n24609 = ~n24593 & ~n24608;
  assign n24610 = ~n4115 & ~n24609;
  assign n24611 = n4115 & ~n24593;
  assign n24612 = ~n24608 & n24611;
  assign n24613 = n4115 & n24609;
  assign n24614 = ~n23805 & ~n23808;
  assign n24615 = ~n23808 & ~n24076;
  assign n24616 = ~n23805 & n24615;
  assign n24617 = ~n24076 & n24614;
  assign n24618 = n23357 & ~n34908;
  assign n24619 = n23806 & n24615;
  assign n24620 = n23357 & ~n23808;
  assign n24621 = ~n23805 & n24620;
  assign n24622 = ~n24076 & n24621;
  assign n24623 = ~n23357 & ~n34908;
  assign n24624 = ~n24622 & ~n24623;
  assign n24625 = ~n24618 & ~n24619;
  assign n24626 = ~n34907 & ~n34909;
  assign n24627 = ~n24610 & ~n24626;
  assign n24628 = ~n3754 & ~n24627;
  assign n24629 = n3754 & ~n24610;
  assign n24630 = ~n24626 & n24629;
  assign n24631 = ~n34803 & ~n23814;
  assign n24632 = ~n23814 & ~n24076;
  assign n24633 = ~n34803 & n24632;
  assign n24634 = ~n24076 & n24631;
  assign n24635 = n23349 & ~n34910;
  assign n24636 = n23813 & n24632;
  assign n24637 = n23349 & ~n34803;
  assign n24638 = ~n23814 & n24637;
  assign n24639 = ~n24076 & n24638;
  assign n24640 = ~n23349 & ~n34910;
  assign n24641 = ~n24639 & ~n24640;
  assign n24642 = ~n24635 & ~n24636;
  assign n24643 = ~n24630 & ~n34911;
  assign n24644 = ~n24628 & ~n24643;
  assign n24645 = ~n3444 & ~n24644;
  assign n24646 = ~n23816 & ~n23831;
  assign n24647 = ~n24076 & n24646;
  assign n24648 = ~n34805 & ~n24647;
  assign n24649 = n34805 & ~n23831;
  assign n24650 = ~n23816 & n24649;
  assign n24651 = n34805 & n24647;
  assign n24652 = ~n24076 & n24650;
  assign n24653 = ~n24648 & ~n34912;
  assign n24654 = n3444 & ~n24628;
  assign n24655 = ~n24643 & n24654;
  assign n24656 = n3444 & n24644;
  assign n24657 = ~n24653 & ~n34913;
  assign n24658 = ~n24645 & ~n24657;
  assign n24659 = ~n3116 & ~n24658;
  assign n24660 = n3116 & ~n24645;
  assign n24661 = ~n24657 & n24660;
  assign n24662 = ~n34806 & ~n23837;
  assign n24663 = ~n23837 & ~n24076;
  assign n24664 = ~n34806 & n24663;
  assign n24665 = ~n24076 & n24662;
  assign n24666 = n23341 & ~n34914;
  assign n24667 = n23836 & n24663;
  assign n24668 = n23341 & ~n34806;
  assign n24669 = ~n23837 & n24668;
  assign n24670 = ~n24076 & n24669;
  assign n24671 = ~n23341 & ~n34914;
  assign n24672 = ~n24670 & ~n24671;
  assign n24673 = ~n24666 & ~n24667;
  assign n24674 = ~n24661 & ~n34915;
  assign n24675 = ~n24659 & ~n24674;
  assign n24676 = ~n2833 & ~n24675;
  assign n24677 = n2833 & ~n24659;
  assign n24678 = ~n24674 & n24677;
  assign n24679 = n2833 & n24675;
  assign n24680 = ~n23839 & ~n23842;
  assign n24681 = ~n23842 & ~n24076;
  assign n24682 = ~n23839 & n24681;
  assign n24683 = ~n24076 & n24680;
  assign n24684 = n23333 & ~n34917;
  assign n24685 = n23840 & n24681;
  assign n24686 = n23333 & ~n23842;
  assign n24687 = ~n23839 & n24686;
  assign n24688 = ~n24076 & n24687;
  assign n24689 = ~n23333 & ~n34917;
  assign n24690 = ~n24688 & ~n24689;
  assign n24691 = ~n24684 & ~n24685;
  assign n24692 = ~n34916 & ~n34918;
  assign n24693 = ~n24676 & ~n24692;
  assign n24694 = ~n2536 & ~n24693;
  assign n24695 = n2536 & ~n24676;
  assign n24696 = ~n24692 & n24695;
  assign n24697 = ~n34807 & ~n23848;
  assign n24698 = ~n23848 & ~n24076;
  assign n24699 = ~n34807 & n24698;
  assign n24700 = ~n24076 & n24697;
  assign n24701 = n23325 & ~n34919;
  assign n24702 = n23847 & n24698;
  assign n24703 = n23325 & ~n34807;
  assign n24704 = ~n23848 & n24703;
  assign n24705 = ~n24076 & n24704;
  assign n24706 = ~n23325 & ~n34919;
  assign n24707 = ~n24705 & ~n24706;
  assign n24708 = ~n24701 & ~n24702;
  assign n24709 = ~n24696 & ~n34920;
  assign n24710 = ~n24694 & ~n24709;
  assign n24711 = ~n2283 & ~n24710;
  assign n24712 = ~n23850 & ~n23865;
  assign n24713 = ~n24076 & n24712;
  assign n24714 = ~n34809 & ~n24713;
  assign n24715 = n34809 & ~n23865;
  assign n24716 = ~n23850 & n24715;
  assign n24717 = n34809 & n24713;
  assign n24718 = ~n24076 & n24716;
  assign n24719 = ~n24714 & ~n34921;
  assign n24720 = n2283 & ~n24694;
  assign n24721 = ~n24709 & n24720;
  assign n24722 = n2283 & n24710;
  assign n24723 = ~n24719 & ~n34922;
  assign n24724 = ~n24711 & ~n24723;
  assign n24725 = ~n2021 & ~n24724;
  assign n24726 = n2021 & ~n24711;
  assign n24727 = ~n24723 & n24726;
  assign n24728 = ~n34810 & ~n23871;
  assign n24729 = ~n23871 & ~n24076;
  assign n24730 = ~n34810 & n24729;
  assign n24731 = ~n24076 & n24728;
  assign n24732 = n23317 & ~n34923;
  assign n24733 = n23870 & n24729;
  assign n24734 = n23317 & ~n34810;
  assign n24735 = ~n23871 & n24734;
  assign n24736 = ~n24076 & n24735;
  assign n24737 = ~n23317 & ~n34923;
  assign n24738 = ~n24736 & ~n24737;
  assign n24739 = ~n24732 & ~n24733;
  assign n24740 = ~n24727 & ~n34924;
  assign n24741 = ~n24725 & ~n24740;
  assign n24742 = ~n1796 & ~n24741;
  assign n24743 = n1796 & ~n24725;
  assign n24744 = ~n24740 & n24743;
  assign n24745 = n1796 & n24741;
  assign n24746 = ~n23873 & ~n23876;
  assign n24747 = ~n23876 & ~n24076;
  assign n24748 = ~n23873 & n24747;
  assign n24749 = ~n24076 & n24746;
  assign n24750 = n23309 & ~n34926;
  assign n24751 = n23874 & n24747;
  assign n24752 = n23309 & ~n23876;
  assign n24753 = ~n23873 & n24752;
  assign n24754 = ~n24076 & n24753;
  assign n24755 = ~n23309 & ~n34926;
  assign n24756 = ~n24754 & ~n24755;
  assign n24757 = ~n24750 & ~n24751;
  assign n24758 = ~n34925 & ~n34927;
  assign n24759 = ~n24742 & ~n24758;
  assign n24760 = ~n1567 & ~n24759;
  assign n24761 = n1567 & ~n24742;
  assign n24762 = ~n24758 & n24761;
  assign n24763 = ~n34811 & ~n23882;
  assign n24764 = ~n23882 & ~n24076;
  assign n24765 = ~n34811 & n24764;
  assign n24766 = ~n24076 & n24763;
  assign n24767 = n23301 & ~n34928;
  assign n24768 = n23881 & n24764;
  assign n24769 = n23301 & ~n34811;
  assign n24770 = ~n23882 & n24769;
  assign n24771 = ~n24076 & n24770;
  assign n24772 = ~n23301 & ~n34928;
  assign n24773 = ~n24771 & ~n24772;
  assign n24774 = ~n24767 & ~n24768;
  assign n24775 = ~n24762 & ~n34929;
  assign n24776 = ~n24760 & ~n24775;
  assign n24777 = ~n1374 & ~n24776;
  assign n24778 = ~n23884 & ~n23899;
  assign n24779 = ~n24076 & n24778;
  assign n24780 = ~n34813 & ~n24779;
  assign n24781 = n34813 & ~n23899;
  assign n24782 = ~n23884 & n24781;
  assign n24783 = n34813 & n24779;
  assign n24784 = ~n24076 & n24782;
  assign n24785 = ~n24780 & ~n34930;
  assign n24786 = n1374 & ~n24760;
  assign n24787 = ~n24775 & n24786;
  assign n24788 = n1374 & n24776;
  assign n24789 = ~n24785 & ~n34931;
  assign n24790 = ~n24777 & ~n24789;
  assign n24791 = ~n1179 & ~n24790;
  assign n24792 = n1179 & ~n24777;
  assign n24793 = ~n24789 & n24792;
  assign n24794 = ~n34814 & ~n23905;
  assign n24795 = ~n23905 & ~n24076;
  assign n24796 = ~n34814 & n24795;
  assign n24797 = ~n24076 & n24794;
  assign n24798 = n23293 & ~n34932;
  assign n24799 = n23904 & n24795;
  assign n24800 = n23293 & ~n34814;
  assign n24801 = ~n23905 & n24800;
  assign n24802 = ~n24076 & n24801;
  assign n24803 = ~n23293 & ~n34932;
  assign n24804 = ~n24802 & ~n24803;
  assign n24805 = ~n24798 & ~n24799;
  assign n24806 = ~n24793 & ~n34933;
  assign n24807 = ~n24791 & ~n24806;
  assign n24808 = ~n1016 & ~n24807;
  assign n24809 = n1016 & ~n24791;
  assign n24810 = ~n24806 & n24809;
  assign n24811 = n1016 & n24807;
  assign n24812 = ~n23907 & ~n23910;
  assign n24813 = ~n23910 & ~n24076;
  assign n24814 = ~n23907 & n24813;
  assign n24815 = ~n24076 & n24812;
  assign n24816 = n23285 & ~n34935;
  assign n24817 = n23908 & n24813;
  assign n24818 = n23285 & ~n23910;
  assign n24819 = ~n23907 & n24818;
  assign n24820 = ~n24076 & n24819;
  assign n24821 = ~n23285 & ~n34935;
  assign n24822 = ~n24820 & ~n24821;
  assign n24823 = ~n24816 & ~n24817;
  assign n24824 = ~n34934 & ~n34936;
  assign n24825 = ~n24808 & ~n24824;
  assign n24826 = ~n855 & ~n24825;
  assign n24827 = n855 & ~n24808;
  assign n24828 = ~n24824 & n24827;
  assign n24829 = ~n34815 & ~n23916;
  assign n24830 = ~n24076 & n24829;
  assign n24831 = n23277 & ~n24830;
  assign n24832 = ~n23277 & n24830;
  assign n24833 = n23277 & ~n34815;
  assign n24834 = ~n23916 & n24833;
  assign n24835 = ~n24076 & n24834;
  assign n24836 = ~n23277 & ~n24830;
  assign n24837 = ~n24835 & ~n24836;
  assign n24838 = ~n24831 & ~n24832;
  assign n24839 = ~n24828 & ~n34937;
  assign n24840 = ~n24826 & ~n24839;
  assign n24841 = ~n720 & ~n24840;
  assign n24842 = ~n23918 & ~n23930;
  assign n24843 = ~n24076 & n24842;
  assign n24844 = ~n34816 & n24843;
  assign n24845 = n34816 & ~n24843;
  assign n24846 = ~n23918 & n34816;
  assign n24847 = ~n23930 & n24846;
  assign n24848 = ~n24076 & n24847;
  assign n24849 = ~n34816 & ~n24843;
  assign n24850 = ~n24848 & ~n24849;
  assign n24851 = ~n24844 & ~n24845;
  assign n24852 = n720 & ~n24826;
  assign n24853 = ~n24839 & n24852;
  assign n24854 = n720 & n24840;
  assign n24855 = ~n34938 & ~n34939;
  assign n24856 = ~n24841 & ~n24855;
  assign n24857 = ~n592 & ~n24856;
  assign n24858 = n592 & ~n24841;
  assign n24859 = ~n24855 & n24858;
  assign n24860 = ~n23933 & ~n34818;
  assign n24861 = ~n23933 & ~n24076;
  assign n24862 = ~n34818 & n24861;
  assign n24863 = ~n24076 & n24860;
  assign n24864 = n23941 & ~n34940;
  assign n24865 = n23945 & n24861;
  assign n24866 = n23941 & ~n34818;
  assign n24867 = ~n23933 & n24866;
  assign n24868 = ~n24076 & n24867;
  assign n24869 = ~n23941 & ~n34940;
  assign n24870 = ~n24868 & ~n24869;
  assign n24871 = ~n24864 & ~n24865;
  assign n24872 = ~n24859 & ~n34941;
  assign n24873 = ~n24857 & ~n24872;
  assign n24874 = ~n487 & ~n24873;
  assign n24875 = ~n23947 & ~n23949;
  assign n24876 = ~n24076 & n24875;
  assign n24877 = ~n34820 & ~n24876;
  assign n24878 = ~n23947 & n34820;
  assign n24879 = ~n23949 & n24878;
  assign n24880 = n34820 & n24876;
  assign n24881 = ~n24076 & n24879;
  assign n24882 = ~n24877 & ~n34942;
  assign n24883 = n487 & ~n24857;
  assign n24884 = ~n24872 & n24883;
  assign n24885 = n487 & n24873;
  assign n24886 = ~n24882 & ~n34943;
  assign n24887 = ~n24874 & ~n24886;
  assign n24888 = ~n393 & ~n24887;
  assign n24889 = n393 & ~n24874;
  assign n24890 = ~n24886 & n24889;
  assign n24891 = ~n23964 & ~n34822;
  assign n24892 = ~n23964 & ~n24076;
  assign n24893 = ~n34822 & n24892;
  assign n24894 = ~n24076 & n24891;
  assign n24895 = n23972 & ~n34944;
  assign n24896 = n23976 & n24892;
  assign n24897 = n23972 & ~n34822;
  assign n24898 = ~n23964 & n24897;
  assign n24899 = ~n24076 & n24898;
  assign n24900 = ~n23972 & ~n34944;
  assign n24901 = ~n24899 & ~n24900;
  assign n24902 = ~n24895 & ~n24896;
  assign n24903 = ~n24890 & ~n34945;
  assign n24904 = ~n24888 & ~n24903;
  assign n24905 = ~n321 & ~n24904;
  assign n24906 = ~n23978 & ~n23980;
  assign n24907 = ~n24076 & n24906;
  assign n24908 = ~n34824 & ~n24907;
  assign n24909 = ~n23978 & n34824;
  assign n24910 = ~n23980 & n24909;
  assign n24911 = n34824 & n24907;
  assign n24912 = ~n24076 & n24910;
  assign n24913 = ~n24908 & ~n34946;
  assign n24914 = n321 & ~n24888;
  assign n24915 = ~n24903 & n24914;
  assign n24916 = n321 & n24904;
  assign n24917 = ~n24913 & ~n34947;
  assign n24918 = ~n24905 & ~n24917;
  assign n24919 = ~n263 & ~n24918;
  assign n24920 = n263 & ~n24905;
  assign n24921 = ~n24917 & n24920;
  assign n24922 = ~n23995 & ~n34826;
  assign n24923 = ~n23995 & ~n24076;
  assign n24924 = ~n34826 & n24923;
  assign n24925 = ~n24076 & n24922;
  assign n24926 = n24003 & ~n34948;
  assign n24927 = n24007 & n24923;
  assign n24928 = n24003 & ~n34826;
  assign n24929 = ~n23995 & n24928;
  assign n24930 = ~n24076 & n24929;
  assign n24931 = ~n24003 & ~n34948;
  assign n24932 = ~n24930 & ~n24931;
  assign n24933 = ~n24926 & ~n24927;
  assign n24934 = ~n24921 & ~n34949;
  assign n24935 = ~n24919 & ~n24934;
  assign n24936 = ~n214 & ~n24935;
  assign n24937 = n214 & ~n24919;
  assign n24938 = ~n24934 & n24937;
  assign n24939 = n214 & n24935;
  assign n24940 = ~n24009 & ~n24019;
  assign n24941 = ~n24009 & ~n24076;
  assign n24942 = ~n24019 & n24941;
  assign n24943 = ~n24076 & n24940;
  assign n24944 = n24017 & ~n34951;
  assign n24945 = n24020 & n24941;
  assign n24946 = ~n24009 & n24017;
  assign n24947 = ~n24019 & n24946;
  assign n24948 = ~n24076 & n24947;
  assign n24949 = ~n24017 & ~n34951;
  assign n24950 = ~n24948 & ~n24949;
  assign n24951 = ~n24944 & ~n24945;
  assign n24952 = ~n34950 & ~n34952;
  assign n24953 = ~n24936 & ~n24952;
  assign n24954 = ~n197 & ~n24953;
  assign n24955 = n197 & ~n24936;
  assign n24956 = ~n24952 & n24955;
  assign n24957 = ~n24022 & ~n34829;
  assign n24958 = ~n24022 & ~n24076;
  assign n24959 = ~n34829 & n24958;
  assign n24960 = ~n24076 & n24957;
  assign n24961 = n24030 & ~n34953;
  assign n24962 = n24034 & n24958;
  assign n24963 = n24030 & ~n34829;
  assign n24964 = ~n24022 & n24963;
  assign n24965 = ~n24076 & n24964;
  assign n24966 = ~n24030 & ~n34953;
  assign n24967 = ~n24965 & ~n24966;
  assign n24968 = ~n24961 & ~n24962;
  assign n24969 = ~n24956 & ~n34954;
  assign n24970 = ~n24954 & ~n24969;
  assign n24971 = ~n24036 & ~n24038;
  assign n24972 = ~n24076 & n24971;
  assign n24973 = ~n34831 & ~n24972;
  assign n24974 = ~n24036 & n34831;
  assign n24975 = ~n24038 & n24974;
  assign n24976 = n34831 & n24972;
  assign n24977 = ~n24076 & n24975;
  assign n24978 = ~n24973 & ~n34955;
  assign n24979 = ~n24052 & ~n24060;
  assign n24980 = ~n24060 & ~n24076;
  assign n24981 = ~n24052 & n24980;
  assign n24982 = ~n24076 & n24979;
  assign n24983 = ~n34834 & ~n34956;
  assign n24984 = ~n24978 & n24983;
  assign n24985 = ~n24970 & n24984;
  assign n24986 = n193 & ~n24985;
  assign n24987 = ~n24954 & n24978;
  assign n24988 = ~n24969 & n24987;
  assign n24989 = n24970 & n24978;
  assign n24990 = n24052 & ~n24980;
  assign n24991 = ~n193 & ~n24979;
  assign n24992 = ~n24990 & n24991;
  assign n24993 = ~n34957 & ~n24992;
  assign n24994 = ~n24986 & n24993;
  assign n24995 = ~n24808 & ~n34934;
  assign n24996 = ~n24994 & n24995;
  assign n24997 = ~n34936 & ~n24996;
  assign n24998 = ~n24808 & n34936;
  assign n24999 = ~n34934 & n24998;
  assign n25000 = n34936 & n24996;
  assign n25001 = ~n24994 & n24999;
  assign n25002 = ~n24997 & ~n34958;
  assign n25003 = ~n24791 & ~n24793;
  assign n25004 = ~n24994 & n25003;
  assign n25005 = ~n34933 & ~n25004;
  assign n25006 = ~n24793 & n34933;
  assign n25007 = ~n24791 & n25006;
  assign n25008 = n34933 & n25004;
  assign n25009 = ~n24994 & n25007;
  assign n25010 = ~n25005 & ~n34959;
  assign n25011 = ~n24760 & ~n24762;
  assign n25012 = ~n24994 & n25011;
  assign n25013 = ~n34929 & ~n25012;
  assign n25014 = ~n24762 & n34929;
  assign n25015 = ~n24760 & n25014;
  assign n25016 = n34929 & n25012;
  assign n25017 = ~n24994 & n25015;
  assign n25018 = ~n25013 & ~n34960;
  assign n25019 = ~n24742 & ~n34925;
  assign n25020 = ~n24994 & n25019;
  assign n25021 = ~n34927 & ~n25020;
  assign n25022 = ~n24742 & n34927;
  assign n25023 = ~n34925 & n25022;
  assign n25024 = n34927 & n25020;
  assign n25025 = ~n24994 & n25023;
  assign n25026 = ~n25021 & ~n34961;
  assign n25027 = ~n24725 & ~n24727;
  assign n25028 = ~n24994 & n25027;
  assign n25029 = ~n34924 & ~n25028;
  assign n25030 = ~n24727 & n34924;
  assign n25031 = ~n24725 & n25030;
  assign n25032 = n34924 & n25028;
  assign n25033 = ~n24994 & n25031;
  assign n25034 = ~n25029 & ~n34962;
  assign n25035 = ~n24694 & ~n24696;
  assign n25036 = ~n24994 & n25035;
  assign n25037 = ~n34920 & ~n25036;
  assign n25038 = ~n24696 & n34920;
  assign n25039 = ~n24694 & n25038;
  assign n25040 = n34920 & n25036;
  assign n25041 = ~n24994 & n25039;
  assign n25042 = ~n25037 & ~n34963;
  assign n25043 = ~n24676 & ~n34916;
  assign n25044 = ~n24994 & n25043;
  assign n25045 = ~n34918 & ~n25044;
  assign n25046 = ~n24676 & n34918;
  assign n25047 = ~n34916 & n25046;
  assign n25048 = n34918 & n25044;
  assign n25049 = ~n24994 & n25047;
  assign n25050 = ~n25045 & ~n34964;
  assign n25051 = ~n24659 & ~n24661;
  assign n25052 = ~n24994 & n25051;
  assign n25053 = ~n34915 & ~n25052;
  assign n25054 = ~n24661 & n34915;
  assign n25055 = ~n24659 & n25054;
  assign n25056 = n34915 & n25052;
  assign n25057 = ~n24994 & n25055;
  assign n25058 = ~n25053 & ~n34965;
  assign n25059 = ~n24628 & ~n24630;
  assign n25060 = ~n24994 & n25059;
  assign n25061 = ~n34911 & ~n25060;
  assign n25062 = ~n24630 & n34911;
  assign n25063 = ~n24628 & n25062;
  assign n25064 = n34911 & n25060;
  assign n25065 = ~n24994 & n25063;
  assign n25066 = ~n25061 & ~n34966;
  assign n25067 = ~n24610 & ~n34907;
  assign n25068 = ~n24994 & n25067;
  assign n25069 = ~n34909 & ~n25068;
  assign n25070 = ~n24610 & n34909;
  assign n25071 = ~n34907 & n25070;
  assign n25072 = n34909 & n25068;
  assign n25073 = ~n24994 & n25071;
  assign n25074 = ~n25069 & ~n34967;
  assign n25075 = ~n24593 & ~n24595;
  assign n25076 = ~n24994 & n25075;
  assign n25077 = ~n34906 & ~n25076;
  assign n25078 = ~n24595 & n34906;
  assign n25079 = ~n24593 & n25078;
  assign n25080 = n34906 & n25076;
  assign n25081 = ~n24994 & n25079;
  assign n25082 = ~n25077 & ~n34968;
  assign n25083 = ~n24562 & ~n24564;
  assign n25084 = ~n24994 & n25083;
  assign n25085 = ~n34902 & ~n25084;
  assign n25086 = ~n24564 & n34902;
  assign n25087 = ~n24562 & n25086;
  assign n25088 = n34902 & n25084;
  assign n25089 = ~n24994 & n25087;
  assign n25090 = ~n25085 & ~n34969;
  assign n25091 = ~n24544 & ~n34898;
  assign n25092 = ~n24994 & n25091;
  assign n25093 = ~n34900 & ~n25092;
  assign n25094 = ~n24544 & n34900;
  assign n25095 = ~n34898 & n25094;
  assign n25096 = n34900 & n25092;
  assign n25097 = ~n24994 & n25095;
  assign n25098 = ~n25093 & ~n34970;
  assign n25099 = ~n24527 & ~n24529;
  assign n25100 = ~n24994 & n25099;
  assign n25101 = ~n34897 & ~n25100;
  assign n25102 = ~n24529 & n34897;
  assign n25103 = ~n24527 & n25102;
  assign n25104 = n34897 & n25100;
  assign n25105 = ~n24994 & n25103;
  assign n25106 = ~n25101 & ~n34971;
  assign n25107 = ~n24496 & ~n24498;
  assign n25108 = ~n24994 & n25107;
  assign n25109 = ~n34893 & ~n25108;
  assign n25110 = ~n24498 & n34893;
  assign n25111 = ~n24496 & n25110;
  assign n25112 = n34893 & n25108;
  assign n25113 = ~n24994 & n25111;
  assign n25114 = ~n25109 & ~n34972;
  assign n25115 = ~n24478 & ~n34889;
  assign n25116 = ~n24994 & n25115;
  assign n25117 = ~n34891 & ~n25116;
  assign n25118 = ~n24478 & n34891;
  assign n25119 = ~n34889 & n25118;
  assign n25120 = n34891 & n25116;
  assign n25121 = ~n24994 & n25119;
  assign n25122 = ~n25117 & ~n34973;
  assign n25123 = ~n24461 & ~n24463;
  assign n25124 = ~n24994 & n25123;
  assign n25125 = ~n34888 & ~n25124;
  assign n25126 = ~n24463 & n34888;
  assign n25127 = ~n24461 & n25126;
  assign n25128 = n34888 & n25124;
  assign n25129 = ~n24994 & n25127;
  assign n25130 = ~n25125 & ~n34974;
  assign n25131 = ~n24430 & ~n24432;
  assign n25132 = ~n24994 & n25131;
  assign n25133 = ~n34884 & ~n25132;
  assign n25134 = ~n24432 & n34884;
  assign n25135 = ~n24430 & n25134;
  assign n25136 = n34884 & n25132;
  assign n25137 = ~n24994 & n25135;
  assign n25138 = ~n25133 & ~n34975;
  assign n25139 = ~n24412 & ~n34880;
  assign n25140 = ~n24994 & n25139;
  assign n25141 = ~n34882 & ~n25140;
  assign n25142 = ~n24412 & n34882;
  assign n25143 = ~n34880 & n25142;
  assign n25144 = n34882 & n25140;
  assign n25145 = ~n24994 & n25143;
  assign n25146 = ~n25141 & ~n34976;
  assign n25147 = ~n24395 & ~n24397;
  assign n25148 = ~n24994 & n25147;
  assign n25149 = ~n34879 & ~n25148;
  assign n25150 = ~n24397 & n34879;
  assign n25151 = ~n24395 & n25150;
  assign n25152 = n34879 & n25148;
  assign n25153 = ~n24994 & n25151;
  assign n25154 = ~n25149 & ~n34977;
  assign n25155 = ~n24364 & ~n24366;
  assign n25156 = ~n24994 & n25155;
  assign n25157 = ~n34875 & ~n25156;
  assign n25158 = ~n24366 & n34875;
  assign n25159 = ~n24364 & n25158;
  assign n25160 = n34875 & n25156;
  assign n25161 = ~n24994 & n25159;
  assign n25162 = ~n25157 & ~n34978;
  assign n25163 = ~n24346 & ~n34871;
  assign n25164 = ~n24994 & n25163;
  assign n25165 = ~n34873 & ~n25164;
  assign n25166 = ~n24346 & n34873;
  assign n25167 = ~n34871 & n25166;
  assign n25168 = n34873 & n25164;
  assign n25169 = ~n24994 & n25167;
  assign n25170 = ~n25165 & ~n34979;
  assign n25171 = ~n24329 & ~n24331;
  assign n25172 = ~n24994 & n25171;
  assign n25173 = ~n34870 & ~n25172;
  assign n25174 = ~n24331 & n34870;
  assign n25175 = ~n24329 & n25174;
  assign n25176 = n34870 & n25172;
  assign n25177 = ~n24994 & n25175;
  assign n25178 = ~n25173 & ~n34980;
  assign n25179 = ~n24298 & ~n24300;
  assign n25180 = ~n24994 & n25179;
  assign n25181 = ~n34866 & ~n25180;
  assign n25182 = ~n24300 & n34866;
  assign n25183 = ~n24298 & n25182;
  assign n25184 = n34866 & n25180;
  assign n25185 = ~n24994 & n25183;
  assign n25186 = ~n25181 & ~n34981;
  assign n25187 = ~n24279 & ~n34861;
  assign n25188 = ~n24994 & n25187;
  assign n25189 = ~n34864 & ~n25188;
  assign n25190 = ~n24279 & n34864;
  assign n25191 = ~n34861 & n25190;
  assign n25192 = n34864 & n25188;
  assign n25193 = ~n24994 & n25191;
  assign n25194 = ~n25189 & ~n34982;
  assign n25195 = ~n24262 & ~n24264;
  assign n25196 = ~n24994 & n25195;
  assign n25197 = ~n34860 & ~n25196;
  assign n25198 = ~n24264 & n34860;
  assign n25199 = ~n24262 & n25198;
  assign n25200 = n34860 & n25196;
  assign n25201 = ~n24994 & n25199;
  assign n25202 = ~n25197 & ~n34983;
  assign n25203 = ~n24228 & ~n24230;
  assign n25204 = ~n24994 & n25203;
  assign n25205 = ~n34855 & ~n25204;
  assign n25206 = ~n24230 & n34855;
  assign n25207 = ~n24228 & n25206;
  assign n25208 = n34855 & n25204;
  assign n25209 = ~n24994 & n25207;
  assign n25210 = ~n25205 & ~n34984;
  assign n25211 = ~n24195 & ~n24197;
  assign n25212 = ~n24994 & n25211;
  assign n25213 = ~n34851 & ~n25212;
  assign n25214 = ~n24197 & n34851;
  assign n25215 = ~n24195 & n25214;
  assign n25216 = n34851 & n25212;
  assign n25217 = ~n24994 & n25215;
  assign n25218 = ~n25213 & ~n34985;
  assign n25219 = ~n24162 & ~n24164;
  assign n25220 = ~n24994 & n25219;
  assign n25221 = ~n34847 & ~n25220;
  assign n25222 = ~n24164 & n34847;
  assign n25223 = ~n24162 & n25222;
  assign n25224 = n34847 & n25220;
  assign n25225 = ~n24994 & n25223;
  assign n25226 = ~n25221 & ~n34986;
  assign n25227 = ~n24128 & ~n24130;
  assign n25228 = ~n24994 & n25227;
  assign n25229 = ~n34842 & ~n25228;
  assign n25230 = ~n24130 & n34842;
  assign n25231 = ~n24128 & n25230;
  assign n25232 = n34842 & n25228;
  assign n25233 = ~n24994 & n25231;
  assign n25234 = ~n25229 & ~n34987;
  assign n25235 = ~n24101 & ~n24103;
  assign n25236 = ~n24994 & n25235;
  assign n25237 = ~n24112 & ~n25236;
  assign n25238 = ~n24103 & n24112;
  assign n25239 = ~n24101 & n25238;
  assign n25240 = n24112 & n25236;
  assign n25241 = ~n24994 & n25239;
  assign n25242 = ~n25237 & ~n34988;
  assign n25243 = ~pi14  & ~n24994;
  assign n25244 = ~pi15  & n25243;
  assign n25245 = n24078 & ~n24994;
  assign n25246 = ~n24076 & ~n24992;
  assign n25247 = ~n34957 & n25246;
  assign n25248 = ~n24986 & n25247;
  assign n25249 = ~n34989 & ~n25248;
  assign n25250 = pi16  & ~n25249;
  assign n25251 = ~pi16  & ~n25248;
  assign n25252 = ~pi16  & n25249;
  assign n25253 = ~n34989 & n25251;
  assign n25254 = ~n25250 & ~n34990;
  assign n25255 = pi14  & ~n24994;
  assign n25256 = ~pi12  & ~pi13 ;
  assign n25257 = ~pi14  & n25256;
  assign n25258 = ~n23250 & ~n34836;
  assign n25259 = ~n23251 & n25258;
  assign n25260 = ~n23267 & n25259;
  assign n25261 = ~n34736 & n25260;
  assign n25262 = n34734 & n23269;
  assign n25263 = ~n23261 & n25261;
  assign n25264 = ~n25257 & ~n34991;
  assign n25265 = ~n24074 & n25264;
  assign n25266 = ~n34834 & n25265;
  assign n25267 = ~n24068 & n25266;
  assign n25268 = ~n25255 & ~n25257;
  assign n25269 = n24076 & n25268;
  assign n25270 = ~n25255 & n25267;
  assign n25271 = pi15  & ~n25243;
  assign n25272 = ~n34989 & ~n25271;
  assign n25273 = ~n34992 & n25272;
  assign n25274 = ~n24076 & ~n25268;
  assign n25275 = n23269 & ~n25274;
  assign n25276 = ~n25273 & ~n25274;
  assign n25277 = n23269 & n25276;
  assign n25278 = ~n25273 & n25275;
  assign n25279 = ~n25254 & ~n34993;
  assign n25280 = ~n23269 & ~n25276;
  assign n25281 = n22386 & ~n25280;
  assign n25282 = ~n25279 & n25281;
  assign n25283 = ~n24081 & ~n34837;
  assign n25284 = ~n24994 & n25283;
  assign n25285 = n24086 & ~n25284;
  assign n25286 = ~n24086 & n25283;
  assign n25287 = ~n24086 & n25284;
  assign n25288 = ~n24994 & n25286;
  assign n25289 = ~n25285 & ~n34994;
  assign n25290 = ~n25282 & ~n25289;
  assign n25291 = ~n25279 & ~n25280;
  assign n25292 = ~n22386 & ~n25291;
  assign n25293 = n21612 & ~n25292;
  assign n25294 = ~n25290 & ~n25292;
  assign n25295 = n21612 & n25294;
  assign n25296 = ~n25290 & n25293;
  assign n25297 = ~n25242 & ~n34995;
  assign n25298 = ~n21612 & ~n25294;
  assign n25299 = n20762 & ~n25298;
  assign n25300 = ~n25297 & n25299;
  assign n25301 = ~n24115 & ~n34839;
  assign n25302 = ~n24994 & n25301;
  assign n25303 = ~n24125 & ~n25302;
  assign n25304 = ~n24115 & n24125;
  assign n25305 = ~n34839 & n25304;
  assign n25306 = n24125 & n25302;
  assign n25307 = ~n24994 & n25305;
  assign n25308 = n24125 & ~n25302;
  assign n25309 = ~n24125 & n25302;
  assign n25310 = ~n25308 & ~n25309;
  assign n25311 = ~n25303 & ~n34996;
  assign n25312 = ~n25300 & n34997;
  assign n25313 = ~n25297 & ~n25298;
  assign n25314 = ~n20762 & ~n25313;
  assign n25315 = n20011 & ~n25314;
  assign n25316 = ~n25312 & ~n25314;
  assign n25317 = n20011 & n25316;
  assign n25318 = ~n25312 & n25315;
  assign n25319 = ~n25234 & ~n34998;
  assign n25320 = ~n20011 & ~n25316;
  assign n25321 = n19190 & ~n25320;
  assign n25322 = ~n25319 & n25321;
  assign n25323 = ~n24145 & ~n34843;
  assign n25324 = ~n24994 & n25323;
  assign n25325 = ~n34845 & ~n25324;
  assign n25326 = n34845 & n25324;
  assign n25327 = ~n24145 & ~n34845;
  assign n25328 = ~n34843 & n25327;
  assign n25329 = ~n24994 & n25328;
  assign n25330 = n34845 & ~n25324;
  assign n25331 = ~n25329 & ~n25330;
  assign n25332 = ~n25325 & ~n25326;
  assign n25333 = ~n25322 & ~n34999;
  assign n25334 = ~n25319 & ~n25320;
  assign n25335 = ~n19190 & ~n25334;
  assign n25336 = n18472 & ~n25335;
  assign n25337 = ~n25333 & ~n25335;
  assign n25338 = n18472 & n25337;
  assign n25339 = ~n25333 & n25336;
  assign n25340 = ~n25226 & ~n35000;
  assign n25341 = ~n18472 & ~n25337;
  assign n25342 = n17690 & ~n25341;
  assign n25343 = ~n25340 & n25342;
  assign n25344 = ~n24179 & ~n34848;
  assign n25345 = ~n24994 & n25344;
  assign n25346 = ~n34849 & n25345;
  assign n25347 = n34849 & ~n25345;
  assign n25348 = ~n24179 & n34849;
  assign n25349 = ~n34848 & n25348;
  assign n25350 = ~n24994 & n25349;
  assign n25351 = ~n34849 & ~n25345;
  assign n25352 = ~n25350 & ~n25351;
  assign n25353 = ~n25346 & ~n25347;
  assign n25354 = ~n25343 & ~n35001;
  assign n25355 = ~n25340 & ~n25341;
  assign n25356 = ~n17690 & ~n25355;
  assign n25357 = n17001 & ~n25356;
  assign n25358 = ~n25354 & ~n25356;
  assign n25359 = n17001 & n25358;
  assign n25360 = ~n25354 & n25357;
  assign n25361 = ~n25218 & ~n35002;
  assign n25362 = ~n17001 & ~n25358;
  assign n25363 = n16248 & ~n25362;
  assign n25364 = ~n25361 & n25363;
  assign n25365 = ~n24212 & ~n34852;
  assign n25366 = ~n24994 & n25365;
  assign n25367 = ~n34853 & n25366;
  assign n25368 = n34853 & ~n25366;
  assign n25369 = ~n34853 & ~n25366;
  assign n25370 = ~n24212 & n34853;
  assign n25371 = ~n34852 & n25370;
  assign n25372 = n34853 & n25366;
  assign n25373 = ~n24994 & n25371;
  assign n25374 = ~n25369 & ~n35003;
  assign n25375 = ~n25367 & ~n25368;
  assign n25376 = ~n25364 & ~n35004;
  assign n25377 = ~n25361 & ~n25362;
  assign n25378 = ~n16248 & ~n25377;
  assign n25379 = n15586 & ~n25378;
  assign n25380 = ~n25376 & ~n25378;
  assign n25381 = n15586 & n25380;
  assign n25382 = ~n25376 & n25379;
  assign n25383 = ~n25210 & ~n35005;
  assign n25384 = ~n15586 & ~n25380;
  assign n25385 = n14866 & ~n25384;
  assign n25386 = ~n25383 & n25385;
  assign n25387 = ~n24245 & ~n34856;
  assign n25388 = ~n24245 & ~n24994;
  assign n25389 = ~n34856 & n25388;
  assign n25390 = ~n24994 & n25387;
  assign n25391 = n34858 & ~n35006;
  assign n25392 = n24260 & n25388;
  assign n25393 = ~n34858 & n35006;
  assign n25394 = ~n24245 & n34858;
  assign n25395 = ~n34856 & n25394;
  assign n25396 = ~n24994 & n25395;
  assign n25397 = ~n34858 & ~n35006;
  assign n25398 = ~n25396 & ~n25397;
  assign n25399 = ~n25391 & ~n35007;
  assign n25400 = ~n25386 & ~n35008;
  assign n25401 = ~n25383 & ~n25384;
  assign n25402 = ~n14866 & ~n25401;
  assign n25403 = n14233 & ~n25402;
  assign n25404 = ~n25400 & ~n25402;
  assign n25405 = n14233 & n25404;
  assign n25406 = ~n25400 & n25403;
  assign n25407 = ~n25202 & ~n35009;
  assign n25408 = ~n14233 & ~n25404;
  assign n25409 = n13548 & ~n25408;
  assign n25410 = ~n25407 & n25409;
  assign n25411 = ~n25194 & ~n25410;
  assign n25412 = ~n25407 & ~n25408;
  assign n25413 = ~n13548 & ~n25412;
  assign n25414 = n12948 & ~n25413;
  assign n25415 = ~n25411 & ~n25413;
  assign n25416 = n12948 & n25415;
  assign n25417 = ~n25411 & n25414;
  assign n25418 = ~n25186 & ~n35010;
  assign n25419 = ~n12948 & ~n25415;
  assign n25420 = n12296 & ~n25419;
  assign n25421 = ~n25418 & n25420;
  assign n25422 = ~n24315 & ~n34868;
  assign n25423 = ~n24315 & ~n24994;
  assign n25424 = ~n34868 & n25423;
  assign n25425 = ~n24994 & n25422;
  assign n25426 = n24323 & ~n35011;
  assign n25427 = n24327 & n25423;
  assign n25428 = ~n24315 & n24323;
  assign n25429 = ~n34868 & n25428;
  assign n25430 = ~n24994 & n25429;
  assign n25431 = ~n24323 & ~n35011;
  assign n25432 = ~n25430 & ~n25431;
  assign n25433 = ~n25426 & ~n25427;
  assign n25434 = ~n25421 & ~n35012;
  assign n25435 = ~n25418 & ~n25419;
  assign n25436 = ~n12296 & ~n25435;
  assign n25437 = n11719 & ~n25436;
  assign n25438 = ~n25434 & ~n25436;
  assign n25439 = n11719 & n25438;
  assign n25440 = ~n25434 & n25437;
  assign n25441 = ~n25178 & ~n35013;
  assign n25442 = ~n11719 & ~n25438;
  assign n25443 = n11097 & ~n25442;
  assign n25444 = ~n25441 & n25443;
  assign n25445 = ~n25170 & ~n25444;
  assign n25446 = ~n25441 & ~n25442;
  assign n25447 = ~n11097 & ~n25446;
  assign n25448 = n10555 & ~n25447;
  assign n25449 = ~n25445 & ~n25447;
  assign n25450 = n10555 & n25449;
  assign n25451 = ~n25445 & n25448;
  assign n25452 = ~n25162 & ~n35014;
  assign n25453 = ~n10555 & ~n25449;
  assign n25454 = n9969 & ~n25453;
  assign n25455 = ~n25452 & n25454;
  assign n25456 = ~n24381 & ~n34877;
  assign n25457 = ~n24381 & ~n24994;
  assign n25458 = ~n34877 & n25457;
  assign n25459 = ~n24994 & n25456;
  assign n25460 = n24389 & ~n35015;
  assign n25461 = n24393 & n25457;
  assign n25462 = ~n24381 & n24389;
  assign n25463 = ~n34877 & n25462;
  assign n25464 = ~n24994 & n25463;
  assign n25465 = ~n24389 & ~n35015;
  assign n25466 = ~n25464 & ~n25465;
  assign n25467 = ~n25460 & ~n25461;
  assign n25468 = ~n25455 & ~n35016;
  assign n25469 = ~n25452 & ~n25453;
  assign n25470 = ~n9969 & ~n25469;
  assign n25471 = n9457 & ~n25470;
  assign n25472 = ~n25468 & ~n25470;
  assign n25473 = n9457 & n25472;
  assign n25474 = ~n25468 & n25471;
  assign n25475 = ~n25154 & ~n35017;
  assign n25476 = ~n9457 & ~n25472;
  assign n25477 = n8896 & ~n25476;
  assign n25478 = ~n25475 & n25477;
  assign n25479 = ~n25146 & ~n25478;
  assign n25480 = ~n25475 & ~n25476;
  assign n25481 = ~n8896 & ~n25480;
  assign n25482 = n8411 & ~n25481;
  assign n25483 = ~n25479 & ~n25481;
  assign n25484 = n8411 & n25483;
  assign n25485 = ~n25479 & n25482;
  assign n25486 = ~n25138 & ~n35018;
  assign n25487 = ~n8411 & ~n25483;
  assign n25488 = n7885 & ~n25487;
  assign n25489 = ~n25486 & n25488;
  assign n25490 = ~n24447 & ~n34886;
  assign n25491 = ~n24447 & ~n24994;
  assign n25492 = ~n34886 & n25491;
  assign n25493 = ~n24994 & n25490;
  assign n25494 = n24455 & ~n35019;
  assign n25495 = n24459 & n25491;
  assign n25496 = ~n24447 & n24455;
  assign n25497 = ~n34886 & n25496;
  assign n25498 = ~n24994 & n25497;
  assign n25499 = ~n24455 & ~n35019;
  assign n25500 = ~n25498 & ~n25499;
  assign n25501 = ~n25494 & ~n25495;
  assign n25502 = ~n25489 & ~n35020;
  assign n25503 = ~n25486 & ~n25487;
  assign n25504 = ~n7885 & ~n25503;
  assign n25505 = n7428 & ~n25504;
  assign n25506 = ~n25502 & ~n25504;
  assign n25507 = n7428 & n25506;
  assign n25508 = ~n25502 & n25505;
  assign n25509 = ~n25130 & ~n35021;
  assign n25510 = ~n7428 & ~n25506;
  assign n25511 = n6937 & ~n25510;
  assign n25512 = ~n25509 & n25511;
  assign n25513 = ~n25122 & ~n25512;
  assign n25514 = ~n25509 & ~n25510;
  assign n25515 = ~n6937 & ~n25514;
  assign n25516 = n6507 & ~n25515;
  assign n25517 = ~n25513 & ~n25515;
  assign n25518 = n6507 & n25517;
  assign n25519 = ~n25513 & n25516;
  assign n25520 = ~n25114 & ~n35022;
  assign n25521 = ~n6507 & ~n25517;
  assign n25522 = n6051 & ~n25521;
  assign n25523 = ~n25520 & n25522;
  assign n25524 = ~n24513 & ~n34895;
  assign n25525 = ~n24513 & ~n24994;
  assign n25526 = ~n34895 & n25525;
  assign n25527 = ~n24994 & n25524;
  assign n25528 = n24521 & ~n35023;
  assign n25529 = n24525 & n25525;
  assign n25530 = ~n24513 & n24521;
  assign n25531 = ~n34895 & n25530;
  assign n25532 = ~n24994 & n25531;
  assign n25533 = ~n24521 & ~n35023;
  assign n25534 = ~n25532 & ~n25533;
  assign n25535 = ~n25528 & ~n25529;
  assign n25536 = ~n25523 & ~n35024;
  assign n25537 = ~n25520 & ~n25521;
  assign n25538 = ~n6051 & ~n25537;
  assign n25539 = n5648 & ~n25538;
  assign n25540 = ~n25536 & ~n25538;
  assign n25541 = n5648 & n25540;
  assign n25542 = ~n25536 & n25539;
  assign n25543 = ~n25106 & ~n35025;
  assign n25544 = ~n5648 & ~n25540;
  assign n25545 = n5223 & ~n25544;
  assign n25546 = ~n25543 & n25545;
  assign n25547 = ~n25098 & ~n25546;
  assign n25548 = ~n25543 & ~n25544;
  assign n25549 = ~n5223 & ~n25548;
  assign n25550 = n4851 & ~n25549;
  assign n25551 = ~n25547 & ~n25549;
  assign n25552 = n4851 & n25551;
  assign n25553 = ~n25547 & n25550;
  assign n25554 = ~n25090 & ~n35026;
  assign n25555 = ~n4851 & ~n25551;
  assign n25556 = n4461 & ~n25555;
  assign n25557 = ~n25554 & n25556;
  assign n25558 = ~n24579 & ~n34904;
  assign n25559 = ~n24579 & ~n24994;
  assign n25560 = ~n34904 & n25559;
  assign n25561 = ~n24994 & n25558;
  assign n25562 = n24587 & ~n35027;
  assign n25563 = n24591 & n25559;
  assign n25564 = ~n24579 & n24587;
  assign n25565 = ~n34904 & n25564;
  assign n25566 = ~n24994 & n25565;
  assign n25567 = ~n24587 & ~n35027;
  assign n25568 = ~n25566 & ~n25567;
  assign n25569 = ~n25562 & ~n25563;
  assign n25570 = ~n25557 & ~n35028;
  assign n25571 = ~n25554 & ~n25555;
  assign n25572 = ~n4461 & ~n25571;
  assign n25573 = n4115 & ~n25572;
  assign n25574 = ~n25570 & ~n25572;
  assign n25575 = n4115 & n25574;
  assign n25576 = ~n25570 & n25573;
  assign n25577 = ~n25082 & ~n35029;
  assign n25578 = ~n4115 & ~n25574;
  assign n25579 = n3754 & ~n25578;
  assign n25580 = ~n25577 & n25579;
  assign n25581 = ~n25074 & ~n25580;
  assign n25582 = ~n25577 & ~n25578;
  assign n25583 = ~n3754 & ~n25582;
  assign n25584 = n3444 & ~n25583;
  assign n25585 = ~n25581 & ~n25583;
  assign n25586 = n3444 & n25585;
  assign n25587 = ~n25581 & n25584;
  assign n25588 = ~n25066 & ~n35030;
  assign n25589 = ~n3444 & ~n25585;
  assign n25590 = n3116 & ~n25589;
  assign n25591 = ~n25588 & n25590;
  assign n25592 = ~n24645 & ~n34913;
  assign n25593 = ~n24645 & ~n24994;
  assign n25594 = ~n34913 & n25593;
  assign n25595 = ~n24994 & n25592;
  assign n25596 = n24653 & ~n35031;
  assign n25597 = n24657 & n25593;
  assign n25598 = ~n24645 & n24653;
  assign n25599 = ~n34913 & n25598;
  assign n25600 = ~n24994 & n25599;
  assign n25601 = ~n24653 & ~n35031;
  assign n25602 = ~n25600 & ~n25601;
  assign n25603 = ~n25596 & ~n25597;
  assign n25604 = ~n25591 & ~n35032;
  assign n25605 = ~n25588 & ~n25589;
  assign n25606 = ~n3116 & ~n25605;
  assign n25607 = n2833 & ~n25606;
  assign n25608 = ~n25604 & ~n25606;
  assign n25609 = n2833 & n25608;
  assign n25610 = ~n25604 & n25607;
  assign n25611 = ~n25058 & ~n35033;
  assign n25612 = ~n2833 & ~n25608;
  assign n25613 = n2536 & ~n25612;
  assign n25614 = ~n25611 & n25613;
  assign n25615 = ~n25050 & ~n25614;
  assign n25616 = ~n25611 & ~n25612;
  assign n25617 = ~n2536 & ~n25616;
  assign n25618 = n2283 & ~n25617;
  assign n25619 = ~n25615 & ~n25617;
  assign n25620 = n2283 & n25619;
  assign n25621 = ~n25615 & n25618;
  assign n25622 = ~n25042 & ~n35034;
  assign n25623 = ~n2283 & ~n25619;
  assign n25624 = n2021 & ~n25623;
  assign n25625 = ~n25622 & n25624;
  assign n25626 = ~n24711 & ~n34922;
  assign n25627 = ~n24711 & ~n24994;
  assign n25628 = ~n34922 & n25627;
  assign n25629 = ~n24994 & n25626;
  assign n25630 = n24719 & ~n35035;
  assign n25631 = n24723 & n25627;
  assign n25632 = ~n24711 & n24719;
  assign n25633 = ~n34922 & n25632;
  assign n25634 = ~n24994 & n25633;
  assign n25635 = ~n24719 & ~n35035;
  assign n25636 = ~n25634 & ~n25635;
  assign n25637 = ~n25630 & ~n25631;
  assign n25638 = ~n25625 & ~n35036;
  assign n25639 = ~n25622 & ~n25623;
  assign n25640 = ~n2021 & ~n25639;
  assign n25641 = n1796 & ~n25640;
  assign n25642 = ~n25638 & ~n25640;
  assign n25643 = n1796 & n25642;
  assign n25644 = ~n25638 & n25641;
  assign n25645 = ~n25034 & ~n35037;
  assign n25646 = ~n1796 & ~n25642;
  assign n25647 = n1567 & ~n25646;
  assign n25648 = ~n25645 & n25647;
  assign n25649 = ~n25026 & ~n25648;
  assign n25650 = ~n25645 & ~n25646;
  assign n25651 = ~n1567 & ~n25650;
  assign n25652 = n1374 & ~n25651;
  assign n25653 = ~n25649 & ~n25651;
  assign n25654 = n1374 & n25653;
  assign n25655 = ~n25649 & n25652;
  assign n25656 = ~n25018 & ~n35038;
  assign n25657 = ~n1374 & ~n25653;
  assign n25658 = n1179 & ~n25657;
  assign n25659 = ~n25656 & n25658;
  assign n25660 = ~n24777 & ~n34931;
  assign n25661 = ~n24777 & ~n24994;
  assign n25662 = ~n34931 & n25661;
  assign n25663 = ~n24994 & n25660;
  assign n25664 = n24785 & ~n35039;
  assign n25665 = n24789 & n25661;
  assign n25666 = ~n24777 & n24785;
  assign n25667 = ~n34931 & n25666;
  assign n25668 = ~n24994 & n25667;
  assign n25669 = ~n24785 & ~n35039;
  assign n25670 = ~n25668 & ~n25669;
  assign n25671 = ~n25664 & ~n25665;
  assign n25672 = ~n25659 & ~n35040;
  assign n25673 = ~n25656 & ~n25657;
  assign n25674 = ~n1179 & ~n25673;
  assign n25675 = n1016 & ~n25674;
  assign n25676 = ~n25672 & ~n25674;
  assign n25677 = n1016 & n25676;
  assign n25678 = ~n25672 & n25675;
  assign n25679 = ~n25010 & ~n35041;
  assign n25680 = ~n1016 & ~n25676;
  assign n25681 = n855 & ~n25680;
  assign n25682 = ~n25679 & n25681;
  assign n25683 = ~n25002 & ~n25682;
  assign n25684 = ~n25679 & ~n25680;
  assign n25685 = ~n855 & ~n25684;
  assign n25686 = n720 & ~n25685;
  assign n25687 = ~n25683 & ~n25685;
  assign n25688 = n720 & n25687;
  assign n25689 = ~n25683 & n25686;
  assign n25690 = ~n24826 & ~n24828;
  assign n25691 = ~n24994 & n25690;
  assign n25692 = ~n34937 & n25691;
  assign n25693 = n34937 & ~n25691;
  assign n25694 = ~n24828 & n34937;
  assign n25695 = ~n24826 & n25694;
  assign n25696 = ~n24994 & n25695;
  assign n25697 = ~n34937 & ~n25691;
  assign n25698 = ~n25696 & ~n25697;
  assign n25699 = ~n25692 & ~n25693;
  assign n25700 = ~n35042 & ~n35043;
  assign n25701 = ~n720 & ~n25687;
  assign n25702 = ~n25700 & ~n25701;
  assign n25703 = ~n592 & ~n25702;
  assign n25704 = ~n24841 & ~n34939;
  assign n25705 = ~n24994 & n25704;
  assign n25706 = n34938 & ~n25705;
  assign n25707 = ~n34938 & n25705;
  assign n25708 = ~n24841 & n34938;
  assign n25709 = ~n34939 & n25708;
  assign n25710 = ~n24994 & n25709;
  assign n25711 = ~n34938 & ~n25705;
  assign n25712 = ~n25710 & ~n25711;
  assign n25713 = ~n25706 & ~n25707;
  assign n25714 = n592 & ~n25701;
  assign n25715 = ~n25700 & n25714;
  assign n25716 = ~n35044 & ~n25715;
  assign n25717 = ~n25703 & ~n25716;
  assign n25718 = ~n487 & ~n25717;
  assign n25719 = ~n24857 & ~n24859;
  assign n25720 = ~n24994 & n25719;
  assign n25721 = ~n34941 & ~n25720;
  assign n25722 = ~n24859 & n34941;
  assign n25723 = ~n24857 & n25722;
  assign n25724 = n34941 & n25720;
  assign n25725 = ~n24994 & n25723;
  assign n25726 = ~n25721 & ~n35045;
  assign n25727 = n487 & ~n25703;
  assign n25728 = n487 & n25717;
  assign n25729 = ~n25716 & n25727;
  assign n25730 = ~n25726 & ~n35046;
  assign n25731 = ~n25718 & ~n25730;
  assign n25732 = ~n393 & ~n25731;
  assign n25733 = n393 & ~n25718;
  assign n25734 = ~n25730 & n25733;
  assign n25735 = ~n24874 & ~n34943;
  assign n25736 = ~n24874 & ~n24994;
  assign n25737 = ~n34943 & n25736;
  assign n25738 = ~n24994 & n25735;
  assign n25739 = n24882 & ~n35047;
  assign n25740 = n24886 & n25736;
  assign n25741 = ~n24874 & n24882;
  assign n25742 = ~n34943 & n25741;
  assign n25743 = ~n24994 & n25742;
  assign n25744 = ~n24882 & ~n35047;
  assign n25745 = ~n25743 & ~n25744;
  assign n25746 = ~n25739 & ~n25740;
  assign n25747 = ~n25734 & ~n35048;
  assign n25748 = ~n25732 & ~n25747;
  assign n25749 = ~n321 & ~n25748;
  assign n25750 = ~n24888 & ~n24890;
  assign n25751 = ~n24994 & n25750;
  assign n25752 = ~n34945 & ~n25751;
  assign n25753 = ~n24890 & n34945;
  assign n25754 = ~n24888 & n25753;
  assign n25755 = n34945 & n25751;
  assign n25756 = ~n24994 & n25754;
  assign n25757 = ~n25752 & ~n35049;
  assign n25758 = n321 & ~n25732;
  assign n25759 = n321 & n25748;
  assign n25760 = ~n25747 & n25758;
  assign n25761 = ~n25757 & ~n35050;
  assign n25762 = ~n25749 & ~n25761;
  assign n25763 = ~n263 & ~n25762;
  assign n25764 = n263 & ~n25749;
  assign n25765 = ~n25761 & n25764;
  assign n25766 = ~n24905 & ~n34947;
  assign n25767 = ~n24905 & ~n24994;
  assign n25768 = ~n34947 & n25767;
  assign n25769 = ~n24994 & n25766;
  assign n25770 = n24913 & ~n35051;
  assign n25771 = n24917 & n25767;
  assign n25772 = ~n24905 & n24913;
  assign n25773 = ~n34947 & n25772;
  assign n25774 = ~n24994 & n25773;
  assign n25775 = ~n24913 & ~n35051;
  assign n25776 = ~n25774 & ~n25775;
  assign n25777 = ~n25770 & ~n25771;
  assign n25778 = ~n25765 & ~n35052;
  assign n25779 = ~n25763 & ~n25778;
  assign n25780 = ~n214 & ~n25779;
  assign n25781 = ~n24919 & ~n24921;
  assign n25782 = ~n24994 & n25781;
  assign n25783 = ~n34949 & ~n25782;
  assign n25784 = ~n24921 & n34949;
  assign n25785 = ~n24919 & n25784;
  assign n25786 = n34949 & n25782;
  assign n25787 = ~n24994 & n25785;
  assign n25788 = ~n25783 & ~n35053;
  assign n25789 = n214 & ~n25763;
  assign n25790 = n214 & n25779;
  assign n25791 = ~n25778 & n25789;
  assign n25792 = ~n25788 & ~n35054;
  assign n25793 = ~n25780 & ~n25792;
  assign n25794 = ~n197 & ~n25793;
  assign n25795 = ~n24936 & ~n34950;
  assign n25796 = ~n24994 & n25795;
  assign n25797 = ~n34952 & ~n25796;
  assign n25798 = ~n24936 & n34952;
  assign n25799 = ~n34950 & n25798;
  assign n25800 = n34952 & n25796;
  assign n25801 = ~n24994 & n25799;
  assign n25802 = ~n25797 & ~n35055;
  assign n25803 = n197 & ~n25780;
  assign n25804 = ~n25792 & n25803;
  assign n25805 = ~n25802 & ~n25804;
  assign n25806 = ~n25794 & ~n25805;
  assign n25807 = ~n24954 & ~n24956;
  assign n25808 = ~n24994 & n25807;
  assign n25809 = ~n34954 & ~n25808;
  assign n25810 = ~n24956 & n34954;
  assign n25811 = ~n24954 & n25810;
  assign n25812 = n34954 & n25808;
  assign n25813 = ~n24994 & n25811;
  assign n25814 = ~n25809 & ~n35056;
  assign n25815 = ~n24970 & ~n24978;
  assign n25816 = ~n24978 & ~n24994;
  assign n25817 = ~n24970 & n25816;
  assign n25818 = ~n24994 & n25815;
  assign n25819 = ~n34957 & ~n35057;
  assign n25820 = ~n25814 & n25819;
  assign n25821 = ~n25806 & n25820;
  assign n25822 = n193 & ~n25821;
  assign n25823 = ~n25794 & n25814;
  assign n25824 = n25806 & n25814;
  assign n25825 = ~n25805 & n25823;
  assign n25826 = n24970 & ~n25816;
  assign n25827 = ~n193 & ~n25815;
  assign n25828 = ~n25826 & n25827;
  assign n25829 = ~n35058 & ~n25828;
  assign n25830 = ~n25822 & n25829;
  assign n25831 = pi12  & ~n25830;
  assign n25832 = ~pi10  & ~pi11 ;
  assign n25833 = ~pi12  & n25832;
  assign n25834 = ~n25831 & ~n25833;
  assign n25835 = ~n24994 & ~n25834;
  assign n25836 = ~pi12  & ~n25830;
  assign n25837 = pi13  & ~n25836;
  assign n25838 = ~pi13  & n25836;
  assign n25839 = n25256 & ~n25830;
  assign n25840 = ~n25837 & ~n35059;
  assign n25841 = ~n34832 & ~n34991;
  assign n25842 = ~n24055 & n25841;
  assign n25843 = ~n24074 & n25842;
  assign n25844 = ~n34834 & n25843;
  assign n25845 = n24060 & n24076;
  assign n25846 = ~n24068 & n25844;
  assign n25847 = ~n25833 & ~n35060;
  assign n25848 = ~n24992 & n25847;
  assign n25849 = ~n34957 & n25848;
  assign n25850 = ~n24986 & n25849;
  assign n25851 = n24994 & n25834;
  assign n25852 = ~n25831 & n25850;
  assign n25853 = n25840 & ~n35061;
  assign n25854 = ~n25835 & ~n25853;
  assign n25855 = ~n24076 & ~n25854;
  assign n25856 = n24076 & ~n25835;
  assign n25857 = ~n25853 & n25856;
  assign n25858 = ~n24994 & ~n25828;
  assign n25859 = ~n35058 & n25858;
  assign n25860 = ~n25822 & n25859;
  assign n25861 = ~n35059 & ~n25860;
  assign n25862 = pi14  & ~n25861;
  assign n25863 = ~pi14  & ~n25860;
  assign n25864 = ~pi14  & n25861;
  assign n25865 = ~n35059 & n25863;
  assign n25866 = ~n25862 & ~n35062;
  assign n25867 = ~n25857 & ~n25866;
  assign n25868 = ~n25855 & ~n25867;
  assign n25869 = ~n23269 & ~n25868;
  assign n25870 = n23269 & ~n25855;
  assign n25871 = ~n25867 & n25870;
  assign n25872 = n23269 & n25868;
  assign n25873 = ~n34992 & ~n25274;
  assign n25874 = ~n25830 & n25873;
  assign n25875 = n25272 & ~n25874;
  assign n25876 = ~n25272 & n25873;
  assign n25877 = ~n25272 & n25874;
  assign n25878 = ~n25830 & n25876;
  assign n25879 = ~n25875 & ~n35064;
  assign n25880 = ~n35063 & ~n25879;
  assign n25881 = ~n25869 & ~n25880;
  assign n25882 = ~n22386 & ~n25881;
  assign n25883 = n22386 & ~n25869;
  assign n25884 = ~n25880 & n25883;
  assign n25885 = ~n34993 & ~n25280;
  assign n25886 = ~n25280 & ~n25830;
  assign n25887 = ~n34993 & n25886;
  assign n25888 = ~n25830 & n25885;
  assign n25889 = n25254 & ~n35065;
  assign n25890 = n25279 & n25886;
  assign n25891 = n25254 & ~n34993;
  assign n25892 = ~n25280 & n25891;
  assign n25893 = ~n25830 & n25892;
  assign n25894 = ~n25254 & ~n35065;
  assign n25895 = ~n25893 & ~n25894;
  assign n25896 = ~n25889 & ~n25890;
  assign n25897 = ~n25884 & ~n35066;
  assign n25898 = ~n25882 & ~n25897;
  assign n25899 = ~n21612 & ~n25898;
  assign n25900 = n21612 & ~n25882;
  assign n25901 = ~n25897 & n25900;
  assign n25902 = n21612 & n25898;
  assign n25903 = ~n25282 & ~n25292;
  assign n25904 = ~n25830 & n25903;
  assign n25905 = ~n25289 & ~n25904;
  assign n25906 = n25289 & ~n25292;
  assign n25907 = ~n25282 & n25906;
  assign n25908 = n25289 & n25904;
  assign n25909 = ~n25830 & n25907;
  assign n25910 = n25289 & ~n25904;
  assign n25911 = ~n25289 & n25904;
  assign n25912 = ~n25910 & ~n25911;
  assign n25913 = ~n25905 & ~n35068;
  assign n25914 = ~n35067 & n35069;
  assign n25915 = ~n25899 & ~n25914;
  assign n25916 = ~n20762 & ~n25915;
  assign n25917 = n20762 & ~n25899;
  assign n25918 = ~n25914 & n25917;
  assign n25919 = ~n34995 & ~n25298;
  assign n25920 = ~n25298 & ~n25830;
  assign n25921 = ~n34995 & n25920;
  assign n25922 = ~n25830 & n25919;
  assign n25923 = n25242 & ~n35070;
  assign n25924 = n25297 & n25920;
  assign n25925 = n25242 & ~n34995;
  assign n25926 = ~n25298 & n25925;
  assign n25927 = ~n25830 & n25926;
  assign n25928 = ~n25242 & ~n35070;
  assign n25929 = ~n25927 & ~n25928;
  assign n25930 = ~n25923 & ~n25924;
  assign n25931 = ~n25918 & ~n35071;
  assign n25932 = ~n25916 & ~n25931;
  assign n25933 = ~n20011 & ~n25932;
  assign n25934 = n20011 & ~n25916;
  assign n25935 = ~n25931 & n25934;
  assign n25936 = n20011 & n25932;
  assign n25937 = ~n25300 & ~n25314;
  assign n25938 = ~n25830 & n25937;
  assign n25939 = ~n34997 & ~n25938;
  assign n25940 = n34997 & n25938;
  assign n25941 = ~n34997 & ~n25314;
  assign n25942 = ~n25300 & n25941;
  assign n25943 = ~n25830 & n25942;
  assign n25944 = n34997 & ~n25938;
  assign n25945 = ~n25943 & ~n25944;
  assign n25946 = ~n25939 & ~n25940;
  assign n25947 = ~n35072 & ~n35073;
  assign n25948 = ~n25933 & ~n25947;
  assign n25949 = ~n19190 & ~n25948;
  assign n25950 = n19190 & ~n25933;
  assign n25951 = ~n25947 & n25950;
  assign n25952 = ~n34998 & ~n25320;
  assign n25953 = ~n25320 & ~n25830;
  assign n25954 = ~n34998 & n25953;
  assign n25955 = ~n25830 & n25952;
  assign n25956 = n25234 & ~n35074;
  assign n25957 = n25319 & n25953;
  assign n25958 = n25234 & ~n34998;
  assign n25959 = ~n25320 & n25958;
  assign n25960 = ~n25830 & n25959;
  assign n25961 = ~n25234 & ~n35074;
  assign n25962 = ~n25960 & ~n25961;
  assign n25963 = ~n25956 & ~n25957;
  assign n25964 = ~n25951 & ~n35075;
  assign n25965 = ~n25949 & ~n25964;
  assign n25966 = ~n18472 & ~n25965;
  assign n25967 = n18472 & ~n25949;
  assign n25968 = ~n25964 & n25967;
  assign n25969 = n18472 & n25965;
  assign n25970 = ~n25322 & ~n25335;
  assign n25971 = ~n25830 & n25970;
  assign n25972 = ~n34999 & n25971;
  assign n25973 = n34999 & ~n25971;
  assign n25974 = n34999 & ~n25335;
  assign n25975 = ~n25322 & n25974;
  assign n25976 = ~n25830 & n25975;
  assign n25977 = ~n34999 & ~n25971;
  assign n25978 = ~n25976 & ~n25977;
  assign n25979 = ~n25972 & ~n25973;
  assign n25980 = ~n35076 & ~n35077;
  assign n25981 = ~n25966 & ~n25980;
  assign n25982 = ~n17690 & ~n25981;
  assign n25983 = n17690 & ~n25966;
  assign n25984 = ~n25980 & n25983;
  assign n25985 = ~n35000 & ~n25341;
  assign n25986 = ~n25341 & ~n25830;
  assign n25987 = ~n35000 & n25986;
  assign n25988 = ~n25830 & n25985;
  assign n25989 = n25226 & ~n35078;
  assign n25990 = n25340 & n25986;
  assign n25991 = n25226 & ~n35000;
  assign n25992 = ~n25341 & n25991;
  assign n25993 = ~n25830 & n25992;
  assign n25994 = ~n25226 & ~n35078;
  assign n25995 = ~n25993 & ~n25994;
  assign n25996 = ~n25989 & ~n25990;
  assign n25997 = ~n25984 & ~n35079;
  assign n25998 = ~n25982 & ~n25997;
  assign n25999 = ~n17001 & ~n25998;
  assign n26000 = n17001 & ~n25982;
  assign n26001 = ~n25997 & n26000;
  assign n26002 = n17001 & n25998;
  assign n26003 = ~n25343 & ~n25356;
  assign n26004 = ~n25830 & n26003;
  assign n26005 = ~n35001 & n26004;
  assign n26006 = n35001 & ~n26004;
  assign n26007 = ~n35001 & ~n26004;
  assign n26008 = n35001 & ~n25356;
  assign n26009 = ~n25343 & n26008;
  assign n26010 = n35001 & n26004;
  assign n26011 = ~n25830 & n26009;
  assign n26012 = ~n26007 & ~n35081;
  assign n26013 = ~n26005 & ~n26006;
  assign n26014 = ~n35080 & ~n35082;
  assign n26015 = ~n25999 & ~n26014;
  assign n26016 = ~n16248 & ~n26015;
  assign n26017 = n16248 & ~n25999;
  assign n26018 = ~n26014 & n26017;
  assign n26019 = ~n35002 & ~n25362;
  assign n26020 = ~n25362 & ~n25830;
  assign n26021 = ~n35002 & n26020;
  assign n26022 = ~n25830 & n26019;
  assign n26023 = n25218 & ~n35083;
  assign n26024 = n25361 & n26020;
  assign n26025 = n25218 & ~n35002;
  assign n26026 = ~n25362 & n26025;
  assign n26027 = ~n25830 & n26026;
  assign n26028 = ~n25218 & ~n35083;
  assign n26029 = ~n26027 & ~n26028;
  assign n26030 = ~n26023 & ~n26024;
  assign n26031 = ~n26018 & ~n35084;
  assign n26032 = ~n26016 & ~n26031;
  assign n26033 = ~n15586 & ~n26032;
  assign n26034 = n15586 & ~n26016;
  assign n26035 = ~n26031 & n26034;
  assign n26036 = n15586 & n26032;
  assign n26037 = ~n25364 & ~n25378;
  assign n26038 = ~n25378 & ~n25830;
  assign n26039 = ~n25364 & n26038;
  assign n26040 = ~n25830 & n26037;
  assign n26041 = n35004 & ~n35086;
  assign n26042 = n25376 & n26038;
  assign n26043 = ~n35004 & n35086;
  assign n26044 = n35004 & ~n25378;
  assign n26045 = ~n25364 & n26044;
  assign n26046 = ~n25830 & n26045;
  assign n26047 = ~n35004 & ~n35086;
  assign n26048 = ~n26046 & ~n26047;
  assign n26049 = ~n26041 & ~n35087;
  assign n26050 = ~n35085 & ~n35088;
  assign n26051 = ~n26033 & ~n26050;
  assign n26052 = ~n14866 & ~n26051;
  assign n26053 = n14866 & ~n26033;
  assign n26054 = ~n26050 & n26053;
  assign n26055 = ~n35005 & ~n25384;
  assign n26056 = ~n25384 & ~n25830;
  assign n26057 = ~n35005 & n26056;
  assign n26058 = ~n25830 & n26055;
  assign n26059 = n25210 & ~n35089;
  assign n26060 = n25383 & n26056;
  assign n26061 = n25210 & ~n35005;
  assign n26062 = ~n25384 & n26061;
  assign n26063 = ~n25830 & n26062;
  assign n26064 = ~n25210 & ~n35089;
  assign n26065 = ~n26063 & ~n26064;
  assign n26066 = ~n26059 & ~n26060;
  assign n26067 = ~n26054 & ~n35090;
  assign n26068 = ~n26052 & ~n26067;
  assign n26069 = ~n14233 & ~n26068;
  assign n26070 = ~n25386 & ~n25402;
  assign n26071 = ~n25830 & n26070;
  assign n26072 = ~n35008 & ~n26071;
  assign n26073 = n35008 & ~n25402;
  assign n26074 = ~n25386 & n26073;
  assign n26075 = n35008 & n26071;
  assign n26076 = ~n25830 & n26074;
  assign n26077 = ~n26072 & ~n35091;
  assign n26078 = n14233 & ~n26052;
  assign n26079 = ~n26067 & n26078;
  assign n26080 = n14233 & n26068;
  assign n26081 = ~n26077 & ~n35092;
  assign n26082 = ~n26069 & ~n26081;
  assign n26083 = ~n13548 & ~n26082;
  assign n26084 = n13548 & ~n26069;
  assign n26085 = ~n26081 & n26084;
  assign n26086 = ~n35009 & ~n25408;
  assign n26087 = ~n25408 & ~n25830;
  assign n26088 = ~n35009 & n26087;
  assign n26089 = ~n25830 & n26086;
  assign n26090 = n25202 & ~n35093;
  assign n26091 = n25407 & n26087;
  assign n26092 = n25202 & ~n35009;
  assign n26093 = ~n25408 & n26092;
  assign n26094 = ~n25830 & n26093;
  assign n26095 = ~n25202 & ~n35093;
  assign n26096 = ~n26094 & ~n26095;
  assign n26097 = ~n26090 & ~n26091;
  assign n26098 = ~n26085 & ~n35094;
  assign n26099 = ~n26083 & ~n26098;
  assign n26100 = ~n12948 & ~n26099;
  assign n26101 = n12948 & ~n26083;
  assign n26102 = ~n26098 & n26101;
  assign n26103 = n12948 & n26099;
  assign n26104 = ~n25410 & ~n25413;
  assign n26105 = ~n25413 & ~n25830;
  assign n26106 = ~n25410 & n26105;
  assign n26107 = ~n25830 & n26104;
  assign n26108 = n25194 & ~n35096;
  assign n26109 = n25411 & n26105;
  assign n26110 = n25194 & ~n25413;
  assign n26111 = ~n25410 & n26110;
  assign n26112 = ~n25830 & n26111;
  assign n26113 = ~n25194 & ~n35096;
  assign n26114 = ~n26112 & ~n26113;
  assign n26115 = ~n26108 & ~n26109;
  assign n26116 = ~n35095 & ~n35097;
  assign n26117 = ~n26100 & ~n26116;
  assign n26118 = ~n12296 & ~n26117;
  assign n26119 = n12296 & ~n26100;
  assign n26120 = ~n26116 & n26119;
  assign n26121 = ~n35010 & ~n25419;
  assign n26122 = ~n25419 & ~n25830;
  assign n26123 = ~n35010 & n26122;
  assign n26124 = ~n25830 & n26121;
  assign n26125 = n25186 & ~n35098;
  assign n26126 = n25418 & n26122;
  assign n26127 = n25186 & ~n35010;
  assign n26128 = ~n25419 & n26127;
  assign n26129 = ~n25830 & n26128;
  assign n26130 = ~n25186 & ~n35098;
  assign n26131 = ~n26129 & ~n26130;
  assign n26132 = ~n26125 & ~n26126;
  assign n26133 = ~n26120 & ~n35099;
  assign n26134 = ~n26118 & ~n26133;
  assign n26135 = ~n11719 & ~n26134;
  assign n26136 = ~n25421 & ~n25436;
  assign n26137 = ~n25830 & n26136;
  assign n26138 = ~n35012 & ~n26137;
  assign n26139 = n35012 & ~n25436;
  assign n26140 = ~n25421 & n26139;
  assign n26141 = n35012 & n26137;
  assign n26142 = ~n25830 & n26140;
  assign n26143 = ~n26138 & ~n35100;
  assign n26144 = n11719 & ~n26118;
  assign n26145 = ~n26133 & n26144;
  assign n26146 = n11719 & n26134;
  assign n26147 = ~n26143 & ~n35101;
  assign n26148 = ~n26135 & ~n26147;
  assign n26149 = ~n11097 & ~n26148;
  assign n26150 = n11097 & ~n26135;
  assign n26151 = ~n26147 & n26150;
  assign n26152 = ~n35013 & ~n25442;
  assign n26153 = ~n25442 & ~n25830;
  assign n26154 = ~n35013 & n26153;
  assign n26155 = ~n25830 & n26152;
  assign n26156 = n25178 & ~n35102;
  assign n26157 = n25441 & n26153;
  assign n26158 = n25178 & ~n35013;
  assign n26159 = ~n25442 & n26158;
  assign n26160 = ~n25830 & n26159;
  assign n26161 = ~n25178 & ~n35102;
  assign n26162 = ~n26160 & ~n26161;
  assign n26163 = ~n26156 & ~n26157;
  assign n26164 = ~n26151 & ~n35103;
  assign n26165 = ~n26149 & ~n26164;
  assign n26166 = ~n10555 & ~n26165;
  assign n26167 = n10555 & ~n26149;
  assign n26168 = ~n26164 & n26167;
  assign n26169 = n10555 & n26165;
  assign n26170 = ~n25444 & ~n25447;
  assign n26171 = ~n25447 & ~n25830;
  assign n26172 = ~n25444 & n26171;
  assign n26173 = ~n25830 & n26170;
  assign n26174 = n25170 & ~n35105;
  assign n26175 = n25445 & n26171;
  assign n26176 = n25170 & ~n25447;
  assign n26177 = ~n25444 & n26176;
  assign n26178 = ~n25830 & n26177;
  assign n26179 = ~n25170 & ~n35105;
  assign n26180 = ~n26178 & ~n26179;
  assign n26181 = ~n26174 & ~n26175;
  assign n26182 = ~n35104 & ~n35106;
  assign n26183 = ~n26166 & ~n26182;
  assign n26184 = ~n9969 & ~n26183;
  assign n26185 = n9969 & ~n26166;
  assign n26186 = ~n26182 & n26185;
  assign n26187 = ~n35014 & ~n25453;
  assign n26188 = ~n25453 & ~n25830;
  assign n26189 = ~n35014 & n26188;
  assign n26190 = ~n25830 & n26187;
  assign n26191 = n25162 & ~n35107;
  assign n26192 = n25452 & n26188;
  assign n26193 = n25162 & ~n35014;
  assign n26194 = ~n25453 & n26193;
  assign n26195 = ~n25830 & n26194;
  assign n26196 = ~n25162 & ~n35107;
  assign n26197 = ~n26195 & ~n26196;
  assign n26198 = ~n26191 & ~n26192;
  assign n26199 = ~n26186 & ~n35108;
  assign n26200 = ~n26184 & ~n26199;
  assign n26201 = ~n9457 & ~n26200;
  assign n26202 = ~n25455 & ~n25470;
  assign n26203 = ~n25830 & n26202;
  assign n26204 = ~n35016 & ~n26203;
  assign n26205 = n35016 & ~n25470;
  assign n26206 = ~n25455 & n26205;
  assign n26207 = n35016 & n26203;
  assign n26208 = ~n25830 & n26206;
  assign n26209 = ~n26204 & ~n35109;
  assign n26210 = n9457 & ~n26184;
  assign n26211 = ~n26199 & n26210;
  assign n26212 = n9457 & n26200;
  assign n26213 = ~n26209 & ~n35110;
  assign n26214 = ~n26201 & ~n26213;
  assign n26215 = ~n8896 & ~n26214;
  assign n26216 = n8896 & ~n26201;
  assign n26217 = ~n26213 & n26216;
  assign n26218 = ~n35017 & ~n25476;
  assign n26219 = ~n25476 & ~n25830;
  assign n26220 = ~n35017 & n26219;
  assign n26221 = ~n25830 & n26218;
  assign n26222 = n25154 & ~n35111;
  assign n26223 = n25475 & n26219;
  assign n26224 = n25154 & ~n35017;
  assign n26225 = ~n25476 & n26224;
  assign n26226 = ~n25830 & n26225;
  assign n26227 = ~n25154 & ~n35111;
  assign n26228 = ~n26226 & ~n26227;
  assign n26229 = ~n26222 & ~n26223;
  assign n26230 = ~n26217 & ~n35112;
  assign n26231 = ~n26215 & ~n26230;
  assign n26232 = ~n8411 & ~n26231;
  assign n26233 = n8411 & ~n26215;
  assign n26234 = ~n26230 & n26233;
  assign n26235 = n8411 & n26231;
  assign n26236 = ~n25478 & ~n25481;
  assign n26237 = ~n25481 & ~n25830;
  assign n26238 = ~n25478 & n26237;
  assign n26239 = ~n25830 & n26236;
  assign n26240 = n25146 & ~n35114;
  assign n26241 = n25479 & n26237;
  assign n26242 = n25146 & ~n25481;
  assign n26243 = ~n25478 & n26242;
  assign n26244 = ~n25830 & n26243;
  assign n26245 = ~n25146 & ~n35114;
  assign n26246 = ~n26244 & ~n26245;
  assign n26247 = ~n26240 & ~n26241;
  assign n26248 = ~n35113 & ~n35115;
  assign n26249 = ~n26232 & ~n26248;
  assign n26250 = ~n7885 & ~n26249;
  assign n26251 = n7885 & ~n26232;
  assign n26252 = ~n26248 & n26251;
  assign n26253 = ~n35018 & ~n25487;
  assign n26254 = ~n25487 & ~n25830;
  assign n26255 = ~n35018 & n26254;
  assign n26256 = ~n25830 & n26253;
  assign n26257 = n25138 & ~n35116;
  assign n26258 = n25486 & n26254;
  assign n26259 = n25138 & ~n35018;
  assign n26260 = ~n25487 & n26259;
  assign n26261 = ~n25830 & n26260;
  assign n26262 = ~n25138 & ~n35116;
  assign n26263 = ~n26261 & ~n26262;
  assign n26264 = ~n26257 & ~n26258;
  assign n26265 = ~n26252 & ~n35117;
  assign n26266 = ~n26250 & ~n26265;
  assign n26267 = ~n7428 & ~n26266;
  assign n26268 = ~n25489 & ~n25504;
  assign n26269 = ~n25830 & n26268;
  assign n26270 = ~n35020 & ~n26269;
  assign n26271 = n35020 & ~n25504;
  assign n26272 = ~n25489 & n26271;
  assign n26273 = n35020 & n26269;
  assign n26274 = ~n25830 & n26272;
  assign n26275 = ~n26270 & ~n35118;
  assign n26276 = n7428 & ~n26250;
  assign n26277 = ~n26265 & n26276;
  assign n26278 = n7428 & n26266;
  assign n26279 = ~n26275 & ~n35119;
  assign n26280 = ~n26267 & ~n26279;
  assign n26281 = ~n6937 & ~n26280;
  assign n26282 = n6937 & ~n26267;
  assign n26283 = ~n26279 & n26282;
  assign n26284 = ~n35021 & ~n25510;
  assign n26285 = ~n25510 & ~n25830;
  assign n26286 = ~n35021 & n26285;
  assign n26287 = ~n25830 & n26284;
  assign n26288 = n25130 & ~n35120;
  assign n26289 = n25509 & n26285;
  assign n26290 = n25130 & ~n35021;
  assign n26291 = ~n25510 & n26290;
  assign n26292 = ~n25830 & n26291;
  assign n26293 = ~n25130 & ~n35120;
  assign n26294 = ~n26292 & ~n26293;
  assign n26295 = ~n26288 & ~n26289;
  assign n26296 = ~n26283 & ~n35121;
  assign n26297 = ~n26281 & ~n26296;
  assign n26298 = ~n6507 & ~n26297;
  assign n26299 = n6507 & ~n26281;
  assign n26300 = ~n26296 & n26299;
  assign n26301 = n6507 & n26297;
  assign n26302 = ~n25512 & ~n25515;
  assign n26303 = ~n25515 & ~n25830;
  assign n26304 = ~n25512 & n26303;
  assign n26305 = ~n25830 & n26302;
  assign n26306 = n25122 & ~n35123;
  assign n26307 = n25513 & n26303;
  assign n26308 = n25122 & ~n25515;
  assign n26309 = ~n25512 & n26308;
  assign n26310 = ~n25830 & n26309;
  assign n26311 = ~n25122 & ~n35123;
  assign n26312 = ~n26310 & ~n26311;
  assign n26313 = ~n26306 & ~n26307;
  assign n26314 = ~n35122 & ~n35124;
  assign n26315 = ~n26298 & ~n26314;
  assign n26316 = ~n6051 & ~n26315;
  assign n26317 = n6051 & ~n26298;
  assign n26318 = ~n26314 & n26317;
  assign n26319 = ~n35022 & ~n25521;
  assign n26320 = ~n25521 & ~n25830;
  assign n26321 = ~n35022 & n26320;
  assign n26322 = ~n25830 & n26319;
  assign n26323 = n25114 & ~n35125;
  assign n26324 = n25520 & n26320;
  assign n26325 = n25114 & ~n35022;
  assign n26326 = ~n25521 & n26325;
  assign n26327 = ~n25830 & n26326;
  assign n26328 = ~n25114 & ~n35125;
  assign n26329 = ~n26327 & ~n26328;
  assign n26330 = ~n26323 & ~n26324;
  assign n26331 = ~n26318 & ~n35126;
  assign n26332 = ~n26316 & ~n26331;
  assign n26333 = ~n5648 & ~n26332;
  assign n26334 = ~n25523 & ~n25538;
  assign n26335 = ~n25830 & n26334;
  assign n26336 = ~n35024 & ~n26335;
  assign n26337 = n35024 & ~n25538;
  assign n26338 = ~n25523 & n26337;
  assign n26339 = n35024 & n26335;
  assign n26340 = ~n25830 & n26338;
  assign n26341 = ~n26336 & ~n35127;
  assign n26342 = n5648 & ~n26316;
  assign n26343 = ~n26331 & n26342;
  assign n26344 = n5648 & n26332;
  assign n26345 = ~n26341 & ~n35128;
  assign n26346 = ~n26333 & ~n26345;
  assign n26347 = ~n5223 & ~n26346;
  assign n26348 = n5223 & ~n26333;
  assign n26349 = ~n26345 & n26348;
  assign n26350 = ~n35025 & ~n25544;
  assign n26351 = ~n25544 & ~n25830;
  assign n26352 = ~n35025 & n26351;
  assign n26353 = ~n25830 & n26350;
  assign n26354 = n25106 & ~n35129;
  assign n26355 = n25543 & n26351;
  assign n26356 = n25106 & ~n35025;
  assign n26357 = ~n25544 & n26356;
  assign n26358 = ~n25830 & n26357;
  assign n26359 = ~n25106 & ~n35129;
  assign n26360 = ~n26358 & ~n26359;
  assign n26361 = ~n26354 & ~n26355;
  assign n26362 = ~n26349 & ~n35130;
  assign n26363 = ~n26347 & ~n26362;
  assign n26364 = ~n4851 & ~n26363;
  assign n26365 = n4851 & ~n26347;
  assign n26366 = ~n26362 & n26365;
  assign n26367 = n4851 & n26363;
  assign n26368 = ~n25546 & ~n25549;
  assign n26369 = ~n25549 & ~n25830;
  assign n26370 = ~n25546 & n26369;
  assign n26371 = ~n25830 & n26368;
  assign n26372 = n25098 & ~n35132;
  assign n26373 = n25547 & n26369;
  assign n26374 = n25098 & ~n25549;
  assign n26375 = ~n25546 & n26374;
  assign n26376 = ~n25830 & n26375;
  assign n26377 = ~n25098 & ~n35132;
  assign n26378 = ~n26376 & ~n26377;
  assign n26379 = ~n26372 & ~n26373;
  assign n26380 = ~n35131 & ~n35133;
  assign n26381 = ~n26364 & ~n26380;
  assign n26382 = ~n4461 & ~n26381;
  assign n26383 = n4461 & ~n26364;
  assign n26384 = ~n26380 & n26383;
  assign n26385 = ~n35026 & ~n25555;
  assign n26386 = ~n25555 & ~n25830;
  assign n26387 = ~n35026 & n26386;
  assign n26388 = ~n25830 & n26385;
  assign n26389 = n25090 & ~n35134;
  assign n26390 = n25554 & n26386;
  assign n26391 = n25090 & ~n35026;
  assign n26392 = ~n25555 & n26391;
  assign n26393 = ~n25830 & n26392;
  assign n26394 = ~n25090 & ~n35134;
  assign n26395 = ~n26393 & ~n26394;
  assign n26396 = ~n26389 & ~n26390;
  assign n26397 = ~n26384 & ~n35135;
  assign n26398 = ~n26382 & ~n26397;
  assign n26399 = ~n4115 & ~n26398;
  assign n26400 = ~n25557 & ~n25572;
  assign n26401 = ~n25830 & n26400;
  assign n26402 = ~n35028 & ~n26401;
  assign n26403 = n35028 & ~n25572;
  assign n26404 = ~n25557 & n26403;
  assign n26405 = n35028 & n26401;
  assign n26406 = ~n25830 & n26404;
  assign n26407 = ~n26402 & ~n35136;
  assign n26408 = n4115 & ~n26382;
  assign n26409 = ~n26397 & n26408;
  assign n26410 = n4115 & n26398;
  assign n26411 = ~n26407 & ~n35137;
  assign n26412 = ~n26399 & ~n26411;
  assign n26413 = ~n3754 & ~n26412;
  assign n26414 = n3754 & ~n26399;
  assign n26415 = ~n26411 & n26414;
  assign n26416 = ~n35029 & ~n25578;
  assign n26417 = ~n25578 & ~n25830;
  assign n26418 = ~n35029 & n26417;
  assign n26419 = ~n25830 & n26416;
  assign n26420 = n25082 & ~n35138;
  assign n26421 = n25577 & n26417;
  assign n26422 = n25082 & ~n35029;
  assign n26423 = ~n25578 & n26422;
  assign n26424 = ~n25830 & n26423;
  assign n26425 = ~n25082 & ~n35138;
  assign n26426 = ~n26424 & ~n26425;
  assign n26427 = ~n26420 & ~n26421;
  assign n26428 = ~n26415 & ~n35139;
  assign n26429 = ~n26413 & ~n26428;
  assign n26430 = ~n3444 & ~n26429;
  assign n26431 = n3444 & ~n26413;
  assign n26432 = ~n26428 & n26431;
  assign n26433 = n3444 & n26429;
  assign n26434 = ~n25580 & ~n25583;
  assign n26435 = ~n25583 & ~n25830;
  assign n26436 = ~n25580 & n26435;
  assign n26437 = ~n25830 & n26434;
  assign n26438 = n25074 & ~n35141;
  assign n26439 = n25581 & n26435;
  assign n26440 = n25074 & ~n25583;
  assign n26441 = ~n25580 & n26440;
  assign n26442 = ~n25830 & n26441;
  assign n26443 = ~n25074 & ~n35141;
  assign n26444 = ~n26442 & ~n26443;
  assign n26445 = ~n26438 & ~n26439;
  assign n26446 = ~n35140 & ~n35142;
  assign n26447 = ~n26430 & ~n26446;
  assign n26448 = ~n3116 & ~n26447;
  assign n26449 = n3116 & ~n26430;
  assign n26450 = ~n26446 & n26449;
  assign n26451 = ~n35030 & ~n25589;
  assign n26452 = ~n25589 & ~n25830;
  assign n26453 = ~n35030 & n26452;
  assign n26454 = ~n25830 & n26451;
  assign n26455 = n25066 & ~n35143;
  assign n26456 = n25588 & n26452;
  assign n26457 = n25066 & ~n35030;
  assign n26458 = ~n25589 & n26457;
  assign n26459 = ~n25830 & n26458;
  assign n26460 = ~n25066 & ~n35143;
  assign n26461 = ~n26459 & ~n26460;
  assign n26462 = ~n26455 & ~n26456;
  assign n26463 = ~n26450 & ~n35144;
  assign n26464 = ~n26448 & ~n26463;
  assign n26465 = ~n2833 & ~n26464;
  assign n26466 = ~n25591 & ~n25606;
  assign n26467 = ~n25830 & n26466;
  assign n26468 = ~n35032 & ~n26467;
  assign n26469 = n35032 & ~n25606;
  assign n26470 = ~n25591 & n26469;
  assign n26471 = n35032 & n26467;
  assign n26472 = ~n25830 & n26470;
  assign n26473 = ~n26468 & ~n35145;
  assign n26474 = n2833 & ~n26448;
  assign n26475 = ~n26463 & n26474;
  assign n26476 = n2833 & n26464;
  assign n26477 = ~n26473 & ~n35146;
  assign n26478 = ~n26465 & ~n26477;
  assign n26479 = ~n2536 & ~n26478;
  assign n26480 = n2536 & ~n26465;
  assign n26481 = ~n26477 & n26480;
  assign n26482 = ~n35033 & ~n25612;
  assign n26483 = ~n25612 & ~n25830;
  assign n26484 = ~n35033 & n26483;
  assign n26485 = ~n25830 & n26482;
  assign n26486 = n25058 & ~n35147;
  assign n26487 = n25611 & n26483;
  assign n26488 = n25058 & ~n35033;
  assign n26489 = ~n25612 & n26488;
  assign n26490 = ~n25830 & n26489;
  assign n26491 = ~n25058 & ~n35147;
  assign n26492 = ~n26490 & ~n26491;
  assign n26493 = ~n26486 & ~n26487;
  assign n26494 = ~n26481 & ~n35148;
  assign n26495 = ~n26479 & ~n26494;
  assign n26496 = ~n2283 & ~n26495;
  assign n26497 = n2283 & ~n26479;
  assign n26498 = ~n26494 & n26497;
  assign n26499 = n2283 & n26495;
  assign n26500 = ~n25614 & ~n25617;
  assign n26501 = ~n25617 & ~n25830;
  assign n26502 = ~n25614 & n26501;
  assign n26503 = ~n25830 & n26500;
  assign n26504 = n25050 & ~n35150;
  assign n26505 = n25615 & n26501;
  assign n26506 = n25050 & ~n25617;
  assign n26507 = ~n25614 & n26506;
  assign n26508 = ~n25830 & n26507;
  assign n26509 = ~n25050 & ~n35150;
  assign n26510 = ~n26508 & ~n26509;
  assign n26511 = ~n26504 & ~n26505;
  assign n26512 = ~n35149 & ~n35151;
  assign n26513 = ~n26496 & ~n26512;
  assign n26514 = ~n2021 & ~n26513;
  assign n26515 = n2021 & ~n26496;
  assign n26516 = ~n26512 & n26515;
  assign n26517 = ~n35034 & ~n25623;
  assign n26518 = ~n25623 & ~n25830;
  assign n26519 = ~n35034 & n26518;
  assign n26520 = ~n25830 & n26517;
  assign n26521 = n25042 & ~n35152;
  assign n26522 = n25622 & n26518;
  assign n26523 = n25042 & ~n35034;
  assign n26524 = ~n25623 & n26523;
  assign n26525 = ~n25830 & n26524;
  assign n26526 = ~n25042 & ~n35152;
  assign n26527 = ~n26525 & ~n26526;
  assign n26528 = ~n26521 & ~n26522;
  assign n26529 = ~n26516 & ~n35153;
  assign n26530 = ~n26514 & ~n26529;
  assign n26531 = ~n1796 & ~n26530;
  assign n26532 = ~n25625 & ~n25640;
  assign n26533 = ~n25830 & n26532;
  assign n26534 = ~n35036 & ~n26533;
  assign n26535 = n35036 & ~n25640;
  assign n26536 = ~n25625 & n26535;
  assign n26537 = n35036 & n26533;
  assign n26538 = ~n25830 & n26536;
  assign n26539 = ~n26534 & ~n35154;
  assign n26540 = n1796 & ~n26514;
  assign n26541 = ~n26529 & n26540;
  assign n26542 = n1796 & n26530;
  assign n26543 = ~n26539 & ~n35155;
  assign n26544 = ~n26531 & ~n26543;
  assign n26545 = ~n1567 & ~n26544;
  assign n26546 = n1567 & ~n26531;
  assign n26547 = ~n26543 & n26546;
  assign n26548 = ~n35037 & ~n25646;
  assign n26549 = ~n25646 & ~n25830;
  assign n26550 = ~n35037 & n26549;
  assign n26551 = ~n25830 & n26548;
  assign n26552 = n25034 & ~n35156;
  assign n26553 = n25645 & n26549;
  assign n26554 = n25034 & ~n35037;
  assign n26555 = ~n25646 & n26554;
  assign n26556 = ~n25830 & n26555;
  assign n26557 = ~n25034 & ~n35156;
  assign n26558 = ~n26556 & ~n26557;
  assign n26559 = ~n26552 & ~n26553;
  assign n26560 = ~n26547 & ~n35157;
  assign n26561 = ~n26545 & ~n26560;
  assign n26562 = ~n1374 & ~n26561;
  assign n26563 = n1374 & ~n26545;
  assign n26564 = ~n26560 & n26563;
  assign n26565 = n1374 & n26561;
  assign n26566 = ~n25648 & ~n25651;
  assign n26567 = ~n25651 & ~n25830;
  assign n26568 = ~n25648 & n26567;
  assign n26569 = ~n25830 & n26566;
  assign n26570 = n25026 & ~n35159;
  assign n26571 = n25649 & n26567;
  assign n26572 = n25026 & ~n25651;
  assign n26573 = ~n25648 & n26572;
  assign n26574 = ~n25830 & n26573;
  assign n26575 = ~n25026 & ~n35159;
  assign n26576 = ~n26574 & ~n26575;
  assign n26577 = ~n26570 & ~n26571;
  assign n26578 = ~n35158 & ~n35160;
  assign n26579 = ~n26562 & ~n26578;
  assign n26580 = ~n1179 & ~n26579;
  assign n26581 = n1179 & ~n26562;
  assign n26582 = ~n26578 & n26581;
  assign n26583 = ~n35038 & ~n25657;
  assign n26584 = ~n25657 & ~n25830;
  assign n26585 = ~n35038 & n26584;
  assign n26586 = ~n25830 & n26583;
  assign n26587 = n25018 & ~n35161;
  assign n26588 = n25656 & n26584;
  assign n26589 = n25018 & ~n35038;
  assign n26590 = ~n25657 & n26589;
  assign n26591 = ~n25830 & n26590;
  assign n26592 = ~n25018 & ~n35161;
  assign n26593 = ~n26591 & ~n26592;
  assign n26594 = ~n26587 & ~n26588;
  assign n26595 = ~n26582 & ~n35162;
  assign n26596 = ~n26580 & ~n26595;
  assign n26597 = ~n1016 & ~n26596;
  assign n26598 = ~n25659 & ~n25674;
  assign n26599 = ~n25830 & n26598;
  assign n26600 = ~n35040 & ~n26599;
  assign n26601 = n35040 & ~n25674;
  assign n26602 = ~n25659 & n26601;
  assign n26603 = n35040 & n26599;
  assign n26604 = ~n25830 & n26602;
  assign n26605 = ~n26600 & ~n35163;
  assign n26606 = n1016 & ~n26580;
  assign n26607 = ~n26595 & n26606;
  assign n26608 = n1016 & n26596;
  assign n26609 = ~n26605 & ~n35164;
  assign n26610 = ~n26597 & ~n26609;
  assign n26611 = ~n855 & ~n26610;
  assign n26612 = n855 & ~n26597;
  assign n26613 = ~n26609 & n26612;
  assign n26614 = ~n35041 & ~n25680;
  assign n26615 = ~n25680 & ~n25830;
  assign n26616 = ~n35041 & n26615;
  assign n26617 = ~n25830 & n26614;
  assign n26618 = n25010 & ~n35165;
  assign n26619 = n25679 & n26615;
  assign n26620 = n25010 & ~n35041;
  assign n26621 = ~n25680 & n26620;
  assign n26622 = ~n25830 & n26621;
  assign n26623 = ~n25010 & ~n35165;
  assign n26624 = ~n26622 & ~n26623;
  assign n26625 = ~n26618 & ~n26619;
  assign n26626 = ~n26613 & ~n35166;
  assign n26627 = ~n26611 & ~n26626;
  assign n26628 = ~n720 & ~n26627;
  assign n26629 = n720 & ~n26611;
  assign n26630 = ~n26626 & n26629;
  assign n26631 = n720 & n26627;
  assign n26632 = ~n25682 & ~n25685;
  assign n26633 = ~n25685 & ~n25830;
  assign n26634 = ~n25682 & n26633;
  assign n26635 = ~n25830 & n26632;
  assign n26636 = n25002 & ~n35168;
  assign n26637 = n25683 & n26633;
  assign n26638 = n25002 & ~n25685;
  assign n26639 = ~n25682 & n26638;
  assign n26640 = ~n25830 & n26639;
  assign n26641 = ~n25002 & ~n35168;
  assign n26642 = ~n26640 & ~n26641;
  assign n26643 = ~n26636 & ~n26637;
  assign n26644 = ~n35167 & ~n35169;
  assign n26645 = ~n26628 & ~n26644;
  assign n26646 = ~n592 & ~n26645;
  assign n26647 = n592 & ~n26628;
  assign n26648 = ~n26644 & n26647;
  assign n26649 = ~n35042 & ~n25701;
  assign n26650 = ~n25830 & n26649;
  assign n26651 = ~n35043 & n26650;
  assign n26652 = n35043 & ~n26650;
  assign n26653 = ~n35042 & n35043;
  assign n26654 = ~n25701 & n26653;
  assign n26655 = ~n25830 & n26654;
  assign n26656 = ~n35043 & ~n26650;
  assign n26657 = ~n26655 & ~n26656;
  assign n26658 = ~n26651 & ~n26652;
  assign n26659 = ~n26648 & ~n35170;
  assign n26660 = ~n26646 & ~n26659;
  assign n26661 = ~n487 & ~n26660;
  assign n26662 = ~n25703 & ~n25715;
  assign n26663 = ~n25830 & n26662;
  assign n26664 = ~n35044 & ~n26663;
  assign n26665 = ~n25703 & n35044;
  assign n26666 = ~n25715 & n26665;
  assign n26667 = n35044 & n26663;
  assign n26668 = ~n25830 & n26666;
  assign n26669 = ~n26664 & ~n35171;
  assign n26670 = n487 & ~n26646;
  assign n26671 = ~n26659 & n26670;
  assign n26672 = n487 & n26660;
  assign n26673 = ~n26669 & ~n35172;
  assign n26674 = ~n26661 & ~n26673;
  assign n26675 = ~n393 & ~n26674;
  assign n26676 = n393 & ~n26661;
  assign n26677 = ~n26673 & n26676;
  assign n26678 = ~n25718 & ~n35046;
  assign n26679 = ~n25718 & ~n25830;
  assign n26680 = ~n35046 & n26679;
  assign n26681 = ~n25830 & n26678;
  assign n26682 = n25726 & ~n35173;
  assign n26683 = n25730 & n26679;
  assign n26684 = n25726 & ~n35046;
  assign n26685 = ~n25718 & n26684;
  assign n26686 = ~n25830 & n26685;
  assign n26687 = ~n25726 & ~n35173;
  assign n26688 = ~n26686 & ~n26687;
  assign n26689 = ~n26682 & ~n26683;
  assign n26690 = ~n26677 & ~n35174;
  assign n26691 = ~n26675 & ~n26690;
  assign n26692 = ~n321 & ~n26691;
  assign n26693 = ~n25732 & ~n25734;
  assign n26694 = ~n25830 & n26693;
  assign n26695 = ~n35048 & ~n26694;
  assign n26696 = ~n25732 & n35048;
  assign n26697 = ~n25734 & n26696;
  assign n26698 = n35048 & n26694;
  assign n26699 = ~n25830 & n26697;
  assign n26700 = ~n26695 & ~n35175;
  assign n26701 = n321 & ~n26675;
  assign n26702 = ~n26690 & n26701;
  assign n26703 = n321 & n26691;
  assign n26704 = ~n26700 & ~n35176;
  assign n26705 = ~n26692 & ~n26704;
  assign n26706 = ~n263 & ~n26705;
  assign n26707 = n263 & ~n26692;
  assign n26708 = ~n26704 & n26707;
  assign n26709 = ~n25749 & ~n35050;
  assign n26710 = ~n25749 & ~n25830;
  assign n26711 = ~n35050 & n26710;
  assign n26712 = ~n25830 & n26709;
  assign n26713 = n25757 & ~n35177;
  assign n26714 = n25761 & n26710;
  assign n26715 = n25757 & ~n35050;
  assign n26716 = ~n25749 & n26715;
  assign n26717 = ~n25830 & n26716;
  assign n26718 = ~n25757 & ~n35177;
  assign n26719 = ~n26717 & ~n26718;
  assign n26720 = ~n26713 & ~n26714;
  assign n26721 = ~n26708 & ~n35178;
  assign n26722 = ~n26706 & ~n26721;
  assign n26723 = ~n214 & ~n26722;
  assign n26724 = ~n25763 & ~n25765;
  assign n26725 = ~n25830 & n26724;
  assign n26726 = ~n35052 & ~n26725;
  assign n26727 = ~n25763 & n35052;
  assign n26728 = ~n25765 & n26727;
  assign n26729 = n35052 & n26725;
  assign n26730 = ~n25830 & n26728;
  assign n26731 = ~n26726 & ~n35179;
  assign n26732 = n214 & ~n26706;
  assign n26733 = ~n26721 & n26732;
  assign n26734 = n214 & n26722;
  assign n26735 = ~n26731 & ~n35180;
  assign n26736 = ~n26723 & ~n26735;
  assign n26737 = ~n197 & ~n26736;
  assign n26738 = n197 & ~n26723;
  assign n26739 = ~n26735 & n26738;
  assign n26740 = ~n25780 & ~n35054;
  assign n26741 = ~n25780 & ~n25830;
  assign n26742 = ~n35054 & n26741;
  assign n26743 = ~n25830 & n26740;
  assign n26744 = n25788 & ~n35181;
  assign n26745 = n25792 & n26741;
  assign n26746 = n25788 & ~n35054;
  assign n26747 = ~n25780 & n26746;
  assign n26748 = ~n25830 & n26747;
  assign n26749 = ~n25788 & ~n35181;
  assign n26750 = ~n26748 & ~n26749;
  assign n26751 = ~n26744 & ~n26745;
  assign n26752 = ~n26739 & ~n35182;
  assign n26753 = ~n26737 & ~n26752;
  assign n26754 = ~n25794 & ~n25804;
  assign n26755 = ~n25794 & ~n25830;
  assign n26756 = ~n25804 & n26755;
  assign n26757 = ~n25830 & n26754;
  assign n26758 = n25802 & ~n35183;
  assign n26759 = n25805 & n26755;
  assign n26760 = ~n25794 & n25802;
  assign n26761 = ~n25804 & n26760;
  assign n26762 = ~n25830 & n26761;
  assign n26763 = ~n25802 & ~n35183;
  assign n26764 = ~n26762 & ~n26763;
  assign n26765 = ~n26758 & ~n26759;
  assign n26766 = ~n25806 & ~n25814;
  assign n26767 = ~n25814 & ~n25830;
  assign n26768 = ~n25806 & n26767;
  assign n26769 = ~n25830 & n26766;
  assign n26770 = ~n35058 & ~n35185;
  assign n26771 = ~n35184 & n26770;
  assign n26772 = ~n26753 & n26771;
  assign n26773 = n193 & ~n26772;
  assign n26774 = ~n26737 & n35184;
  assign n26775 = ~n26752 & n26774;
  assign n26776 = n26753 & n35184;
  assign n26777 = n25806 & ~n26767;
  assign n26778 = ~n193 & ~n26766;
  assign n26779 = ~n26777 & n26778;
  assign n26780 = ~n35186 & ~n26779;
  assign n26781 = ~n26773 & n26780;
  assign n26782 = ~n26661 & n26669;
  assign n26783 = ~n35172 & n26782;
  assign n26784 = ~n26661 & ~n35172;
  assign n26785 = ~n26781 & n26784;
  assign n26786 = n26669 & n26785;
  assign n26787 = ~n26781 & n26783;
  assign n26788 = ~n26669 & ~n26785;
  assign n26789 = ~n35187 & ~n26788;
  assign n26790 = ~n26646 & ~n26648;
  assign n26791 = ~n26781 & n26790;
  assign n26792 = ~n35170 & ~n26791;
  assign n26793 = ~n26648 & n35170;
  assign n26794 = ~n26646 & n26793;
  assign n26795 = n35170 & n26791;
  assign n26796 = ~n26781 & n26794;
  assign n26797 = ~n26792 & ~n35188;
  assign n26798 = ~n26628 & ~n35167;
  assign n26799 = ~n26781 & n26798;
  assign n26800 = ~n35169 & ~n26799;
  assign n26801 = ~n26628 & n35169;
  assign n26802 = ~n35167 & n26801;
  assign n26803 = n35169 & n26799;
  assign n26804 = ~n26781 & n26802;
  assign n26805 = ~n26800 & ~n35189;
  assign n26806 = ~n26611 & ~n26613;
  assign n26807 = ~n26781 & n26806;
  assign n26808 = ~n35166 & ~n26807;
  assign n26809 = ~n26613 & n35166;
  assign n26810 = ~n26611 & n26809;
  assign n26811 = n35166 & n26807;
  assign n26812 = ~n26781 & n26810;
  assign n26813 = ~n26808 & ~n35190;
  assign n26814 = ~n26580 & ~n26582;
  assign n26815 = ~n26781 & n26814;
  assign n26816 = ~n35162 & ~n26815;
  assign n26817 = ~n26582 & n35162;
  assign n26818 = ~n26580 & n26817;
  assign n26819 = n35162 & n26815;
  assign n26820 = ~n26781 & n26818;
  assign n26821 = ~n26816 & ~n35191;
  assign n26822 = ~n26562 & ~n35158;
  assign n26823 = ~n26781 & n26822;
  assign n26824 = ~n35160 & ~n26823;
  assign n26825 = ~n26562 & n35160;
  assign n26826 = ~n35158 & n26825;
  assign n26827 = n35160 & n26823;
  assign n26828 = ~n26781 & n26826;
  assign n26829 = ~n26824 & ~n35192;
  assign n26830 = ~n26545 & ~n26547;
  assign n26831 = ~n26781 & n26830;
  assign n26832 = ~n35157 & ~n26831;
  assign n26833 = ~n26547 & n35157;
  assign n26834 = ~n26545 & n26833;
  assign n26835 = n35157 & n26831;
  assign n26836 = ~n26781 & n26834;
  assign n26837 = ~n26832 & ~n35193;
  assign n26838 = ~n26514 & ~n26516;
  assign n26839 = ~n26781 & n26838;
  assign n26840 = ~n35153 & ~n26839;
  assign n26841 = ~n26516 & n35153;
  assign n26842 = ~n26514 & n26841;
  assign n26843 = n35153 & n26839;
  assign n26844 = ~n26781 & n26842;
  assign n26845 = ~n26840 & ~n35194;
  assign n26846 = ~n26496 & ~n35149;
  assign n26847 = ~n26781 & n26846;
  assign n26848 = ~n35151 & ~n26847;
  assign n26849 = ~n26496 & n35151;
  assign n26850 = ~n35149 & n26849;
  assign n26851 = n35151 & n26847;
  assign n26852 = ~n26781 & n26850;
  assign n26853 = ~n26848 & ~n35195;
  assign n26854 = ~n26479 & ~n26481;
  assign n26855 = ~n26781 & n26854;
  assign n26856 = ~n35148 & ~n26855;
  assign n26857 = ~n26481 & n35148;
  assign n26858 = ~n26479 & n26857;
  assign n26859 = n35148 & n26855;
  assign n26860 = ~n26781 & n26858;
  assign n26861 = ~n26856 & ~n35196;
  assign n26862 = ~n26448 & ~n26450;
  assign n26863 = ~n26781 & n26862;
  assign n26864 = ~n35144 & ~n26863;
  assign n26865 = ~n26450 & n35144;
  assign n26866 = ~n26448 & n26865;
  assign n26867 = n35144 & n26863;
  assign n26868 = ~n26781 & n26866;
  assign n26869 = ~n26864 & ~n35197;
  assign n26870 = ~n26430 & ~n35140;
  assign n26871 = ~n26781 & n26870;
  assign n26872 = ~n35142 & ~n26871;
  assign n26873 = ~n26430 & n35142;
  assign n26874 = ~n35140 & n26873;
  assign n26875 = n35142 & n26871;
  assign n26876 = ~n26781 & n26874;
  assign n26877 = ~n26872 & ~n35198;
  assign n26878 = ~n26413 & ~n26415;
  assign n26879 = ~n26781 & n26878;
  assign n26880 = ~n35139 & ~n26879;
  assign n26881 = ~n26415 & n35139;
  assign n26882 = ~n26413 & n26881;
  assign n26883 = n35139 & n26879;
  assign n26884 = ~n26781 & n26882;
  assign n26885 = ~n26880 & ~n35199;
  assign n26886 = ~n26382 & ~n26384;
  assign n26887 = ~n26781 & n26886;
  assign n26888 = ~n35135 & ~n26887;
  assign n26889 = ~n26384 & n35135;
  assign n26890 = ~n26382 & n26889;
  assign n26891 = n35135 & n26887;
  assign n26892 = ~n26781 & n26890;
  assign n26893 = ~n26888 & ~n35200;
  assign n26894 = ~n26364 & ~n35131;
  assign n26895 = ~n26781 & n26894;
  assign n26896 = ~n35133 & ~n26895;
  assign n26897 = ~n26364 & n35133;
  assign n26898 = ~n35131 & n26897;
  assign n26899 = n35133 & n26895;
  assign n26900 = ~n26781 & n26898;
  assign n26901 = ~n26896 & ~n35201;
  assign n26902 = ~n26347 & ~n26349;
  assign n26903 = ~n26781 & n26902;
  assign n26904 = ~n35130 & ~n26903;
  assign n26905 = ~n26349 & n35130;
  assign n26906 = ~n26347 & n26905;
  assign n26907 = n35130 & n26903;
  assign n26908 = ~n26781 & n26906;
  assign n26909 = ~n26904 & ~n35202;
  assign n26910 = ~n26316 & ~n26318;
  assign n26911 = ~n26781 & n26910;
  assign n26912 = ~n35126 & ~n26911;
  assign n26913 = ~n26318 & n35126;
  assign n26914 = ~n26316 & n26913;
  assign n26915 = n35126 & n26911;
  assign n26916 = ~n26781 & n26914;
  assign n26917 = ~n26912 & ~n35203;
  assign n26918 = ~n26298 & ~n35122;
  assign n26919 = ~n26781 & n26918;
  assign n26920 = ~n35124 & ~n26919;
  assign n26921 = ~n26298 & n35124;
  assign n26922 = ~n35122 & n26921;
  assign n26923 = n35124 & n26919;
  assign n26924 = ~n26781 & n26922;
  assign n26925 = ~n26920 & ~n35204;
  assign n26926 = ~n26281 & ~n26283;
  assign n26927 = ~n26781 & n26926;
  assign n26928 = ~n35121 & ~n26927;
  assign n26929 = ~n26283 & n35121;
  assign n26930 = ~n26281 & n26929;
  assign n26931 = n35121 & n26927;
  assign n26932 = ~n26781 & n26930;
  assign n26933 = ~n26928 & ~n35205;
  assign n26934 = ~n26250 & ~n26252;
  assign n26935 = ~n26781 & n26934;
  assign n26936 = ~n35117 & ~n26935;
  assign n26937 = ~n26252 & n35117;
  assign n26938 = ~n26250 & n26937;
  assign n26939 = n35117 & n26935;
  assign n26940 = ~n26781 & n26938;
  assign n26941 = ~n26936 & ~n35206;
  assign n26942 = ~n26232 & ~n35113;
  assign n26943 = ~n26781 & n26942;
  assign n26944 = ~n35115 & ~n26943;
  assign n26945 = ~n26232 & n35115;
  assign n26946 = ~n35113 & n26945;
  assign n26947 = n35115 & n26943;
  assign n26948 = ~n26781 & n26946;
  assign n26949 = ~n26944 & ~n35207;
  assign n26950 = ~n26215 & ~n26217;
  assign n26951 = ~n26781 & n26950;
  assign n26952 = ~n35112 & ~n26951;
  assign n26953 = ~n26217 & n35112;
  assign n26954 = ~n26215 & n26953;
  assign n26955 = n35112 & n26951;
  assign n26956 = ~n26781 & n26954;
  assign n26957 = ~n26952 & ~n35208;
  assign n26958 = ~n26184 & ~n26186;
  assign n26959 = ~n26781 & n26958;
  assign n26960 = ~n35108 & ~n26959;
  assign n26961 = ~n26186 & n35108;
  assign n26962 = ~n26184 & n26961;
  assign n26963 = n35108 & n26959;
  assign n26964 = ~n26781 & n26962;
  assign n26965 = ~n26960 & ~n35209;
  assign n26966 = ~n26166 & ~n35104;
  assign n26967 = ~n26781 & n26966;
  assign n26968 = ~n35106 & ~n26967;
  assign n26969 = ~n26166 & n35106;
  assign n26970 = ~n35104 & n26969;
  assign n26971 = n35106 & n26967;
  assign n26972 = ~n26781 & n26970;
  assign n26973 = ~n26968 & ~n35210;
  assign n26974 = ~n26149 & ~n26151;
  assign n26975 = ~n26781 & n26974;
  assign n26976 = ~n35103 & ~n26975;
  assign n26977 = ~n26151 & n35103;
  assign n26978 = ~n26149 & n26977;
  assign n26979 = n35103 & n26975;
  assign n26980 = ~n26781 & n26978;
  assign n26981 = ~n26976 & ~n35211;
  assign n26982 = ~n26118 & ~n26120;
  assign n26983 = ~n26781 & n26982;
  assign n26984 = ~n35099 & ~n26983;
  assign n26985 = ~n26120 & n35099;
  assign n26986 = ~n26118 & n26985;
  assign n26987 = n35099 & n26983;
  assign n26988 = ~n26781 & n26986;
  assign n26989 = ~n26984 & ~n35212;
  assign n26990 = ~n26100 & ~n35095;
  assign n26991 = ~n26781 & n26990;
  assign n26992 = ~n35097 & ~n26991;
  assign n26993 = ~n26100 & n35097;
  assign n26994 = ~n35095 & n26993;
  assign n26995 = n35097 & n26991;
  assign n26996 = ~n26781 & n26994;
  assign n26997 = ~n26992 & ~n35213;
  assign n26998 = ~n26083 & ~n26085;
  assign n26999 = ~n26781 & n26998;
  assign n27000 = ~n35094 & ~n26999;
  assign n27001 = ~n26085 & n35094;
  assign n27002 = ~n26083 & n27001;
  assign n27003 = n35094 & n26999;
  assign n27004 = ~n26781 & n27002;
  assign n27005 = ~n27000 & ~n35214;
  assign n27006 = ~n26052 & ~n26054;
  assign n27007 = ~n26781 & n27006;
  assign n27008 = ~n35090 & ~n27007;
  assign n27009 = ~n26054 & n35090;
  assign n27010 = ~n26052 & n27009;
  assign n27011 = n35090 & n27007;
  assign n27012 = ~n26781 & n27010;
  assign n27013 = ~n27008 & ~n35215;
  assign n27014 = ~n26033 & ~n35085;
  assign n27015 = ~n26781 & n27014;
  assign n27016 = ~n35088 & ~n27015;
  assign n27017 = ~n26033 & n35088;
  assign n27018 = ~n35085 & n27017;
  assign n27019 = n35088 & n27015;
  assign n27020 = ~n26781 & n27018;
  assign n27021 = ~n27016 & ~n35216;
  assign n27022 = ~n26016 & ~n26018;
  assign n27023 = ~n26781 & n27022;
  assign n27024 = ~n35084 & ~n27023;
  assign n27025 = ~n26018 & n35084;
  assign n27026 = ~n26016 & n27025;
  assign n27027 = n35084 & n27023;
  assign n27028 = ~n26781 & n27026;
  assign n27029 = ~n27024 & ~n35217;
  assign n27030 = ~n25982 & ~n25984;
  assign n27031 = ~n26781 & n27030;
  assign n27032 = ~n35079 & ~n27031;
  assign n27033 = ~n25984 & n35079;
  assign n27034 = ~n25982 & n27033;
  assign n27035 = n35079 & n27031;
  assign n27036 = ~n26781 & n27034;
  assign n27037 = ~n27032 & ~n35218;
  assign n27038 = ~n25949 & ~n25951;
  assign n27039 = ~n26781 & n27038;
  assign n27040 = ~n35075 & ~n27039;
  assign n27041 = ~n25951 & n35075;
  assign n27042 = ~n25949 & n27041;
  assign n27043 = n35075 & n27039;
  assign n27044 = ~n26781 & n27042;
  assign n27045 = ~n27040 & ~n35219;
  assign n27046 = ~n25916 & ~n25918;
  assign n27047 = ~n26781 & n27046;
  assign n27048 = ~n35071 & ~n27047;
  assign n27049 = ~n25918 & n35071;
  assign n27050 = ~n25916 & n27049;
  assign n27051 = n35071 & n27047;
  assign n27052 = ~n26781 & n27050;
  assign n27053 = ~n27048 & ~n35220;
  assign n27054 = ~n25882 & ~n25884;
  assign n27055 = ~n26781 & n27054;
  assign n27056 = ~n35066 & ~n27055;
  assign n27057 = ~n25884 & n35066;
  assign n27058 = ~n25882 & n27057;
  assign n27059 = n35066 & n27055;
  assign n27060 = ~n26781 & n27058;
  assign n27061 = ~n27056 & ~n35221;
  assign n27062 = ~n25855 & ~n25857;
  assign n27063 = ~n26781 & n27062;
  assign n27064 = ~n25866 & ~n27063;
  assign n27065 = ~n25857 & n25866;
  assign n27066 = ~n25855 & n27065;
  assign n27067 = n25866 & n27063;
  assign n27068 = ~n26781 & n27066;
  assign n27069 = ~n27064 & ~n35222;
  assign n27070 = ~pi10  & ~n26781;
  assign n27071 = ~pi11  & n27070;
  assign n27072 = n25832 & ~n26781;
  assign n27073 = ~n25830 & ~n26779;
  assign n27074 = ~n35186 & n27073;
  assign n27075 = ~n25830 & n26781;
  assign n27076 = ~n26773 & n27074;
  assign n27077 = ~n35223 & ~n35224;
  assign n27078 = pi12  & ~n27077;
  assign n27079 = ~pi12  & ~n35224;
  assign n27080 = ~pi12  & n27077;
  assign n27081 = ~n35223 & n27079;
  assign n27082 = ~n27078 & ~n35225;
  assign n27083 = pi10  & ~n26781;
  assign n27084 = ~pi8  & ~pi9 ;
  assign n27085 = ~pi10  & n27084;
  assign n27086 = ~n34955 & ~n35060;
  assign n27087 = ~n24973 & n27086;
  assign n27088 = ~n24992 & n27087;
  assign n27089 = ~n34957 & n27088;
  assign n27090 = n24978 & n24994;
  assign n27091 = ~n24986 & n27089;
  assign n27092 = ~n27085 & ~n35226;
  assign n27093 = ~n25828 & n27092;
  assign n27094 = ~n35058 & n27093;
  assign n27095 = ~n25822 & n27094;
  assign n27096 = ~pi10  & ~n27084;
  assign n27097 = pi10  & n26781;
  assign n27098 = ~n27096 & ~n27097;
  assign n27099 = ~n27083 & ~n27085;
  assign n27100 = n25830 & ~n35227;
  assign n27101 = ~n27083 & n27095;
  assign n27102 = pi11  & ~n27070;
  assign n27103 = ~n35223 & ~n27102;
  assign n27104 = ~n35228 & n27103;
  assign n27105 = ~n25830 & n35227;
  assign n27106 = n24994 & ~n27105;
  assign n27107 = ~n27104 & ~n27105;
  assign n27108 = n24994 & n27107;
  assign n27109 = ~n27104 & n27106;
  assign n27110 = ~n27082 & ~n35229;
  assign n27111 = ~n24994 & ~n27107;
  assign n27112 = n24076 & ~n27111;
  assign n27113 = ~n27110 & n27112;
  assign n27114 = ~n25835 & ~n35061;
  assign n27115 = ~n26781 & n27114;
  assign n27116 = n25840 & ~n27115;
  assign n27117 = ~n25840 & n27114;
  assign n27118 = ~n25840 & n27115;
  assign n27119 = ~n26781 & n27117;
  assign n27120 = ~n27116 & ~n35230;
  assign n27121 = ~n27113 & ~n27120;
  assign n27122 = ~n27110 & ~n27111;
  assign n27123 = ~n24076 & ~n27122;
  assign n27124 = n23269 & ~n27123;
  assign n27125 = ~n27121 & ~n27123;
  assign n27126 = n23269 & n27125;
  assign n27127 = ~n27121 & n27124;
  assign n27128 = ~n27069 & ~n35231;
  assign n27129 = ~n23269 & ~n27125;
  assign n27130 = n22386 & ~n27129;
  assign n27131 = ~n27128 & n27130;
  assign n27132 = ~n25869 & ~n35063;
  assign n27133 = ~n26781 & n27132;
  assign n27134 = ~n25879 & ~n27133;
  assign n27135 = ~n25869 & n25879;
  assign n27136 = ~n35063 & n27135;
  assign n27137 = n25879 & n27133;
  assign n27138 = ~n26781 & n27136;
  assign n27139 = n25879 & ~n27133;
  assign n27140 = ~n25879 & n27133;
  assign n27141 = ~n27139 & ~n27140;
  assign n27142 = ~n27134 & ~n35232;
  assign n27143 = ~n27131 & n35233;
  assign n27144 = ~n27128 & ~n27129;
  assign n27145 = ~n22386 & ~n27144;
  assign n27146 = n21612 & ~n27145;
  assign n27147 = ~n27143 & ~n27145;
  assign n27148 = n21612 & n27147;
  assign n27149 = ~n27143 & n27146;
  assign n27150 = ~n27061 & ~n35234;
  assign n27151 = ~n21612 & ~n27147;
  assign n27152 = n20762 & ~n27151;
  assign n27153 = ~n27150 & n27152;
  assign n27154 = ~n25899 & ~n35067;
  assign n27155 = ~n26781 & n27154;
  assign n27156 = ~n35069 & ~n27155;
  assign n27157 = n35069 & n27155;
  assign n27158 = ~n25899 & ~n35069;
  assign n27159 = ~n35067 & n27158;
  assign n27160 = ~n26781 & n27159;
  assign n27161 = n35069 & ~n27155;
  assign n27162 = ~n27160 & ~n27161;
  assign n27163 = ~n27156 & ~n27157;
  assign n27164 = ~n27153 & ~n35235;
  assign n27165 = ~n27150 & ~n27151;
  assign n27166 = ~n20762 & ~n27165;
  assign n27167 = n20011 & ~n27166;
  assign n27168 = ~n27164 & ~n27166;
  assign n27169 = n20011 & n27168;
  assign n27170 = ~n27164 & n27167;
  assign n27171 = ~n27053 & ~n35236;
  assign n27172 = ~n20011 & ~n27168;
  assign n27173 = n19190 & ~n27172;
  assign n27174 = ~n27171 & n27173;
  assign n27175 = ~n25933 & ~n35072;
  assign n27176 = ~n26781 & n27175;
  assign n27177 = ~n35073 & n27176;
  assign n27178 = n35073 & ~n27176;
  assign n27179 = ~n25933 & n35073;
  assign n27180 = ~n35072 & n27179;
  assign n27181 = ~n26781 & n27180;
  assign n27182 = ~n35073 & ~n27176;
  assign n27183 = ~n27181 & ~n27182;
  assign n27184 = ~n27177 & ~n27178;
  assign n27185 = ~n27174 & ~n35237;
  assign n27186 = ~n27171 & ~n27172;
  assign n27187 = ~n19190 & ~n27186;
  assign n27188 = n18472 & ~n27187;
  assign n27189 = ~n27185 & ~n27187;
  assign n27190 = n18472 & n27189;
  assign n27191 = ~n27185 & n27188;
  assign n27192 = ~n27045 & ~n35238;
  assign n27193 = ~n18472 & ~n27189;
  assign n27194 = n17690 & ~n27193;
  assign n27195 = ~n27192 & n27194;
  assign n27196 = ~n25966 & ~n35076;
  assign n27197 = ~n26781 & n27196;
  assign n27198 = ~n35077 & n27197;
  assign n27199 = n35077 & ~n27197;
  assign n27200 = ~n35077 & ~n27197;
  assign n27201 = ~n25966 & n35077;
  assign n27202 = ~n35076 & n27201;
  assign n27203 = n35077 & n27197;
  assign n27204 = ~n26781 & n27202;
  assign n27205 = ~n27200 & ~n35239;
  assign n27206 = ~n27198 & ~n27199;
  assign n27207 = ~n27195 & ~n35240;
  assign n27208 = ~n27192 & ~n27193;
  assign n27209 = ~n17690 & ~n27208;
  assign n27210 = n17001 & ~n27209;
  assign n27211 = ~n27207 & ~n27209;
  assign n27212 = n17001 & n27211;
  assign n27213 = ~n27207 & n27210;
  assign n27214 = ~n27037 & ~n35241;
  assign n27215 = ~n17001 & ~n27211;
  assign n27216 = n16248 & ~n27215;
  assign n27217 = ~n27214 & n27216;
  assign n27218 = ~n25999 & ~n35080;
  assign n27219 = ~n25999 & ~n26781;
  assign n27220 = ~n35080 & n27219;
  assign n27221 = ~n26781 & n27218;
  assign n27222 = n35082 & ~n35242;
  assign n27223 = n26014 & n27219;
  assign n27224 = ~n35082 & n35242;
  assign n27225 = ~n25999 & n35082;
  assign n27226 = ~n35080 & n27225;
  assign n27227 = ~n26781 & n27226;
  assign n27228 = ~n35082 & ~n35242;
  assign n27229 = ~n27227 & ~n27228;
  assign n27230 = ~n27222 & ~n35243;
  assign n27231 = ~n27217 & ~n35244;
  assign n27232 = ~n27214 & ~n27215;
  assign n27233 = ~n16248 & ~n27232;
  assign n27234 = n15586 & ~n27233;
  assign n27235 = ~n27231 & ~n27233;
  assign n27236 = n15586 & n27235;
  assign n27237 = ~n27231 & n27234;
  assign n27238 = ~n27029 & ~n35245;
  assign n27239 = ~n15586 & ~n27235;
  assign n27240 = n14866 & ~n27239;
  assign n27241 = ~n27238 & n27240;
  assign n27242 = ~n27021 & ~n27241;
  assign n27243 = ~n27238 & ~n27239;
  assign n27244 = ~n14866 & ~n27243;
  assign n27245 = n14233 & ~n27244;
  assign n27246 = ~n27242 & ~n27244;
  assign n27247 = n14233 & n27246;
  assign n27248 = ~n27242 & n27245;
  assign n27249 = ~n27013 & ~n35246;
  assign n27250 = ~n14233 & ~n27246;
  assign n27251 = n13548 & ~n27250;
  assign n27252 = ~n27249 & n27251;
  assign n27253 = ~n26069 & ~n35092;
  assign n27254 = ~n26069 & ~n26781;
  assign n27255 = ~n35092 & n27254;
  assign n27256 = ~n26781 & n27253;
  assign n27257 = n26077 & ~n35247;
  assign n27258 = n26081 & n27254;
  assign n27259 = ~n26069 & n26077;
  assign n27260 = ~n35092 & n27259;
  assign n27261 = ~n26781 & n27260;
  assign n27262 = ~n26077 & ~n35247;
  assign n27263 = ~n27261 & ~n27262;
  assign n27264 = ~n27257 & ~n27258;
  assign n27265 = ~n27252 & ~n35248;
  assign n27266 = ~n27249 & ~n27250;
  assign n27267 = ~n13548 & ~n27266;
  assign n27268 = n12948 & ~n27267;
  assign n27269 = ~n27265 & ~n27267;
  assign n27270 = n12948 & n27269;
  assign n27271 = ~n27265 & n27268;
  assign n27272 = ~n27005 & ~n35249;
  assign n27273 = ~n12948 & ~n27269;
  assign n27274 = n12296 & ~n27273;
  assign n27275 = ~n27272 & n27274;
  assign n27276 = ~n26997 & ~n27275;
  assign n27277 = ~n27272 & ~n27273;
  assign n27278 = ~n12296 & ~n27277;
  assign n27279 = n11719 & ~n27278;
  assign n27280 = ~n27276 & ~n27278;
  assign n27281 = n11719 & n27280;
  assign n27282 = ~n27276 & n27279;
  assign n27283 = ~n26989 & ~n35250;
  assign n27284 = ~n11719 & ~n27280;
  assign n27285 = n11097 & ~n27284;
  assign n27286 = ~n27283 & n27285;
  assign n27287 = ~n26135 & ~n35101;
  assign n27288 = ~n26135 & ~n26781;
  assign n27289 = ~n35101 & n27288;
  assign n27290 = ~n26781 & n27287;
  assign n27291 = n26143 & ~n35251;
  assign n27292 = n26147 & n27288;
  assign n27293 = ~n26135 & n26143;
  assign n27294 = ~n35101 & n27293;
  assign n27295 = ~n26781 & n27294;
  assign n27296 = ~n26143 & ~n35251;
  assign n27297 = ~n27295 & ~n27296;
  assign n27298 = ~n27291 & ~n27292;
  assign n27299 = ~n27286 & ~n35252;
  assign n27300 = ~n27283 & ~n27284;
  assign n27301 = ~n11097 & ~n27300;
  assign n27302 = n10555 & ~n27301;
  assign n27303 = ~n27299 & ~n27301;
  assign n27304 = n10555 & n27303;
  assign n27305 = ~n27299 & n27302;
  assign n27306 = ~n26981 & ~n35253;
  assign n27307 = ~n10555 & ~n27303;
  assign n27308 = n9969 & ~n27307;
  assign n27309 = ~n27306 & n27308;
  assign n27310 = ~n26973 & ~n27309;
  assign n27311 = ~n27306 & ~n27307;
  assign n27312 = ~n9969 & ~n27311;
  assign n27313 = n9457 & ~n27312;
  assign n27314 = ~n27310 & ~n27312;
  assign n27315 = n9457 & n27314;
  assign n27316 = ~n27310 & n27313;
  assign n27317 = ~n26965 & ~n35254;
  assign n27318 = ~n9457 & ~n27314;
  assign n27319 = n8896 & ~n27318;
  assign n27320 = ~n27317 & n27319;
  assign n27321 = ~n26201 & ~n35110;
  assign n27322 = ~n26201 & ~n26781;
  assign n27323 = ~n35110 & n27322;
  assign n27324 = ~n26781 & n27321;
  assign n27325 = n26209 & ~n35255;
  assign n27326 = n26213 & n27322;
  assign n27327 = ~n26201 & n26209;
  assign n27328 = ~n35110 & n27327;
  assign n27329 = ~n26781 & n27328;
  assign n27330 = ~n26209 & ~n35255;
  assign n27331 = ~n27329 & ~n27330;
  assign n27332 = ~n27325 & ~n27326;
  assign n27333 = ~n27320 & ~n35256;
  assign n27334 = ~n27317 & ~n27318;
  assign n27335 = ~n8896 & ~n27334;
  assign n27336 = n8411 & ~n27335;
  assign n27337 = ~n27333 & ~n27335;
  assign n27338 = n8411 & n27337;
  assign n27339 = ~n27333 & n27336;
  assign n27340 = ~n26957 & ~n35257;
  assign n27341 = ~n8411 & ~n27337;
  assign n27342 = n7885 & ~n27341;
  assign n27343 = ~n27340 & n27342;
  assign n27344 = ~n26949 & ~n27343;
  assign n27345 = ~n27340 & ~n27341;
  assign n27346 = ~n7885 & ~n27345;
  assign n27347 = n7428 & ~n27346;
  assign n27348 = ~n27344 & ~n27346;
  assign n27349 = n7428 & n27348;
  assign n27350 = ~n27344 & n27347;
  assign n27351 = ~n26941 & ~n35258;
  assign n27352 = ~n7428 & ~n27348;
  assign n27353 = n6937 & ~n27352;
  assign n27354 = ~n27351 & n27353;
  assign n27355 = ~n26267 & ~n35119;
  assign n27356 = ~n26267 & ~n26781;
  assign n27357 = ~n35119 & n27356;
  assign n27358 = ~n26781 & n27355;
  assign n27359 = n26275 & ~n35259;
  assign n27360 = n26279 & n27356;
  assign n27361 = ~n26267 & n26275;
  assign n27362 = ~n35119 & n27361;
  assign n27363 = ~n26781 & n27362;
  assign n27364 = ~n26275 & ~n35259;
  assign n27365 = ~n27363 & ~n27364;
  assign n27366 = ~n27359 & ~n27360;
  assign n27367 = ~n27354 & ~n35260;
  assign n27368 = ~n27351 & ~n27352;
  assign n27369 = ~n6937 & ~n27368;
  assign n27370 = n6507 & ~n27369;
  assign n27371 = ~n27367 & ~n27369;
  assign n27372 = n6507 & n27371;
  assign n27373 = ~n27367 & n27370;
  assign n27374 = ~n26933 & ~n35261;
  assign n27375 = ~n6507 & ~n27371;
  assign n27376 = n6051 & ~n27375;
  assign n27377 = ~n27374 & n27376;
  assign n27378 = ~n26925 & ~n27377;
  assign n27379 = ~n27374 & ~n27375;
  assign n27380 = ~n6051 & ~n27379;
  assign n27381 = n5648 & ~n27380;
  assign n27382 = ~n27378 & ~n27380;
  assign n27383 = n5648 & n27382;
  assign n27384 = ~n27378 & n27381;
  assign n27385 = ~n26917 & ~n35262;
  assign n27386 = ~n5648 & ~n27382;
  assign n27387 = n5223 & ~n27386;
  assign n27388 = ~n27385 & n27387;
  assign n27389 = ~n26333 & ~n35128;
  assign n27390 = ~n26333 & ~n26781;
  assign n27391 = ~n35128 & n27390;
  assign n27392 = ~n26781 & n27389;
  assign n27393 = n26341 & ~n35263;
  assign n27394 = n26345 & n27390;
  assign n27395 = ~n26333 & n26341;
  assign n27396 = ~n35128 & n27395;
  assign n27397 = ~n26781 & n27396;
  assign n27398 = ~n26341 & ~n35263;
  assign n27399 = ~n27397 & ~n27398;
  assign n27400 = ~n27393 & ~n27394;
  assign n27401 = ~n27388 & ~n35264;
  assign n27402 = ~n27385 & ~n27386;
  assign n27403 = ~n5223 & ~n27402;
  assign n27404 = n4851 & ~n27403;
  assign n27405 = ~n27401 & ~n27403;
  assign n27406 = n4851 & n27405;
  assign n27407 = ~n27401 & n27404;
  assign n27408 = ~n26909 & ~n35265;
  assign n27409 = ~n4851 & ~n27405;
  assign n27410 = n4461 & ~n27409;
  assign n27411 = ~n27408 & n27410;
  assign n27412 = ~n26901 & ~n27411;
  assign n27413 = ~n27408 & ~n27409;
  assign n27414 = ~n4461 & ~n27413;
  assign n27415 = n4115 & ~n27414;
  assign n27416 = ~n27412 & ~n27414;
  assign n27417 = n4115 & n27416;
  assign n27418 = ~n27412 & n27415;
  assign n27419 = ~n26893 & ~n35266;
  assign n27420 = ~n4115 & ~n27416;
  assign n27421 = n3754 & ~n27420;
  assign n27422 = ~n27419 & n27421;
  assign n27423 = ~n26399 & ~n35137;
  assign n27424 = ~n26399 & ~n26781;
  assign n27425 = ~n35137 & n27424;
  assign n27426 = ~n26781 & n27423;
  assign n27427 = n26407 & ~n35267;
  assign n27428 = n26411 & n27424;
  assign n27429 = ~n26399 & n26407;
  assign n27430 = ~n35137 & n27429;
  assign n27431 = ~n26781 & n27430;
  assign n27432 = ~n26407 & ~n35267;
  assign n27433 = ~n27431 & ~n27432;
  assign n27434 = ~n27427 & ~n27428;
  assign n27435 = ~n27422 & ~n35268;
  assign n27436 = ~n27419 & ~n27420;
  assign n27437 = ~n3754 & ~n27436;
  assign n27438 = n3444 & ~n27437;
  assign n27439 = ~n27435 & ~n27437;
  assign n27440 = n3444 & n27439;
  assign n27441 = ~n27435 & n27438;
  assign n27442 = ~n26885 & ~n35269;
  assign n27443 = ~n3444 & ~n27439;
  assign n27444 = n3116 & ~n27443;
  assign n27445 = ~n27442 & n27444;
  assign n27446 = ~n26877 & ~n27445;
  assign n27447 = ~n27442 & ~n27443;
  assign n27448 = ~n3116 & ~n27447;
  assign n27449 = n2833 & ~n27448;
  assign n27450 = ~n27446 & ~n27448;
  assign n27451 = n2833 & n27450;
  assign n27452 = ~n27446 & n27449;
  assign n27453 = ~n26869 & ~n35270;
  assign n27454 = ~n2833 & ~n27450;
  assign n27455 = n2536 & ~n27454;
  assign n27456 = ~n27453 & n27455;
  assign n27457 = ~n26465 & ~n35146;
  assign n27458 = ~n26465 & ~n26781;
  assign n27459 = ~n35146 & n27458;
  assign n27460 = ~n26781 & n27457;
  assign n27461 = n26473 & ~n35271;
  assign n27462 = n26477 & n27458;
  assign n27463 = ~n26465 & n26473;
  assign n27464 = ~n35146 & n27463;
  assign n27465 = ~n26781 & n27464;
  assign n27466 = ~n26473 & ~n35271;
  assign n27467 = ~n27465 & ~n27466;
  assign n27468 = ~n27461 & ~n27462;
  assign n27469 = ~n27456 & ~n35272;
  assign n27470 = ~n27453 & ~n27454;
  assign n27471 = ~n2536 & ~n27470;
  assign n27472 = n2283 & ~n27471;
  assign n27473 = ~n27469 & ~n27471;
  assign n27474 = n2283 & n27473;
  assign n27475 = ~n27469 & n27472;
  assign n27476 = ~n26861 & ~n35273;
  assign n27477 = ~n2283 & ~n27473;
  assign n27478 = n2021 & ~n27477;
  assign n27479 = ~n27476 & n27478;
  assign n27480 = ~n26853 & ~n27479;
  assign n27481 = ~n27476 & ~n27477;
  assign n27482 = ~n2021 & ~n27481;
  assign n27483 = n1796 & ~n27482;
  assign n27484 = ~n27480 & ~n27482;
  assign n27485 = n1796 & n27484;
  assign n27486 = ~n27480 & n27483;
  assign n27487 = ~n26845 & ~n35274;
  assign n27488 = ~n1796 & ~n27484;
  assign n27489 = n1567 & ~n27488;
  assign n27490 = ~n27487 & n27489;
  assign n27491 = ~n26531 & ~n35155;
  assign n27492 = ~n26531 & ~n26781;
  assign n27493 = ~n35155 & n27492;
  assign n27494 = ~n26781 & n27491;
  assign n27495 = n26539 & ~n35275;
  assign n27496 = n26543 & n27492;
  assign n27497 = ~n26531 & n26539;
  assign n27498 = ~n35155 & n27497;
  assign n27499 = ~n26781 & n27498;
  assign n27500 = ~n26539 & ~n35275;
  assign n27501 = ~n27499 & ~n27500;
  assign n27502 = ~n27495 & ~n27496;
  assign n27503 = ~n27490 & ~n35276;
  assign n27504 = ~n27487 & ~n27488;
  assign n27505 = ~n1567 & ~n27504;
  assign n27506 = n1374 & ~n27505;
  assign n27507 = ~n27503 & ~n27505;
  assign n27508 = n1374 & n27507;
  assign n27509 = ~n27503 & n27506;
  assign n27510 = ~n26837 & ~n35277;
  assign n27511 = ~n1374 & ~n27507;
  assign n27512 = n1179 & ~n27511;
  assign n27513 = ~n27510 & n27512;
  assign n27514 = ~n26829 & ~n27513;
  assign n27515 = ~n27510 & ~n27511;
  assign n27516 = ~n1179 & ~n27515;
  assign n27517 = n1016 & ~n27516;
  assign n27518 = ~n27514 & ~n27516;
  assign n27519 = n1016 & n27518;
  assign n27520 = ~n27514 & n27517;
  assign n27521 = ~n26821 & ~n35278;
  assign n27522 = ~n1016 & ~n27518;
  assign n27523 = n855 & ~n27522;
  assign n27524 = ~n27521 & n27523;
  assign n27525 = ~n26597 & ~n35164;
  assign n27526 = ~n26597 & ~n26781;
  assign n27527 = ~n35164 & n27526;
  assign n27528 = ~n26781 & n27525;
  assign n27529 = n26605 & ~n35279;
  assign n27530 = n26609 & n27526;
  assign n27531 = ~n26597 & n26605;
  assign n27532 = ~n35164 & n27531;
  assign n27533 = ~n26781 & n27532;
  assign n27534 = ~n26605 & ~n35279;
  assign n27535 = ~n27533 & ~n27534;
  assign n27536 = ~n27529 & ~n27530;
  assign n27537 = ~n27524 & ~n35280;
  assign n27538 = ~n27521 & ~n27522;
  assign n27539 = ~n855 & ~n27538;
  assign n27540 = n720 & ~n27539;
  assign n27541 = ~n27537 & ~n27539;
  assign n27542 = n720 & n27541;
  assign n27543 = ~n27537 & n27540;
  assign n27544 = ~n26813 & ~n35281;
  assign n27545 = ~n720 & ~n27541;
  assign n27546 = n592 & ~n27545;
  assign n27547 = ~n27544 & n27546;
  assign n27548 = ~n26805 & ~n27547;
  assign n27549 = ~n27544 & ~n27545;
  assign n27550 = ~n592 & ~n27549;
  assign n27551 = n487 & ~n27550;
  assign n27552 = ~n27548 & ~n27550;
  assign n27553 = n487 & n27552;
  assign n27554 = ~n27548 & n27551;
  assign n27555 = ~n26797 & ~n35282;
  assign n27556 = ~n487 & ~n27552;
  assign n27557 = ~n27555 & ~n27556;
  assign n27558 = ~n393 & ~n27557;
  assign n27559 = n393 & ~n27556;
  assign n27560 = ~n27555 & n27559;
  assign n27561 = ~n26789 & ~n27560;
  assign n27562 = ~n27558 & ~n27561;
  assign n27563 = ~n321 & ~n27562;
  assign n27564 = ~n26675 & ~n26677;
  assign n27565 = ~n26781 & n27564;
  assign n27566 = ~n35174 & ~n27565;
  assign n27567 = ~n26677 & n35174;
  assign n27568 = ~n26675 & n27567;
  assign n27569 = n35174 & n27565;
  assign n27570 = ~n26781 & n27568;
  assign n27571 = ~n27566 & ~n35283;
  assign n27572 = n321 & ~n27558;
  assign n27573 = n321 & n27562;
  assign n27574 = ~n27561 & n27572;
  assign n27575 = ~n27571 & ~n35284;
  assign n27576 = ~n27563 & ~n27575;
  assign n27577 = ~n263 & ~n27576;
  assign n27578 = n263 & ~n27563;
  assign n27579 = ~n27575 & n27578;
  assign n27580 = ~n26692 & ~n35176;
  assign n27581 = ~n26692 & ~n26781;
  assign n27582 = ~n35176 & n27581;
  assign n27583 = ~n26781 & n27580;
  assign n27584 = n26700 & ~n35285;
  assign n27585 = n26704 & n27581;
  assign n27586 = ~n26692 & n26700;
  assign n27587 = ~n35176 & n27586;
  assign n27588 = ~n26781 & n27587;
  assign n27589 = ~n26700 & ~n35285;
  assign n27590 = ~n27588 & ~n27589;
  assign n27591 = ~n27584 & ~n27585;
  assign n27592 = ~n27579 & ~n35286;
  assign n27593 = ~n27577 & ~n27592;
  assign n27594 = ~n214 & ~n27593;
  assign n27595 = ~n26706 & ~n26708;
  assign n27596 = ~n26781 & n27595;
  assign n27597 = ~n35178 & ~n27596;
  assign n27598 = ~n26708 & n35178;
  assign n27599 = ~n26706 & n27598;
  assign n27600 = n35178 & n27596;
  assign n27601 = ~n26781 & n27599;
  assign n27602 = ~n27597 & ~n35287;
  assign n27603 = n214 & ~n27577;
  assign n27604 = n214 & n27593;
  assign n27605 = ~n27592 & n27603;
  assign n27606 = ~n27602 & ~n35288;
  assign n27607 = ~n27594 & ~n27606;
  assign n27608 = ~n197 & ~n27607;
  assign n27609 = n197 & ~n27594;
  assign n27610 = ~n27606 & n27609;
  assign n27611 = ~n26723 & ~n35180;
  assign n27612 = ~n26723 & ~n26781;
  assign n27613 = ~n35180 & n27612;
  assign n27614 = ~n26781 & n27611;
  assign n27615 = n26731 & ~n35289;
  assign n27616 = n26735 & n27612;
  assign n27617 = ~n26723 & n26731;
  assign n27618 = ~n35180 & n27617;
  assign n27619 = ~n26781 & n27618;
  assign n27620 = ~n26731 & ~n35289;
  assign n27621 = ~n27619 & ~n27620;
  assign n27622 = ~n27615 & ~n27616;
  assign n27623 = ~n27610 & ~n35290;
  assign n27624 = ~n27608 & ~n27623;
  assign n27625 = ~n26737 & ~n26739;
  assign n27626 = ~n26781 & n27625;
  assign n27627 = ~n35182 & ~n27626;
  assign n27628 = ~n26739 & n35182;
  assign n27629 = ~n26737 & n27628;
  assign n27630 = n35182 & n27626;
  assign n27631 = ~n26781 & n27629;
  assign n27632 = ~n27627 & ~n35291;
  assign n27633 = ~n26753 & ~n35184;
  assign n27634 = ~n35184 & ~n26781;
  assign n27635 = ~n26753 & n27634;
  assign n27636 = ~n26781 & n27633;
  assign n27637 = ~n35186 & ~n35292;
  assign n27638 = ~n27632 & n27637;
  assign n27639 = ~n27624 & n27638;
  assign n27640 = n193 & ~n27639;
  assign n27641 = ~n27608 & n27632;
  assign n27642 = n27624 & n27632;
  assign n27643 = ~n27623 & n27641;
  assign n27644 = n26753 & ~n27634;
  assign n27645 = ~n193 & ~n27633;
  assign n27646 = ~n27644 & n27645;
  assign n27647 = ~n35293 & ~n27646;
  assign n27648 = ~n27640 & n27647;
  assign n27649 = ~n27558 & ~n27560;
  assign n27650 = ~n27648 & n27649;
  assign n27651 = ~n26789 & ~n27650;
  assign n27652 = n26789 & ~n27558;
  assign n27653 = ~n27560 & n27652;
  assign n27654 = n26789 & n27650;
  assign n27655 = ~n27648 & n27653;
  assign n27656 = ~n27651 & ~n35294;
  assign n27657 = pi8  & ~n27648;
  assign n27658 = ~pi6  & ~pi7 ;
  assign n27659 = ~pi8  & n27658;
  assign n27660 = ~pi8  & ~n27658;
  assign n27661 = pi8  & n27648;
  assign n27662 = ~n27660 & ~n27661;
  assign n27663 = ~n27657 & ~n27659;
  assign n27664 = ~n26781 & n35295;
  assign n27665 = ~pi8  & ~n27648;
  assign n27666 = pi9  & ~n27665;
  assign n27667 = ~pi9  & n27665;
  assign n27668 = n27084 & ~n27648;
  assign n27669 = ~n27666 & ~n35296;
  assign n27670 = ~n26779 & ~n27659;
  assign n27671 = ~n35186 & n27670;
  assign n27672 = ~n26773 & n27671;
  assign n27673 = n26781 & ~n35295;
  assign n27674 = ~n27657 & n27672;
  assign n27675 = n27669 & ~n35297;
  assign n27676 = ~n27664 & ~n27675;
  assign n27677 = ~n25830 & ~n27676;
  assign n27678 = n25830 & ~n27664;
  assign n27679 = ~n27675 & n27678;
  assign n27680 = ~n26781 & ~n27646;
  assign n27681 = ~n35293 & n27680;
  assign n27682 = ~n26781 & n27648;
  assign n27683 = ~n27640 & n27681;
  assign n27684 = ~n35296 & ~n35298;
  assign n27685 = pi10  & ~n27684;
  assign n27686 = ~pi10  & ~n35298;
  assign n27687 = ~pi10  & n27684;
  assign n27688 = ~n35296 & n27686;
  assign n27689 = ~n27685 & ~n35299;
  assign n27690 = ~n27679 & ~n27689;
  assign n27691 = ~n27677 & ~n27690;
  assign n27692 = ~n24994 & ~n27691;
  assign n27693 = n24994 & ~n27677;
  assign n27694 = ~n27690 & n27693;
  assign n27695 = n24994 & n27691;
  assign n27696 = ~n35228 & ~n27105;
  assign n27697 = ~n27648 & n27696;
  assign n27698 = n27103 & ~n27697;
  assign n27699 = ~n27103 & n27696;
  assign n27700 = ~n27103 & n27697;
  assign n27701 = ~n27648 & n27699;
  assign n27702 = ~n27698 & ~n35301;
  assign n27703 = ~n35300 & ~n27702;
  assign n27704 = ~n27692 & ~n27703;
  assign n27705 = ~n24076 & ~n27704;
  assign n27706 = n24076 & ~n27692;
  assign n27707 = ~n27703 & n27706;
  assign n27708 = ~n35229 & ~n27111;
  assign n27709 = ~n27111 & ~n27648;
  assign n27710 = ~n35229 & n27709;
  assign n27711 = ~n27648 & n27708;
  assign n27712 = n27082 & ~n35302;
  assign n27713 = n27110 & n27709;
  assign n27714 = n27082 & ~n35229;
  assign n27715 = ~n27111 & n27714;
  assign n27716 = ~n27648 & n27715;
  assign n27717 = ~n27082 & ~n35302;
  assign n27718 = ~n27716 & ~n27717;
  assign n27719 = ~n27712 & ~n27713;
  assign n27720 = ~n27707 & ~n35303;
  assign n27721 = ~n27705 & ~n27720;
  assign n27722 = ~n23269 & ~n27721;
  assign n27723 = n23269 & ~n27705;
  assign n27724 = ~n27720 & n27723;
  assign n27725 = n23269 & n27721;
  assign n27726 = ~n27113 & ~n27123;
  assign n27727 = ~n27648 & n27726;
  assign n27728 = ~n27120 & ~n27727;
  assign n27729 = n27120 & ~n27123;
  assign n27730 = ~n27113 & n27729;
  assign n27731 = n27120 & n27727;
  assign n27732 = ~n27648 & n27730;
  assign n27733 = n27120 & ~n27727;
  assign n27734 = ~n27120 & n27727;
  assign n27735 = ~n27733 & ~n27734;
  assign n27736 = ~n27728 & ~n35305;
  assign n27737 = ~n35304 & n35306;
  assign n27738 = ~n27722 & ~n27737;
  assign n27739 = ~n22386 & ~n27738;
  assign n27740 = n22386 & ~n27722;
  assign n27741 = ~n27737 & n27740;
  assign n27742 = ~n35231 & ~n27129;
  assign n27743 = ~n27129 & ~n27648;
  assign n27744 = ~n35231 & n27743;
  assign n27745 = ~n27648 & n27742;
  assign n27746 = n27069 & ~n35307;
  assign n27747 = n27128 & n27743;
  assign n27748 = n27069 & ~n35231;
  assign n27749 = ~n27129 & n27748;
  assign n27750 = ~n27648 & n27749;
  assign n27751 = ~n27069 & ~n35307;
  assign n27752 = ~n27750 & ~n27751;
  assign n27753 = ~n27746 & ~n27747;
  assign n27754 = ~n27741 & ~n35308;
  assign n27755 = ~n27739 & ~n27754;
  assign n27756 = ~n21612 & ~n27755;
  assign n27757 = n21612 & ~n27739;
  assign n27758 = ~n27754 & n27757;
  assign n27759 = n21612 & n27755;
  assign n27760 = ~n27131 & ~n27145;
  assign n27761 = ~n27648 & n27760;
  assign n27762 = ~n35233 & ~n27761;
  assign n27763 = n35233 & n27761;
  assign n27764 = ~n35233 & ~n27145;
  assign n27765 = ~n27131 & n27764;
  assign n27766 = ~n27648 & n27765;
  assign n27767 = n35233 & ~n27761;
  assign n27768 = ~n27766 & ~n27767;
  assign n27769 = ~n27762 & ~n27763;
  assign n27770 = ~n35309 & ~n35310;
  assign n27771 = ~n27756 & ~n27770;
  assign n27772 = ~n20762 & ~n27771;
  assign n27773 = n20762 & ~n27756;
  assign n27774 = ~n27770 & n27773;
  assign n27775 = ~n35234 & ~n27151;
  assign n27776 = ~n27151 & ~n27648;
  assign n27777 = ~n35234 & n27776;
  assign n27778 = ~n27648 & n27775;
  assign n27779 = n27061 & ~n35311;
  assign n27780 = n27150 & n27776;
  assign n27781 = n27061 & ~n35234;
  assign n27782 = ~n27151 & n27781;
  assign n27783 = ~n27648 & n27782;
  assign n27784 = ~n27061 & ~n35311;
  assign n27785 = ~n27783 & ~n27784;
  assign n27786 = ~n27779 & ~n27780;
  assign n27787 = ~n27774 & ~n35312;
  assign n27788 = ~n27772 & ~n27787;
  assign n27789 = ~n20011 & ~n27788;
  assign n27790 = n20011 & ~n27772;
  assign n27791 = ~n27787 & n27790;
  assign n27792 = n20011 & n27788;
  assign n27793 = ~n27153 & ~n27166;
  assign n27794 = ~n27648 & n27793;
  assign n27795 = ~n35235 & n27794;
  assign n27796 = n35235 & ~n27794;
  assign n27797 = n35235 & ~n27166;
  assign n27798 = ~n27153 & n27797;
  assign n27799 = ~n27648 & n27798;
  assign n27800 = ~n35235 & ~n27794;
  assign n27801 = ~n27799 & ~n27800;
  assign n27802 = ~n27795 & ~n27796;
  assign n27803 = ~n35313 & ~n35314;
  assign n27804 = ~n27789 & ~n27803;
  assign n27805 = ~n19190 & ~n27804;
  assign n27806 = n19190 & ~n27789;
  assign n27807 = ~n27803 & n27806;
  assign n27808 = ~n35236 & ~n27172;
  assign n27809 = ~n27172 & ~n27648;
  assign n27810 = ~n35236 & n27809;
  assign n27811 = ~n27648 & n27808;
  assign n27812 = n27053 & ~n35315;
  assign n27813 = n27171 & n27809;
  assign n27814 = n27053 & ~n35236;
  assign n27815 = ~n27172 & n27814;
  assign n27816 = ~n27648 & n27815;
  assign n27817 = ~n27053 & ~n35315;
  assign n27818 = ~n27816 & ~n27817;
  assign n27819 = ~n27812 & ~n27813;
  assign n27820 = ~n27807 & ~n35316;
  assign n27821 = ~n27805 & ~n27820;
  assign n27822 = ~n18472 & ~n27821;
  assign n27823 = n18472 & ~n27805;
  assign n27824 = ~n27820 & n27823;
  assign n27825 = n18472 & n27821;
  assign n27826 = ~n27174 & ~n27187;
  assign n27827 = ~n27648 & n27826;
  assign n27828 = ~n35237 & n27827;
  assign n27829 = n35237 & ~n27827;
  assign n27830 = ~n35237 & ~n27827;
  assign n27831 = n35237 & ~n27187;
  assign n27832 = ~n27174 & n27831;
  assign n27833 = n35237 & n27827;
  assign n27834 = ~n27648 & n27832;
  assign n27835 = ~n27830 & ~n35318;
  assign n27836 = ~n27828 & ~n27829;
  assign n27837 = ~n35317 & ~n35319;
  assign n27838 = ~n27822 & ~n27837;
  assign n27839 = ~n17690 & ~n27838;
  assign n27840 = n17690 & ~n27822;
  assign n27841 = ~n27837 & n27840;
  assign n27842 = ~n35238 & ~n27193;
  assign n27843 = ~n27193 & ~n27648;
  assign n27844 = ~n35238 & n27843;
  assign n27845 = ~n27648 & n27842;
  assign n27846 = n27045 & ~n35320;
  assign n27847 = n27192 & n27843;
  assign n27848 = n27045 & ~n35238;
  assign n27849 = ~n27193 & n27848;
  assign n27850 = ~n27648 & n27849;
  assign n27851 = ~n27045 & ~n35320;
  assign n27852 = ~n27850 & ~n27851;
  assign n27853 = ~n27846 & ~n27847;
  assign n27854 = ~n27841 & ~n35321;
  assign n27855 = ~n27839 & ~n27854;
  assign n27856 = ~n17001 & ~n27855;
  assign n27857 = n17001 & ~n27839;
  assign n27858 = ~n27854 & n27857;
  assign n27859 = n17001 & n27855;
  assign n27860 = ~n27195 & ~n27209;
  assign n27861 = ~n27209 & ~n27648;
  assign n27862 = ~n27195 & n27861;
  assign n27863 = ~n27648 & n27860;
  assign n27864 = n35240 & ~n35323;
  assign n27865 = n27207 & n27861;
  assign n27866 = ~n35240 & n35323;
  assign n27867 = n35240 & ~n27209;
  assign n27868 = ~n27195 & n27867;
  assign n27869 = ~n27648 & n27868;
  assign n27870 = ~n35240 & ~n35323;
  assign n27871 = ~n27869 & ~n27870;
  assign n27872 = ~n27864 & ~n35324;
  assign n27873 = ~n35322 & ~n35325;
  assign n27874 = ~n27856 & ~n27873;
  assign n27875 = ~n16248 & ~n27874;
  assign n27876 = n16248 & ~n27856;
  assign n27877 = ~n27873 & n27876;
  assign n27878 = ~n35241 & ~n27215;
  assign n27879 = ~n27215 & ~n27648;
  assign n27880 = ~n35241 & n27879;
  assign n27881 = ~n27648 & n27878;
  assign n27882 = n27037 & ~n35326;
  assign n27883 = n27214 & n27879;
  assign n27884 = n27037 & ~n35241;
  assign n27885 = ~n27215 & n27884;
  assign n27886 = ~n27648 & n27885;
  assign n27887 = ~n27037 & ~n35326;
  assign n27888 = ~n27886 & ~n27887;
  assign n27889 = ~n27882 & ~n27883;
  assign n27890 = ~n27877 & ~n35327;
  assign n27891 = ~n27875 & ~n27890;
  assign n27892 = ~n15586 & ~n27891;
  assign n27893 = ~n27217 & ~n27233;
  assign n27894 = ~n27648 & n27893;
  assign n27895 = ~n35244 & ~n27894;
  assign n27896 = n35244 & ~n27233;
  assign n27897 = ~n27217 & n27896;
  assign n27898 = n35244 & n27894;
  assign n27899 = ~n27648 & n27897;
  assign n27900 = ~n27895 & ~n35328;
  assign n27901 = n15586 & ~n27875;
  assign n27902 = ~n27890 & n27901;
  assign n27903 = n15586 & n27891;
  assign n27904 = ~n27900 & ~n35329;
  assign n27905 = ~n27892 & ~n27904;
  assign n27906 = ~n14866 & ~n27905;
  assign n27907 = n14866 & ~n27892;
  assign n27908 = ~n27904 & n27907;
  assign n27909 = ~n35245 & ~n27239;
  assign n27910 = ~n27239 & ~n27648;
  assign n27911 = ~n35245 & n27910;
  assign n27912 = ~n27648 & n27909;
  assign n27913 = n27029 & ~n35330;
  assign n27914 = n27238 & n27910;
  assign n27915 = n27029 & ~n35245;
  assign n27916 = ~n27239 & n27915;
  assign n27917 = ~n27648 & n27916;
  assign n27918 = ~n27029 & ~n35330;
  assign n27919 = ~n27917 & ~n27918;
  assign n27920 = ~n27913 & ~n27914;
  assign n27921 = ~n27908 & ~n35331;
  assign n27922 = ~n27906 & ~n27921;
  assign n27923 = ~n14233 & ~n27922;
  assign n27924 = n14233 & ~n27906;
  assign n27925 = ~n27921 & n27924;
  assign n27926 = n14233 & n27922;
  assign n27927 = ~n27241 & ~n27244;
  assign n27928 = ~n27244 & ~n27648;
  assign n27929 = ~n27241 & n27928;
  assign n27930 = ~n27648 & n27927;
  assign n27931 = n27021 & ~n35333;
  assign n27932 = n27242 & n27928;
  assign n27933 = n27021 & ~n27244;
  assign n27934 = ~n27241 & n27933;
  assign n27935 = ~n27648 & n27934;
  assign n27936 = ~n27021 & ~n35333;
  assign n27937 = ~n27935 & ~n27936;
  assign n27938 = ~n27931 & ~n27932;
  assign n27939 = ~n35332 & ~n35334;
  assign n27940 = ~n27923 & ~n27939;
  assign n27941 = ~n13548 & ~n27940;
  assign n27942 = n13548 & ~n27923;
  assign n27943 = ~n27939 & n27942;
  assign n27944 = ~n35246 & ~n27250;
  assign n27945 = ~n27250 & ~n27648;
  assign n27946 = ~n35246 & n27945;
  assign n27947 = ~n27648 & n27944;
  assign n27948 = n27013 & ~n35335;
  assign n27949 = n27249 & n27945;
  assign n27950 = n27013 & ~n35246;
  assign n27951 = ~n27250 & n27950;
  assign n27952 = ~n27648 & n27951;
  assign n27953 = ~n27013 & ~n35335;
  assign n27954 = ~n27952 & ~n27953;
  assign n27955 = ~n27948 & ~n27949;
  assign n27956 = ~n27943 & ~n35336;
  assign n27957 = ~n27941 & ~n27956;
  assign n27958 = ~n12948 & ~n27957;
  assign n27959 = ~n27252 & ~n27267;
  assign n27960 = ~n27648 & n27959;
  assign n27961 = ~n35248 & ~n27960;
  assign n27962 = n35248 & ~n27267;
  assign n27963 = ~n27252 & n27962;
  assign n27964 = n35248 & n27960;
  assign n27965 = ~n27648 & n27963;
  assign n27966 = ~n27961 & ~n35337;
  assign n27967 = n12948 & ~n27941;
  assign n27968 = ~n27956 & n27967;
  assign n27969 = n12948 & n27957;
  assign n27970 = ~n27966 & ~n35338;
  assign n27971 = ~n27958 & ~n27970;
  assign n27972 = ~n12296 & ~n27971;
  assign n27973 = n12296 & ~n27958;
  assign n27974 = ~n27970 & n27973;
  assign n27975 = ~n35249 & ~n27273;
  assign n27976 = ~n27273 & ~n27648;
  assign n27977 = ~n35249 & n27976;
  assign n27978 = ~n27648 & n27975;
  assign n27979 = n27005 & ~n35339;
  assign n27980 = n27272 & n27976;
  assign n27981 = n27005 & ~n35249;
  assign n27982 = ~n27273 & n27981;
  assign n27983 = ~n27648 & n27982;
  assign n27984 = ~n27005 & ~n35339;
  assign n27985 = ~n27983 & ~n27984;
  assign n27986 = ~n27979 & ~n27980;
  assign n27987 = ~n27974 & ~n35340;
  assign n27988 = ~n27972 & ~n27987;
  assign n27989 = ~n11719 & ~n27988;
  assign n27990 = n11719 & ~n27972;
  assign n27991 = ~n27987 & n27990;
  assign n27992 = n11719 & n27988;
  assign n27993 = ~n27275 & ~n27278;
  assign n27994 = ~n27278 & ~n27648;
  assign n27995 = ~n27275 & n27994;
  assign n27996 = ~n27648 & n27993;
  assign n27997 = n26997 & ~n35342;
  assign n27998 = n27276 & n27994;
  assign n27999 = n26997 & ~n27278;
  assign n28000 = ~n27275 & n27999;
  assign n28001 = ~n27648 & n28000;
  assign n28002 = ~n26997 & ~n35342;
  assign n28003 = ~n28001 & ~n28002;
  assign n28004 = ~n27997 & ~n27998;
  assign n28005 = ~n35341 & ~n35343;
  assign n28006 = ~n27989 & ~n28005;
  assign n28007 = ~n11097 & ~n28006;
  assign n28008 = n11097 & ~n27989;
  assign n28009 = ~n28005 & n28008;
  assign n28010 = ~n35250 & ~n27284;
  assign n28011 = ~n27284 & ~n27648;
  assign n28012 = ~n35250 & n28011;
  assign n28013 = ~n27648 & n28010;
  assign n28014 = n26989 & ~n35344;
  assign n28015 = n27283 & n28011;
  assign n28016 = n26989 & ~n35250;
  assign n28017 = ~n27284 & n28016;
  assign n28018 = ~n27648 & n28017;
  assign n28019 = ~n26989 & ~n35344;
  assign n28020 = ~n28018 & ~n28019;
  assign n28021 = ~n28014 & ~n28015;
  assign n28022 = ~n28009 & ~n35345;
  assign n28023 = ~n28007 & ~n28022;
  assign n28024 = ~n10555 & ~n28023;
  assign n28025 = ~n27286 & ~n27301;
  assign n28026 = ~n27648 & n28025;
  assign n28027 = ~n35252 & ~n28026;
  assign n28028 = n35252 & ~n27301;
  assign n28029 = ~n27286 & n28028;
  assign n28030 = n35252 & n28026;
  assign n28031 = ~n27648 & n28029;
  assign n28032 = ~n28027 & ~n35346;
  assign n28033 = n10555 & ~n28007;
  assign n28034 = ~n28022 & n28033;
  assign n28035 = n10555 & n28023;
  assign n28036 = ~n28032 & ~n35347;
  assign n28037 = ~n28024 & ~n28036;
  assign n28038 = ~n9969 & ~n28037;
  assign n28039 = n9969 & ~n28024;
  assign n28040 = ~n28036 & n28039;
  assign n28041 = ~n35253 & ~n27307;
  assign n28042 = ~n27307 & ~n27648;
  assign n28043 = ~n35253 & n28042;
  assign n28044 = ~n27648 & n28041;
  assign n28045 = n26981 & ~n35348;
  assign n28046 = n27306 & n28042;
  assign n28047 = n26981 & ~n35253;
  assign n28048 = ~n27307 & n28047;
  assign n28049 = ~n27648 & n28048;
  assign n28050 = ~n26981 & ~n35348;
  assign n28051 = ~n28049 & ~n28050;
  assign n28052 = ~n28045 & ~n28046;
  assign n28053 = ~n28040 & ~n35349;
  assign n28054 = ~n28038 & ~n28053;
  assign n28055 = ~n9457 & ~n28054;
  assign n28056 = n9457 & ~n28038;
  assign n28057 = ~n28053 & n28056;
  assign n28058 = n9457 & n28054;
  assign n28059 = ~n27309 & ~n27312;
  assign n28060 = ~n27312 & ~n27648;
  assign n28061 = ~n27309 & n28060;
  assign n28062 = ~n27648 & n28059;
  assign n28063 = n26973 & ~n35351;
  assign n28064 = n27310 & n28060;
  assign n28065 = n26973 & ~n27312;
  assign n28066 = ~n27309 & n28065;
  assign n28067 = ~n27648 & n28066;
  assign n28068 = ~n26973 & ~n35351;
  assign n28069 = ~n28067 & ~n28068;
  assign n28070 = ~n28063 & ~n28064;
  assign n28071 = ~n35350 & ~n35352;
  assign n28072 = ~n28055 & ~n28071;
  assign n28073 = ~n8896 & ~n28072;
  assign n28074 = n8896 & ~n28055;
  assign n28075 = ~n28071 & n28074;
  assign n28076 = ~n35254 & ~n27318;
  assign n28077 = ~n27318 & ~n27648;
  assign n28078 = ~n35254 & n28077;
  assign n28079 = ~n27648 & n28076;
  assign n28080 = n26965 & ~n35353;
  assign n28081 = n27317 & n28077;
  assign n28082 = n26965 & ~n35254;
  assign n28083 = ~n27318 & n28082;
  assign n28084 = ~n27648 & n28083;
  assign n28085 = ~n26965 & ~n35353;
  assign n28086 = ~n28084 & ~n28085;
  assign n28087 = ~n28080 & ~n28081;
  assign n28088 = ~n28075 & ~n35354;
  assign n28089 = ~n28073 & ~n28088;
  assign n28090 = ~n8411 & ~n28089;
  assign n28091 = ~n27320 & ~n27335;
  assign n28092 = ~n27648 & n28091;
  assign n28093 = ~n35256 & ~n28092;
  assign n28094 = n35256 & ~n27335;
  assign n28095 = ~n27320 & n28094;
  assign n28096 = n35256 & n28092;
  assign n28097 = ~n27648 & n28095;
  assign n28098 = ~n28093 & ~n35355;
  assign n28099 = n8411 & ~n28073;
  assign n28100 = ~n28088 & n28099;
  assign n28101 = n8411 & n28089;
  assign n28102 = ~n28098 & ~n35356;
  assign n28103 = ~n28090 & ~n28102;
  assign n28104 = ~n7885 & ~n28103;
  assign n28105 = n7885 & ~n28090;
  assign n28106 = ~n28102 & n28105;
  assign n28107 = ~n35257 & ~n27341;
  assign n28108 = ~n27341 & ~n27648;
  assign n28109 = ~n35257 & n28108;
  assign n28110 = ~n27648 & n28107;
  assign n28111 = n26957 & ~n35357;
  assign n28112 = n27340 & n28108;
  assign n28113 = n26957 & ~n35257;
  assign n28114 = ~n27341 & n28113;
  assign n28115 = ~n27648 & n28114;
  assign n28116 = ~n26957 & ~n35357;
  assign n28117 = ~n28115 & ~n28116;
  assign n28118 = ~n28111 & ~n28112;
  assign n28119 = ~n28106 & ~n35358;
  assign n28120 = ~n28104 & ~n28119;
  assign n28121 = ~n7428 & ~n28120;
  assign n28122 = n7428 & ~n28104;
  assign n28123 = ~n28119 & n28122;
  assign n28124 = n7428 & n28120;
  assign n28125 = ~n27343 & ~n27346;
  assign n28126 = ~n27346 & ~n27648;
  assign n28127 = ~n27343 & n28126;
  assign n28128 = ~n27648 & n28125;
  assign n28129 = n26949 & ~n35360;
  assign n28130 = n27344 & n28126;
  assign n28131 = n26949 & ~n27346;
  assign n28132 = ~n27343 & n28131;
  assign n28133 = ~n27648 & n28132;
  assign n28134 = ~n26949 & ~n35360;
  assign n28135 = ~n28133 & ~n28134;
  assign n28136 = ~n28129 & ~n28130;
  assign n28137 = ~n35359 & ~n35361;
  assign n28138 = ~n28121 & ~n28137;
  assign n28139 = ~n6937 & ~n28138;
  assign n28140 = n6937 & ~n28121;
  assign n28141 = ~n28137 & n28140;
  assign n28142 = ~n35258 & ~n27352;
  assign n28143 = ~n27352 & ~n27648;
  assign n28144 = ~n35258 & n28143;
  assign n28145 = ~n27648 & n28142;
  assign n28146 = n26941 & ~n35362;
  assign n28147 = n27351 & n28143;
  assign n28148 = n26941 & ~n35258;
  assign n28149 = ~n27352 & n28148;
  assign n28150 = ~n27648 & n28149;
  assign n28151 = ~n26941 & ~n35362;
  assign n28152 = ~n28150 & ~n28151;
  assign n28153 = ~n28146 & ~n28147;
  assign n28154 = ~n28141 & ~n35363;
  assign n28155 = ~n28139 & ~n28154;
  assign n28156 = ~n6507 & ~n28155;
  assign n28157 = ~n27354 & ~n27369;
  assign n28158 = ~n27648 & n28157;
  assign n28159 = ~n35260 & ~n28158;
  assign n28160 = n35260 & ~n27369;
  assign n28161 = ~n27354 & n28160;
  assign n28162 = n35260 & n28158;
  assign n28163 = ~n27648 & n28161;
  assign n28164 = ~n28159 & ~n35364;
  assign n28165 = n6507 & ~n28139;
  assign n28166 = ~n28154 & n28165;
  assign n28167 = n6507 & n28155;
  assign n28168 = ~n28164 & ~n35365;
  assign n28169 = ~n28156 & ~n28168;
  assign n28170 = ~n6051 & ~n28169;
  assign n28171 = n6051 & ~n28156;
  assign n28172 = ~n28168 & n28171;
  assign n28173 = ~n35261 & ~n27375;
  assign n28174 = ~n27375 & ~n27648;
  assign n28175 = ~n35261 & n28174;
  assign n28176 = ~n27648 & n28173;
  assign n28177 = n26933 & ~n35366;
  assign n28178 = n27374 & n28174;
  assign n28179 = n26933 & ~n35261;
  assign n28180 = ~n27375 & n28179;
  assign n28181 = ~n27648 & n28180;
  assign n28182 = ~n26933 & ~n35366;
  assign n28183 = ~n28181 & ~n28182;
  assign n28184 = ~n28177 & ~n28178;
  assign n28185 = ~n28172 & ~n35367;
  assign n28186 = ~n28170 & ~n28185;
  assign n28187 = ~n5648 & ~n28186;
  assign n28188 = n5648 & ~n28170;
  assign n28189 = ~n28185 & n28188;
  assign n28190 = n5648 & n28186;
  assign n28191 = ~n27377 & ~n27380;
  assign n28192 = ~n27380 & ~n27648;
  assign n28193 = ~n27377 & n28192;
  assign n28194 = ~n27648 & n28191;
  assign n28195 = n26925 & ~n35369;
  assign n28196 = n27378 & n28192;
  assign n28197 = n26925 & ~n27380;
  assign n28198 = ~n27377 & n28197;
  assign n28199 = ~n27648 & n28198;
  assign n28200 = ~n26925 & ~n35369;
  assign n28201 = ~n28199 & ~n28200;
  assign n28202 = ~n28195 & ~n28196;
  assign n28203 = ~n35368 & ~n35370;
  assign n28204 = ~n28187 & ~n28203;
  assign n28205 = ~n5223 & ~n28204;
  assign n28206 = n5223 & ~n28187;
  assign n28207 = ~n28203 & n28206;
  assign n28208 = ~n35262 & ~n27386;
  assign n28209 = ~n27386 & ~n27648;
  assign n28210 = ~n35262 & n28209;
  assign n28211 = ~n27648 & n28208;
  assign n28212 = n26917 & ~n35371;
  assign n28213 = n27385 & n28209;
  assign n28214 = n26917 & ~n35262;
  assign n28215 = ~n27386 & n28214;
  assign n28216 = ~n27648 & n28215;
  assign n28217 = ~n26917 & ~n35371;
  assign n28218 = ~n28216 & ~n28217;
  assign n28219 = ~n28212 & ~n28213;
  assign n28220 = ~n28207 & ~n35372;
  assign n28221 = ~n28205 & ~n28220;
  assign n28222 = ~n4851 & ~n28221;
  assign n28223 = ~n27388 & ~n27403;
  assign n28224 = ~n27648 & n28223;
  assign n28225 = ~n35264 & ~n28224;
  assign n28226 = n35264 & ~n27403;
  assign n28227 = ~n27388 & n28226;
  assign n28228 = n35264 & n28224;
  assign n28229 = ~n27648 & n28227;
  assign n28230 = ~n28225 & ~n35373;
  assign n28231 = n4851 & ~n28205;
  assign n28232 = ~n28220 & n28231;
  assign n28233 = n4851 & n28221;
  assign n28234 = ~n28230 & ~n35374;
  assign n28235 = ~n28222 & ~n28234;
  assign n28236 = ~n4461 & ~n28235;
  assign n28237 = n4461 & ~n28222;
  assign n28238 = ~n28234 & n28237;
  assign n28239 = ~n35265 & ~n27409;
  assign n28240 = ~n27409 & ~n27648;
  assign n28241 = ~n35265 & n28240;
  assign n28242 = ~n27648 & n28239;
  assign n28243 = n26909 & ~n35375;
  assign n28244 = n27408 & n28240;
  assign n28245 = n26909 & ~n35265;
  assign n28246 = ~n27409 & n28245;
  assign n28247 = ~n27648 & n28246;
  assign n28248 = ~n26909 & ~n35375;
  assign n28249 = ~n28247 & ~n28248;
  assign n28250 = ~n28243 & ~n28244;
  assign n28251 = ~n28238 & ~n35376;
  assign n28252 = ~n28236 & ~n28251;
  assign n28253 = ~n4115 & ~n28252;
  assign n28254 = n4115 & ~n28236;
  assign n28255 = ~n28251 & n28254;
  assign n28256 = n4115 & n28252;
  assign n28257 = ~n27411 & ~n27414;
  assign n28258 = ~n27414 & ~n27648;
  assign n28259 = ~n27411 & n28258;
  assign n28260 = ~n27648 & n28257;
  assign n28261 = n26901 & ~n35378;
  assign n28262 = n27412 & n28258;
  assign n28263 = n26901 & ~n27414;
  assign n28264 = ~n27411 & n28263;
  assign n28265 = ~n27648 & n28264;
  assign n28266 = ~n26901 & ~n35378;
  assign n28267 = ~n28265 & ~n28266;
  assign n28268 = ~n28261 & ~n28262;
  assign n28269 = ~n35377 & ~n35379;
  assign n28270 = ~n28253 & ~n28269;
  assign n28271 = ~n3754 & ~n28270;
  assign n28272 = n3754 & ~n28253;
  assign n28273 = ~n28269 & n28272;
  assign n28274 = ~n35266 & ~n27420;
  assign n28275 = ~n27420 & ~n27648;
  assign n28276 = ~n35266 & n28275;
  assign n28277 = ~n27648 & n28274;
  assign n28278 = n26893 & ~n35380;
  assign n28279 = n27419 & n28275;
  assign n28280 = n26893 & ~n35266;
  assign n28281 = ~n27420 & n28280;
  assign n28282 = ~n27648 & n28281;
  assign n28283 = ~n26893 & ~n35380;
  assign n28284 = ~n28282 & ~n28283;
  assign n28285 = ~n28278 & ~n28279;
  assign n28286 = ~n28273 & ~n35381;
  assign n28287 = ~n28271 & ~n28286;
  assign n28288 = ~n3444 & ~n28287;
  assign n28289 = ~n27422 & ~n27437;
  assign n28290 = ~n27648 & n28289;
  assign n28291 = ~n35268 & ~n28290;
  assign n28292 = n35268 & ~n27437;
  assign n28293 = ~n27422 & n28292;
  assign n28294 = n35268 & n28290;
  assign n28295 = ~n27648 & n28293;
  assign n28296 = ~n28291 & ~n35382;
  assign n28297 = n3444 & ~n28271;
  assign n28298 = ~n28286 & n28297;
  assign n28299 = n3444 & n28287;
  assign n28300 = ~n28296 & ~n35383;
  assign n28301 = ~n28288 & ~n28300;
  assign n28302 = ~n3116 & ~n28301;
  assign n28303 = n3116 & ~n28288;
  assign n28304 = ~n28300 & n28303;
  assign n28305 = ~n35269 & ~n27443;
  assign n28306 = ~n27443 & ~n27648;
  assign n28307 = ~n35269 & n28306;
  assign n28308 = ~n27648 & n28305;
  assign n28309 = n26885 & ~n35384;
  assign n28310 = n27442 & n28306;
  assign n28311 = n26885 & ~n35269;
  assign n28312 = ~n27443 & n28311;
  assign n28313 = ~n27648 & n28312;
  assign n28314 = ~n26885 & ~n35384;
  assign n28315 = ~n28313 & ~n28314;
  assign n28316 = ~n28309 & ~n28310;
  assign n28317 = ~n28304 & ~n35385;
  assign n28318 = ~n28302 & ~n28317;
  assign n28319 = ~n2833 & ~n28318;
  assign n28320 = n2833 & ~n28302;
  assign n28321 = ~n28317 & n28320;
  assign n28322 = n2833 & n28318;
  assign n28323 = ~n27445 & ~n27448;
  assign n28324 = ~n27448 & ~n27648;
  assign n28325 = ~n27445 & n28324;
  assign n28326 = ~n27648 & n28323;
  assign n28327 = n26877 & ~n35387;
  assign n28328 = n27446 & n28324;
  assign n28329 = n26877 & ~n27448;
  assign n28330 = ~n27445 & n28329;
  assign n28331 = ~n27648 & n28330;
  assign n28332 = ~n26877 & ~n35387;
  assign n28333 = ~n28331 & ~n28332;
  assign n28334 = ~n28327 & ~n28328;
  assign n28335 = ~n35386 & ~n35388;
  assign n28336 = ~n28319 & ~n28335;
  assign n28337 = ~n2536 & ~n28336;
  assign n28338 = n2536 & ~n28319;
  assign n28339 = ~n28335 & n28338;
  assign n28340 = ~n35270 & ~n27454;
  assign n28341 = ~n27454 & ~n27648;
  assign n28342 = ~n35270 & n28341;
  assign n28343 = ~n27648 & n28340;
  assign n28344 = n26869 & ~n35389;
  assign n28345 = n27453 & n28341;
  assign n28346 = n26869 & ~n35270;
  assign n28347 = ~n27454 & n28346;
  assign n28348 = ~n27648 & n28347;
  assign n28349 = ~n26869 & ~n35389;
  assign n28350 = ~n28348 & ~n28349;
  assign n28351 = ~n28344 & ~n28345;
  assign n28352 = ~n28339 & ~n35390;
  assign n28353 = ~n28337 & ~n28352;
  assign n28354 = ~n2283 & ~n28353;
  assign n28355 = ~n27456 & ~n27471;
  assign n28356 = ~n27648 & n28355;
  assign n28357 = ~n35272 & ~n28356;
  assign n28358 = n35272 & ~n27471;
  assign n28359 = ~n27456 & n28358;
  assign n28360 = n35272 & n28356;
  assign n28361 = ~n27648 & n28359;
  assign n28362 = ~n28357 & ~n35391;
  assign n28363 = n2283 & ~n28337;
  assign n28364 = ~n28352 & n28363;
  assign n28365 = n2283 & n28353;
  assign n28366 = ~n28362 & ~n35392;
  assign n28367 = ~n28354 & ~n28366;
  assign n28368 = ~n2021 & ~n28367;
  assign n28369 = n2021 & ~n28354;
  assign n28370 = ~n28366 & n28369;
  assign n28371 = ~n35273 & ~n27477;
  assign n28372 = ~n27477 & ~n27648;
  assign n28373 = ~n35273 & n28372;
  assign n28374 = ~n27648 & n28371;
  assign n28375 = n26861 & ~n35393;
  assign n28376 = n27476 & n28372;
  assign n28377 = n26861 & ~n35273;
  assign n28378 = ~n27477 & n28377;
  assign n28379 = ~n27648 & n28378;
  assign n28380 = ~n26861 & ~n35393;
  assign n28381 = ~n28379 & ~n28380;
  assign n28382 = ~n28375 & ~n28376;
  assign n28383 = ~n28370 & ~n35394;
  assign n28384 = ~n28368 & ~n28383;
  assign n28385 = ~n1796 & ~n28384;
  assign n28386 = n1796 & ~n28368;
  assign n28387 = ~n28383 & n28386;
  assign n28388 = n1796 & n28384;
  assign n28389 = ~n27479 & ~n27482;
  assign n28390 = ~n27482 & ~n27648;
  assign n28391 = ~n27479 & n28390;
  assign n28392 = ~n27648 & n28389;
  assign n28393 = n26853 & ~n35396;
  assign n28394 = n27480 & n28390;
  assign n28395 = n26853 & ~n27482;
  assign n28396 = ~n27479 & n28395;
  assign n28397 = ~n27648 & n28396;
  assign n28398 = ~n26853 & ~n35396;
  assign n28399 = ~n28397 & ~n28398;
  assign n28400 = ~n28393 & ~n28394;
  assign n28401 = ~n35395 & ~n35397;
  assign n28402 = ~n28385 & ~n28401;
  assign n28403 = ~n1567 & ~n28402;
  assign n28404 = n1567 & ~n28385;
  assign n28405 = ~n28401 & n28404;
  assign n28406 = ~n35274 & ~n27488;
  assign n28407 = ~n27488 & ~n27648;
  assign n28408 = ~n35274 & n28407;
  assign n28409 = ~n27648 & n28406;
  assign n28410 = n26845 & ~n35398;
  assign n28411 = n27487 & n28407;
  assign n28412 = n26845 & ~n35274;
  assign n28413 = ~n27488 & n28412;
  assign n28414 = ~n27648 & n28413;
  assign n28415 = ~n26845 & ~n35398;
  assign n28416 = ~n28414 & ~n28415;
  assign n28417 = ~n28410 & ~n28411;
  assign n28418 = ~n28405 & ~n35399;
  assign n28419 = ~n28403 & ~n28418;
  assign n28420 = ~n1374 & ~n28419;
  assign n28421 = ~n27490 & ~n27505;
  assign n28422 = ~n27648 & n28421;
  assign n28423 = ~n35276 & ~n28422;
  assign n28424 = n35276 & ~n27505;
  assign n28425 = ~n27490 & n28424;
  assign n28426 = n35276 & n28422;
  assign n28427 = ~n27648 & n28425;
  assign n28428 = ~n28423 & ~n35400;
  assign n28429 = n1374 & ~n28403;
  assign n28430 = ~n28418 & n28429;
  assign n28431 = n1374 & n28419;
  assign n28432 = ~n28428 & ~n35401;
  assign n28433 = ~n28420 & ~n28432;
  assign n28434 = ~n1179 & ~n28433;
  assign n28435 = n1179 & ~n28420;
  assign n28436 = ~n28432 & n28435;
  assign n28437 = ~n35277 & ~n27511;
  assign n28438 = ~n27511 & ~n27648;
  assign n28439 = ~n35277 & n28438;
  assign n28440 = ~n27648 & n28437;
  assign n28441 = n26837 & ~n35402;
  assign n28442 = n27510 & n28438;
  assign n28443 = n26837 & ~n35277;
  assign n28444 = ~n27511 & n28443;
  assign n28445 = ~n27648 & n28444;
  assign n28446 = ~n26837 & ~n35402;
  assign n28447 = ~n28445 & ~n28446;
  assign n28448 = ~n28441 & ~n28442;
  assign n28449 = ~n28436 & ~n35403;
  assign n28450 = ~n28434 & ~n28449;
  assign n28451 = ~n1016 & ~n28450;
  assign n28452 = n1016 & ~n28434;
  assign n28453 = ~n28449 & n28452;
  assign n28454 = n1016 & n28450;
  assign n28455 = ~n27513 & ~n27516;
  assign n28456 = ~n27516 & ~n27648;
  assign n28457 = ~n27513 & n28456;
  assign n28458 = ~n27648 & n28455;
  assign n28459 = n26829 & ~n35405;
  assign n28460 = n27514 & n28456;
  assign n28461 = n26829 & ~n27516;
  assign n28462 = ~n27513 & n28461;
  assign n28463 = ~n27648 & n28462;
  assign n28464 = ~n26829 & ~n35405;
  assign n28465 = ~n28463 & ~n28464;
  assign n28466 = ~n28459 & ~n28460;
  assign n28467 = ~n35404 & ~n35406;
  assign n28468 = ~n28451 & ~n28467;
  assign n28469 = ~n855 & ~n28468;
  assign n28470 = n855 & ~n28451;
  assign n28471 = ~n28467 & n28470;
  assign n28472 = ~n35278 & ~n27522;
  assign n28473 = ~n27522 & ~n27648;
  assign n28474 = ~n35278 & n28473;
  assign n28475 = ~n27648 & n28472;
  assign n28476 = n26821 & ~n35407;
  assign n28477 = n27521 & n28473;
  assign n28478 = n26821 & ~n35278;
  assign n28479 = ~n27522 & n28478;
  assign n28480 = ~n27648 & n28479;
  assign n28481 = ~n26821 & ~n35407;
  assign n28482 = ~n28480 & ~n28481;
  assign n28483 = ~n28476 & ~n28477;
  assign n28484 = ~n28471 & ~n35408;
  assign n28485 = ~n28469 & ~n28484;
  assign n28486 = ~n720 & ~n28485;
  assign n28487 = ~n27524 & ~n27539;
  assign n28488 = ~n27648 & n28487;
  assign n28489 = ~n35280 & ~n28488;
  assign n28490 = n35280 & ~n27539;
  assign n28491 = ~n27524 & n28490;
  assign n28492 = n35280 & n28488;
  assign n28493 = ~n27648 & n28491;
  assign n28494 = ~n28489 & ~n35409;
  assign n28495 = n720 & ~n28469;
  assign n28496 = ~n28484 & n28495;
  assign n28497 = n720 & n28485;
  assign n28498 = ~n28494 & ~n35410;
  assign n28499 = ~n28486 & ~n28498;
  assign n28500 = ~n592 & ~n28499;
  assign n28501 = n592 & ~n28486;
  assign n28502 = ~n28498 & n28501;
  assign n28503 = ~n35281 & ~n27545;
  assign n28504 = ~n27545 & ~n27648;
  assign n28505 = ~n35281 & n28504;
  assign n28506 = ~n27648 & n28503;
  assign n28507 = n26813 & ~n35411;
  assign n28508 = n27544 & n28504;
  assign n28509 = n26813 & ~n35281;
  assign n28510 = ~n27545 & n28509;
  assign n28511 = ~n27648 & n28510;
  assign n28512 = ~n26813 & ~n35411;
  assign n28513 = ~n28511 & ~n28512;
  assign n28514 = ~n28507 & ~n28508;
  assign n28515 = ~n28502 & ~n35412;
  assign n28516 = ~n28500 & ~n28515;
  assign n28517 = ~n487 & ~n28516;
  assign n28518 = n487 & ~n28500;
  assign n28519 = ~n28515 & n28518;
  assign n28520 = n487 & n28516;
  assign n28521 = ~n27547 & ~n27550;
  assign n28522 = ~n27550 & ~n27648;
  assign n28523 = ~n27547 & n28522;
  assign n28524 = ~n27648 & n28521;
  assign n28525 = n26805 & ~n35414;
  assign n28526 = n27548 & n28522;
  assign n28527 = n26805 & ~n27550;
  assign n28528 = ~n27547 & n28527;
  assign n28529 = ~n27648 & n28528;
  assign n28530 = ~n26805 & ~n35414;
  assign n28531 = ~n28529 & ~n28530;
  assign n28532 = ~n28525 & ~n28526;
  assign n28533 = ~n35413 & ~n35415;
  assign n28534 = ~n28517 & ~n28533;
  assign n28535 = ~n393 & ~n28534;
  assign n28536 = n393 & ~n28517;
  assign n28537 = ~n28533 & n28536;
  assign n28538 = n26797 & ~n35282;
  assign n28539 = ~n27556 & n28538;
  assign n28540 = ~n35282 & ~n27556;
  assign n28541 = ~n27648 & n28540;
  assign n28542 = n26797 & n28541;
  assign n28543 = ~n27648 & n28539;
  assign n28544 = ~n26797 & ~n28541;
  assign n28545 = ~n35416 & ~n28544;
  assign n28546 = ~n28537 & ~n28545;
  assign n28547 = ~n28535 & ~n28546;
  assign n28548 = ~n321 & ~n28547;
  assign n28549 = n321 & ~n28535;
  assign n28550 = ~n28546 & n28549;
  assign n28551 = n321 & n28547;
  assign n28552 = ~n27656 & ~n35417;
  assign n28553 = ~n28548 & ~n28552;
  assign n28554 = ~n263 & ~n28553;
  assign n28555 = n263 & ~n28548;
  assign n28556 = ~n28552 & n28555;
  assign n28557 = ~n27563 & ~n35284;
  assign n28558 = ~n27563 & ~n27648;
  assign n28559 = ~n35284 & n28558;
  assign n28560 = ~n27648 & n28557;
  assign n28561 = n27571 & ~n35418;
  assign n28562 = n27575 & n28558;
  assign n28563 = n27571 & ~n35284;
  assign n28564 = ~n27563 & n28563;
  assign n28565 = ~n27648 & n28564;
  assign n28566 = ~n27571 & ~n35418;
  assign n28567 = ~n28565 & ~n28566;
  assign n28568 = ~n28561 & ~n28562;
  assign n28569 = ~n28556 & ~n35419;
  assign n28570 = ~n28554 & ~n28569;
  assign n28571 = ~n214 & ~n28570;
  assign n28572 = ~n27577 & ~n27579;
  assign n28573 = ~n27648 & n28572;
  assign n28574 = ~n35286 & ~n28573;
  assign n28575 = ~n27577 & n35286;
  assign n28576 = ~n27579 & n28575;
  assign n28577 = n35286 & n28573;
  assign n28578 = ~n27648 & n28576;
  assign n28579 = ~n28574 & ~n35420;
  assign n28580 = n214 & ~n28554;
  assign n28581 = ~n28569 & n28580;
  assign n28582 = n214 & n28570;
  assign n28583 = ~n28579 & ~n35421;
  assign n28584 = ~n28571 & ~n28583;
  assign n28585 = ~n197 & ~n28584;
  assign n28586 = n197 & ~n28571;
  assign n28587 = ~n28583 & n28586;
  assign n28588 = ~n27594 & ~n35288;
  assign n28589 = ~n27594 & ~n27648;
  assign n28590 = ~n35288 & n28589;
  assign n28591 = ~n27648 & n28588;
  assign n28592 = n27602 & ~n35422;
  assign n28593 = n27606 & n28589;
  assign n28594 = n27602 & ~n35288;
  assign n28595 = ~n27594 & n28594;
  assign n28596 = ~n27648 & n28595;
  assign n28597 = ~n27602 & ~n35422;
  assign n28598 = ~n28596 & ~n28597;
  assign n28599 = ~n28592 & ~n28593;
  assign n28600 = ~n28587 & ~n35423;
  assign n28601 = ~n28585 & ~n28600;
  assign n28602 = ~n27608 & ~n27610;
  assign n28603 = ~n27648 & n28602;
  assign n28604 = ~n35290 & ~n28603;
  assign n28605 = ~n27608 & n35290;
  assign n28606 = ~n27610 & n28605;
  assign n28607 = n35290 & n28603;
  assign n28608 = ~n27648 & n28606;
  assign n28609 = ~n28604 & ~n35424;
  assign n28610 = ~n27624 & ~n27632;
  assign n28611 = ~n27632 & ~n27648;
  assign n28612 = ~n27624 & n28611;
  assign n28613 = ~n27648 & n28610;
  assign n28614 = ~n35293 & ~n35425;
  assign n28615 = ~n28609 & n28614;
  assign n28616 = ~n28601 & n28615;
  assign n28617 = n193 & ~n28616;
  assign n28618 = ~n28585 & n28609;
  assign n28619 = ~n28600 & n28618;
  assign n28620 = n28601 & n28609;
  assign n28621 = n27624 & ~n28611;
  assign n28622 = ~n193 & ~n28610;
  assign n28623 = ~n28621 & n28622;
  assign n28624 = ~n35426 & ~n28623;
  assign n28625 = ~n28617 & n28624;
  assign n28626 = ~n28548 & ~n35417;
  assign n28627 = ~n28625 & n28626;
  assign n28628 = n27656 & ~n28627;
  assign n28629 = ~n27656 & n28627;
  assign n28630 = n27656 & ~n28548;
  assign n28631 = ~n35417 & n28630;
  assign n28632 = ~n28625 & n28631;
  assign n28633 = ~n27656 & ~n28627;
  assign n28634 = ~n28632 & ~n28633;
  assign n28635 = ~n28628 & ~n28629;
  assign n28636 = ~n28535 & ~n28537;
  assign n28637 = ~n28625 & n28636;
  assign n28638 = ~n28545 & ~n28637;
  assign n28639 = ~n28537 & n28545;
  assign n28640 = ~n28535 & n28639;
  assign n28641 = n28545 & n28637;
  assign n28642 = ~n28625 & n28640;
  assign n28643 = ~n28638 & ~n35428;
  assign n28644 = ~n28517 & ~n35413;
  assign n28645 = ~n28625 & n28644;
  assign n28646 = ~n35415 & ~n28645;
  assign n28647 = ~n28517 & n35415;
  assign n28648 = ~n35413 & n28647;
  assign n28649 = n35415 & n28645;
  assign n28650 = ~n28625 & n28648;
  assign n28651 = ~n28646 & ~n35429;
  assign n28652 = ~n28500 & ~n28502;
  assign n28653 = ~n28625 & n28652;
  assign n28654 = ~n35412 & ~n28653;
  assign n28655 = ~n28502 & n35412;
  assign n28656 = ~n28500 & n28655;
  assign n28657 = n35412 & n28653;
  assign n28658 = ~n28625 & n28656;
  assign n28659 = ~n28654 & ~n35430;
  assign n28660 = ~n28469 & ~n28471;
  assign n28661 = ~n28625 & n28660;
  assign n28662 = ~n35408 & ~n28661;
  assign n28663 = ~n28471 & n35408;
  assign n28664 = ~n28469 & n28663;
  assign n28665 = n35408 & n28661;
  assign n28666 = ~n28625 & n28664;
  assign n28667 = ~n28662 & ~n35431;
  assign n28668 = ~n28451 & ~n35404;
  assign n28669 = ~n28625 & n28668;
  assign n28670 = ~n35406 & ~n28669;
  assign n28671 = ~n28451 & n35406;
  assign n28672 = ~n35404 & n28671;
  assign n28673 = n35406 & n28669;
  assign n28674 = ~n28625 & n28672;
  assign n28675 = ~n28670 & ~n35432;
  assign n28676 = ~n28434 & ~n28436;
  assign n28677 = ~n28625 & n28676;
  assign n28678 = ~n35403 & ~n28677;
  assign n28679 = ~n28436 & n35403;
  assign n28680 = ~n28434 & n28679;
  assign n28681 = n35403 & n28677;
  assign n28682 = ~n28625 & n28680;
  assign n28683 = ~n28678 & ~n35433;
  assign n28684 = ~n28403 & ~n28405;
  assign n28685 = ~n28625 & n28684;
  assign n28686 = ~n35399 & ~n28685;
  assign n28687 = ~n28405 & n35399;
  assign n28688 = ~n28403 & n28687;
  assign n28689 = n35399 & n28685;
  assign n28690 = ~n28625 & n28688;
  assign n28691 = ~n28686 & ~n35434;
  assign n28692 = ~n28385 & ~n35395;
  assign n28693 = ~n28625 & n28692;
  assign n28694 = ~n35397 & ~n28693;
  assign n28695 = ~n28385 & n35397;
  assign n28696 = ~n35395 & n28695;
  assign n28697 = n35397 & n28693;
  assign n28698 = ~n28625 & n28696;
  assign n28699 = ~n28694 & ~n35435;
  assign n28700 = ~n28368 & ~n28370;
  assign n28701 = ~n28625 & n28700;
  assign n28702 = ~n35394 & ~n28701;
  assign n28703 = ~n28370 & n35394;
  assign n28704 = ~n28368 & n28703;
  assign n28705 = n35394 & n28701;
  assign n28706 = ~n28625 & n28704;
  assign n28707 = ~n28702 & ~n35436;
  assign n28708 = ~n28337 & ~n28339;
  assign n28709 = ~n28625 & n28708;
  assign n28710 = ~n35390 & ~n28709;
  assign n28711 = ~n28339 & n35390;
  assign n28712 = ~n28337 & n28711;
  assign n28713 = n35390 & n28709;
  assign n28714 = ~n28625 & n28712;
  assign n28715 = ~n28710 & ~n35437;
  assign n28716 = ~n28319 & ~n35386;
  assign n28717 = ~n28625 & n28716;
  assign n28718 = ~n35388 & ~n28717;
  assign n28719 = ~n28319 & n35388;
  assign n28720 = ~n35386 & n28719;
  assign n28721 = n35388 & n28717;
  assign n28722 = ~n28625 & n28720;
  assign n28723 = ~n28718 & ~n35438;
  assign n28724 = ~n28302 & ~n28304;
  assign n28725 = ~n28625 & n28724;
  assign n28726 = ~n35385 & ~n28725;
  assign n28727 = ~n28304 & n35385;
  assign n28728 = ~n28302 & n28727;
  assign n28729 = n35385 & n28725;
  assign n28730 = ~n28625 & n28728;
  assign n28731 = ~n28726 & ~n35439;
  assign n28732 = ~n28271 & ~n28273;
  assign n28733 = ~n28625 & n28732;
  assign n28734 = ~n35381 & ~n28733;
  assign n28735 = ~n28273 & n35381;
  assign n28736 = ~n28271 & n28735;
  assign n28737 = n35381 & n28733;
  assign n28738 = ~n28625 & n28736;
  assign n28739 = ~n28734 & ~n35440;
  assign n28740 = ~n28253 & ~n35377;
  assign n28741 = ~n28625 & n28740;
  assign n28742 = ~n35379 & ~n28741;
  assign n28743 = ~n28253 & n35379;
  assign n28744 = ~n35377 & n28743;
  assign n28745 = n35379 & n28741;
  assign n28746 = ~n28625 & n28744;
  assign n28747 = ~n28742 & ~n35441;
  assign n28748 = ~n28236 & ~n28238;
  assign n28749 = ~n28625 & n28748;
  assign n28750 = ~n35376 & ~n28749;
  assign n28751 = ~n28238 & n35376;
  assign n28752 = ~n28236 & n28751;
  assign n28753 = n35376 & n28749;
  assign n28754 = ~n28625 & n28752;
  assign n28755 = ~n28750 & ~n35442;
  assign n28756 = ~n28205 & ~n28207;
  assign n28757 = ~n28625 & n28756;
  assign n28758 = ~n35372 & ~n28757;
  assign n28759 = ~n28207 & n35372;
  assign n28760 = ~n28205 & n28759;
  assign n28761 = n35372 & n28757;
  assign n28762 = ~n28625 & n28760;
  assign n28763 = ~n28758 & ~n35443;
  assign n28764 = ~n28187 & ~n35368;
  assign n28765 = ~n28625 & n28764;
  assign n28766 = ~n35370 & ~n28765;
  assign n28767 = ~n28187 & n35370;
  assign n28768 = ~n35368 & n28767;
  assign n28769 = n35370 & n28765;
  assign n28770 = ~n28625 & n28768;
  assign n28771 = ~n28766 & ~n35444;
  assign n28772 = ~n28170 & ~n28172;
  assign n28773 = ~n28625 & n28772;
  assign n28774 = ~n35367 & ~n28773;
  assign n28775 = ~n28172 & n35367;
  assign n28776 = ~n28170 & n28775;
  assign n28777 = n35367 & n28773;
  assign n28778 = ~n28625 & n28776;
  assign n28779 = ~n28774 & ~n35445;
  assign n28780 = ~n28139 & ~n28141;
  assign n28781 = ~n28625 & n28780;
  assign n28782 = ~n35363 & ~n28781;
  assign n28783 = ~n28141 & n35363;
  assign n28784 = ~n28139 & n28783;
  assign n28785 = n35363 & n28781;
  assign n28786 = ~n28625 & n28784;
  assign n28787 = ~n28782 & ~n35446;
  assign n28788 = ~n28121 & ~n35359;
  assign n28789 = ~n28625 & n28788;
  assign n28790 = ~n35361 & ~n28789;
  assign n28791 = ~n28121 & n35361;
  assign n28792 = ~n35359 & n28791;
  assign n28793 = n35361 & n28789;
  assign n28794 = ~n28625 & n28792;
  assign n28795 = ~n28790 & ~n35447;
  assign n28796 = ~n28104 & ~n28106;
  assign n28797 = ~n28625 & n28796;
  assign n28798 = ~n35358 & ~n28797;
  assign n28799 = ~n28106 & n35358;
  assign n28800 = ~n28104 & n28799;
  assign n28801 = n35358 & n28797;
  assign n28802 = ~n28625 & n28800;
  assign n28803 = ~n28798 & ~n35448;
  assign n28804 = ~n28073 & ~n28075;
  assign n28805 = ~n28625 & n28804;
  assign n28806 = ~n35354 & ~n28805;
  assign n28807 = ~n28075 & n35354;
  assign n28808 = ~n28073 & n28807;
  assign n28809 = n35354 & n28805;
  assign n28810 = ~n28625 & n28808;
  assign n28811 = ~n28806 & ~n35449;
  assign n28812 = ~n28055 & ~n35350;
  assign n28813 = ~n28625 & n28812;
  assign n28814 = ~n35352 & ~n28813;
  assign n28815 = ~n28055 & n35352;
  assign n28816 = ~n35350 & n28815;
  assign n28817 = n35352 & n28813;
  assign n28818 = ~n28625 & n28816;
  assign n28819 = ~n28814 & ~n35450;
  assign n28820 = ~n28038 & ~n28040;
  assign n28821 = ~n28625 & n28820;
  assign n28822 = ~n35349 & ~n28821;
  assign n28823 = ~n28040 & n35349;
  assign n28824 = ~n28038 & n28823;
  assign n28825 = n35349 & n28821;
  assign n28826 = ~n28625 & n28824;
  assign n28827 = ~n28822 & ~n35451;
  assign n28828 = ~n28007 & ~n28009;
  assign n28829 = ~n28625 & n28828;
  assign n28830 = ~n35345 & ~n28829;
  assign n28831 = ~n28009 & n35345;
  assign n28832 = ~n28007 & n28831;
  assign n28833 = n35345 & n28829;
  assign n28834 = ~n28625 & n28832;
  assign n28835 = ~n28830 & ~n35452;
  assign n28836 = ~n27989 & ~n35341;
  assign n28837 = ~n28625 & n28836;
  assign n28838 = ~n35343 & ~n28837;
  assign n28839 = ~n27989 & n35343;
  assign n28840 = ~n35341 & n28839;
  assign n28841 = n35343 & n28837;
  assign n28842 = ~n28625 & n28840;
  assign n28843 = ~n28838 & ~n35453;
  assign n28844 = ~n27972 & ~n27974;
  assign n28845 = ~n28625 & n28844;
  assign n28846 = ~n35340 & ~n28845;
  assign n28847 = ~n27974 & n35340;
  assign n28848 = ~n27972 & n28847;
  assign n28849 = n35340 & n28845;
  assign n28850 = ~n28625 & n28848;
  assign n28851 = ~n28846 & ~n35454;
  assign n28852 = ~n27941 & ~n27943;
  assign n28853 = ~n28625 & n28852;
  assign n28854 = ~n35336 & ~n28853;
  assign n28855 = ~n27943 & n35336;
  assign n28856 = ~n27941 & n28855;
  assign n28857 = n35336 & n28853;
  assign n28858 = ~n28625 & n28856;
  assign n28859 = ~n28854 & ~n35455;
  assign n28860 = ~n27923 & ~n35332;
  assign n28861 = ~n28625 & n28860;
  assign n28862 = ~n35334 & ~n28861;
  assign n28863 = ~n27923 & n35334;
  assign n28864 = ~n35332 & n28863;
  assign n28865 = n35334 & n28861;
  assign n28866 = ~n28625 & n28864;
  assign n28867 = ~n28862 & ~n35456;
  assign n28868 = ~n27906 & ~n27908;
  assign n28869 = ~n28625 & n28868;
  assign n28870 = ~n35331 & ~n28869;
  assign n28871 = ~n27908 & n35331;
  assign n28872 = ~n27906 & n28871;
  assign n28873 = n35331 & n28869;
  assign n28874 = ~n28625 & n28872;
  assign n28875 = ~n28870 & ~n35457;
  assign n28876 = ~n27875 & ~n27877;
  assign n28877 = ~n28625 & n28876;
  assign n28878 = ~n35327 & ~n28877;
  assign n28879 = ~n27877 & n35327;
  assign n28880 = ~n27875 & n28879;
  assign n28881 = n35327 & n28877;
  assign n28882 = ~n28625 & n28880;
  assign n28883 = ~n28878 & ~n35458;
  assign n28884 = ~n27856 & ~n35322;
  assign n28885 = ~n28625 & n28884;
  assign n28886 = ~n35325 & ~n28885;
  assign n28887 = ~n27856 & n35325;
  assign n28888 = ~n35322 & n28887;
  assign n28889 = n35325 & n28885;
  assign n28890 = ~n28625 & n28888;
  assign n28891 = ~n28886 & ~n35459;
  assign n28892 = ~n27839 & ~n27841;
  assign n28893 = ~n28625 & n28892;
  assign n28894 = ~n35321 & ~n28893;
  assign n28895 = ~n27841 & n35321;
  assign n28896 = ~n27839 & n28895;
  assign n28897 = n35321 & n28893;
  assign n28898 = ~n28625 & n28896;
  assign n28899 = ~n28894 & ~n35460;
  assign n28900 = ~n27805 & ~n27807;
  assign n28901 = ~n28625 & n28900;
  assign n28902 = ~n35316 & ~n28901;
  assign n28903 = ~n27807 & n35316;
  assign n28904 = ~n27805 & n28903;
  assign n28905 = n35316 & n28901;
  assign n28906 = ~n28625 & n28904;
  assign n28907 = ~n28902 & ~n35461;
  assign n28908 = ~n27772 & ~n27774;
  assign n28909 = ~n28625 & n28908;
  assign n28910 = ~n35312 & ~n28909;
  assign n28911 = ~n27774 & n35312;
  assign n28912 = ~n27772 & n28911;
  assign n28913 = n35312 & n28909;
  assign n28914 = ~n28625 & n28912;
  assign n28915 = ~n28910 & ~n35462;
  assign n28916 = ~n27739 & ~n27741;
  assign n28917 = ~n28625 & n28916;
  assign n28918 = ~n35308 & ~n28917;
  assign n28919 = ~n27741 & n35308;
  assign n28920 = ~n27739 & n28919;
  assign n28921 = n35308 & n28917;
  assign n28922 = ~n28625 & n28920;
  assign n28923 = ~n28918 & ~n35463;
  assign n28924 = ~n27705 & ~n27707;
  assign n28925 = ~n28625 & n28924;
  assign n28926 = ~n35303 & ~n28925;
  assign n28927 = ~n27707 & n35303;
  assign n28928 = ~n27705 & n28927;
  assign n28929 = n35303 & n28925;
  assign n28930 = ~n28625 & n28928;
  assign n28931 = ~n28926 & ~n35464;
  assign n28932 = ~n27677 & ~n27679;
  assign n28933 = ~n28625 & n28932;
  assign n28934 = ~n27689 & ~n28933;
  assign n28935 = ~n27679 & n27689;
  assign n28936 = ~n27677 & n28935;
  assign n28937 = n27689 & n28933;
  assign n28938 = ~n28625 & n28936;
  assign n28939 = ~n28934 & ~n35465;
  assign n28940 = ~pi6  & ~n28625;
  assign n28941 = ~pi7  & n28940;
  assign n28942 = n27658 & ~n28625;
  assign n28943 = ~n27648 & ~n28623;
  assign n28944 = ~n35426 & n28943;
  assign n28945 = ~n27648 & n28625;
  assign n28946 = ~n28617 & n28944;
  assign n28947 = ~n35466 & ~n35467;
  assign n28948 = pi8  & ~n28947;
  assign n28949 = ~pi8  & ~n35467;
  assign n28950 = ~pi8  & n28947;
  assign n28951 = ~n35466 & n28949;
  assign n28952 = ~n28948 & ~n35468;
  assign n28953 = pi6  & ~n28625;
  assign n28954 = ~pi4  & ~pi5 ;
  assign n28955 = ~pi6  & n28954;
  assign n28956 = ~n27646 & ~n28955;
  assign n28957 = ~n35293 & n28956;
  assign n28958 = ~n27640 & n28957;
  assign n28959 = ~pi6  & ~n28954;
  assign n28960 = pi6  & n28625;
  assign n28961 = ~n28959 & ~n28960;
  assign n28962 = ~n28953 & ~n28955;
  assign n28963 = n27648 & ~n35469;
  assign n28964 = ~n28953 & n28958;
  assign n28965 = pi7  & ~n28940;
  assign n28966 = ~n35466 & ~n28965;
  assign n28967 = ~n35470 & n28966;
  assign n28968 = ~n27648 & n35469;
  assign n28969 = n26781 & ~n28968;
  assign n28970 = ~n28967 & ~n28968;
  assign n28971 = n26781 & n28970;
  assign n28972 = ~n28967 & n28969;
  assign n28973 = ~n28952 & ~n35471;
  assign n28974 = ~n26781 & ~n28970;
  assign n28975 = n25830 & ~n28974;
  assign n28976 = ~n28973 & n28975;
  assign n28977 = ~n27664 & ~n35297;
  assign n28978 = ~n28625 & n28977;
  assign n28979 = n27669 & ~n28978;
  assign n28980 = ~n27669 & n28977;
  assign n28981 = ~n27669 & n28978;
  assign n28982 = ~n28625 & n28980;
  assign n28983 = ~n28979 & ~n35472;
  assign n28984 = ~n28976 & ~n28983;
  assign n28985 = ~n28973 & ~n28974;
  assign n28986 = ~n25830 & ~n28985;
  assign n28987 = n24994 & ~n28986;
  assign n28988 = ~n28984 & ~n28986;
  assign n28989 = n24994 & n28988;
  assign n28990 = ~n28984 & n28987;
  assign n28991 = ~n28939 & ~n35473;
  assign n28992 = ~n24994 & ~n28988;
  assign n28993 = n24076 & ~n28992;
  assign n28994 = ~n28991 & n28993;
  assign n28995 = ~n27692 & ~n35300;
  assign n28996 = ~n28625 & n28995;
  assign n28997 = ~n27702 & ~n28996;
  assign n28998 = ~n27692 & n27702;
  assign n28999 = ~n35300 & n28998;
  assign n29000 = n27702 & n28996;
  assign n29001 = ~n28625 & n28999;
  assign n29002 = n27702 & ~n28996;
  assign n29003 = ~n27702 & n28996;
  assign n29004 = ~n29002 & ~n29003;
  assign n29005 = ~n28997 & ~n35474;
  assign n29006 = ~n28994 & n35475;
  assign n29007 = ~n28991 & ~n28992;
  assign n29008 = ~n24076 & ~n29007;
  assign n29009 = n23269 & ~n29008;
  assign n29010 = ~n29006 & ~n29008;
  assign n29011 = n23269 & n29010;
  assign n29012 = ~n29006 & n29009;
  assign n29013 = ~n28931 & ~n35476;
  assign n29014 = ~n23269 & ~n29010;
  assign n29015 = n22386 & ~n29014;
  assign n29016 = ~n29013 & n29015;
  assign n29017 = ~n27722 & ~n35304;
  assign n29018 = ~n28625 & n29017;
  assign n29019 = ~n35306 & ~n29018;
  assign n29020 = n35306 & n29018;
  assign n29021 = ~n27722 & ~n35306;
  assign n29022 = ~n35304 & n29021;
  assign n29023 = ~n28625 & n29022;
  assign n29024 = n35306 & ~n29018;
  assign n29025 = ~n29023 & ~n29024;
  assign n29026 = ~n29019 & ~n29020;
  assign n29027 = ~n29016 & ~n35477;
  assign n29028 = ~n29013 & ~n29014;
  assign n29029 = ~n22386 & ~n29028;
  assign n29030 = n21612 & ~n29029;
  assign n29031 = ~n29027 & ~n29029;
  assign n29032 = n21612 & n29031;
  assign n29033 = ~n29027 & n29030;
  assign n29034 = ~n28923 & ~n35478;
  assign n29035 = ~n21612 & ~n29031;
  assign n29036 = n20762 & ~n29035;
  assign n29037 = ~n29034 & n29036;
  assign n29038 = ~n27756 & ~n35309;
  assign n29039 = ~n28625 & n29038;
  assign n29040 = ~n35310 & n29039;
  assign n29041 = n35310 & ~n29039;
  assign n29042 = ~n27756 & n35310;
  assign n29043 = ~n35309 & n29042;
  assign n29044 = ~n28625 & n29043;
  assign n29045 = ~n35310 & ~n29039;
  assign n29046 = ~n29044 & ~n29045;
  assign n29047 = ~n29040 & ~n29041;
  assign n29048 = ~n29037 & ~n35479;
  assign n29049 = ~n29034 & ~n29035;
  assign n29050 = ~n20762 & ~n29049;
  assign n29051 = n20011 & ~n29050;
  assign n29052 = ~n29048 & ~n29050;
  assign n29053 = n20011 & n29052;
  assign n29054 = ~n29048 & n29051;
  assign n29055 = ~n28915 & ~n35480;
  assign n29056 = ~n20011 & ~n29052;
  assign n29057 = n19190 & ~n29056;
  assign n29058 = ~n29055 & n29057;
  assign n29059 = ~n27789 & ~n35313;
  assign n29060 = ~n28625 & n29059;
  assign n29061 = ~n35314 & n29060;
  assign n29062 = n35314 & ~n29060;
  assign n29063 = ~n35314 & ~n29060;
  assign n29064 = ~n27789 & n35314;
  assign n29065 = ~n35313 & n29064;
  assign n29066 = n35314 & n29060;
  assign n29067 = ~n28625 & n29065;
  assign n29068 = ~n29063 & ~n35481;
  assign n29069 = ~n29061 & ~n29062;
  assign n29070 = ~n29058 & ~n35482;
  assign n29071 = ~n29055 & ~n29056;
  assign n29072 = ~n19190 & ~n29071;
  assign n29073 = n18472 & ~n29072;
  assign n29074 = ~n29070 & ~n29072;
  assign n29075 = n18472 & n29074;
  assign n29076 = ~n29070 & n29073;
  assign n29077 = ~n28907 & ~n35483;
  assign n29078 = ~n18472 & ~n29074;
  assign n29079 = n17690 & ~n29078;
  assign n29080 = ~n29077 & n29079;
  assign n29081 = ~n27822 & ~n35317;
  assign n29082 = ~n27822 & ~n28625;
  assign n29083 = ~n35317 & n29082;
  assign n29084 = ~n28625 & n29081;
  assign n29085 = n35319 & ~n35484;
  assign n29086 = n27837 & n29082;
  assign n29087 = ~n35319 & n35484;
  assign n29088 = ~n27822 & n35319;
  assign n29089 = ~n35317 & n29088;
  assign n29090 = ~n28625 & n29089;
  assign n29091 = ~n35319 & ~n35484;
  assign n29092 = ~n29090 & ~n29091;
  assign n29093 = ~n29085 & ~n35485;
  assign n29094 = ~n29080 & ~n35486;
  assign n29095 = ~n29077 & ~n29078;
  assign n29096 = ~n17690 & ~n29095;
  assign n29097 = n17001 & ~n29096;
  assign n29098 = ~n29094 & ~n29096;
  assign n29099 = n17001 & n29098;
  assign n29100 = ~n29094 & n29097;
  assign n29101 = ~n28899 & ~n35487;
  assign n29102 = ~n17001 & ~n29098;
  assign n29103 = n16248 & ~n29102;
  assign n29104 = ~n29101 & n29103;
  assign n29105 = ~n28891 & ~n29104;
  assign n29106 = ~n29101 & ~n29102;
  assign n29107 = ~n16248 & ~n29106;
  assign n29108 = n15586 & ~n29107;
  assign n29109 = ~n29105 & ~n29107;
  assign n29110 = n15586 & n29109;
  assign n29111 = ~n29105 & n29108;
  assign n29112 = ~n28883 & ~n35488;
  assign n29113 = ~n15586 & ~n29109;
  assign n29114 = n14866 & ~n29113;
  assign n29115 = ~n29112 & n29114;
  assign n29116 = ~n27892 & ~n35329;
  assign n29117 = ~n27892 & ~n28625;
  assign n29118 = ~n35329 & n29117;
  assign n29119 = ~n28625 & n29116;
  assign n29120 = n27900 & ~n35489;
  assign n29121 = n27904 & n29117;
  assign n29122 = ~n27892 & n27900;
  assign n29123 = ~n35329 & n29122;
  assign n29124 = ~n28625 & n29123;
  assign n29125 = ~n27900 & ~n35489;
  assign n29126 = ~n29124 & ~n29125;
  assign n29127 = ~n29120 & ~n29121;
  assign n29128 = ~n29115 & ~n35490;
  assign n29129 = ~n29112 & ~n29113;
  assign n29130 = ~n14866 & ~n29129;
  assign n29131 = n14233 & ~n29130;
  assign n29132 = ~n29128 & ~n29130;
  assign n29133 = n14233 & n29132;
  assign n29134 = ~n29128 & n29131;
  assign n29135 = ~n28875 & ~n35491;
  assign n29136 = ~n14233 & ~n29132;
  assign n29137 = n13548 & ~n29136;
  assign n29138 = ~n29135 & n29137;
  assign n29139 = ~n28867 & ~n29138;
  assign n29140 = ~n29135 & ~n29136;
  assign n29141 = ~n13548 & ~n29140;
  assign n29142 = n12948 & ~n29141;
  assign n29143 = ~n29139 & ~n29141;
  assign n29144 = n12948 & n29143;
  assign n29145 = ~n29139 & n29142;
  assign n29146 = ~n28859 & ~n35492;
  assign n29147 = ~n12948 & ~n29143;
  assign n29148 = n12296 & ~n29147;
  assign n29149 = ~n29146 & n29148;
  assign n29150 = ~n27958 & ~n35338;
  assign n29151 = ~n27958 & ~n28625;
  assign n29152 = ~n35338 & n29151;
  assign n29153 = ~n28625 & n29150;
  assign n29154 = n27966 & ~n35493;
  assign n29155 = n27970 & n29151;
  assign n29156 = ~n27958 & n27966;
  assign n29157 = ~n35338 & n29156;
  assign n29158 = ~n28625 & n29157;
  assign n29159 = ~n27966 & ~n35493;
  assign n29160 = ~n29158 & ~n29159;
  assign n29161 = ~n29154 & ~n29155;
  assign n29162 = ~n29149 & ~n35494;
  assign n29163 = ~n29146 & ~n29147;
  assign n29164 = ~n12296 & ~n29163;
  assign n29165 = n11719 & ~n29164;
  assign n29166 = ~n29162 & ~n29164;
  assign n29167 = n11719 & n29166;
  assign n29168 = ~n29162 & n29165;
  assign n29169 = ~n28851 & ~n35495;
  assign n29170 = ~n11719 & ~n29166;
  assign n29171 = n11097 & ~n29170;
  assign n29172 = ~n29169 & n29171;
  assign n29173 = ~n28843 & ~n29172;
  assign n29174 = ~n29169 & ~n29170;
  assign n29175 = ~n11097 & ~n29174;
  assign n29176 = n10555 & ~n29175;
  assign n29177 = ~n29173 & ~n29175;
  assign n29178 = n10555 & n29177;
  assign n29179 = ~n29173 & n29176;
  assign n29180 = ~n28835 & ~n35496;
  assign n29181 = ~n10555 & ~n29177;
  assign n29182 = n9969 & ~n29181;
  assign n29183 = ~n29180 & n29182;
  assign n29184 = ~n28024 & ~n35347;
  assign n29185 = ~n28024 & ~n28625;
  assign n29186 = ~n35347 & n29185;
  assign n29187 = ~n28625 & n29184;
  assign n29188 = n28032 & ~n35497;
  assign n29189 = n28036 & n29185;
  assign n29190 = ~n28024 & n28032;
  assign n29191 = ~n35347 & n29190;
  assign n29192 = ~n28625 & n29191;
  assign n29193 = ~n28032 & ~n35497;
  assign n29194 = ~n29192 & ~n29193;
  assign n29195 = ~n29188 & ~n29189;
  assign n29196 = ~n29183 & ~n35498;
  assign n29197 = ~n29180 & ~n29181;
  assign n29198 = ~n9969 & ~n29197;
  assign n29199 = n9457 & ~n29198;
  assign n29200 = ~n29196 & ~n29198;
  assign n29201 = n9457 & n29200;
  assign n29202 = ~n29196 & n29199;
  assign n29203 = ~n28827 & ~n35499;
  assign n29204 = ~n9457 & ~n29200;
  assign n29205 = n8896 & ~n29204;
  assign n29206 = ~n29203 & n29205;
  assign n29207 = ~n28819 & ~n29206;
  assign n29208 = ~n29203 & ~n29204;
  assign n29209 = ~n8896 & ~n29208;
  assign n29210 = n8411 & ~n29209;
  assign n29211 = ~n29207 & ~n29209;
  assign n29212 = n8411 & n29211;
  assign n29213 = ~n29207 & n29210;
  assign n29214 = ~n28811 & ~n35500;
  assign n29215 = ~n8411 & ~n29211;
  assign n29216 = n7885 & ~n29215;
  assign n29217 = ~n29214 & n29216;
  assign n29218 = ~n28090 & ~n35356;
  assign n29219 = ~n28090 & ~n28625;
  assign n29220 = ~n35356 & n29219;
  assign n29221 = ~n28625 & n29218;
  assign n29222 = n28098 & ~n35501;
  assign n29223 = n28102 & n29219;
  assign n29224 = ~n28090 & n28098;
  assign n29225 = ~n35356 & n29224;
  assign n29226 = ~n28625 & n29225;
  assign n29227 = ~n28098 & ~n35501;
  assign n29228 = ~n29226 & ~n29227;
  assign n29229 = ~n29222 & ~n29223;
  assign n29230 = ~n29217 & ~n35502;
  assign n29231 = ~n29214 & ~n29215;
  assign n29232 = ~n7885 & ~n29231;
  assign n29233 = n7428 & ~n29232;
  assign n29234 = ~n29230 & ~n29232;
  assign n29235 = n7428 & n29234;
  assign n29236 = ~n29230 & n29233;
  assign n29237 = ~n28803 & ~n35503;
  assign n29238 = ~n7428 & ~n29234;
  assign n29239 = n6937 & ~n29238;
  assign n29240 = ~n29237 & n29239;
  assign n29241 = ~n28795 & ~n29240;
  assign n29242 = ~n29237 & ~n29238;
  assign n29243 = ~n6937 & ~n29242;
  assign n29244 = n6507 & ~n29243;
  assign n29245 = ~n29241 & ~n29243;
  assign n29246 = n6507 & n29245;
  assign n29247 = ~n29241 & n29244;
  assign n29248 = ~n28787 & ~n35504;
  assign n29249 = ~n6507 & ~n29245;
  assign n29250 = n6051 & ~n29249;
  assign n29251 = ~n29248 & n29250;
  assign n29252 = ~n28156 & ~n35365;
  assign n29253 = ~n28156 & ~n28625;
  assign n29254 = ~n35365 & n29253;
  assign n29255 = ~n28625 & n29252;
  assign n29256 = n28164 & ~n35505;
  assign n29257 = n28168 & n29253;
  assign n29258 = ~n28156 & n28164;
  assign n29259 = ~n35365 & n29258;
  assign n29260 = ~n28625 & n29259;
  assign n29261 = ~n28164 & ~n35505;
  assign n29262 = ~n29260 & ~n29261;
  assign n29263 = ~n29256 & ~n29257;
  assign n29264 = ~n29251 & ~n35506;
  assign n29265 = ~n29248 & ~n29249;
  assign n29266 = ~n6051 & ~n29265;
  assign n29267 = n5648 & ~n29266;
  assign n29268 = ~n29264 & ~n29266;
  assign n29269 = n5648 & n29268;
  assign n29270 = ~n29264 & n29267;
  assign n29271 = ~n28779 & ~n35507;
  assign n29272 = ~n5648 & ~n29268;
  assign n29273 = n5223 & ~n29272;
  assign n29274 = ~n29271 & n29273;
  assign n29275 = ~n28771 & ~n29274;
  assign n29276 = ~n29271 & ~n29272;
  assign n29277 = ~n5223 & ~n29276;
  assign n29278 = n4851 & ~n29277;
  assign n29279 = ~n29275 & ~n29277;
  assign n29280 = n4851 & n29279;
  assign n29281 = ~n29275 & n29278;
  assign n29282 = ~n28763 & ~n35508;
  assign n29283 = ~n4851 & ~n29279;
  assign n29284 = n4461 & ~n29283;
  assign n29285 = ~n29282 & n29284;
  assign n29286 = ~n28222 & ~n35374;
  assign n29287 = ~n28222 & ~n28625;
  assign n29288 = ~n35374 & n29287;
  assign n29289 = ~n28625 & n29286;
  assign n29290 = n28230 & ~n35509;
  assign n29291 = n28234 & n29287;
  assign n29292 = ~n28222 & n28230;
  assign n29293 = ~n35374 & n29292;
  assign n29294 = ~n28625 & n29293;
  assign n29295 = ~n28230 & ~n35509;
  assign n29296 = ~n29294 & ~n29295;
  assign n29297 = ~n29290 & ~n29291;
  assign n29298 = ~n29285 & ~n35510;
  assign n29299 = ~n29282 & ~n29283;
  assign n29300 = ~n4461 & ~n29299;
  assign n29301 = n4115 & ~n29300;
  assign n29302 = ~n29298 & ~n29300;
  assign n29303 = n4115 & n29302;
  assign n29304 = ~n29298 & n29301;
  assign n29305 = ~n28755 & ~n35511;
  assign n29306 = ~n4115 & ~n29302;
  assign n29307 = n3754 & ~n29306;
  assign n29308 = ~n29305 & n29307;
  assign n29309 = ~n28747 & ~n29308;
  assign n29310 = ~n29305 & ~n29306;
  assign n29311 = ~n3754 & ~n29310;
  assign n29312 = n3444 & ~n29311;
  assign n29313 = ~n29309 & ~n29311;
  assign n29314 = n3444 & n29313;
  assign n29315 = ~n29309 & n29312;
  assign n29316 = ~n28739 & ~n35512;
  assign n29317 = ~n3444 & ~n29313;
  assign n29318 = n3116 & ~n29317;
  assign n29319 = ~n29316 & n29318;
  assign n29320 = ~n28288 & ~n35383;
  assign n29321 = ~n28288 & ~n28625;
  assign n29322 = ~n35383 & n29321;
  assign n29323 = ~n28625 & n29320;
  assign n29324 = n28296 & ~n35513;
  assign n29325 = n28300 & n29321;
  assign n29326 = ~n28288 & n28296;
  assign n29327 = ~n35383 & n29326;
  assign n29328 = ~n28625 & n29327;
  assign n29329 = ~n28296 & ~n35513;
  assign n29330 = ~n29328 & ~n29329;
  assign n29331 = ~n29324 & ~n29325;
  assign n29332 = ~n29319 & ~n35514;
  assign n29333 = ~n29316 & ~n29317;
  assign n29334 = ~n3116 & ~n29333;
  assign n29335 = n2833 & ~n29334;
  assign n29336 = ~n29332 & ~n29334;
  assign n29337 = n2833 & n29336;
  assign n29338 = ~n29332 & n29335;
  assign n29339 = ~n28731 & ~n35515;
  assign n29340 = ~n2833 & ~n29336;
  assign n29341 = n2536 & ~n29340;
  assign n29342 = ~n29339 & n29341;
  assign n29343 = ~n28723 & ~n29342;
  assign n29344 = ~n29339 & ~n29340;
  assign n29345 = ~n2536 & ~n29344;
  assign n29346 = n2283 & ~n29345;
  assign n29347 = ~n29343 & ~n29345;
  assign n29348 = n2283 & n29347;
  assign n29349 = ~n29343 & n29346;
  assign n29350 = ~n28715 & ~n35516;
  assign n29351 = ~n2283 & ~n29347;
  assign n29352 = n2021 & ~n29351;
  assign n29353 = ~n29350 & n29352;
  assign n29354 = ~n28354 & ~n35392;
  assign n29355 = ~n28354 & ~n28625;
  assign n29356 = ~n35392 & n29355;
  assign n29357 = ~n28625 & n29354;
  assign n29358 = n28362 & ~n35517;
  assign n29359 = n28366 & n29355;
  assign n29360 = ~n28354 & n28362;
  assign n29361 = ~n35392 & n29360;
  assign n29362 = ~n28625 & n29361;
  assign n29363 = ~n28362 & ~n35517;
  assign n29364 = ~n29362 & ~n29363;
  assign n29365 = ~n29358 & ~n29359;
  assign n29366 = ~n29353 & ~n35518;
  assign n29367 = ~n29350 & ~n29351;
  assign n29368 = ~n2021 & ~n29367;
  assign n29369 = n1796 & ~n29368;
  assign n29370 = ~n29366 & ~n29368;
  assign n29371 = n1796 & n29370;
  assign n29372 = ~n29366 & n29369;
  assign n29373 = ~n28707 & ~n35519;
  assign n29374 = ~n1796 & ~n29370;
  assign n29375 = n1567 & ~n29374;
  assign n29376 = ~n29373 & n29375;
  assign n29377 = ~n28699 & ~n29376;
  assign n29378 = ~n29373 & ~n29374;
  assign n29379 = ~n1567 & ~n29378;
  assign n29380 = n1374 & ~n29379;
  assign n29381 = ~n29377 & ~n29379;
  assign n29382 = n1374 & n29381;
  assign n29383 = ~n29377 & n29380;
  assign n29384 = ~n28691 & ~n35520;
  assign n29385 = ~n1374 & ~n29381;
  assign n29386 = n1179 & ~n29385;
  assign n29387 = ~n29384 & n29386;
  assign n29388 = ~n28420 & ~n35401;
  assign n29389 = ~n28420 & ~n28625;
  assign n29390 = ~n35401 & n29389;
  assign n29391 = ~n28625 & n29388;
  assign n29392 = n28428 & ~n35521;
  assign n29393 = n28432 & n29389;
  assign n29394 = ~n28420 & n28428;
  assign n29395 = ~n35401 & n29394;
  assign n29396 = ~n28625 & n29395;
  assign n29397 = ~n28428 & ~n35521;
  assign n29398 = ~n29396 & ~n29397;
  assign n29399 = ~n29392 & ~n29393;
  assign n29400 = ~n29387 & ~n35522;
  assign n29401 = ~n29384 & ~n29385;
  assign n29402 = ~n1179 & ~n29401;
  assign n29403 = n1016 & ~n29402;
  assign n29404 = ~n29400 & ~n29402;
  assign n29405 = n1016 & n29404;
  assign n29406 = ~n29400 & n29403;
  assign n29407 = ~n28683 & ~n35523;
  assign n29408 = ~n1016 & ~n29404;
  assign n29409 = n855 & ~n29408;
  assign n29410 = ~n29407 & n29409;
  assign n29411 = ~n28675 & ~n29410;
  assign n29412 = ~n29407 & ~n29408;
  assign n29413 = ~n855 & ~n29412;
  assign n29414 = n720 & ~n29413;
  assign n29415 = ~n29411 & ~n29413;
  assign n29416 = n720 & n29415;
  assign n29417 = ~n29411 & n29414;
  assign n29418 = ~n28667 & ~n35524;
  assign n29419 = ~n720 & ~n29415;
  assign n29420 = n592 & ~n29419;
  assign n29421 = ~n29418 & n29420;
  assign n29422 = ~n28486 & ~n35410;
  assign n29423 = ~n28486 & ~n28625;
  assign n29424 = ~n35410 & n29423;
  assign n29425 = ~n28625 & n29422;
  assign n29426 = n28494 & ~n35525;
  assign n29427 = n28498 & n29423;
  assign n29428 = ~n28486 & n28494;
  assign n29429 = ~n35410 & n29428;
  assign n29430 = ~n28625 & n29429;
  assign n29431 = ~n28494 & ~n35525;
  assign n29432 = ~n29430 & ~n29431;
  assign n29433 = ~n29426 & ~n29427;
  assign n29434 = ~n29421 & ~n35526;
  assign n29435 = ~n29418 & ~n29419;
  assign n29436 = ~n592 & ~n29435;
  assign n29437 = n487 & ~n29436;
  assign n29438 = ~n29434 & ~n29436;
  assign n29439 = n487 & n29438;
  assign n29440 = ~n29434 & n29437;
  assign n29441 = ~n28659 & ~n35527;
  assign n29442 = ~n487 & ~n29438;
  assign n29443 = n393 & ~n29442;
  assign n29444 = ~n29441 & n29443;
  assign n29445 = ~n28651 & ~n29444;
  assign n29446 = ~n29441 & ~n29442;
  assign n29447 = ~n393 & ~n29446;
  assign n29448 = n321 & ~n29447;
  assign n29449 = ~n29445 & ~n29447;
  assign n29450 = n321 & n29449;
  assign n29451 = ~n29445 & n29448;
  assign n29452 = ~n28643 & ~n35528;
  assign n29453 = ~n321 & ~n29449;
  assign n29454 = ~n29452 & ~n29453;
  assign n29455 = ~n263 & ~n29454;
  assign n29456 = n263 & ~n29453;
  assign n29457 = ~n29452 & n29456;
  assign n29458 = ~n35427 & ~n29457;
  assign n29459 = ~n29455 & ~n29458;
  assign n29460 = ~n214 & ~n29459;
  assign n29461 = ~n28554 & ~n28556;
  assign n29462 = ~n28625 & n29461;
  assign n29463 = ~n35419 & ~n29462;
  assign n29464 = ~n28556 & n35419;
  assign n29465 = ~n28554 & n29464;
  assign n29466 = n35419 & n29462;
  assign n29467 = ~n28625 & n29465;
  assign n29468 = ~n29463 & ~n35529;
  assign n29469 = n214 & ~n29455;
  assign n29470 = n214 & n29459;
  assign n29471 = ~n29458 & n29469;
  assign n29472 = ~n29468 & ~n35530;
  assign n29473 = ~n29460 & ~n29472;
  assign n29474 = ~n197 & ~n29473;
  assign n29475 = n197 & ~n29460;
  assign n29476 = ~n29472 & n29475;
  assign n29477 = ~n28571 & ~n35421;
  assign n29478 = ~n28571 & ~n28625;
  assign n29479 = ~n35421 & n29478;
  assign n29480 = ~n28625 & n29477;
  assign n29481 = n28579 & ~n35531;
  assign n29482 = n28583 & n29478;
  assign n29483 = ~n28571 & n28579;
  assign n29484 = ~n35421 & n29483;
  assign n29485 = ~n28625 & n29484;
  assign n29486 = ~n28579 & ~n35531;
  assign n29487 = ~n29485 & ~n29486;
  assign n29488 = ~n29481 & ~n29482;
  assign n29489 = ~n29476 & ~n35532;
  assign n29490 = ~n29474 & ~n29489;
  assign n29491 = ~n28585 & ~n28587;
  assign n29492 = ~n28625 & n29491;
  assign n29493 = ~n35423 & ~n29492;
  assign n29494 = ~n28587 & n35423;
  assign n29495 = ~n28585 & n29494;
  assign n29496 = n35423 & n29492;
  assign n29497 = ~n28625 & n29495;
  assign n29498 = ~n29493 & ~n35533;
  assign n29499 = ~n28601 & ~n28609;
  assign n29500 = ~n28609 & ~n28625;
  assign n29501 = ~n28601 & n29500;
  assign n29502 = ~n28625 & n29499;
  assign n29503 = ~n35426 & ~n35534;
  assign n29504 = ~n29498 & n29503;
  assign n29505 = ~n29490 & n29504;
  assign n29506 = n193 & ~n29505;
  assign n29507 = ~n29474 & n29498;
  assign n29508 = n29490 & n29498;
  assign n29509 = ~n29489 & n29507;
  assign n29510 = n28601 & ~n29500;
  assign n29511 = ~n193 & ~n29499;
  assign n29512 = ~n29510 & n29511;
  assign n29513 = ~n35535 & ~n29512;
  assign n29514 = ~n29506 & n29513;
  assign n29515 = ~n29455 & ~n29457;
  assign n29516 = ~n29514 & n29515;
  assign n29517 = ~n35427 & n29516;
  assign n29518 = n35427 & ~n29516;
  assign n29519 = n35427 & ~n29455;
  assign n29520 = ~n29457 & n29519;
  assign n29521 = ~n29514 & n29520;
  assign n29522 = ~n35427 & ~n29516;
  assign n29523 = ~n29521 & ~n29522;
  assign n29524 = ~n29517 & ~n29518;
  assign n29525 = pi4  & ~n29514;
  assign n29526 = ~pi2  & ~pi3 ;
  assign n29527 = ~pi4  & n29526;
  assign n29528 = ~pi4  & ~n29526;
  assign n29529 = pi4  & n29514;
  assign n29530 = ~n29528 & ~n29529;
  assign n29531 = ~n29525 & ~n29527;
  assign n29532 = ~n28625 & n35537;
  assign n29533 = ~pi4  & ~n29514;
  assign n29534 = pi5  & ~n29533;
  assign n29535 = ~pi5  & n29533;
  assign n29536 = n28954 & ~n29514;
  assign n29537 = ~n29534 & ~n35538;
  assign n29538 = ~n28623 & ~n29527;
  assign n29539 = ~n35426 & n29538;
  assign n29540 = ~n28617 & n29539;
  assign n29541 = n28625 & ~n35537;
  assign n29542 = ~n29525 & n29540;
  assign n29543 = n29537 & ~n35539;
  assign n29544 = ~n29532 & ~n29543;
  assign n29545 = ~n27648 & ~n29544;
  assign n29546 = n27648 & ~n29532;
  assign n29547 = ~n29543 & n29546;
  assign n29548 = ~n28625 & ~n29512;
  assign n29549 = ~n35535 & n29548;
  assign n29550 = ~n28625 & n29514;
  assign n29551 = ~n29506 & n29549;
  assign n29552 = ~n35538 & ~n35540;
  assign n29553 = pi6  & ~n29552;
  assign n29554 = ~pi6  & ~n35540;
  assign n29555 = ~pi6  & n29552;
  assign n29556 = ~n35538 & n29554;
  assign n29557 = ~n29553 & ~n35541;
  assign n29558 = ~n29547 & ~n29557;
  assign n29559 = ~n29545 & ~n29558;
  assign n29560 = ~n26781 & ~n29559;
  assign n29561 = n26781 & ~n29545;
  assign n29562 = ~n29558 & n29561;
  assign n29563 = n26781 & n29559;
  assign n29564 = ~n35470 & ~n28968;
  assign n29565 = ~n29514 & n29564;
  assign n29566 = n28966 & ~n29565;
  assign n29567 = ~n28966 & n29564;
  assign n29568 = ~n28966 & n29565;
  assign n29569 = ~n29514 & n29567;
  assign n29570 = ~n29566 & ~n35543;
  assign n29571 = ~n35542 & ~n29570;
  assign n29572 = ~n29560 & ~n29571;
  assign n29573 = ~n25830 & ~n29572;
  assign n29574 = n25830 & ~n29560;
  assign n29575 = ~n29571 & n29574;
  assign n29576 = ~n35471 & ~n28974;
  assign n29577 = ~n28974 & ~n29514;
  assign n29578 = ~n35471 & n29577;
  assign n29579 = ~n29514 & n29576;
  assign n29580 = n28952 & ~n35544;
  assign n29581 = n28973 & n29577;
  assign n29582 = n28952 & ~n35471;
  assign n29583 = ~n28974 & n29582;
  assign n29584 = ~n29514 & n29583;
  assign n29585 = ~n28952 & ~n35544;
  assign n29586 = ~n29584 & ~n29585;
  assign n29587 = ~n29580 & ~n29581;
  assign n29588 = ~n29575 & ~n35545;
  assign n29589 = ~n29573 & ~n29588;
  assign n29590 = ~n24994 & ~n29589;
  assign n29591 = n24994 & ~n29573;
  assign n29592 = ~n29588 & n29591;
  assign n29593 = n24994 & n29589;
  assign n29594 = ~n28976 & ~n28986;
  assign n29595 = ~n29514 & n29594;
  assign n29596 = ~n28983 & ~n29595;
  assign n29597 = n28983 & ~n28986;
  assign n29598 = ~n28976 & n29597;
  assign n29599 = n28983 & n29595;
  assign n29600 = ~n29514 & n29598;
  assign n29601 = n28983 & ~n29595;
  assign n29602 = ~n28983 & n29595;
  assign n29603 = ~n29601 & ~n29602;
  assign n29604 = ~n29596 & ~n35547;
  assign n29605 = ~n35546 & n35548;
  assign n29606 = ~n29590 & ~n29605;
  assign n29607 = ~n24076 & ~n29606;
  assign n29608 = n24076 & ~n29590;
  assign n29609 = ~n29605 & n29608;
  assign n29610 = ~n35473 & ~n28992;
  assign n29611 = ~n28992 & ~n29514;
  assign n29612 = ~n35473 & n29611;
  assign n29613 = ~n29514 & n29610;
  assign n29614 = n28939 & ~n35549;
  assign n29615 = n28991 & n29611;
  assign n29616 = n28939 & ~n35473;
  assign n29617 = ~n28992 & n29616;
  assign n29618 = ~n29514 & n29617;
  assign n29619 = ~n28939 & ~n35549;
  assign n29620 = ~n29618 & ~n29619;
  assign n29621 = ~n29614 & ~n29615;
  assign n29622 = ~n29609 & ~n35550;
  assign n29623 = ~n29607 & ~n29622;
  assign n29624 = ~n23269 & ~n29623;
  assign n29625 = n23269 & ~n29607;
  assign n29626 = ~n29622 & n29625;
  assign n29627 = n23269 & n29623;
  assign n29628 = ~n28994 & ~n29008;
  assign n29629 = ~n29514 & n29628;
  assign n29630 = ~n35475 & ~n29629;
  assign n29631 = n35475 & n29629;
  assign n29632 = ~n35475 & ~n29008;
  assign n29633 = ~n28994 & n29632;
  assign n29634 = ~n29514 & n29633;
  assign n29635 = n35475 & ~n29629;
  assign n29636 = ~n29634 & ~n29635;
  assign n29637 = ~n29630 & ~n29631;
  assign n29638 = ~n35551 & ~n35552;
  assign n29639 = ~n29624 & ~n29638;
  assign n29640 = ~n22386 & ~n29639;
  assign n29641 = n22386 & ~n29624;
  assign n29642 = ~n29638 & n29641;
  assign n29643 = ~n35476 & ~n29014;
  assign n29644 = ~n29014 & ~n29514;
  assign n29645 = ~n35476 & n29644;
  assign n29646 = ~n29514 & n29643;
  assign n29647 = n28931 & ~n35553;
  assign n29648 = n29013 & n29644;
  assign n29649 = n28931 & ~n35476;
  assign n29650 = ~n29014 & n29649;
  assign n29651 = ~n29514 & n29650;
  assign n29652 = ~n28931 & ~n35553;
  assign n29653 = ~n29651 & ~n29652;
  assign n29654 = ~n29647 & ~n29648;
  assign n29655 = ~n29642 & ~n35554;
  assign n29656 = ~n29640 & ~n29655;
  assign n29657 = ~n21612 & ~n29656;
  assign n29658 = n21612 & ~n29640;
  assign n29659 = ~n29655 & n29658;
  assign n29660 = n21612 & n29656;
  assign n29661 = ~n29016 & ~n29029;
  assign n29662 = ~n29514 & n29661;
  assign n29663 = ~n35477 & n29662;
  assign n29664 = n35477 & ~n29662;
  assign n29665 = n35477 & ~n29029;
  assign n29666 = ~n29016 & n29665;
  assign n29667 = ~n29514 & n29666;
  assign n29668 = ~n35477 & ~n29662;
  assign n29669 = ~n29667 & ~n29668;
  assign n29670 = ~n29663 & ~n29664;
  assign n29671 = ~n35555 & ~n35556;
  assign n29672 = ~n29657 & ~n29671;
  assign n29673 = ~n20762 & ~n29672;
  assign n29674 = n20762 & ~n29657;
  assign n29675 = ~n29671 & n29674;
  assign n29676 = ~n35478 & ~n29035;
  assign n29677 = ~n29035 & ~n29514;
  assign n29678 = ~n35478 & n29677;
  assign n29679 = ~n29514 & n29676;
  assign n29680 = n28923 & ~n35557;
  assign n29681 = n29034 & n29677;
  assign n29682 = n28923 & ~n35478;
  assign n29683 = ~n29035 & n29682;
  assign n29684 = ~n29514 & n29683;
  assign n29685 = ~n28923 & ~n35557;
  assign n29686 = ~n29684 & ~n29685;
  assign n29687 = ~n29680 & ~n29681;
  assign n29688 = ~n29675 & ~n35558;
  assign n29689 = ~n29673 & ~n29688;
  assign n29690 = ~n20011 & ~n29689;
  assign n29691 = n20011 & ~n29673;
  assign n29692 = ~n29688 & n29691;
  assign n29693 = n20011 & n29689;
  assign n29694 = ~n29037 & ~n29050;
  assign n29695 = ~n29514 & n29694;
  assign n29696 = ~n35479 & n29695;
  assign n29697 = n35479 & ~n29695;
  assign n29698 = ~n35479 & ~n29695;
  assign n29699 = n35479 & ~n29050;
  assign n29700 = ~n29037 & n29699;
  assign n29701 = n35479 & n29695;
  assign n29702 = ~n29514 & n29700;
  assign n29703 = ~n29698 & ~n35560;
  assign n29704 = ~n29696 & ~n29697;
  assign n29705 = ~n35559 & ~n35561;
  assign n29706 = ~n29690 & ~n29705;
  assign n29707 = ~n19190 & ~n29706;
  assign n29708 = n19190 & ~n29690;
  assign n29709 = ~n29705 & n29708;
  assign n29710 = ~n35480 & ~n29056;
  assign n29711 = ~n29056 & ~n29514;
  assign n29712 = ~n35480 & n29711;
  assign n29713 = ~n29514 & n29710;
  assign n29714 = n28915 & ~n35562;
  assign n29715 = n29055 & n29711;
  assign n29716 = n28915 & ~n35480;
  assign n29717 = ~n29056 & n29716;
  assign n29718 = ~n29514 & n29717;
  assign n29719 = ~n28915 & ~n35562;
  assign n29720 = ~n29718 & ~n29719;
  assign n29721 = ~n29714 & ~n29715;
  assign n29722 = ~n29709 & ~n35563;
  assign n29723 = ~n29707 & ~n29722;
  assign n29724 = ~n18472 & ~n29723;
  assign n29725 = n18472 & ~n29707;
  assign n29726 = ~n29722 & n29725;
  assign n29727 = n18472 & n29723;
  assign n29728 = ~n29058 & ~n29072;
  assign n29729 = ~n29072 & ~n29514;
  assign n29730 = ~n29058 & n29729;
  assign n29731 = ~n29514 & n29728;
  assign n29732 = n35482 & ~n35565;
  assign n29733 = n29070 & n29729;
  assign n29734 = ~n35482 & n35565;
  assign n29735 = n35482 & ~n29072;
  assign n29736 = ~n29058 & n29735;
  assign n29737 = ~n29514 & n29736;
  assign n29738 = ~n35482 & ~n35565;
  assign n29739 = ~n29737 & ~n29738;
  assign n29740 = ~n29732 & ~n35566;
  assign n29741 = ~n35564 & ~n35567;
  assign n29742 = ~n29724 & ~n29741;
  assign n29743 = ~n17690 & ~n29742;
  assign n29744 = n17690 & ~n29724;
  assign n29745 = ~n29741 & n29744;
  assign n29746 = ~n35483 & ~n29078;
  assign n29747 = ~n29078 & ~n29514;
  assign n29748 = ~n35483 & n29747;
  assign n29749 = ~n29514 & n29746;
  assign n29750 = n28907 & ~n35568;
  assign n29751 = n29077 & n29747;
  assign n29752 = n28907 & ~n35483;
  assign n29753 = ~n29078 & n29752;
  assign n29754 = ~n29514 & n29753;
  assign n29755 = ~n28907 & ~n35568;
  assign n29756 = ~n29754 & ~n29755;
  assign n29757 = ~n29750 & ~n29751;
  assign n29758 = ~n29745 & ~n35569;
  assign n29759 = ~n29743 & ~n29758;
  assign n29760 = ~n17001 & ~n29759;
  assign n29761 = ~n29080 & ~n29096;
  assign n29762 = ~n29514 & n29761;
  assign n29763 = ~n35486 & ~n29762;
  assign n29764 = n35486 & ~n29096;
  assign n29765 = ~n29080 & n29764;
  assign n29766 = n35486 & n29762;
  assign n29767 = ~n29514 & n29765;
  assign n29768 = ~n29763 & ~n35570;
  assign n29769 = n17001 & ~n29743;
  assign n29770 = ~n29758 & n29769;
  assign n29771 = n17001 & n29759;
  assign n29772 = ~n29768 & ~n35571;
  assign n29773 = ~n29760 & ~n29772;
  assign n29774 = ~n16248 & ~n29773;
  assign n29775 = n16248 & ~n29760;
  assign n29776 = ~n29772 & n29775;
  assign n29777 = ~n35487 & ~n29102;
  assign n29778 = ~n29102 & ~n29514;
  assign n29779 = ~n35487 & n29778;
  assign n29780 = ~n29514 & n29777;
  assign n29781 = n28899 & ~n35572;
  assign n29782 = n29101 & n29778;
  assign n29783 = n28899 & ~n35487;
  assign n29784 = ~n29102 & n29783;
  assign n29785 = ~n29514 & n29784;
  assign n29786 = ~n28899 & ~n35572;
  assign n29787 = ~n29785 & ~n29786;
  assign n29788 = ~n29781 & ~n29782;
  assign n29789 = ~n29776 & ~n35573;
  assign n29790 = ~n29774 & ~n29789;
  assign n29791 = ~n15586 & ~n29790;
  assign n29792 = n15586 & ~n29774;
  assign n29793 = ~n29789 & n29792;
  assign n29794 = n15586 & n29790;
  assign n29795 = ~n29104 & ~n29107;
  assign n29796 = ~n29107 & ~n29514;
  assign n29797 = ~n29104 & n29796;
  assign n29798 = ~n29514 & n29795;
  assign n29799 = n28891 & ~n35575;
  assign n29800 = n29105 & n29796;
  assign n29801 = n28891 & ~n29107;
  assign n29802 = ~n29104 & n29801;
  assign n29803 = ~n29514 & n29802;
  assign n29804 = ~n28891 & ~n35575;
  assign n29805 = ~n29803 & ~n29804;
  assign n29806 = ~n29799 & ~n29800;
  assign n29807 = ~n35574 & ~n35576;
  assign n29808 = ~n29791 & ~n29807;
  assign n29809 = ~n14866 & ~n29808;
  assign n29810 = n14866 & ~n29791;
  assign n29811 = ~n29807 & n29810;
  assign n29812 = ~n35488 & ~n29113;
  assign n29813 = ~n29113 & ~n29514;
  assign n29814 = ~n35488 & n29813;
  assign n29815 = ~n29514 & n29812;
  assign n29816 = n28883 & ~n35577;
  assign n29817 = n29112 & n29813;
  assign n29818 = n28883 & ~n35488;
  assign n29819 = ~n29113 & n29818;
  assign n29820 = ~n29514 & n29819;
  assign n29821 = ~n28883 & ~n35577;
  assign n29822 = ~n29820 & ~n29821;
  assign n29823 = ~n29816 & ~n29817;
  assign n29824 = ~n29811 & ~n35578;
  assign n29825 = ~n29809 & ~n29824;
  assign n29826 = ~n14233 & ~n29825;
  assign n29827 = ~n29115 & ~n29130;
  assign n29828 = ~n29514 & n29827;
  assign n29829 = ~n35490 & ~n29828;
  assign n29830 = n35490 & ~n29130;
  assign n29831 = ~n29115 & n29830;
  assign n29832 = n35490 & n29828;
  assign n29833 = ~n29514 & n29831;
  assign n29834 = ~n29829 & ~n35579;
  assign n29835 = n14233 & ~n29809;
  assign n29836 = ~n29824 & n29835;
  assign n29837 = n14233 & n29825;
  assign n29838 = ~n29834 & ~n35580;
  assign n29839 = ~n29826 & ~n29838;
  assign n29840 = ~n13548 & ~n29839;
  assign n29841 = n13548 & ~n29826;
  assign n29842 = ~n29838 & n29841;
  assign n29843 = ~n35491 & ~n29136;
  assign n29844 = ~n29136 & ~n29514;
  assign n29845 = ~n35491 & n29844;
  assign n29846 = ~n29514 & n29843;
  assign n29847 = n28875 & ~n35581;
  assign n29848 = n29135 & n29844;
  assign n29849 = n28875 & ~n35491;
  assign n29850 = ~n29136 & n29849;
  assign n29851 = ~n29514 & n29850;
  assign n29852 = ~n28875 & ~n35581;
  assign n29853 = ~n29851 & ~n29852;
  assign n29854 = ~n29847 & ~n29848;
  assign n29855 = ~n29842 & ~n35582;
  assign n29856 = ~n29840 & ~n29855;
  assign n29857 = ~n12948 & ~n29856;
  assign n29858 = n12948 & ~n29840;
  assign n29859 = ~n29855 & n29858;
  assign n29860 = n12948 & n29856;
  assign n29861 = ~n29138 & ~n29141;
  assign n29862 = ~n29141 & ~n29514;
  assign n29863 = ~n29138 & n29862;
  assign n29864 = ~n29514 & n29861;
  assign n29865 = n28867 & ~n35584;
  assign n29866 = n29139 & n29862;
  assign n29867 = n28867 & ~n29141;
  assign n29868 = ~n29138 & n29867;
  assign n29869 = ~n29514 & n29868;
  assign n29870 = ~n28867 & ~n35584;
  assign n29871 = ~n29869 & ~n29870;
  assign n29872 = ~n29865 & ~n29866;
  assign n29873 = ~n35583 & ~n35585;
  assign n29874 = ~n29857 & ~n29873;
  assign n29875 = ~n12296 & ~n29874;
  assign n29876 = n12296 & ~n29857;
  assign n29877 = ~n29873 & n29876;
  assign n29878 = ~n35492 & ~n29147;
  assign n29879 = ~n29147 & ~n29514;
  assign n29880 = ~n35492 & n29879;
  assign n29881 = ~n29514 & n29878;
  assign n29882 = n28859 & ~n35586;
  assign n29883 = n29146 & n29879;
  assign n29884 = n28859 & ~n35492;
  assign n29885 = ~n29147 & n29884;
  assign n29886 = ~n29514 & n29885;
  assign n29887 = ~n28859 & ~n35586;
  assign n29888 = ~n29886 & ~n29887;
  assign n29889 = ~n29882 & ~n29883;
  assign n29890 = ~n29877 & ~n35587;
  assign n29891 = ~n29875 & ~n29890;
  assign n29892 = ~n11719 & ~n29891;
  assign n29893 = ~n29149 & ~n29164;
  assign n29894 = ~n29514 & n29893;
  assign n29895 = ~n35494 & ~n29894;
  assign n29896 = n35494 & ~n29164;
  assign n29897 = ~n29149 & n29896;
  assign n29898 = n35494 & n29894;
  assign n29899 = ~n29514 & n29897;
  assign n29900 = ~n29895 & ~n35588;
  assign n29901 = n11719 & ~n29875;
  assign n29902 = ~n29890 & n29901;
  assign n29903 = n11719 & n29891;
  assign n29904 = ~n29900 & ~n35589;
  assign n29905 = ~n29892 & ~n29904;
  assign n29906 = ~n11097 & ~n29905;
  assign n29907 = n11097 & ~n29892;
  assign n29908 = ~n29904 & n29907;
  assign n29909 = ~n35495 & ~n29170;
  assign n29910 = ~n29170 & ~n29514;
  assign n29911 = ~n35495 & n29910;
  assign n29912 = ~n29514 & n29909;
  assign n29913 = n28851 & ~n35590;
  assign n29914 = n29169 & n29910;
  assign n29915 = n28851 & ~n35495;
  assign n29916 = ~n29170 & n29915;
  assign n29917 = ~n29514 & n29916;
  assign n29918 = ~n28851 & ~n35590;
  assign n29919 = ~n29917 & ~n29918;
  assign n29920 = ~n29913 & ~n29914;
  assign n29921 = ~n29908 & ~n35591;
  assign n29922 = ~n29906 & ~n29921;
  assign n29923 = ~n10555 & ~n29922;
  assign n29924 = n10555 & ~n29906;
  assign n29925 = ~n29921 & n29924;
  assign n29926 = n10555 & n29922;
  assign n29927 = ~n29172 & ~n29175;
  assign n29928 = ~n29175 & ~n29514;
  assign n29929 = ~n29172 & n29928;
  assign n29930 = ~n29514 & n29927;
  assign n29931 = n28843 & ~n35593;
  assign n29932 = n29173 & n29928;
  assign n29933 = n28843 & ~n29175;
  assign n29934 = ~n29172 & n29933;
  assign n29935 = ~n29514 & n29934;
  assign n29936 = ~n28843 & ~n35593;
  assign n29937 = ~n29935 & ~n29936;
  assign n29938 = ~n29931 & ~n29932;
  assign n29939 = ~n35592 & ~n35594;
  assign n29940 = ~n29923 & ~n29939;
  assign n29941 = ~n9969 & ~n29940;
  assign n29942 = n9969 & ~n29923;
  assign n29943 = ~n29939 & n29942;
  assign n29944 = ~n35496 & ~n29181;
  assign n29945 = ~n29181 & ~n29514;
  assign n29946 = ~n35496 & n29945;
  assign n29947 = ~n29514 & n29944;
  assign n29948 = n28835 & ~n35595;
  assign n29949 = n29180 & n29945;
  assign n29950 = n28835 & ~n35496;
  assign n29951 = ~n29181 & n29950;
  assign n29952 = ~n29514 & n29951;
  assign n29953 = ~n28835 & ~n35595;
  assign n29954 = ~n29952 & ~n29953;
  assign n29955 = ~n29948 & ~n29949;
  assign n29956 = ~n29943 & ~n35596;
  assign n29957 = ~n29941 & ~n29956;
  assign n29958 = ~n9457 & ~n29957;
  assign n29959 = ~n29183 & ~n29198;
  assign n29960 = ~n29514 & n29959;
  assign n29961 = ~n35498 & ~n29960;
  assign n29962 = n35498 & ~n29198;
  assign n29963 = ~n29183 & n29962;
  assign n29964 = n35498 & n29960;
  assign n29965 = ~n29514 & n29963;
  assign n29966 = ~n29961 & ~n35597;
  assign n29967 = n9457 & ~n29941;
  assign n29968 = ~n29956 & n29967;
  assign n29969 = n9457 & n29957;
  assign n29970 = ~n29966 & ~n35598;
  assign n29971 = ~n29958 & ~n29970;
  assign n29972 = ~n8896 & ~n29971;
  assign n29973 = n8896 & ~n29958;
  assign n29974 = ~n29970 & n29973;
  assign n29975 = ~n35499 & ~n29204;
  assign n29976 = ~n29204 & ~n29514;
  assign n29977 = ~n35499 & n29976;
  assign n29978 = ~n29514 & n29975;
  assign n29979 = n28827 & ~n35599;
  assign n29980 = n29203 & n29976;
  assign n29981 = n28827 & ~n35499;
  assign n29982 = ~n29204 & n29981;
  assign n29983 = ~n29514 & n29982;
  assign n29984 = ~n28827 & ~n35599;
  assign n29985 = ~n29983 & ~n29984;
  assign n29986 = ~n29979 & ~n29980;
  assign n29987 = ~n29974 & ~n35600;
  assign n29988 = ~n29972 & ~n29987;
  assign n29989 = ~n8411 & ~n29988;
  assign n29990 = n8411 & ~n29972;
  assign n29991 = ~n29987 & n29990;
  assign n29992 = n8411 & n29988;
  assign n29993 = ~n29206 & ~n29209;
  assign n29994 = ~n29209 & ~n29514;
  assign n29995 = ~n29206 & n29994;
  assign n29996 = ~n29514 & n29993;
  assign n29997 = n28819 & ~n35602;
  assign n29998 = n29207 & n29994;
  assign n29999 = n28819 & ~n29209;
  assign n30000 = ~n29206 & n29999;
  assign n30001 = ~n29514 & n30000;
  assign n30002 = ~n28819 & ~n35602;
  assign n30003 = ~n30001 & ~n30002;
  assign n30004 = ~n29997 & ~n29998;
  assign n30005 = ~n35601 & ~n35603;
  assign n30006 = ~n29989 & ~n30005;
  assign n30007 = ~n7885 & ~n30006;
  assign n30008 = n7885 & ~n29989;
  assign n30009 = ~n30005 & n30008;
  assign n30010 = ~n35500 & ~n29215;
  assign n30011 = ~n29215 & ~n29514;
  assign n30012 = ~n35500 & n30011;
  assign n30013 = ~n29514 & n30010;
  assign n30014 = n28811 & ~n35604;
  assign n30015 = n29214 & n30011;
  assign n30016 = n28811 & ~n35500;
  assign n30017 = ~n29215 & n30016;
  assign n30018 = ~n29514 & n30017;
  assign n30019 = ~n28811 & ~n35604;
  assign n30020 = ~n30018 & ~n30019;
  assign n30021 = ~n30014 & ~n30015;
  assign n30022 = ~n30009 & ~n35605;
  assign n30023 = ~n30007 & ~n30022;
  assign n30024 = ~n7428 & ~n30023;
  assign n30025 = ~n29217 & ~n29232;
  assign n30026 = ~n29514 & n30025;
  assign n30027 = ~n35502 & ~n30026;
  assign n30028 = n35502 & ~n29232;
  assign n30029 = ~n29217 & n30028;
  assign n30030 = n35502 & n30026;
  assign n30031 = ~n29514 & n30029;
  assign n30032 = ~n30027 & ~n35606;
  assign n30033 = n7428 & ~n30007;
  assign n30034 = ~n30022 & n30033;
  assign n30035 = n7428 & n30023;
  assign n30036 = ~n30032 & ~n35607;
  assign n30037 = ~n30024 & ~n30036;
  assign n30038 = ~n6937 & ~n30037;
  assign n30039 = n6937 & ~n30024;
  assign n30040 = ~n30036 & n30039;
  assign n30041 = ~n35503 & ~n29238;
  assign n30042 = ~n29238 & ~n29514;
  assign n30043 = ~n35503 & n30042;
  assign n30044 = ~n29514 & n30041;
  assign n30045 = n28803 & ~n35608;
  assign n30046 = n29237 & n30042;
  assign n30047 = n28803 & ~n35503;
  assign n30048 = ~n29238 & n30047;
  assign n30049 = ~n29514 & n30048;
  assign n30050 = ~n28803 & ~n35608;
  assign n30051 = ~n30049 & ~n30050;
  assign n30052 = ~n30045 & ~n30046;
  assign n30053 = ~n30040 & ~n35609;
  assign n30054 = ~n30038 & ~n30053;
  assign n30055 = ~n6507 & ~n30054;
  assign n30056 = n6507 & ~n30038;
  assign n30057 = ~n30053 & n30056;
  assign n30058 = n6507 & n30054;
  assign n30059 = ~n29240 & ~n29243;
  assign n30060 = ~n29243 & ~n29514;
  assign n30061 = ~n29240 & n30060;
  assign n30062 = ~n29514 & n30059;
  assign n30063 = n28795 & ~n35611;
  assign n30064 = n29241 & n30060;
  assign n30065 = n28795 & ~n29243;
  assign n30066 = ~n29240 & n30065;
  assign n30067 = ~n29514 & n30066;
  assign n30068 = ~n28795 & ~n35611;
  assign n30069 = ~n30067 & ~n30068;
  assign n30070 = ~n30063 & ~n30064;
  assign n30071 = ~n35610 & ~n35612;
  assign n30072 = ~n30055 & ~n30071;
  assign n30073 = ~n6051 & ~n30072;
  assign n30074 = n6051 & ~n30055;
  assign n30075 = ~n30071 & n30074;
  assign n30076 = ~n35504 & ~n29249;
  assign n30077 = ~n29249 & ~n29514;
  assign n30078 = ~n35504 & n30077;
  assign n30079 = ~n29514 & n30076;
  assign n30080 = n28787 & ~n35613;
  assign n30081 = n29248 & n30077;
  assign n30082 = n28787 & ~n35504;
  assign n30083 = ~n29249 & n30082;
  assign n30084 = ~n29514 & n30083;
  assign n30085 = ~n28787 & ~n35613;
  assign n30086 = ~n30084 & ~n30085;
  assign n30087 = ~n30080 & ~n30081;
  assign n30088 = ~n30075 & ~n35614;
  assign n30089 = ~n30073 & ~n30088;
  assign n30090 = ~n5648 & ~n30089;
  assign n30091 = ~n29251 & ~n29266;
  assign n30092 = ~n29514 & n30091;
  assign n30093 = ~n35506 & ~n30092;
  assign n30094 = n35506 & ~n29266;
  assign n30095 = ~n29251 & n30094;
  assign n30096 = n35506 & n30092;
  assign n30097 = ~n29514 & n30095;
  assign n30098 = ~n30093 & ~n35615;
  assign n30099 = n5648 & ~n30073;
  assign n30100 = ~n30088 & n30099;
  assign n30101 = n5648 & n30089;
  assign n30102 = ~n30098 & ~n35616;
  assign n30103 = ~n30090 & ~n30102;
  assign n30104 = ~n5223 & ~n30103;
  assign n30105 = n5223 & ~n30090;
  assign n30106 = ~n30102 & n30105;
  assign n30107 = ~n35507 & ~n29272;
  assign n30108 = ~n29272 & ~n29514;
  assign n30109 = ~n35507 & n30108;
  assign n30110 = ~n29514 & n30107;
  assign n30111 = n28779 & ~n35617;
  assign n30112 = n29271 & n30108;
  assign n30113 = n28779 & ~n35507;
  assign n30114 = ~n29272 & n30113;
  assign n30115 = ~n29514 & n30114;
  assign n30116 = ~n28779 & ~n35617;
  assign n30117 = ~n30115 & ~n30116;
  assign n30118 = ~n30111 & ~n30112;
  assign n30119 = ~n30106 & ~n35618;
  assign n30120 = ~n30104 & ~n30119;
  assign n30121 = ~n4851 & ~n30120;
  assign n30122 = n4851 & ~n30104;
  assign n30123 = ~n30119 & n30122;
  assign n30124 = n4851 & n30120;
  assign n30125 = ~n29274 & ~n29277;
  assign n30126 = ~n29277 & ~n29514;
  assign n30127 = ~n29274 & n30126;
  assign n30128 = ~n29514 & n30125;
  assign n30129 = n28771 & ~n35620;
  assign n30130 = n29275 & n30126;
  assign n30131 = n28771 & ~n29277;
  assign n30132 = ~n29274 & n30131;
  assign n30133 = ~n29514 & n30132;
  assign n30134 = ~n28771 & ~n35620;
  assign n30135 = ~n30133 & ~n30134;
  assign n30136 = ~n30129 & ~n30130;
  assign n30137 = ~n35619 & ~n35621;
  assign n30138 = ~n30121 & ~n30137;
  assign n30139 = ~n4461 & ~n30138;
  assign n30140 = n4461 & ~n30121;
  assign n30141 = ~n30137 & n30140;
  assign n30142 = ~n35508 & ~n29283;
  assign n30143 = ~n29283 & ~n29514;
  assign n30144 = ~n35508 & n30143;
  assign n30145 = ~n29514 & n30142;
  assign n30146 = n28763 & ~n35622;
  assign n30147 = n29282 & n30143;
  assign n30148 = n28763 & ~n35508;
  assign n30149 = ~n29283 & n30148;
  assign n30150 = ~n29514 & n30149;
  assign n30151 = ~n28763 & ~n35622;
  assign n30152 = ~n30150 & ~n30151;
  assign n30153 = ~n30146 & ~n30147;
  assign n30154 = ~n30141 & ~n35623;
  assign n30155 = ~n30139 & ~n30154;
  assign n30156 = ~n4115 & ~n30155;
  assign n30157 = ~n29285 & ~n29300;
  assign n30158 = ~n29514 & n30157;
  assign n30159 = ~n35510 & ~n30158;
  assign n30160 = n35510 & ~n29300;
  assign n30161 = ~n29285 & n30160;
  assign n30162 = n35510 & n30158;
  assign n30163 = ~n29514 & n30161;
  assign n30164 = ~n30159 & ~n35624;
  assign n30165 = n4115 & ~n30139;
  assign n30166 = ~n30154 & n30165;
  assign n30167 = n4115 & n30155;
  assign n30168 = ~n30164 & ~n35625;
  assign n30169 = ~n30156 & ~n30168;
  assign n30170 = ~n3754 & ~n30169;
  assign n30171 = n3754 & ~n30156;
  assign n30172 = ~n30168 & n30171;
  assign n30173 = ~n35511 & ~n29306;
  assign n30174 = ~n29306 & ~n29514;
  assign n30175 = ~n35511 & n30174;
  assign n30176 = ~n29514 & n30173;
  assign n30177 = n28755 & ~n35626;
  assign n30178 = n29305 & n30174;
  assign n30179 = n28755 & ~n35511;
  assign n30180 = ~n29306 & n30179;
  assign n30181 = ~n29514 & n30180;
  assign n30182 = ~n28755 & ~n35626;
  assign n30183 = ~n30181 & ~n30182;
  assign n30184 = ~n30177 & ~n30178;
  assign n30185 = ~n30172 & ~n35627;
  assign n30186 = ~n30170 & ~n30185;
  assign n30187 = ~n3444 & ~n30186;
  assign n30188 = n3444 & ~n30170;
  assign n30189 = ~n30185 & n30188;
  assign n30190 = n3444 & n30186;
  assign n30191 = ~n29308 & ~n29311;
  assign n30192 = ~n29311 & ~n29514;
  assign n30193 = ~n29308 & n30192;
  assign n30194 = ~n29514 & n30191;
  assign n30195 = n28747 & ~n35629;
  assign n30196 = n29309 & n30192;
  assign n30197 = n28747 & ~n29311;
  assign n30198 = ~n29308 & n30197;
  assign n30199 = ~n29514 & n30198;
  assign n30200 = ~n28747 & ~n35629;
  assign n30201 = ~n30199 & ~n30200;
  assign n30202 = ~n30195 & ~n30196;
  assign n30203 = ~n35628 & ~n35630;
  assign n30204 = ~n30187 & ~n30203;
  assign n30205 = ~n3116 & ~n30204;
  assign n30206 = n3116 & ~n30187;
  assign n30207 = ~n30203 & n30206;
  assign n30208 = ~n35512 & ~n29317;
  assign n30209 = ~n29317 & ~n29514;
  assign n30210 = ~n35512 & n30209;
  assign n30211 = ~n29514 & n30208;
  assign n30212 = n28739 & ~n35631;
  assign n30213 = n29316 & n30209;
  assign n30214 = n28739 & ~n35512;
  assign n30215 = ~n29317 & n30214;
  assign n30216 = ~n29514 & n30215;
  assign n30217 = ~n28739 & ~n35631;
  assign n30218 = ~n30216 & ~n30217;
  assign n30219 = ~n30212 & ~n30213;
  assign n30220 = ~n30207 & ~n35632;
  assign n30221 = ~n30205 & ~n30220;
  assign n30222 = ~n2833 & ~n30221;
  assign n30223 = ~n29319 & ~n29334;
  assign n30224 = ~n29514 & n30223;
  assign n30225 = ~n35514 & ~n30224;
  assign n30226 = n35514 & ~n29334;
  assign n30227 = ~n29319 & n30226;
  assign n30228 = n35514 & n30224;
  assign n30229 = ~n29514 & n30227;
  assign n30230 = ~n30225 & ~n35633;
  assign n30231 = n2833 & ~n30205;
  assign n30232 = ~n30220 & n30231;
  assign n30233 = n2833 & n30221;
  assign n30234 = ~n30230 & ~n35634;
  assign n30235 = ~n30222 & ~n30234;
  assign n30236 = ~n2536 & ~n30235;
  assign n30237 = n2536 & ~n30222;
  assign n30238 = ~n30234 & n30237;
  assign n30239 = ~n35515 & ~n29340;
  assign n30240 = ~n29340 & ~n29514;
  assign n30241 = ~n35515 & n30240;
  assign n30242 = ~n29514 & n30239;
  assign n30243 = n28731 & ~n35635;
  assign n30244 = n29339 & n30240;
  assign n30245 = n28731 & ~n35515;
  assign n30246 = ~n29340 & n30245;
  assign n30247 = ~n29514 & n30246;
  assign n30248 = ~n28731 & ~n35635;
  assign n30249 = ~n30247 & ~n30248;
  assign n30250 = ~n30243 & ~n30244;
  assign n30251 = ~n30238 & ~n35636;
  assign n30252 = ~n30236 & ~n30251;
  assign n30253 = ~n2283 & ~n30252;
  assign n30254 = n2283 & ~n30236;
  assign n30255 = ~n30251 & n30254;
  assign n30256 = n2283 & n30252;
  assign n30257 = ~n29342 & ~n29345;
  assign n30258 = ~n29345 & ~n29514;
  assign n30259 = ~n29342 & n30258;
  assign n30260 = ~n29514 & n30257;
  assign n30261 = n28723 & ~n35638;
  assign n30262 = n29343 & n30258;
  assign n30263 = n28723 & ~n29345;
  assign n30264 = ~n29342 & n30263;
  assign n30265 = ~n29514 & n30264;
  assign n30266 = ~n28723 & ~n35638;
  assign n30267 = ~n30265 & ~n30266;
  assign n30268 = ~n30261 & ~n30262;
  assign n30269 = ~n35637 & ~n35639;
  assign n30270 = ~n30253 & ~n30269;
  assign n30271 = ~n2021 & ~n30270;
  assign n30272 = n2021 & ~n30253;
  assign n30273 = ~n30269 & n30272;
  assign n30274 = ~n35516 & ~n29351;
  assign n30275 = ~n29351 & ~n29514;
  assign n30276 = ~n35516 & n30275;
  assign n30277 = ~n29514 & n30274;
  assign n30278 = n28715 & ~n35640;
  assign n30279 = n29350 & n30275;
  assign n30280 = n28715 & ~n35516;
  assign n30281 = ~n29351 & n30280;
  assign n30282 = ~n29514 & n30281;
  assign n30283 = ~n28715 & ~n35640;
  assign n30284 = ~n30282 & ~n30283;
  assign n30285 = ~n30278 & ~n30279;
  assign n30286 = ~n30273 & ~n35641;
  assign n30287 = ~n30271 & ~n30286;
  assign n30288 = ~n1796 & ~n30287;
  assign n30289 = ~n29353 & ~n29368;
  assign n30290 = ~n29514 & n30289;
  assign n30291 = ~n35518 & ~n30290;
  assign n30292 = n35518 & ~n29368;
  assign n30293 = ~n29353 & n30292;
  assign n30294 = n35518 & n30290;
  assign n30295 = ~n29514 & n30293;
  assign n30296 = ~n30291 & ~n35642;
  assign n30297 = n1796 & ~n30271;
  assign n30298 = ~n30286 & n30297;
  assign n30299 = n1796 & n30287;
  assign n30300 = ~n30296 & ~n35643;
  assign n30301 = ~n30288 & ~n30300;
  assign n30302 = ~n1567 & ~n30301;
  assign n30303 = n1567 & ~n30288;
  assign n30304 = ~n30300 & n30303;
  assign n30305 = ~n35519 & ~n29374;
  assign n30306 = ~n29374 & ~n29514;
  assign n30307 = ~n35519 & n30306;
  assign n30308 = ~n29514 & n30305;
  assign n30309 = n28707 & ~n35644;
  assign n30310 = n29373 & n30306;
  assign n30311 = n28707 & ~n35519;
  assign n30312 = ~n29374 & n30311;
  assign n30313 = ~n29514 & n30312;
  assign n30314 = ~n28707 & ~n35644;
  assign n30315 = ~n30313 & ~n30314;
  assign n30316 = ~n30309 & ~n30310;
  assign n30317 = ~n30304 & ~n35645;
  assign n30318 = ~n30302 & ~n30317;
  assign n30319 = ~n1374 & ~n30318;
  assign n30320 = n1374 & ~n30302;
  assign n30321 = ~n30317 & n30320;
  assign n30322 = n1374 & n30318;
  assign n30323 = ~n29376 & ~n29379;
  assign n30324 = ~n29379 & ~n29514;
  assign n30325 = ~n29376 & n30324;
  assign n30326 = ~n29514 & n30323;
  assign n30327 = n28699 & ~n35647;
  assign n30328 = n29377 & n30324;
  assign n30329 = n28699 & ~n29379;
  assign n30330 = ~n29376 & n30329;
  assign n30331 = ~n29514 & n30330;
  assign n30332 = ~n28699 & ~n35647;
  assign n30333 = ~n30331 & ~n30332;
  assign n30334 = ~n30327 & ~n30328;
  assign n30335 = ~n35646 & ~n35648;
  assign n30336 = ~n30319 & ~n30335;
  assign n30337 = ~n1179 & ~n30336;
  assign n30338 = n1179 & ~n30319;
  assign n30339 = ~n30335 & n30338;
  assign n30340 = ~n35520 & ~n29385;
  assign n30341 = ~n29385 & ~n29514;
  assign n30342 = ~n35520 & n30341;
  assign n30343 = ~n29514 & n30340;
  assign n30344 = n28691 & ~n35649;
  assign n30345 = n29384 & n30341;
  assign n30346 = n28691 & ~n35520;
  assign n30347 = ~n29385 & n30346;
  assign n30348 = ~n29514 & n30347;
  assign n30349 = ~n28691 & ~n35649;
  assign n30350 = ~n30348 & ~n30349;
  assign n30351 = ~n30344 & ~n30345;
  assign n30352 = ~n30339 & ~n35650;
  assign n30353 = ~n30337 & ~n30352;
  assign n30354 = ~n1016 & ~n30353;
  assign n30355 = ~n29387 & ~n29402;
  assign n30356 = ~n29514 & n30355;
  assign n30357 = ~n35522 & ~n30356;
  assign n30358 = n35522 & ~n29402;
  assign n30359 = ~n29387 & n30358;
  assign n30360 = n35522 & n30356;
  assign n30361 = ~n29514 & n30359;
  assign n30362 = ~n30357 & ~n35651;
  assign n30363 = n1016 & ~n30337;
  assign n30364 = ~n30352 & n30363;
  assign n30365 = n1016 & n30353;
  assign n30366 = ~n30362 & ~n35652;
  assign n30367 = ~n30354 & ~n30366;
  assign n30368 = ~n855 & ~n30367;
  assign n30369 = n855 & ~n30354;
  assign n30370 = ~n30366 & n30369;
  assign n30371 = ~n35523 & ~n29408;
  assign n30372 = ~n29408 & ~n29514;
  assign n30373 = ~n35523 & n30372;
  assign n30374 = ~n29514 & n30371;
  assign n30375 = n28683 & ~n35653;
  assign n30376 = n29407 & n30372;
  assign n30377 = n28683 & ~n35523;
  assign n30378 = ~n29408 & n30377;
  assign n30379 = ~n29514 & n30378;
  assign n30380 = ~n28683 & ~n35653;
  assign n30381 = ~n30379 & ~n30380;
  assign n30382 = ~n30375 & ~n30376;
  assign n30383 = ~n30370 & ~n35654;
  assign n30384 = ~n30368 & ~n30383;
  assign n30385 = ~n720 & ~n30384;
  assign n30386 = n720 & ~n30368;
  assign n30387 = ~n30383 & n30386;
  assign n30388 = n720 & n30384;
  assign n30389 = ~n29410 & ~n29413;
  assign n30390 = ~n29413 & ~n29514;
  assign n30391 = ~n29410 & n30390;
  assign n30392 = ~n29514 & n30389;
  assign n30393 = n28675 & ~n35656;
  assign n30394 = n29411 & n30390;
  assign n30395 = n28675 & ~n29413;
  assign n30396 = ~n29410 & n30395;
  assign n30397 = ~n29514 & n30396;
  assign n30398 = ~n28675 & ~n35656;
  assign n30399 = ~n30397 & ~n30398;
  assign n30400 = ~n30393 & ~n30394;
  assign n30401 = ~n35655 & ~n35657;
  assign n30402 = ~n30385 & ~n30401;
  assign n30403 = ~n592 & ~n30402;
  assign n30404 = n592 & ~n30385;
  assign n30405 = ~n30401 & n30404;
  assign n30406 = ~n35524 & ~n29419;
  assign n30407 = ~n29419 & ~n29514;
  assign n30408 = ~n35524 & n30407;
  assign n30409 = ~n29514 & n30406;
  assign n30410 = n28667 & ~n35658;
  assign n30411 = n29418 & n30407;
  assign n30412 = n28667 & ~n35524;
  assign n30413 = ~n29419 & n30412;
  assign n30414 = ~n29514 & n30413;
  assign n30415 = ~n28667 & ~n35658;
  assign n30416 = ~n30414 & ~n30415;
  assign n30417 = ~n30410 & ~n30411;
  assign n30418 = ~n30405 & ~n35659;
  assign n30419 = ~n30403 & ~n30418;
  assign n30420 = ~n487 & ~n30419;
  assign n30421 = ~n29421 & ~n29436;
  assign n30422 = ~n29514 & n30421;
  assign n30423 = ~n35526 & ~n30422;
  assign n30424 = n35526 & ~n29436;
  assign n30425 = ~n29421 & n30424;
  assign n30426 = n35526 & n30422;
  assign n30427 = ~n29514 & n30425;
  assign n30428 = ~n30423 & ~n35660;
  assign n30429 = n487 & ~n30403;
  assign n30430 = ~n30418 & n30429;
  assign n30431 = n487 & n30419;
  assign n30432 = ~n30428 & ~n35661;
  assign n30433 = ~n30420 & ~n30432;
  assign n30434 = ~n393 & ~n30433;
  assign n30435 = n393 & ~n30420;
  assign n30436 = ~n30432 & n30435;
  assign n30437 = ~n35527 & ~n29442;
  assign n30438 = ~n29442 & ~n29514;
  assign n30439 = ~n35527 & n30438;
  assign n30440 = ~n29514 & n30437;
  assign n30441 = n28659 & ~n35662;
  assign n30442 = n29441 & n30438;
  assign n30443 = n28659 & ~n35527;
  assign n30444 = ~n29442 & n30443;
  assign n30445 = ~n29514 & n30444;
  assign n30446 = ~n28659 & ~n35662;
  assign n30447 = ~n30445 & ~n30446;
  assign n30448 = ~n30441 & ~n30442;
  assign n30449 = ~n30436 & ~n35663;
  assign n30450 = ~n30434 & ~n30449;
  assign n30451 = ~n321 & ~n30450;
  assign n30452 = n321 & ~n30434;
  assign n30453 = ~n30449 & n30452;
  assign n30454 = n321 & n30450;
  assign n30455 = ~n29444 & ~n29447;
  assign n30456 = ~n29447 & ~n29514;
  assign n30457 = ~n29444 & n30456;
  assign n30458 = ~n29514 & n30455;
  assign n30459 = n28651 & ~n35665;
  assign n30460 = n29445 & n30456;
  assign n30461 = n28651 & ~n29447;
  assign n30462 = ~n29444 & n30461;
  assign n30463 = ~n29514 & n30462;
  assign n30464 = ~n28651 & ~n35665;
  assign n30465 = ~n30463 & ~n30464;
  assign n30466 = ~n30459 & ~n30460;
  assign n30467 = ~n35664 & ~n35666;
  assign n30468 = ~n30451 & ~n30467;
  assign n30469 = ~n263 & ~n30468;
  assign n30470 = n263 & ~n30451;
  assign n30471 = ~n30467 & n30470;
  assign n30472 = ~n35528 & ~n29453;
  assign n30473 = ~n29514 & n30472;
  assign n30474 = n28643 & ~n30473;
  assign n30475 = ~n28643 & n30473;
  assign n30476 = n28643 & ~n35528;
  assign n30477 = ~n29453 & n30476;
  assign n30478 = ~n29514 & n30477;
  assign n30479 = ~n28643 & ~n30473;
  assign n30480 = ~n30478 & ~n30479;
  assign n30481 = ~n30474 & ~n30475;
  assign n30482 = ~n30471 & ~n35667;
  assign n30483 = ~n30469 & ~n30482;
  assign n30484 = ~n214 & ~n30483;
  assign n30485 = n214 & ~n30469;
  assign n30486 = ~n30482 & n30485;
  assign n30487 = n214 & n30483;
  assign n30488 = ~n35536 & ~n35668;
  assign n30489 = ~n30484 & ~n30488;
  assign n30490 = ~n197 & ~n30489;
  assign n30491 = n197 & ~n30484;
  assign n30492 = ~n30488 & n30491;
  assign n30493 = ~n29460 & ~n35530;
  assign n30494 = ~n29460 & ~n29514;
  assign n30495 = ~n35530 & n30494;
  assign n30496 = ~n29514 & n30493;
  assign n30497 = n29468 & ~n35669;
  assign n30498 = n29472 & n30494;
  assign n30499 = n29468 & ~n35530;
  assign n30500 = ~n29460 & n30499;
  assign n30501 = ~n29514 & n30500;
  assign n30502 = ~n29468 & ~n35669;
  assign n30503 = ~n30501 & ~n30502;
  assign n30504 = ~n30497 & ~n30498;
  assign n30505 = ~n30492 & ~n35670;
  assign n30506 = ~n30490 & ~n30505;
  assign n30507 = ~n29474 & ~n29476;
  assign n30508 = ~n29514 & n30507;
  assign n30509 = ~n35532 & ~n30508;
  assign n30510 = ~n29474 & n35532;
  assign n30511 = ~n29476 & n30510;
  assign n30512 = n35532 & n30508;
  assign n30513 = ~n29514 & n30511;
  assign n30514 = ~n30509 & ~n35671;
  assign n30515 = ~n29490 & ~n29498;
  assign n30516 = ~n29498 & ~n29514;
  assign n30517 = ~n29490 & n30516;
  assign n30518 = ~n29514 & n30515;
  assign n30519 = ~n35535 & ~n35672;
  assign n30520 = ~n30514 & n30519;
  assign n30521 = ~n30506 & n30520;
  assign n30522 = n193 & ~n30521;
  assign n30523 = ~n30490 & n30514;
  assign n30524 = ~n30505 & n30523;
  assign n30525 = n30506 & n30514;
  assign n30526 = n29490 & ~n30516;
  assign n30527 = ~n193 & ~n30515;
  assign n30528 = ~n30526 & n30527;
  assign n30529 = ~n35673 & ~n30528;
  assign n30530 = ~n30522 & n30529;
  assign n30531 = ~n30484 & ~n35668;
  assign n30532 = ~n30530 & n30531;
  assign n30533 = n35536 & ~n30532;
  assign n30534 = ~n35536 & n30532;
  assign n30535 = ~n35536 & ~n30532;
  assign n30536 = n35536 & ~n30484;
  assign n30537 = ~n35668 & n30536;
  assign n30538 = ~n30530 & n30537;
  assign n30539 = ~n30535 & ~n30538;
  assign n30540 = ~n30533 & ~n30534;
  assign n30541 = n197 & n35674;
  assign n30542 = ~n197 & ~n35674;
  assign n30543 = ~n30469 & ~n30471;
  assign n30544 = ~n30530 & n30543;
  assign n30545 = ~n35667 & n30544;
  assign n30546 = n35667 & ~n30544;
  assign n30547 = ~n35667 & ~n30544;
  assign n30548 = ~n30471 & n35667;
  assign n30549 = ~n30469 & n30548;
  assign n30550 = ~n30530 & n30549;
  assign n30551 = ~n30547 & ~n30550;
  assign n30552 = ~n30545 & ~n30546;
  assign n30553 = n214 & n35675;
  assign n30554 = ~n30434 & ~n30436;
  assign n30555 = ~n30530 & n30554;
  assign n30556 = ~n35663 & ~n30555;
  assign n30557 = ~n30436 & n35663;
  assign n30558 = ~n30434 & n30557;
  assign n30559 = n35663 & n30555;
  assign n30560 = ~n30530 & n30558;
  assign n30561 = ~n30556 & ~n35676;
  assign n30562 = ~n321 & ~n30561;
  assign n30563 = ~n30420 & ~n35661;
  assign n30564 = ~n30420 & ~n30530;
  assign n30565 = ~n35661 & n30564;
  assign n30566 = ~n30530 & n30563;
  assign n30567 = n30428 & ~n35677;
  assign n30568 = n30432 & n30564;
  assign n30569 = ~n30428 & ~n35677;
  assign n30570 = ~n30420 & n30428;
  assign n30571 = ~n35661 & n30570;
  assign n30572 = ~n30530 & n30571;
  assign n30573 = ~n30569 & ~n30572;
  assign n30574 = ~n30567 & ~n30568;
  assign n30575 = n393 & n35678;
  assign n30576 = ~n393 & ~n35678;
  assign n30577 = ~n30403 & ~n30405;
  assign n30578 = ~n30530 & n30577;
  assign n30579 = ~n35659 & ~n30578;
  assign n30580 = ~n30405 & n35659;
  assign n30581 = ~n30403 & n30580;
  assign n30582 = n35659 & n30578;
  assign n30583 = ~n30530 & n30581;
  assign n30584 = ~n30579 & ~n35679;
  assign n30585 = n487 & n30584;
  assign n30586 = ~n487 & ~n30584;
  assign n30587 = ~n30385 & ~n35655;
  assign n30588 = ~n30530 & n30587;
  assign n30589 = ~n35657 & ~n30588;
  assign n30590 = ~n30385 & n35657;
  assign n30591 = ~n35655 & n30590;
  assign n30592 = n35657 & n30588;
  assign n30593 = ~n30530 & n30591;
  assign n30594 = ~n30589 & ~n35680;
  assign n30595 = n592 & n30594;
  assign n30596 = ~n592 & ~n30594;
  assign n30597 = ~n30368 & ~n30370;
  assign n30598 = ~n30530 & n30597;
  assign n30599 = ~n35654 & ~n30598;
  assign n30600 = ~n30370 & n35654;
  assign n30601 = ~n30368 & n30600;
  assign n30602 = n35654 & n30598;
  assign n30603 = ~n30530 & n30601;
  assign n30604 = ~n30599 & ~n35681;
  assign n30605 = n720 & n30604;
  assign n30606 = ~n720 & ~n30604;
  assign n30607 = ~n30354 & ~n35652;
  assign n30608 = ~n30354 & ~n30530;
  assign n30609 = ~n35652 & n30608;
  assign n30610 = ~n30530 & n30607;
  assign n30611 = n30362 & ~n35682;
  assign n30612 = n30366 & n30608;
  assign n30613 = ~n30362 & ~n35682;
  assign n30614 = ~n30354 & n30362;
  assign n30615 = ~n35652 & n30614;
  assign n30616 = ~n30530 & n30615;
  assign n30617 = ~n30613 & ~n30616;
  assign n30618 = ~n30611 & ~n30612;
  assign n30619 = n855 & n35683;
  assign n30620 = ~n855 & ~n35683;
  assign n30621 = ~n30337 & ~n30339;
  assign n30622 = ~n30530 & n30621;
  assign n30623 = ~n35650 & ~n30622;
  assign n30624 = ~n30339 & n35650;
  assign n30625 = ~n30337 & n30624;
  assign n30626 = n35650 & n30622;
  assign n30627 = ~n30530 & n30625;
  assign n30628 = ~n30623 & ~n35684;
  assign n30629 = n1016 & n30628;
  assign n30630 = ~n1016 & ~n30628;
  assign n30631 = ~n30319 & ~n35646;
  assign n30632 = ~n30530 & n30631;
  assign n30633 = ~n35648 & ~n30632;
  assign n30634 = ~n30319 & n35648;
  assign n30635 = ~n35646 & n30634;
  assign n30636 = n35648 & n30632;
  assign n30637 = ~n30530 & n30635;
  assign n30638 = ~n30633 & ~n35685;
  assign n30639 = n1179 & n30638;
  assign n30640 = ~n1179 & ~n30638;
  assign n30641 = ~n30302 & ~n30304;
  assign n30642 = ~n30530 & n30641;
  assign n30643 = ~n35645 & ~n30642;
  assign n30644 = ~n30304 & n35645;
  assign n30645 = ~n30302 & n30644;
  assign n30646 = n35645 & n30642;
  assign n30647 = ~n30530 & n30645;
  assign n30648 = ~n30643 & ~n35686;
  assign n30649 = n1374 & n30648;
  assign n30650 = ~n1374 & ~n30648;
  assign n30651 = ~n30288 & ~n35643;
  assign n30652 = ~n30288 & ~n30530;
  assign n30653 = ~n35643 & n30652;
  assign n30654 = ~n30530 & n30651;
  assign n30655 = n30296 & ~n35687;
  assign n30656 = n30300 & n30652;
  assign n30657 = ~n30296 & ~n35687;
  assign n30658 = ~n30288 & n30296;
  assign n30659 = ~n35643 & n30658;
  assign n30660 = ~n30530 & n30659;
  assign n30661 = ~n30657 & ~n30660;
  assign n30662 = ~n30655 & ~n30656;
  assign n30663 = n1567 & n35688;
  assign n30664 = ~n1567 & ~n35688;
  assign n30665 = ~n30271 & ~n30273;
  assign n30666 = ~n30530 & n30665;
  assign n30667 = ~n35641 & ~n30666;
  assign n30668 = ~n30273 & n35641;
  assign n30669 = ~n30271 & n30668;
  assign n30670 = n35641 & n30666;
  assign n30671 = ~n30530 & n30669;
  assign n30672 = ~n30667 & ~n35689;
  assign n30673 = n1796 & n30672;
  assign n30674 = ~n1796 & ~n30672;
  assign n30675 = ~n30253 & ~n35637;
  assign n30676 = ~n30530 & n30675;
  assign n30677 = ~n35639 & ~n30676;
  assign n30678 = ~n30253 & n35639;
  assign n30679 = ~n35637 & n30678;
  assign n30680 = n35639 & n30676;
  assign n30681 = ~n30530 & n30679;
  assign n30682 = ~n30677 & ~n35690;
  assign n30683 = n2021 & n30682;
  assign n30684 = ~n2021 & ~n30682;
  assign n30685 = ~n30236 & ~n30238;
  assign n30686 = ~n30530 & n30685;
  assign n30687 = ~n35636 & ~n30686;
  assign n30688 = ~n30238 & n35636;
  assign n30689 = ~n30236 & n30688;
  assign n30690 = n35636 & n30686;
  assign n30691 = ~n30530 & n30689;
  assign n30692 = ~n30687 & ~n35691;
  assign n30693 = n2283 & n30692;
  assign n30694 = ~n2283 & ~n30692;
  assign n30695 = ~n30222 & ~n35634;
  assign n30696 = ~n30222 & ~n30530;
  assign n30697 = ~n35634 & n30696;
  assign n30698 = ~n30530 & n30695;
  assign n30699 = n30230 & ~n35692;
  assign n30700 = n30234 & n30696;
  assign n30701 = ~n30230 & ~n35692;
  assign n30702 = ~n30222 & n30230;
  assign n30703 = ~n35634 & n30702;
  assign n30704 = ~n30530 & n30703;
  assign n30705 = ~n30701 & ~n30704;
  assign n30706 = ~n30699 & ~n30700;
  assign n30707 = n2536 & n35693;
  assign n30708 = ~n2536 & ~n35693;
  assign n30709 = ~n30205 & ~n30207;
  assign n30710 = ~n30530 & n30709;
  assign n30711 = ~n35632 & ~n30710;
  assign n30712 = ~n30207 & n35632;
  assign n30713 = ~n30205 & n30712;
  assign n30714 = n35632 & n30710;
  assign n30715 = ~n30530 & n30713;
  assign n30716 = ~n30711 & ~n35694;
  assign n30717 = n2833 & n30716;
  assign n30718 = ~n2833 & ~n30716;
  assign n30719 = ~n30187 & ~n35628;
  assign n30720 = ~n30530 & n30719;
  assign n30721 = ~n35630 & ~n30720;
  assign n30722 = ~n30187 & n35630;
  assign n30723 = ~n35628 & n30722;
  assign n30724 = n35630 & n30720;
  assign n30725 = ~n30530 & n30723;
  assign n30726 = ~n30721 & ~n35695;
  assign n30727 = n3116 & n30726;
  assign n30728 = ~n3116 & ~n30726;
  assign n30729 = ~n30170 & ~n30172;
  assign n30730 = ~n30530 & n30729;
  assign n30731 = ~n35627 & ~n30730;
  assign n30732 = ~n30172 & n35627;
  assign n30733 = ~n30170 & n30732;
  assign n30734 = n35627 & n30730;
  assign n30735 = ~n30530 & n30733;
  assign n30736 = ~n30731 & ~n35696;
  assign n30737 = n3444 & n30736;
  assign n30738 = ~n3444 & ~n30736;
  assign n30739 = ~n30156 & ~n35625;
  assign n30740 = ~n30156 & ~n30530;
  assign n30741 = ~n35625 & n30740;
  assign n30742 = ~n30530 & n30739;
  assign n30743 = n30164 & ~n35697;
  assign n30744 = n30168 & n30740;
  assign n30745 = ~n30164 & ~n35697;
  assign n30746 = ~n30156 & n30164;
  assign n30747 = ~n35625 & n30746;
  assign n30748 = ~n30530 & n30747;
  assign n30749 = ~n30745 & ~n30748;
  assign n30750 = ~n30743 & ~n30744;
  assign n30751 = n3754 & n35698;
  assign n30752 = ~n3754 & ~n35698;
  assign n30753 = ~n30139 & ~n30141;
  assign n30754 = ~n30530 & n30753;
  assign n30755 = ~n35623 & ~n30754;
  assign n30756 = ~n30141 & n35623;
  assign n30757 = ~n30139 & n30756;
  assign n30758 = n35623 & n30754;
  assign n30759 = ~n30530 & n30757;
  assign n30760 = ~n30755 & ~n35699;
  assign n30761 = n4115 & n30760;
  assign n30762 = ~n4115 & ~n30760;
  assign n30763 = ~n30121 & ~n35619;
  assign n30764 = ~n30530 & n30763;
  assign n30765 = ~n35621 & ~n30764;
  assign n30766 = ~n30121 & n35621;
  assign n30767 = ~n35619 & n30766;
  assign n30768 = n35621 & n30764;
  assign n30769 = ~n30530 & n30767;
  assign n30770 = ~n30765 & ~n35700;
  assign n30771 = n4461 & n30770;
  assign n30772 = ~n4461 & ~n30770;
  assign n30773 = ~n30104 & ~n30106;
  assign n30774 = ~n30530 & n30773;
  assign n30775 = ~n35618 & ~n30774;
  assign n30776 = ~n30106 & n35618;
  assign n30777 = ~n30104 & n30776;
  assign n30778 = n35618 & n30774;
  assign n30779 = ~n30530 & n30777;
  assign n30780 = ~n30775 & ~n35701;
  assign n30781 = n4851 & n30780;
  assign n30782 = ~n4851 & ~n30780;
  assign n30783 = ~n30090 & ~n35616;
  assign n30784 = ~n30090 & ~n30530;
  assign n30785 = ~n35616 & n30784;
  assign n30786 = ~n30530 & n30783;
  assign n30787 = n30098 & ~n35702;
  assign n30788 = n30102 & n30784;
  assign n30789 = ~n30098 & ~n35702;
  assign n30790 = ~n30090 & n30098;
  assign n30791 = ~n35616 & n30790;
  assign n30792 = ~n30530 & n30791;
  assign n30793 = ~n30789 & ~n30792;
  assign n30794 = ~n30787 & ~n30788;
  assign n30795 = n5223 & n35703;
  assign n30796 = ~n5223 & ~n35703;
  assign n30797 = ~n30073 & ~n30075;
  assign n30798 = ~n30530 & n30797;
  assign n30799 = ~n35614 & ~n30798;
  assign n30800 = ~n30075 & n35614;
  assign n30801 = ~n30073 & n30800;
  assign n30802 = n35614 & n30798;
  assign n30803 = ~n30530 & n30801;
  assign n30804 = ~n30799 & ~n35704;
  assign n30805 = n5648 & n30804;
  assign n30806 = ~n5648 & ~n30804;
  assign n30807 = ~n30055 & ~n35610;
  assign n30808 = ~n30530 & n30807;
  assign n30809 = ~n35612 & ~n30808;
  assign n30810 = ~n30055 & n35612;
  assign n30811 = ~n35610 & n30810;
  assign n30812 = n35612 & n30808;
  assign n30813 = ~n30530 & n30811;
  assign n30814 = ~n30809 & ~n35705;
  assign n30815 = n6051 & n30814;
  assign n30816 = ~n6051 & ~n30814;
  assign n30817 = ~n30038 & ~n30040;
  assign n30818 = ~n30530 & n30817;
  assign n30819 = ~n35609 & ~n30818;
  assign n30820 = ~n30040 & n35609;
  assign n30821 = ~n30038 & n30820;
  assign n30822 = n35609 & n30818;
  assign n30823 = ~n30530 & n30821;
  assign n30824 = ~n30819 & ~n35706;
  assign n30825 = n6507 & n30824;
  assign n30826 = ~n6507 & ~n30824;
  assign n30827 = ~n30024 & ~n35607;
  assign n30828 = ~n30024 & ~n30530;
  assign n30829 = ~n35607 & n30828;
  assign n30830 = ~n30530 & n30827;
  assign n30831 = n30032 & ~n35707;
  assign n30832 = n30036 & n30828;
  assign n30833 = ~n30032 & ~n35707;
  assign n30834 = ~n30024 & n30032;
  assign n30835 = ~n35607 & n30834;
  assign n30836 = ~n30530 & n30835;
  assign n30837 = ~n30833 & ~n30836;
  assign n30838 = ~n30831 & ~n30832;
  assign n30839 = n6937 & n35708;
  assign n30840 = ~n6937 & ~n35708;
  assign n30841 = ~n30007 & ~n30009;
  assign n30842 = ~n30530 & n30841;
  assign n30843 = ~n35605 & ~n30842;
  assign n30844 = ~n30009 & n35605;
  assign n30845 = ~n30007 & n30844;
  assign n30846 = n35605 & n30842;
  assign n30847 = ~n30530 & n30845;
  assign n30848 = ~n30843 & ~n35709;
  assign n30849 = n7428 & n30848;
  assign n30850 = ~n7428 & ~n30848;
  assign n30851 = ~n29989 & ~n35601;
  assign n30852 = ~n30530 & n30851;
  assign n30853 = ~n35603 & ~n30852;
  assign n30854 = ~n29989 & n35603;
  assign n30855 = ~n35601 & n30854;
  assign n30856 = n35603 & n30852;
  assign n30857 = ~n30530 & n30855;
  assign n30858 = ~n30853 & ~n35710;
  assign n30859 = n7885 & n30858;
  assign n30860 = ~n7885 & ~n30858;
  assign n30861 = ~n29972 & ~n29974;
  assign n30862 = ~n30530 & n30861;
  assign n30863 = ~n35600 & ~n30862;
  assign n30864 = ~n29974 & n35600;
  assign n30865 = ~n29972 & n30864;
  assign n30866 = n35600 & n30862;
  assign n30867 = ~n30530 & n30865;
  assign n30868 = ~n30863 & ~n35711;
  assign n30869 = n8411 & n30868;
  assign n30870 = ~n8411 & ~n30868;
  assign n30871 = ~n29958 & ~n35598;
  assign n30872 = ~n29958 & ~n30530;
  assign n30873 = ~n35598 & n30872;
  assign n30874 = ~n30530 & n30871;
  assign n30875 = n29966 & ~n35712;
  assign n30876 = n29970 & n30872;
  assign n30877 = ~n29966 & ~n35712;
  assign n30878 = ~n29958 & n29966;
  assign n30879 = ~n35598 & n30878;
  assign n30880 = ~n30530 & n30879;
  assign n30881 = ~n30877 & ~n30880;
  assign n30882 = ~n30875 & ~n30876;
  assign n30883 = n8896 & n35713;
  assign n30884 = ~n8896 & ~n35713;
  assign n30885 = ~n29941 & ~n29943;
  assign n30886 = ~n30530 & n30885;
  assign n30887 = ~n35596 & ~n30886;
  assign n30888 = ~n29943 & n35596;
  assign n30889 = ~n29941 & n30888;
  assign n30890 = n35596 & n30886;
  assign n30891 = ~n30530 & n30889;
  assign n30892 = ~n30887 & ~n35714;
  assign n30893 = n9457 & n30892;
  assign n30894 = ~n9457 & ~n30892;
  assign n30895 = ~n29923 & ~n35592;
  assign n30896 = ~n30530 & n30895;
  assign n30897 = ~n35594 & ~n30896;
  assign n30898 = ~n29923 & n35594;
  assign n30899 = ~n35592 & n30898;
  assign n30900 = n35594 & n30896;
  assign n30901 = ~n30530 & n30899;
  assign n30902 = ~n30897 & ~n35715;
  assign n30903 = n9969 & n30902;
  assign n30904 = ~n9969 & ~n30902;
  assign n30905 = ~n29906 & ~n29908;
  assign n30906 = ~n30530 & n30905;
  assign n30907 = ~n35591 & ~n30906;
  assign n30908 = ~n29908 & n35591;
  assign n30909 = ~n29906 & n30908;
  assign n30910 = n35591 & n30906;
  assign n30911 = ~n30530 & n30909;
  assign n30912 = ~n30907 & ~n35716;
  assign n30913 = n10555 & n30912;
  assign n30914 = ~n10555 & ~n30912;
  assign n30915 = ~n29892 & ~n35589;
  assign n30916 = ~n29892 & ~n30530;
  assign n30917 = ~n35589 & n30916;
  assign n30918 = ~n30530 & n30915;
  assign n30919 = n29900 & ~n35717;
  assign n30920 = n29904 & n30916;
  assign n30921 = ~n29900 & ~n35717;
  assign n30922 = ~n29892 & n29900;
  assign n30923 = ~n35589 & n30922;
  assign n30924 = ~n30530 & n30923;
  assign n30925 = ~n30921 & ~n30924;
  assign n30926 = ~n30919 & ~n30920;
  assign n30927 = n11097 & n35718;
  assign n30928 = ~n11097 & ~n35718;
  assign n30929 = ~n29875 & ~n29877;
  assign n30930 = ~n30530 & n30929;
  assign n30931 = ~n35587 & ~n30930;
  assign n30932 = ~n29877 & n35587;
  assign n30933 = ~n29875 & n30932;
  assign n30934 = n35587 & n30930;
  assign n30935 = ~n30530 & n30933;
  assign n30936 = ~n30931 & ~n35719;
  assign n30937 = n11719 & n30936;
  assign n30938 = ~n11719 & ~n30936;
  assign n30939 = ~n29857 & ~n35583;
  assign n30940 = ~n30530 & n30939;
  assign n30941 = ~n35585 & ~n30940;
  assign n30942 = ~n29857 & n35585;
  assign n30943 = ~n35583 & n30942;
  assign n30944 = n35585 & n30940;
  assign n30945 = ~n30530 & n30943;
  assign n30946 = ~n30941 & ~n35720;
  assign n30947 = n12296 & n30946;
  assign n30948 = ~n12296 & ~n30946;
  assign n30949 = ~n29840 & ~n29842;
  assign n30950 = ~n30530 & n30949;
  assign n30951 = ~n35582 & ~n30950;
  assign n30952 = ~n29842 & n35582;
  assign n30953 = ~n29840 & n30952;
  assign n30954 = n35582 & n30950;
  assign n30955 = ~n30530 & n30953;
  assign n30956 = ~n30951 & ~n35721;
  assign n30957 = n12948 & n30956;
  assign n30958 = ~n12948 & ~n30956;
  assign n30959 = ~n29826 & ~n35580;
  assign n30960 = ~n29826 & ~n30530;
  assign n30961 = ~n35580 & n30960;
  assign n30962 = ~n30530 & n30959;
  assign n30963 = n29834 & ~n35722;
  assign n30964 = n29838 & n30960;
  assign n30965 = ~n29834 & ~n35722;
  assign n30966 = ~n29826 & n29834;
  assign n30967 = ~n35580 & n30966;
  assign n30968 = ~n30530 & n30967;
  assign n30969 = ~n30965 & ~n30968;
  assign n30970 = ~n30963 & ~n30964;
  assign n30971 = n13548 & n35723;
  assign n30972 = ~n13548 & ~n35723;
  assign n30973 = ~n29809 & ~n29811;
  assign n30974 = ~n30530 & n30973;
  assign n30975 = ~n35578 & ~n30974;
  assign n30976 = ~n29811 & n35578;
  assign n30977 = ~n29809 & n30976;
  assign n30978 = n35578 & n30974;
  assign n30979 = ~n30530 & n30977;
  assign n30980 = ~n30975 & ~n35724;
  assign n30981 = n14233 & n30980;
  assign n30982 = ~n14233 & ~n30980;
  assign n30983 = ~n29791 & ~n35574;
  assign n30984 = ~n30530 & n30983;
  assign n30985 = ~n35576 & ~n30984;
  assign n30986 = ~n29791 & n35576;
  assign n30987 = ~n35574 & n30986;
  assign n30988 = n35576 & n30984;
  assign n30989 = ~n30530 & n30987;
  assign n30990 = ~n30985 & ~n35725;
  assign n30991 = n14866 & n30990;
  assign n30992 = ~n14866 & ~n30990;
  assign n30993 = ~n29774 & ~n29776;
  assign n30994 = ~n30530 & n30993;
  assign n30995 = ~n35573 & ~n30994;
  assign n30996 = ~n29776 & n35573;
  assign n30997 = ~n29774 & n30996;
  assign n30998 = n35573 & n30994;
  assign n30999 = ~n30530 & n30997;
  assign n31000 = ~n30995 & ~n35726;
  assign n31001 = n15586 & n31000;
  assign n31002 = ~n15586 & ~n31000;
  assign n31003 = ~n29760 & ~n35571;
  assign n31004 = ~n29760 & ~n30530;
  assign n31005 = ~n35571 & n31004;
  assign n31006 = ~n30530 & n31003;
  assign n31007 = n29768 & ~n35727;
  assign n31008 = n29772 & n31004;
  assign n31009 = ~n29768 & ~n35727;
  assign n31010 = ~n29760 & n29768;
  assign n31011 = ~n35571 & n31010;
  assign n31012 = ~n30530 & n31011;
  assign n31013 = ~n31009 & ~n31012;
  assign n31014 = ~n31007 & ~n31008;
  assign n31015 = n16248 & n35728;
  assign n31016 = ~n16248 & ~n35728;
  assign n31017 = ~n29743 & ~n29745;
  assign n31018 = ~n30530 & n31017;
  assign n31019 = ~n35569 & ~n31018;
  assign n31020 = ~n29745 & n35569;
  assign n31021 = ~n29743 & n31020;
  assign n31022 = n35569 & n31018;
  assign n31023 = ~n30530 & n31021;
  assign n31024 = ~n31019 & ~n35729;
  assign n31025 = n17001 & n31024;
  assign n31026 = ~n17001 & ~n31024;
  assign n31027 = ~n29724 & ~n35564;
  assign n31028 = ~n30530 & n31027;
  assign n31029 = ~n35567 & ~n31028;
  assign n31030 = ~n29724 & n35567;
  assign n31031 = ~n35564 & n31030;
  assign n31032 = n35567 & n31028;
  assign n31033 = ~n30530 & n31031;
  assign n31034 = ~n31029 & ~n35730;
  assign n31035 = n17690 & n31034;
  assign n31036 = ~n17690 & ~n31034;
  assign n31037 = ~n29707 & ~n29709;
  assign n31038 = ~n30530 & n31037;
  assign n31039 = ~n35563 & ~n31038;
  assign n31040 = ~n29709 & n35563;
  assign n31041 = ~n29707 & n31040;
  assign n31042 = n35563 & n31038;
  assign n31043 = ~n30530 & n31041;
  assign n31044 = ~n31039 & ~n35731;
  assign n31045 = n18472 & n31044;
  assign n31046 = ~n18472 & ~n31044;
  assign n31047 = ~n29690 & ~n35559;
  assign n31048 = ~n29690 & ~n30530;
  assign n31049 = ~n35559 & n31048;
  assign n31050 = ~n30530 & n31047;
  assign n31051 = n35561 & ~n35732;
  assign n31052 = n29705 & n31048;
  assign n31053 = ~n35561 & n35732;
  assign n31054 = ~n35561 & ~n35732;
  assign n31055 = ~n29690 & n35561;
  assign n31056 = ~n35559 & n31055;
  assign n31057 = ~n30530 & n31056;
  assign n31058 = ~n31054 & ~n31057;
  assign n31059 = ~n31051 & ~n35733;
  assign n31060 = n19190 & n35734;
  assign n31061 = ~n19190 & ~n35734;
  assign n31062 = ~n29673 & ~n29675;
  assign n31063 = ~n30530 & n31062;
  assign n31064 = ~n35558 & ~n31063;
  assign n31065 = ~n29675 & n35558;
  assign n31066 = ~n29673 & n31065;
  assign n31067 = n35558 & n31063;
  assign n31068 = ~n30530 & n31066;
  assign n31069 = ~n31064 & ~n35735;
  assign n31070 = n20011 & n31069;
  assign n31071 = ~n20011 & ~n31069;
  assign n31072 = ~n29657 & ~n35555;
  assign n31073 = ~n30530 & n31072;
  assign n31074 = ~n35556 & n31073;
  assign n31075 = n35556 & ~n31073;
  assign n31076 = ~n35556 & ~n31073;
  assign n31077 = ~n29657 & n35556;
  assign n31078 = ~n35555 & n31077;
  assign n31079 = n35556 & n31073;
  assign n31080 = ~n30530 & n31078;
  assign n31081 = ~n31076 & ~n35736;
  assign n31082 = ~n31074 & ~n31075;
  assign n31083 = n20762 & n35737;
  assign n31084 = ~n20762 & ~n35737;
  assign n31085 = ~n29640 & ~n29642;
  assign n31086 = ~n30530 & n31085;
  assign n31087 = ~n35554 & ~n31086;
  assign n31088 = ~n29642 & n35554;
  assign n31089 = ~n29640 & n31088;
  assign n31090 = n35554 & n31086;
  assign n31091 = ~n30530 & n31089;
  assign n31092 = ~n31087 & ~n35738;
  assign n31093 = n21612 & n31092;
  assign n31094 = ~n21612 & ~n31092;
  assign n31095 = ~n29624 & ~n35551;
  assign n31096 = ~n30530 & n31095;
  assign n31097 = ~n35552 & n31096;
  assign n31098 = n35552 & ~n31096;
  assign n31099 = ~n35552 & ~n31096;
  assign n31100 = ~n29624 & n35552;
  assign n31101 = ~n35551 & n31100;
  assign n31102 = ~n30530 & n31101;
  assign n31103 = ~n31099 & ~n31102;
  assign n31104 = ~n31097 & ~n31098;
  assign n31105 = n22386 & n35739;
  assign n31106 = ~n22386 & ~n35739;
  assign n31107 = ~n29607 & ~n29609;
  assign n31108 = ~n30530 & n31107;
  assign n31109 = ~n35550 & ~n31108;
  assign n31110 = ~n29609 & n35550;
  assign n31111 = ~n29607 & n31110;
  assign n31112 = n35550 & n31108;
  assign n31113 = ~n30530 & n31111;
  assign n31114 = ~n31109 & ~n35740;
  assign n31115 = n23269 & n31114;
  assign n31116 = ~n23269 & ~n31114;
  assign n31117 = ~n29590 & ~n35546;
  assign n31118 = ~n30530 & n31117;
  assign n31119 = ~n35548 & ~n31118;
  assign n31120 = n35548 & n31118;
  assign n31121 = n35548 & ~n31118;
  assign n31122 = ~n29590 & ~n35548;
  assign n31123 = ~n35546 & n31122;
  assign n31124 = ~n30530 & n31123;
  assign n31125 = ~n31121 & ~n31124;
  assign n31126 = ~n31119 & ~n31120;
  assign n31127 = n24076 & n35741;
  assign n31128 = ~n24076 & ~n35741;
  assign n31129 = ~n29573 & ~n29575;
  assign n31130 = ~n30530 & n31129;
  assign n31131 = ~n35545 & ~n31130;
  assign n31132 = ~n29575 & n35545;
  assign n31133 = ~n29573 & n31132;
  assign n31134 = n35545 & n31130;
  assign n31135 = ~n30530 & n31133;
  assign n31136 = ~n31131 & ~n35742;
  assign n31137 = n24994 & n31136;
  assign n31138 = ~n24994 & ~n31136;
  assign n31139 = ~n29560 & ~n35542;
  assign n31140 = ~n30530 & n31139;
  assign n31141 = ~n29570 & ~n31140;
  assign n31142 = ~n29560 & n29570;
  assign n31143 = ~n35542 & n31142;
  assign n31144 = n29570 & n31140;
  assign n31145 = ~n30530 & n31143;
  assign n31146 = n29570 & ~n31140;
  assign n31147 = ~n29570 & n31140;
  assign n31148 = ~n31146 & ~n31147;
  assign n31149 = ~n31141 & ~n35743;
  assign n31150 = n25830 & ~n35744;
  assign n31151 = ~n25830 & n35744;
  assign n31152 = ~n29545 & ~n29547;
  assign n31153 = ~n30530 & n31152;
  assign n31154 = ~n29557 & ~n31153;
  assign n31155 = ~n29547 & n29557;
  assign n31156 = ~n29545 & n31155;
  assign n31157 = n29557 & n31153;
  assign n31158 = ~n30530 & n31156;
  assign n31159 = ~n31154 & ~n35745;
  assign n31160 = n26781 & n31159;
  assign n31161 = ~pi0  & ~pi1 ;
  assign n31162 = ~pi2  & ~n31161;
  assign n31163 = pi2  & ~n30528;
  assign n31164 = ~n35673 & n31163;
  assign n31165 = pi2  & n30530;
  assign n31166 = ~n30522 & n31164;
  assign n31167 = ~n31162 & ~n35746;
  assign n31168 = ~pi2  & ~n30530;
  assign n31169 = ~pi3  & n31168;
  assign n31170 = n29526 & ~n30530;
  assign n31171 = pi3  & ~n31168;
  assign n31172 = ~n35747 & ~n31171;
  assign n31173 = ~n31167 & ~n31172;
  assign n31174 = n31167 & ~n35747;
  assign n31175 = n31167 & n31172;
  assign n31176 = ~n31171 & n31174;
  assign n31177 = n29514 & ~n35748;
  assign n31178 = ~n29514 & ~n31173;
  assign n31179 = ~n35748 & ~n31178;
  assign n31180 = n29514 & ~n31167;
  assign n31181 = ~n29514 & n31167;
  assign n31182 = ~n31172 & ~n31181;
  assign n31183 = ~n31180 & ~n31182;
  assign n31184 = ~n31173 & ~n31177;
  assign n31185 = ~n28625 & ~n35749;
  assign n31186 = ~n29514 & ~n30528;
  assign n31187 = ~n35673 & n31186;
  assign n31188 = ~n29514 & n30530;
  assign n31189 = ~n30522 & n31187;
  assign n31190 = ~n35747 & ~n35750;
  assign n31191 = pi4  & ~n31190;
  assign n31192 = ~pi4  & ~n35750;
  assign n31193 = ~pi4  & n31190;
  assign n31194 = ~n35747 & n31192;
  assign n31195 = ~n31191 & ~n35751;
  assign n31196 = ~n31185 & n31195;
  assign n31197 = ~n29532 & ~n35539;
  assign n31198 = ~n30530 & n31197;
  assign n31199 = n29537 & ~n31198;
  assign n31200 = ~n29537 & n31197;
  assign n31201 = ~n29537 & n31198;
  assign n31202 = ~n30530 & n31200;
  assign n31203 = ~n31199 & ~n35752;
  assign n31204 = n27648 & n31203;
  assign n31205 = n28625 & n35749;
  assign n31206 = ~n31204 & ~n31205;
  assign n31207 = ~n31196 & n31206;
  assign n31208 = ~n27648 & ~n31203;
  assign n31209 = ~n26781 & ~n31159;
  assign n31210 = ~n31208 & ~n31209;
  assign n31211 = ~n31207 & n31210;
  assign n31212 = ~n35749 & ~n31195;
  assign n31213 = n28625 & ~n31212;
  assign n31214 = n35749 & n31195;
  assign n31215 = ~n31213 & ~n31214;
  assign n31216 = ~n31196 & ~n31205;
  assign n31217 = n31203 & ~n35753;
  assign n31218 = ~n31203 & ~n31214;
  assign n31219 = ~n31213 & n31218;
  assign n31220 = n27648 & ~n31219;
  assign n31221 = ~n31159 & ~n31220;
  assign n31222 = ~n31217 & n31221;
  assign n31223 = n26781 & ~n31222;
  assign n31224 = ~n31208 & ~n35753;
  assign n31225 = ~n31217 & ~n31220;
  assign n31226 = ~n31204 & ~n31224;
  assign n31227 = n31159 & ~n35754;
  assign n31228 = ~n31223 & ~n31227;
  assign n31229 = ~n26781 & n35754;
  assign n31230 = n31159 & ~n31229;
  assign n31231 = n26781 & ~n35754;
  assign n31232 = ~n31230 & ~n31231;
  assign n31233 = ~n31160 & ~n31211;
  assign n31234 = ~n31151 & ~n35755;
  assign n31235 = ~n35744 & ~n35755;
  assign n31236 = n35744 & ~n31227;
  assign n31237 = ~n31223 & n31236;
  assign n31238 = n25830 & ~n31237;
  assign n31239 = ~n31235 & ~n31238;
  assign n31240 = ~n31150 & ~n31234;
  assign n31241 = ~n31138 & ~n35756;
  assign n31242 = ~n31136 & ~n31238;
  assign n31243 = ~n31235 & n31242;
  assign n31244 = n24994 & ~n31243;
  assign n31245 = n31136 & ~n35756;
  assign n31246 = ~n31244 & ~n31245;
  assign n31247 = ~n24994 & n35756;
  assign n31248 = n31136 & ~n31247;
  assign n31249 = n24994 & ~n35756;
  assign n31250 = ~n31248 & ~n31249;
  assign n31251 = ~n31137 & ~n31241;
  assign n31252 = ~n31128 & ~n35757;
  assign n31253 = n35741 & ~n35757;
  assign n31254 = ~n35741 & ~n31245;
  assign n31255 = ~n31244 & n31254;
  assign n31256 = n24076 & ~n31255;
  assign n31257 = ~n31253 & ~n31256;
  assign n31258 = ~n31127 & ~n31252;
  assign n31259 = ~n31116 & ~n35758;
  assign n31260 = ~n31114 & ~n31256;
  assign n31261 = ~n31253 & n31260;
  assign n31262 = n23269 & ~n31261;
  assign n31263 = n31114 & ~n35758;
  assign n31264 = ~n31262 & ~n31263;
  assign n31265 = ~n23269 & n35758;
  assign n31266 = n31114 & ~n31265;
  assign n31267 = n23269 & ~n35758;
  assign n31268 = ~n31266 & ~n31267;
  assign n31269 = ~n31115 & ~n31259;
  assign n31270 = ~n31106 & ~n35759;
  assign n31271 = n35739 & ~n35759;
  assign n31272 = ~n35739 & ~n31263;
  assign n31273 = ~n31262 & n31272;
  assign n31274 = n22386 & ~n31273;
  assign n31275 = ~n31271 & ~n31274;
  assign n31276 = ~n31105 & ~n31270;
  assign n31277 = ~n31094 & ~n35760;
  assign n31278 = ~n31092 & ~n31274;
  assign n31279 = ~n31271 & n31278;
  assign n31280 = n21612 & ~n31279;
  assign n31281 = n31092 & ~n35760;
  assign n31282 = ~n31280 & ~n31281;
  assign n31283 = ~n21612 & n35760;
  assign n31284 = n31092 & ~n31283;
  assign n31285 = n21612 & ~n35760;
  assign n31286 = ~n31284 & ~n31285;
  assign n31287 = ~n31093 & ~n31277;
  assign n31288 = ~n31084 & ~n35761;
  assign n31289 = n35737 & ~n35761;
  assign n31290 = ~n35737 & ~n31281;
  assign n31291 = ~n31280 & n31290;
  assign n31292 = n20762 & ~n31291;
  assign n31293 = ~n31289 & ~n31292;
  assign n31294 = ~n31083 & ~n31288;
  assign n31295 = ~n31071 & ~n35762;
  assign n31296 = ~n31069 & ~n31292;
  assign n31297 = ~n31289 & n31296;
  assign n31298 = n20011 & ~n31297;
  assign n31299 = n31069 & ~n35762;
  assign n31300 = ~n31298 & ~n31299;
  assign n31301 = ~n20011 & n35762;
  assign n31302 = n31069 & ~n31301;
  assign n31303 = n20011 & ~n35762;
  assign n31304 = ~n31302 & ~n31303;
  assign n31305 = ~n31070 & ~n31295;
  assign n31306 = ~n31061 & ~n35763;
  assign n31307 = n35734 & ~n35763;
  assign n31308 = ~n35734 & ~n31299;
  assign n31309 = ~n31298 & n31308;
  assign n31310 = n19190 & ~n31309;
  assign n31311 = ~n31307 & ~n31310;
  assign n31312 = ~n31060 & ~n31306;
  assign n31313 = ~n31046 & ~n35764;
  assign n31314 = ~n31044 & ~n31310;
  assign n31315 = ~n31307 & n31314;
  assign n31316 = n18472 & ~n31315;
  assign n31317 = n31044 & ~n35764;
  assign n31318 = ~n31316 & ~n31317;
  assign n31319 = ~n18472 & n35764;
  assign n31320 = n31044 & ~n31319;
  assign n31321 = n18472 & ~n35764;
  assign n31322 = ~n31320 & ~n31321;
  assign n31323 = ~n31045 & ~n31313;
  assign n31324 = ~n31036 & ~n35765;
  assign n31325 = n31034 & ~n35765;
  assign n31326 = ~n31034 & ~n31317;
  assign n31327 = ~n31316 & n31326;
  assign n31328 = n17690 & ~n31327;
  assign n31329 = ~n31325 & ~n31328;
  assign n31330 = ~n31035 & ~n31324;
  assign n31331 = ~n31026 & ~n35766;
  assign n31332 = ~n31024 & ~n31328;
  assign n31333 = ~n31325 & n31332;
  assign n31334 = n17001 & ~n31333;
  assign n31335 = n31024 & ~n35766;
  assign n31336 = ~n31334 & ~n31335;
  assign n31337 = ~n17001 & n35766;
  assign n31338 = n31024 & ~n31337;
  assign n31339 = n17001 & ~n35766;
  assign n31340 = ~n31338 & ~n31339;
  assign n31341 = ~n31025 & ~n31331;
  assign n31342 = ~n31016 & ~n35767;
  assign n31343 = n35728 & ~n35767;
  assign n31344 = ~n35728 & ~n31335;
  assign n31345 = ~n31334 & n31344;
  assign n31346 = n16248 & ~n31345;
  assign n31347 = ~n31343 & ~n31346;
  assign n31348 = ~n31015 & ~n31342;
  assign n31349 = ~n31002 & ~n35768;
  assign n31350 = ~n31000 & ~n31346;
  assign n31351 = ~n31343 & n31350;
  assign n31352 = n15586 & ~n31351;
  assign n31353 = n31000 & ~n35768;
  assign n31354 = ~n31352 & ~n31353;
  assign n31355 = ~n15586 & n35768;
  assign n31356 = n31000 & ~n31355;
  assign n31357 = n15586 & ~n35768;
  assign n31358 = ~n31356 & ~n31357;
  assign n31359 = ~n31001 & ~n31349;
  assign n31360 = ~n30992 & ~n35769;
  assign n31361 = n30990 & ~n35769;
  assign n31362 = ~n30990 & ~n31353;
  assign n31363 = ~n31352 & n31362;
  assign n31364 = n14866 & ~n31363;
  assign n31365 = ~n31361 & ~n31364;
  assign n31366 = ~n30991 & ~n31360;
  assign n31367 = ~n30982 & ~n35770;
  assign n31368 = ~n30980 & ~n31364;
  assign n31369 = ~n31361 & n31368;
  assign n31370 = n14233 & ~n31369;
  assign n31371 = n30980 & ~n35770;
  assign n31372 = ~n31370 & ~n31371;
  assign n31373 = ~n14233 & n35770;
  assign n31374 = n30980 & ~n31373;
  assign n31375 = n14233 & ~n35770;
  assign n31376 = ~n31374 & ~n31375;
  assign n31377 = ~n30981 & ~n31367;
  assign n31378 = ~n30972 & ~n35771;
  assign n31379 = n35723 & ~n35771;
  assign n31380 = ~n35723 & ~n31371;
  assign n31381 = ~n31370 & n31380;
  assign n31382 = n13548 & ~n31381;
  assign n31383 = ~n31379 & ~n31382;
  assign n31384 = ~n30971 & ~n31378;
  assign n31385 = ~n30958 & ~n35772;
  assign n31386 = ~n30956 & ~n31382;
  assign n31387 = ~n31379 & n31386;
  assign n31388 = n12948 & ~n31387;
  assign n31389 = n30956 & ~n35772;
  assign n31390 = ~n31388 & ~n31389;
  assign n31391 = ~n12948 & n35772;
  assign n31392 = n30956 & ~n31391;
  assign n31393 = n12948 & ~n35772;
  assign n31394 = ~n31392 & ~n31393;
  assign n31395 = ~n30957 & ~n31385;
  assign n31396 = ~n30948 & ~n35773;
  assign n31397 = n30946 & ~n35773;
  assign n31398 = ~n30946 & ~n31389;
  assign n31399 = ~n31388 & n31398;
  assign n31400 = n12296 & ~n31399;
  assign n31401 = ~n31397 & ~n31400;
  assign n31402 = ~n30947 & ~n31396;
  assign n31403 = ~n30938 & ~n35774;
  assign n31404 = ~n30936 & ~n31400;
  assign n31405 = ~n31397 & n31404;
  assign n31406 = n11719 & ~n31405;
  assign n31407 = n30936 & ~n35774;
  assign n31408 = ~n31406 & ~n31407;
  assign n31409 = ~n11719 & n35774;
  assign n31410 = n30936 & ~n31409;
  assign n31411 = n11719 & ~n35774;
  assign n31412 = ~n31410 & ~n31411;
  assign n31413 = ~n30937 & ~n31403;
  assign n31414 = ~n30928 & ~n35775;
  assign n31415 = n35718 & ~n35775;
  assign n31416 = ~n35718 & ~n31407;
  assign n31417 = ~n31406 & n31416;
  assign n31418 = n11097 & ~n31417;
  assign n31419 = ~n31415 & ~n31418;
  assign n31420 = ~n30927 & ~n31414;
  assign n31421 = ~n30914 & ~n35776;
  assign n31422 = ~n30912 & ~n31418;
  assign n31423 = ~n31415 & n31422;
  assign n31424 = n10555 & ~n31423;
  assign n31425 = n30912 & ~n35776;
  assign n31426 = ~n31424 & ~n31425;
  assign n31427 = ~n10555 & n35776;
  assign n31428 = n30912 & ~n31427;
  assign n31429 = n10555 & ~n35776;
  assign n31430 = ~n31428 & ~n31429;
  assign n31431 = ~n30913 & ~n31421;
  assign n31432 = ~n30904 & ~n35777;
  assign n31433 = n30902 & ~n35777;
  assign n31434 = ~n30902 & ~n31425;
  assign n31435 = ~n31424 & n31434;
  assign n31436 = n9969 & ~n31435;
  assign n31437 = ~n31433 & ~n31436;
  assign n31438 = ~n30903 & ~n31432;
  assign n31439 = ~n30894 & ~n35778;
  assign n31440 = ~n30892 & ~n31436;
  assign n31441 = ~n31433 & n31440;
  assign n31442 = n9457 & ~n31441;
  assign n31443 = n30892 & ~n35778;
  assign n31444 = ~n31442 & ~n31443;
  assign n31445 = ~n9457 & n35778;
  assign n31446 = n30892 & ~n31445;
  assign n31447 = n9457 & ~n35778;
  assign n31448 = ~n31446 & ~n31447;
  assign n31449 = ~n30893 & ~n31439;
  assign n31450 = ~n30884 & ~n35779;
  assign n31451 = n35713 & ~n35779;
  assign n31452 = ~n35713 & ~n31443;
  assign n31453 = ~n31442 & n31452;
  assign n31454 = n8896 & ~n31453;
  assign n31455 = ~n31451 & ~n31454;
  assign n31456 = ~n30883 & ~n31450;
  assign n31457 = ~n30870 & ~n35780;
  assign n31458 = ~n30868 & ~n31454;
  assign n31459 = ~n31451 & n31458;
  assign n31460 = n8411 & ~n31459;
  assign n31461 = n30868 & ~n35780;
  assign n31462 = ~n31460 & ~n31461;
  assign n31463 = ~n8411 & n35780;
  assign n31464 = n30868 & ~n31463;
  assign n31465 = n8411 & ~n35780;
  assign n31466 = ~n31464 & ~n31465;
  assign n31467 = ~n30869 & ~n31457;
  assign n31468 = ~n30860 & ~n35781;
  assign n31469 = n30858 & ~n35781;
  assign n31470 = ~n30858 & ~n31461;
  assign n31471 = ~n31460 & n31470;
  assign n31472 = n7885 & ~n31471;
  assign n31473 = ~n31469 & ~n31472;
  assign n31474 = ~n30859 & ~n31468;
  assign n31475 = ~n30850 & ~n35782;
  assign n31476 = ~n30848 & ~n31472;
  assign n31477 = ~n31469 & n31476;
  assign n31478 = n7428 & ~n31477;
  assign n31479 = n30848 & ~n35782;
  assign n31480 = ~n31478 & ~n31479;
  assign n31481 = ~n7428 & n35782;
  assign n31482 = n30848 & ~n31481;
  assign n31483 = n7428 & ~n35782;
  assign n31484 = ~n31482 & ~n31483;
  assign n31485 = ~n30849 & ~n31475;
  assign n31486 = ~n30840 & ~n35783;
  assign n31487 = n35708 & ~n35783;
  assign n31488 = ~n35708 & ~n31479;
  assign n31489 = ~n31478 & n31488;
  assign n31490 = n6937 & ~n31489;
  assign n31491 = ~n31487 & ~n31490;
  assign n31492 = ~n30839 & ~n31486;
  assign n31493 = ~n30826 & ~n35784;
  assign n31494 = ~n30824 & ~n31490;
  assign n31495 = ~n31487 & n31494;
  assign n31496 = n6507 & ~n31495;
  assign n31497 = n30824 & ~n35784;
  assign n31498 = ~n31496 & ~n31497;
  assign n31499 = ~n6507 & n35784;
  assign n31500 = n30824 & ~n31499;
  assign n31501 = n6507 & ~n35784;
  assign n31502 = ~n31500 & ~n31501;
  assign n31503 = ~n30825 & ~n31493;
  assign n31504 = ~n30816 & ~n35785;
  assign n31505 = n30814 & ~n35785;
  assign n31506 = ~n30814 & ~n31497;
  assign n31507 = ~n31496 & n31506;
  assign n31508 = n6051 & ~n31507;
  assign n31509 = ~n31505 & ~n31508;
  assign n31510 = ~n30815 & ~n31504;
  assign n31511 = ~n30806 & ~n35786;
  assign n31512 = ~n30804 & ~n31508;
  assign n31513 = ~n31505 & n31512;
  assign n31514 = n5648 & ~n31513;
  assign n31515 = n30804 & ~n35786;
  assign n31516 = ~n31514 & ~n31515;
  assign n31517 = ~n5648 & n35786;
  assign n31518 = n30804 & ~n31517;
  assign n31519 = n5648 & ~n35786;
  assign n31520 = ~n31518 & ~n31519;
  assign n31521 = ~n30805 & ~n31511;
  assign n31522 = ~n30796 & ~n35787;
  assign n31523 = n35703 & ~n35787;
  assign n31524 = ~n35703 & ~n31515;
  assign n31525 = ~n31514 & n31524;
  assign n31526 = n5223 & ~n31525;
  assign n31527 = ~n31523 & ~n31526;
  assign n31528 = ~n30795 & ~n31522;
  assign n31529 = ~n30782 & ~n35788;
  assign n31530 = ~n30780 & ~n31526;
  assign n31531 = ~n31523 & n31530;
  assign n31532 = n4851 & ~n31531;
  assign n31533 = n30780 & ~n35788;
  assign n31534 = ~n31532 & ~n31533;
  assign n31535 = ~n4851 & n35788;
  assign n31536 = n30780 & ~n31535;
  assign n31537 = n4851 & ~n35788;
  assign n31538 = ~n31536 & ~n31537;
  assign n31539 = ~n30781 & ~n31529;
  assign n31540 = ~n30772 & ~n35789;
  assign n31541 = n30770 & ~n35789;
  assign n31542 = ~n30770 & ~n31533;
  assign n31543 = ~n31532 & n31542;
  assign n31544 = n4461 & ~n31543;
  assign n31545 = ~n31541 & ~n31544;
  assign n31546 = ~n30771 & ~n31540;
  assign n31547 = ~n30762 & ~n35790;
  assign n31548 = ~n30760 & ~n31544;
  assign n31549 = ~n31541 & n31548;
  assign n31550 = n4115 & ~n31549;
  assign n31551 = n30760 & ~n35790;
  assign n31552 = ~n31550 & ~n31551;
  assign n31553 = ~n4115 & n35790;
  assign n31554 = n30760 & ~n31553;
  assign n31555 = n4115 & ~n35790;
  assign n31556 = ~n31554 & ~n31555;
  assign n31557 = ~n30761 & ~n31547;
  assign n31558 = ~n30752 & ~n35791;
  assign n31559 = n35698 & ~n35791;
  assign n31560 = ~n35698 & ~n31551;
  assign n31561 = ~n31550 & n31560;
  assign n31562 = n3754 & ~n31561;
  assign n31563 = ~n31559 & ~n31562;
  assign n31564 = ~n30751 & ~n31558;
  assign n31565 = ~n30738 & ~n35792;
  assign n31566 = ~n30736 & ~n31562;
  assign n31567 = ~n31559 & n31566;
  assign n31568 = n3444 & ~n31567;
  assign n31569 = n30736 & ~n35792;
  assign n31570 = ~n31568 & ~n31569;
  assign n31571 = ~n3444 & n35792;
  assign n31572 = n30736 & ~n31571;
  assign n31573 = n3444 & ~n35792;
  assign n31574 = ~n31572 & ~n31573;
  assign n31575 = ~n30737 & ~n31565;
  assign n31576 = ~n30728 & ~n35793;
  assign n31577 = n30726 & ~n35793;
  assign n31578 = ~n30726 & ~n31569;
  assign n31579 = ~n31568 & n31578;
  assign n31580 = n3116 & ~n31579;
  assign n31581 = ~n31577 & ~n31580;
  assign n31582 = ~n30727 & ~n31576;
  assign n31583 = ~n30718 & ~n35794;
  assign n31584 = ~n30716 & ~n31580;
  assign n31585 = ~n31577 & n31584;
  assign n31586 = n2833 & ~n31585;
  assign n31587 = n30716 & ~n35794;
  assign n31588 = ~n31586 & ~n31587;
  assign n31589 = ~n2833 & n35794;
  assign n31590 = n30716 & ~n31589;
  assign n31591 = n2833 & ~n35794;
  assign n31592 = ~n31590 & ~n31591;
  assign n31593 = ~n30717 & ~n31583;
  assign n31594 = ~n30708 & ~n35795;
  assign n31595 = n35693 & ~n35795;
  assign n31596 = ~n35693 & ~n31587;
  assign n31597 = ~n31586 & n31596;
  assign n31598 = n2536 & ~n31597;
  assign n31599 = ~n31595 & ~n31598;
  assign n31600 = ~n30707 & ~n31594;
  assign n31601 = ~n30694 & ~n35796;
  assign n31602 = ~n30692 & ~n31598;
  assign n31603 = ~n31595 & n31602;
  assign n31604 = n2283 & ~n31603;
  assign n31605 = n30692 & ~n35796;
  assign n31606 = ~n31604 & ~n31605;
  assign n31607 = ~n2283 & n35796;
  assign n31608 = n30692 & ~n31607;
  assign n31609 = n2283 & ~n35796;
  assign n31610 = ~n31608 & ~n31609;
  assign n31611 = ~n30693 & ~n31601;
  assign n31612 = ~n30684 & ~n35797;
  assign n31613 = n30682 & ~n35797;
  assign n31614 = ~n30682 & ~n31605;
  assign n31615 = ~n31604 & n31614;
  assign n31616 = n2021 & ~n31615;
  assign n31617 = ~n31613 & ~n31616;
  assign n31618 = ~n30683 & ~n31612;
  assign n31619 = ~n30674 & ~n35798;
  assign n31620 = ~n30672 & ~n31616;
  assign n31621 = ~n31613 & n31620;
  assign n31622 = n1796 & ~n31621;
  assign n31623 = n30672 & ~n35798;
  assign n31624 = ~n31622 & ~n31623;
  assign n31625 = ~n1796 & n35798;
  assign n31626 = n30672 & ~n31625;
  assign n31627 = n1796 & ~n35798;
  assign n31628 = ~n31626 & ~n31627;
  assign n31629 = ~n30673 & ~n31619;
  assign n31630 = ~n30664 & ~n35799;
  assign n31631 = n35688 & ~n35799;
  assign n31632 = ~n35688 & ~n31623;
  assign n31633 = ~n31622 & n31632;
  assign n31634 = n1567 & ~n31633;
  assign n31635 = ~n31631 & ~n31634;
  assign n31636 = ~n30663 & ~n31630;
  assign n31637 = ~n30650 & ~n35800;
  assign n31638 = ~n30648 & ~n31634;
  assign n31639 = ~n31631 & n31638;
  assign n31640 = n1374 & ~n31639;
  assign n31641 = n30648 & ~n35800;
  assign n31642 = ~n31640 & ~n31641;
  assign n31643 = ~n1374 & n35800;
  assign n31644 = n30648 & ~n31643;
  assign n31645 = n1374 & ~n35800;
  assign n31646 = ~n31644 & ~n31645;
  assign n31647 = ~n30649 & ~n31637;
  assign n31648 = ~n30640 & ~n35801;
  assign n31649 = n30638 & ~n35801;
  assign n31650 = ~n30638 & ~n31641;
  assign n31651 = ~n31640 & n31650;
  assign n31652 = n1179 & ~n31651;
  assign n31653 = ~n31649 & ~n31652;
  assign n31654 = ~n30639 & ~n31648;
  assign n31655 = ~n30630 & ~n35802;
  assign n31656 = ~n30628 & ~n31652;
  assign n31657 = ~n31649 & n31656;
  assign n31658 = n1016 & ~n31657;
  assign n31659 = n30628 & ~n35802;
  assign n31660 = ~n31658 & ~n31659;
  assign n31661 = ~n1016 & n35802;
  assign n31662 = n30628 & ~n31661;
  assign n31663 = n1016 & ~n35802;
  assign n31664 = ~n31662 & ~n31663;
  assign n31665 = ~n30629 & ~n31655;
  assign n31666 = ~n30620 & ~n35803;
  assign n31667 = n35683 & ~n35803;
  assign n31668 = ~n35683 & ~n31659;
  assign n31669 = ~n31658 & n31668;
  assign n31670 = n855 & ~n31669;
  assign n31671 = ~n31667 & ~n31670;
  assign n31672 = ~n30619 & ~n31666;
  assign n31673 = ~n30606 & ~n35804;
  assign n31674 = ~n30604 & ~n31670;
  assign n31675 = ~n31667 & n31674;
  assign n31676 = n720 & ~n31675;
  assign n31677 = n30604 & ~n35804;
  assign n31678 = ~n31676 & ~n31677;
  assign n31679 = ~n720 & n35804;
  assign n31680 = n30604 & ~n31679;
  assign n31681 = n720 & ~n35804;
  assign n31682 = ~n31680 & ~n31681;
  assign n31683 = ~n30605 & ~n31673;
  assign n31684 = ~n30596 & ~n35805;
  assign n31685 = n30594 & ~n35805;
  assign n31686 = ~n30594 & ~n31677;
  assign n31687 = ~n31676 & n31686;
  assign n31688 = n592 & ~n31687;
  assign n31689 = ~n31685 & ~n31688;
  assign n31690 = ~n30595 & ~n31684;
  assign n31691 = ~n30586 & ~n35806;
  assign n31692 = ~n30584 & ~n31688;
  assign n31693 = ~n31685 & n31692;
  assign n31694 = n487 & ~n31693;
  assign n31695 = n30584 & ~n35806;
  assign n31696 = ~n31694 & ~n31695;
  assign n31697 = ~n487 & n35806;
  assign n31698 = n30584 & ~n31697;
  assign n31699 = n487 & ~n35806;
  assign n31700 = ~n31698 & ~n31699;
  assign n31701 = ~n30585 & ~n31691;
  assign n31702 = ~n30576 & ~n35807;
  assign n31703 = n35678 & ~n35807;
  assign n31704 = ~n35678 & ~n31695;
  assign n31705 = ~n31694 & n31704;
  assign n31706 = n393 & ~n31705;
  assign n31707 = ~n31703 & ~n31706;
  assign n31708 = ~n30575 & ~n31702;
  assign n31709 = ~n30562 & ~n35808;
  assign n31710 = n321 & n30561;
  assign n31711 = ~n30451 & ~n35664;
  assign n31712 = ~n30530 & n31711;
  assign n31713 = ~n35666 & ~n31712;
  assign n31714 = ~n30451 & n35666;
  assign n31715 = ~n35664 & n31714;
  assign n31716 = n35666 & n31712;
  assign n31717 = ~n30530 & n31715;
  assign n31718 = ~n31713 & ~n35809;
  assign n31719 = n263 & n31718;
  assign n31720 = ~n31710 & ~n31719;
  assign n31721 = ~n31709 & n31720;
  assign n31722 = ~n263 & ~n31718;
  assign n31723 = ~n214 & ~n35675;
  assign n31724 = ~n31722 & ~n31723;
  assign n31725 = ~n31721 & n31724;
  assign n31726 = ~n321 & n35808;
  assign n31727 = n30561 & ~n31726;
  assign n31728 = n321 & ~n35808;
  assign n31729 = ~n30561 & ~n31706;
  assign n31730 = ~n31703 & n31729;
  assign n31731 = n321 & ~n31730;
  assign n31732 = n30561 & ~n35808;
  assign n31733 = ~n31731 & ~n31732;
  assign n31734 = ~n31727 & ~n31728;
  assign n31735 = ~n31722 & ~n35810;
  assign n31736 = n31718 & ~n35810;
  assign n31737 = ~n31718 & ~n31732;
  assign n31738 = ~n31731 & n31737;
  assign n31739 = n263 & ~n31738;
  assign n31740 = ~n31736 & ~n31739;
  assign n31741 = ~n31719 & ~n31735;
  assign n31742 = ~n35675 & ~n31739;
  assign n31743 = ~n31736 & n31742;
  assign n31744 = ~n35675 & n35811;
  assign n31745 = n214 & ~n35812;
  assign n31746 = n35675 & ~n35811;
  assign n31747 = ~n31745 & ~n31746;
  assign n31748 = ~n30553 & ~n31725;
  assign n31749 = ~n30542 & ~n35813;
  assign n31750 = n35674 & ~n35813;
  assign n31751 = ~n35674 & ~n31746;
  assign n31752 = ~n31745 & n31751;
  assign n31753 = n197 & ~n31752;
  assign n31754 = ~n31750 & ~n31753;
  assign n31755 = ~n30541 & ~n31749;
  assign n31756 = ~n30490 & ~n30492;
  assign n31757 = ~n30530 & n31756;
  assign n31758 = ~n35670 & ~n31757;
  assign n31759 = ~n30492 & n35670;
  assign n31760 = ~n30490 & n31759;
  assign n31761 = n35670 & n31757;
  assign n31762 = ~n30530 & n31760;
  assign n31763 = ~n31758 & ~n35815;
  assign n31764 = ~n30506 & ~n30514;
  assign n31765 = ~n30514 & ~n30530;
  assign n31766 = ~n30506 & n31765;
  assign n31767 = ~n30530 & n31764;
  assign n31768 = ~n35673 & ~n35816;
  assign n31769 = ~n31763 & n31768;
  assign n31770 = ~n31753 & n31769;
  assign n31771 = ~n31750 & n31770;
  assign n31772 = n35814 & n31769;
  assign n31773 = n193 & ~n35817;
  assign n31774 = ~n35814 & n31763;
  assign n31775 = n30506 & ~n31765;
  assign n31776 = ~n193 & ~n31764;
  assign n31777 = ~n31775 & n31776;
  assign n31778 = ~n31774 & ~n31777;
  assign n31779 = ~n31773 & n31778;
  assign n31780 = n200 | n201;
  assign n31781 = n222 | ~n223;
  assign n31782 = n224 | n225;
  assign n31783 = n228 | n229;
  assign n31784 = n234 | ~n235;
  assign n31785 = n238 | n239;
  assign n31786 = n243 | n244;
  assign n31787 = n246 | n247;
  assign n31788 = n251 | n252;
  assign n31789 = n260 | n261;
  assign n31790 = n271 | n272;
  assign n31791 = n277 | n278;
  assign n31792 = n284 | n285;
  assign n31793 = n291 | n292;
  assign n31794 = n300 | n301;
  assign n31795 = n309 | n310;
  assign n31796 = n318 | n319;
  assign n31797 = n329 | n330;
  assign n31798 = n335 | n336;
  assign n31799 = n339 | n340;
  assign n31800 = n350 | n351;
  assign n31801 = n354 | n355;
  assign n31802 = n366 | n367;
  assign n31803 = n376 | n377;
  assign n31804 = n386 | n387;
  assign n31805 = n401 | n402;
  assign n31806 = n413 | n414;
  assign n31807 = n426 | n427;
  assign n31808 = n433 | n434;
  assign n31809 = n439 | n440;
  assign n31810 = n449 | n450;
  assign n31811 = n457 | ~n458;
  assign n31812 = n466 | n467;
  assign n31813 = n470 | ~n471;
  assign n31814 = n474 | n475;
  assign n31815 = n481 | n482;
  assign n31816 = n497 | n498;
  assign n31817 = n503 | n504;
  assign n31818 = n507 | n508;
  assign n31819 = n519 | n520;
  assign n31820 = n523 | n524;
  assign n31821 = n534 | n535;
  assign n31822 = n545 | n546;
  assign n31823 = n549 | n550;
  assign n31824 = n561 | n562;
  assign n31825 = n565 | ~n566;
  assign n31826 = n574 | n575;
  assign n31827 = n579 | n580;
  assign n31828 = n586 | n587;
  assign n31829 = n600 | n601;
  assign n31830 = n607 | n608;
  assign n31831 = n613 | n614;
  assign n31832 = n626 | n627;
  assign n31833 = n633 | n634;
  assign n31834 = n639 | n640;
  assign n31835 = n649 | n650;
  assign n31836 = n657 | ~n658;
  assign n31837 = n663 | n664;
  assign n31838 = n670 | n671;
  assign n31839 = n674 | ~n675;
  assign n31840 = n683 | n684;
  assign n31841 = n691 | ~n692;
  assign n31842 = n703 | ~n704;
  assign n31843 = n707 | n708;
  assign n31844 = n714 | n715;
  assign n31845 = n730 | n731;
  assign n31846 = n736 | n737;
  assign n31847 = n740 | n741;
  assign n31848 = n752 | n753;
  assign n31849 = n756 | n757;
  assign n31850 = n768 | n769;
  assign n31851 = n779 | n780;
  assign n31852 = n783 | n784;
  assign n31853 = n795 | n796;
  assign n31854 = n799 | ~n800;
  assign n31855 = n809 | n810;
  assign n31856 = n813 | n814;
  assign n31857 = n828 | ~n829;
  assign n31858 = n837 | n838;
  assign n31859 = n842 | n843;
  assign n31860 = n849 | n850;
  assign n31861 = n863 | n864;
  assign n31862 = n870 | n871;
  assign n31863 = n876 | n877;
  assign n31864 = n889 | n890;
  assign n31865 = n896 | n897;
  assign n31866 = n902 | n903;
  assign n31867 = n912 | n913;
  assign n31868 = n920 | ~n921;
  assign n31869 = n926 | n927;
  assign n31870 = n933 | n934;
  assign n31871 = n937 | ~n938;
  assign n31872 = n946 | n947;
  assign n31873 = n954 | ~n955;
  assign n31874 = n960 | n961;
  assign n31875 = n970 | ~n971;
  assign n31876 = n979 | n980;
  assign n31877 = n987 | ~n988;
  assign n31878 = n999 | ~n1000;
  assign n31879 = n1003 | n1004;
  assign n31880 = n1010 | n1011;
  assign n31881 = n1026 | n1027;
  assign n31882 = n1032 | n1033;
  assign n31883 = n1036 | n1037;
  assign n31884 = n1048 | n1049;
  assign n31885 = n1052 | n1053;
  assign n31886 = n1063 | n1064;
  assign n31887 = n1074 | n1075;
  assign n31888 = n1078 | n1079;
  assign n31889 = n1090 | n1091;
  assign n31890 = n1094 | ~n1095;
  assign n31891 = n1104 | n1105;
  assign n31892 = n1108 | n1109;
  assign n31893 = n1123 | ~n1124;
  assign n31894 = n1133 | n1134;
  assign n31895 = n1137 | n1138;
  assign n31896 = n1152 | ~n1153;
  assign n31897 = n1161 | n1162;
  assign n31898 = n1166 | n1167;
  assign n31899 = n1173 | n1174;
  assign n31900 = n1187 | n1188;
  assign n31901 = n1194 | n1195;
  assign n31902 = n1200 | n1201;
  assign n31903 = n1213 | n1214;
  assign n31904 = n1220 | n1221;
  assign n31905 = n1226 | n1227;
  assign n31906 = n1236 | n1237;
  assign n31907 = n1244 | ~n1245;
  assign n31908 = n1250 | n1251;
  assign n31909 = n1257 | n1258;
  assign n31910 = n1261 | ~n1262;
  assign n31911 = n1270 | n1271;
  assign n31912 = n1278 | ~n1279;
  assign n31913 = n1284 | n1285;
  assign n31914 = n1294 | ~n1295;
  assign n31915 = n1303 | n1304;
  assign n31916 = n1311 | ~n1312;
  assign n31917 = n1317 | n1318;
  assign n31918 = n1327 | ~n1328;
  assign n31919 = n1336 | n1337;
  assign n31920 = n1344 | ~n1345;
  assign n31921 = n1355 | n1356;
  assign n31922 = n1357 | ~n1358;
  assign n31923 = n1361 | n1362;
  assign n31924 = n1368 | n1369;
  assign n31925 = n1384 | n1385;
  assign n31926 = n1390 | n1391;
  assign n31927 = n1394 | n1395;
  assign n31928 = n1406 | n1407;
  assign n31929 = n1410 | n1411;
  assign n31930 = n1421 | n1422;
  assign n31931 = n1432 | n1433;
  assign n31932 = n1436 | n1437;
  assign n31933 = n1448 | n1449;
  assign n31934 = n1452 | ~n1453;
  assign n31935 = n1462 | n1463;
  assign n31936 = n1466 | n1467;
  assign n31937 = n1481 | ~n1482;
  assign n31938 = n1491 | n1492;
  assign n31939 = n1495 | n1496;
  assign n31940 = n1510 | ~n1511;
  assign n31941 = n1520 | n1521;
  assign n31942 = n1524 | n1525;
  assign n31943 = n1536 | n1537;
  assign n31944 = n1540 | ~n1541;
  assign n31945 = n1549 | n1550;
  assign n31946 = n1554 | n1555;
  assign n31947 = n1561 | n1562;
  assign n31948 = n1575 | n1576;
  assign n31949 = n1582 | n1583;
  assign n31950 = n1588 | n1589;
  assign n31951 = n1601 | n1602;
  assign n31952 = n1608 | n1609;
  assign n31953 = n1614 | n1615;
  assign n31954 = n1624 | n1625;
  assign n31955 = n1632 | ~n1633;
  assign n31956 = n1638 | n1639;
  assign n31957 = n1645 | n1646;
  assign n31958 = n1649 | ~n1650;
  assign n31959 = n1658 | n1659;
  assign n31960 = n1666 | ~n1667;
  assign n31961 = n1672 | n1673;
  assign n31962 = n1682 | ~n1683;
  assign n31963 = n1691 | n1692;
  assign n31964 = n1699 | ~n1700;
  assign n31965 = n1705 | n1706;
  assign n31966 = n1715 | ~n1716;
  assign n31967 = n1724 | n1725;
  assign n31968 = n1732 | ~n1733;
  assign n31969 = n1738 | n1739;
  assign n31970 = n1747 | n1748;
  assign n31971 = n1749 | ~n1750;
  assign n31972 = n1758 | n1759;
  assign n31973 = n1766 | ~n1767;
  assign n31974 = n1777 | n1778;
  assign n31975 = n1779 | ~n1780;
  assign n31976 = n1783 | n1784;
  assign n31977 = n1790 | n1791;
  assign n31978 = n1806 | n1807;
  assign n31979 = n1812 | n1813;
  assign n31980 = n1816 | n1817;
  assign n31981 = n1828 | n1829;
  assign n31982 = n1832 | n1833;
  assign n31983 = n1843 | n1844;
  assign n31984 = n1854 | n1855;
  assign n31985 = n1858 | n1859;
  assign n31986 = n1870 | n1871;
  assign n31987 = n1874 | ~n1875;
  assign n31988 = n1884 | n1885;
  assign n31989 = n1888 | n1889;
  assign n31990 = n1903 | ~n1904;
  assign n31991 = n1913 | n1914;
  assign n31992 = n1917 | n1918;
  assign n31993 = n1932 | ~n1933;
  assign n31994 = n1942 | n1943;
  assign n31995 = n1946 | n1947;
  assign n31996 = n1960 | n1961;
  assign n31997 = n1962 | ~n1963;
  assign n31998 = n1972 | n1973;
  assign n31999 = n1976 | n1977;
  assign n32000 = n1985 | n1986;
  assign n32001 = n1988 | n1989;
  assign n32002 = n1994 | ~n1995;
  assign n32003 = n2003 | n2004;
  assign n32004 = n2008 | n2009;
  assign n32005 = n2015 | n2016;
  assign n32006 = n2029 | n2030;
  assign n32007 = n2036 | n2037;
  assign n32008 = n2042 | n2043;
  assign n32009 = n2055 | n2056;
  assign n32010 = n2062 | n2063;
  assign n32011 = n2068 | n2069;
  assign n32012 = n2078 | n2079;
  assign n32013 = n2086 | ~n2087;
  assign n32014 = n2092 | n2093;
  assign n32015 = n2099 | n2100;
  assign n32016 = n2103 | ~n2104;
  assign n32017 = n2112 | n2113;
  assign n32018 = n2120 | ~n2121;
  assign n32019 = n2126 | n2127;
  assign n32020 = n2136 | ~n2137;
  assign n32021 = n2145 | n2146;
  assign n32022 = n2153 | ~n2154;
  assign n32023 = n2159 | n2160;
  assign n32024 = n2169 | ~n2170;
  assign n32025 = n2178 | n2179;
  assign n32026 = n2186 | ~n2187;
  assign n32027 = n2192 | n2193;
  assign n32028 = n2201 | n2202;
  assign n32029 = n2203 | ~n2204;
  assign n32030 = n2212 | n2213;
  assign n32031 = n2220 | ~n2221;
  assign n32032 = n2226 | n2227;
  assign n32033 = n2230 | n2231;
  assign n32034 = n2233 | n2234;
  assign n32035 = n2239 | ~n2240;
  assign n32036 = n2248 | n2249;
  assign n32037 = n2256 | ~n2257;
  assign n32038 = n2265 | n2266;
  assign n32039 = n2270 | n2271;
  assign n32040 = n2277 | n2278;
  assign n32041 = n2293 | n2294;
  assign n32042 = n2299 | n2300;
  assign n32043 = n2303 | n2304;
  assign n32044 = n2315 | n2316;
  assign n32045 = n2319 | n2320;
  assign n32046 = n2331 | n2332;
  assign n32047 = n2342 | n2343;
  assign n32048 = n2346 | n2347;
  assign n32049 = n2358 | n2359;
  assign n32050 = n2362 | ~n2363;
  assign n32051 = n2372 | n2373;
  assign n32052 = n2376 | n2377;
  assign n32053 = n2391 | ~n2392;
  assign n32054 = n2401 | n2402;
  assign n32055 = n2405 | n2406;
  assign n32056 = n2420 | ~n2421;
  assign n32057 = n2430 | n2431;
  assign n32058 = n2434 | n2435;
  assign n32059 = n2448 | n2449;
  assign n32060 = n2450 | ~n2451;
  assign n32061 = n2460 | n2461;
  assign n32062 = n2464 | n2465;
  assign n32063 = n2473 | n2474;
  assign n32064 = n2476 | n2477;
  assign n32065 = n2482 | ~n2483;
  assign n32066 = n2492 | n2493;
  assign n32067 = n2496 | n2497;
  assign n32068 = n2506 | n2507;
  assign n32069 = n2518 | n2519;
  assign n32070 = n2523 | n2524;
  assign n32071 = n2530 | n2531;
  assign n32072 = n2544 | n2545;
  assign n32073 = n2551 | n2552;
  assign n32074 = n2557 | n2558;
  assign n32075 = n2570 | n2571;
  assign n32076 = n2577 | n2578;
  assign n32077 = n2583 | n2584;
  assign n32078 = n2593 | n2594;
  assign n32079 = n2601 | ~n2602;
  assign n32080 = n2607 | n2608;
  assign n32081 = n2614 | n2615;
  assign n32082 = n2618 | ~n2619;
  assign n32083 = n2627 | n2628;
  assign n32084 = n2635 | ~n2636;
  assign n32085 = n2641 | n2642;
  assign n32086 = n2651 | ~n2652;
  assign n32087 = n2660 | n2661;
  assign n32088 = n2668 | ~n2669;
  assign n32089 = n2674 | n2675;
  assign n32090 = n2684 | ~n2685;
  assign n32091 = n2693 | n2694;
  assign n32092 = n2701 | ~n2702;
  assign n32093 = n2707 | n2708;
  assign n32094 = n2716 | n2717;
  assign n32095 = n2718 | ~n2719;
  assign n32096 = n2727 | n2728;
  assign n32097 = n2735 | ~n2736;
  assign n32098 = n2741 | n2742;
  assign n32099 = n2745 | n2746;
  assign n32100 = n2748 | n2749;
  assign n32101 = n2754 | ~n2755;
  assign n32102 = n2763 | n2764;
  assign n32103 = n2771 | ~n2772;
  assign n32104 = n2781 | n2782;
  assign n32105 = n2785 | n2786;
  assign n32106 = n2794 | n2795;
  assign n32107 = n2802 | ~n2803;
  assign n32108 = n2808 | n2809;
  assign n32109 = n2816 | ~n2817;
  assign n32110 = n2820 | n2821;
  assign n32111 = n2827 | n2828;
  assign n32112 = n2843 | n2844;
  assign n32113 = n2849 | n2850;
  assign n32114 = n2853 | n2854;
  assign n32115 = n2865 | n2866;
  assign n32116 = n2869 | n2870;
  assign n32117 = n2880 | n2881;
  assign n32118 = n2891 | n2892;
  assign n32119 = n2895 | n2896;
  assign n32120 = n2907 | n2908;
  assign n32121 = n2911 | ~n2912;
  assign n32122 = n2921 | n2922;
  assign n32123 = n2925 | n2926;
  assign n32124 = n2940 | ~n2941;
  assign n32125 = n2950 | n2951;
  assign n32126 = n2954 | n2955;
  assign n32127 = n2969 | ~n2970;
  assign n32128 = n2979 | n2980;
  assign n32129 = n2983 | n2984;
  assign n32130 = n2997 | n2998;
  assign n32131 = n2999 | ~n3000;
  assign n32132 = n3009 | n3010;
  assign n32133 = n3013 | n3014;
  assign n32134 = n3022 | n3023;
  assign n32135 = n3025 | n3026;
  assign n32136 = n3031 | ~n3032;
  assign n32137 = n3041 | n3042;
  assign n32138 = n3045 | n3046;
  assign n32139 = n3055 | n3056;
  assign n32140 = n3068 | n3069;
  assign n32141 = n3072 | n3073;
  assign n32142 = n3081 | n3082;
  assign n32143 = n3089 | ~n3090;
  assign n32144 = n3098 | n3099;
  assign n32145 = n3103 | n3104;
  assign n32146 = n3110 | n3111;
  assign n32147 = n3124 | n3125;
  assign n32148 = n3131 | n3132;
  assign n32149 = n3137 | n3138;
  assign n32150 = n3150 | n3151;
  assign n32151 = n3157 | n3158;
  assign n32152 = n3163 | n3164;
  assign n32153 = n3173 | n3174;
  assign n32154 = n3181 | ~n3182;
  assign n32155 = n3187 | n3188;
  assign n32156 = n3194 | n3195;
  assign n32157 = n3198 | ~n3199;
  assign n32158 = n3207 | n3208;
  assign n32159 = n3215 | ~n3216;
  assign n32160 = n3221 | n3222;
  assign n32161 = n3231 | ~n3232;
  assign n32162 = n3240 | n3241;
  assign n32163 = n3248 | ~n3249;
  assign n32164 = n3254 | n3255;
  assign n32165 = n3264 | ~n3265;
  assign n32166 = n3273 | n3274;
  assign n32167 = n3281 | ~n3282;
  assign n32168 = n3287 | n3288;
  assign n32169 = n3296 | n3297;
  assign n32170 = n3298 | ~n3299;
  assign n32171 = n3307 | n3308;
  assign n32172 = n3315 | ~n3316;
  assign n32173 = n3321 | n3322;
  assign n32174 = n3325 | n3326;
  assign n32175 = n3328 | n3329;
  assign n32176 = n3334 | ~n3335;
  assign n32177 = n3343 | n3344;
  assign n32178 = n3351 | ~n3352;
  assign n32179 = n3361 | n3362;
  assign n32180 = n3365 | n3366;
  assign n32181 = n3374 | n3375;
  assign n32182 = n3382 | ~n3383;
  assign n32183 = n3388 | n3389;
  assign n32184 = n3392 | n3393;
  assign n32185 = n3400 | ~n3401;
  assign n32186 = n3409 | n3410;
  assign n32187 = n3417 | ~n3418;
  assign n32188 = n3426 | n3427;
  assign n32189 = n3431 | n3432;
  assign n32190 = n3438 | n3439;
  assign n32191 = n3454 | n3455;
  assign n32192 = n3460 | n3461;
  assign n32193 = n3464 | n3465;
  assign n32194 = n3476 | n3477;
  assign n32195 = n3480 | n3481;
  assign n32196 = n3491 | n3492;
  assign n32197 = n3502 | n3503;
  assign n32198 = n3506 | n3507;
  assign n32199 = n3518 | n3519;
  assign n32200 = n3522 | ~n3523;
  assign n32201 = n3532 | n3533;
  assign n32202 = n3536 | n3537;
  assign n32203 = n3551 | ~n3552;
  assign n32204 = n3561 | n3562;
  assign n32205 = n3565 | n3566;
  assign n32206 = n3580 | ~n3581;
  assign n32207 = n3590 | n3591;
  assign n32208 = n3594 | n3595;
  assign n32209 = n3606 | n3607;
  assign n32210 = n3610 | ~n3611;
  assign n32211 = n3620 | n3621;
  assign n32212 = n3624 | n3625;
  assign n32213 = n3633 | n3634;
  assign n32214 = n3636 | n3637;
  assign n32215 = n3642 | ~n3643;
  assign n32216 = n3652 | n3653;
  assign n32217 = n3656 | n3657;
  assign n32218 = n3666 | n3667;
  assign n32219 = n3679 | n3680;
  assign n32220 = n3683 | n3684;
  assign n32221 = n3692 | n3693;
  assign n32222 = n3700 | ~n3701;
  assign n32223 = n3710 | n3711;
  assign n32224 = n3714 | n3715;
  assign n32225 = n3724 | n3725;
  assign n32226 = n3736 | n3737;
  assign n32227 = n3741 | n3742;
  assign n32228 = n3748 | n3749;
  assign n32229 = n3762 | n3763;
  assign n32230 = n3769 | n3770;
  assign n32231 = n3775 | n3776;
  assign n32232 = n3788 | n3789;
  assign n32233 = n3795 | n3796;
  assign n32234 = n3801 | n3802;
  assign n32235 = n3811 | n3812;
  assign n32236 = n3819 | ~n3820;
  assign n32237 = n3825 | n3826;
  assign n32238 = n3832 | n3833;
  assign n32239 = n3836 | ~n3837;
  assign n32240 = n3845 | n3846;
  assign n32241 = n3853 | ~n3854;
  assign n32242 = n3859 | n3860;
  assign n32243 = n3869 | ~n3870;
  assign n32244 = n3878 | n3879;
  assign n32245 = n3886 | ~n3887;
  assign n32246 = n3892 | n3893;
  assign n32247 = n3902 | ~n3903;
  assign n32248 = n3911 | n3912;
  assign n32249 = n3919 | ~n3920;
  assign n32250 = n3925 | n3926;
  assign n32251 = n3934 | n3935;
  assign n32252 = n3936 | ~n3937;
  assign n32253 = n3945 | n3946;
  assign n32254 = n3953 | ~n3954;
  assign n32255 = n3959 | n3960;
  assign n32256 = n3968 | n3969;
  assign n32257 = n3970 | ~n3971;
  assign n32258 = n3979 | n3980;
  assign n32259 = n3987 | ~n3988;
  assign n32260 = n3997 | n3998;
  assign n32261 = n4001 | n4002;
  assign n32262 = n4010 | n4011;
  assign n32263 = n4018 | ~n4019;
  assign n32264 = n4024 | n4025;
  assign n32265 = n4028 | n4029;
  assign n32266 = n4036 | ~n4037;
  assign n32267 = n4045 | n4046;
  assign n32268 = n4053 | ~n4054;
  assign n32269 = n4063 | n4064;
  assign n32270 = n4067 | n4068;
  assign n32271 = n4076 | n4077;
  assign n32272 = n4084 | ~n4085;
  assign n32273 = n4090 | n4091;
  assign n32274 = n4098 | ~n4099;
  assign n32275 = n4102 | n4103;
  assign n32276 = n4109 | n4110;
  assign n32277 = n4125 | n4126;
  assign n32278 = n4131 | n4132;
  assign n32279 = n4135 | n4136;
  assign n32280 = n4147 | n4148;
  assign n32281 = n4151 | n4152;
  assign n32282 = n4162 | n4163;
  assign n32283 = n4173 | n4174;
  assign n32284 = n4177 | n4178;
  assign n32285 = n4189 | n4190;
  assign n32286 = n4193 | ~n4194;
  assign n32287 = n4203 | n4204;
  assign n32288 = n4207 | n4208;
  assign n32289 = n4222 | ~n4223;
  assign n32290 = n4232 | n4233;
  assign n32291 = n4236 | n4237;
  assign n32292 = n4251 | ~n4252;
  assign n32293 = n4261 | n4262;
  assign n32294 = n4265 | n4266;
  assign n32295 = n4279 | n4280;
  assign n32296 = n4281 | ~n4282;
  assign n32297 = n4291 | n4292;
  assign n32298 = n4295 | n4296;
  assign n32299 = n4304 | n4305;
  assign n32300 = n4307 | n4308;
  assign n32301 = n4313 | ~n4314;
  assign n32302 = n4323 | n4324;
  assign n32303 = n4327 | n4328;
  assign n32304 = n4336 | n4337;
  assign n32305 = n4341 | n4342;
  assign n32306 = n4345 | ~n4346;
  assign n32307 = n4355 | n4356;
  assign n32308 = n4359 | n4360;
  assign n32309 = n4368 | n4369;
  assign n32310 = n4376 | ~n4377;
  assign n32311 = n4386 | n4387;
  assign n32312 = n4390 | n4391;
  assign n32313 = n4400 | n4401;
  assign n32314 = n4413 | n4414;
  assign n32315 = n4417 | n4418;
  assign n32316 = n4426 | n4427;
  assign n32317 = n4434 | ~n4435;
  assign n32318 = n4443 | n4444;
  assign n32319 = n4448 | n4449;
  assign n32320 = n4455 | n4456;
  assign n32321 = n4469 | n4470;
  assign n32322 = n4476 | n4477;
  assign n32323 = n4482 | n4483;
  assign n32324 = n4495 | n4496;
  assign n32325 = n4502 | n4503;
  assign n32326 = n4508 | n4509;
  assign n32327 = n4518 | n4519;
  assign n32328 = n4526 | ~n4527;
  assign n32329 = n4532 | n4533;
  assign n32330 = n4539 | n4540;
  assign n32331 = n4543 | ~n4544;
  assign n32332 = n4552 | n4553;
  assign n32333 = n4560 | ~n4561;
  assign n32334 = n4566 | n4567;
  assign n32335 = n4576 | ~n4577;
  assign n32336 = n4585 | n4586;
  assign n32337 = n4593 | ~n4594;
  assign n32338 = n4599 | n4600;
  assign n32339 = n4609 | ~n4610;
  assign n32340 = n4618 | n4619;
  assign n32341 = n4626 | ~n4627;
  assign n32342 = n4632 | n4633;
  assign n32343 = n4641 | n4642;
  assign n32344 = n4643 | ~n4644;
  assign n32345 = n4652 | n4653;
  assign n32346 = n4660 | ~n4661;
  assign n32347 = n4666 | n4667;
  assign n32348 = n4670 | n4671;
  assign n32349 = n4673 | n4674;
  assign n32350 = n4679 | ~n4680;
  assign n32351 = n4688 | n4689;
  assign n32352 = n4696 | ~n4697;
  assign n32353 = n4706 | n4707;
  assign n32354 = n4710 | n4711;
  assign n32355 = n4719 | n4720;
  assign n32356 = n4727 | ~n4728;
  assign n32357 = n4737 | n4738;
  assign n32358 = n4741 | n4742;
  assign n32359 = n4750 | n4751;
  assign n32360 = n4758 | ~n4759;
  assign n32361 = n4768 | n4769;
  assign n32362 = n4772 | n4773;
  assign n32363 = n4781 | n4782;
  assign n32364 = n4789 | ~n4790;
  assign n32365 = n4795 | n4796;
  assign n32366 = n4799 | n4800;
  assign n32367 = n4807 | ~n4808;
  assign n32368 = n4816 | n4817;
  assign n32369 = n4824 | ~n4825;
  assign n32370 = n4833 | n4834;
  assign n32371 = n4838 | n4839;
  assign n32372 = n4845 | n4846;
  assign n32373 = n4861 | n4862;
  assign n32374 = n4867 | n4868;
  assign n32375 = n4871 | n4872;
  assign n32376 = n4883 | n4884;
  assign n32377 = n4887 | n4888;
  assign n32378 = n4898 | n4899;
  assign n32379 = n4909 | n4910;
  assign n32380 = n4913 | n4914;
  assign n32381 = n4925 | n4926;
  assign n32382 = n4929 | ~n4930;
  assign n32383 = n4939 | n4940;
  assign n32384 = n4943 | n4944;
  assign n32385 = n4958 | ~n4959;
  assign n32386 = n4968 | n4969;
  assign n32387 = n4972 | n4973;
  assign n32388 = n4987 | ~n4988;
  assign n32389 = n4997 | n4998;
  assign n32390 = n5001 | n5002;
  assign n32391 = n5015 | n5016;
  assign n32392 = n5017 | ~n5018;
  assign n32393 = n5027 | n5028;
  assign n32394 = n5031 | n5032;
  assign n32395 = n5040 | n5041;
  assign n32396 = n5043 | n5044;
  assign n32397 = n5049 | ~n5050;
  assign n32398 = n5059 | n5060;
  assign n32399 = n5063 | n5064;
  assign n32400 = n5073 | n5074;
  assign n32401 = n5086 | n5087;
  assign n32402 = n5090 | n5091;
  assign n32403 = n5099 | n5100;
  assign n32404 = n5107 | ~n5108;
  assign n32405 = n5117 | n5118;
  assign n32406 = n5121 | n5122;
  assign n32407 = n5130 | n5131;
  assign n32408 = n5138 | ~n5139;
  assign n32409 = n5148 | n5149;
  assign n32410 = n5152 | n5153;
  assign n32411 = n5161 | n5162;
  assign n32412 = n5169 | ~n5170;
  assign n32413 = n5179 | n5180;
  assign n32414 = n5183 | n5184;
  assign n32415 = n5193 | n5194;
  assign n32416 = n5205 | n5206;
  assign n32417 = n5210 | n5211;
  assign n32418 = n5217 | n5218;
  assign n32419 = n5231 | n5232;
  assign n32420 = n5238 | n5239;
  assign n32421 = n5244 | n5245;
  assign n32422 = n5257 | n5258;
  assign n32423 = n5264 | n5265;
  assign n32424 = n5270 | n5271;
  assign n32425 = n5280 | n5281;
  assign n32426 = n5288 | ~n5289;
  assign n32427 = n5294 | n5295;
  assign n32428 = n5301 | n5302;
  assign n32429 = n5305 | ~n5306;
  assign n32430 = n5314 | n5315;
  assign n32431 = n5322 | ~n5323;
  assign n32432 = n5328 | n5329;
  assign n32433 = n5338 | ~n5339;
  assign n32434 = n5347 | n5348;
  assign n32435 = n5355 | ~n5356;
  assign n32436 = n5361 | n5362;
  assign n32437 = n5371 | ~n5372;
  assign n32438 = n5380 | n5381;
  assign n32439 = n5388 | ~n5389;
  assign n32440 = n5394 | n5395;
  assign n32441 = n5403 | n5404;
  assign n32442 = n5405 | ~n5406;
  assign n32443 = n5414 | n5415;
  assign n32444 = n5422 | ~n5423;
  assign n32445 = n5428 | n5429;
  assign n32446 = n5432 | n5433;
  assign n32447 = n5435 | n5436;
  assign n32448 = n5441 | ~n5442;
  assign n32449 = n5450 | n5451;
  assign n32450 = n5458 | ~n5459;
  assign n32451 = n5468 | n5469;
  assign n32452 = n5472 | n5473;
  assign n32453 = n5481 | n5482;
  assign n32454 = n5489 | ~n5490;
  assign n32455 = n5495 | n5496;
  assign n32456 = n5499 | n5500;
  assign n32457 = n5507 | ~n5508;
  assign n32458 = n5516 | n5517;
  assign n32459 = n5524 | ~n5525;
  assign n32460 = n5534 | n5535;
  assign n32461 = n5538 | n5539;
  assign n32462 = n5547 | n5548;
  assign n32463 = n5555 | ~n5556;
  assign n32464 = n5565 | n5566;
  assign n32465 = n5569 | n5570;
  assign n32466 = n5578 | n5579;
  assign n32467 = n5586 | ~n5587;
  assign n32468 = n5596 | n5597;
  assign n32469 = n5600 | n5601;
  assign n32470 = n5609 | n5610;
  assign n32471 = n5617 | ~n5618;
  assign n32472 = n5623 | n5624;
  assign n32473 = n5631 | ~n5632;
  assign n32474 = n5635 | n5636;
  assign n32475 = n5642 | n5643;
  assign n32476 = n5658 | n5659;
  assign n32477 = n5664 | n5665;
  assign n32478 = n5668 | n5669;
  assign n32479 = n5680 | n5681;
  assign n32480 = n5684 | n5685;
  assign n32481 = n5695 | n5696;
  assign n32482 = n5706 | n5707;
  assign n32483 = n5710 | n5711;
  assign n32484 = n5722 | n5723;
  assign n32485 = n5726 | ~n5727;
  assign n32486 = n5736 | n5737;
  assign n32487 = n5740 | n5741;
  assign n32488 = n5755 | ~n5756;
  assign n32489 = n5765 | n5766;
  assign n32490 = n5769 | n5770;
  assign n32491 = n5784 | ~n5785;
  assign n32492 = n5794 | n5795;
  assign n32493 = n5798 | n5799;
  assign n32494 = n5812 | n5813;
  assign n32495 = n5814 | ~n5815;
  assign n32496 = n5824 | n5825;
  assign n32497 = n5828 | n5829;
  assign n32498 = n5837 | n5838;
  assign n32499 = n5840 | n5841;
  assign n32500 = n5846 | ~n5847;
  assign n32501 = n5856 | n5857;
  assign n32502 = n5860 | n5861;
  assign n32503 = n5870 | n5871;
  assign n32504 = n5883 | n5884;
  assign n32505 = n5887 | n5888;
  assign n32506 = n5896 | n5897;
  assign n32507 = n5904 | ~n5905;
  assign n32508 = n5914 | n5915;
  assign n32509 = n5918 | n5919;
  assign n32510 = n5928 | n5929;
  assign n32511 = n5941 | n5942;
  assign n32512 = n5945 | n5946;
  assign n32513 = n5954 | n5955;
  assign n32514 = n5962 | ~n5963;
  assign n32515 = n5972 | n5973;
  assign n32516 = n5976 | n5977;
  assign n32517 = n5985 | n5986;
  assign n32518 = n5993 | ~n5994;
  assign n32519 = n6003 | n6004;
  assign n32520 = n6007 | n6008;
  assign n32521 = n6016 | n6017;
  assign n32522 = n6024 | ~n6025;
  assign n32523 = n6033 | n6034;
  assign n32524 = n6038 | n6039;
  assign n32525 = n6045 | n6046;
  assign n32526 = n6059 | n6060;
  assign n32527 = n6066 | n6067;
  assign n32528 = n6072 | n6073;
  assign n32529 = n6085 | n6086;
  assign n32530 = n6092 | n6093;
  assign n32531 = n6098 | n6099;
  assign n32532 = n6108 | n6109;
  assign n32533 = n6116 | ~n6117;
  assign n32534 = n6122 | n6123;
  assign n32535 = n6129 | n6130;
  assign n32536 = n6133 | ~n6134;
  assign n32537 = n6142 | n6143;
  assign n32538 = n6150 | ~n6151;
  assign n32539 = n6156 | n6157;
  assign n32540 = n6166 | ~n6167;
  assign n32541 = n6175 | n6176;
  assign n32542 = n6183 | ~n6184;
  assign n32543 = n6189 | n6190;
  assign n32544 = n6199 | ~n6200;
  assign n32545 = n6208 | n6209;
  assign n32546 = n6216 | ~n6217;
  assign n32547 = n6222 | n6223;
  assign n32548 = n6231 | n6232;
  assign n32549 = n6233 | ~n6234;
  assign n32550 = n6242 | n6243;
  assign n32551 = n6250 | ~n6251;
  assign n32552 = n6256 | n6257;
  assign n32553 = n6260 | n6261;
  assign n32554 = n6263 | n6264;
  assign n32555 = n6269 | ~n6270;
  assign n32556 = n6278 | n6279;
  assign n32557 = n6286 | ~n6287;
  assign n32558 = n6296 | n6297;
  assign n32559 = n6300 | n6301;
  assign n32560 = n6309 | n6310;
  assign n32561 = n6317 | ~n6318;
  assign n32562 = n6323 | n6324;
  assign n32563 = n6327 | n6328;
  assign n32564 = n6335 | ~n6336;
  assign n32565 = n6344 | n6345;
  assign n32566 = n6352 | ~n6353;
  assign n32567 = n6362 | n6363;
  assign n32568 = n6366 | n6367;
  assign n32569 = n6375 | n6376;
  assign n32570 = n6383 | ~n6384;
  assign n32571 = n6389 | n6390;
  assign n32572 = n6393 | n6394;
  assign n32573 = n6401 | ~n6402;
  assign n32574 = n6410 | n6411;
  assign n32575 = n6418 | ~n6419;
  assign n32576 = n6428 | n6429;
  assign n32577 = n6432 | n6433;
  assign n32578 = n6441 | n6442;
  assign n32579 = n6449 | ~n6450;
  assign n32580 = n6459 | n6460;
  assign n32581 = n6463 | n6464;
  assign n32582 = n6472 | n6473;
  assign n32583 = n6480 | ~n6481;
  assign n32584 = n6489 | n6490;
  assign n32585 = n6494 | n6495;
  assign n32586 = n6501 | n6502;
  assign n32587 = n6517 | n6518;
  assign n32588 = n6523 | n6524;
  assign n32589 = n6527 | n6528;
  assign n32590 = n6539 | n6540;
  assign n32591 = n6543 | n6544;
  assign n32592 = n6554 | n6555;
  assign n32593 = n6565 | n6566;
  assign n32594 = n6569 | n6570;
  assign n32595 = n6581 | n6582;
  assign n32596 = n6585 | ~n6586;
  assign n32597 = n6595 | n6596;
  assign n32598 = n6599 | n6600;
  assign n32599 = n6614 | ~n6615;
  assign n32600 = n6624 | n6625;
  assign n32601 = n6628 | n6629;
  assign n32602 = n6643 | ~n6644;
  assign n32603 = n6653 | n6654;
  assign n32604 = n6657 | n6658;
  assign n32605 = n6671 | n6672;
  assign n32606 = n6673 | ~n6674;
  assign n32607 = n6683 | n6684;
  assign n32608 = n6687 | n6688;
  assign n32609 = n6696 | n6697;
  assign n32610 = n6699 | n6700;
  assign n32611 = n6705 | ~n6706;
  assign n32612 = n6715 | n6716;
  assign n32613 = n6719 | n6720;
  assign n32614 = n6729 | n6730;
  assign n32615 = n6742 | n6743;
  assign n32616 = n6746 | n6747;
  assign n32617 = n6755 | n6756;
  assign n32618 = n6763 | ~n6764;
  assign n32619 = n6773 | n6774;
  assign n32620 = n6777 | n6778;
  assign n32621 = n6787 | n6788;
  assign n32622 = n6800 | n6801;
  assign n32623 = n6804 | n6805;
  assign n32624 = n6813 | n6814;
  assign n32625 = n6821 | ~n6822;
  assign n32626 = n6831 | n6832;
  assign n32627 = n6835 | n6836;
  assign n32628 = n6845 | n6846;
  assign n32629 = n6858 | n6859;
  assign n32630 = n6862 | n6863;
  assign n32631 = n6871 | n6872;
  assign n32632 = n6879 | ~n6880;
  assign n32633 = n6889 | n6890;
  assign n32634 = n6893 | n6894;
  assign n32635 = n6902 | n6903;
  assign n32636 = n6910 | ~n6911;
  assign n32637 = n6919 | n6920;
  assign n32638 = n6924 | n6925;
  assign n32639 = n6931 | n6932;
  assign n32640 = n6945 | n6946;
  assign n32641 = n6952 | n6953;
  assign n32642 = n6958 | n6959;
  assign n32643 = n6971 | n6972;
  assign n32644 = n6978 | n6979;
  assign n32645 = n6984 | n6985;
  assign n32646 = n6994 | n6995;
  assign n32647 = n7002 | ~n7003;
  assign n32648 = n7008 | n7009;
  assign n32649 = n7015 | n7016;
  assign n32650 = n7019 | ~n7020;
  assign n32651 = n7028 | n7029;
  assign n32652 = n7036 | ~n7037;
  assign n32653 = n7042 | n7043;
  assign n32654 = n7052 | ~n7053;
  assign n32655 = n7061 | n7062;
  assign n32656 = n7069 | ~n7070;
  assign n32657 = n7075 | n7076;
  assign n32658 = n7085 | ~n7086;
  assign n32659 = n7094 | n7095;
  assign n32660 = n7102 | ~n7103;
  assign n32661 = n7108 | n7109;
  assign n32662 = n7117 | n7118;
  assign n32663 = n7119 | ~n7120;
  assign n32664 = n7128 | n7129;
  assign n32665 = n7136 | ~n7137;
  assign n32666 = n7142 | n7143;
  assign n32667 = n7146 | n7147;
  assign n32668 = n7149 | n7150;
  assign n32669 = n7155 | ~n7156;
  assign n32670 = n7164 | n7165;
  assign n32671 = n7172 | ~n7173;
  assign n32672 = n7182 | n7183;
  assign n32673 = n7186 | n7187;
  assign n32674 = n7195 | n7196;
  assign n32675 = n7203 | ~n7204;
  assign n32676 = n7209 | n7210;
  assign n32677 = n7213 | n7214;
  assign n32678 = n7221 | ~n7222;
  assign n32679 = n7230 | n7231;
  assign n32680 = n7238 | ~n7239;
  assign n32681 = n7248 | n7249;
  assign n32682 = n7252 | n7253;
  assign n32683 = n7261 | n7262;
  assign n32684 = n7269 | ~n7270;
  assign n32685 = n7275 | n7276;
  assign n32686 = n7279 | n7280;
  assign n32687 = n7287 | ~n7288;
  assign n32688 = n7296 | n7297;
  assign n32689 = n7304 | ~n7305;
  assign n32690 = n7314 | n7315;
  assign n32691 = n7318 | n7319;
  assign n32692 = n7327 | n7328;
  assign n32693 = n7335 | ~n7336;
  assign n32694 = n7341 | n7342;
  assign n32695 = n7345 | n7346;
  assign n32696 = n7353 | ~n7354;
  assign n32697 = n7362 | n7363;
  assign n32698 = n7370 | ~n7371;
  assign n32699 = n7380 | n7381;
  assign n32700 = n7384 | n7385;
  assign n32701 = n7393 | n7394;
  assign n32702 = n7401 | ~n7402;
  assign n32703 = n7410 | n7411;
  assign n32704 = n7415 | n7416;
  assign n32705 = n7422 | n7423;
  assign n32706 = n7438 | n7439;
  assign n32707 = n7444 | n7445;
  assign n32708 = n7448 | n7449;
  assign n32709 = n7460 | n7461;
  assign n32710 = n7464 | n7465;
  assign n32711 = n7475 | n7476;
  assign n32712 = n7486 | n7487;
  assign n32713 = n7490 | n7491;
  assign n32714 = n7502 | n7503;
  assign n32715 = n7506 | ~n7507;
  assign n32716 = n7516 | n7517;
  assign n32717 = n7520 | n7521;
  assign n32718 = n7535 | ~n7536;
  assign n32719 = n7545 | n7546;
  assign n32720 = n7549 | n7550;
  assign n32721 = n7564 | ~n7565;
  assign n32722 = n7574 | n7575;
  assign n32723 = n7578 | n7579;
  assign n32724 = n7592 | n7593;
  assign n32725 = n7594 | ~n7595;
  assign n32726 = n7604 | n7605;
  assign n32727 = n7608 | n7609;
  assign n32728 = n7617 | n7618;
  assign n32729 = n7620 | n7621;
  assign n32730 = n7626 | ~n7627;
  assign n32731 = n7636 | n7637;
  assign n32732 = n7640 | n7641;
  assign n32733 = n7650 | n7651;
  assign n32734 = n7663 | n7664;
  assign n32735 = n7667 | n7668;
  assign n32736 = n7676 | n7677;
  assign n32737 = n7684 | ~n7685;
  assign n32738 = n7694 | n7695;
  assign n32739 = n7698 | n7699;
  assign n32740 = n7708 | n7709;
  assign n32741 = n7721 | n7722;
  assign n32742 = n7725 | n7726;
  assign n32743 = n7734 | n7735;
  assign n32744 = n7742 | ~n7743;
  assign n32745 = n7752 | n7753;
  assign n32746 = n7756 | n7757;
  assign n32747 = n7766 | n7767;
  assign n32748 = n7779 | n7780;
  assign n32749 = n7783 | n7784;
  assign n32750 = n7792 | n7793;
  assign n32751 = n7800 | ~n7801;
  assign n32752 = n7810 | n7811;
  assign n32753 = n7814 | n7815;
  assign n32754 = n7824 | n7825;
  assign n32755 = n7837 | n7838;
  assign n32756 = n7841 | n7842;
  assign n32757 = n7850 | n7851;
  assign n32758 = n7858 | ~n7859;
  assign n32759 = n7867 | n7868;
  assign n32760 = n7872 | n7873;
  assign n32761 = n7879 | n7880;
  assign n32762 = n7893 | n7894;
  assign n32763 = n7900 | n7901;
  assign n32764 = n7906 | n7907;
  assign n32765 = n7919 | n7920;
  assign n32766 = n7926 | n7927;
  assign n32767 = n7932 | n7933;
  assign n32768 = n7942 | n7943;
  assign n32769 = n7950 | ~n7951;
  assign n32770 = n7956 | n7957;
  assign n32771 = n7963 | n7964;
  assign n32772 = n7967 | ~n7968;
  assign n32773 = n7976 | n7977;
  assign n32774 = n7984 | ~n7985;
  assign n32775 = n7990 | n7991;
  assign n32776 = n8000 | ~n8001;
  assign n32777 = n8009 | n8010;
  assign n32778 = n8017 | ~n8018;
  assign n32779 = n8023 | n8024;
  assign n32780 = n8033 | ~n8034;
  assign n32781 = n8042 | n8043;
  assign n32782 = n8050 | ~n8051;
  assign n32783 = n8056 | n8057;
  assign n32784 = n8065 | n8066;
  assign n32785 = n8067 | ~n8068;
  assign n32786 = n8076 | n8077;
  assign n32787 = n8084 | ~n8085;
  assign n32788 = n8090 | n8091;
  assign n32789 = n8094 | n8095;
  assign n32790 = n8097 | n8098;
  assign n32791 = n8103 | ~n8104;
  assign n32792 = n8112 | n8113;
  assign n32793 = n8120 | ~n8121;
  assign n32794 = n8130 | n8131;
  assign n32795 = n8134 | n8135;
  assign n32796 = n8143 | n8144;
  assign n32797 = n8151 | ~n8152;
  assign n32798 = n8157 | n8158;
  assign n32799 = n8161 | n8162;
  assign n32800 = n8169 | ~n8170;
  assign n32801 = n8178 | n8179;
  assign n32802 = n8186 | ~n8187;
  assign n32803 = n8196 | n8197;
  assign n32804 = n8200 | n8201;
  assign n32805 = n8209 | n8210;
  assign n32806 = n8217 | ~n8218;
  assign n32807 = n8223 | n8224;
  assign n32808 = n8227 | n8228;
  assign n32809 = n8235 | ~n8236;
  assign n32810 = n8244 | n8245;
  assign n32811 = n8252 | ~n8253;
  assign n32812 = n8262 | n8263;
  assign n32813 = n8266 | n8267;
  assign n32814 = n8275 | n8276;
  assign n32815 = n8283 | ~n8284;
  assign n32816 = n8289 | n8290;
  assign n32817 = n8293 | n8294;
  assign n32818 = n8301 | ~n8302;
  assign n32819 = n8310 | n8311;
  assign n32820 = n8318 | ~n8319;
  assign n32821 = n8328 | n8329;
  assign n32822 = n8332 | n8333;
  assign n32823 = n8341 | n8342;
  assign n32824 = n8349 | ~n8350;
  assign n32825 = n8355 | n8356;
  assign n32826 = n8359 | n8360;
  assign n32827 = n8367 | ~n8368;
  assign n32828 = n8376 | n8377;
  assign n32829 = n8384 | ~n8385;
  assign n32830 = n8393 | n8394;
  assign n32831 = n8398 | n8399;
  assign n32832 = n8405 | n8406;
  assign n32833 = n8418 | n8419;
  assign n32834 = n8426 | n8427;
  assign n32835 = n8432 | n8433;
  assign n32836 = n8443 | n8444;
  assign n32837 = n8447 | n8448;
  assign n32838 = n8459 | n8460;
  assign n32839 = n8470 | n8471;
  assign n32840 = n8474 | n8475;
  assign n32841 = n8486 | n8487;
  assign n32842 = n8490 | ~n8491;
  assign n32843 = n8500 | n8501;
  assign n32844 = n8504 | n8505;
  assign n32845 = n8519 | ~n8520;
  assign n32846 = n8529 | n8530;
  assign n32847 = n8533 | n8534;
  assign n32848 = n8548 | ~n8549;
  assign n32849 = n8558 | n8559;
  assign n32850 = n8562 | n8563;
  assign n32851 = n8576 | n8577;
  assign n32852 = n8578 | ~n8579;
  assign n32853 = n8588 | n8589;
  assign n32854 = n8592 | n8593;
  assign n32855 = n8601 | n8602;
  assign n32856 = n8604 | n8605;
  assign n32857 = n8610 | ~n8611;
  assign n32858 = n8620 | n8621;
  assign n32859 = n8624 | n8625;
  assign n32860 = n8634 | n8635;
  assign n32861 = n8647 | n8648;
  assign n32862 = n8651 | n8652;
  assign n32863 = n8660 | n8661;
  assign n32864 = n8668 | ~n8669;
  assign n32865 = n8678 | n8679;
  assign n32866 = n8682 | n8683;
  assign n32867 = n8692 | n8693;
  assign n32868 = n8705 | n8706;
  assign n32869 = n8709 | n8710;
  assign n32870 = n8718 | n8719;
  assign n32871 = n8726 | ~n8727;
  assign n32872 = n8736 | n8737;
  assign n32873 = n8740 | n8741;
  assign n32874 = n8750 | n8751;
  assign n32875 = n8763 | n8764;
  assign n32876 = n8767 | n8768;
  assign n32877 = n8776 | n8777;
  assign n32878 = n8784 | ~n8785;
  assign n32879 = n8794 | n8795;
  assign n32880 = n8798 | n8799;
  assign n32881 = n8808 | n8809;
  assign n32882 = n8821 | n8822;
  assign n32883 = n8825 | n8826;
  assign n32884 = n8834 | n8835;
  assign n32885 = n8842 | ~n8843;
  assign n32886 = n8852 | n8853;
  assign n32887 = n8856 | n8857;
  assign n32888 = n8866 | n8867;
  assign n32889 = n8878 | n8879;
  assign n32890 = n8883 | n8884;
  assign n32891 = n8890 | n8891;
  assign n32892 = n8904 | n8905;
  assign n32893 = n8911 | n8912;
  assign n32894 = n8917 | n8918;
  assign n32895 = n8930 | n8931;
  assign n32896 = n8940 | n8941;
  assign n32897 = n8944 | n8945;
  assign n32898 = n8953 | n8954;
  assign n32899 = n8961 | ~n8962;
  assign n32900 = n8967 | n8968;
  assign n32901 = n8974 | n8975;
  assign n32902 = n8978 | ~n8979;
  assign n32903 = n8987 | n8988;
  assign n32904 = n8995 | ~n8996;
  assign n32905 = n9001 | n9002;
  assign n32906 = n9011 | ~n9012;
  assign n32907 = n9020 | n9021;
  assign n32908 = n9028 | ~n9029;
  assign n32909 = n9034 | n9035;
  assign n32910 = n9044 | ~n9045;
  assign n32911 = n9053 | n9054;
  assign n32912 = n9061 | ~n9062;
  assign n32913 = n9067 | n9068;
  assign n32914 = n9076 | n9077;
  assign n32915 = n9078 | ~n9079;
  assign n32916 = n9087 | n9088;
  assign n32917 = n9095 | ~n9096;
  assign n32918 = n9101 | n9102;
  assign n32919 = n9105 | n9106;
  assign n32920 = n9108 | n9109;
  assign n32921 = n9114 | ~n9115;
  assign n32922 = n9123 | n9124;
  assign n32923 = n9131 | ~n9132;
  assign n32924 = n9141 | n9142;
  assign n32925 = n9145 | n9146;
  assign n32926 = n9154 | n9155;
  assign n32927 = n9162 | ~n9163;
  assign n32928 = n9168 | n9169;
  assign n32929 = n9172 | n9173;
  assign n32930 = n9180 | ~n9181;
  assign n32931 = n9189 | n9190;
  assign n32932 = n9197 | ~n9198;
  assign n32933 = n9207 | n9208;
  assign n32934 = n9211 | n9212;
  assign n32935 = n9220 | n9221;
  assign n32936 = n9228 | ~n9229;
  assign n32937 = n9234 | n9235;
  assign n32938 = n9238 | n9239;
  assign n32939 = n9246 | ~n9247;
  assign n32940 = n9255 | n9256;
  assign n32941 = n9263 | ~n9264;
  assign n32942 = n9273 | n9274;
  assign n32943 = n9277 | n9278;
  assign n32944 = n9286 | n9287;
  assign n32945 = n9294 | ~n9295;
  assign n32946 = n9300 | n9301;
  assign n32947 = n9304 | n9305;
  assign n32948 = n9312 | ~n9313;
  assign n32949 = n9321 | n9322;
  assign n32950 = n9329 | ~n9330;
  assign n32951 = n9339 | n9340;
  assign n32952 = n9343 | n9344;
  assign n32953 = n9352 | n9353;
  assign n32954 = n9360 | ~n9361;
  assign n32955 = n9366 | n9367;
  assign n32956 = n9370 | n9371;
  assign n32957 = n9378 | ~n9379;
  assign n32958 = n9387 | n9388;
  assign n32959 = n9395 | ~n9396;
  assign n32960 = n9405 | n9406;
  assign n32961 = n9409 | n9410;
  assign n32962 = n9418 | n9419;
  assign n32963 = n9426 | ~n9427;
  assign n32964 = n9432 | n9433;
  assign n32965 = n9440 | ~n9441;
  assign n32966 = n9444 | n9445;
  assign n32967 = n9451 | n9452;
  assign n32968 = n9463 | n9464;
  assign n32969 = n9467 | n9468;
  assign n32970 = n9475 | n9476;
  assign n32971 = n9485 | n9486;
  assign n32972 = n9492 | n9493;
  assign n32973 = n9500 | n9501;
  assign n32974 = n9510 | n9511;
  assign n32975 = n9518 | n9519;
  assign n32976 = n9528 | n9529;
  assign n32977 = n9542 | n9543;
  assign n32978 = n9546 | n9547;
  assign n32979 = n9561 | ~n9562;
  assign n32980 = n9571 | n9572;
  assign n32981 = n9575 | n9576;
  assign n32982 = n9590 | ~n9591;
  assign n32983 = n9600 | n9601;
  assign n32984 = n9604 | n9605;
  assign n32985 = n9618 | n9619;
  assign n32986 = n9620 | ~n9621;
  assign n32987 = n9630 | n9631;
  assign n32988 = n9634 | n9635;
  assign n32989 = n9643 | n9644;
  assign n32990 = n9646 | n9647;
  assign n32991 = n9652 | ~n9653;
  assign n32992 = n9662 | n9663;
  assign n32993 = n9666 | n9667;
  assign n32994 = n9676 | n9677;
  assign n32995 = n9689 | n9690;
  assign n32996 = n9693 | n9694;
  assign n32997 = n9702 | n9703;
  assign n32998 = n9710 | ~n9711;
  assign n32999 = n9720 | n9721;
  assign n33000 = n9724 | n9725;
  assign n33001 = n9734 | n9735;
  assign n33002 = n9747 | n9748;
  assign n33003 = n9751 | n9752;
  assign n33004 = n9760 | n9761;
  assign n33005 = n9768 | ~n9769;
  assign n33006 = n9778 | n9779;
  assign n33007 = n9782 | n9783;
  assign n33008 = n9792 | n9793;
  assign n33009 = n9805 | n9806;
  assign n33010 = n9809 | n9810;
  assign n33011 = n9818 | n9819;
  assign n33012 = n9826 | ~n9827;
  assign n33013 = n9836 | n9837;
  assign n33014 = n9840 | n9841;
  assign n33015 = n9850 | n9851;
  assign n33016 = n9863 | n9864;
  assign n33017 = n9867 | n9868;
  assign n33018 = n9876 | n9877;
  assign n33019 = n9884 | ~n9885;
  assign n33020 = n9894 | n9895;
  assign n33021 = n9898 | n9899;
  assign n33022 = n9908 | n9909;
  assign n33023 = n9921 | n9922;
  assign n33024 = n9925 | n9926;
  assign n33025 = n9934 | n9935;
  assign n33026 = n9942 | ~n9943;
  assign n33027 = n9951 | n9952;
  assign n33028 = n9956 | n9957;
  assign n33029 = n9963 | n9964;
  assign n33030 = n9977 | n9978;
  assign n33031 = n9984 | n9985;
  assign n33032 = n9990 | n9991;
  assign n33033 = n10003 | n10004;
  assign n33034 = n10010 | n10011;
  assign n33035 = n10016 | n10017;
  assign n33036 = n10026 | n10027;
  assign n33037 = n10034 | ~n10035;
  assign n33038 = n10040 | n10041;
  assign n33039 = n10047 | n10048;
  assign n33040 = n10051 | ~n10052;
  assign n33041 = n10062 | n10063;
  assign n33042 = n10074 | n10075;
  assign n33043 = n10078 | n10079;
  assign n33044 = n10087 | n10088;
  assign n33045 = n10095 | ~n10096;
  assign n33046 = n10101 | n10102;
  assign n33047 = n10111 | ~n10112;
  assign n33048 = n10120 | n10121;
  assign n33049 = n10128 | ~n10129;
  assign n33050 = n10134 | n10135;
  assign n33051 = n10143 | n10144;
  assign n33052 = n10145 | ~n10146;
  assign n33053 = n10154 | n10155;
  assign n33054 = n10162 | ~n10163;
  assign n33055 = n10168 | n10169;
  assign n33056 = n10172 | n10173;
  assign n33057 = n10175 | n10176;
  assign n33058 = n10181 | ~n10182;
  assign n33059 = n10190 | n10191;
  assign n33060 = n10198 | ~n10199;
  assign n33061 = n10208 | n10209;
  assign n33062 = n10212 | n10213;
  assign n33063 = n10221 | n10222;
  assign n33064 = n10229 | ~n10230;
  assign n33065 = n10235 | n10236;
  assign n33066 = n10239 | n10240;
  assign n33067 = n10247 | ~n10248;
  assign n33068 = n10256 | n10257;
  assign n33069 = n10264 | ~n10265;
  assign n33070 = n10274 | n10275;
  assign n33071 = n10278 | n10279;
  assign n33072 = n10287 | n10288;
  assign n33073 = n10295 | ~n10296;
  assign n33074 = n10301 | n10302;
  assign n33075 = n10305 | n10306;
  assign n33076 = n10313 | ~n10314;
  assign n33077 = n10322 | n10323;
  assign n33078 = n10330 | ~n10331;
  assign n33079 = n10340 | n10341;
  assign n33080 = n10344 | n10345;
  assign n33081 = n10353 | n10354;
  assign n33082 = n10361 | ~n10362;
  assign n33083 = n10367 | n10368;
  assign n33084 = n10371 | n10372;
  assign n33085 = n10379 | ~n10380;
  assign n33086 = n10388 | n10389;
  assign n33087 = n10396 | ~n10397;
  assign n33088 = n10406 | n10407;
  assign n33089 = n10410 | n10411;
  assign n33090 = n10419 | n10420;
  assign n33091 = n10427 | ~n10428;
  assign n33092 = n10433 | n10434;
  assign n33093 = n10437 | n10438;
  assign n33094 = n10445 | ~n10446;
  assign n33095 = n10454 | n10455;
  assign n33096 = n10462 | ~n10463;
  assign n33097 = n10472 | n10473;
  assign n33098 = n10476 | n10477;
  assign n33099 = n10485 | n10486;
  assign n33100 = n10493 | ~n10494;
  assign n33101 = n10499 | n10500;
  assign n33102 = n10503 | n10504;
  assign n33103 = n10511 | ~n10512;
  assign n33104 = n10520 | n10521;
  assign n33105 = n10528 | ~n10529;
  assign n33106 = n10537 | n10538;
  assign n33107 = n10542 | n10543;
  assign n33108 = n10549 | n10550;
  assign n33109 = n10561 | n10562;
  assign n33110 = n10569 | n10570;
  assign n33111 = n10577 | n10578;
  assign n33112 = n10581 | n10582;
  assign n33113 = n10589 | n10590;
  assign n33114 = n10599 | n10600;
  assign n33115 = n10606 | n10607;
  assign n33116 = n10614 | n10615;
  assign n33117 = n10624 | n10625;
  assign n33118 = n10632 | n10633;
  assign n33119 = n10643 | n10644;
  assign n33120 = n10647 | ~n10648;
  assign n33121 = n10654 | n10655;
  assign n33122 = n10668 | ~n10669;
  assign n33123 = n10675 | n10676;
  assign n33124 = n10689 | ~n10690;
  assign n33125 = n10701 | n10702;
  assign n33126 = n10705 | n10706;
  assign n33127 = n10717 | n10718;
  assign n33128 = n10721 | ~n10722;
  assign n33129 = n10731 | n10732;
  assign n33130 = n10735 | n10736;
  assign n33131 = n10744 | n10745;
  assign n33132 = n10747 | n10748;
  assign n33133 = n10753 | ~n10754;
  assign n33134 = n10763 | n10764;
  assign n33135 = n10767 | n10768;
  assign n33136 = n10777 | n10778;
  assign n33137 = n10790 | n10791;
  assign n33138 = n10794 | n10795;
  assign n33139 = n10803 | n10804;
  assign n33140 = n10811 | ~n10812;
  assign n33141 = n10821 | n10822;
  assign n33142 = n10825 | n10826;
  assign n33143 = n10835 | n10836;
  assign n33144 = n10848 | n10849;
  assign n33145 = n10852 | n10853;
  assign n33146 = n10861 | n10862;
  assign n33147 = n10869 | ~n10870;
  assign n33148 = n10879 | n10880;
  assign n33149 = n10883 | n10884;
  assign n33150 = n10893 | n10894;
  assign n33151 = n10906 | n10907;
  assign n33152 = n10910 | n10911;
  assign n33153 = n10919 | n10920;
  assign n33154 = n10927 | ~n10928;
  assign n33155 = n10937 | n10938;
  assign n33156 = n10941 | n10942;
  assign n33157 = n10951 | n10952;
  assign n33158 = n10964 | n10965;
  assign n33159 = n10968 | n10969;
  assign n33160 = n10977 | n10978;
  assign n33161 = n10985 | ~n10986;
  assign n33162 = n10995 | n10996;
  assign n33163 = n10999 | n11000;
  assign n33164 = n11009 | n11010;
  assign n33165 = n11022 | n11023;
  assign n33166 = n11026 | n11027;
  assign n33167 = n11035 | n11036;
  assign n33168 = n11043 | ~n11044;
  assign n33169 = n11053 | n11054;
  assign n33170 = n11057 | n11058;
  assign n33171 = n11067 | n11068;
  assign n33172 = n11079 | n11080;
  assign n33173 = n11084 | n11085;
  assign n33174 = n11091 | n11092;
  assign n33175 = n11105 | n11106;
  assign n33176 = n11112 | n11113;
  assign n33177 = n11118 | n11119;
  assign n33178 = n11131 | n11132;
  assign n33179 = n11138 | n11139;
  assign n33180 = n11144 | n11145;
  assign n33181 = n11154 | n11155;
  assign n33182 = n11162 | ~n11163;
  assign n33183 = n11168 | n11169;
  assign n33184 = n11175 | n11176;
  assign n33185 = n11179 | ~n11180;
  assign n33186 = n11188 | n11189;
  assign n33187 = n11196 | ~n11197;
  assign n33188 = n11202 | n11203;
  assign n33189 = n11212 | ~n11213;
  assign n33190 = n11221 | n11222;
  assign n33191 = n11229 | ~n11230;
  assign n33192 = n11235 | n11236;
  assign n33193 = n11245 | ~n11246;
  assign n33194 = n11260 | ~n11261;
  assign n33195 = n11273 | ~n11274;
  assign n33196 = n11276 | n11277;
  assign n33197 = n11285 | n11286;
  assign n33198 = n11293 | ~n11294;
  assign n33199 = n11299 | n11300;
  assign n33200 = n11308 | n11309;
  assign n33201 = n11310 | ~n11311;
  assign n33202 = n11319 | n11320;
  assign n33203 = n11327 | ~n11328;
  assign n33204 = n11337 | n11338;
  assign n33205 = n11341 | n11342;
  assign n33206 = n11350 | n11351;
  assign n33207 = n11358 | ~n11359;
  assign n33208 = n11364 | n11365;
  assign n33209 = n11368 | n11369;
  assign n33210 = n11376 | ~n11377;
  assign n33211 = n11385 | n11386;
  assign n33212 = n11393 | ~n11394;
  assign n33213 = n11403 | n11404;
  assign n33214 = n11407 | n11408;
  assign n33215 = n11416 | n11417;
  assign n33216 = n11424 | ~n11425;
  assign n33217 = n11430 | n11431;
  assign n33218 = n11434 | n11435;
  assign n33219 = n11442 | ~n11443;
  assign n33220 = n11451 | n11452;
  assign n33221 = n11459 | ~n11460;
  assign n33222 = n11469 | n11470;
  assign n33223 = n11473 | n11474;
  assign n33224 = n11482 | n11483;
  assign n33225 = n11490 | ~n11491;
  assign n33226 = n11496 | n11497;
  assign n33227 = n11500 | n11501;
  assign n33228 = n11508 | ~n11509;
  assign n33229 = n11517 | n11518;
  assign n33230 = n11525 | ~n11526;
  assign n33231 = n11535 | n11536;
  assign n33232 = n11539 | n11540;
  assign n33233 = n11548 | n11549;
  assign n33234 = n11556 | ~n11557;
  assign n33235 = n11562 | n11563;
  assign n33236 = n11566 | n11567;
  assign n33237 = n11574 | ~n11575;
  assign n33238 = n11583 | n11584;
  assign n33239 = n11591 | ~n11592;
  assign n33240 = n11601 | n11602;
  assign n33241 = n11605 | n11606;
  assign n33242 = n11614 | n11615;
  assign n33243 = n11622 | ~n11623;
  assign n33244 = n11628 | n11629;
  assign n33245 = n11632 | n11633;
  assign n33246 = n11640 | ~n11641;
  assign n33247 = n11649 | n11650;
  assign n33248 = n11657 | ~n11658;
  assign n33249 = n11667 | n11668;
  assign n33250 = n11671 | n11672;
  assign n33251 = n11680 | n11681;
  assign n33252 = n11688 | ~n11689;
  assign n33253 = n11694 | n11695;
  assign n33254 = n11702 | ~n11703;
  assign n33255 = n11706 | n11707;
  assign n33256 = n11713 | n11714;
  assign n33257 = n11725 | n11726;
  assign n33258 = n11733 | n11734;
  assign n33259 = n11741 | n11742;
  assign n33260 = n11749 | n11750;
  assign n33261 = n11753 | n11754;
  assign n33262 = n11761 | n11762;
  assign n33263 = n11771 | n11772;
  assign n33264 = n11778 | n11779;
  assign n33265 = n11786 | n11787;
  assign n33266 = n11796 | n11797;
  assign n33267 = n11804 | n11805;
  assign n33268 = n11815 | n11816;
  assign n33269 = n11819 | ~n11820;
  assign n33270 = n11826 | n11827;
  assign n33271 = n11840 | ~n11841;
  assign n33272 = n11847 | n11848;
  assign n33273 = n11861 | ~n11862;
  assign n33274 = n11868 | n11869;
  assign n33275 = n11881 | n11882;
  assign n33276 = n11883 | ~n11884;
  assign n33277 = n11890 | n11891;
  assign n33278 = n11900 | ~n11901;
  assign n33279 = n11914 | ~n11915;
  assign n33280 = n11926 | n11927;
  assign n33281 = n11930 | n11931;
  assign n33282 = n11939 | n11940;
  assign n33283 = n11944 | n11945;
  assign n33284 = n11948 | ~n11949;
  assign n33285 = n11958 | n11959;
  assign n33286 = n11962 | n11963;
  assign n33287 = n11971 | n11972;
  assign n33288 = n11979 | ~n11980;
  assign n33289 = n11989 | n11990;
  assign n33290 = n11993 | n11994;
  assign n33291 = n12003 | n12004;
  assign n33292 = n12016 | n12017;
  assign n33293 = n12020 | n12021;
  assign n33294 = n12029 | n12030;
  assign n33295 = n12037 | ~n12038;
  assign n33296 = n12047 | n12048;
  assign n33297 = n12051 | n12052;
  assign n33298 = n12061 | n12062;
  assign n33299 = n12074 | n12075;
  assign n33300 = n12078 | n12079;
  assign n33301 = n12087 | n12088;
  assign n33302 = n12095 | ~n12096;
  assign n33303 = n12105 | n12106;
  assign n33304 = n12109 | n12110;
  assign n33305 = n12119 | n12120;
  assign n33306 = n12132 | n12133;
  assign n33307 = n12136 | n12137;
  assign n33308 = n12145 | n12146;
  assign n33309 = n12153 | ~n12154;
  assign n33310 = n12163 | n12164;
  assign n33311 = n12167 | n12168;
  assign n33312 = n12177 | n12178;
  assign n33313 = n12190 | n12191;
  assign n33314 = n12194 | n12195;
  assign n33315 = n12203 | n12204;
  assign n33316 = n12211 | ~n12212;
  assign n33317 = n12221 | n12222;
  assign n33318 = n12225 | n12226;
  assign n33319 = n12235 | n12236;
  assign n33320 = n12248 | n12249;
  assign n33321 = n12252 | n12253;
  assign n33322 = n12261 | n12262;
  assign n33323 = n12269 | ~n12270;
  assign n33324 = n12278 | n12279;
  assign n33325 = n12283 | n12284;
  assign n33326 = n12290 | n12291;
  assign n33327 = n12304 | n12305;
  assign n33328 = n12311 | n12312;
  assign n33329 = n12317 | n12318;
  assign n33330 = n12330 | n12331;
  assign n33331 = n12337 | n12338;
  assign n33332 = n12343 | n12344;
  assign n33333 = n12353 | n12354;
  assign n33334 = n12361 | ~n12362;
  assign n33335 = n12367 | n12368;
  assign n33336 = n12374 | n12375;
  assign n33337 = n12378 | ~n12379;
  assign n33338 = n12387 | n12388;
  assign n33339 = n12395 | ~n12396;
  assign n33340 = n12401 | n12402;
  assign n33341 = n12411 | ~n12412;
  assign n33342 = n12420 | n12421;
  assign n33343 = n12428 | ~n12429;
  assign n33344 = n12434 | n12435;
  assign n33345 = n12444 | ~n12445;
  assign n33346 = n12453 | n12454;
  assign n33347 = n12461 | ~n12462;
  assign n33348 = n12467 | n12468;
  assign n33349 = n12476 | n12477;
  assign n33350 = n12478 | ~n12479;
  assign n33351 = n12487 | n12488;
  assign n33352 = n12495 | ~n12496;
  assign n33353 = n12501 | n12502;
  assign n33354 = n12505 | n12506;
  assign n33355 = n12508 | n12509;
  assign n33356 = n12514 | ~n12515;
  assign n33357 = n12529 | ~n12530;
  assign n33358 = n12539 | n12540;
  assign n33359 = n12543 | n12544;
  assign n33360 = n12552 | n12553;
  assign n33361 = n12560 | ~n12561;
  assign n33362 = n12570 | n12571;
  assign n33363 = n12574 | n12575;
  assign n33364 = n12583 | n12584;
  assign n33365 = n12591 | ~n12592;
  assign n33366 = n12601 | n12602;
  assign n33367 = n12605 | n12606;
  assign n33368 = n12614 | n12615;
  assign n33369 = n12622 | ~n12623;
  assign n33370 = n12628 | n12629;
  assign n33371 = n12632 | n12633;
  assign n33372 = n12640 | ~n12641;
  assign n33373 = n12649 | n12650;
  assign n33374 = n12657 | ~n12658;
  assign n33375 = n12667 | n12668;
  assign n33376 = n12671 | n12672;
  assign n33377 = n12680 | n12681;
  assign n33378 = n12688 | ~n12689;
  assign n33379 = n12694 | n12695;
  assign n33380 = n12698 | n12699;
  assign n33381 = n12706 | ~n12707;
  assign n33382 = n12715 | n12716;
  assign n33383 = n12723 | ~n12724;
  assign n33384 = n12733 | n12734;
  assign n33385 = n12737 | n12738;
  assign n33386 = n12746 | n12747;
  assign n33387 = n12754 | ~n12755;
  assign n33388 = n12760 | n12761;
  assign n33389 = n12764 | n12765;
  assign n33390 = n12772 | ~n12773;
  assign n33391 = n12781 | n12782;
  assign n33392 = n12789 | ~n12790;
  assign n33393 = n12799 | n12800;
  assign n33394 = n12803 | n12804;
  assign n33395 = n12812 | n12813;
  assign n33396 = n12820 | ~n12821;
  assign n33397 = n12826 | n12827;
  assign n33398 = n12830 | n12831;
  assign n33399 = n12838 | ~n12839;
  assign n33400 = n12847 | n12848;
  assign n33401 = n12855 | ~n12856;
  assign n33402 = n12865 | n12866;
  assign n33403 = n12869 | n12870;
  assign n33404 = n12878 | n12879;
  assign n33405 = n12886 | ~n12887;
  assign n33406 = n12892 | n12893;
  assign n33407 = n12896 | n12897;
  assign n33408 = n12904 | ~n12905;
  assign n33409 = n12913 | n12914;
  assign n33410 = n12921 | ~n12922;
  assign n33411 = n12930 | n12931;
  assign n33412 = n12935 | n12936;
  assign n33413 = n12942 | n12943;
  assign n33414 = n12954 | n12955;
  assign n33415 = n12962 | n12963;
  assign n33416 = n12970 | n12971;
  assign n33417 = n12978 | n12979;
  assign n33418 = n12986 | n12987;
  assign n33419 = n12994 | n12995;
  assign n33420 = n13002 | n13003;
  assign n33421 = n13010 | n13011;
  assign n33422 = n13014 | n13015;
  assign n33423 = n13022 | n13023;
  assign n33424 = n13032 | n13033;
  assign n33425 = n13039 | n13040;
  assign n33426 = n13047 | n13048;
  assign n33427 = n13057 | n13058;
  assign n33428 = n13065 | n13066;
  assign n33429 = n13076 | n13077;
  assign n33430 = n13080 | ~n13081;
  assign n33431 = n13087 | n13088;
  assign n33432 = n13101 | ~n13102;
  assign n33433 = n13108 | n13109;
  assign n33434 = n13122 | ~n13123;
  assign n33435 = n13129 | n13130;
  assign n33436 = n13142 | n13143;
  assign n33437 = n13144 | ~n13145;
  assign n33438 = n13151 | n13152;
  assign n33439 = n13159 | n13160;
  assign n33440 = n13162 | n13163;
  assign n33441 = n13168 | ~n13169;
  assign n33442 = n13175 | n13176;
  assign n33443 = n13186 | n13187;
  assign n33444 = n13196 | n13197;
  assign n33445 = n13210 | n13211;
  assign n33446 = n13214 | n13215;
  assign n33447 = n13223 | n13224;
  assign n33448 = n13231 | ~n13232;
  assign n33449 = n13241 | n13242;
  assign n33450 = n13245 | n13246;
  assign n33451 = n13254 | n13255;
  assign n33452 = n13262 | ~n13263;
  assign n33453 = n13272 | n13273;
  assign n33454 = n13276 | n13277;
  assign n33455 = n13286 | n13287;
  assign n33456 = n13299 | n13300;
  assign n33457 = n13303 | n13304;
  assign n33458 = n13312 | n13313;
  assign n33459 = n13320 | ~n13321;
  assign n33460 = n13330 | n13331;
  assign n33461 = n13334 | n13335;
  assign n33462 = n13344 | n13345;
  assign n33463 = n13357 | n13358;
  assign n33464 = n13361 | n13362;
  assign n33465 = n13370 | n13371;
  assign n33466 = n13378 | ~n13379;
  assign n33467 = n13388 | n13389;
  assign n33468 = n13392 | n13393;
  assign n33469 = n13402 | n13403;
  assign n33470 = n13415 | n13416;
  assign n33471 = n13419 | n13420;
  assign n33472 = n13428 | n13429;
  assign n33473 = n13436 | ~n13437;
  assign n33474 = n13446 | n13447;
  assign n33475 = n13450 | n13451;
  assign n33476 = n13460 | n13461;
  assign n33477 = n13473 | n13474;
  assign n33478 = n13477 | n13478;
  assign n33479 = n13486 | n13487;
  assign n33480 = n13494 | ~n13495;
  assign n33481 = n13504 | n13505;
  assign n33482 = n13508 | n13509;
  assign n33483 = n13518 | n13519;
  assign n33484 = n13530 | n13531;
  assign n33485 = n13535 | n13536;
  assign n33486 = n13542 | n13543;
  assign n33487 = n13556 | n13557;
  assign n33488 = n13563 | n13564;
  assign n33489 = n13569 | n13570;
  assign n33490 = n13582 | n13583;
  assign n33491 = n13589 | n13590;
  assign n33492 = n13595 | n13596;
  assign n33493 = n13605 | n13606;
  assign n33494 = n13613 | ~n13614;
  assign n33495 = n13619 | n13620;
  assign n33496 = n13626 | n13627;
  assign n33497 = n13630 | ~n13631;
  assign n33498 = n13639 | n13640;
  assign n33499 = n13647 | ~n13648;
  assign n33500 = n13653 | n13654;
  assign n33501 = n13663 | ~n13664;
  assign n33502 = n13672 | n13673;
  assign n33503 = n13680 | ~n13681;
  assign n33504 = n13686 | n13687;
  assign n33505 = n13696 | ~n13697;
  assign n33506 = n13705 | n13706;
  assign n33507 = n13713 | ~n13714;
  assign n33508 = n13719 | n13720;
  assign n33509 = n13728 | n13729;
  assign n33510 = n13730 | ~n13731;
  assign n33511 = n13739 | n13740;
  assign n33512 = n13747 | ~n13748;
  assign n33513 = n13753 | n13754;
  assign n33514 = n13757 | n13758;
  assign n33515 = n13760 | n13761;
  assign n33516 = n13766 | ~n13767;
  assign n33517 = n13775 | n13776;
  assign n33518 = n13783 | ~n13784;
  assign n33519 = n13793 | n13794;
  assign n33520 = n13797 | n13798;
  assign n33521 = n13806 | n13807;
  assign n33522 = n13814 | ~n13815;
  assign n33523 = n13820 | n13821;
  assign n33524 = n13824 | n13825;
  assign n33525 = n13832 | ~n13833;
  assign n33526 = n13843 | n13844;
  assign n33527 = n13855 | n13856;
  assign n33528 = n13859 | n13860;
  assign n33529 = n13868 | n13869;
  assign n33530 = n13876 | ~n13877;
  assign n33531 = n13886 | n13887;
  assign n33532 = n13890 | n13891;
  assign n33533 = n13899 | n13900;
  assign n33534 = n13907 | ~n13908;
  assign n33535 = n13917 | n13918;
  assign n33536 = n13921 | n13922;
  assign n33537 = n13930 | n13931;
  assign n33538 = n13938 | ~n13939;
  assign n33539 = n13944 | n13945;
  assign n33540 = n13948 | n13949;
  assign n33541 = n13956 | ~n13957;
  assign n33542 = n13965 | n13966;
  assign n33543 = n13973 | ~n13974;
  assign n33544 = n13983 | n13984;
  assign n33545 = n13987 | n13988;
  assign n33546 = n13996 | n13997;
  assign n33547 = n14004 | ~n14005;
  assign n33548 = n14010 | n14011;
  assign n33549 = n14014 | n14015;
  assign n33550 = n14022 | ~n14023;
  assign n33551 = n14031 | n14032;
  assign n33552 = n14039 | ~n14040;
  assign n33553 = n14049 | n14050;
  assign n33554 = n14053 | n14054;
  assign n33555 = n14062 | n14063;
  assign n33556 = n14070 | ~n14071;
  assign n33557 = n14076 | n14077;
  assign n33558 = n14080 | n14081;
  assign n33559 = n14088 | ~n14089;
  assign n33560 = n14097 | n14098;
  assign n33561 = n14105 | ~n14106;
  assign n33562 = n14115 | n14116;
  assign n33563 = n14119 | n14120;
  assign n33564 = n14128 | n14129;
  assign n33565 = n14136 | ~n14137;
  assign n33566 = n14142 | n14143;
  assign n33567 = n14146 | n14147;
  assign n33568 = n14154 | ~n14155;
  assign n33569 = n14163 | n14164;
  assign n33570 = n14171 | ~n14172;
  assign n33571 = n14181 | n14182;
  assign n33572 = n14185 | n14186;
  assign n33573 = n14194 | n14195;
  assign n33574 = n14202 | ~n14203;
  assign n33575 = n14208 | n14209;
  assign n33576 = n14216 | ~n14217;
  assign n33577 = n14220 | n14221;
  assign n33578 = n14227 | n14228;
  assign n33579 = n14239 | n14240;
  assign n33580 = n14247 | n14248;
  assign n33581 = n14255 | n14256;
  assign n33582 = n14263 | n14264;
  assign n33583 = n14271 | n14272;
  assign n33584 = n14279 | n14280;
  assign n33585 = n14287 | n14288;
  assign n33586 = n14295 | n14296;
  assign n33587 = n14303 | n14304;
  assign n33588 = n14311 | n14312;
  assign n33589 = n14319 | n14320;
  assign n33590 = n14323 | n14324;
  assign n33591 = n14331 | n14332;
  assign n33592 = n14341 | n14342;
  assign n33593 = n14348 | n14349;
  assign n33594 = n14356 | n14357;
  assign n33595 = n14366 | n14367;
  assign n33596 = n14374 | n14375;
  assign n33597 = n14385 | n14386;
  assign n33598 = n14389 | ~n14390;
  assign n33599 = n14396 | n14397;
  assign n33600 = n14410 | ~n14411;
  assign n33601 = n14417 | n14418;
  assign n33602 = n14431 | ~n14432;
  assign n33603 = n14438 | n14439;
  assign n33604 = n14451 | n14452;
  assign n33605 = n14453 | ~n14454;
  assign n33606 = n14460 | n14461;
  assign n33607 = n14468 | n14469;
  assign n33608 = n14471 | n14472;
  assign n33609 = n14477 | ~n14478;
  assign n33610 = n14484 | n14485;
  assign n33611 = n14495 | n14496;
  assign n33612 = n14503 | n14504;
  assign n33613 = n14511 | ~n14512;
  assign n33614 = n14518 | n14519;
  assign n33615 = n14529 | n14530;
  assign n33616 = n14543 | ~n14544;
  assign n33617 = n14555 | n14556;
  assign n33618 = n14559 | n14560;
  assign n33619 = n14568 | n14569;
  assign n33620 = n14576 | ~n14577;
  assign n33621 = n14586 | n14587;
  assign n33622 = n14590 | n14591;
  assign n33623 = n14599 | n14600;
  assign n33624 = n14607 | ~n14608;
  assign n33625 = n14617 | n14618;
  assign n33626 = n14621 | n14622;
  assign n33627 = n14631 | n14632;
  assign n33628 = n14644 | n14645;
  assign n33629 = n14648 | n14649;
  assign n33630 = n14657 | n14658;
  assign n33631 = n14665 | ~n14666;
  assign n33632 = n14675 | n14676;
  assign n33633 = n14679 | n14680;
  assign n33634 = n14689 | n14690;
  assign n33635 = n14702 | n14703;
  assign n33636 = n14706 | n14707;
  assign n33637 = n14715 | n14716;
  assign n33638 = n14723 | ~n14724;
  assign n33639 = n14733 | n14734;
  assign n33640 = n14737 | n14738;
  assign n33641 = n14747 | n14748;
  assign n33642 = n14760 | n14761;
  assign n33643 = n14764 | n14765;
  assign n33644 = n14773 | n14774;
  assign n33645 = n14781 | ~n14782;
  assign n33646 = n14791 | n14792;
  assign n33647 = n14795 | n14796;
  assign n33648 = n14805 | n14806;
  assign n33649 = n14818 | n14819;
  assign n33650 = n14822 | n14823;
  assign n33651 = n14831 | n14832;
  assign n33652 = n14839 | ~n14840;
  assign n33653 = n14848 | n14849;
  assign n33654 = n14853 | n14854;
  assign n33655 = n14860 | n14861;
  assign n33656 = n14874 | n14875;
  assign n33657 = n14881 | n14882;
  assign n33658 = n14887 | n14888;
  assign n33659 = n14900 | n14901;
  assign n33660 = n14907 | n14908;
  assign n33661 = n14913 | n14914;
  assign n33662 = n14923 | n14924;
  assign n33663 = n14931 | ~n14932;
  assign n33664 = n14937 | n14938;
  assign n33665 = n14944 | n14945;
  assign n33666 = n14948 | ~n14949;
  assign n33667 = n14957 | n14958;
  assign n33668 = n14965 | ~n14966;
  assign n33669 = n14971 | n14972;
  assign n33670 = n14981 | ~n14982;
  assign n33671 = n14990 | n14991;
  assign n33672 = n14998 | ~n14999;
  assign n33673 = n15004 | n15005;
  assign n33674 = n15014 | ~n15015;
  assign n33675 = n15023 | n15024;
  assign n33676 = n15031 | ~n15032;
  assign n33677 = n15037 | n15038;
  assign n33678 = n15046 | n15047;
  assign n33679 = n15048 | ~n15049;
  assign n33680 = n15057 | n15058;
  assign n33681 = n15065 | ~n15066;
  assign n33682 = n15071 | n15072;
  assign n33683 = n15075 | n15076;
  assign n33684 = n15078 | n15079;
  assign n33685 = n15084 | ~n15085;
  assign n33686 = n15093 | n15094;
  assign n33687 = n15101 | ~n15102;
  assign n33688 = n15111 | n15112;
  assign n33689 = n15115 | n15116;
  assign n33690 = n15124 | n15125;
  assign n33691 = n15132 | ~n15133;
  assign n33692 = n15138 | n15139;
  assign n33693 = n15142 | n15143;
  assign n33694 = n15150 | ~n15151;
  assign n33695 = n15159 | n15160;
  assign n33696 = n15167 | ~n15168;
  assign n33697 = n15177 | n15178;
  assign n33698 = n15181 | n15182;
  assign n33699 = n15190 | n15191;
  assign n33700 = n15198 | ~n15199;
  assign n33701 = n15204 | n15205;
  assign n33702 = n15208 | n15209;
  assign n33703 = n15216 | ~n15217;
  assign n33704 = n15231 | ~n15232;
  assign n33705 = n15244 | ~n15245;
  assign n33706 = n15247 | n15248;
  assign n33707 = n15256 | n15257;
  assign n33708 = n15264 | ~n15265;
  assign n33709 = n15274 | n15275;
  assign n33710 = n15278 | n15279;
  assign n33711 = n15287 | n15288;
  assign n33712 = n15295 | ~n15296;
  assign n33713 = n15305 | n15306;
  assign n33714 = n15309 | n15310;
  assign n33715 = n15318 | n15319;
  assign n33716 = n15326 | ~n15327;
  assign n33717 = n15332 | n15333;
  assign n33718 = n15336 | n15337;
  assign n33719 = n15344 | ~n15345;
  assign n33720 = n15353 | n15354;
  assign n33721 = n15361 | ~n15362;
  assign n33722 = n15371 | n15372;
  assign n33723 = n15375 | n15376;
  assign n33724 = n15384 | n15385;
  assign n33725 = n15392 | ~n15393;
  assign n33726 = n15398 | n15399;
  assign n33727 = n15402 | n15403;
  assign n33728 = n15410 | ~n15411;
  assign n33729 = n15419 | n15420;
  assign n33730 = n15427 | ~n15428;
  assign n33731 = n15437 | n15438;
  assign n33732 = n15441 | n15442;
  assign n33733 = n15450 | n15451;
  assign n33734 = n15458 | ~n15459;
  assign n33735 = n15464 | n15465;
  assign n33736 = n15468 | n15469;
  assign n33737 = n15476 | ~n15477;
  assign n33738 = n15485 | n15486;
  assign n33739 = n15493 | ~n15494;
  assign n33740 = n15503 | n15504;
  assign n33741 = n15507 | n15508;
  assign n33742 = n15516 | n15517;
  assign n33743 = n15524 | ~n15525;
  assign n33744 = n15530 | n15531;
  assign n33745 = n15534 | n15535;
  assign n33746 = n15542 | ~n15543;
  assign n33747 = n15551 | n15552;
  assign n33748 = n15559 | ~n15560;
  assign n33749 = n15568 | n15569;
  assign n33750 = n15573 | n15574;
  assign n33751 = n15580 | n15581;
  assign n33752 = n15592 | n15593;
  assign n33753 = n15600 | n15601;
  assign n33754 = n15608 | n15609;
  assign n33755 = n15616 | n15617;
  assign n33756 = n15624 | n15625;
  assign n33757 = n15632 | n15633;
  assign n33758 = n15640 | n15641;
  assign n33759 = n15648 | n15649;
  assign n33760 = n15656 | n15657;
  assign n33761 = n15664 | n15665;
  assign n33762 = n15672 | n15673;
  assign n33763 = n15680 | n15681;
  assign n33764 = n15688 | n15689;
  assign n33765 = n15692 | n15693;
  assign n33766 = n15700 | n15701;
  assign n33767 = n15710 | n15711;
  assign n33768 = n15717 | n15718;
  assign n33769 = n15725 | n15726;
  assign n33770 = n15735 | n15736;
  assign n33771 = n15743 | n15744;
  assign n33772 = n15754 | n15755;
  assign n33773 = n15758 | ~n15759;
  assign n33774 = n15765 | n15766;
  assign n33775 = n15779 | ~n15780;
  assign n33776 = n15786 | n15787;
  assign n33777 = n15800 | ~n15801;
  assign n33778 = n15807 | n15808;
  assign n33779 = n15820 | n15821;
  assign n33780 = n15822 | ~n15823;
  assign n33781 = n15829 | n15830;
  assign n33782 = n15837 | n15838;
  assign n33783 = n15840 | n15841;
  assign n33784 = n15846 | ~n15847;
  assign n33785 = n15853 | n15854;
  assign n33786 = n15864 | n15865;
  assign n33787 = n15872 | n15873;
  assign n33788 = n15880 | ~n15881;
  assign n33789 = n15887 | n15888;
  assign n33790 = n15898 | n15899;
  assign n33791 = n15906 | n15907;
  assign n33792 = n15914 | ~n15915;
  assign n33793 = n15921 | n15922;
  assign n33794 = n15932 | n15933;
  assign n33795 = n15942 | ~n15943;
  assign n33796 = n15956 | ~n15957;
  assign n33797 = n15968 | n15969;
  assign n33798 = n15972 | n15973;
  assign n33799 = n15981 | n15982;
  assign n33800 = n15989 | ~n15990;
  assign n33801 = n15999 | n16000;
  assign n33802 = n16003 | n16004;
  assign n33803 = n16012 | n16013;
  assign n33804 = n16020 | ~n16021;
  assign n33805 = n16030 | n16031;
  assign n33806 = n16034 | n16035;
  assign n33807 = n16044 | n16045;
  assign n33808 = n16057 | n16058;
  assign n33809 = n16061 | n16062;
  assign n33810 = n16070 | n16071;
  assign n33811 = n16078 | ~n16079;
  assign n33812 = n16088 | n16089;
  assign n33813 = n16092 | n16093;
  assign n33814 = n16102 | n16103;
  assign n33815 = n16115 | n16116;
  assign n33816 = n16119 | n16120;
  assign n33817 = n16128 | n16129;
  assign n33818 = n16136 | ~n16137;
  assign n33819 = n16146 | n16147;
  assign n33820 = n16150 | n16151;
  assign n33821 = n16160 | n16161;
  assign n33822 = n16173 | n16174;
  assign n33823 = n16177 | n16178;
  assign n33824 = n16186 | n16187;
  assign n33825 = n16194 | ~n16195;
  assign n33826 = n16204 | n16205;
  assign n33827 = n16208 | n16209;
  assign n33828 = n16218 | n16219;
  assign n33829 = n16230 | n16231;
  assign n33830 = n16235 | n16236;
  assign n33831 = n16242 | n16243;
  assign n33832 = n16256 | n16257;
  assign n33833 = n16263 | n16264;
  assign n33834 = n16269 | n16270;
  assign n33835 = n16282 | n16283;
  assign n33836 = n16289 | n16290;
  assign n33837 = n16295 | n16296;
  assign n33838 = n16305 | n16306;
  assign n33839 = n16313 | ~n16314;
  assign n33840 = n16319 | n16320;
  assign n33841 = n16326 | n16327;
  assign n33842 = n16330 | ~n16331;
  assign n33843 = n16339 | n16340;
  assign n33844 = n16347 | ~n16348;
  assign n33845 = n16353 | n16354;
  assign n33846 = n16363 | ~n16364;
  assign n33847 = n16372 | n16373;
  assign n33848 = n16380 | ~n16381;
  assign n33849 = n16386 | n16387;
  assign n33850 = n16396 | ~n16397;
  assign n33851 = n16405 | n16406;
  assign n33852 = n16413 | ~n16414;
  assign n33853 = n16419 | n16420;
  assign n33854 = n16428 | n16429;
  assign n33855 = n16430 | ~n16431;
  assign n33856 = n16439 | n16440;
  assign n33857 = n16447 | ~n16448;
  assign n33858 = n16453 | n16454;
  assign n33859 = n16457 | n16458;
  assign n33860 = n16460 | n16461;
  assign n33861 = n16466 | ~n16467;
  assign n33862 = n16475 | n16476;
  assign n33863 = n16483 | ~n16484;
  assign n33864 = n16493 | n16494;
  assign n33865 = n16497 | n16498;
  assign n33866 = n16506 | n16507;
  assign n33867 = n16514 | ~n16515;
  assign n33868 = n16520 | n16521;
  assign n33869 = n16524 | n16525;
  assign n33870 = n16532 | ~n16533;
  assign n33871 = n16541 | n16542;
  assign n33872 = n16549 | ~n16550;
  assign n33873 = n16559 | n16560;
  assign n33874 = n16563 | n16564;
  assign n33875 = n16572 | n16573;
  assign n33876 = n16580 | ~n16581;
  assign n33877 = n16586 | n16587;
  assign n33878 = n16590 | n16591;
  assign n33879 = n16598 | ~n16599;
  assign n33880 = n16607 | n16608;
  assign n33881 = n16615 | ~n16616;
  assign n33882 = n16625 | n16626;
  assign n33883 = n16629 | n16630;
  assign n33884 = n16638 | n16639;
  assign n33885 = n16646 | ~n16647;
  assign n33886 = n16652 | n16653;
  assign n33887 = n16656 | n16657;
  assign n33888 = n16664 | ~n16665;
  assign n33889 = n16679 | ~n16680;
  assign n33890 = n16689 | n16690;
  assign n33891 = n16693 | n16694;
  assign n33892 = n16702 | n16703;
  assign n33893 = n16710 | ~n16711;
  assign n33894 = n16720 | n16721;
  assign n33895 = n16724 | n16725;
  assign n33896 = n16733 | n16734;
  assign n33897 = n16741 | ~n16742;
  assign n33898 = n16751 | n16752;
  assign n33899 = n16755 | n16756;
  assign n33900 = n16764 | n16765;
  assign n33901 = n16772 | ~n16773;
  assign n33902 = n16778 | n16779;
  assign n33903 = n16782 | n16783;
  assign n33904 = n16790 | ~n16791;
  assign n33905 = n16799 | n16800;
  assign n33906 = n16807 | ~n16808;
  assign n33907 = n16817 | n16818;
  assign n33908 = n16821 | n16822;
  assign n33909 = n16830 | n16831;
  assign n33910 = n16838 | ~n16839;
  assign n33911 = n16844 | n16845;
  assign n33912 = n16848 | n16849;
  assign n33913 = n16856 | ~n16857;
  assign n33914 = n16865 | n16866;
  assign n33915 = n16873 | ~n16874;
  assign n33916 = n16883 | n16884;
  assign n33917 = n16887 | n16888;
  assign n33918 = n16896 | n16897;
  assign n33919 = n16904 | ~n16905;
  assign n33920 = n16910 | n16911;
  assign n33921 = n16914 | n16915;
  assign n33922 = n16922 | ~n16923;
  assign n33923 = n16931 | n16932;
  assign n33924 = n16939 | ~n16940;
  assign n33925 = n16949 | n16950;
  assign n33926 = n16953 | n16954;
  assign n33927 = n16962 | n16963;
  assign n33928 = n16970 | ~n16971;
  assign n33929 = n16976 | n16977;
  assign n33930 = n16984 | ~n16985;
  assign n33931 = n16988 | n16989;
  assign n33932 = n16995 | n16996;
  assign n33933 = n17007 | n17008;
  assign n33934 = n17015 | n17016;
  assign n33935 = n17023 | n17024;
  assign n33936 = n17031 | n17032;
  assign n33937 = n17039 | n17040;
  assign n33938 = n17047 | n17048;
  assign n33939 = n17055 | n17056;
  assign n33940 = n17063 | n17064;
  assign n33941 = n17071 | n17072;
  assign n33942 = n17079 | n17080;
  assign n33943 = n17087 | n17088;
  assign n33944 = n17095 | n17096;
  assign n33945 = n17103 | n17104;
  assign n33946 = n17111 | n17112;
  assign n33947 = n17119 | n17120;
  assign n33948 = n17127 | n17128;
  assign n33949 = n17135 | n17136;
  assign n33950 = n17139 | n17140;
  assign n33951 = n17147 | n17148;
  assign n33952 = n17157 | n17158;
  assign n33953 = n17164 | n17165;
  assign n33954 = n17172 | n17173;
  assign n33955 = n17182 | n17183;
  assign n33956 = n17190 | n17191;
  assign n33957 = n17201 | n17202;
  assign n33958 = n17205 | ~n17206;
  assign n33959 = n17212 | n17213;
  assign n33960 = n17226 | ~n17227;
  assign n33961 = n17233 | n17234;
  assign n33962 = n17247 | ~n17248;
  assign n33963 = n17254 | n17255;
  assign n33964 = n17267 | n17268;
  assign n33965 = n17269 | ~n17270;
  assign n33966 = n17276 | n17277;
  assign n33967 = n17284 | n17285;
  assign n33968 = n17287 | n17288;
  assign n33969 = n17293 | ~n17294;
  assign n33970 = n17300 | n17301;
  assign n33971 = n17311 | n17312;
  assign n33972 = n17319 | n17320;
  assign n33973 = n17327 | ~n17328;
  assign n33974 = n17334 | n17335;
  assign n33975 = n17345 | n17346;
  assign n33976 = n17353 | n17354;
  assign n33977 = n17361 | ~n17362;
  assign n33978 = n17368 | n17369;
  assign n33979 = n17379 | n17380;
  assign n33980 = n17387 | n17388;
  assign n33981 = n17395 | ~n17396;
  assign n33982 = n17402 | n17403;
  assign n33983 = n17413 | n17414;
  assign n33984 = n17423 | n17424;
  assign n33985 = n17437 | n17438;
  assign n33986 = n17441 | n17442;
  assign n33987 = n17450 | n17451;
  assign n33988 = n17458 | ~n17459;
  assign n33989 = n17468 | n17469;
  assign n33990 = n17472 | n17473;
  assign n33991 = n17481 | n17482;
  assign n33992 = n17489 | ~n17490;
  assign n33993 = n17499 | n17500;
  assign n33994 = n17503 | n17504;
  assign n33995 = n17513 | n17514;
  assign n33996 = n17526 | n17527;
  assign n33997 = n17530 | n17531;
  assign n33998 = n17539 | n17540;
  assign n33999 = n17547 | ~n17548;
  assign n34000 = n17557 | n17558;
  assign n34001 = n17561 | n17562;
  assign n34002 = n17571 | n17572;
  assign n34003 = n17584 | n17585;
  assign n34004 = n17588 | n17589;
  assign n34005 = n17597 | n17598;
  assign n34006 = n17605 | ~n17606;
  assign n34007 = n17615 | n17616;
  assign n34008 = n17619 | n17620;
  assign n34009 = n17629 | n17630;
  assign n34010 = n17642 | n17643;
  assign n34011 = n17646 | n17647;
  assign n34012 = n17655 | n17656;
  assign n34013 = n17663 | ~n17664;
  assign n34014 = n17672 | n17673;
  assign n34015 = n17677 | n17678;
  assign n34016 = n17684 | n17685;
  assign n34017 = n17698 | n17699;
  assign n34018 = n17705 | n17706;
  assign n34019 = n17711 | n17712;
  assign n34020 = n17724 | n17725;
  assign n34021 = n17731 | n17732;
  assign n34022 = n17737 | n17738;
  assign n34023 = n17747 | n17748;
  assign n34024 = n17755 | ~n17756;
  assign n34025 = n17761 | n17762;
  assign n34026 = n17768 | n17769;
  assign n34027 = n17772 | ~n17773;
  assign n34028 = n17781 | n17782;
  assign n34029 = n17789 | ~n17790;
  assign n34030 = n17795 | n17796;
  assign n34031 = n17805 | ~n17806;
  assign n34032 = n17814 | n17815;
  assign n34033 = n17822 | ~n17823;
  assign n34034 = n17828 | n17829;
  assign n34035 = n17838 | ~n17839;
  assign n34036 = n17847 | n17848;
  assign n34037 = n17855 | ~n17856;
  assign n34038 = n17861 | n17862;
  assign n34039 = n17870 | n17871;
  assign n34040 = n17872 | ~n17873;
  assign n34041 = n17881 | n17882;
  assign n34042 = n17889 | ~n17890;
  assign n34043 = n17895 | n17896;
  assign n34044 = n17899 | n17900;
  assign n34045 = n17902 | n17903;
  assign n34046 = n17908 | ~n17909;
  assign n34047 = n17917 | n17918;
  assign n34048 = n17925 | ~n17926;
  assign n34049 = n17935 | n17936;
  assign n34050 = n17939 | n17940;
  assign n34051 = n17948 | n17949;
  assign n34052 = n17956 | ~n17957;
  assign n34053 = n17962 | n17963;
  assign n34054 = n17966 | n17967;
  assign n34055 = n17974 | ~n17975;
  assign n34056 = n17983 | n17984;
  assign n34057 = n17991 | ~n17992;
  assign n34058 = n18001 | n18002;
  assign n34059 = n18005 | n18006;
  assign n34060 = n18014 | n18015;
  assign n34061 = n18022 | ~n18023;
  assign n34062 = n18028 | n18029;
  assign n34063 = n18032 | n18033;
  assign n34064 = n18040 | ~n18041;
  assign n34065 = n18049 | n18050;
  assign n34066 = n18057 | ~n18058;
  assign n34067 = n18067 | n18068;
  assign n34068 = n18071 | n18072;
  assign n34069 = n18080 | n18081;
  assign n34070 = n18088 | ~n18089;
  assign n34071 = n18094 | n18095;
  assign n34072 = n18098 | n18099;
  assign n34073 = n18106 | ~n18107;
  assign n34074 = n18115 | n18116;
  assign n34075 = n18123 | ~n18124;
  assign n34076 = n18133 | n18134;
  assign n34077 = n18137 | n18138;
  assign n34078 = n18146 | n18147;
  assign n34079 = n18154 | ~n18155;
  assign n34080 = n18160 | n18161;
  assign n34081 = n18164 | n18165;
  assign n34082 = n18172 | ~n18173;
  assign n34083 = n18183 | n18184;
  assign n34084 = n18195 | n18196;
  assign n34085 = n18199 | n18200;
  assign n34086 = n18208 | n18209;
  assign n34087 = n18216 | ~n18217;
  assign n34088 = n18226 | n18227;
  assign n34089 = n18230 | n18231;
  assign n34090 = n18239 | n18240;
  assign n34091 = n18247 | ~n18248;
  assign n34092 = n18257 | n18258;
  assign n34093 = n18261 | n18262;
  assign n34094 = n18270 | n18271;
  assign n34095 = n18278 | ~n18279;
  assign n34096 = n18284 | n18285;
  assign n34097 = n18288 | n18289;
  assign n34098 = n18296 | ~n18297;
  assign n34099 = n18305 | n18306;
  assign n34100 = n18313 | ~n18314;
  assign n34101 = n18323 | n18324;
  assign n34102 = n18327 | n18328;
  assign n34103 = n18336 | n18337;
  assign n34104 = n18344 | ~n18345;
  assign n34105 = n18350 | n18351;
  assign n34106 = n18354 | n18355;
  assign n34107 = n18362 | ~n18363;
  assign n34108 = n18371 | n18372;
  assign n34109 = n18379 | ~n18380;
  assign n34110 = n18389 | n18390;
  assign n34111 = n18393 | n18394;
  assign n34112 = n18402 | n18403;
  assign n34113 = n18410 | ~n18411;
  assign n34114 = n18416 | n18417;
  assign n34115 = n18420 | n18421;
  assign n34116 = n18428 | ~n18429;
  assign n34117 = n18437 | n18438;
  assign n34118 = n18445 | ~n18446;
  assign n34119 = n18454 | n18455;
  assign n34120 = n18459 | n18460;
  assign n34121 = n18466 | n18467;
  assign n34122 = n18478 | n18479;
  assign n34123 = n18486 | n18487;
  assign n34124 = n18494 | n18495;
  assign n34125 = n18502 | n18503;
  assign n34126 = n18510 | n18511;
  assign n34127 = n18518 | n18519;
  assign n34128 = n18526 | n18527;
  assign n34129 = n18534 | n18535;
  assign n34130 = n18542 | n18543;
  assign n34131 = n18550 | n18551;
  assign n34132 = n18558 | n18559;
  assign n34133 = n18566 | n18567;
  assign n34134 = n18574 | n18575;
  assign n34135 = n18582 | n18583;
  assign n34136 = n18590 | n18591;
  assign n34137 = n18598 | n18599;
  assign n34138 = n18606 | n18607;
  assign n34139 = n18614 | n18615;
  assign n34140 = n18622 | n18623;
  assign n34141 = n18630 | n18631;
  assign n34142 = n18634 | n18635;
  assign n34143 = n18642 | n18643;
  assign n34144 = n18652 | n18653;
  assign n34145 = n18659 | n18660;
  assign n34146 = n18667 | n18668;
  assign n34147 = n18677 | n18678;
  assign n34148 = n18685 | n18686;
  assign n34149 = n18696 | n18697;
  assign n34150 = n18700 | ~n18701;
  assign n34151 = n18707 | n18708;
  assign n34152 = n18721 | ~n18722;
  assign n34153 = n18728 | n18729;
  assign n34154 = n18742 | ~n18743;
  assign n34155 = n18749 | n18750;
  assign n34156 = n18762 | n18763;
  assign n34157 = n18764 | ~n18765;
  assign n34158 = n18771 | n18772;
  assign n34159 = n18779 | n18780;
  assign n34160 = n18782 | n18783;
  assign n34161 = n18788 | ~n18789;
  assign n34162 = n18795 | n18796;
  assign n34163 = n18806 | n18807;
  assign n34164 = n18814 | n18815;
  assign n34165 = n18822 | ~n18823;
  assign n34166 = n18829 | n18830;
  assign n34167 = n18840 | n18841;
  assign n34168 = n18848 | n18849;
  assign n34169 = n18856 | ~n18857;
  assign n34170 = n18863 | n18864;
  assign n34171 = n18874 | n18875;
  assign n34172 = n18882 | n18883;
  assign n34173 = n18890 | ~n18891;
  assign n34174 = n18897 | n18898;
  assign n34175 = n18908 | n18909;
  assign n34176 = n18916 | n18917;
  assign n34177 = n18924 | ~n18925;
  assign n34178 = n18931 | n18932;
  assign n34179 = n18942 | n18943;
  assign n34180 = n18956 | ~n18957;
  assign n34181 = n18968 | n18969;
  assign n34182 = n18972 | n18973;
  assign n34183 = n18981 | n18982;
  assign n34184 = n18989 | ~n18990;
  assign n34185 = n18999 | n19000;
  assign n34186 = n19003 | n19004;
  assign n34187 = n19012 | n19013;
  assign n34188 = n19020 | ~n19021;
  assign n34189 = n19030 | n19031;
  assign n34190 = n19034 | n19035;
  assign n34191 = n19044 | n19045;
  assign n34192 = n19057 | n19058;
  assign n34193 = n19061 | n19062;
  assign n34194 = n19070 | n19071;
  assign n34195 = n19078 | ~n19079;
  assign n34196 = n19088 | n19089;
  assign n34197 = n19092 | n19093;
  assign n34198 = n19102 | n19103;
  assign n34199 = n19115 | n19116;
  assign n34200 = n19119 | n19120;
  assign n34201 = n19128 | n19129;
  assign n34202 = n19136 | ~n19137;
  assign n34203 = n19146 | n19147;
  assign n34204 = n19150 | n19151;
  assign n34205 = n19160 | n19161;
  assign n34206 = n19172 | n19173;
  assign n34207 = n19177 | n19178;
  assign n34208 = n19184 | n19185;
  assign n34209 = n19198 | n19199;
  assign n34210 = n19205 | n19206;
  assign n34211 = n19211 | n19212;
  assign n34212 = n19224 | n19225;
  assign n34213 = n19231 | n19232;
  assign n34214 = n19237 | n19238;
  assign n34215 = n19247 | n19248;
  assign n34216 = n19255 | ~n19256;
  assign n34217 = n19261 | n19262;
  assign n34218 = n19268 | n19269;
  assign n34219 = n19272 | ~n19273;
  assign n34220 = n19281 | n19282;
  assign n34221 = n19289 | ~n19290;
  assign n34222 = n19295 | n19296;
  assign n34223 = n19305 | ~n19306;
  assign n34224 = n19314 | n19315;
  assign n34225 = n19322 | ~n19323;
  assign n34226 = n19328 | n19329;
  assign n34227 = n19338 | ~n19339;
  assign n34228 = n19347 | n19348;
  assign n34229 = n19355 | ~n19356;
  assign n34230 = n19361 | n19362;
  assign n34231 = n19370 | n19371;
  assign n34232 = n19372 | ~n19373;
  assign n34233 = n19381 | n19382;
  assign n34234 = n19389 | ~n19390;
  assign n34235 = n19395 | n19396;
  assign n34236 = n19399 | n19400;
  assign n34237 = n19402 | n19403;
  assign n34238 = n19408 | ~n19409;
  assign n34239 = n19417 | n19418;
  assign n34240 = n19425 | ~n19426;
  assign n34241 = n19435 | n19436;
  assign n34242 = n19439 | n19440;
  assign n34243 = n19448 | n19449;
  assign n34244 = n19456 | ~n19457;
  assign n34245 = n19462 | n19463;
  assign n34246 = n19466 | n19467;
  assign n34247 = n19474 | ~n19475;
  assign n34248 = n19483 | n19484;
  assign n34249 = n19491 | ~n19492;
  assign n34250 = n19501 | n19502;
  assign n34251 = n19505 | n19506;
  assign n34252 = n19514 | n19515;
  assign n34253 = n19522 | ~n19523;
  assign n34254 = n19528 | n19529;
  assign n34255 = n19532 | n19533;
  assign n34256 = n19540 | ~n19541;
  assign n34257 = n19549 | n19550;
  assign n34258 = n19557 | ~n19558;
  assign n34259 = n19567 | n19568;
  assign n34260 = n19571 | n19572;
  assign n34261 = n19580 | n19581;
  assign n34262 = n19588 | ~n19589;
  assign n34263 = n19594 | n19595;
  assign n34264 = n19598 | n19599;
  assign n34265 = n19606 | ~n19607;
  assign n34266 = n19615 | n19616;
  assign n34267 = n19623 | ~n19624;
  assign n34268 = n19633 | n19634;
  assign n34269 = n19637 | n19638;
  assign n34270 = n19646 | n19647;
  assign n34271 = n19654 | ~n19655;
  assign n34272 = n19660 | n19661;
  assign n34273 = n19664 | n19665;
  assign n34274 = n19672 | ~n19673;
  assign n34275 = n19681 | n19682;
  assign n34276 = n19689 | ~n19690;
  assign n34277 = n19699 | n19700;
  assign n34278 = n19703 | n19704;
  assign n34279 = n19712 | n19713;
  assign n34280 = n19720 | ~n19721;
  assign n34281 = n19726 | n19727;
  assign n34282 = n19730 | n19731;
  assign n34283 = n19738 | ~n19739;
  assign n34284 = n19753 | ~n19754;
  assign n34285 = n19766 | ~n19767;
  assign n34286 = n19769 | n19770;
  assign n34287 = n19778 | n19779;
  assign n34288 = n19786 | ~n19787;
  assign n34289 = n19796 | n19797;
  assign n34290 = n19800 | n19801;
  assign n34291 = n19809 | n19810;
  assign n34292 = n19817 | ~n19818;
  assign n34293 = n19827 | n19828;
  assign n34294 = n19831 | n19832;
  assign n34295 = n19840 | n19841;
  assign n34296 = n19848 | ~n19849;
  assign n34297 = n19854 | n19855;
  assign n34298 = n19858 | n19859;
  assign n34299 = n19866 | ~n19867;
  assign n34300 = n19875 | n19876;
  assign n34301 = n19883 | ~n19884;
  assign n34302 = n19893 | n19894;
  assign n34303 = n19897 | n19898;
  assign n34304 = n19906 | n19907;
  assign n34305 = n19914 | ~n19915;
  assign n34306 = n19920 | n19921;
  assign n34307 = n19924 | n19925;
  assign n34308 = n19932 | ~n19933;
  assign n34309 = n19941 | n19942;
  assign n34310 = n19949 | ~n19950;
  assign n34311 = n19959 | n19960;
  assign n34312 = n19963 | n19964;
  assign n34313 = n19972 | n19973;
  assign n34314 = n19980 | ~n19981;
  assign n34315 = n19986 | n19987;
  assign n34316 = n19994 | ~n19995;
  assign n34317 = n19998 | n19999;
  assign n34318 = n20005 | n20006;
  assign n34319 = n20017 | n20018;
  assign n34320 = n20025 | n20026;
  assign n34321 = n20033 | n20034;
  assign n34322 = n20041 | n20042;
  assign n34323 = n20049 | n20050;
  assign n34324 = n20057 | n20058;
  assign n34325 = n20065 | n20066;
  assign n34326 = n20073 | n20074;
  assign n34327 = n20081 | n20082;
  assign n34328 = n20089 | n20090;
  assign n34329 = n20097 | n20098;
  assign n34330 = n20105 | n20106;
  assign n34331 = n20113 | n20114;
  assign n34332 = n20121 | n20122;
  assign n34333 = n20129 | n20130;
  assign n34334 = n20137 | n20138;
  assign n34335 = n20145 | n20146;
  assign n34336 = n20153 | n20154;
  assign n34337 = n20161 | n20162;
  assign n34338 = n20169 | n20170;
  assign n34339 = n20177 | n20178;
  assign n34340 = n20185 | n20186;
  assign n34341 = n20189 | n20190;
  assign n34342 = n20197 | n20198;
  assign n34343 = n20207 | n20208;
  assign n34344 = n20214 | n20215;
  assign n34345 = n20222 | n20223;
  assign n34346 = n20232 | n20233;
  assign n34347 = n20240 | n20241;
  assign n34348 = n20251 | n20252;
  assign n34349 = n20255 | ~n20256;
  assign n34350 = n20262 | n20263;
  assign n34351 = n20276 | ~n20277;
  assign n34352 = n20283 | n20284;
  assign n34353 = n20297 | ~n20298;
  assign n34354 = n20304 | n20305;
  assign n34355 = n20317 | n20318;
  assign n34356 = n20319 | ~n20320;
  assign n34357 = n20326 | n20327;
  assign n34358 = n20334 | n20335;
  assign n34359 = n20337 | n20338;
  assign n34360 = n20343 | ~n20344;
  assign n34361 = n20350 | n20351;
  assign n34362 = n20361 | n20362;
  assign n34363 = n20369 | n20370;
  assign n34364 = n20377 | ~n20378;
  assign n34365 = n20384 | n20385;
  assign n34366 = n20395 | n20396;
  assign n34367 = n20403 | n20404;
  assign n34368 = n20411 | ~n20412;
  assign n34369 = n20418 | n20419;
  assign n34370 = n20429 | n20430;
  assign n34371 = n20437 | n20438;
  assign n34372 = n20445 | ~n20446;
  assign n34373 = n20452 | n20453;
  assign n34374 = n20463 | n20464;
  assign n34375 = n20471 | n20472;
  assign n34376 = n20479 | ~n20480;
  assign n34377 = n20486 | n20487;
  assign n34378 = n20497 | n20498;
  assign n34379 = n20505 | n20506;
  assign n34380 = n20513 | ~n20514;
  assign n34381 = n20520 | n20521;
  assign n34382 = n20531 | n20532;
  assign n34383 = n20541 | ~n20542;
  assign n34384 = n20555 | ~n20556;
  assign n34385 = n20567 | n20568;
  assign n34386 = n20571 | n20572;
  assign n34387 = n20580 | n20581;
  assign n34388 = n20588 | ~n20589;
  assign n34389 = n20598 | n20599;
  assign n34390 = n20602 | n20603;
  assign n34391 = n20611 | n20612;
  assign n34392 = n20619 | ~n20620;
  assign n34393 = n20629 | n20630;
  assign n34394 = n20633 | n20634;
  assign n34395 = n20643 | n20644;
  assign n34396 = n20656 | n20657;
  assign n34397 = n20660 | n20661;
  assign n34398 = n20669 | n20670;
  assign n34399 = n20677 | ~n20678;
  assign n34400 = n20687 | n20688;
  assign n34401 = n20691 | n20692;
  assign n34402 = n20701 | n20702;
  assign n34403 = n20714 | n20715;
  assign n34404 = n20718 | n20719;
  assign n34405 = n20727 | n20728;
  assign n34406 = n20735 | ~n20736;
  assign n34407 = n20744 | n20745;
  assign n34408 = n20749 | n20750;
  assign n34409 = n20756 | n20757;
  assign n34410 = n20770 | n20771;
  assign n34411 = n20777 | n20778;
  assign n34412 = n20783 | n20784;
  assign n34413 = n20796 | n20797;
  assign n34414 = n20803 | n20804;
  assign n34415 = n20809 | n20810;
  assign n34416 = n20819 | n20820;
  assign n34417 = n20827 | ~n20828;
  assign n34418 = n20833 | n20834;
  assign n34419 = n20840 | n20841;
  assign n34420 = n20844 | ~n20845;
  assign n34421 = n20853 | n20854;
  assign n34422 = n20861 | ~n20862;
  assign n34423 = n20867 | n20868;
  assign n34424 = n20877 | ~n20878;
  assign n34425 = n20886 | n20887;
  assign n34426 = n20894 | ~n20895;
  assign n34427 = n20900 | n20901;
  assign n34428 = n20910 | ~n20911;
  assign n34429 = n20919 | n20920;
  assign n34430 = n20927 | ~n20928;
  assign n34431 = n20933 | n20934;
  assign n34432 = n20942 | n20943;
  assign n34433 = n20944 | ~n20945;
  assign n34434 = n20953 | n20954;
  assign n34435 = n20961 | ~n20962;
  assign n34436 = n20967 | n20968;
  assign n34437 = n20971 | n20972;
  assign n34438 = n20974 | n20975;
  assign n34439 = n20980 | ~n20981;
  assign n34440 = n20989 | n20990;
  assign n34441 = n20997 | ~n20998;
  assign n34442 = n21007 | n21008;
  assign n34443 = n21011 | n21012;
  assign n34444 = n21020 | n21021;
  assign n34445 = n21028 | ~n21029;
  assign n34446 = n21034 | n21035;
  assign n34447 = n21038 | n21039;
  assign n34448 = n21046 | ~n21047;
  assign n34449 = n21055 | n21056;
  assign n34450 = n21063 | ~n21064;
  assign n34451 = n21073 | n21074;
  assign n34452 = n21077 | n21078;
  assign n34453 = n21086 | n21087;
  assign n34454 = n21094 | ~n21095;
  assign n34455 = n21100 | n21101;
  assign n34456 = n21104 | n21105;
  assign n34457 = n21112 | ~n21113;
  assign n34458 = n21121 | n21122;
  assign n34459 = n21129 | ~n21130;
  assign n34460 = n21139 | n21140;
  assign n34461 = n21143 | n21144;
  assign n34462 = n21152 | n21153;
  assign n34463 = n21160 | ~n21161;
  assign n34464 = n21166 | n21167;
  assign n34465 = n21170 | n21171;
  assign n34466 = n21178 | ~n21179;
  assign n34467 = n21187 | n21188;
  assign n34468 = n21195 | ~n21196;
  assign n34469 = n21205 | n21206;
  assign n34470 = n21209 | n21210;
  assign n34471 = n21218 | n21219;
  assign n34472 = n21226 | ~n21227;
  assign n34473 = n21232 | n21233;
  assign n34474 = n21236 | n21237;
  assign n34475 = n21244 | ~n21245;
  assign n34476 = n21253 | n21254;
  assign n34477 = n21261 | ~n21262;
  assign n34478 = n21271 | n21272;
  assign n34479 = n21275 | n21276;
  assign n34480 = n21284 | n21285;
  assign n34481 = n21292 | ~n21293;
  assign n34482 = n21298 | n21299;
  assign n34483 = n21302 | n21303;
  assign n34484 = n21310 | ~n21311;
  assign n34485 = n21319 | n21320;
  assign n34486 = n21327 | ~n21328;
  assign n34487 = n21337 | n21338;
  assign n34488 = n21341 | n21342;
  assign n34489 = n21350 | n21351;
  assign n34490 = n21358 | ~n21359;
  assign n34491 = n21364 | n21365;
  assign n34492 = n21368 | n21369;
  assign n34493 = n21376 | ~n21377;
  assign n34494 = n21391 | ~n21392;
  assign n34495 = n21401 | n21402;
  assign n34496 = n21405 | n21406;
  assign n34497 = n21414 | n21415;
  assign n34498 = n21422 | ~n21423;
  assign n34499 = n21432 | n21433;
  assign n34500 = n21436 | n21437;
  assign n34501 = n21445 | n21446;
  assign n34502 = n21453 | ~n21454;
  assign n34503 = n21463 | n21464;
  assign n34504 = n21467 | n21468;
  assign n34505 = n21476 | n21477;
  assign n34506 = n21484 | ~n21485;
  assign n34507 = n21490 | n21491;
  assign n34508 = n21494 | n21495;
  assign n34509 = n21502 | ~n21503;
  assign n34510 = n21511 | n21512;
  assign n34511 = n21519 | ~n21520;
  assign n34512 = n21529 | n21530;
  assign n34513 = n21533 | n21534;
  assign n34514 = n21542 | n21543;
  assign n34515 = n21550 | ~n21551;
  assign n34516 = n21556 | n21557;
  assign n34517 = n21560 | n21561;
  assign n34518 = n21568 | ~n21569;
  assign n34519 = n21577 | n21578;
  assign n34520 = n21585 | ~n21586;
  assign n34521 = n21594 | n21595;
  assign n34522 = n21599 | n21600;
  assign n34523 = n21606 | n21607;
  assign n34524 = n21618 | n21619;
  assign n34525 = n21626 | n21627;
  assign n34526 = n21634 | n21635;
  assign n34527 = n21642 | n21643;
  assign n34528 = n21650 | n21651;
  assign n34529 = n21658 | n21659;
  assign n34530 = n21666 | n21667;
  assign n34531 = n21674 | n21675;
  assign n34532 = n21682 | n21683;
  assign n34533 = n21690 | n21691;
  assign n34534 = n21698 | n21699;
  assign n34535 = n21706 | n21707;
  assign n34536 = n21714 | n21715;
  assign n34537 = n21722 | n21723;
  assign n34538 = n21730 | n21731;
  assign n34539 = n21738 | n21739;
  assign n34540 = n21746 | n21747;
  assign n34541 = n21754 | n21755;
  assign n34542 = n21762 | n21763;
  assign n34543 = n21770 | n21771;
  assign n34544 = n21778 | n21779;
  assign n34545 = n21786 | n21787;
  assign n34546 = n21794 | n21795;
  assign n34547 = n21802 | n21803;
  assign n34548 = n21810 | n21811;
  assign n34549 = n21818 | n21819;
  assign n34550 = n21822 | n21823;
  assign n34551 = n21830 | n21831;
  assign n34552 = n21840 | n21841;
  assign n34553 = n21847 | n21848;
  assign n34554 = n21855 | n21856;
  assign n34555 = n21865 | n21866;
  assign n34556 = n21873 | n21874;
  assign n34557 = n21884 | n21885;
  assign n34558 = n21888 | ~n21889;
  assign n34559 = n21895 | n21896;
  assign n34560 = n21909 | ~n21910;
  assign n34561 = n21916 | n21917;
  assign n34562 = n21930 | ~n21931;
  assign n34563 = n21937 | n21938;
  assign n34564 = n21950 | n21951;
  assign n34565 = n21952 | ~n21953;
  assign n34566 = n21959 | n21960;
  assign n34567 = n21967 | n21968;
  assign n34568 = n21970 | n21971;
  assign n34569 = n21976 | ~n21977;
  assign n34570 = n21983 | n21984;
  assign n34571 = n21994 | n21995;
  assign n34572 = n22002 | n22003;
  assign n34573 = n22010 | ~n22011;
  assign n34574 = n22017 | n22018;
  assign n34575 = n22028 | n22029;
  assign n34576 = n22036 | n22037;
  assign n34577 = n22044 | ~n22045;
  assign n34578 = n22051 | n22052;
  assign n34579 = n22062 | n22063;
  assign n34580 = n22070 | n22071;
  assign n34581 = n22078 | ~n22079;
  assign n34582 = n22085 | n22086;
  assign n34583 = n22096 | n22097;
  assign n34584 = n22104 | n22105;
  assign n34585 = n22112 | ~n22113;
  assign n34586 = n22119 | n22120;
  assign n34587 = n22130 | n22131;
  assign n34588 = n22138 | n22139;
  assign n34589 = n22146 | ~n22147;
  assign n34590 = n22153 | n22154;
  assign n34591 = n22164 | n22165;
  assign n34592 = n22172 | n22173;
  assign n34593 = n22180 | ~n22181;
  assign n34594 = n22187 | n22188;
  assign n34595 = n22198 | n22199;
  assign n34596 = n22208 | n22209;
  assign n34597 = n22222 | n22223;
  assign n34598 = n22226 | n22227;
  assign n34599 = n22235 | n22236;
  assign n34600 = n22243 | ~n22244;
  assign n34601 = n22253 | n22254;
  assign n34602 = n22257 | n22258;
  assign n34603 = n22266 | n22267;
  assign n34604 = n22274 | ~n22275;
  assign n34605 = n22284 | n22285;
  assign n34606 = n22288 | n22289;
  assign n34607 = n22298 | n22299;
  assign n34608 = n22311 | n22312;
  assign n34609 = n22315 | n22316;
  assign n34610 = n22324 | n22325;
  assign n34611 = n22332 | ~n22333;
  assign n34612 = n22342 | n22343;
  assign n34613 = n22346 | n22347;
  assign n34614 = n22356 | n22357;
  assign n34615 = n22368 | n22369;
  assign n34616 = n22373 | n22374;
  assign n34617 = n22380 | n22381;
  assign n34618 = n22394 | n22395;
  assign n34619 = n22401 | n22402;
  assign n34620 = n22407 | n22408;
  assign n34621 = n22420 | n22421;
  assign n34622 = n22427 | n22428;
  assign n34623 = n22433 | n22434;
  assign n34624 = n22443 | n22444;
  assign n34625 = n22451 | ~n22452;
  assign n34626 = n22457 | n22458;
  assign n34627 = n22464 | n22465;
  assign n34628 = n22468 | ~n22469;
  assign n34629 = n22477 | n22478;
  assign n34630 = n22485 | ~n22486;
  assign n34631 = n22491 | n22492;
  assign n34632 = n22501 | ~n22502;
  assign n34633 = n22510 | n22511;
  assign n34634 = n22518 | ~n22519;
  assign n34635 = n22524 | n22525;
  assign n34636 = n22534 | ~n22535;
  assign n34637 = n22543 | n22544;
  assign n34638 = n22551 | ~n22552;
  assign n34639 = n22557 | n22558;
  assign n34640 = n22566 | n22567;
  assign n34641 = n22568 | ~n22569;
  assign n34642 = n22577 | n22578;
  assign n34643 = n22585 | ~n22586;
  assign n34644 = n22591 | n22592;
  assign n34645 = n22595 | n22596;
  assign n34646 = n22598 | n22599;
  assign n34647 = n22604 | ~n22605;
  assign n34648 = n22613 | n22614;
  assign n34649 = n22621 | ~n22622;
  assign n34650 = n22631 | n22632;
  assign n34651 = n22635 | n22636;
  assign n34652 = n22644 | n22645;
  assign n34653 = n22652 | ~n22653;
  assign n34654 = n22658 | n22659;
  assign n34655 = n22662 | n22663;
  assign n34656 = n22670 | ~n22671;
  assign n34657 = n22679 | n22680;
  assign n34658 = n22687 | ~n22688;
  assign n34659 = n22697 | n22698;
  assign n34660 = n22701 | n22702;
  assign n34661 = n22710 | n22711;
  assign n34662 = n22718 | ~n22719;
  assign n34663 = n22724 | n22725;
  assign n34664 = n22728 | n22729;
  assign n34665 = n22736 | ~n22737;
  assign n34666 = n22745 | n22746;
  assign n34667 = n22753 | ~n22754;
  assign n34668 = n22763 | n22764;
  assign n34669 = n22767 | n22768;
  assign n34670 = n22776 | n22777;
  assign n34671 = n22784 | ~n22785;
  assign n34672 = n22790 | n22791;
  assign n34673 = n22794 | n22795;
  assign n34674 = n22802 | ~n22803;
  assign n34675 = n22811 | n22812;
  assign n34676 = n22819 | ~n22820;
  assign n34677 = n22829 | n22830;
  assign n34678 = n22833 | n22834;
  assign n34679 = n22842 | n22843;
  assign n34680 = n22850 | ~n22851;
  assign n34681 = n22856 | n22857;
  assign n34682 = n22860 | n22861;
  assign n34683 = n22868 | ~n22869;
  assign n34684 = n22877 | n22878;
  assign n34685 = n22885 | ~n22886;
  assign n34686 = n22895 | n22896;
  assign n34687 = n22899 | n22900;
  assign n34688 = n22908 | n22909;
  assign n34689 = n22916 | ~n22917;
  assign n34690 = n22922 | n22923;
  assign n34691 = n22926 | n22927;
  assign n34692 = n22934 | ~n22935;
  assign n34693 = n22943 | n22944;
  assign n34694 = n22951 | ~n22952;
  assign n34695 = n22961 | n22962;
  assign n34696 = n22965 | n22966;
  assign n34697 = n22974 | n22975;
  assign n34698 = n22982 | ~n22983;
  assign n34699 = n22988 | n22989;
  assign n34700 = n22992 | n22993;
  assign n34701 = n23000 | ~n23001;
  assign n34702 = n23009 | n23010;
  assign n34703 = n23017 | ~n23018;
  assign n34704 = n23027 | n23028;
  assign n34705 = n23031 | n23032;
  assign n34706 = n23040 | n23041;
  assign n34707 = n23048 | ~n23049;
  assign n34708 = n23054 | n23055;
  assign n34709 = n23058 | n23059;
  assign n34710 = n23066 | ~n23067;
  assign n34711 = n23077 | n23078;
  assign n34712 = n23089 | n23090;
  assign n34713 = n23093 | n23094;
  assign n34714 = n23102 | n23103;
  assign n34715 = n23110 | ~n23111;
  assign n34716 = n23120 | n23121;
  assign n34717 = n23124 | n23125;
  assign n34718 = n23133 | n23134;
  assign n34719 = n23141 | ~n23142;
  assign n34720 = n23151 | n23152;
  assign n34721 = n23155 | n23156;
  assign n34722 = n23164 | n23165;
  assign n34723 = n23172 | ~n23173;
  assign n34724 = n23178 | n23179;
  assign n34725 = n23182 | n23183;
  assign n34726 = n23190 | ~n23191;
  assign n34727 = n23199 | n23200;
  assign n34728 = n23207 | ~n23208;
  assign n34729 = n23217 | n23218;
  assign n34730 = n23221 | n23222;
  assign n34731 = n23230 | n23231;
  assign n34732 = n23238 | ~n23239;
  assign n34733 = n23244 | n23245;
  assign n34734 = n23252 | ~n23253;
  assign n34735 = n23256 | n23257;
  assign n34736 = n23263 | n23264;
  assign n34737 = n23275 | n23276;
  assign n34738 = n23283 | n23284;
  assign n34739 = n23291 | n23292;
  assign n34740 = n23299 | n23300;
  assign n34741 = n23307 | n23308;
  assign n34742 = n23315 | n23316;
  assign n34743 = n23323 | n23324;
  assign n34744 = n23331 | n23332;
  assign n34745 = n23339 | n23340;
  assign n34746 = n23347 | n23348;
  assign n34747 = n23355 | n23356;
  assign n34748 = n23363 | n23364;
  assign n34749 = n23371 | n23372;
  assign n34750 = n23379 | n23380;
  assign n34751 = n23387 | n23388;
  assign n34752 = n23395 | n23396;
  assign n34753 = n23403 | n23404;
  assign n34754 = n23411 | n23412;
  assign n34755 = n23419 | n23420;
  assign n34756 = n23427 | n23428;
  assign n34757 = n23435 | n23436;
  assign n34758 = n23443 | n23444;
  assign n34759 = n23451 | n23452;
  assign n34760 = n23459 | n23460;
  assign n34761 = n23467 | n23468;
  assign n34762 = n23475 | n23476;
  assign n34763 = n23483 | n23484;
  assign n34764 = n23491 | n23492;
  assign n34765 = n23499 | n23500;
  assign n34766 = n23503 | n23504;
  assign n34767 = n23511 | n23512;
  assign n34768 = n23521 | n23522;
  assign n34769 = n23528 | n23529;
  assign n34770 = n23536 | n23537;
  assign n34771 = n23546 | n23547;
  assign n34772 = n23554 | n23555;
  assign n34773 = n23565 | n23566;
  assign n34774 = n23569 | ~n23570;
  assign n34775 = n23576 | n23577;
  assign n34776 = n23590 | ~n23591;
  assign n34777 = n23597 | n23598;
  assign n34778 = n23611 | ~n23612;
  assign n34779 = n23618 | n23619;
  assign n34780 = n23631 | n23632;
  assign n34781 = n23633 | ~n23634;
  assign n34782 = n23640 | n23641;
  assign n34783 = n23648 | n23649;
  assign n34784 = n23651 | n23652;
  assign n34785 = n23657 | ~n23658;
  assign n34786 = n23664 | n23665;
  assign n34787 = n23675 | n23676;
  assign n34788 = n23683 | n23684;
  assign n34789 = n23691 | ~n23692;
  assign n34790 = n23698 | n23699;
  assign n34791 = n23709 | n23710;
  assign n34792 = n23717 | n23718;
  assign n34793 = n23725 | ~n23726;
  assign n34794 = n23732 | n23733;
  assign n34795 = n23743 | n23744;
  assign n34796 = n23751 | n23752;
  assign n34797 = n23759 | ~n23760;
  assign n34798 = n23766 | n23767;
  assign n34799 = n23777 | n23778;
  assign n34800 = n23785 | n23786;
  assign n34801 = n23793 | ~n23794;
  assign n34802 = n23800 | n23801;
  assign n34803 = n23811 | n23812;
  assign n34804 = n23819 | n23820;
  assign n34805 = n23827 | ~n23828;
  assign n34806 = n23834 | n23835;
  assign n34807 = n23845 | n23846;
  assign n34808 = n23853 | n23854;
  assign n34809 = n23861 | ~n23862;
  assign n34810 = n23868 | n23869;
  assign n34811 = n23879 | n23880;
  assign n34812 = n23887 | n23888;
  assign n34813 = n23895 | ~n23896;
  assign n34814 = n23902 | n23903;
  assign n34815 = n23913 | n23914;
  assign n34816 = n23927 | ~n23928;
  assign n34817 = n23939 | n23940;
  assign n34818 = n23943 | n23944;
  assign n34819 = n23952 | n23953;
  assign n34820 = n23960 | ~n23961;
  assign n34821 = n23970 | n23971;
  assign n34822 = n23974 | n23975;
  assign n34823 = n23983 | n23984;
  assign n34824 = n23991 | ~n23992;
  assign n34825 = n24001 | n24002;
  assign n34826 = n24005 | n24006;
  assign n34827 = n24015 | n24016;
  assign n34828 = n24028 | n24029;
  assign n34829 = n24032 | n24033;
  assign n34830 = n24041 | n24042;
  assign n34831 = n24049 | ~n24050;
  assign n34832 = n24058 | n24059;
  assign n34833 = n24063 | n24064;
  assign n34834 = n24070 | n24071;
  assign n34835 = n24084 | n24085;
  assign n34836 = n24091 | n24092;
  assign n34837 = n24097 | n24098;
  assign n34838 = n24110 | n24111;
  assign n34839 = n24117 | n24118;
  assign n34840 = n24123 | n24124;
  assign n34841 = n24133 | n24134;
  assign n34842 = n24141 | ~n24142;
  assign n34843 = n24147 | n24148;
  assign n34844 = n24154 | n24155;
  assign n34845 = n24158 | ~n24159;
  assign n34846 = n24167 | n24168;
  assign n34847 = n24175 | ~n24176;
  assign n34848 = n24181 | n24182;
  assign n34849 = n24191 | ~n24192;
  assign n34850 = n24200 | n24201;
  assign n34851 = n24208 | ~n24209;
  assign n34852 = n24214 | n24215;
  assign n34853 = n24224 | ~n24225;
  assign n34854 = n24233 | n24234;
  assign n34855 = n24241 | ~n24242;
  assign n34856 = n24247 | n24248;
  assign n34857 = n24256 | n24257;
  assign n34858 = n24258 | ~n24259;
  assign n34859 = n24267 | n24268;
  assign n34860 = n24275 | ~n24276;
  assign n34861 = n24281 | n24282;
  assign n34862 = n24285 | n24286;
  assign n34863 = n24288 | n24289;
  assign n34864 = n24294 | ~n24295;
  assign n34865 = n24303 | n24304;
  assign n34866 = n24311 | ~n24312;
  assign n34867 = n24321 | n24322;
  assign n34868 = n24325 | n24326;
  assign n34869 = n24334 | n24335;
  assign n34870 = n24342 | ~n24343;
  assign n34871 = n24348 | n24349;
  assign n34872 = n24352 | n24353;
  assign n34873 = n24360 | ~n24361;
  assign n34874 = n24369 | n24370;
  assign n34875 = n24377 | ~n24378;
  assign n34876 = n24387 | n24388;
  assign n34877 = n24391 | n24392;
  assign n34878 = n24400 | n24401;
  assign n34879 = n24408 | ~n24409;
  assign n34880 = n24414 | n24415;
  assign n34881 = n24418 | n24419;
  assign n34882 = n24426 | ~n24427;
  assign n34883 = n24435 | n24436;
  assign n34884 = n24443 | ~n24444;
  assign n34885 = n24453 | n24454;
  assign n34886 = n24457 | n24458;
  assign n34887 = n24466 | n24467;
  assign n34888 = n24474 | ~n24475;
  assign n34889 = n24480 | n24481;
  assign n34890 = n24484 | n24485;
  assign n34891 = n24492 | ~n24493;
  assign n34892 = n24501 | n24502;
  assign n34893 = n24509 | ~n24510;
  assign n34894 = n24519 | n24520;
  assign n34895 = n24523 | n24524;
  assign n34896 = n24532 | n24533;
  assign n34897 = n24540 | ~n24541;
  assign n34898 = n24546 | n24547;
  assign n34899 = n24550 | n24551;
  assign n34900 = n24558 | ~n24559;
  assign n34901 = n24567 | n24568;
  assign n34902 = n24575 | ~n24576;
  assign n34903 = n24585 | n24586;
  assign n34904 = n24589 | n24590;
  assign n34905 = n24598 | n24599;
  assign n34906 = n24606 | ~n24607;
  assign n34907 = n24612 | n24613;
  assign n34908 = n24616 | n24617;
  assign n34909 = n24624 | ~n24625;
  assign n34910 = n24633 | n24634;
  assign n34911 = n24641 | ~n24642;
  assign n34912 = n24651 | n24652;
  assign n34913 = n24655 | n24656;
  assign n34914 = n24664 | n24665;
  assign n34915 = n24672 | ~n24673;
  assign n34916 = n24678 | n24679;
  assign n34917 = n24682 | n24683;
  assign n34918 = n24690 | ~n24691;
  assign n34919 = n24699 | n24700;
  assign n34920 = n24707 | ~n24708;
  assign n34921 = n24717 | n24718;
  assign n34922 = n24721 | n24722;
  assign n34923 = n24730 | n24731;
  assign n34924 = n24738 | ~n24739;
  assign n34925 = n24744 | n24745;
  assign n34926 = n24748 | n24749;
  assign n34927 = n24756 | ~n24757;
  assign n34928 = n24765 | n24766;
  assign n34929 = n24773 | ~n24774;
  assign n34930 = n24783 | n24784;
  assign n34931 = n24787 | n24788;
  assign n34932 = n24796 | n24797;
  assign n34933 = n24804 | ~n24805;
  assign n34934 = n24810 | n24811;
  assign n34935 = n24814 | n24815;
  assign n34936 = n24822 | ~n24823;
  assign n34937 = n24837 | ~n24838;
  assign n34938 = n24850 | ~n24851;
  assign n34939 = n24853 | n24854;
  assign n34940 = n24862 | n24863;
  assign n34941 = n24870 | ~n24871;
  assign n34942 = n24880 | n24881;
  assign n34943 = n24884 | n24885;
  assign n34944 = n24893 | n24894;
  assign n34945 = n24901 | ~n24902;
  assign n34946 = n24911 | n24912;
  assign n34947 = n24915 | n24916;
  assign n34948 = n24924 | n24925;
  assign n34949 = n24932 | ~n24933;
  assign n34950 = n24938 | n24939;
  assign n34951 = n24942 | n24943;
  assign n34952 = n24950 | ~n24951;
  assign n34953 = n24959 | n24960;
  assign n34954 = n24967 | ~n24968;
  assign n34955 = n24976 | n24977;
  assign n34956 = n24981 | n24982;
  assign n34957 = n24988 | n24989;
  assign n34958 = n25000 | n25001;
  assign n34959 = n25008 | n25009;
  assign n34960 = n25016 | n25017;
  assign n34961 = n25024 | n25025;
  assign n34962 = n25032 | n25033;
  assign n34963 = n25040 | n25041;
  assign n34964 = n25048 | n25049;
  assign n34965 = n25056 | n25057;
  assign n34966 = n25064 | n25065;
  assign n34967 = n25072 | n25073;
  assign n34968 = n25080 | n25081;
  assign n34969 = n25088 | n25089;
  assign n34970 = n25096 | n25097;
  assign n34971 = n25104 | n25105;
  assign n34972 = n25112 | n25113;
  assign n34973 = n25120 | n25121;
  assign n34974 = n25128 | n25129;
  assign n34975 = n25136 | n25137;
  assign n34976 = n25144 | n25145;
  assign n34977 = n25152 | n25153;
  assign n34978 = n25160 | n25161;
  assign n34979 = n25168 | n25169;
  assign n34980 = n25176 | n25177;
  assign n34981 = n25184 | n25185;
  assign n34982 = n25192 | n25193;
  assign n34983 = n25200 | n25201;
  assign n34984 = n25208 | n25209;
  assign n34985 = n25216 | n25217;
  assign n34986 = n25224 | n25225;
  assign n34987 = n25232 | n25233;
  assign n34988 = n25240 | n25241;
  assign n34989 = n25244 | n25245;
  assign n34990 = n25252 | n25253;
  assign n34991 = n25262 | n25263;
  assign n34992 = n25269 | n25270;
  assign n34993 = n25277 | n25278;
  assign n34994 = n25287 | n25288;
  assign n34995 = n25295 | n25296;
  assign n34996 = n25306 | n25307;
  assign n34997 = n25310 | ~n25311;
  assign n34998 = n25317 | n25318;
  assign n34999 = n25331 | ~n25332;
  assign n35000 = n25338 | n25339;
  assign n35001 = n25352 | ~n25353;
  assign n35002 = n25359 | n25360;
  assign n35003 = n25372 | n25373;
  assign n35004 = n25374 | ~n25375;
  assign n35005 = n25381 | n25382;
  assign n35006 = n25389 | n25390;
  assign n35007 = n25392 | n25393;
  assign n35008 = n25398 | ~n25399;
  assign n35009 = n25405 | n25406;
  assign n35010 = n25416 | n25417;
  assign n35011 = n25424 | n25425;
  assign n35012 = n25432 | ~n25433;
  assign n35013 = n25439 | n25440;
  assign n35014 = n25450 | n25451;
  assign n35015 = n25458 | n25459;
  assign n35016 = n25466 | ~n25467;
  assign n35017 = n25473 | n25474;
  assign n35018 = n25484 | n25485;
  assign n35019 = n25492 | n25493;
  assign n35020 = n25500 | ~n25501;
  assign n35021 = n25507 | n25508;
  assign n35022 = n25518 | n25519;
  assign n35023 = n25526 | n25527;
  assign n35024 = n25534 | ~n25535;
  assign n35025 = n25541 | n25542;
  assign n35026 = n25552 | n25553;
  assign n35027 = n25560 | n25561;
  assign n35028 = n25568 | ~n25569;
  assign n35029 = n25575 | n25576;
  assign n35030 = n25586 | n25587;
  assign n35031 = n25594 | n25595;
  assign n35032 = n25602 | ~n25603;
  assign n35033 = n25609 | n25610;
  assign n35034 = n25620 | n25621;
  assign n35035 = n25628 | n25629;
  assign n35036 = n25636 | ~n25637;
  assign n35037 = n25643 | n25644;
  assign n35038 = n25654 | n25655;
  assign n35039 = n25662 | n25663;
  assign n35040 = n25670 | ~n25671;
  assign n35041 = n25677 | n25678;
  assign n35042 = n25688 | n25689;
  assign n35043 = n25698 | ~n25699;
  assign n35044 = n25712 | ~n25713;
  assign n35045 = n25724 | n25725;
  assign n35046 = n25728 | n25729;
  assign n35047 = n25737 | n25738;
  assign n35048 = n25745 | ~n25746;
  assign n35049 = n25755 | n25756;
  assign n35050 = n25759 | n25760;
  assign n35051 = n25768 | n25769;
  assign n35052 = n25776 | ~n25777;
  assign n35053 = n25786 | n25787;
  assign n35054 = n25790 | n25791;
  assign n35055 = n25800 | n25801;
  assign n35056 = n25812 | n25813;
  assign n35057 = n25817 | n25818;
  assign n35058 = n25824 | n25825;
  assign n35059 = n25838 | n25839;
  assign n35060 = n25845 | n25846;
  assign n35061 = n25851 | n25852;
  assign n35062 = n25864 | n25865;
  assign n35063 = n25871 | n25872;
  assign n35064 = n25877 | n25878;
  assign n35065 = n25887 | n25888;
  assign n35066 = n25895 | ~n25896;
  assign n35067 = n25901 | n25902;
  assign n35068 = n25908 | n25909;
  assign n35069 = n25912 | ~n25913;
  assign n35070 = n25921 | n25922;
  assign n35071 = n25929 | ~n25930;
  assign n35072 = n25935 | n25936;
  assign n35073 = n25945 | ~n25946;
  assign n35074 = n25954 | n25955;
  assign n35075 = n25962 | ~n25963;
  assign n35076 = n25968 | n25969;
  assign n35077 = n25978 | ~n25979;
  assign n35078 = n25987 | n25988;
  assign n35079 = n25995 | ~n25996;
  assign n35080 = n26001 | n26002;
  assign n35081 = n26010 | n26011;
  assign n35082 = n26012 | ~n26013;
  assign n35083 = n26021 | n26022;
  assign n35084 = n26029 | ~n26030;
  assign n35085 = n26035 | n26036;
  assign n35086 = n26039 | n26040;
  assign n35087 = n26042 | n26043;
  assign n35088 = n26048 | ~n26049;
  assign n35089 = n26057 | n26058;
  assign n35090 = n26065 | ~n26066;
  assign n35091 = n26075 | n26076;
  assign n35092 = n26079 | n26080;
  assign n35093 = n26088 | n26089;
  assign n35094 = n26096 | ~n26097;
  assign n35095 = n26102 | n26103;
  assign n35096 = n26106 | n26107;
  assign n35097 = n26114 | ~n26115;
  assign n35098 = n26123 | n26124;
  assign n35099 = n26131 | ~n26132;
  assign n35100 = n26141 | n26142;
  assign n35101 = n26145 | n26146;
  assign n35102 = n26154 | n26155;
  assign n35103 = n26162 | ~n26163;
  assign n35104 = n26168 | n26169;
  assign n35105 = n26172 | n26173;
  assign n35106 = n26180 | ~n26181;
  assign n35107 = n26189 | n26190;
  assign n35108 = n26197 | ~n26198;
  assign n35109 = n26207 | n26208;
  assign n35110 = n26211 | n26212;
  assign n35111 = n26220 | n26221;
  assign n35112 = n26228 | ~n26229;
  assign n35113 = n26234 | n26235;
  assign n35114 = n26238 | n26239;
  assign n35115 = n26246 | ~n26247;
  assign n35116 = n26255 | n26256;
  assign n35117 = n26263 | ~n26264;
  assign n35118 = n26273 | n26274;
  assign n35119 = n26277 | n26278;
  assign n35120 = n26286 | n26287;
  assign n35121 = n26294 | ~n26295;
  assign n35122 = n26300 | n26301;
  assign n35123 = n26304 | n26305;
  assign n35124 = n26312 | ~n26313;
  assign n35125 = n26321 | n26322;
  assign n35126 = n26329 | ~n26330;
  assign n35127 = n26339 | n26340;
  assign n35128 = n26343 | n26344;
  assign n35129 = n26352 | n26353;
  assign n35130 = n26360 | ~n26361;
  assign n35131 = n26366 | n26367;
  assign n35132 = n26370 | n26371;
  assign n35133 = n26378 | ~n26379;
  assign n35134 = n26387 | n26388;
  assign n35135 = n26395 | ~n26396;
  assign n35136 = n26405 | n26406;
  assign n35137 = n26409 | n26410;
  assign n35138 = n26418 | n26419;
  assign n35139 = n26426 | ~n26427;
  assign n35140 = n26432 | n26433;
  assign n35141 = n26436 | n26437;
  assign n35142 = n26444 | ~n26445;
  assign n35143 = n26453 | n26454;
  assign n35144 = n26461 | ~n26462;
  assign n35145 = n26471 | n26472;
  assign n35146 = n26475 | n26476;
  assign n35147 = n26484 | n26485;
  assign n35148 = n26492 | ~n26493;
  assign n35149 = n26498 | n26499;
  assign n35150 = n26502 | n26503;
  assign n35151 = n26510 | ~n26511;
  assign n35152 = n26519 | n26520;
  assign n35153 = n26527 | ~n26528;
  assign n35154 = n26537 | n26538;
  assign n35155 = n26541 | n26542;
  assign n35156 = n26550 | n26551;
  assign n35157 = n26558 | ~n26559;
  assign n35158 = n26564 | n26565;
  assign n35159 = n26568 | n26569;
  assign n35160 = n26576 | ~n26577;
  assign n35161 = n26585 | n26586;
  assign n35162 = n26593 | ~n26594;
  assign n35163 = n26603 | n26604;
  assign n35164 = n26607 | n26608;
  assign n35165 = n26616 | n26617;
  assign n35166 = n26624 | ~n26625;
  assign n35167 = n26630 | n26631;
  assign n35168 = n26634 | n26635;
  assign n35169 = n26642 | ~n26643;
  assign n35170 = n26657 | ~n26658;
  assign n35171 = n26667 | n26668;
  assign n35172 = n26671 | n26672;
  assign n35173 = n26680 | n26681;
  assign n35174 = n26688 | ~n26689;
  assign n35175 = n26698 | n26699;
  assign n35176 = n26702 | n26703;
  assign n35177 = n26711 | n26712;
  assign n35178 = n26719 | ~n26720;
  assign n35179 = n26729 | n26730;
  assign n35180 = n26733 | n26734;
  assign n35181 = n26742 | n26743;
  assign n35182 = n26750 | ~n26751;
  assign n35183 = n26756 | n26757;
  assign n35184 = n26764 | ~n26765;
  assign n35185 = n26768 | n26769;
  assign n35186 = n26775 | n26776;
  assign n35187 = n26786 | n26787;
  assign n35188 = n26795 | n26796;
  assign n35189 = n26803 | n26804;
  assign n35190 = n26811 | n26812;
  assign n35191 = n26819 | n26820;
  assign n35192 = n26827 | n26828;
  assign n35193 = n26835 | n26836;
  assign n35194 = n26843 | n26844;
  assign n35195 = n26851 | n26852;
  assign n35196 = n26859 | n26860;
  assign n35197 = n26867 | n26868;
  assign n35198 = n26875 | n26876;
  assign n35199 = n26883 | n26884;
  assign n35200 = n26891 | n26892;
  assign n35201 = n26899 | n26900;
  assign n35202 = n26907 | n26908;
  assign n35203 = n26915 | n26916;
  assign n35204 = n26923 | n26924;
  assign n35205 = n26931 | n26932;
  assign n35206 = n26939 | n26940;
  assign n35207 = n26947 | n26948;
  assign n35208 = n26955 | n26956;
  assign n35209 = n26963 | n26964;
  assign n35210 = n26971 | n26972;
  assign n35211 = n26979 | n26980;
  assign n35212 = n26987 | n26988;
  assign n35213 = n26995 | n26996;
  assign n35214 = n27003 | n27004;
  assign n35215 = n27011 | n27012;
  assign n35216 = n27019 | n27020;
  assign n35217 = n27027 | n27028;
  assign n35218 = n27035 | n27036;
  assign n35219 = n27043 | n27044;
  assign n35220 = n27051 | n27052;
  assign n35221 = n27059 | n27060;
  assign n35222 = n27067 | n27068;
  assign n35223 = n27071 | n27072;
  assign n35224 = n27075 | n27076;
  assign n35225 = n27080 | n27081;
  assign n35226 = n27090 | n27091;
  assign n35227 = n27098 | ~n27099;
  assign n35228 = n27100 | n27101;
  assign n35229 = n27108 | n27109;
  assign n35230 = n27118 | n27119;
  assign n35231 = n27126 | n27127;
  assign n35232 = n27137 | n27138;
  assign n35233 = n27141 | ~n27142;
  assign n35234 = n27148 | n27149;
  assign n35235 = n27162 | ~n27163;
  assign n35236 = n27169 | n27170;
  assign n35237 = n27183 | ~n27184;
  assign n35238 = n27190 | n27191;
  assign n35239 = n27203 | n27204;
  assign n35240 = n27205 | ~n27206;
  assign n35241 = n27212 | n27213;
  assign n35242 = n27220 | n27221;
  assign n35243 = n27223 | n27224;
  assign n35244 = n27229 | ~n27230;
  assign n35245 = n27236 | n27237;
  assign n35246 = n27247 | n27248;
  assign n35247 = n27255 | n27256;
  assign n35248 = n27263 | ~n27264;
  assign n35249 = n27270 | n27271;
  assign n35250 = n27281 | n27282;
  assign n35251 = n27289 | n27290;
  assign n35252 = n27297 | ~n27298;
  assign n35253 = n27304 | n27305;
  assign n35254 = n27315 | n27316;
  assign n35255 = n27323 | n27324;
  assign n35256 = n27331 | ~n27332;
  assign n35257 = n27338 | n27339;
  assign n35258 = n27349 | n27350;
  assign n35259 = n27357 | n27358;
  assign n35260 = n27365 | ~n27366;
  assign n35261 = n27372 | n27373;
  assign n35262 = n27383 | n27384;
  assign n35263 = n27391 | n27392;
  assign n35264 = n27399 | ~n27400;
  assign n35265 = n27406 | n27407;
  assign n35266 = n27417 | n27418;
  assign n35267 = n27425 | n27426;
  assign n35268 = n27433 | ~n27434;
  assign n35269 = n27440 | n27441;
  assign n35270 = n27451 | n27452;
  assign n35271 = n27459 | n27460;
  assign n35272 = n27467 | ~n27468;
  assign n35273 = n27474 | n27475;
  assign n35274 = n27485 | n27486;
  assign n35275 = n27493 | n27494;
  assign n35276 = n27501 | ~n27502;
  assign n35277 = n27508 | n27509;
  assign n35278 = n27519 | n27520;
  assign n35279 = n27527 | n27528;
  assign n35280 = n27535 | ~n27536;
  assign n35281 = n27542 | n27543;
  assign n35282 = n27553 | n27554;
  assign n35283 = n27569 | n27570;
  assign n35284 = n27573 | n27574;
  assign n35285 = n27582 | n27583;
  assign n35286 = n27590 | ~n27591;
  assign n35287 = n27600 | n27601;
  assign n35288 = n27604 | n27605;
  assign n35289 = n27613 | n27614;
  assign n35290 = n27621 | ~n27622;
  assign n35291 = n27630 | n27631;
  assign n35292 = n27635 | n27636;
  assign n35293 = n27642 | n27643;
  assign n35294 = n27654 | n27655;
  assign n35295 = n27662 | ~n27663;
  assign n35296 = n27667 | n27668;
  assign n35297 = n27673 | n27674;
  assign n35298 = n27682 | n27683;
  assign n35299 = n27687 | n27688;
  assign n35300 = n27694 | n27695;
  assign n35301 = n27700 | n27701;
  assign n35302 = n27710 | n27711;
  assign n35303 = n27718 | ~n27719;
  assign n35304 = n27724 | n27725;
  assign n35305 = n27731 | n27732;
  assign n35306 = n27735 | ~n27736;
  assign n35307 = n27744 | n27745;
  assign n35308 = n27752 | ~n27753;
  assign n35309 = n27758 | n27759;
  assign n35310 = n27768 | ~n27769;
  assign n35311 = n27777 | n27778;
  assign n35312 = n27785 | ~n27786;
  assign n35313 = n27791 | n27792;
  assign n35314 = n27801 | ~n27802;
  assign n35315 = n27810 | n27811;
  assign n35316 = n27818 | ~n27819;
  assign n35317 = n27824 | n27825;
  assign n35318 = n27833 | n27834;
  assign n35319 = n27835 | ~n27836;
  assign n35320 = n27844 | n27845;
  assign n35321 = n27852 | ~n27853;
  assign n35322 = n27858 | n27859;
  assign n35323 = n27862 | n27863;
  assign n35324 = n27865 | n27866;
  assign n35325 = n27871 | ~n27872;
  assign n35326 = n27880 | n27881;
  assign n35327 = n27888 | ~n27889;
  assign n35328 = n27898 | n27899;
  assign n35329 = n27902 | n27903;
  assign n35330 = n27911 | n27912;
  assign n35331 = n27919 | ~n27920;
  assign n35332 = n27925 | n27926;
  assign n35333 = n27929 | n27930;
  assign n35334 = n27937 | ~n27938;
  assign n35335 = n27946 | n27947;
  assign n35336 = n27954 | ~n27955;
  assign n35337 = n27964 | n27965;
  assign n35338 = n27968 | n27969;
  assign n35339 = n27977 | n27978;
  assign n35340 = n27985 | ~n27986;
  assign n35341 = n27991 | n27992;
  assign n35342 = n27995 | n27996;
  assign n35343 = n28003 | ~n28004;
  assign n35344 = n28012 | n28013;
  assign n35345 = n28020 | ~n28021;
  assign n35346 = n28030 | n28031;
  assign n35347 = n28034 | n28035;
  assign n35348 = n28043 | n28044;
  assign n35349 = n28051 | ~n28052;
  assign n35350 = n28057 | n28058;
  assign n35351 = n28061 | n28062;
  assign n35352 = n28069 | ~n28070;
  assign n35353 = n28078 | n28079;
  assign n35354 = n28086 | ~n28087;
  assign n35355 = n28096 | n28097;
  assign n35356 = n28100 | n28101;
  assign n35357 = n28109 | n28110;
  assign n35358 = n28117 | ~n28118;
  assign n35359 = n28123 | n28124;
  assign n35360 = n28127 | n28128;
  assign n35361 = n28135 | ~n28136;
  assign n35362 = n28144 | n28145;
  assign n35363 = n28152 | ~n28153;
  assign n35364 = n28162 | n28163;
  assign n35365 = n28166 | n28167;
  assign n35366 = n28175 | n28176;
  assign n35367 = n28183 | ~n28184;
  assign n35368 = n28189 | n28190;
  assign n35369 = n28193 | n28194;
  assign n35370 = n28201 | ~n28202;
  assign n35371 = n28210 | n28211;
  assign n35372 = n28218 | ~n28219;
  assign n35373 = n28228 | n28229;
  assign n35374 = n28232 | n28233;
  assign n35375 = n28241 | n28242;
  assign n35376 = n28249 | ~n28250;
  assign n35377 = n28255 | n28256;
  assign n35378 = n28259 | n28260;
  assign n35379 = n28267 | ~n28268;
  assign n35380 = n28276 | n28277;
  assign n35381 = n28284 | ~n28285;
  assign n35382 = n28294 | n28295;
  assign n35383 = n28298 | n28299;
  assign n35384 = n28307 | n28308;
  assign n35385 = n28315 | ~n28316;
  assign n35386 = n28321 | n28322;
  assign n35387 = n28325 | n28326;
  assign n35388 = n28333 | ~n28334;
  assign n35389 = n28342 | n28343;
  assign n35390 = n28350 | ~n28351;
  assign n35391 = n28360 | n28361;
  assign n35392 = n28364 | n28365;
  assign n35393 = n28373 | n28374;
  assign n35394 = n28381 | ~n28382;
  assign n35395 = n28387 | n28388;
  assign n35396 = n28391 | n28392;
  assign n35397 = n28399 | ~n28400;
  assign n35398 = n28408 | n28409;
  assign n35399 = n28416 | ~n28417;
  assign n35400 = n28426 | n28427;
  assign n35401 = n28430 | n28431;
  assign n35402 = n28439 | n28440;
  assign n35403 = n28447 | ~n28448;
  assign n35404 = n28453 | n28454;
  assign n35405 = n28457 | n28458;
  assign n35406 = n28465 | ~n28466;
  assign n35407 = n28474 | n28475;
  assign n35408 = n28482 | ~n28483;
  assign n35409 = n28492 | n28493;
  assign n35410 = n28496 | n28497;
  assign n35411 = n28505 | n28506;
  assign n35412 = n28513 | ~n28514;
  assign n35413 = n28519 | n28520;
  assign n35414 = n28523 | n28524;
  assign n35415 = n28531 | ~n28532;
  assign n35416 = n28542 | n28543;
  assign n35417 = n28550 | n28551;
  assign n35418 = n28559 | n28560;
  assign n35419 = n28567 | ~n28568;
  assign n35420 = n28577 | n28578;
  assign n35421 = n28581 | n28582;
  assign n35422 = n28590 | n28591;
  assign n35423 = n28598 | ~n28599;
  assign n35424 = n28607 | n28608;
  assign n35425 = n28612 | n28613;
  assign n35426 = n28619 | n28620;
  assign n35427 = n28634 | ~n28635;
  assign n35428 = n28641 | n28642;
  assign n35429 = n28649 | n28650;
  assign n35430 = n28657 | n28658;
  assign n35431 = n28665 | n28666;
  assign n35432 = n28673 | n28674;
  assign n35433 = n28681 | n28682;
  assign n35434 = n28689 | n28690;
  assign n35435 = n28697 | n28698;
  assign n35436 = n28705 | n28706;
  assign n35437 = n28713 | n28714;
  assign n35438 = n28721 | n28722;
  assign n35439 = n28729 | n28730;
  assign n35440 = n28737 | n28738;
  assign n35441 = n28745 | n28746;
  assign n35442 = n28753 | n28754;
  assign n35443 = n28761 | n28762;
  assign n35444 = n28769 | n28770;
  assign n35445 = n28777 | n28778;
  assign n35446 = n28785 | n28786;
  assign n35447 = n28793 | n28794;
  assign n35448 = n28801 | n28802;
  assign n35449 = n28809 | n28810;
  assign n35450 = n28817 | n28818;
  assign n35451 = n28825 | n28826;
  assign n35452 = n28833 | n28834;
  assign n35453 = n28841 | n28842;
  assign n35454 = n28849 | n28850;
  assign n35455 = n28857 | n28858;
  assign n35456 = n28865 | n28866;
  assign n35457 = n28873 | n28874;
  assign n35458 = n28881 | n28882;
  assign n35459 = n28889 | n28890;
  assign n35460 = n28897 | n28898;
  assign n35461 = n28905 | n28906;
  assign n35462 = n28913 | n28914;
  assign n35463 = n28921 | n28922;
  assign n35464 = n28929 | n28930;
  assign n35465 = n28937 | n28938;
  assign n35466 = n28941 | n28942;
  assign n35467 = n28945 | n28946;
  assign n35468 = n28950 | n28951;
  assign n35469 = n28961 | ~n28962;
  assign n35470 = n28963 | n28964;
  assign n35471 = n28971 | n28972;
  assign n35472 = n28981 | n28982;
  assign n35473 = n28989 | n28990;
  assign n35474 = n29000 | n29001;
  assign n35475 = n29004 | ~n29005;
  assign n35476 = n29011 | n29012;
  assign n35477 = n29025 | ~n29026;
  assign n35478 = n29032 | n29033;
  assign n35479 = n29046 | ~n29047;
  assign n35480 = n29053 | n29054;
  assign n35481 = n29066 | n29067;
  assign n35482 = n29068 | ~n29069;
  assign n35483 = n29075 | n29076;
  assign n35484 = n29083 | n29084;
  assign n35485 = n29086 | n29087;
  assign n35486 = n29092 | ~n29093;
  assign n35487 = n29099 | n29100;
  assign n35488 = n29110 | n29111;
  assign n35489 = n29118 | n29119;
  assign n35490 = n29126 | ~n29127;
  assign n35491 = n29133 | n29134;
  assign n35492 = n29144 | n29145;
  assign n35493 = n29152 | n29153;
  assign n35494 = n29160 | ~n29161;
  assign n35495 = n29167 | n29168;
  assign n35496 = n29178 | n29179;
  assign n35497 = n29186 | n29187;
  assign n35498 = n29194 | ~n29195;
  assign n35499 = n29201 | n29202;
  assign n35500 = n29212 | n29213;
  assign n35501 = n29220 | n29221;
  assign n35502 = n29228 | ~n29229;
  assign n35503 = n29235 | n29236;
  assign n35504 = n29246 | n29247;
  assign n35505 = n29254 | n29255;
  assign n35506 = n29262 | ~n29263;
  assign n35507 = n29269 | n29270;
  assign n35508 = n29280 | n29281;
  assign n35509 = n29288 | n29289;
  assign n35510 = n29296 | ~n29297;
  assign n35511 = n29303 | n29304;
  assign n35512 = n29314 | n29315;
  assign n35513 = n29322 | n29323;
  assign n35514 = n29330 | ~n29331;
  assign n35515 = n29337 | n29338;
  assign n35516 = n29348 | n29349;
  assign n35517 = n29356 | n29357;
  assign n35518 = n29364 | ~n29365;
  assign n35519 = n29371 | n29372;
  assign n35520 = n29382 | n29383;
  assign n35521 = n29390 | n29391;
  assign n35522 = n29398 | ~n29399;
  assign n35523 = n29405 | n29406;
  assign n35524 = n29416 | n29417;
  assign n35525 = n29424 | n29425;
  assign n35526 = n29432 | ~n29433;
  assign n35527 = n29439 | n29440;
  assign n35528 = n29450 | n29451;
  assign n35529 = n29466 | n29467;
  assign n35530 = n29470 | n29471;
  assign n35531 = n29479 | n29480;
  assign n35532 = n29487 | ~n29488;
  assign n35533 = n29496 | n29497;
  assign n35534 = n29501 | n29502;
  assign n35535 = n29508 | n29509;
  assign n35536 = n29523 | ~n29524;
  assign n35537 = n29530 | ~n29531;
  assign n35538 = n29535 | n29536;
  assign n35539 = n29541 | n29542;
  assign n35540 = n29550 | n29551;
  assign n35541 = n29555 | n29556;
  assign n35542 = n29562 | n29563;
  assign n35543 = n29568 | n29569;
  assign n35544 = n29578 | n29579;
  assign n35545 = n29586 | ~n29587;
  assign n35546 = n29592 | n29593;
  assign n35547 = n29599 | n29600;
  assign n35548 = n29603 | ~n29604;
  assign n35549 = n29612 | n29613;
  assign n35550 = n29620 | ~n29621;
  assign n35551 = n29626 | n29627;
  assign n35552 = n29636 | ~n29637;
  assign n35553 = n29645 | n29646;
  assign n35554 = n29653 | ~n29654;
  assign n35555 = n29659 | n29660;
  assign n35556 = n29669 | ~n29670;
  assign n35557 = n29678 | n29679;
  assign n35558 = n29686 | ~n29687;
  assign n35559 = n29692 | n29693;
  assign n35560 = n29701 | n29702;
  assign n35561 = n29703 | ~n29704;
  assign n35562 = n29712 | n29713;
  assign n35563 = n29720 | ~n29721;
  assign n35564 = n29726 | n29727;
  assign n35565 = n29730 | n29731;
  assign n35566 = n29733 | n29734;
  assign n35567 = n29739 | ~n29740;
  assign n35568 = n29748 | n29749;
  assign n35569 = n29756 | ~n29757;
  assign n35570 = n29766 | n29767;
  assign n35571 = n29770 | n29771;
  assign n35572 = n29779 | n29780;
  assign n35573 = n29787 | ~n29788;
  assign n35574 = n29793 | n29794;
  assign n35575 = n29797 | n29798;
  assign n35576 = n29805 | ~n29806;
  assign n35577 = n29814 | n29815;
  assign n35578 = n29822 | ~n29823;
  assign n35579 = n29832 | n29833;
  assign n35580 = n29836 | n29837;
  assign n35581 = n29845 | n29846;
  assign n35582 = n29853 | ~n29854;
  assign n35583 = n29859 | n29860;
  assign n35584 = n29863 | n29864;
  assign n35585 = n29871 | ~n29872;
  assign n35586 = n29880 | n29881;
  assign n35587 = n29888 | ~n29889;
  assign n35588 = n29898 | n29899;
  assign n35589 = n29902 | n29903;
  assign n35590 = n29911 | n29912;
  assign n35591 = n29919 | ~n29920;
  assign n35592 = n29925 | n29926;
  assign n35593 = n29929 | n29930;
  assign n35594 = n29937 | ~n29938;
  assign n35595 = n29946 | n29947;
  assign n35596 = n29954 | ~n29955;
  assign n35597 = n29964 | n29965;
  assign n35598 = n29968 | n29969;
  assign n35599 = n29977 | n29978;
  assign n35600 = n29985 | ~n29986;
  assign n35601 = n29991 | n29992;
  assign n35602 = n29995 | n29996;
  assign n35603 = n30003 | ~n30004;
  assign n35604 = n30012 | n30013;
  assign n35605 = n30020 | ~n30021;
  assign n35606 = n30030 | n30031;
  assign n35607 = n30034 | n30035;
  assign n35608 = n30043 | n30044;
  assign n35609 = n30051 | ~n30052;
  assign n35610 = n30057 | n30058;
  assign n35611 = n30061 | n30062;
  assign n35612 = n30069 | ~n30070;
  assign n35613 = n30078 | n30079;
  assign n35614 = n30086 | ~n30087;
  assign n35615 = n30096 | n30097;
  assign n35616 = n30100 | n30101;
  assign n35617 = n30109 | n30110;
  assign n35618 = n30117 | ~n30118;
  assign n35619 = n30123 | n30124;
  assign n35620 = n30127 | n30128;
  assign n35621 = n30135 | ~n30136;
  assign n35622 = n30144 | n30145;
  assign n35623 = n30152 | ~n30153;
  assign n35624 = n30162 | n30163;
  assign n35625 = n30166 | n30167;
  assign n35626 = n30175 | n30176;
  assign n35627 = n30183 | ~n30184;
  assign n35628 = n30189 | n30190;
  assign n35629 = n30193 | n30194;
  assign n35630 = n30201 | ~n30202;
  assign n35631 = n30210 | n30211;
  assign n35632 = n30218 | ~n30219;
  assign n35633 = n30228 | n30229;
  assign n35634 = n30232 | n30233;
  assign n35635 = n30241 | n30242;
  assign n35636 = n30249 | ~n30250;
  assign n35637 = n30255 | n30256;
  assign n35638 = n30259 | n30260;
  assign n35639 = n30267 | ~n30268;
  assign n35640 = n30276 | n30277;
  assign n35641 = n30284 | ~n30285;
  assign n35642 = n30294 | n30295;
  assign n35643 = n30298 | n30299;
  assign n35644 = n30307 | n30308;
  assign n35645 = n30315 | ~n30316;
  assign n35646 = n30321 | n30322;
  assign n35647 = n30325 | n30326;
  assign n35648 = n30333 | ~n30334;
  assign n35649 = n30342 | n30343;
  assign n35650 = n30350 | ~n30351;
  assign n35651 = n30360 | n30361;
  assign n35652 = n30364 | n30365;
  assign n35653 = n30373 | n30374;
  assign n35654 = n30381 | ~n30382;
  assign n35655 = n30387 | n30388;
  assign n35656 = n30391 | n30392;
  assign n35657 = n30399 | ~n30400;
  assign n35658 = n30408 | n30409;
  assign n35659 = n30416 | ~n30417;
  assign n35660 = n30426 | n30427;
  assign n35661 = n30430 | n30431;
  assign n35662 = n30439 | n30440;
  assign n35663 = n30447 | ~n30448;
  assign n35664 = n30453 | n30454;
  assign n35665 = n30457 | n30458;
  assign n35666 = n30465 | ~n30466;
  assign n35667 = n30480 | ~n30481;
  assign n35668 = n30486 | n30487;
  assign n35669 = n30495 | n30496;
  assign n35670 = n30503 | ~n30504;
  assign n35671 = n30512 | n30513;
  assign n35672 = n30517 | n30518;
  assign n35673 = n30524 | n30525;
  assign n35674 = n30539 | ~n30540;
  assign n35675 = n30551 | ~n30552;
  assign n35676 = n30559 | n30560;
  assign n35677 = n30565 | n30566;
  assign n35678 = n30573 | ~n30574;
  assign n35679 = n30582 | n30583;
  assign n35680 = n30592 | n30593;
  assign n35681 = n30602 | n30603;
  assign n35682 = n30609 | n30610;
  assign n35683 = n30617 | ~n30618;
  assign n35684 = n30626 | n30627;
  assign n35685 = n30636 | n30637;
  assign n35686 = n30646 | n30647;
  assign n35687 = n30653 | n30654;
  assign n35688 = n30661 | ~n30662;
  assign n35689 = n30670 | n30671;
  assign n35690 = n30680 | n30681;
  assign n35691 = n30690 | n30691;
  assign n35692 = n30697 | n30698;
  assign n35693 = n30705 | ~n30706;
  assign n35694 = n30714 | n30715;
  assign n35695 = n30724 | n30725;
  assign n35696 = n30734 | n30735;
  assign n35697 = n30741 | n30742;
  assign n35698 = n30749 | ~n30750;
  assign n35699 = n30758 | n30759;
  assign n35700 = n30768 | n30769;
  assign n35701 = n30778 | n30779;
  assign n35702 = n30785 | n30786;
  assign n35703 = n30793 | ~n30794;
  assign n35704 = n30802 | n30803;
  assign n35705 = n30812 | n30813;
  assign n35706 = n30822 | n30823;
  assign n35707 = n30829 | n30830;
  assign n35708 = n30837 | ~n30838;
  assign n35709 = n30846 | n30847;
  assign n35710 = n30856 | n30857;
  assign n35711 = n30866 | n30867;
  assign n35712 = n30873 | n30874;
  assign n35713 = n30881 | ~n30882;
  assign n35714 = n30890 | n30891;
  assign n35715 = n30900 | n30901;
  assign n35716 = n30910 | n30911;
  assign n35717 = n30917 | n30918;
  assign n35718 = n30925 | ~n30926;
  assign n35719 = n30934 | n30935;
  assign n35720 = n30944 | n30945;
  assign n35721 = n30954 | n30955;
  assign n35722 = n30961 | n30962;
  assign n35723 = n30969 | ~n30970;
  assign n35724 = n30978 | n30979;
  assign n35725 = n30988 | n30989;
  assign n35726 = n30998 | n30999;
  assign n35727 = n31005 | n31006;
  assign n35728 = n31013 | ~n31014;
  assign n35729 = n31022 | n31023;
  assign n35730 = n31032 | n31033;
  assign n35731 = n31042 | n31043;
  assign n35732 = n31049 | n31050;
  assign n35733 = n31052 | n31053;
  assign n35734 = n31058 | ~n31059;
  assign n35735 = n31067 | n31068;
  assign n35736 = n31079 | n31080;
  assign n35737 = n31081 | ~n31082;
  assign n35738 = n31090 | n31091;
  assign n35739 = n31103 | ~n31104;
  assign n35740 = n31112 | n31113;
  assign n35741 = n31125 | ~n31126;
  assign n35742 = n31134 | n31135;
  assign n35743 = n31144 | n31145;
  assign n35744 = n31148 | ~n31149;
  assign n35745 = n31157 | n31158;
  assign n35746 = n31165 | n31166;
  assign n35747 = n31169 | n31170;
  assign n35748 = n31175 | n31176;
  assign n35749 = ~n31184 | n31179 | ~n31183;
  assign n35750 = n31188 | n31189;
  assign n35751 = n31193 | n31194;
  assign n35752 = n31201 | n31202;
  assign n35753 = n31215 | n31216;
  assign n35754 = n31225 | n31226;
  assign n35755 = n31233 | n31228 | n31232;
  assign n35756 = n31239 | n31240;
  assign n35757 = n31251 | n31246 | n31250;
  assign n35758 = n31257 | n31258;
  assign n35759 = n31269 | n31264 | n31268;
  assign n35760 = n31275 | n31276;
  assign n35761 = n31287 | n31282 | n31286;
  assign n35762 = n31293 | n31294;
  assign n35763 = n31305 | n31300 | n31304;
  assign n35764 = n31311 | n31312;
  assign n35765 = n31323 | n31318 | n31322;
  assign n35766 = n31329 | n31330;
  assign n35767 = n31341 | n31336 | n31340;
  assign n35768 = n31347 | n31348;
  assign n35769 = n31359 | n31354 | n31358;
  assign n35770 = n31365 | n31366;
  assign n35771 = n31377 | n31372 | n31376;
  assign n35772 = n31383 | n31384;
  assign n35773 = n31395 | n31390 | n31394;
  assign n35774 = n31401 | n31402;
  assign n35775 = n31413 | n31408 | n31412;
  assign n35776 = n31419 | n31420;
  assign n35777 = n31431 | n31426 | n31430;
  assign n35778 = n31437 | n31438;
  assign n35779 = n31449 | n31444 | n31448;
  assign n35780 = n31455 | n31456;
  assign n35781 = n31467 | n31462 | n31466;
  assign n35782 = n31473 | n31474;
  assign n35783 = n31485 | n31480 | n31484;
  assign n35784 = n31491 | n31492;
  assign n35785 = n31503 | n31498 | n31502;
  assign n35786 = n31509 | n31510;
  assign n35787 = n31521 | n31516 | n31520;
  assign n35788 = n31527 | n31528;
  assign n35789 = n31539 | n31534 | n31538;
  assign n35790 = n31545 | n31546;
  assign n35791 = n31557 | n31552 | n31556;
  assign n35792 = n31563 | n31564;
  assign n35793 = n31575 | n31570 | n31574;
  assign n35794 = n31581 | n31582;
  assign n35795 = n31593 | n31588 | n31592;
  assign n35796 = n31599 | n31600;
  assign n35797 = n31611 | n31606 | n31610;
  assign n35798 = n31617 | n31618;
  assign n35799 = n31629 | n31624 | n31628;
  assign n35800 = n31635 | n31636;
  assign n35801 = n31647 | n31642 | n31646;
  assign n35802 = n31653 | n31654;
  assign n35803 = n31665 | n31660 | n31664;
  assign n35804 = n31671 | n31672;
  assign n35805 = n31683 | n31678 | n31682;
  assign n35806 = n31689 | n31690;
  assign n35807 = n31701 | n31696 | n31700;
  assign n35808 = n31707 | n31708;
  assign n35809 = n31716 | n31717;
  assign n35810 = n31733 | n31734;
  assign n35811 = n31740 | n31741;
  assign n35812 = n31743 | n31744;
  assign n35813 = n31747 | n31748;
  assign n35814 = n31754 | n31755;
  assign n35815 = n31761 | n31762;
  assign n35816 = n31766 | n31767;
  assign n35817 = n31771 | n31772;
  assign po0  = ~n31779;
  assign po1  = ~n30530;
  assign po2  = ~n29514;
  assign po3  = ~n28625;
  assign po4  = ~n27648;
  assign po5  = ~n26781;
  assign po6  = ~n25830;
  assign po7  = ~n24994;
  assign po8  = ~n24076;
  assign po9  = ~n23269;
  assign po10  = ~n22386;
  assign po11  = ~n21612;
  assign po12  = ~n20762;
  assign po13  = ~n20011;
  assign po14  = ~n19190;
  assign po15  = ~n18472;
  assign po16  = ~n17690;
  assign po17  = ~n17001;
  assign po18  = ~n16248;
  assign po19  = ~n15586;
  assign po20  = ~n14866;
  assign po21  = ~n14233;
  assign po22  = ~n13548;
  assign po23  = ~n12948;
  assign po24  = ~n12296;
  assign po25  = ~n11719;
  assign po26  = ~n11097;
  assign po27  = ~n10555;
  assign po28  = ~n9969;
  assign po29  = ~n9457;
  assign po30  = ~n8896;
  assign po31  = ~n8411;
  assign po32  = ~n7885;
  assign po33  = ~n7428;
  assign po34  = ~n6937;
  assign po35  = ~n6507;
  assign po36  = ~n6051;
  assign po37  = ~n5648;
  assign po38  = ~n5223;
  assign po39  = ~n4851;
  assign po40  = ~n4461;
  assign po41  = ~n4115;
  assign po42  = ~n3754;
  assign po43  = ~n3444;
  assign po44  = ~n3116;
  assign po45  = ~n2833;
  assign po46  = ~n2536;
  assign po47  = ~n2283;
  assign po48  = ~n2021;
  assign po49  = ~n1796;
  assign po50  = ~n1567;
  assign po51  = ~n1374;
  assign po52  = ~n1179;
  assign po53  = ~n1016;
  assign po54  = ~n855;
  assign po55  = ~n720;
  assign po56  = ~n592;
  assign po57  = ~n487;
  assign po58  = ~n393;
  assign po59  = ~n321;
  assign po60  = ~n263;
  assign po61  = ~n214;
  assign po62  = ~n197;
  assign po63  = ~n193;
endmodule
