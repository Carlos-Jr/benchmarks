module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379,
    n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414,
    n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463,
    n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n625,
    n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667,
    n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681,
    n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730,
    n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n758,
    n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885,
    n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1186;
  assign n22 = ~pi5  & pi7 ;
  assign n23 = pi7  & pi8 ;
  assign n24 = ~pi5  & n23;
  assign n25 = pi8  & n22;
  assign n26 = ~pi0  & ~pi1 ;
  assign n27 = pi2  & ~pi9 ;
  assign n28 = n26 & n27;
  assign n29 = n1062 & n28;
  assign n30 = ~pi7  & pi9 ;
  assign n31 = ~n1062 & ~n30;
  assign n32 = pi1  & ~n31;
  assign n33 = pi1  & ~pi7 ;
  assign n34 = ~pi5  & ~pi9 ;
  assign n35 = ~n33 & n34;
  assign n36 = ~n32 & ~n35;
  assign n37 = pi0  & ~pi2 ;
  assign n38 = ~n36 & n37;
  assign n39 = ~n29 & ~n38;
  assign n40 = ~pi3  & ~n39;
  assign n41 = ~pi0  & pi9 ;
  assign n42 = pi1  & ~n41;
  assign n43 = ~pi3  & ~pi5 ;
  assign n44 = ~pi1  & pi9 ;
  assign n45 = n43 & ~n44;
  assign n46 = ~n42 & ~n44;
  assign n47 = n43 & n46;
  assign n48 = ~n42 & n45;
  assign n49 = pi0  & ~pi9 ;
  assign n50 = ~pi1  & ~n49;
  assign n51 = pi1  & ~pi9 ;
  assign n52 = ~pi7  & ~n51;
  assign n53 = ~n50 & n52;
  assign n54 = ~n1063 & ~n53;
  assign n55 = ~pi2  & ~n54;
  assign n56 = ~pi0  & pi5 ;
  assign n57 = pi0  & ~pi1 ;
  assign n58 = pi2  & ~n57;
  assign n59 = pi1  & pi2 ;
  assign n60 = ~pi2  & ~pi5 ;
  assign n61 = ~pi0  & ~n60;
  assign n62 = ~n59 & ~n61;
  assign n63 = ~n56 & ~n58;
  assign n64 = ~pi9  & ~n1064;
  assign n65 = ~pi2  & ~pi3 ;
  assign n66 = pi9  & ~n65;
  assign n67 = pi0  & pi3 ;
  assign n68 = ~n66 & ~n67;
  assign n69 = ~pi1  & ~n68;
  assign n70 = pi1  & ~pi3 ;
  assign n71 = ~n69 & ~n70;
  assign n72 = ~n64 & ~n70;
  assign n73 = ~n69 & n72;
  assign n74 = ~n64 & n71;
  assign n75 = ~pi7  & ~n1065;
  assign n76 = ~n55 & ~n75;
  assign n77 = ~pi8  & ~n76;
  assign n78 = ~n40 & ~n77;
  assign n79 = ~pi6  & ~n78;
  assign n80 = ~pi0  & ~pi2 ;
  assign n81 = n44 & n80;
  assign n82 = ~pi5  & ~n81;
  assign n83 = pi6  & ~n82;
  assign n84 = ~pi0  & ~pi9 ;
  assign n85 = pi0  & pi9 ;
  assign n86 = ~n84 & ~n85;
  assign n87 = ~n41 & ~n49;
  assign n88 = pi1  & pi5 ;
  assign n89 = pi2  & n88;
  assign n90 = pi1  & ~n1066;
  assign n91 = pi2  & n90;
  assign n92 = pi5  & n91;
  assign n93 = pi2  & pi5 ;
  assign n94 = n90 & n93;
  assign n95 = ~n1066 & n89;
  assign n96 = ~n83 & ~n1067;
  assign n97 = pi3  & ~n96;
  assign n98 = ~pi2  & ~n49;
  assign n99 = ~pi3  & n42;
  assign n100 = n98 & ~n99;
  assign n101 = ~pi6  & ~n98;
  assign n102 = pi5  & ~n101;
  assign n103 = pi6  & ~n98;
  assign n104 = pi1  & n65;
  assign n105 = n65 & n90;
  assign n106 = ~n1066 & n104;
  assign n107 = ~n103 & ~n1068;
  assign n108 = pi5  & ~n107;
  assign n109 = ~n100 & n102;
  assign n110 = pi2  & pi9 ;
  assign n111 = ~pi2  & n51;
  assign n112 = ~n110 & ~n111;
  assign n113 = ~pi0  & ~pi3 ;
  assign n114 = pi6  & n113;
  assign n115 = ~n112 & n113;
  assign n116 = pi6  & n115;
  assign n117 = ~n112 & n114;
  assign n118 = ~n1069 & ~n1070;
  assign n119 = ~n97 & n118;
  assign n120 = pi8  & ~n119;
  assign n121 = ~pi1  & ~pi9 ;
  assign n122 = ~pi2  & pi6 ;
  assign n123 = pi3  & ~n122;
  assign n124 = n121 & ~n123;
  assign n125 = ~n110 & ~n124;
  assign n126 = ~pi8  & ~n125;
  assign n127 = ~pi1  & ~n41;
  assign n128 = ~pi8  & ~n127;
  assign n129 = ~pi1  & pi2 ;
  assign n130 = n49 & n129;
  assign n131 = n27 & n57;
  assign n132 = ~n128 & ~n1071;
  assign n133 = pi3  & ~n132;
  assign n134 = pi1  & ~pi8 ;
  assign n135 = pi2  & ~pi3 ;
  assign n136 = n44 & n135;
  assign n137 = ~n134 & ~n136;
  assign n138 = ~pi0  & ~n137;
  assign n139 = ~n133 & ~n138;
  assign n140 = ~n126 & ~n138;
  assign n141 = ~n133 & n140;
  assign n142 = ~n126 & n139;
  assign n143 = ~pi5  & ~n1072;
  assign n144 = ~pi8  & n121;
  assign n145 = ~pi0  & n65;
  assign n146 = ~pi3  & n80;
  assign n147 = n144 & n1073;
  assign n148 = ~n143 & ~n147;
  assign n149 = pi8  & ~n96;
  assign n150 = ~pi5  & ~n132;
  assign n151 = ~n149 & ~n150;
  assign n152 = pi3  & ~n151;
  assign n153 = ~pi5  & ~n140;
  assign n154 = pi8  & ~n118;
  assign n155 = ~n147 & ~n154;
  assign n156 = ~n147 & ~n153;
  assign n157 = ~n154 & n156;
  assign n158 = ~n153 & n155;
  assign n159 = ~n152 & n1074;
  assign n160 = ~n152 & n156;
  assign n161 = ~n154 & n160;
  assign n162 = ~n120 & n148;
  assign n163 = ~pi7  & ~n1075;
  assign n164 = ~n79 & ~n163;
  assign n165 = ~pi4  & ~n164;
  assign n166 = pi4  & pi8 ;
  assign n167 = ~pi6  & ~pi9 ;
  assign n168 = ~n166 & ~n167;
  assign n169 = ~pi6  & pi8 ;
  assign n170 = pi5  & ~n169;
  assign n171 = ~pi8  & ~pi9 ;
  assign n172 = ~pi6  & n171;
  assign n173 = pi6  & n166;
  assign n174 = ~n172 & ~n173;
  assign n175 = pi5  & ~n174;
  assign n176 = ~n168 & n170;
  assign n177 = pi6  & ~pi9 ;
  assign n178 = pi4  & pi9 ;
  assign n179 = ~n177 & ~n178;
  assign n180 = pi5  & pi6 ;
  assign n181 = ~pi8  & ~n180;
  assign n182 = ~n179 & ~n180;
  assign n183 = ~pi8  & n182;
  assign n184 = ~n179 & n181;
  assign n185 = ~n1076 & ~n1077;
  assign n186 = ~pi1  & ~pi3 ;
  assign n187 = ~pi7  & n80;
  assign n188 = ~pi2  & n186;
  assign n189 = ~pi0  & ~pi7 ;
  assign n190 = n188 & n189;
  assign n191 = n186 & n187;
  assign n192 = ~pi7  & ~n185;
  assign n193 = n188 & n192;
  assign n194 = ~pi0  & n193;
  assign n195 = ~n185 & n1078;
  assign n196 = ~n165 & ~n1079;
  assign n197 = ~pi2  & ~pi8 ;
  assign n198 = n84 & n197;
  assign n199 = n80 & n171;
  assign n200 = pi0  & pi8 ;
  assign n201 = pi8  & n85;
  assign n202 = pi9  & n200;
  assign n203 = pi2  & n1081;
  assign n204 = n110 & n200;
  assign n205 = ~n1080 & ~n1082;
  assign n206 = pi5  & ~n205;
  assign n207 = ~pi5  & pi8 ;
  assign n208 = pi6  & pi9 ;
  assign n209 = ~n207 & ~n208;
  assign n210 = ~pi0  & ~n209;
  assign n211 = pi8  & pi9 ;
  assign n212 = ~pi8  & pi9 ;
  assign n213 = pi8  & ~pi9 ;
  assign n214 = ~n212 & ~n213;
  assign n215 = ~n171 & ~n211;
  assign n216 = pi5  & ~pi8 ;
  assign n217 = ~pi6  & pi9 ;
  assign n218 = ~n216 & ~n217;
  assign n219 = pi8  & n208;
  assign n220 = ~pi8  & n34;
  assign n221 = ~n219 & ~n220;
  assign n222 = n1083 & n218;
  assign n223 = ~n210 & n1084;
  assign n224 = pi2  & ~n223;
  assign n225 = ~n206 & ~n224;
  assign n226 = ~pi4  & ~n225;
  assign n227 = ~n166 & ~n216;
  assign n228 = ~pi6  & ~n227;
  assign n229 = ~n178 & ~n228;
  assign n230 = n80 & ~n217;
  assign n231 = ~n217 & ~n229;
  assign n232 = n80 & n231;
  assign n233 = ~n229 & n230;
  assign n234 = ~n226 & ~n1085;
  assign n235 = ~pi1  & ~n234;
  assign n236 = n56 & n212;
  assign n237 = pi6  & pi8 ;
  assign n238 = pi0  & ~n237;
  assign n239 = ~n209 & ~n237;
  assign n240 = pi0  & n239;
  assign n241 = ~n209 & n238;
  assign n242 = ~n236 & ~n1086;
  assign n243 = ~pi2  & ~n242;
  assign n244 = ~pi6  & ~pi8 ;
  assign n245 = ~pi0  & pi6 ;
  assign n246 = ~pi2  & ~n245;
  assign n247 = n207 & ~n246;
  assign n248 = ~n244 & ~n247;
  assign n249 = ~pi9  & ~n248;
  assign n250 = ~n243 & ~n249;
  assign n251 = pi1  & ~n250;
  assign n252 = n27 & n169;
  assign n253 = ~n251 & ~n252;
  assign n254 = ~pi4  & ~n253;
  assign n255 = ~pi1  & ~n225;
  assign n256 = ~n252 & ~n255;
  assign n257 = ~n251 & n256;
  assign n258 = ~pi4  & ~n257;
  assign n259 = ~pi1  & n80;
  assign n260 = ~pi1  & ~pi2 ;
  assign n261 = ~pi0  & n260;
  assign n262 = ~pi2  & n26;
  assign n263 = ~n217 & n1087;
  assign n264 = ~n229 & n263;
  assign n265 = ~n258 & ~n264;
  assign n266 = ~n235 & ~n254;
  assign n267 = ~pi3  & ~n1088;
  assign n268 = pi5  & n197;
  assign n269 = ~pi3  & ~pi8 ;
  assign n270 = pi0  & ~n207;
  assign n271 = ~n207 & ~n269;
  assign n272 = pi0  & n271;
  assign n273 = ~n269 & n270;
  assign n274 = ~n268 & ~n1089;
  assign n275 = ~pi1  & ~n274;
  assign n276 = pi3  & pi8 ;
  assign n277 = ~pi2  & ~n276;
  assign n278 = ~pi0  & ~n277;
  assign n279 = ~pi2  & pi8 ;
  assign n280 = pi0  & n279;
  assign n281 = pi0  & ~pi5 ;
  assign n282 = ~n56 & ~n281;
  assign n283 = ~n280 & n282;
  assign n284 = pi1  & ~n283;
  assign n285 = ~n278 & ~n284;
  assign n286 = ~n275 & n285;
  assign n287 = ~pi6  & ~n286;
  assign n288 = ~pi1  & pi6 ;
  assign n289 = pi2  & ~n288;
  assign n290 = ~pi1  & ~pi8 ;
  assign n291 = pi3  & ~n290;
  assign n292 = ~pi2  & ~n290;
  assign n293 = ~pi1  & pi8 ;
  assign n294 = pi6  & n293;
  assign n295 = ~n289 & ~n290;
  assign n296 = ~n292 & ~n294;
  assign n297 = pi3  & n1090;
  assign n298 = ~n289 & n291;
  assign n299 = ~pi0  & pi8 ;
  assign n300 = ~pi2  & ~n299;
  assign n301 = pi0  & pi1 ;
  assign n302 = ~pi1  & ~pi6 ;
  assign n303 = ~n301 & ~n302;
  assign n304 = ~n299 & n303;
  assign n305 = ~pi2  & n304;
  assign n306 = n300 & n303;
  assign n307 = ~n1091 & ~n1092;
  assign n308 = ~pi5  & ~n307;
  assign n309 = ~pi9  & ~n308;
  assign n310 = ~n287 & n309;
  assign n311 = ~pi1  & pi3 ;
  assign n312 = pi3  & ~pi8 ;
  assign n313 = n260 & n312;
  assign n314 = n197 & n311;
  assign n315 = ~n88 & ~n1093;
  assign n316 = pi0  & ~n315;
  assign n317 = pi3  & n59;
  assign n318 = pi5  & ~n65;
  assign n319 = ~pi5  & ~n317;
  assign n320 = ~n65 & ~n319;
  assign n321 = ~n317 & ~n318;
  assign n322 = ~n316 & ~n1094;
  assign n323 = pi6  & ~n322;
  assign n324 = n216 & n317;
  assign n325 = pi9  & ~n324;
  assign n326 = ~n323 & n325;
  assign n327 = ~pi4  & ~n326;
  assign n328 = ~n287 & ~n308;
  assign n329 = ~pi9  & ~n328;
  assign n330 = ~n323 & ~n324;
  assign n331 = pi9  & ~n330;
  assign n332 = ~n329 & ~n331;
  assign n333 = ~pi4  & ~n332;
  assign n334 = ~n310 & n327;
  assign n335 = ~n267 & ~n1095;
  assign n336 = ~pi7  & ~n335;
  assign n337 = n51 & n279;
  assign n338 = n98 & ~n301;
  assign n339 = pi2  & ~n26;
  assign n340 = ~pi8  & ~n339;
  assign n341 = ~n338 & ~n339;
  assign n342 = ~pi8  & n341;
  assign n343 = ~n338 & n340;
  assign n344 = ~n337 & ~n1096;
  assign n345 = pi7  & ~n344;
  assign n346 = ~n28 & ~n345;
  assign n347 = ~pi4  & ~pi6 ;
  assign n348 = ~pi6  & n43;
  assign n349 = ~pi4  & n348;
  assign n350 = n43 & n347;
  assign n351 = ~pi4  & ~n346;
  assign n352 = ~pi6  & n351;
  assign n353 = n43 & n352;
  assign n354 = ~n346 & n1097;
  assign n355 = ~n336 & ~n1098;
  assign n356 = ~n121 & n1083;
  assign n357 = n1083 & ~n290;
  assign n358 = pi2  & ~n1099;
  assign n359 = pi5  & ~n171;
  assign n360 = n1083 & ~n299;
  assign n361 = ~n171 & ~n1081;
  assign n362 = pi5  & ~n1100;
  assign n363 = ~n1081 & n359;
  assign n364 = ~pi5  & ~n110;
  assign n365 = pi1  & ~n364;
  assign n366 = pi5  & ~n299;
  assign n367 = pi5  & n1100;
  assign n368 = n1083 & n366;
  assign n369 = ~pi5  & n110;
  assign n370 = ~n1102 & ~n369;
  assign n371 = pi1  & ~n370;
  assign n372 = ~n1101 & n365;
  assign n373 = ~n358 & ~n1103;
  assign n374 = ~pi3  & ~n373;
  assign n375 = n66 & n293;
  assign n376 = pi5  & ~n311;
  assign n377 = ~pi2  & n171;
  assign n378 = ~n376 & n377;
  assign n379 = ~n375 & ~n378;
  assign n380 = pi0  & ~n379;
  assign n381 = ~n374 & ~n380;
  assign n382 = ~pi6  & ~n381;
  assign n383 = pi6  & ~n44;
  assign n384 = ~n51 & ~n383;
  assign n385 = pi8  & ~n384;
  assign n386 = pi1  & pi9 ;
  assign n387 = ~n121 & ~n386;
  assign n388 = n269 & ~n387;
  assign n389 = ~n385 & ~n388;
  assign n390 = ~pi2  & ~n389;
  assign n391 = pi2  & n386;
  assign n392 = ~n293 & ~n391;
  assign n393 = pi6  & ~n392;
  assign n394 = pi8  & ~n27;
  assign n395 = pi2  & n171;
  assign n396 = ~n394 & ~n395;
  assign n397 = ~n393 & n396;
  assign n398 = pi3  & ~n397;
  assign n399 = ~n390 & ~n398;
  assign n400 = n281 & ~n399;
  assign n401 = ~n382 & ~n400;
  assign n402 = ~pi4  & ~n401;
  assign n403 = pi3  & ~n279;
  assign n404 = pi5  & ~n403;
  assign n405 = pi2  & ~pi5 ;
  assign n406 = pi3  & ~n405;
  assign n407 = pi8  & ~n406;
  assign n408 = ~n404 & ~n407;
  assign n409 = pi1  & ~n408;
  assign n410 = ~pi5  & pi6 ;
  assign n411 = ~pi3  & n410;
  assign n412 = ~pi8  & n410;
  assign n413 = n186 & n412;
  assign n414 = n290 & n411;
  assign n415 = ~n409 & ~n1104;
  assign n416 = ~pi9  & ~n415;
  assign n417 = pi1  & pi8 ;
  assign n418 = pi6  & ~n417;
  assign n419 = ~pi9  & ~n418;
  assign n420 = ~pi2  & ~n419;
  assign n421 = ~pi1  & n212;
  assign n422 = ~pi8  & n44;
  assign n423 = ~n420 & ~n1105;
  assign n424 = pi3  & ~n423;
  assign n425 = pi2  & ~n169;
  assign n426 = pi1  & ~n425;
  assign n427 = pi5  & ~n277;
  assign n428 = ~pi1  & ~n277;
  assign n429 = ~n425 & ~n428;
  assign n430 = pi5  & ~n429;
  assign n431 = ~n426 & n427;
  assign n432 = ~n70 & ~n212;
  assign n433 = ~pi3  & pi9 ;
  assign n434 = ~pi6  & ~n433;
  assign n435 = ~n432 & ~n433;
  assign n436 = ~pi6  & n435;
  assign n437 = ~n432 & n434;
  assign n438 = pi6  & ~pi8 ;
  assign n439 = pi1  & n433;
  assign n440 = n438 & n439;
  assign n441 = ~pi4  & ~n440;
  assign n442 = ~pi4  & ~n1107;
  assign n443 = ~n440 & n442;
  assign n444 = ~n1107 & n441;
  assign n445 = ~n1106 & n1108;
  assign n446 = ~n424 & n445;
  assign n447 = ~n416 & n446;
  assign n448 = ~pi5  & ~n213;
  assign n449 = ~n213 & ~n244;
  assign n450 = ~n211 & ~n438;
  assign n451 = ~pi5  & n1109;
  assign n452 = ~pi5  & ~n244;
  assign n453 = ~n213 & n452;
  assign n454 = ~n244 & n448;
  assign n455 = n188 & ~n1110;
  assign n456 = pi4  & ~n455;
  assign n457 = ~pi0  & ~n456;
  assign n458 = ~n1107 & ~n440;
  assign n459 = ~n1106 & n458;
  assign n460 = ~n424 & n459;
  assign n461 = ~n424 & ~n440;
  assign n462 = ~n1106 & n461;
  assign n463 = ~n416 & n462;
  assign n464 = ~n1107 & n463;
  assign n465 = ~n416 & n460;
  assign n466 = ~pi4  & ~n1111;
  assign n467 = ~pi3  & pi4 ;
  assign n468 = pi4  & n65;
  assign n469 = ~pi2  & n467;
  assign n470 = ~pi1  & n1112;
  assign n471 = n260 & n467;
  assign n472 = ~pi1  & n467;
  assign n473 = ~n1110 & n472;
  assign n474 = ~pi2  & n473;
  assign n475 = ~n1110 & n1113;
  assign n476 = ~n466 & ~n1114;
  assign n477 = ~pi0  & ~n476;
  assign n478 = ~n447 & n457;
  assign n479 = ~n402 & ~n1115;
  assign n480 = ~pi7  & ~n479;
  assign n481 = pi7  & n211;
  assign n482 = pi0  & ~n481;
  assign n483 = n23 & n85;
  assign n484 = ~n84 & ~n483;
  assign n485 = pi1  & ~n484;
  assign n486 = n42 & ~n482;
  assign n487 = n49 & n290;
  assign n488 = ~n1116 & ~n487;
  assign n489 = ~pi5  & ~pi6 ;
  assign n490 = ~pi4  & n65;
  assign n491 = n489 & n490;
  assign n492 = ~pi4  & ~n488;
  assign n493 = n65 & n492;
  assign n494 = n489 & n493;
  assign n495 = ~n488 & n491;
  assign n496 = ~n480 & ~n1117;
  assign n497 = pi5  & pi9 ;
  assign n498 = ~n171 & ~n497;
  assign n499 = pi2  & ~n498;
  assign n500 = ~pi3  & ~n438;
  assign n501 = ~n499 & n500;
  assign n502 = pi1  & ~n170;
  assign n503 = pi5  & pi8 ;
  assign n504 = n217 & n503;
  assign n505 = ~n220 & ~n504;
  assign n506 = pi2  & ~n505;
  assign n507 = pi3  & ~n170;
  assign n508 = ~n412 & ~n507;
  assign n509 = ~n506 & n508;
  assign n510 = pi1  & ~n509;
  assign n511 = ~n501 & n502;
  assign n512 = pi6  & n405;
  assign n513 = pi2  & n410;
  assign n514 = pi3  & ~n217;
  assign n515 = pi2  & pi6 ;
  assign n516 = pi3  & ~pi9 ;
  assign n517 = pi6  & ~n65;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n514 & ~n515;
  assign n520 = ~pi1  & ~n1120;
  assign n521 = ~n1119 & ~n520;
  assign n522 = ~pi3  & ~n499;
  assign n523 = pi1  & ~n522;
  assign n524 = ~pi6  & ~n516;
  assign n525 = ~n523 & n524;
  assign n526 = n65 & ~n134;
  assign n527 = n88 & ~n169;
  assign n528 = ~n526 & ~n527;
  assign n529 = ~n525 & n528;
  assign n530 = ~n1118 & n521;
  assign n531 = ~pi0  & ~n1121;
  assign n532 = ~n433 & ~n503;
  assign n533 = ~pi6  & ~n532;
  assign n534 = pi3  & n448;
  assign n535 = ~n533 & ~n534;
  assign n536 = pi2  & ~n535;
  assign n537 = ~pi2  & ~n359;
  assign n538 = ~n211 & ~n537;
  assign n539 = ~pi3  & ~pi6 ;
  assign n540 = ~n538 & n539;
  assign n541 = pi1  & ~n540;
  assign n542 = pi2  & ~n271;
  assign n543 = ~pi2  & pi5 ;
  assign n544 = pi8  & n543;
  assign n545 = pi5  & n279;
  assign n546 = ~pi2  & n503;
  assign n547 = ~n542 & ~n1122;
  assign n548 = ~pi9  & ~n547;
  assign n549 = pi5  & n212;
  assign n550 = ~pi8  & n497;
  assign n551 = ~pi3  & ~n1123;
  assign n552 = ~pi2  & ~n551;
  assign n553 = pi3  & ~pi5 ;
  assign n554 = ~pi6  & ~n312;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~n552 & ~n555;
  assign n557 = ~n548 & n556;
  assign n558 = pi1  & ~n557;
  assign n559 = ~n536 & n541;
  assign n560 = n268 & n302;
  assign n561 = ~n411 & ~n560;
  assign n562 = ~pi9  & ~n561;
  assign n563 = pi0  & ~n562;
  assign n564 = ~n1124 & n563;
  assign n565 = ~n531 & ~n564;
  assign n566 = pi3  & ~pi6 ;
  assign n567 = pi2  & n566;
  assign n568 = ~n65 & n410;
  assign n569 = ~n567 & ~n568;
  assign n570 = pi9  & ~n569;
  assign n571 = ~pi9  & n410;
  assign n572 = ~n566 & ~n571;
  assign n573 = ~pi8  & ~n572;
  assign n574 = ~n570 & ~n573;
  assign n575 = ~pi1  & ~n574;
  assign n576 = pi1  & n213;
  assign n577 = n410 & n576;
  assign n578 = pi1  & n410;
  assign n579 = n213 & n578;
  assign n580 = n417 & n571;
  assign n581 = ~n34 & ~n244;
  assign n582 = ~pi2  & ~n581;
  assign n583 = ~pi6  & ~n497;
  assign n584 = ~n386 & ~n503;
  assign n585 = n583 & ~n584;
  assign n586 = ~n582 & ~n585;
  assign n587 = pi3  & ~n586;
  assign n588 = ~n1125 & ~n587;
  assign n589 = ~n575 & n588;
  assign n590 = ~n1124 & ~n562;
  assign n591 = pi0  & ~n590;
  assign n592 = ~pi0  & n1121;
  assign n593 = n589 & ~n592;
  assign n594 = ~n591 & n593;
  assign n595 = ~n565 & n589;
  assign n596 = ~pi4  & ~n1126;
  assign n597 = n26 & n1112;
  assign n598 = ~pi1  & pi4 ;
  assign n599 = n1073 & n598;
  assign n600 = n1087 & n467;
  assign n601 = ~n180 & ~n489;
  assign n602 = ~pi5  & ~n211;
  assign n603 = n211 & n489;
  assign n604 = ~n180 & ~n603;
  assign n605 = ~n601 & ~n602;
  assign n606 = n467 & ~n601;
  assign n607 = n1087 & ~n602;
  assign n608 = n606 & n607;
  assign n609 = n1127 & ~n1128;
  assign n610 = ~pi4  & ~n1120;
  assign n611 = n1112 & ~n602;
  assign n612 = ~n601 & n611;
  assign n613 = n1112 & ~n1128;
  assign n614 = ~n610 & ~n1130;
  assign n615 = ~pi1  & ~n614;
  assign n616 = ~n1118 & ~n1119;
  assign n617 = ~pi4  & ~n616;
  assign n618 = ~n615 & ~n617;
  assign n619 = ~pi0  & ~n618;
  assign n620 = n589 & ~n591;
  assign n621 = ~pi4  & ~n620;
  assign n622 = ~n619 & ~n621;
  assign n623 = ~n596 & ~n1129;
  assign po3  = ~pi7  & ~n1131;
  assign n625 = ~n180 & ~n1127;
  assign n626 = ~pi7  & ~n625;
  assign n627 = pi7  & ~pi9 ;
  assign n628 = pi8  & ~n627;
  assign n629 = n129 & ~n628;
  assign n630 = ~n111 & ~n629;
  assign n631 = ~pi0  & ~n630;
  assign n632 = pi1  & n1081;
  assign n633 = n200 & n386;
  assign n634 = ~n171 & ~n1132;
  assign n635 = ~pi2  & pi7 ;
  assign n636 = pi7  & ~n634;
  assign n637 = ~pi2  & n636;
  assign n638 = ~n634 & n635;
  assign n639 = ~n631 & ~n1133;
  assign n640 = n348 & ~n639;
  assign n641 = ~pi1  & ~pi5 ;
  assign n642 = pi2  & ~n641;
  assign n643 = ~pi9  & ~n642;
  assign n644 = ~pi6  & n643;
  assign n645 = n167 & ~n642;
  assign n646 = pi5  & n386;
  assign n647 = ~n1134 & ~n646;
  assign n648 = pi0  & ~n647;
  assign n649 = ~pi0  & pi2 ;
  assign n650 = ~pi0  & ~n34;
  assign n651 = pi2  & n650;
  assign n652 = ~n34 & n649;
  assign n653 = ~n648 & ~n1135;
  assign n654 = pi8  & ~n653;
  assign n655 = pi2  & n41;
  assign n656 = pi9  & n649;
  assign n657 = ~n144 & ~n1136;
  assign n658 = pi5  & ~n657;
  assign n659 = ~pi2  & ~pi9 ;
  assign n660 = ~pi2  & pi9 ;
  assign n661 = ~n27 & ~n660;
  assign n662 = ~n110 & ~n659;
  assign n663 = pi2  & pi8 ;
  assign n664 = ~n197 & ~n663;
  assign n665 = pi6  & ~n664;
  assign n666 = pi6  & n1137;
  assign n667 = ~n664 & n666;
  assign n668 = pi6  & n1083;
  assign n669 = n1137 & n668;
  assign n670 = n1137 & n665;
  assign n671 = ~n658 & ~n1138;
  assign n672 = ~n654 & ~n658;
  assign n673 = ~n1138 & n672;
  assign n674 = ~n654 & n671;
  assign n675 = ~pi3  & ~n1139;
  assign n676 = pi8  & ~n281;
  assign n677 = ~pi0  & ~pi6 ;
  assign n678 = n659 & ~n677;
  assign n679 = ~pi8  & ~n677;
  assign n680 = ~n281 & ~n679;
  assign n681 = ~pi9  & ~n680;
  assign n682 = ~pi2  & n681;
  assign n683 = ~pi0  & ~n438;
  assign n684 = ~n503 & n659;
  assign n685 = ~n683 & n684;
  assign n686 = n659 & ~n680;
  assign n687 = ~n676 & n678;
  assign n688 = n41 & n663;
  assign n689 = ~pi1  & ~n688;
  assign n690 = ~n1140 & n689;
  assign n691 = ~n1066 & n543;
  assign n692 = ~pi6  & ~n405;
  assign n693 = n41 & ~n692;
  assign n694 = ~n691 & ~n693;
  assign n695 = ~pi8  & ~n694;
  assign n696 = pi2  & ~n171;
  assign n697 = ~n1081 & ~n696;
  assign n698 = pi6  & ~n697;
  assign n699 = pi1  & ~n698;
  assign n700 = ~n695 & n699;
  assign n701 = ~n695 & ~n698;
  assign n702 = pi1  & ~n701;
  assign n703 = ~n1140 & ~n688;
  assign n704 = ~pi1  & ~n703;
  assign n705 = ~n702 & ~n704;
  assign n706 = ~n690 & ~n700;
  assign n707 = ~pi1  & ~n171;
  assign n708 = pi0  & ~n51;
  assign n709 = pi0  & ~n707;
  assign n710 = ~n51 & n709;
  assign n711 = ~n144 & ~n386;
  assign n712 = pi0  & ~n711;
  assign n713 = ~n707 & n708;
  assign n714 = ~n290 & n677;
  assign n715 = ~n59 & ~n714;
  assign n716 = pi2  & n51;
  assign n717 = ~n290 & n387;
  assign n718 = n677 & n717;
  assign n719 = n387 & n714;
  assign n720 = ~n716 & ~n1143;
  assign n721 = n387 & ~n715;
  assign n722 = ~n1142 & ~n716;
  assign n723 = ~n1143 & n722;
  assign n724 = ~n1142 & n1144;
  assign n725 = ~pi5  & ~n1145;
  assign n726 = pi0  & n237;
  assign n727 = ~pi2  & n726;
  assign n728 = n134 & ~n649;
  assign n729 = ~pi8  & n301;
  assign n730 = ~n134 & ~n726;
  assign n731 = ~pi2  & ~n730;
  assign n732 = ~n729 & ~n731;
  assign n733 = ~n727 & ~n728;
  assign n734 = ~n134 & ~n727;
  assign n735 = pi9  & ~n649;
  assign n736 = ~n734 & n735;
  assign n737 = pi9  & ~n1146;
  assign n738 = ~pi0  & ~pi8 ;
  assign n739 = n51 & ~n281;
  assign n740 = ~n281 & ~n738;
  assign n741 = n51 & n740;
  assign n742 = ~n738 & n739;
  assign n743 = ~n1147 & ~n1148;
  assign n744 = ~n725 & ~n1148;
  assign n745 = ~n1147 & n744;
  assign n746 = ~n725 & n743;
  assign n747 = pi3  & ~n1149;
  assign n748 = n1141 & ~n747;
  assign n749 = ~n675 & n748;
  assign n750 = ~pi7  & ~n749;
  assign n751 = ~pi7  & ~n1139;
  assign n752 = n489 & ~n639;
  assign n753 = ~n751 & ~n752;
  assign n754 = ~pi3  & ~n753;
  assign n755 = ~pi7  & ~n748;
  assign n756 = ~n754 & ~n755;
  assign n757 = ~n640 & ~n750;
  assign n758 = ~pi4  & ~n1150;
  assign po6  = ~n626 & ~n758;
  assign n760 = n299 & n566;
  assign n761 = ~n438 & ~n760;
  assign n762 = pi9  & ~n761;
  assign n763 = ~pi8  & ~n208;
  assign n764 = pi0  & ~n566;
  assign n765 = ~n177 & ~n764;
  assign n766 = ~pi3  & pi8 ;
  assign n767 = ~n208 & ~n766;
  assign n768 = pi0  & ~n767;
  assign n769 = ~pi9  & n237;
  assign n770 = ~n768 & ~n769;
  assign n771 = ~n763 & ~n765;
  assign n772 = ~n762 & ~n769;
  assign n773 = ~n768 & n772;
  assign n774 = ~n762 & n1151;
  assign n775 = ~pi2  & ~n1152;
  assign n776 = ~pi3  & n172;
  assign n777 = n167 & n269;
  assign n778 = pi3  & ~n211;
  assign n779 = ~n200 & ~n778;
  assign n780 = ~pi6  & ~n779;
  assign n781 = ~pi3  & n211;
  assign n782 = ~n780 & ~n781;
  assign n783 = pi2  & ~n782;
  assign n784 = ~n1153 & ~n783;
  assign n785 = ~n775 & ~n1153;
  assign n786 = ~n783 & n785;
  assign n787 = ~n775 & n784;
  assign n788 = pi1  & ~n1154;
  assign n789 = ~pi0  & n668;
  assign n790 = n1083 & n245;
  assign n791 = ~pi6  & ~n211;
  assign n792 = ~n84 & ~n212;
  assign n793 = ~pi6  & ~n792;
  assign n794 = ~pi2  & n793;
  assign n795 = ~pi2  & ~pi6 ;
  assign n796 = ~n792 & n795;
  assign n797 = n98 & n791;
  assign n798 = ~n1155 & ~n1156;
  assign n799 = pi3  & ~n798;
  assign n800 = ~pi0  & n197;
  assign n801 = ~n726 & ~n800;
  assign n802 = ~pi9  & ~n801;
  assign n803 = ~pi6  & ~n269;
  assign n804 = n696 & ~n803;
  assign n805 = ~n802 & ~n804;
  assign n806 = ~n799 & n805;
  assign n807 = ~pi1  & ~n806;
  assign n808 = pi6  & n197;
  assign n809 = ~pi8  & n122;
  assign n810 = pi3  & n197;
  assign n811 = n177 & n810;
  assign n812 = ~pi2  & pi3 ;
  assign n813 = ~pi9  & n438;
  assign n814 = n812 & n813;
  assign n815 = n516 & n1157;
  assign n816 = ~n807 & ~n1158;
  assign n817 = ~n788 & n816;
  assign n818 = ~pi5  & ~n817;
  assign n819 = pi0  & ~n1137;
  assign n820 = pi5  & ~pi9 ;
  assign n821 = ~pi0  & n820;
  assign n822 = ~pi9  & n56;
  assign n823 = ~n819 & ~n1159;
  assign n824 = pi8  & ~n823;
  assign n825 = pi2  & n1123;
  assign n826 = n110 & n216;
  assign n827 = ~n824 & ~n1160;
  assign n828 = ~pi3  & ~n827;
  assign n829 = pi3  & pi5 ;
  assign n830 = ~n27 & ~n829;
  assign n831 = pi2  & ~n738;
  assign n832 = ~n211 & ~n831;
  assign n833 = pi3  & n543;
  assign n834 = n738 & ~n830;
  assign n835 = ~n833 & ~n834;
  assign n836 = ~n211 & ~n835;
  assign n837 = ~pi0  & ~n830;
  assign n838 = ~n833 & ~n837;
  assign n839 = ~pi8  & ~n838;
  assign n840 = n812 & n820;
  assign n841 = ~n839 & ~n840;
  assign n842 = ~n830 & n832;
  assign n843 = ~n828 & ~n1161;
  assign n844 = pi1  & ~n843;
  assign n845 = n67 & n395;
  assign n846 = pi2  & pi3 ;
  assign n847 = ~n1083 & ~n846;
  assign n848 = ~pi2  & ~n67;
  assign n849 = pi5  & ~n848;
  assign n850 = n1083 & ~n848;
  assign n851 = ~n846 & ~n850;
  assign n852 = pi5  & ~n851;
  assign n853 = ~n847 & n849;
  assign n854 = ~n845 & ~n1162;
  assign n855 = ~pi1  & ~n854;
  assign n856 = pi8  & n497;
  assign n857 = n846 & n856;
  assign n858 = ~n855 & ~n857;
  assign n859 = ~n844 & n858;
  assign n860 = ~pi6  & ~n859;
  assign n861 = ~n818 & ~n860;
  assign n862 = ~pi7  & ~n861;
  assign n863 = pi2  & ~n1083;
  assign n864 = ~pi0  & n863;
  assign n865 = ~n1083 & n649;
  assign n866 = ~pi9  & n23;
  assign n867 = n37 & n866;
  assign n868 = n280 & n627;
  assign n869 = ~n1163 & ~n1164;
  assign n870 = n186 & n489;
  assign n871 = n43 & n302;
  assign n872 = n302 & ~n869;
  assign n873 = n43 & n872;
  assign n874 = ~n869 & n1165;
  assign n875 = ~n862 & ~n1166;
  assign n876 = ~pi4  & ~n875;
  assign n877 = n60 & n113;
  assign n878 = pi4  & ~pi7 ;
  assign n879 = n302 & n878;
  assign n880 = n43 & n878;
  assign n881 = ~pi5  & ~pi7 ;
  assign n882 = n1127 & n881;
  assign n883 = n1087 & n880;
  assign n884 = ~pi6  & n1167;
  assign n885 = n877 & n879;
  assign po7  = ~n876 & ~n1168;
  assign n887 = ~pi1  & pi5 ;
  assign n888 = ~n43 & ~n887;
  assign n889 = ~pi2  & ~n113;
  assign n890 = ~pi2  & ~n88;
  assign n891 = ~n553 & n890;
  assign n892 = ~n113 & n891;
  assign n893 = ~n113 & ~n888;
  assign n894 = ~pi2  & n893;
  assign n895 = ~n888 & n889;
  assign n896 = n186 & n281;
  assign n897 = n43 & n57;
  assign n898 = ~n1169 & ~n1170;
  assign n899 = pi8  & ~n898;
  assign n900 = ~pi5  & ~n299;
  assign n901 = n59 & ~n829;
  assign n902 = ~n829 & ~n900;
  assign n903 = n59 & n902;
  assign n904 = ~n900 & n901;
  assign n905 = ~n899 & ~n1171;
  assign n906 = ~pi9  & ~n905;
  assign n907 = ~n405 & ~n829;
  assign n908 = pi1  & ~n403;
  assign n909 = ~n403 & ~n907;
  assign n910 = pi1  & n909;
  assign n911 = ~n907 & n908;
  assign n912 = ~n56 & n279;
  assign n913 = ~n56 & n311;
  assign n914 = n279 & n913;
  assign n915 = n311 & n912;
  assign n916 = ~n1172 & ~n1173;
  assign n917 = pi9  & ~n916;
  assign n918 = ~n121 & ~n433;
  assign n919 = ~n888 & n918;
  assign n920 = ~pi2  & n919;
  assign n921 = ~pi2  & ~n121;
  assign n922 = ~n433 & n921;
  assign n923 = ~n888 & n922;
  assign n924 = n891 & n918;
  assign n925 = n387 & ~n641;
  assign n926 = n135 & ~n925;
  assign n927 = n260 & n820;
  assign n928 = n121 & n543;
  assign n929 = ~n439 & ~n1175;
  assign n930 = ~pi0  & ~n929;
  assign n931 = ~n926 & ~n930;
  assign n932 = ~n1174 & ~n926;
  assign n933 = ~n930 & n932;
  assign n934 = ~n1174 & ~n930;
  assign n935 = ~n926 & n934;
  assign n936 = ~n1174 & n931;
  assign n937 = ~pi8  & ~n1176;
  assign n938 = ~n917 & ~n937;
  assign n939 = ~n906 & ~n917;
  assign n940 = ~n937 & n939;
  assign n941 = ~n906 & n938;
  assign n942 = ~pi6  & ~n1177;
  assign n943 = ~n51 & n299;
  assign n944 = n383 & ~n943;
  assign n945 = ~pi2  & ~n944;
  assign n946 = ~pi6  & ~n134;
  assign n947 = ~n709 & n946;
  assign n948 = n553 & ~n947;
  assign n949 = pi2  & ~n707;
  assign n950 = ~n383 & ~n949;
  assign n951 = pi0  & ~n950;
  assign n952 = pi2  & ~n946;
  assign n953 = pi8  & ~n51;
  assign n954 = pi6  & ~n211;
  assign n955 = ~n707 & n954;
  assign n956 = n383 & ~n953;
  assign n957 = ~n952 & ~n1178;
  assign n958 = ~n951 & n957;
  assign n959 = n553 & ~n958;
  assign n960 = ~n945 & n948;
  assign n961 = ~n942 & ~n1179;
  assign n962 = ~pi7  & ~n961;
  assign n963 = ~pi0  & ~n664;
  assign n964 = ~n280 & ~n963;
  assign n965 = ~pi9  & ~n964;
  assign n966 = ~pi8  & n1136;
  assign n967 = n110 & n738;
  assign n968 = ~n965 & ~n1180;
  assign n969 = ~pi1  & ~n968;
  assign n970 = n386 & n800;
  assign n971 = ~n969 & ~n970;
  assign n972 = n43 & ~n971;
  assign n973 = ~pi6  & n972;
  assign n974 = n348 & ~n971;
  assign n975 = ~n962 & ~n1181;
  assign n976 = ~pi4  & ~n975;
  assign po8  = ~n1167 & ~n976;
  assign n978 = pi3  & ~n208;
  assign n979 = n299 & ~n583;
  assign n980 = n978 & ~n979;
  assign n981 = n467 & ~n489;
  assign n982 = ~pi2  & ~n981;
  assign n983 = ~n208 & ~n979;
  assign n984 = pi3  & ~n983;
  assign n985 = pi4  & ~n489;
  assign n986 = ~pi3  & ~n985;
  assign n987 = ~n984 & ~n986;
  assign n988 = ~pi2  & ~n987;
  assign n989 = ~n980 & n982;
  assign n990 = n135 & ~n171;
  assign n991 = ~pi3  & ~n602;
  assign n992 = n696 & n991;
  assign n993 = ~pi3  & ~n34;
  assign n994 = ~pi8  & ~n497;
  assign n995 = n993 & ~n994;
  assign n996 = pi2  & n995;
  assign n997 = pi2  & n993;
  assign n998 = ~n994 & n997;
  assign n999 = ~n602 & n990;
  assign n1000 = ~n1182 & ~n1183;
  assign n1001 = ~pi1  & ~n1000;
  assign n1002 = n299 & ~n978;
  assign n1003 = ~n993 & ~n1002;
  assign n1004 = ~pi2  & ~n1003;
  assign n1005 = ~n211 & n567;
  assign n1006 = ~pi5  & n1005;
  assign n1007 = n567 & n602;
  assign n1008 = ~pi6  & ~n856;
  assign n1009 = ~pi3  & ~n1008;
  assign n1010 = ~n1184 & ~n1009;
  assign n1011 = ~n1004 & n1010;
  assign n1012 = pi1  & ~n1011;
  assign n1013 = n281 & n567;
  assign n1014 = ~pi7  & ~n1013;
  assign n1015 = ~n707 & ~n1014;
  assign n1016 = ~pi7  & ~n188;
  assign n1017 = pi0  & ~n1016;
  assign n1018 = ~pi5  & ~n135;
  assign n1019 = pi6  & ~n1018;
  assign n1020 = pi4  & ~n188;
  assign n1021 = pi7  & ~n135;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n1019 & n1022;
  assign n1024 = ~n1017 & n1023;
  assign n1025 = ~n1015 & n1024;
  assign n1026 = ~n1012 & n1025;
  assign n1027 = ~n1001 & ~n1019;
  assign n1028 = ~n1012 & n1027;
  assign n1029 = ~n1021 & n1028;
  assign n1030 = ~n1017 & n1029;
  assign n1031 = ~n1015 & n1030;
  assign n1032 = ~n1020 & n1031;
  assign n1033 = ~n1001 & n1026;
  assign n1034 = pi8  & ~n42;
  assign n1035 = pi3  & ~pi4 ;
  assign n1036 = pi2  & n1035;
  assign n1037 = ~n50 & n1036;
  assign n1038 = ~pi8  & ~n50;
  assign n1039 = ~n42 & ~n1038;
  assign n1040 = n1035 & ~n1039;
  assign n1041 = pi2  & n1040;
  assign n1042 = n1036 & ~n1039;
  assign n1043 = ~n1034 & n1037;
  assign n1044 = ~n1127 & ~n1186;
  assign n1045 = ~pi7  & n489;
  assign n1046 = ~pi7  & ~n1044;
  assign n1047 = n489 & n1046;
  assign n1048 = ~n1044 & n1045;
  assign n1049 = ~pi4  & n339;
  assign n1050 = ~n467 & ~n1035;
  assign n1051 = n1087 & ~n1050;
  assign n1052 = ~n1049 & ~n1051;
  assign n1053 = ~pi7  & n180;
  assign n1054 = ~pi7  & ~n1052;
  assign n1055 = n180 & n1054;
  assign n1056 = ~n1052 & n1053;
  assign n1057 = ~n1087 & n1035;
  assign n1058 = ~n1127 & ~n1057;
  assign n1059 = ~pi7  & ~n1058;
  assign n1060 = n180 & n1059;
  assign n1061 = n1053 & ~n1058;
  assign n1062 = n24 | n25;
  assign n1063 = n47 | n48;
  assign n1064 = n62 | n63;
  assign n1065 = n73 | n74;
  assign n1066 = n86 | ~n87;
  assign n1067 = n95 | n92 | n94;
  assign n1068 = n105 | n106;
  assign n1069 = n108 | n109;
  assign n1070 = n116 | n117;
  assign n1071 = n130 | n131;
  assign n1072 = n141 | n142;
  assign n1073 = n145 | n146;
  assign n1074 = n157 | n158;
  assign n1075 = n162 | n159 | n161;
  assign n1076 = n175 | n176;
  assign n1077 = n183 | n184;
  assign n1078 = n190 | n191;
  assign n1079 = n194 | n195;
  assign n1080 = n198 | n199;
  assign n1081 = n201 | n202;
  assign n1082 = n203 | n204;
  assign n1083 = n214 | ~n215;
  assign n1084 = n221 | ~n222;
  assign n1085 = n232 | n233;
  assign n1086 = n240 | n241;
  assign n1087 = n262 | n259 | n261;
  assign n1088 = n265 | n266;
  assign n1089 = n272 | n273;
  assign n1090 = n295 | ~n296;
  assign n1091 = n297 | n298;
  assign n1092 = n305 | n306;
  assign n1093 = n313 | n314;
  assign n1094 = n320 | ~n321;
  assign n1095 = n333 | n334;
  assign n1096 = n342 | n343;
  assign n1097 = n349 | n350;
  assign n1098 = n353 | n354;
  assign n1099 = n356 | n357;
  assign n1100 = n360 | ~n361;
  assign n1101 = n362 | n363;
  assign n1102 = n367 | n368;
  assign n1103 = n371 | n372;
  assign n1104 = n413 | n414;
  assign n1105 = n421 | n422;
  assign n1106 = n430 | n431;
  assign n1107 = n436 | n437;
  assign n1108 = n443 | n444;
  assign n1109 = n449 | ~n450;
  assign n1110 = n454 | n451 | n453;
  assign n1111 = n464 | n465;
  assign n1112 = n468 | n469;
  assign n1113 = n470 | n471;
  assign n1114 = n474 | n475;
  assign n1115 = n477 | n478;
  assign n1116 = n485 | n486;
  assign n1117 = n494 | n495;
  assign n1118 = n510 | n511;
  assign n1119 = n512 | n513;
  assign n1120 = n518 | n519;
  assign n1121 = n529 | ~n530;
  assign n1122 = n546 | n544 | n545;
  assign n1123 = n549 | n550;
  assign n1124 = n558 | n559;
  assign n1125 = n580 | n577 | n579;
  assign n1126 = n594 | n595;
  assign n1127 = n600 | n597 | n599;
  assign n1128 = n604 | ~n605;
  assign n1129 = n608 | n609;
  assign n1130 = n612 | n613;
  assign n1131 = n622 | n623;
  assign n1132 = n632 | n633;
  assign n1133 = n637 | n638;
  assign n1134 = n644 | n645;
  assign n1135 = n651 | n652;
  assign n1136 = n655 | n656;
  assign n1137 = n661 | ~n662;
  assign n1138 = n670 | n667 | n669;
  assign n1139 = n673 | n674;
  assign n1140 = n682 | n685 | n686 | n687;
  assign n1141 = n705 | ~n706;
  assign n1142 = n713 | n710 | n712;
  assign n1143 = n718 | n719;
  assign n1144 = n720 | ~n721;
  assign n1145 = n723 | n724;
  assign n1146 = n732 | n733;
  assign n1147 = n736 | n737;
  assign n1148 = n741 | n742;
  assign n1149 = n745 | n746;
  assign n1150 = n756 | n757;
  assign n1151 = n770 | ~n771;
  assign n1152 = n773 | n774;
  assign n1153 = n776 | n777;
  assign n1154 = n786 | n787;
  assign n1155 = n789 | n790;
  assign n1156 = n797 | n794 | n796;
  assign n1157 = n808 | n809;
  assign n1158 = n815 | n811 | n814;
  assign n1159 = n821 | n822;
  assign n1160 = n825 | n826;
  assign n1161 = n842 | n836 | ~n841;
  assign n1162 = n852 | n853;
  assign n1163 = n864 | n865;
  assign n1164 = n867 | n868;
  assign n1165 = n870 | n871;
  assign n1166 = n873 | n874;
  assign n1167 = n882 | n883;
  assign n1168 = n884 | n885;
  assign n1169 = n895 | n892 | n894;
  assign n1170 = n896 | n897;
  assign n1171 = n903 | n904;
  assign n1172 = n910 | n911;
  assign n1173 = n914 | n915;
  assign n1174 = n924 | n920 | n923;
  assign n1175 = n927 | n928;
  assign n1176 = n936 | n933 | n935;
  assign n1177 = n940 | n941;
  assign n1178 = n955 | n956;
  assign n1179 = n959 | n960;
  assign n1180 = n966 | n967;
  assign n1181 = n973 | n974;
  assign n1182 = n988 | n989;
  assign n1183 = n992 | n996 | n998 | n999;
  assign n1184 = n1006 | n1007;
  assign po9  = n1032 | n1033;
  assign n1186 = n1043 | n1041 | n1042;
  assign po10  = n1047 | n1048;
  assign po4  = n1055 | n1056;
  assign po5  = n1060 | n1061;
  assign po0  = ~n196;
  assign po1  = ~n355;
  assign po2  = ~n496;
endmodule
