module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 ,
    pi131 , pi132 , pi133 , pi134 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 ,
    pi130 , pi131 , pi132 , pi133 , pi134 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ;
  wire n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n635,
    n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108,
    n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168,
    n1169, n1170, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361,
    n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391,
    n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421,
    n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451,
    n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542,
    n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1813, n1814, n1815, n1816,
    n1817, n1818, n1819, n1820, n1821, n1822,
    n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834,
    n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852,
    n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882,
    n1883, n1884, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901,
    n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931,
    n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1959, n1960, n1961, n1962,
    n1963, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1992,
    n1993, n1994, n1995, n1996, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016,
    n2017, n2018, n2019, n2020, n2021, n2022,
    n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101,
    n2102, n2103, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2251, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266,
    n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278,
    n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296,
    n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2324, n2325, n2326, n2327,
    n2328, n2329, n2330, n2331, n2332, n2333,
    n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351,
    n2352, n2353, n2354, n2355, n2356, n2357,
    n2358, n2359, n2360, n2361, n2362, n2363,
    n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381,
    n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393,
    n2394, n2395, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412,
    n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2479, n2480, n2482, n2483,
    n2484, n2485, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514,
    n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2567, n2568, n2569, n2570, n2571, n2572,
    n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597,
    n2598, n2599, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616,
    n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2693,
    n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718,
    n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731,
    n2732, n2733, n2734, n2735, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801,
    n2802, n2803, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820,
    n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2837, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884,
    n2885, n2886, n2887, n2888, n2890, n2891,
    n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922,
    n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986,
    n2987, n2988, n2989, n2990, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3007, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024,
    n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075,
    n3077, n3078, n3079, n3080, n3081, n3082,
    n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101,
    n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3109, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177,
    n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3186, n3187, n3188, n3189, n3190,
    n3191, n3192, n3193, n3194, n3196, n3197,
    n3198, n3199, n3200, n3201, n3202, n3203,
    n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3213, n3214, n3216, n3217,
    n3219, n3220, n3222, n3223, n3225, n3226,
    n3228, n3229, n3231, n3232, n3234, n3235,
    n3237, n3238, n3240, n3241, n3243, n3244,
    n3246, n3247, n3249, n3250, n3252, n3253,
    n3255, n3256, n3258, n3259, n3261, n3262,
    n3264, n3265, n3267, n3268, n3270, n3271,
    n3273, n3274, n3276, n3277, n3279, n3280,
    n3282, n3283, n3285, n3286, n3288, n3289,
    n3291, n3292, n3294, n3295, n3297, n3298,
    n3300, n3301, n3303, n3304, n3306, n3307,
    n3309, n3310, n3312, n3313, n3315, n3316,
    n3318, n3319, n3321, n3322, n3324, n3325,
    n3327, n3328, n3330, n3331, n3333, n3334,
    n3336, n3337, n3339, n3340, n3342, n3343,
    n3345, n3346, n3348, n3349, n3351, n3352,
    n3354, n3355, n3357, n3358, n3360, n3361,
    n3363, n3364, n3366, n3367, n3369, n3370,
    n3372, n3373, n3375, n3376, n3378, n3379,
    n3381, n3382, n3384, n3385, n3387, n3388,
    n3390, n3391, n3393, n3394, n3396, n3397,
    n3399, n3400, n3402, n3403;
  assign n264 = pi77  & pi128 ;
  assign n265 = pi78  & ~pi128 ;
  assign n266 = ~n264 & ~n265;
  assign n267 = pi129  & ~n266;
  assign n268 = pi80  & ~pi128 ;
  assign n269 = pi79  & pi128 ;
  assign n270 = ~n268 & ~n269;
  assign n271 = ~pi129  & ~n270;
  assign n272 = ~n267 & ~n271;
  assign n273 = ~pi130  & ~pi131 ;
  assign n274 = ~n272 & n273;
  assign n275 = pi73  & pi128 ;
  assign n276 = pi74  & ~pi128 ;
  assign n277 = ~n275 & ~n276;
  assign n278 = pi129  & ~n277;
  assign n279 = pi76  & ~pi128 ;
  assign n280 = pi75  & pi128 ;
  assign n281 = ~n279 & ~n280;
  assign n282 = ~pi129  & ~n281;
  assign n283 = ~n278 & ~n282;
  assign n284 = pi130  & ~pi131 ;
  assign n285 = ~n283 & n284;
  assign n286 = ~n274 & ~n285;
  assign n287 = pi65  & pi128 ;
  assign n288 = pi66  & ~pi128 ;
  assign n289 = ~n287 & ~n288;
  assign n290 = pi129  & ~n289;
  assign n291 = pi68  & ~pi128 ;
  assign n292 = pi67  & pi128 ;
  assign n293 = ~n291 & ~n292;
  assign n294 = ~pi129  & ~n293;
  assign n295 = ~n290 & ~n294;
  assign n296 = pi130  & pi131 ;
  assign n297 = ~n295 & n296;
  assign n298 = pi69  & pi128 ;
  assign n299 = pi70  & ~pi128 ;
  assign n300 = ~n298 & ~n299;
  assign n301 = pi129  & ~n300;
  assign n302 = pi72  & ~pi128 ;
  assign n303 = pi71  & pi128 ;
  assign n304 = ~n302 & ~n303;
  assign n305 = ~pi129  & ~n304;
  assign n306 = ~n301 & ~n305;
  assign n307 = ~pi130  & pi131 ;
  assign n308 = ~n306 & n307;
  assign n309 = ~n297 & ~n308;
  assign n310 = n286 & n309;
  assign n311 = pi132  & pi133 ;
  assign n312 = ~n310 & n311;
  assign n313 = pi93  & pi128 ;
  assign n314 = pi94  & ~pi128 ;
  assign n315 = ~n313 & ~n314;
  assign n316 = pi129  & ~n315;
  assign n317 = pi96  & ~pi128 ;
  assign n318 = pi95  & pi128 ;
  assign n319 = ~n317 & ~n318;
  assign n320 = ~pi129  & ~n319;
  assign n321 = ~n316 & ~n320;
  assign n322 = n273 & ~n321;
  assign n323 = pi89  & pi128 ;
  assign n324 = pi90  & ~pi128 ;
  assign n325 = ~n323 & ~n324;
  assign n326 = pi129  & ~n325;
  assign n327 = pi92  & ~pi128 ;
  assign n328 = pi91  & pi128 ;
  assign n329 = ~n327 & ~n328;
  assign n330 = ~pi129  & ~n329;
  assign n331 = ~n326 & ~n330;
  assign n332 = n284 & ~n331;
  assign n333 = ~n322 & ~n332;
  assign n334 = pi81  & pi128 ;
  assign n335 = pi82  & ~pi128 ;
  assign n336 = ~n334 & ~n335;
  assign n337 = pi129  & ~n336;
  assign n338 = pi84  & ~pi128 ;
  assign n339 = pi83  & pi128 ;
  assign n340 = ~n338 & ~n339;
  assign n341 = ~pi129  & ~n340;
  assign n342 = ~n337 & ~n341;
  assign n343 = n296 & ~n342;
  assign n344 = pi85  & pi128 ;
  assign n345 = pi86  & ~pi128 ;
  assign n346 = ~n344 & ~n345;
  assign n347 = pi129  & ~n346;
  assign n348 = pi88  & ~pi128 ;
  assign n349 = pi87  & pi128 ;
  assign n350 = ~n348 & ~n349;
  assign n351 = ~pi129  & ~n350;
  assign n352 = ~n347 & ~n351;
  assign n353 = n307 & ~n352;
  assign n354 = ~n343 & ~n353;
  assign n355 = n333 & n354;
  assign n356 = ~pi132  & pi133 ;
  assign n357 = ~n355 & n356;
  assign n358 = ~n312 & ~n357;
  assign n359 = pi125  & pi128 ;
  assign n360 = pi126  & ~pi128 ;
  assign n361 = ~n359 & ~n360;
  assign n362 = pi129  & ~n361;
  assign n363 = pi0  & ~pi128 ;
  assign n364 = pi127  & pi128 ;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~pi129  & ~n365;
  assign n367 = ~n362 & ~n366;
  assign n368 = n273 & ~n367;
  assign n369 = pi121  & pi128 ;
  assign n370 = pi122  & ~pi128 ;
  assign n371 = ~n369 & ~n370;
  assign n372 = pi129  & ~n371;
  assign n373 = pi124  & ~pi128 ;
  assign n374 = pi123  & pi128 ;
  assign n375 = ~n373 & ~n374;
  assign n376 = ~pi129  & ~n375;
  assign n377 = ~n372 & ~n376;
  assign n378 = n284 & ~n377;
  assign n379 = ~n368 & ~n378;
  assign n380 = pi113  & pi128 ;
  assign n381 = pi114  & ~pi128 ;
  assign n382 = ~n380 & ~n381;
  assign n383 = pi129  & ~n382;
  assign n384 = pi116  & ~pi128 ;
  assign n385 = pi115  & pi128 ;
  assign n386 = ~n384 & ~n385;
  assign n387 = ~pi129  & ~n386;
  assign n388 = ~n383 & ~n387;
  assign n389 = n296 & ~n388;
  assign n390 = pi117  & pi128 ;
  assign n391 = pi118  & ~pi128 ;
  assign n392 = ~n390 & ~n391;
  assign n393 = pi129  & ~n392;
  assign n394 = pi120  & ~pi128 ;
  assign n395 = pi119  & pi128 ;
  assign n396 = ~n394 & ~n395;
  assign n397 = ~pi129  & ~n396;
  assign n398 = ~n393 & ~n397;
  assign n399 = n307 & ~n398;
  assign n400 = ~n389 & ~n399;
  assign n401 = n379 & n400;
  assign n402 = ~pi132  & ~pi133 ;
  assign n403 = ~n401 & n402;
  assign n404 = pi109  & pi128 ;
  assign n405 = pi110  & ~pi128 ;
  assign n406 = ~n404 & ~n405;
  assign n407 = pi129  & ~n406;
  assign n408 = pi112  & ~pi128 ;
  assign n409 = pi111  & pi128 ;
  assign n410 = ~n408 & ~n409;
  assign n411 = ~pi129  & ~n410;
  assign n412 = ~n407 & ~n411;
  assign n413 = n273 & ~n412;
  assign n414 = pi105  & pi128 ;
  assign n415 = pi106  & ~pi128 ;
  assign n416 = ~n414 & ~n415;
  assign n417 = pi129  & ~n416;
  assign n418 = pi108  & ~pi128 ;
  assign n419 = pi107  & pi128 ;
  assign n420 = ~n418 & ~n419;
  assign n421 = ~pi129  & ~n420;
  assign n422 = ~n417 & ~n421;
  assign n423 = n284 & ~n422;
  assign n424 = ~n413 & ~n423;
  assign n425 = pi97  & pi128 ;
  assign n426 = pi98  & ~pi128 ;
  assign n427 = ~n425 & ~n426;
  assign n428 = pi129  & ~n427;
  assign n429 = pi100  & ~pi128 ;
  assign n430 = pi99  & pi128 ;
  assign n431 = ~n429 & ~n430;
  assign n432 = ~pi129  & ~n431;
  assign n433 = ~n428 & ~n432;
  assign n434 = n296 & ~n433;
  assign n435 = pi101  & pi128 ;
  assign n436 = pi102  & ~pi128 ;
  assign n437 = ~n435 & ~n436;
  assign n438 = pi129  & ~n437;
  assign n439 = pi104  & ~pi128 ;
  assign n440 = pi103  & pi128 ;
  assign n441 = ~n439 & ~n440;
  assign n442 = ~pi129  & ~n441;
  assign n443 = ~n438 & ~n442;
  assign n444 = n307 & ~n443;
  assign n445 = ~n434 & ~n444;
  assign n446 = n424 & n445;
  assign n447 = pi132  & ~pi133 ;
  assign n448 = ~n446 & n447;
  assign n449 = ~n403 & ~n448;
  assign n450 = n358 & n449;
  assign n451 = ~pi134  & ~n450;
  assign n452 = pi13  & pi128 ;
  assign n453 = pi14  & ~pi128 ;
  assign n454 = ~n452 & ~n453;
  assign n455 = pi129  & ~n454;
  assign n456 = pi16  & ~pi128 ;
  assign n457 = pi15  & pi128 ;
  assign n458 = ~n456 & ~n457;
  assign n459 = ~pi129  & ~n458;
  assign n460 = ~n455 & ~n459;
  assign n461 = n273 & ~n460;
  assign n462 = pi9  & pi128 ;
  assign n463 = pi10  & ~pi128 ;
  assign n464 = ~n462 & ~n463;
  assign n465 = pi129  & ~n464;
  assign n466 = pi12  & ~pi128 ;
  assign n467 = pi11  & pi128 ;
  assign n468 = ~n466 & ~n467;
  assign n469 = ~pi129  & ~n468;
  assign n470 = ~n465 & ~n469;
  assign n471 = n284 & ~n470;
  assign n472 = ~n461 & ~n471;
  assign n473 = pi1  & pi128 ;
  assign n474 = pi2  & ~pi128 ;
  assign n475 = ~n473 & ~n474;
  assign n476 = pi129  & ~n475;
  assign n477 = pi4  & ~pi128 ;
  assign n478 = pi3  & pi128 ;
  assign n479 = ~n477 & ~n478;
  assign n480 = ~pi129  & ~n479;
  assign n481 = ~n476 & ~n480;
  assign n482 = n296 & ~n481;
  assign n483 = pi5  & pi128 ;
  assign n484 = pi6  & ~pi128 ;
  assign n485 = ~n483 & ~n484;
  assign n486 = pi129  & ~n485;
  assign n487 = pi8  & ~pi128 ;
  assign n488 = pi7  & pi128 ;
  assign n489 = ~n487 & ~n488;
  assign n490 = ~pi129  & ~n489;
  assign n491 = ~n486 & ~n490;
  assign n492 = n307 & ~n491;
  assign n493 = ~n482 & ~n492;
  assign n494 = n472 & n493;
  assign n495 = n311 & ~n494;
  assign n496 = pi29  & pi128 ;
  assign n497 = pi30  & ~pi128 ;
  assign n498 = ~n496 & ~n497;
  assign n499 = pi129  & ~n498;
  assign n500 = pi32  & ~pi128 ;
  assign n501 = pi31  & pi128 ;
  assign n502 = ~n500 & ~n501;
  assign n503 = ~pi129  & ~n502;
  assign n504 = ~n499 & ~n503;
  assign n505 = n273 & ~n504;
  assign n506 = pi25  & pi128 ;
  assign n507 = pi26  & ~pi128 ;
  assign n508 = ~n506 & ~n507;
  assign n509 = pi129  & ~n508;
  assign n510 = pi28  & ~pi128 ;
  assign n511 = pi27  & pi128 ;
  assign n512 = ~n510 & ~n511;
  assign n513 = ~pi129  & ~n512;
  assign n514 = ~n509 & ~n513;
  assign n515 = n284 & ~n514;
  assign n516 = ~n505 & ~n515;
  assign n517 = pi17  & pi128 ;
  assign n518 = pi18  & ~pi128 ;
  assign n519 = ~n517 & ~n518;
  assign n520 = pi129  & ~n519;
  assign n521 = pi20  & ~pi128 ;
  assign n522 = pi19  & pi128 ;
  assign n523 = ~n521 & ~n522;
  assign n524 = ~pi129  & ~n523;
  assign n525 = ~n520 & ~n524;
  assign n526 = n296 & ~n525;
  assign n527 = pi21  & pi128 ;
  assign n528 = pi22  & ~pi128 ;
  assign n529 = ~n527 & ~n528;
  assign n530 = pi129  & ~n529;
  assign n531 = pi24  & ~pi128 ;
  assign n532 = pi23  & pi128 ;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~pi129  & ~n533;
  assign n535 = ~n530 & ~n534;
  assign n536 = n307 & ~n535;
  assign n537 = ~n526 & ~n536;
  assign n538 = n516 & n537;
  assign n539 = n356 & ~n538;
  assign n540 = ~n495 & ~n539;
  assign n541 = pi61  & pi128 ;
  assign n542 = pi62  & ~pi128 ;
  assign n543 = ~n541 & ~n542;
  assign n544 = pi129  & ~n543;
  assign n545 = pi64  & ~pi128 ;
  assign n546 = pi63  & pi128 ;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~pi129  & ~n547;
  assign n549 = ~n544 & ~n548;
  assign n550 = n273 & ~n549;
  assign n551 = pi57  & pi128 ;
  assign n552 = pi58  & ~pi128 ;
  assign n553 = ~n551 & ~n552;
  assign n554 = pi129  & ~n553;
  assign n555 = pi60  & ~pi128 ;
  assign n556 = pi59  & pi128 ;
  assign n557 = ~n555 & ~n556;
  assign n558 = ~pi129  & ~n557;
  assign n559 = ~n554 & ~n558;
  assign n560 = n284 & ~n559;
  assign n561 = ~n550 & ~n560;
  assign n562 = pi49  & pi128 ;
  assign n563 = pi50  & ~pi128 ;
  assign n564 = ~n562 & ~n563;
  assign n565 = pi129  & ~n564;
  assign n566 = pi52  & ~pi128 ;
  assign n567 = pi51  & pi128 ;
  assign n568 = ~n566 & ~n567;
  assign n569 = ~pi129  & ~n568;
  assign n570 = ~n565 & ~n569;
  assign n571 = n296 & ~n570;
  assign n572 = pi53  & pi128 ;
  assign n573 = pi54  & ~pi128 ;
  assign n574 = ~n572 & ~n573;
  assign n575 = pi129  & ~n574;
  assign n576 = pi56  & ~pi128 ;
  assign n577 = pi55  & pi128 ;
  assign n578 = ~n576 & ~n577;
  assign n579 = ~pi129  & ~n578;
  assign n580 = ~n575 & ~n579;
  assign n581 = n307 & ~n580;
  assign n582 = ~n571 & ~n581;
  assign n583 = n561 & n582;
  assign n584 = n402 & ~n583;
  assign n585 = pi45  & pi128 ;
  assign n586 = pi46  & ~pi128 ;
  assign n587 = ~n585 & ~n586;
  assign n588 = pi129  & ~n587;
  assign n589 = pi48  & ~pi128 ;
  assign n590 = pi47  & pi128 ;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~pi129  & ~n591;
  assign n593 = ~n588 & ~n592;
  assign n594 = n273 & ~n593;
  assign n595 = pi41  & pi128 ;
  assign n596 = pi42  & ~pi128 ;
  assign n597 = ~n595 & ~n596;
  assign n598 = pi129  & ~n597;
  assign n599 = pi44  & ~pi128 ;
  assign n600 = pi43  & pi128 ;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~pi129  & ~n601;
  assign n603 = ~n598 & ~n602;
  assign n604 = n284 & ~n603;
  assign n605 = ~n594 & ~n604;
  assign n606 = pi33  & pi128 ;
  assign n607 = pi34  & ~pi128 ;
  assign n608 = ~n606 & ~n607;
  assign n609 = pi129  & ~n608;
  assign n610 = pi36  & ~pi128 ;
  assign n611 = pi35  & pi128 ;
  assign n612 = ~n610 & ~n611;
  assign n613 = ~pi129  & ~n612;
  assign n614 = ~n609 & ~n613;
  assign n615 = n296 & ~n614;
  assign n616 = pi40  & ~pi128 ;
  assign n617 = ~pi129  & n616;
  assign n618 = pi37  & pi128 ;
  assign n619 = pi129  & n618;
  assign n620 = ~n617 & ~n619;
  assign n621 = pi39  & pi128 ;
  assign n622 = ~pi129  & n621;
  assign n623 = pi38  & ~pi128 ;
  assign n624 = pi129  & n623;
  assign n625 = ~n622 & ~n624;
  assign n626 = n620 & n625;
  assign n627 = n307 & ~n626;
  assign n628 = ~n615 & ~n627;
  assign n629 = n605 & n628;
  assign n630 = n447 & ~n629;
  assign n631 = ~n584 & ~n630;
  assign n632 = n540 & n631;
  assign n633 = pi134  & ~n632;
  assign po0  = n451 | n633;
  assign n635 = pi81  & ~pi128 ;
  assign n636 = ~pi129  & n635;
  assign n637 = pi78  & pi128 ;
  assign n638 = pi129  & n637;
  assign n639 = ~n636 & ~n638;
  assign n640 = pi80  & pi128 ;
  assign n641 = ~pi129  & n640;
  assign n642 = pi79  & ~pi128 ;
  assign n643 = pi129  & n642;
  assign n644 = ~n641 & ~n643;
  assign n645 = n639 & n644;
  assign n646 = n273 & ~n645;
  assign n647 = pi77  & ~pi128 ;
  assign n648 = ~pi129  & n647;
  assign n649 = pi74  & pi128 ;
  assign n650 = pi129  & n649;
  assign n651 = ~n648 & ~n650;
  assign n652 = pi76  & pi128 ;
  assign n653 = ~pi129  & n652;
  assign n654 = pi75  & ~pi128 ;
  assign n655 = pi129  & n654;
  assign n656 = ~n653 & ~n655;
  assign n657 = n651 & n656;
  assign n658 = n284 & ~n657;
  assign n659 = ~n646 & ~n658;
  assign n660 = pi69  & ~pi128 ;
  assign n661 = ~pi129  & n660;
  assign n662 = pi66  & pi128 ;
  assign n663 = pi129  & n662;
  assign n664 = ~n661 & ~n663;
  assign n665 = pi68  & pi128 ;
  assign n666 = ~pi129  & n665;
  assign n667 = pi67  & ~pi128 ;
  assign n668 = pi129  & n667;
  assign n669 = ~n666 & ~n668;
  assign n670 = n664 & n669;
  assign n671 = n296 & ~n670;
  assign n672 = pi73  & ~pi128 ;
  assign n673 = ~pi129  & n672;
  assign n674 = pi70  & pi128 ;
  assign n675 = pi129  & n674;
  assign n676 = ~n673 & ~n675;
  assign n677 = pi72  & pi128 ;
  assign n678 = ~pi129  & n677;
  assign n679 = pi71  & ~pi128 ;
  assign n680 = pi129  & n679;
  assign n681 = ~n678 & ~n680;
  assign n682 = n676 & n681;
  assign n683 = n307 & ~n682;
  assign n684 = ~n671 & ~n683;
  assign n685 = n659 & n684;
  assign n686 = n311 & ~n685;
  assign n687 = pi97  & ~pi128 ;
  assign n688 = ~pi129  & n687;
  assign n689 = pi94  & pi128 ;
  assign n690 = pi129  & n689;
  assign n691 = ~n688 & ~n690;
  assign n692 = pi96  & pi128 ;
  assign n693 = ~pi129  & n692;
  assign n694 = pi95  & ~pi128 ;
  assign n695 = pi129  & n694;
  assign n696 = ~n693 & ~n695;
  assign n697 = n691 & n696;
  assign n698 = n273 & ~n697;
  assign n699 = pi93  & ~pi128 ;
  assign n700 = ~pi129  & n699;
  assign n701 = pi90  & pi128 ;
  assign n702 = pi129  & n701;
  assign n703 = ~n700 & ~n702;
  assign n704 = pi92  & pi128 ;
  assign n705 = ~pi129  & n704;
  assign n706 = pi91  & ~pi128 ;
  assign n707 = pi129  & n706;
  assign n708 = ~n705 & ~n707;
  assign n709 = n703 & n708;
  assign n710 = n284 & ~n709;
  assign n711 = ~n698 & ~n710;
  assign n712 = pi85  & ~pi128 ;
  assign n713 = ~pi129  & n712;
  assign n714 = pi82  & pi128 ;
  assign n715 = pi129  & n714;
  assign n716 = ~n713 & ~n715;
  assign n717 = pi84  & pi128 ;
  assign n718 = ~pi129  & n717;
  assign n719 = pi83  & ~pi128 ;
  assign n720 = pi129  & n719;
  assign n721 = ~n718 & ~n720;
  assign n722 = n716 & n721;
  assign n723 = n296 & ~n722;
  assign n724 = pi89  & ~pi128 ;
  assign n725 = ~pi129  & n724;
  assign n726 = pi86  & pi128 ;
  assign n727 = pi129  & n726;
  assign n728 = ~n725 & ~n727;
  assign n729 = pi88  & pi128 ;
  assign n730 = ~pi129  & n729;
  assign n731 = pi87  & ~pi128 ;
  assign n732 = pi129  & n731;
  assign n733 = ~n730 & ~n732;
  assign n734 = n728 & n733;
  assign n735 = n307 & ~n734;
  assign n736 = ~n723 & ~n735;
  assign n737 = n711 & n736;
  assign n738 = n356 & ~n737;
  assign n739 = ~n686 & ~n738;
  assign n740 = pi1  & ~pi128 ;
  assign n741 = ~pi129  & n740;
  assign n742 = pi126  & pi128 ;
  assign n743 = pi129  & n742;
  assign n744 = ~n741 & ~n743;
  assign n745 = pi0  & pi128 ;
  assign n746 = ~pi129  & n745;
  assign n747 = pi127  & ~pi128 ;
  assign n748 = pi129  & n747;
  assign n749 = ~n746 & ~n748;
  assign n750 = n744 & n749;
  assign n751 = n273 & ~n750;
  assign n752 = pi125  & ~pi128 ;
  assign n753 = ~pi129  & n752;
  assign n754 = pi122  & pi128 ;
  assign n755 = pi129  & n754;
  assign n756 = ~n753 & ~n755;
  assign n757 = pi124  & pi128 ;
  assign n758 = ~pi129  & n757;
  assign n759 = pi123  & ~pi128 ;
  assign n760 = pi129  & n759;
  assign n761 = ~n758 & ~n760;
  assign n762 = n756 & n761;
  assign n763 = n284 & ~n762;
  assign n764 = ~n751 & ~n763;
  assign n765 = pi117  & ~pi128 ;
  assign n766 = ~pi129  & n765;
  assign n767 = pi114  & pi128 ;
  assign n768 = pi129  & n767;
  assign n769 = ~n766 & ~n768;
  assign n770 = pi116  & pi128 ;
  assign n771 = ~pi129  & n770;
  assign n772 = pi115  & ~pi128 ;
  assign n773 = pi129  & n772;
  assign n774 = ~n771 & ~n773;
  assign n775 = n769 & n774;
  assign n776 = n296 & ~n775;
  assign n777 = pi121  & ~pi128 ;
  assign n778 = ~pi129  & n777;
  assign n779 = pi118  & pi128 ;
  assign n780 = pi129  & n779;
  assign n781 = ~n778 & ~n780;
  assign n782 = pi120  & pi128 ;
  assign n783 = ~pi129  & n782;
  assign n784 = pi119  & ~pi128 ;
  assign n785 = pi129  & n784;
  assign n786 = ~n783 & ~n785;
  assign n787 = n781 & n786;
  assign n788 = n307 & ~n787;
  assign n789 = ~n776 & ~n788;
  assign n790 = n764 & n789;
  assign n791 = n402 & ~n790;
  assign n792 = pi113  & ~pi128 ;
  assign n793 = ~pi129  & n792;
  assign n794 = pi110  & pi128 ;
  assign n795 = pi129  & n794;
  assign n796 = ~n793 & ~n795;
  assign n797 = pi112  & pi128 ;
  assign n798 = ~pi129  & n797;
  assign n799 = pi111  & ~pi128 ;
  assign n800 = pi129  & n799;
  assign n801 = ~n798 & ~n800;
  assign n802 = n796 & n801;
  assign n803 = n273 & ~n802;
  assign n804 = pi109  & ~pi128 ;
  assign n805 = ~pi129  & n804;
  assign n806 = pi106  & pi128 ;
  assign n807 = pi129  & n806;
  assign n808 = ~n805 & ~n807;
  assign n809 = pi108  & pi128 ;
  assign n810 = ~pi129  & n809;
  assign n811 = pi107  & ~pi128 ;
  assign n812 = pi129  & n811;
  assign n813 = ~n810 & ~n812;
  assign n814 = n808 & n813;
  assign n815 = n284 & ~n814;
  assign n816 = ~n803 & ~n815;
  assign n817 = pi101  & ~pi128 ;
  assign n818 = ~pi129  & n817;
  assign n819 = pi98  & pi128 ;
  assign n820 = pi129  & n819;
  assign n821 = ~n818 & ~n820;
  assign n822 = pi100  & pi128 ;
  assign n823 = ~pi129  & n822;
  assign n824 = pi99  & ~pi128 ;
  assign n825 = pi129  & n824;
  assign n826 = ~n823 & ~n825;
  assign n827 = n821 & n826;
  assign n828 = n296 & ~n827;
  assign n829 = pi105  & ~pi128 ;
  assign n830 = ~pi129  & n829;
  assign n831 = pi102  & pi128 ;
  assign n832 = pi129  & n831;
  assign n833 = ~n830 & ~n832;
  assign n834 = pi104  & pi128 ;
  assign n835 = ~pi129  & n834;
  assign n836 = pi103  & ~pi128 ;
  assign n837 = pi129  & n836;
  assign n838 = ~n835 & ~n837;
  assign n839 = n833 & n838;
  assign n840 = n307 & ~n839;
  assign n841 = ~n828 & ~n840;
  assign n842 = n816 & n841;
  assign n843 = n447 & ~n842;
  assign n844 = ~n791 & ~n843;
  assign n845 = n739 & n844;
  assign n846 = ~pi134  & ~n845;
  assign n847 = pi65  & ~pi128 ;
  assign n848 = ~pi129  & n847;
  assign n849 = pi62  & pi128 ;
  assign n850 = pi129  & n849;
  assign n851 = ~n848 & ~n850;
  assign n852 = pi64  & pi128 ;
  assign n853 = ~pi129  & n852;
  assign n854 = pi63  & ~pi128 ;
  assign n855 = pi129  & n854;
  assign n856 = ~n853 & ~n855;
  assign n857 = n851 & n856;
  assign n858 = n273 & ~n857;
  assign n859 = pi61  & ~pi128 ;
  assign n860 = ~pi129  & n859;
  assign n861 = pi58  & pi128 ;
  assign n862 = pi129  & n861;
  assign n863 = ~n860 & ~n862;
  assign n864 = pi60  & pi128 ;
  assign n865 = ~pi129  & n864;
  assign n866 = pi59  & ~pi128 ;
  assign n867 = pi129  & n866;
  assign n868 = ~n865 & ~n867;
  assign n869 = n863 & n868;
  assign n870 = n284 & ~n869;
  assign n871 = ~n858 & ~n870;
  assign n872 = pi53  & ~pi128 ;
  assign n873 = ~pi129  & n872;
  assign n874 = pi50  & pi128 ;
  assign n875 = pi129  & n874;
  assign n876 = ~n873 & ~n875;
  assign n877 = pi52  & pi128 ;
  assign n878 = ~pi129  & n877;
  assign n879 = pi51  & ~pi128 ;
  assign n880 = pi129  & n879;
  assign n881 = ~n878 & ~n880;
  assign n882 = n876 & n881;
  assign n883 = n296 & ~n882;
  assign n884 = pi57  & ~pi128 ;
  assign n885 = ~pi129  & n884;
  assign n886 = pi54  & pi128 ;
  assign n887 = pi129  & n886;
  assign n888 = ~n885 & ~n887;
  assign n889 = pi56  & pi128 ;
  assign n890 = ~pi129  & n889;
  assign n891 = pi55  & ~pi128 ;
  assign n892 = pi129  & n891;
  assign n893 = ~n890 & ~n892;
  assign n894 = n888 & n893;
  assign n895 = n307 & ~n894;
  assign n896 = ~n883 & ~n895;
  assign n897 = n871 & n896;
  assign n898 = n402 & ~n897;
  assign n899 = pi17  & ~pi128 ;
  assign n900 = ~pi129  & n899;
  assign n901 = pi14  & pi128 ;
  assign n902 = pi129  & n901;
  assign n903 = ~n900 & ~n902;
  assign n904 = pi16  & pi128 ;
  assign n905 = ~pi129  & n904;
  assign n906 = pi15  & ~pi128 ;
  assign n907 = pi129  & n906;
  assign n908 = ~n905 & ~n907;
  assign n909 = n903 & n908;
  assign n910 = n273 & ~n909;
  assign n911 = pi13  & ~pi128 ;
  assign n912 = ~pi129  & n911;
  assign n913 = pi10  & pi128 ;
  assign n914 = pi129  & n913;
  assign n915 = ~n912 & ~n914;
  assign n916 = pi12  & pi128 ;
  assign n917 = ~pi129  & n916;
  assign n918 = pi11  & ~pi128 ;
  assign n919 = pi129  & n918;
  assign n920 = ~n917 & ~n919;
  assign n921 = n915 & n920;
  assign n922 = n284 & ~n921;
  assign n923 = ~n910 & ~n922;
  assign n924 = pi5  & ~pi128 ;
  assign n925 = ~pi129  & n924;
  assign n926 = pi2  & pi128 ;
  assign n927 = pi129  & n926;
  assign n928 = ~n925 & ~n927;
  assign n929 = pi4  & pi128 ;
  assign n930 = ~pi129  & n929;
  assign n931 = pi3  & ~pi128 ;
  assign n932 = pi129  & n931;
  assign n933 = ~n930 & ~n932;
  assign n934 = n928 & n933;
  assign n935 = n296 & ~n934;
  assign n936 = pi9  & ~pi128 ;
  assign n937 = ~pi129  & n936;
  assign n938 = pi6  & pi128 ;
  assign n939 = pi129  & n938;
  assign n940 = ~n937 & ~n939;
  assign n941 = pi8  & pi128 ;
  assign n942 = ~pi129  & n941;
  assign n943 = pi7  & ~pi128 ;
  assign n944 = pi129  & n943;
  assign n945 = ~n942 & ~n944;
  assign n946 = n940 & n945;
  assign n947 = n307 & ~n946;
  assign n948 = ~n935 & ~n947;
  assign n949 = n923 & n948;
  assign n950 = n311 & ~n949;
  assign n951 = ~n898 & ~n950;
  assign n952 = pi49  & ~pi128 ;
  assign n953 = ~pi129  & n952;
  assign n954 = pi46  & pi128 ;
  assign n955 = pi129  & n954;
  assign n956 = ~n953 & ~n955;
  assign n957 = pi48  & pi128 ;
  assign n958 = ~pi129  & n957;
  assign n959 = pi47  & ~pi128 ;
  assign n960 = pi129  & n959;
  assign n961 = ~n958 & ~n960;
  assign n962 = n956 & n961;
  assign n963 = n273 & ~n962;
  assign n964 = pi42  & pi128 ;
  assign n965 = pi43  & ~pi128 ;
  assign n966 = ~n964 & ~n965;
  assign n967 = pi129  & ~n966;
  assign n968 = pi45  & ~pi128 ;
  assign n969 = pi44  & pi128 ;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~pi129  & ~n970;
  assign n972 = ~n967 & ~n971;
  assign n973 = n284 & ~n972;
  assign n974 = ~n963 & ~n973;
  assign n975 = pi37  & ~pi128 ;
  assign n976 = ~pi129  & n975;
  assign n977 = pi34  & pi128 ;
  assign n978 = pi129  & n977;
  assign n979 = ~n976 & ~n978;
  assign n980 = pi36  & pi128 ;
  assign n981 = ~pi129  & n980;
  assign n982 = pi35  & ~pi128 ;
  assign n983 = pi129  & n982;
  assign n984 = ~n981 & ~n983;
  assign n985 = n979 & n984;
  assign n986 = n296 & ~n985;
  assign n987 = pi41  & ~pi128 ;
  assign n988 = pi40  & pi128 ;
  assign n989 = ~n987 & ~n988;
  assign n990 = ~pi129  & ~n989;
  assign n991 = pi39  & ~pi128 ;
  assign n992 = pi38  & pi128 ;
  assign n993 = ~n991 & ~n992;
  assign n994 = pi129  & ~n993;
  assign n995 = ~n990 & ~n994;
  assign n996 = n307 & ~n995;
  assign n997 = ~n986 & ~n996;
  assign n998 = n974 & n997;
  assign n999 = n447 & ~n998;
  assign n1000 = pi33  & ~pi128 ;
  assign n1001 = ~pi129  & n1000;
  assign n1002 = pi30  & pi128 ;
  assign n1003 = pi129  & n1002;
  assign n1004 = ~n1001 & ~n1003;
  assign n1005 = pi32  & pi128 ;
  assign n1006 = ~pi129  & n1005;
  assign n1007 = pi31  & ~pi128 ;
  assign n1008 = pi129  & n1007;
  assign n1009 = ~n1006 & ~n1008;
  assign n1010 = n1004 & n1009;
  assign n1011 = n273 & ~n1010;
  assign n1012 = pi29  & ~pi128 ;
  assign n1013 = ~pi129  & n1012;
  assign n1014 = pi26  & pi128 ;
  assign n1015 = pi129  & n1014;
  assign n1016 = ~n1013 & ~n1015;
  assign n1017 = pi28  & pi128 ;
  assign n1018 = ~pi129  & n1017;
  assign n1019 = pi27  & ~pi128 ;
  assign n1020 = pi129  & n1019;
  assign n1021 = ~n1018 & ~n1020;
  assign n1022 = n1016 & n1021;
  assign n1023 = n284 & ~n1022;
  assign n1024 = ~n1011 & ~n1023;
  assign n1025 = pi21  & ~pi128 ;
  assign n1026 = ~pi129  & n1025;
  assign n1027 = pi18  & pi128 ;
  assign n1028 = pi129  & n1027;
  assign n1029 = ~n1026 & ~n1028;
  assign n1030 = pi20  & pi128 ;
  assign n1031 = ~pi129  & n1030;
  assign n1032 = pi19  & ~pi128 ;
  assign n1033 = pi129  & n1032;
  assign n1034 = ~n1031 & ~n1033;
  assign n1035 = n1029 & n1034;
  assign n1036 = n296 & ~n1035;
  assign n1037 = pi25  & ~pi128 ;
  assign n1038 = ~pi129  & n1037;
  assign n1039 = pi22  & pi128 ;
  assign n1040 = pi129  & n1039;
  assign n1041 = ~n1038 & ~n1040;
  assign n1042 = pi24  & pi128 ;
  assign n1043 = ~pi129  & n1042;
  assign n1044 = pi23  & ~pi128 ;
  assign n1045 = pi129  & n1044;
  assign n1046 = ~n1043 & ~n1045;
  assign n1047 = n1041 & n1046;
  assign n1048 = n307 & ~n1047;
  assign n1049 = ~n1036 & ~n1048;
  assign n1050 = n1024 & n1049;
  assign n1051 = n356 & ~n1050;
  assign n1052 = ~n999 & ~n1051;
  assign n1053 = n951 & n1052;
  assign n1054 = pi134  & ~n1053;
  assign po1  = n846 | n1054;
  assign n1056 = ~n336 & ~n337;
  assign n1057 = pi129  & ~n270;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = n273 & ~n1058;
  assign n1060 = ~n266 & ~n267;
  assign n1061 = pi129  & ~n281;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = n284 & ~n1062;
  assign n1064 = ~n1059 & ~n1063;
  assign n1065 = ~n300 & ~n301;
  assign n1066 = pi129  & ~n293;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = n296 & ~n1067;
  assign n1069 = ~n277 & ~n278;
  assign n1070 = pi129  & ~n304;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = n307 & ~n1071;
  assign n1073 = ~n1068 & ~n1072;
  assign n1074 = n1064 & n1073;
  assign n1075 = n311 & ~n1074;
  assign n1076 = ~n427 & ~n428;
  assign n1077 = pi129  & ~n319;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = n273 & ~n1078;
  assign n1080 = ~n315 & ~n316;
  assign n1081 = pi129  & ~n329;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = n284 & ~n1082;
  assign n1084 = ~n1079 & ~n1083;
  assign n1085 = ~n346 & ~n347;
  assign n1086 = pi129  & ~n340;
  assign n1087 = ~n1085 & ~n1086;
  assign n1088 = n296 & ~n1087;
  assign n1089 = ~n325 & ~n326;
  assign n1090 = pi129  & ~n350;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = n307 & ~n1091;
  assign n1093 = ~n1088 & ~n1092;
  assign n1094 = n1084 & n1093;
  assign n1095 = n356 & ~n1094;
  assign n1096 = ~n1075 & ~n1095;
  assign n1097 = ~n475 & ~n476;
  assign n1098 = pi129  & ~n365;
  assign n1099 = ~n1097 & ~n1098;
  assign n1100 = n273 & ~n1099;
  assign n1101 = ~n361 & ~n362;
  assign n1102 = pi129  & ~n375;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = n284 & ~n1103;
  assign n1105 = ~n1100 & ~n1104;
  assign n1106 = ~n392 & ~n393;
  assign n1107 = pi129  & ~n386;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = n296 & ~n1108;
  assign n1110 = ~n371 & ~n372;
  assign n1111 = pi129  & ~n396;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = n307 & ~n1112;
  assign n1114 = ~n1109 & ~n1113;
  assign n1115 = n1105 & n1114;
  assign n1116 = n402 & ~n1115;
  assign n1117 = ~n382 & ~n383;
  assign n1118 = pi129  & ~n410;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = n273 & ~n1119;
  assign n1121 = ~n406 & ~n407;
  assign n1122 = pi129  & ~n420;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = n284 & ~n1123;
  assign n1125 = ~n1120 & ~n1124;
  assign n1126 = ~n437 & ~n438;
  assign n1127 = pi129  & ~n431;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = n296 & ~n1128;
  assign n1130 = ~n416 & ~n417;
  assign n1131 = pi129  & ~n441;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = n307 & ~n1132;
  assign n1134 = ~n1129 & ~n1133;
  assign n1135 = n1125 & n1134;
  assign n1136 = n447 & ~n1135;
  assign n1137 = ~n1116 & ~n1136;
  assign n1138 = n1096 & n1137;
  assign n1139 = ~pi134  & ~n1138;
  assign n1140 = ~n289 & ~n290;
  assign n1141 = pi129  & ~n547;
  assign n1142 = ~n1140 & ~n1141;
  assign n1143 = n273 & ~n1142;
  assign n1144 = ~n543 & ~n544;
  assign n1145 = pi129  & ~n557;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = n284 & ~n1146;
  assign n1148 = ~n1143 & ~n1147;
  assign n1149 = ~n574 & ~n575;
  assign n1150 = pi129  & ~n568;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = n296 & ~n1151;
  assign n1153 = ~n553 & ~n554;
  assign n1154 = pi129  & ~n578;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = n307 & ~n1155;
  assign n1157 = ~n1152 & ~n1156;
  assign n1158 = n1148 & n1157;
  assign n1159 = n402 & ~n1158;
  assign n1160 = ~n519 & ~n520;
  assign n1161 = pi129  & ~n458;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = n273 & ~n1162;
  assign n1164 = ~n454 & ~n455;
  assign n1165 = pi129  & ~n468;
  assign n1166 = ~n1164 & ~n1165;
  assign n1167 = n284 & ~n1166;
  assign n1168 = ~n1163 & ~n1167;
  assign n1169 = ~n485 & ~n486;
  assign n1170 = pi129  & ~n479;
  assign n1171 = ~n1169 & ~n1170;
  assign n1172 = n296 & ~n1171;
  assign n1173 = ~n464 & ~n465;
  assign n1174 = pi129  & ~n489;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = n307 & ~n1175;
  assign n1177 = ~n1172 & ~n1176;
  assign n1178 = n1168 & n1177;
  assign n1179 = n311 & ~n1178;
  assign n1180 = ~n1159 & ~n1179;
  assign n1181 = ~n564 & ~n565;
  assign n1182 = pi129  & ~n591;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = n273 & ~n1183;
  assign n1185 = pi129  & ~n601;
  assign n1186 = ~n587 & ~n588;
  assign n1187 = ~n1185 & ~n1186;
  assign n1188 = n284 & ~n1187;
  assign n1189 = ~n1184 & ~n1188;
  assign n1190 = ~n618 & ~n623;
  assign n1191 = ~pi129  & ~n1190;
  assign n1192 = pi129  & ~n612;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = n296 & ~n1193;
  assign n1195 = ~n597 & ~n598;
  assign n1196 = ~n616 & ~n621;
  assign n1197 = pi129  & ~n1196;
  assign n1198 = ~n1195 & ~n1197;
  assign n1199 = n307 & ~n1198;
  assign n1200 = ~n1194 & ~n1199;
  assign n1201 = n1189 & n1200;
  assign n1202 = n447 & ~n1201;
  assign n1203 = ~n608 & ~n609;
  assign n1204 = pi129  & ~n502;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = n273 & ~n1205;
  assign n1207 = ~n498 & ~n499;
  assign n1208 = pi129  & ~n512;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = n284 & ~n1209;
  assign n1211 = ~n1206 & ~n1210;
  assign n1212 = ~n529 & ~n530;
  assign n1213 = pi129  & ~n523;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = n296 & ~n1214;
  assign n1216 = ~n508 & ~n509;
  assign n1217 = pi129  & ~n533;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = n307 & ~n1218;
  assign n1220 = ~n1215 & ~n1219;
  assign n1221 = n1211 & n1220;
  assign n1222 = n356 & ~n1221;
  assign n1223 = ~n1202 & ~n1222;
  assign n1224 = n1180 & n1223;
  assign n1225 = pi134  & ~n1224;
  assign po2  = n1139 | n1225;
  assign n1227 = pi129  & n792;
  assign n1228 = ~pi129  & n767;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = pi129  & n797;
  assign n1231 = ~pi129  & n772;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = n1229 & n1232;
  assign n1234 = n273 & ~n1233;
  assign n1235 = pi129  & n804;
  assign n1236 = ~pi129  & n794;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = pi129  & n809;
  assign n1239 = ~pi129  & n799;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = n1237 & n1240;
  assign n1242 = n284 & ~n1241;
  assign n1243 = ~n1234 & ~n1242;
  assign n1244 = pi129  & n817;
  assign n1245 = ~pi129  & n831;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = pi129  & n822;
  assign n1248 = ~pi129  & n836;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = n1246 & n1249;
  assign n1251 = n296 & ~n1250;
  assign n1252 = pi129  & n829;
  assign n1253 = ~pi129  & n806;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = pi129  & n834;
  assign n1256 = ~pi129  & n811;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = n1254 & n1257;
  assign n1259 = n307 & ~n1258;
  assign n1260 = ~n1251 & ~n1259;
  assign n1261 = n1243 & n1260;
  assign n1262 = n447 & ~n1261;
  assign n1263 = pi129  & n687;
  assign n1264 = ~pi129  & n819;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = pi129  & n692;
  assign n1267 = ~pi129  & n824;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = n1265 & n1268;
  assign n1270 = n273 & ~n1269;
  assign n1271 = pi129  & n699;
  assign n1272 = ~pi129  & n689;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = pi129  & n704;
  assign n1275 = ~pi129  & n694;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = n1273 & n1276;
  assign n1278 = n284 & ~n1277;
  assign n1279 = ~n1270 & ~n1278;
  assign n1280 = pi129  & n712;
  assign n1281 = ~pi129  & n726;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = pi129  & n717;
  assign n1284 = ~pi129  & n731;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = n1282 & n1285;
  assign n1287 = n296 & ~n1286;
  assign n1288 = pi129  & n724;
  assign n1289 = ~pi129  & n701;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = pi129  & n729;
  assign n1292 = ~pi129  & n706;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = n1290 & n1293;
  assign n1295 = n307 & ~n1294;
  assign n1296 = ~n1287 & ~n1295;
  assign n1297 = n1279 & n1296;
  assign n1298 = n356 & ~n1297;
  assign n1299 = ~n1262 & ~n1298;
  assign n1300 = pi129  & n740;
  assign n1301 = ~pi129  & n926;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = pi129  & n745;
  assign n1304 = ~pi129  & n931;
  assign n1305 = ~n1303 & ~n1304;
  assign n1306 = n1302 & n1305;
  assign n1307 = n273 & ~n1306;
  assign n1308 = pi129  & n752;
  assign n1309 = ~pi129  & n742;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = pi129  & n757;
  assign n1312 = ~pi129  & n747;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = n1310 & n1313;
  assign n1315 = n284 & ~n1314;
  assign n1316 = ~n1307 & ~n1315;
  assign n1317 = pi129  & n765;
  assign n1318 = ~pi129  & n779;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = pi129  & n770;
  assign n1321 = ~pi129  & n784;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = n1319 & n1322;
  assign n1324 = n296 & ~n1323;
  assign n1325 = pi129  & n777;
  assign n1326 = ~pi129  & n754;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = pi129  & n782;
  assign n1329 = ~pi129  & n759;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = n1327 & n1330;
  assign n1332 = n307 & ~n1331;
  assign n1333 = ~n1324 & ~n1332;
  assign n1334 = n1316 & n1333;
  assign n1335 = n402 & ~n1334;
  assign n1336 = pi129  & n635;
  assign n1337 = ~pi129  & n714;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = pi129  & n640;
  assign n1340 = ~pi129  & n719;
  assign n1341 = ~n1339 & ~n1340;
  assign n1342 = n1338 & n1341;
  assign n1343 = n273 & ~n1342;
  assign n1344 = pi129  & n647;
  assign n1345 = ~pi129  & n637;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = pi129  & n652;
  assign n1348 = ~pi129  & n642;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = n1346 & n1349;
  assign n1351 = n284 & ~n1350;
  assign n1352 = ~n1343 & ~n1351;
  assign n1353 = pi129  & n660;
  assign n1354 = ~pi129  & n674;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = pi129  & n665;
  assign n1357 = ~pi129  & n679;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = n1355 & n1358;
  assign n1360 = n296 & ~n1359;
  assign n1361 = pi129  & n672;
  assign n1362 = ~pi129  & n649;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = pi129  & n677;
  assign n1365 = ~pi129  & n654;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = n1363 & n1366;
  assign n1368 = n307 & ~n1367;
  assign n1369 = ~n1360 & ~n1368;
  assign n1370 = n1352 & n1369;
  assign n1371 = n311 & ~n1370;
  assign n1372 = ~n1335 & ~n1371;
  assign n1373 = n1299 & n1372;
  assign n1374 = ~pi134  & ~n1373;
  assign n1375 = pi129  & n847;
  assign n1376 = ~pi129  & n662;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = pi129  & n852;
  assign n1379 = ~pi129  & n667;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = n1377 & n1380;
  assign n1382 = n273 & ~n1381;
  assign n1383 = pi129  & n859;
  assign n1384 = ~pi129  & n849;
  assign n1385 = ~n1383 & ~n1384;
  assign n1386 = pi129  & n864;
  assign n1387 = ~pi129  & n854;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = n1385 & n1388;
  assign n1390 = n284 & ~n1389;
  assign n1391 = ~n1382 & ~n1390;
  assign n1392 = pi129  & n872;
  assign n1393 = ~pi129  & n886;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = pi129  & n877;
  assign n1396 = ~pi129  & n891;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = n1394 & n1397;
  assign n1399 = n296 & ~n1398;
  assign n1400 = pi129  & n884;
  assign n1401 = ~pi129  & n861;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = pi129  & n889;
  assign n1404 = ~pi129  & n866;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = n1402 & n1405;
  assign n1407 = n307 & ~n1406;
  assign n1408 = ~n1399 & ~n1407;
  assign n1409 = n1391 & n1408;
  assign n1410 = n402 & ~n1409;
  assign n1411 = pi129  & n952;
  assign n1412 = ~pi129  & n874;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = pi129  & n957;
  assign n1415 = ~pi129  & n879;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = n1413 & n1416;
  assign n1418 = n273 & ~n1417;
  assign n1419 = pi129  & ~n970;
  assign n1420 = ~n954 & ~n959;
  assign n1421 = ~pi129  & ~n1420;
  assign n1422 = ~n1419 & ~n1421;
  assign n1423 = n284 & ~n1422;
  assign n1424 = ~n1418 & ~n1423;
  assign n1425 = pi129  & n975;
  assign n1426 = ~pi129  & n992;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = pi129  & n980;
  assign n1429 = ~pi129  & n991;
  assign n1430 = ~n1428 & ~n1429;
  assign n1431 = n1427 & n1430;
  assign n1432 = n296 & ~n1431;
  assign n1433 = pi129  & n987;
  assign n1434 = ~pi129  & n964;
  assign n1435 = ~n1433 & ~n1434;
  assign n1436 = pi129  & n988;
  assign n1437 = ~pi129  & n965;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = n1435 & n1438;
  assign n1440 = n307 & ~n1439;
  assign n1441 = ~n1432 & ~n1440;
  assign n1442 = n1424 & n1441;
  assign n1443 = n447 & ~n1442;
  assign n1444 = ~n1410 & ~n1443;
  assign n1445 = pi129  & n899;
  assign n1446 = ~pi129  & n1027;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = pi129  & n904;
  assign n1449 = ~pi129  & n1032;
  assign n1450 = ~n1448 & ~n1449;
  assign n1451 = n1447 & n1450;
  assign n1452 = n273 & ~n1451;
  assign n1453 = pi129  & n911;
  assign n1454 = ~pi129  & n901;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = pi129  & n916;
  assign n1457 = ~pi129  & n906;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = n1455 & n1458;
  assign n1460 = n284 & ~n1459;
  assign n1461 = ~n1452 & ~n1460;
  assign n1462 = pi129  & n924;
  assign n1463 = ~pi129  & n938;
  assign n1464 = ~n1462 & ~n1463;
  assign n1465 = pi129  & n929;
  assign n1466 = ~pi129  & n943;
  assign n1467 = ~n1465 & ~n1466;
  assign n1468 = n1464 & n1467;
  assign n1469 = n296 & ~n1468;
  assign n1470 = pi129  & n936;
  assign n1471 = ~pi129  & n913;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = pi129  & n941;
  assign n1474 = ~pi129  & n918;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = n1472 & n1475;
  assign n1477 = n307 & ~n1476;
  assign n1478 = ~n1469 & ~n1477;
  assign n1479 = n1461 & n1478;
  assign n1480 = n311 & ~n1479;
  assign n1481 = pi129  & n1000;
  assign n1482 = ~pi129  & n977;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = pi129  & n1005;
  assign n1485 = ~pi129  & n982;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = n1483 & n1486;
  assign n1488 = n273 & ~n1487;
  assign n1489 = pi129  & n1012;
  assign n1490 = ~pi129  & n1002;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = pi129  & n1017;
  assign n1493 = ~pi129  & n1007;
  assign n1494 = ~n1492 & ~n1493;
  assign n1495 = n1491 & n1494;
  assign n1496 = n284 & ~n1495;
  assign n1497 = ~n1488 & ~n1496;
  assign n1498 = pi129  & n1025;
  assign n1499 = ~pi129  & n1039;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = pi129  & n1030;
  assign n1502 = ~pi129  & n1044;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = n1500 & n1503;
  assign n1505 = n296 & ~n1504;
  assign n1506 = pi129  & n1037;
  assign n1507 = ~pi129  & n1014;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = pi129  & n1042;
  assign n1510 = ~pi129  & n1019;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = n1508 & n1511;
  assign n1513 = n307 & ~n1512;
  assign n1514 = ~n1505 & ~n1513;
  assign n1515 = n1497 & n1514;
  assign n1516 = n356 & ~n1515;
  assign n1517 = ~n1480 & ~n1516;
  assign n1518 = n1444 & n1517;
  assign n1519 = pi134  & ~n1518;
  assign po3  = n1374 | n1519;
  assign n1521 = n273 & ~n342;
  assign n1522 = ~n272 & n284;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = n296 & ~n306;
  assign n1525 = ~n283 & n307;
  assign n1526 = ~n1524 & ~n1525;
  assign n1527 = n1523 & n1526;
  assign n1528 = n311 & ~n1527;
  assign n1529 = n273 & ~n433;
  assign n1530 = n284 & ~n321;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = n296 & ~n352;
  assign n1533 = n307 & ~n331;
  assign n1534 = ~n1532 & ~n1533;
  assign n1535 = n1531 & n1534;
  assign n1536 = n356 & ~n1535;
  assign n1537 = ~n1528 & ~n1536;
  assign n1538 = n273 & ~n481;
  assign n1539 = n284 & ~n367;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = n296 & ~n398;
  assign n1542 = n307 & ~n377;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = n1540 & n1543;
  assign n1545 = n402 & ~n1544;
  assign n1546 = n273 & ~n388;
  assign n1547 = n284 & ~n412;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = n296 & ~n443;
  assign n1550 = n307 & ~n422;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = n1548 & n1551;
  assign n1553 = n447 & ~n1552;
  assign n1554 = ~n1545 & ~n1553;
  assign n1555 = n1537 & n1554;
  assign n1556 = ~pi134  & ~n1555;
  assign n1557 = n273 & ~n570;
  assign n1558 = n284 & ~n593;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = n296 & ~n626;
  assign n1561 = n307 & ~n603;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = n1559 & n1562;
  assign n1564 = n447 & ~n1563;
  assign n1565 = n273 & ~n295;
  assign n1566 = n284 & ~n549;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = n296 & ~n580;
  assign n1569 = n307 & ~n559;
  assign n1570 = ~n1568 & ~n1569;
  assign n1571 = n1567 & n1570;
  assign n1572 = n402 & ~n1571;
  assign n1573 = ~n1564 & ~n1572;
  assign n1574 = n273 & ~n614;
  assign n1575 = n284 & ~n504;
  assign n1576 = ~n1574 & ~n1575;
  assign n1577 = n296 & ~n535;
  assign n1578 = n307 & ~n514;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = n1576 & n1579;
  assign n1581 = n356 & ~n1580;
  assign n1582 = n273 & ~n525;
  assign n1583 = n284 & ~n460;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = n296 & ~n491;
  assign n1586 = n307 & ~n470;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = n1584 & n1587;
  assign n1589 = n311 & ~n1588;
  assign n1590 = ~n1581 & ~n1589;
  assign n1591 = n1573 & n1590;
  assign n1592 = pi134  & ~n1591;
  assign po4  = n1556 | n1592;
  assign n1594 = n273 & ~n722;
  assign n1595 = n284 & ~n645;
  assign n1596 = ~n1594 & ~n1595;
  assign n1597 = n296 & ~n682;
  assign n1598 = n307 & ~n657;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = n1596 & n1599;
  assign n1601 = n311 & ~n1600;
  assign n1602 = n273 & ~n827;
  assign n1603 = n284 & ~n697;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = n296 & ~n734;
  assign n1606 = n307 & ~n709;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = n1604 & n1607;
  assign n1609 = n356 & ~n1608;
  assign n1610 = ~n1601 & ~n1609;
  assign n1611 = n273 & ~n934;
  assign n1612 = n284 & ~n750;
  assign n1613 = ~n1611 & ~n1612;
  assign n1614 = n296 & ~n787;
  assign n1615 = n307 & ~n762;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = n1613 & n1616;
  assign n1618 = n402 & ~n1617;
  assign n1619 = n273 & ~n775;
  assign n1620 = n284 & ~n802;
  assign n1621 = ~n1619 & ~n1620;
  assign n1622 = n296 & ~n839;
  assign n1623 = n307 & ~n814;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = n1621 & n1624;
  assign n1626 = n447 & ~n1625;
  assign n1627 = ~n1618 & ~n1626;
  assign n1628 = n1610 & n1627;
  assign n1629 = ~pi134  & ~n1628;
  assign n1630 = n273 & ~n882;
  assign n1631 = n284 & ~n962;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = n296 & ~n995;
  assign n1634 = n307 & ~n972;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = n1632 & n1635;
  assign n1637 = n447 & ~n1636;
  assign n1638 = n273 & ~n670;
  assign n1639 = n284 & ~n857;
  assign n1640 = ~n1638 & ~n1639;
  assign n1641 = n296 & ~n894;
  assign n1642 = n307 & ~n869;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = n1640 & n1643;
  assign n1645 = n402 & ~n1644;
  assign n1646 = ~n1637 & ~n1645;
  assign n1647 = n273 & ~n985;
  assign n1648 = n284 & ~n1010;
  assign n1649 = ~n1647 & ~n1648;
  assign n1650 = n296 & ~n1047;
  assign n1651 = n307 & ~n1022;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = n1649 & n1652;
  assign n1654 = n356 & ~n1653;
  assign n1655 = n273 & ~n1035;
  assign n1656 = n284 & ~n909;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = n296 & ~n946;
  assign n1659 = n307 & ~n921;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = n1657 & n1660;
  assign n1662 = n311 & ~n1661;
  assign n1663 = ~n1654 & ~n1662;
  assign n1664 = n1646 & n1663;
  assign n1665 = pi134  & ~n1664;
  assign po5  = n1629 | n1665;
  assign n1667 = n273 & ~n1087;
  assign n1668 = n284 & ~n1058;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = n296 & ~n1071;
  assign n1671 = n307 & ~n1062;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = n1669 & n1672;
  assign n1674 = n311 & ~n1673;
  assign n1675 = n273 & ~n1128;
  assign n1676 = n284 & ~n1078;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = n296 & ~n1091;
  assign n1679 = n307 & ~n1082;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = n1677 & n1680;
  assign n1682 = n356 & ~n1681;
  assign n1683 = ~n1674 & ~n1682;
  assign n1684 = n273 & ~n1171;
  assign n1685 = n284 & ~n1099;
  assign n1686 = ~n1684 & ~n1685;
  assign n1687 = n296 & ~n1112;
  assign n1688 = n307 & ~n1103;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = n1686 & n1689;
  assign n1691 = n402 & ~n1690;
  assign n1692 = n273 & ~n1108;
  assign n1693 = n284 & ~n1119;
  assign n1694 = ~n1692 & ~n1693;
  assign n1695 = n296 & ~n1132;
  assign n1696 = n307 & ~n1123;
  assign n1697 = ~n1695 & ~n1696;
  assign n1698 = n1694 & n1697;
  assign n1699 = n447 & ~n1698;
  assign n1700 = ~n1691 & ~n1699;
  assign n1701 = n1683 & n1700;
  assign n1702 = ~pi134  & ~n1701;
  assign n1703 = n273 & ~n1151;
  assign n1704 = n284 & ~n1183;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = n296 & ~n1198;
  assign n1707 = n307 & ~n1187;
  assign n1708 = ~n1706 & ~n1707;
  assign n1709 = n1705 & n1708;
  assign n1710 = n447 & ~n1709;
  assign n1711 = n273 & ~n1067;
  assign n1712 = n284 & ~n1142;
  assign n1713 = ~n1711 & ~n1712;
  assign n1714 = n296 & ~n1155;
  assign n1715 = n307 & ~n1146;
  assign n1716 = ~n1714 & ~n1715;
  assign n1717 = n1713 & n1716;
  assign n1718 = n402 & ~n1717;
  assign n1719 = ~n1710 & ~n1718;
  assign n1720 = n273 & ~n1193;
  assign n1721 = n284 & ~n1205;
  assign n1722 = ~n1720 & ~n1721;
  assign n1723 = n296 & ~n1218;
  assign n1724 = n307 & ~n1209;
  assign n1725 = ~n1723 & ~n1724;
  assign n1726 = n1722 & n1725;
  assign n1727 = n356 & ~n1726;
  assign n1728 = n273 & ~n1214;
  assign n1729 = n284 & ~n1162;
  assign n1730 = ~n1728 & ~n1729;
  assign n1731 = n296 & ~n1175;
  assign n1732 = n307 & ~n1166;
  assign n1733 = ~n1731 & ~n1732;
  assign n1734 = n1730 & n1733;
  assign n1735 = n311 & ~n1734;
  assign n1736 = ~n1727 & ~n1735;
  assign n1737 = n1719 & n1736;
  assign n1738 = pi134  & ~n1737;
  assign po6  = n1702 | n1738;
  assign n1740 = n273 & ~n1286;
  assign n1741 = n284 & ~n1342;
  assign n1742 = ~n1740 & ~n1741;
  assign n1743 = n296 & ~n1367;
  assign n1744 = n307 & ~n1350;
  assign n1745 = ~n1743 & ~n1744;
  assign n1746 = n1742 & n1745;
  assign n1747 = n311 & ~n1746;
  assign n1748 = n273 & ~n1250;
  assign n1749 = n284 & ~n1269;
  assign n1750 = ~n1748 & ~n1749;
  assign n1751 = n296 & ~n1294;
  assign n1752 = n307 & ~n1277;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = n1750 & n1753;
  assign n1755 = n356 & ~n1754;
  assign n1756 = ~n1747 & ~n1755;
  assign n1757 = n273 & ~n1468;
  assign n1758 = n284 & ~n1306;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = n296 & ~n1331;
  assign n1761 = n307 & ~n1314;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = n1759 & n1762;
  assign n1764 = n402 & ~n1763;
  assign n1765 = n273 & ~n1323;
  assign n1766 = n284 & ~n1233;
  assign n1767 = ~n1765 & ~n1766;
  assign n1768 = n296 & ~n1258;
  assign n1769 = n307 & ~n1241;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = n1767 & n1770;
  assign n1772 = n447 & ~n1771;
  assign n1773 = ~n1764 & ~n1772;
  assign n1774 = n1756 & n1773;
  assign n1775 = ~pi134  & ~n1774;
  assign n1776 = n284 & ~n1417;
  assign n1777 = n307 & ~n1422;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = n296 & ~n1439;
  assign n1780 = n273 & ~n1398;
  assign n1781 = ~n1779 & ~n1780;
  assign n1782 = n1778 & n1781;
  assign n1783 = n447 & ~n1782;
  assign n1784 = n273 & ~n1359;
  assign n1785 = n284 & ~n1381;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = n296 & ~n1406;
  assign n1788 = n307 & ~n1389;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = n1786 & n1789;
  assign n1791 = n402 & ~n1790;
  assign n1792 = ~n1783 & ~n1791;
  assign n1793 = n273 & ~n1431;
  assign n1794 = n284 & ~n1487;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = n296 & ~n1512;
  assign n1797 = n307 & ~n1495;
  assign n1798 = ~n1796 & ~n1797;
  assign n1799 = n1795 & n1798;
  assign n1800 = n356 & ~n1799;
  assign n1801 = n273 & ~n1504;
  assign n1802 = n284 & ~n1451;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = n296 & ~n1476;
  assign n1805 = n307 & ~n1459;
  assign n1806 = ~n1804 & ~n1805;
  assign n1807 = n1803 & n1806;
  assign n1808 = n311 & ~n1807;
  assign n1809 = ~n1800 & ~n1808;
  assign n1810 = n1792 & n1809;
  assign n1811 = pi134  & ~n1810;
  assign po7  = n1775 | n1811;
  assign n1813 = n273 & ~n352;
  assign n1814 = n284 & ~n342;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = ~n283 & n296;
  assign n1817 = ~n272 & n307;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = n1815 & n1818;
  assign n1820 = n311 & ~n1819;
  assign n1821 = n273 & ~n443;
  assign n1822 = n284 & ~n433;
  assign n1823 = ~n1821 & ~n1822;
  assign n1824 = n296 & ~n331;
  assign n1825 = n307 & ~n321;
  assign n1826 = ~n1824 & ~n1825;
  assign n1827 = n1823 & n1826;
  assign n1828 = n356 & ~n1827;
  assign n1829 = ~n1820 & ~n1828;
  assign n1830 = n273 & ~n491;
  assign n1831 = n284 & ~n481;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = n296 & ~n377;
  assign n1834 = n307 & ~n367;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = n1832 & n1835;
  assign n1837 = n402 & ~n1836;
  assign n1838 = n273 & ~n398;
  assign n1839 = n284 & ~n388;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = n296 & ~n422;
  assign n1842 = n307 & ~n412;
  assign n1843 = ~n1841 & ~n1842;
  assign n1844 = n1840 & n1843;
  assign n1845 = n447 & ~n1844;
  assign n1846 = ~n1837 & ~n1845;
  assign n1847 = n1829 & n1846;
  assign n1848 = ~pi134  & ~n1847;
  assign n1849 = n273 & ~n580;
  assign n1850 = n284 & ~n570;
  assign n1851 = ~n1849 & ~n1850;
  assign n1852 = n296 & ~n603;
  assign n1853 = n307 & ~n593;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = n1851 & n1854;
  assign n1856 = n447 & ~n1855;
  assign n1857 = n273 & ~n306;
  assign n1858 = n284 & ~n295;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = n296 & ~n559;
  assign n1861 = n307 & ~n549;
  assign n1862 = ~n1860 & ~n1861;
  assign n1863 = n1859 & n1862;
  assign n1864 = n402 & ~n1863;
  assign n1865 = ~n1856 & ~n1864;
  assign n1866 = n273 & ~n626;
  assign n1867 = n284 & ~n614;
  assign n1868 = ~n1866 & ~n1867;
  assign n1869 = n296 & ~n514;
  assign n1870 = n307 & ~n504;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = n1868 & n1871;
  assign n1873 = n356 & ~n1872;
  assign n1874 = n273 & ~n535;
  assign n1875 = n284 & ~n525;
  assign n1876 = ~n1874 & ~n1875;
  assign n1877 = n296 & ~n470;
  assign n1878 = n307 & ~n460;
  assign n1879 = ~n1877 & ~n1878;
  assign n1880 = n1876 & n1879;
  assign n1881 = n311 & ~n1880;
  assign n1882 = ~n1873 & ~n1881;
  assign n1883 = n1865 & n1882;
  assign n1884 = pi134  & ~n1883;
  assign po8  = n1848 | n1884;
  assign n1886 = n273 & ~n734;
  assign n1887 = n284 & ~n722;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = n296 & ~n657;
  assign n1890 = n307 & ~n645;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = n1888 & n1891;
  assign n1893 = n311 & ~n1892;
  assign n1894 = n273 & ~n839;
  assign n1895 = n284 & ~n827;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = n296 & ~n709;
  assign n1898 = n307 & ~n697;
  assign n1899 = ~n1897 & ~n1898;
  assign n1900 = n1896 & n1899;
  assign n1901 = n356 & ~n1900;
  assign n1902 = ~n1893 & ~n1901;
  assign n1903 = n273 & ~n946;
  assign n1904 = n284 & ~n934;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = n296 & ~n762;
  assign n1907 = n307 & ~n750;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = n1905 & n1908;
  assign n1910 = n402 & ~n1909;
  assign n1911 = n273 & ~n787;
  assign n1912 = n284 & ~n775;
  assign n1913 = ~n1911 & ~n1912;
  assign n1914 = n296 & ~n814;
  assign n1915 = n307 & ~n802;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = n1913 & n1916;
  assign n1918 = n447 & ~n1917;
  assign n1919 = ~n1910 & ~n1918;
  assign n1920 = n1902 & n1919;
  assign n1921 = ~pi134  & ~n1920;
  assign n1922 = n273 & ~n894;
  assign n1923 = n284 & ~n882;
  assign n1924 = ~n1922 & ~n1923;
  assign n1925 = n296 & ~n972;
  assign n1926 = n307 & ~n962;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = n1924 & n1927;
  assign n1929 = n447 & ~n1928;
  assign n1930 = n273 & ~n682;
  assign n1931 = n284 & ~n670;
  assign n1932 = ~n1930 & ~n1931;
  assign n1933 = n296 & ~n869;
  assign n1934 = n307 & ~n857;
  assign n1935 = ~n1933 & ~n1934;
  assign n1936 = n1932 & n1935;
  assign n1937 = n402 & ~n1936;
  assign n1938 = ~n1929 & ~n1937;
  assign n1939 = n273 & ~n995;
  assign n1940 = n284 & ~n985;
  assign n1941 = ~n1939 & ~n1940;
  assign n1942 = n296 & ~n1022;
  assign n1943 = n307 & ~n1010;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = n1941 & n1944;
  assign n1946 = n356 & ~n1945;
  assign n1947 = n273 & ~n1047;
  assign n1948 = n284 & ~n1035;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = n296 & ~n921;
  assign n1951 = n307 & ~n909;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = n1949 & n1952;
  assign n1954 = n311 & ~n1953;
  assign n1955 = ~n1946 & ~n1954;
  assign n1956 = n1938 & n1955;
  assign n1957 = pi134  & ~n1956;
  assign po9  = n1921 | n1957;
  assign n1959 = n273 & ~n1091;
  assign n1960 = n284 & ~n1087;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = n296 & ~n1062;
  assign n1963 = n307 & ~n1058;
  assign n1964 = ~n1962 & ~n1963;
  assign n1965 = n1961 & n1964;
  assign n1966 = n311 & ~n1965;
  assign n1967 = n273 & ~n1132;
  assign n1968 = n284 & ~n1128;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = n296 & ~n1082;
  assign n1971 = n307 & ~n1078;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = n1969 & n1972;
  assign n1974 = n356 & ~n1973;
  assign n1975 = ~n1966 & ~n1974;
  assign n1976 = n273 & ~n1175;
  assign n1977 = n284 & ~n1171;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = n296 & ~n1103;
  assign n1980 = n307 & ~n1099;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = n1978 & n1981;
  assign n1983 = n402 & ~n1982;
  assign n1984 = n273 & ~n1112;
  assign n1985 = n284 & ~n1108;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = n296 & ~n1123;
  assign n1988 = n307 & ~n1119;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = n1986 & n1989;
  assign n1991 = n447 & ~n1990;
  assign n1992 = ~n1983 & ~n1991;
  assign n1993 = n1975 & n1992;
  assign n1994 = ~pi134  & ~n1993;
  assign n1995 = n273 & ~n1155;
  assign n1996 = n284 & ~n1151;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = n296 & ~n1187;
  assign n1999 = n307 & ~n1183;
  assign n2000 = ~n1998 & ~n1999;
  assign n2001 = n1997 & n2000;
  assign n2002 = n447 & ~n2001;
  assign n2003 = n273 & ~n1071;
  assign n2004 = n284 & ~n1067;
  assign n2005 = ~n2003 & ~n2004;
  assign n2006 = n296 & ~n1146;
  assign n2007 = n307 & ~n1142;
  assign n2008 = ~n2006 & ~n2007;
  assign n2009 = n2005 & n2008;
  assign n2010 = n402 & ~n2009;
  assign n2011 = ~n2002 & ~n2010;
  assign n2012 = n273 & ~n1198;
  assign n2013 = n284 & ~n1193;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = n296 & ~n1209;
  assign n2016 = n307 & ~n1205;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = n2014 & n2017;
  assign n2019 = n356 & ~n2018;
  assign n2020 = n273 & ~n1218;
  assign n2021 = n284 & ~n1214;
  assign n2022 = ~n2020 & ~n2021;
  assign n2023 = n296 & ~n1166;
  assign n2024 = n307 & ~n1162;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = n2022 & n2025;
  assign n2027 = n311 & ~n2026;
  assign n2028 = ~n2019 & ~n2027;
  assign n2029 = n2011 & n2028;
  assign n2030 = pi134  & ~n2029;
  assign po10  = n1994 | n2030;
  assign n2032 = n273 & ~n1294;
  assign n2033 = n284 & ~n1286;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = n296 & ~n1350;
  assign n2036 = n307 & ~n1342;
  assign n2037 = ~n2035 & ~n2036;
  assign n2038 = n2034 & n2037;
  assign n2039 = n311 & ~n2038;
  assign n2040 = n273 & ~n1258;
  assign n2041 = n284 & ~n1250;
  assign n2042 = ~n2040 & ~n2041;
  assign n2043 = n296 & ~n1277;
  assign n2044 = n307 & ~n1269;
  assign n2045 = ~n2043 & ~n2044;
  assign n2046 = n2042 & n2045;
  assign n2047 = n356 & ~n2046;
  assign n2048 = ~n2039 & ~n2047;
  assign n2049 = n273 & ~n1476;
  assign n2050 = n284 & ~n1468;
  assign n2051 = ~n2049 & ~n2050;
  assign n2052 = n296 & ~n1314;
  assign n2053 = n307 & ~n1306;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = n2051 & n2054;
  assign n2056 = n402 & ~n2055;
  assign n2057 = n273 & ~n1331;
  assign n2058 = n284 & ~n1323;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = n296 & ~n1241;
  assign n2061 = n307 & ~n1233;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = n2059 & n2062;
  assign n2064 = n447 & ~n2063;
  assign n2065 = ~n2056 & ~n2064;
  assign n2066 = n2048 & n2065;
  assign n2067 = ~pi134  & ~n2066;
  assign n2068 = n273 & ~n1406;
  assign n2069 = n307 & ~n1417;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = n296 & ~n1422;
  assign n2072 = n284 & ~n1398;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = n2070 & n2073;
  assign n2075 = n447 & ~n2074;
  assign n2076 = n273 & ~n1367;
  assign n2077 = n284 & ~n1359;
  assign n2078 = ~n2076 & ~n2077;
  assign n2079 = n296 & ~n1389;
  assign n2080 = n307 & ~n1381;
  assign n2081 = ~n2079 & ~n2080;
  assign n2082 = n2078 & n2081;
  assign n2083 = n402 & ~n2082;
  assign n2084 = ~n2075 & ~n2083;
  assign n2085 = n273 & ~n1439;
  assign n2086 = n284 & ~n1431;
  assign n2087 = ~n2085 & ~n2086;
  assign n2088 = n296 & ~n1495;
  assign n2089 = n307 & ~n1487;
  assign n2090 = ~n2088 & ~n2089;
  assign n2091 = n2087 & n2090;
  assign n2092 = n356 & ~n2091;
  assign n2093 = n273 & ~n1512;
  assign n2094 = n284 & ~n1504;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = n296 & ~n1459;
  assign n2097 = n307 & ~n1451;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = n2095 & n2098;
  assign n2100 = n311 & ~n2099;
  assign n2101 = ~n2092 & ~n2100;
  assign n2102 = n2084 & n2101;
  assign n2103 = pi134  & ~n2102;
  assign po11  = n2067 | n2103;
  assign n2105 = n273 & ~n331;
  assign n2106 = n284 & ~n352;
  assign n2107 = ~n2105 & ~n2106;
  assign n2108 = ~n272 & n296;
  assign n2109 = n307 & ~n342;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = n2107 & n2110;
  assign n2112 = n311 & ~n2111;
  assign n2113 = n273 & ~n422;
  assign n2114 = n284 & ~n443;
  assign n2115 = ~n2113 & ~n2114;
  assign n2116 = n296 & ~n321;
  assign n2117 = n307 & ~n433;
  assign n2118 = ~n2116 & ~n2117;
  assign n2119 = n2115 & n2118;
  assign n2120 = n356 & ~n2119;
  assign n2121 = ~n2112 & ~n2120;
  assign n2122 = n273 & ~n470;
  assign n2123 = n284 & ~n491;
  assign n2124 = ~n2122 & ~n2123;
  assign n2125 = n296 & ~n367;
  assign n2126 = n307 & ~n481;
  assign n2127 = ~n2125 & ~n2126;
  assign n2128 = n2124 & n2127;
  assign n2129 = n402 & ~n2128;
  assign n2130 = n273 & ~n377;
  assign n2131 = n284 & ~n398;
  assign n2132 = ~n2130 & ~n2131;
  assign n2133 = n296 & ~n412;
  assign n2134 = n307 & ~n388;
  assign n2135 = ~n2133 & ~n2134;
  assign n2136 = n2132 & n2135;
  assign n2137 = n447 & ~n2136;
  assign n2138 = ~n2129 & ~n2137;
  assign n2139 = n2121 & n2138;
  assign n2140 = ~pi134  & ~n2139;
  assign n2141 = n273 & ~n559;
  assign n2142 = n284 & ~n580;
  assign n2143 = ~n2141 & ~n2142;
  assign n2144 = n296 & ~n593;
  assign n2145 = n307 & ~n570;
  assign n2146 = ~n2144 & ~n2145;
  assign n2147 = n2143 & n2146;
  assign n2148 = n447 & ~n2147;
  assign n2149 = n273 & ~n283;
  assign n2150 = n284 & ~n306;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = n296 & ~n549;
  assign n2153 = ~n295 & n307;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = n2151 & n2154;
  assign n2156 = n402 & ~n2155;
  assign n2157 = ~n2148 & ~n2156;
  assign n2158 = n273 & ~n603;
  assign n2159 = n284 & ~n626;
  assign n2160 = ~n2158 & ~n2159;
  assign n2161 = n296 & ~n504;
  assign n2162 = n307 & ~n614;
  assign n2163 = ~n2161 & ~n2162;
  assign n2164 = n2160 & n2163;
  assign n2165 = n356 & ~n2164;
  assign n2166 = n273 & ~n514;
  assign n2167 = n284 & ~n535;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = n296 & ~n460;
  assign n2170 = n307 & ~n525;
  assign n2171 = ~n2169 & ~n2170;
  assign n2172 = n2168 & n2171;
  assign n2173 = n311 & ~n2172;
  assign n2174 = ~n2165 & ~n2173;
  assign n2175 = n2157 & n2174;
  assign n2176 = pi134  & ~n2175;
  assign po12  = n2140 | n2176;
  assign n2178 = n273 & ~n709;
  assign n2179 = n284 & ~n734;
  assign n2180 = ~n2178 & ~n2179;
  assign n2181 = n296 & ~n645;
  assign n2182 = n307 & ~n722;
  assign n2183 = ~n2181 & ~n2182;
  assign n2184 = n2180 & n2183;
  assign n2185 = n311 & ~n2184;
  assign n2186 = n273 & ~n814;
  assign n2187 = n284 & ~n839;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = n296 & ~n697;
  assign n2190 = n307 & ~n827;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = n2188 & n2191;
  assign n2193 = n356 & ~n2192;
  assign n2194 = ~n2185 & ~n2193;
  assign n2195 = n273 & ~n921;
  assign n2196 = n284 & ~n946;
  assign n2197 = ~n2195 & ~n2196;
  assign n2198 = n296 & ~n750;
  assign n2199 = n307 & ~n934;
  assign n2200 = ~n2198 & ~n2199;
  assign n2201 = n2197 & n2200;
  assign n2202 = n402 & ~n2201;
  assign n2203 = n273 & ~n762;
  assign n2204 = n284 & ~n787;
  assign n2205 = ~n2203 & ~n2204;
  assign n2206 = n296 & ~n802;
  assign n2207 = n307 & ~n775;
  assign n2208 = ~n2206 & ~n2207;
  assign n2209 = n2205 & n2208;
  assign n2210 = n447 & ~n2209;
  assign n2211 = ~n2202 & ~n2210;
  assign n2212 = n2194 & n2211;
  assign n2213 = ~pi134  & ~n2212;
  assign n2214 = n273 & ~n869;
  assign n2215 = n284 & ~n894;
  assign n2216 = ~n2214 & ~n2215;
  assign n2217 = n296 & ~n962;
  assign n2218 = n307 & ~n882;
  assign n2219 = ~n2217 & ~n2218;
  assign n2220 = n2216 & n2219;
  assign n2221 = n447 & ~n2220;
  assign n2222 = n273 & ~n657;
  assign n2223 = n284 & ~n682;
  assign n2224 = ~n2222 & ~n2223;
  assign n2225 = n296 & ~n857;
  assign n2226 = n307 & ~n670;
  assign n2227 = ~n2225 & ~n2226;
  assign n2228 = n2224 & n2227;
  assign n2229 = n402 & ~n2228;
  assign n2230 = ~n2221 & ~n2229;
  assign n2231 = n273 & ~n972;
  assign n2232 = n284 & ~n995;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = n296 & ~n1010;
  assign n2235 = n307 & ~n985;
  assign n2236 = ~n2234 & ~n2235;
  assign n2237 = n2233 & n2236;
  assign n2238 = n356 & ~n2237;
  assign n2239 = n273 & ~n1022;
  assign n2240 = n284 & ~n1047;
  assign n2241 = ~n2239 & ~n2240;
  assign n2242 = n296 & ~n909;
  assign n2243 = n307 & ~n1035;
  assign n2244 = ~n2242 & ~n2243;
  assign n2245 = n2241 & n2244;
  assign n2246 = n311 & ~n2245;
  assign n2247 = ~n2238 & ~n2246;
  assign n2248 = n2230 & n2247;
  assign n2249 = pi134  & ~n2248;
  assign po13  = n2213 | n2249;
  assign n2251 = n273 & ~n1082;
  assign n2252 = n284 & ~n1091;
  assign n2253 = ~n2251 & ~n2252;
  assign n2254 = n296 & ~n1058;
  assign n2255 = n307 & ~n1087;
  assign n2256 = ~n2254 & ~n2255;
  assign n2257 = n2253 & n2256;
  assign n2258 = n311 & ~n2257;
  assign n2259 = n273 & ~n1123;
  assign n2260 = n284 & ~n1132;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = n296 & ~n1078;
  assign n2263 = n307 & ~n1128;
  assign n2264 = ~n2262 & ~n2263;
  assign n2265 = n2261 & n2264;
  assign n2266 = n356 & ~n2265;
  assign n2267 = ~n2258 & ~n2266;
  assign n2268 = n273 & ~n1166;
  assign n2269 = n284 & ~n1175;
  assign n2270 = ~n2268 & ~n2269;
  assign n2271 = n296 & ~n1099;
  assign n2272 = n307 & ~n1171;
  assign n2273 = ~n2271 & ~n2272;
  assign n2274 = n2270 & n2273;
  assign n2275 = n402 & ~n2274;
  assign n2276 = n273 & ~n1103;
  assign n2277 = n284 & ~n1112;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = n296 & ~n1119;
  assign n2280 = n307 & ~n1108;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = n2278 & n2281;
  assign n2283 = n447 & ~n2282;
  assign n2284 = ~n2275 & ~n2283;
  assign n2285 = n2267 & n2284;
  assign n2286 = ~pi134  & ~n2285;
  assign n2287 = n273 & ~n1146;
  assign n2288 = n284 & ~n1155;
  assign n2289 = ~n2287 & ~n2288;
  assign n2290 = n296 & ~n1183;
  assign n2291 = n307 & ~n1151;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = n2289 & n2292;
  assign n2294 = n447 & ~n2293;
  assign n2295 = n273 & ~n1062;
  assign n2296 = n284 & ~n1071;
  assign n2297 = ~n2295 & ~n2296;
  assign n2298 = n296 & ~n1142;
  assign n2299 = n307 & ~n1067;
  assign n2300 = ~n2298 & ~n2299;
  assign n2301 = n2297 & n2300;
  assign n2302 = n402 & ~n2301;
  assign n2303 = ~n2294 & ~n2302;
  assign n2304 = n273 & ~n1187;
  assign n2305 = n284 & ~n1198;
  assign n2306 = ~n2304 & ~n2305;
  assign n2307 = n296 & ~n1205;
  assign n2308 = n307 & ~n1193;
  assign n2309 = ~n2307 & ~n2308;
  assign n2310 = n2306 & n2309;
  assign n2311 = n356 & ~n2310;
  assign n2312 = n273 & ~n1209;
  assign n2313 = n284 & ~n1218;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = n296 & ~n1162;
  assign n2316 = n307 & ~n1214;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = n2314 & n2317;
  assign n2319 = n311 & ~n2318;
  assign n2320 = ~n2311 & ~n2319;
  assign n2321 = n2303 & n2320;
  assign n2322 = pi134  & ~n2321;
  assign po14  = n2286 | n2322;
  assign n2324 = n273 & ~n1277;
  assign n2325 = n284 & ~n1294;
  assign n2326 = ~n2324 & ~n2325;
  assign n2327 = n296 & ~n1342;
  assign n2328 = n307 & ~n1286;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = n2326 & n2329;
  assign n2331 = n311 & ~n2330;
  assign n2332 = n273 & ~n1241;
  assign n2333 = n284 & ~n1258;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = n296 & ~n1269;
  assign n2336 = n307 & ~n1250;
  assign n2337 = ~n2335 & ~n2336;
  assign n2338 = n2334 & n2337;
  assign n2339 = n356 & ~n2338;
  assign n2340 = ~n2331 & ~n2339;
  assign n2341 = n273 & ~n1459;
  assign n2342 = n284 & ~n1476;
  assign n2343 = ~n2341 & ~n2342;
  assign n2344 = n296 & ~n1306;
  assign n2345 = n307 & ~n1468;
  assign n2346 = ~n2344 & ~n2345;
  assign n2347 = n2343 & n2346;
  assign n2348 = n402 & ~n2347;
  assign n2349 = n273 & ~n1314;
  assign n2350 = n284 & ~n1331;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = n296 & ~n1233;
  assign n2353 = n307 & ~n1323;
  assign n2354 = ~n2352 & ~n2353;
  assign n2355 = n2351 & n2354;
  assign n2356 = n447 & ~n2355;
  assign n2357 = ~n2348 & ~n2356;
  assign n2358 = n2340 & n2357;
  assign n2359 = ~pi134  & ~n2358;
  assign n2360 = n273 & ~n1389;
  assign n2361 = n284 & ~n1406;
  assign n2362 = ~n2360 & ~n2361;
  assign n2363 = n296 & ~n1417;
  assign n2364 = n307 & ~n1398;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = n2362 & n2365;
  assign n2367 = n447 & ~n2366;
  assign n2368 = n273 & ~n1350;
  assign n2369 = n284 & ~n1367;
  assign n2370 = ~n2368 & ~n2369;
  assign n2371 = n296 & ~n1381;
  assign n2372 = n307 & ~n1359;
  assign n2373 = ~n2371 & ~n2372;
  assign n2374 = n2370 & n2373;
  assign n2375 = n402 & ~n2374;
  assign n2376 = ~n2367 & ~n2375;
  assign n2377 = n273 & ~n1422;
  assign n2378 = n284 & ~n1439;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = n296 & ~n1487;
  assign n2381 = n307 & ~n1431;
  assign n2382 = ~n2380 & ~n2381;
  assign n2383 = n2379 & n2382;
  assign n2384 = n356 & ~n2383;
  assign n2385 = n273 & ~n1495;
  assign n2386 = n284 & ~n1512;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = n296 & ~n1451;
  assign n2389 = n307 & ~n1504;
  assign n2390 = ~n2388 & ~n2389;
  assign n2391 = n2387 & n2390;
  assign n2392 = n311 & ~n2391;
  assign n2393 = ~n2384 & ~n2392;
  assign n2394 = n2376 & n2393;
  assign n2395 = pi134  & ~n2394;
  assign po15  = n2359 | n2395;
  assign n2397 = n311 & ~n355;
  assign n2398 = n356 & ~n446;
  assign n2399 = ~n2397 & ~n2398;
  assign n2400 = n402 & ~n494;
  assign n2401 = ~n401 & n447;
  assign n2402 = ~n2400 & ~n2401;
  assign n2403 = n2399 & n2402;
  assign n2404 = ~pi134  & ~n2403;
  assign n2405 = ~n310 & n402;
  assign n2406 = n311 & ~n538;
  assign n2407 = ~n2405 & ~n2406;
  assign n2408 = n447 & ~n583;
  assign n2409 = n356 & ~n629;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = n2407 & n2410;
  assign n2412 = pi134  & ~n2411;
  assign po16  = n2404 | n2412;
  assign n2414 = n311 & ~n737;
  assign n2415 = n356 & ~n842;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = n402 & ~n949;
  assign n2418 = n447 & ~n790;
  assign n2419 = ~n2417 & ~n2418;
  assign n2420 = n2416 & n2419;
  assign n2421 = ~pi134  & ~n2420;
  assign n2422 = n447 & ~n897;
  assign n2423 = n402 & ~n685;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = n356 & ~n998;
  assign n2426 = n311 & ~n1050;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = n2424 & n2427;
  assign n2429 = pi134  & ~n2428;
  assign po17  = n2421 | n2429;
  assign n2431 = n311 & ~n1094;
  assign n2432 = n356 & ~n1135;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = n402 & ~n1178;
  assign n2435 = n447 & ~n1115;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = n2433 & n2436;
  assign n2438 = ~pi134  & ~n2437;
  assign n2439 = n447 & ~n1158;
  assign n2440 = n402 & ~n1074;
  assign n2441 = ~n2439 & ~n2440;
  assign n2442 = n356 & ~n1201;
  assign n2443 = n311 & ~n1221;
  assign n2444 = ~n2442 & ~n2443;
  assign n2445 = n2441 & n2444;
  assign n2446 = pi134  & ~n2445;
  assign po18  = n2438 | n2446;
  assign n2448 = n356 & ~n1261;
  assign n2449 = n311 & ~n1297;
  assign n2450 = ~n2448 & ~n2449;
  assign n2451 = n447 & ~n1334;
  assign n2452 = n402 & ~n1479;
  assign n2453 = ~n2451 & ~n2452;
  assign n2454 = n2450 & n2453;
  assign n2455 = ~pi134  & ~n2454;
  assign n2456 = n447 & ~n1409;
  assign n2457 = n402 & ~n1370;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = n311 & ~n1515;
  assign n2460 = n356 & ~n1442;
  assign n2461 = ~n2459 & ~n2460;
  assign n2462 = n2458 & n2461;
  assign n2463 = pi134  & ~n2462;
  assign po19  = n2455 | n2463;
  assign n2465 = n311 & ~n1535;
  assign n2466 = n356 & ~n1552;
  assign n2467 = ~n2465 & ~n2466;
  assign n2468 = n402 & ~n1588;
  assign n2469 = n447 & ~n1544;
  assign n2470 = ~n2468 & ~n2469;
  assign n2471 = n2467 & n2470;
  assign n2472 = ~pi134  & ~n2471;
  assign n2473 = n402 & ~n1527;
  assign n2474 = n356 & ~n1563;
  assign n2475 = ~n2473 & ~n2474;
  assign n2476 = n311 & ~n1580;
  assign n2477 = n447 & ~n1571;
  assign n2478 = ~n2476 & ~n2477;
  assign n2479 = n2475 & n2478;
  assign n2480 = pi134  & ~n2479;
  assign po20  = n2472 | n2480;
  assign n2482 = n311 & ~n1608;
  assign n2483 = n356 & ~n1625;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = n402 & ~n1661;
  assign n2486 = n447 & ~n1617;
  assign n2487 = ~n2485 & ~n2486;
  assign n2488 = n2484 & n2487;
  assign n2489 = ~pi134  & ~n2488;
  assign n2490 = n402 & ~n1600;
  assign n2491 = n356 & ~n1636;
  assign n2492 = ~n2490 & ~n2491;
  assign n2493 = n311 & ~n1653;
  assign n2494 = n447 & ~n1644;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = n2492 & n2495;
  assign n2497 = pi134  & ~n2496;
  assign po21  = n2489 | n2497;
  assign n2499 = n311 & ~n1681;
  assign n2500 = n356 & ~n1698;
  assign n2501 = ~n2499 & ~n2500;
  assign n2502 = n402 & ~n1734;
  assign n2503 = n447 & ~n1690;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = n2501 & n2504;
  assign n2506 = ~pi134  & ~n2505;
  assign n2507 = n402 & ~n1673;
  assign n2508 = n356 & ~n1709;
  assign n2509 = ~n2507 & ~n2508;
  assign n2510 = n311 & ~n1726;
  assign n2511 = n447 & ~n1717;
  assign n2512 = ~n2510 & ~n2511;
  assign n2513 = n2509 & n2512;
  assign n2514 = pi134  & ~n2513;
  assign po22  = n2506 | n2514;
  assign n2516 = n311 & ~n1754;
  assign n2517 = n402 & ~n1807;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = n447 & ~n1763;
  assign n2520 = n356 & ~n1771;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = n2518 & n2521;
  assign n2523 = ~pi134  & ~n2522;
  assign n2524 = n356 & ~n1782;
  assign n2525 = n447 & ~n1790;
  assign n2526 = ~n2524 & ~n2525;
  assign n2527 = n311 & ~n1799;
  assign n2528 = n402 & ~n1746;
  assign n2529 = ~n2527 & ~n2528;
  assign n2530 = n2526 & n2529;
  assign n2531 = pi134  & ~n2530;
  assign po23  = n2523 | n2531;
  assign n2533 = n311 & ~n1827;
  assign n2534 = n402 & ~n1880;
  assign n2535 = ~n2533 & ~n2534;
  assign n2536 = n447 & ~n1836;
  assign n2537 = n356 & ~n1844;
  assign n2538 = ~n2536 & ~n2537;
  assign n2539 = n2535 & n2538;
  assign n2540 = ~pi134  & ~n2539;
  assign n2541 = n356 & ~n1855;
  assign n2542 = n447 & ~n1863;
  assign n2543 = ~n2541 & ~n2542;
  assign n2544 = n311 & ~n1872;
  assign n2545 = n402 & ~n1819;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = n2543 & n2546;
  assign n2548 = pi134  & ~n2547;
  assign po24  = n2540 | n2548;
  assign n2550 = n311 & ~n1900;
  assign n2551 = n402 & ~n1953;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = n447 & ~n1909;
  assign n2554 = n356 & ~n1917;
  assign n2555 = ~n2553 & ~n2554;
  assign n2556 = n2552 & n2555;
  assign n2557 = ~pi134  & ~n2556;
  assign n2558 = n356 & ~n1928;
  assign n2559 = n447 & ~n1936;
  assign n2560 = ~n2558 & ~n2559;
  assign n2561 = n311 & ~n1945;
  assign n2562 = n402 & ~n1892;
  assign n2563 = ~n2561 & ~n2562;
  assign n2564 = n2560 & n2563;
  assign n2565 = pi134  & ~n2564;
  assign po25  = n2557 | n2565;
  assign n2567 = n311 & ~n1973;
  assign n2568 = n356 & ~n1990;
  assign n2569 = ~n2567 & ~n2568;
  assign n2570 = n402 & ~n2026;
  assign n2571 = n447 & ~n1982;
  assign n2572 = ~n2570 & ~n2571;
  assign n2573 = n2569 & n2572;
  assign n2574 = ~pi134  & ~n2573;
  assign n2575 = n356 & ~n2001;
  assign n2576 = n447 & ~n2009;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = n311 & ~n2018;
  assign n2579 = n402 & ~n1965;
  assign n2580 = ~n2578 & ~n2579;
  assign n2581 = n2577 & n2580;
  assign n2582 = pi134  & ~n2581;
  assign po26  = n2574 | n2582;
  assign n2584 = n311 & ~n2046;
  assign n2585 = n356 & ~n2063;
  assign n2586 = ~n2584 & ~n2585;
  assign n2587 = n402 & ~n2099;
  assign n2588 = n447 & ~n2055;
  assign n2589 = ~n2587 & ~n2588;
  assign n2590 = n2586 & n2589;
  assign n2591 = ~pi134  & ~n2590;
  assign n2592 = n356 & ~n2074;
  assign n2593 = n447 & ~n2082;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = n311 & ~n2091;
  assign n2596 = n402 & ~n2038;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = n2594 & n2597;
  assign n2599 = pi134  & ~n2598;
  assign po27  = n2591 | n2599;
  assign n2601 = n311 & ~n2119;
  assign n2602 = n356 & ~n2136;
  assign n2603 = ~n2601 & ~n2602;
  assign n2604 = n402 & ~n2172;
  assign n2605 = n447 & ~n2128;
  assign n2606 = ~n2604 & ~n2605;
  assign n2607 = n2603 & n2606;
  assign n2608 = ~pi134  & ~n2607;
  assign n2609 = n356 & ~n2147;
  assign n2610 = n447 & ~n2155;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = n311 & ~n2164;
  assign n2613 = n402 & ~n2111;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = n2611 & n2614;
  assign n2616 = pi134  & ~n2615;
  assign po28  = n2608 | n2616;
  assign n2618 = n311 & ~n2192;
  assign n2619 = n356 & ~n2209;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = n402 & ~n2245;
  assign n2622 = n447 & ~n2201;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = n2620 & n2623;
  assign n2625 = ~pi134  & ~n2624;
  assign n2626 = n356 & ~n2220;
  assign n2627 = n447 & ~n2228;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = n311 & ~n2237;
  assign n2630 = n402 & ~n2184;
  assign n2631 = ~n2629 & ~n2630;
  assign n2632 = n2628 & n2631;
  assign n2633 = pi134  & ~n2632;
  assign po29  = n2625 | n2633;
  assign n2635 = n311 & ~n2265;
  assign n2636 = n356 & ~n2282;
  assign n2637 = ~n2635 & ~n2636;
  assign n2638 = n402 & ~n2318;
  assign n2639 = n447 & ~n2274;
  assign n2640 = ~n2638 & ~n2639;
  assign n2641 = n2637 & n2640;
  assign n2642 = ~pi134  & ~n2641;
  assign n2643 = n356 & ~n2293;
  assign n2644 = n447 & ~n2301;
  assign n2645 = ~n2643 & ~n2644;
  assign n2646 = n311 & ~n2310;
  assign n2647 = n402 & ~n2257;
  assign n2648 = ~n2646 & ~n2647;
  assign n2649 = n2645 & n2648;
  assign n2650 = pi134  & ~n2649;
  assign po30  = n2642 | n2650;
  assign n2652 = n311 & ~n2338;
  assign n2653 = n356 & ~n2355;
  assign n2654 = ~n2652 & ~n2653;
  assign n2655 = n402 & ~n2391;
  assign n2656 = n447 & ~n2347;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = n2654 & n2657;
  assign n2659 = ~pi134  & ~n2658;
  assign n2660 = n356 & ~n2366;
  assign n2661 = n447 & ~n2374;
  assign n2662 = ~n2660 & ~n2661;
  assign n2663 = n311 & ~n2383;
  assign n2664 = n402 & ~n2330;
  assign n2665 = ~n2663 & ~n2664;
  assign n2666 = n2662 & n2665;
  assign n2667 = pi134  & ~n2666;
  assign po31  = n2659 | n2667;
  assign n2669 = n311 & ~n446;
  assign n2670 = n356 & ~n401;
  assign n2671 = ~n2669 & ~n2670;
  assign n2672 = n402 & ~n538;
  assign n2673 = n447 & ~n494;
  assign n2674 = ~n2672 & ~n2673;
  assign n2675 = n2671 & n2674;
  assign n2676 = ~pi134  & ~n2675;
  assign n2677 = ~n310 & n447;
  assign n2678 = ~n355 & n402;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = n356 & ~n583;
  assign n2681 = n311 & ~n629;
  assign n2682 = ~n2680 & ~n2681;
  assign n2683 = n2679 & n2682;
  assign n2684 = pi134  & ~n2683;
  assign po32  = n2676 | n2684;
  assign n2686 = n311 & ~n842;
  assign n2687 = n356 & ~n790;
  assign n2688 = ~n2686 & ~n2687;
  assign n2689 = n402 & ~n1050;
  assign n2690 = n447 & ~n949;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = n2688 & n2691;
  assign n2693 = ~pi134  & ~n2692;
  assign n2694 = n356 & ~n897;
  assign n2695 = n447 & ~n685;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = n311 & ~n998;
  assign n2698 = n402 & ~n737;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = n2696 & n2699;
  assign n2701 = pi134  & ~n2700;
  assign po33  = n2693 | n2701;
  assign n2703 = n311 & ~n1135;
  assign n2704 = n356 & ~n1115;
  assign n2705 = ~n2703 & ~n2704;
  assign n2706 = n402 & ~n1221;
  assign n2707 = n447 & ~n1178;
  assign n2708 = ~n2706 & ~n2707;
  assign n2709 = n2705 & n2708;
  assign n2710 = ~pi134  & ~n2709;
  assign n2711 = n356 & ~n1158;
  assign n2712 = n447 & ~n1074;
  assign n2713 = ~n2711 & ~n2712;
  assign n2714 = n311 & ~n1201;
  assign n2715 = n402 & ~n1094;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = n2713 & n2716;
  assign n2718 = pi134  & ~n2717;
  assign po34  = n2710 | n2718;
  assign n2720 = n311 & ~n1261;
  assign n2721 = n402 & ~n1515;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = n356 & ~n1334;
  assign n2724 = n447 & ~n1479;
  assign n2725 = ~n2723 & ~n2724;
  assign n2726 = n2722 & n2725;
  assign n2727 = ~pi134  & ~n2726;
  assign n2728 = n356 & ~n1409;
  assign n2729 = n402 & ~n1297;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = n311 & ~n1442;
  assign n2732 = n447 & ~n1370;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = n2730 & n2733;
  assign n2735 = pi134  & ~n2734;
  assign po35  = n2727 | n2735;
  assign n2737 = n311 & ~n1552;
  assign n2738 = n356 & ~n1544;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = n402 & ~n1580;
  assign n2741 = n447 & ~n1588;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = n2739 & n2742;
  assign n2744 = ~pi134  & ~n2743;
  assign n2745 = n447 & ~n1527;
  assign n2746 = n402 & ~n1535;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = n356 & ~n1571;
  assign n2749 = n311 & ~n1563;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = n2747 & n2750;
  assign n2752 = pi134  & ~n2751;
  assign po36  = n2744 | n2752;
  assign n2754 = n311 & ~n1625;
  assign n2755 = n356 & ~n1617;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = n402 & ~n1653;
  assign n2758 = n447 & ~n1661;
  assign n2759 = ~n2757 & ~n2758;
  assign n2760 = n2756 & n2759;
  assign n2761 = ~pi134  & ~n2760;
  assign n2762 = n447 & ~n1600;
  assign n2763 = n402 & ~n1608;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = n356 & ~n1644;
  assign n2766 = n311 & ~n1636;
  assign n2767 = ~n2765 & ~n2766;
  assign n2768 = n2764 & n2767;
  assign n2769 = pi134  & ~n2768;
  assign po37  = n2761 | n2769;
  assign n2771 = n311 & ~n1698;
  assign n2772 = n356 & ~n1690;
  assign n2773 = ~n2771 & ~n2772;
  assign n2774 = n402 & ~n1726;
  assign n2775 = n447 & ~n1734;
  assign n2776 = ~n2774 & ~n2775;
  assign n2777 = n2773 & n2776;
  assign n2778 = ~pi134  & ~n2777;
  assign n2779 = n447 & ~n1673;
  assign n2780 = n402 & ~n1681;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = n356 & ~n1717;
  assign n2783 = n311 & ~n1709;
  assign n2784 = ~n2782 & ~n2783;
  assign n2785 = n2781 & n2784;
  assign n2786 = pi134  & ~n2785;
  assign po38  = n2778 | n2786;
  assign n2788 = n447 & ~n1807;
  assign n2789 = n402 & ~n1799;
  assign n2790 = ~n2788 & ~n2789;
  assign n2791 = n356 & ~n1763;
  assign n2792 = n311 & ~n1771;
  assign n2793 = ~n2791 & ~n2792;
  assign n2794 = n2790 & n2793;
  assign n2795 = ~pi134  & ~n2794;
  assign n2796 = n311 & ~n1782;
  assign n2797 = n356 & ~n1790;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = n402 & ~n1754;
  assign n2800 = n447 & ~n1746;
  assign n2801 = ~n2799 & ~n2800;
  assign n2802 = n2798 & n2801;
  assign n2803 = pi134  & ~n2802;
  assign po39  = n2795 | n2803;
  assign n2805 = n447 & ~n1880;
  assign n2806 = n402 & ~n1872;
  assign n2807 = ~n2805 & ~n2806;
  assign n2808 = n356 & ~n1836;
  assign n2809 = n311 & ~n1844;
  assign n2810 = ~n2808 & ~n2809;
  assign n2811 = n2807 & n2810;
  assign n2812 = ~pi134  & ~n2811;
  assign n2813 = n311 & ~n1855;
  assign n2814 = n356 & ~n1863;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = n402 & ~n1827;
  assign n2817 = n447 & ~n1819;
  assign n2818 = ~n2816 & ~n2817;
  assign n2819 = n2815 & n2818;
  assign n2820 = pi134  & ~n2819;
  assign po40  = n2812 | n2820;
  assign n2822 = n447 & ~n1953;
  assign n2823 = n402 & ~n1945;
  assign n2824 = ~n2822 & ~n2823;
  assign n2825 = n356 & ~n1909;
  assign n2826 = n311 & ~n1917;
  assign n2827 = ~n2825 & ~n2826;
  assign n2828 = n2824 & n2827;
  assign n2829 = ~pi134  & ~n2828;
  assign n2830 = n311 & ~n1928;
  assign n2831 = n356 & ~n1936;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = n402 & ~n1900;
  assign n2834 = n447 & ~n1892;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = n2832 & n2835;
  assign n2837 = pi134  & ~n2836;
  assign po41  = n2829 | n2837;
  assign n2839 = n311 & ~n1990;
  assign n2840 = n356 & ~n1982;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = n402 & ~n2018;
  assign n2843 = n447 & ~n2026;
  assign n2844 = ~n2842 & ~n2843;
  assign n2845 = n2841 & n2844;
  assign n2846 = ~pi134  & ~n2845;
  assign n2847 = n311 & ~n2001;
  assign n2848 = n356 & ~n2009;
  assign n2849 = ~n2847 & ~n2848;
  assign n2850 = n402 & ~n1973;
  assign n2851 = n447 & ~n1965;
  assign n2852 = ~n2850 & ~n2851;
  assign n2853 = n2849 & n2852;
  assign n2854 = pi134  & ~n2853;
  assign po42  = n2846 | n2854;
  assign n2856 = n311 & ~n2063;
  assign n2857 = n356 & ~n2055;
  assign n2858 = ~n2856 & ~n2857;
  assign n2859 = n402 & ~n2091;
  assign n2860 = n447 & ~n2099;
  assign n2861 = ~n2859 & ~n2860;
  assign n2862 = n2858 & n2861;
  assign n2863 = ~pi134  & ~n2862;
  assign n2864 = n311 & ~n2074;
  assign n2865 = n356 & ~n2082;
  assign n2866 = ~n2864 & ~n2865;
  assign n2867 = n402 & ~n2046;
  assign n2868 = n447 & ~n2038;
  assign n2869 = ~n2867 & ~n2868;
  assign n2870 = n2866 & n2869;
  assign n2871 = pi134  & ~n2870;
  assign po43  = n2863 | n2871;
  assign n2873 = n311 & ~n2136;
  assign n2874 = n356 & ~n2128;
  assign n2875 = ~n2873 & ~n2874;
  assign n2876 = n402 & ~n2164;
  assign n2877 = n447 & ~n2172;
  assign n2878 = ~n2876 & ~n2877;
  assign n2879 = n2875 & n2878;
  assign n2880 = ~pi134  & ~n2879;
  assign n2881 = n311 & ~n2147;
  assign n2882 = n356 & ~n2155;
  assign n2883 = ~n2881 & ~n2882;
  assign n2884 = n402 & ~n2119;
  assign n2885 = n447 & ~n2111;
  assign n2886 = ~n2884 & ~n2885;
  assign n2887 = n2883 & n2886;
  assign n2888 = pi134  & ~n2887;
  assign po44  = n2880 | n2888;
  assign n2890 = n311 & ~n2209;
  assign n2891 = n356 & ~n2201;
  assign n2892 = ~n2890 & ~n2891;
  assign n2893 = n402 & ~n2237;
  assign n2894 = n447 & ~n2245;
  assign n2895 = ~n2893 & ~n2894;
  assign n2896 = n2892 & n2895;
  assign n2897 = ~pi134  & ~n2896;
  assign n2898 = n311 & ~n2220;
  assign n2899 = n356 & ~n2228;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = n402 & ~n2192;
  assign n2902 = n447 & ~n2184;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = n2900 & n2903;
  assign n2905 = pi134  & ~n2904;
  assign po45  = n2897 | n2905;
  assign n2907 = n311 & ~n2282;
  assign n2908 = n356 & ~n2274;
  assign n2909 = ~n2907 & ~n2908;
  assign n2910 = n402 & ~n2310;
  assign n2911 = n447 & ~n2318;
  assign n2912 = ~n2910 & ~n2911;
  assign n2913 = n2909 & n2912;
  assign n2914 = ~pi134  & ~n2913;
  assign n2915 = n311 & ~n2293;
  assign n2916 = n356 & ~n2301;
  assign n2917 = ~n2915 & ~n2916;
  assign n2918 = n402 & ~n2265;
  assign n2919 = n447 & ~n2257;
  assign n2920 = ~n2918 & ~n2919;
  assign n2921 = n2917 & n2920;
  assign n2922 = pi134  & ~n2921;
  assign po46  = n2914 | n2922;
  assign n2924 = n311 & ~n2355;
  assign n2925 = n356 & ~n2347;
  assign n2926 = ~n2924 & ~n2925;
  assign n2927 = n402 & ~n2383;
  assign n2928 = n447 & ~n2391;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = n2926 & n2929;
  assign n2931 = ~pi134  & ~n2930;
  assign n2932 = n311 & ~n2366;
  assign n2933 = n356 & ~n2374;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = n402 & ~n2338;
  assign n2936 = n447 & ~n2330;
  assign n2937 = ~n2935 & ~n2936;
  assign n2938 = n2934 & n2937;
  assign n2939 = pi134  & ~n2938;
  assign po47  = n2931 | n2939;
  assign n2941 = n311 & ~n401;
  assign n2942 = n356 & ~n494;
  assign n2943 = ~n2941 & ~n2942;
  assign n2944 = n402 & ~n629;
  assign n2945 = n447 & ~n538;
  assign n2946 = ~n2944 & ~n2945;
  assign n2947 = n2943 & n2946;
  assign n2948 = ~pi134  & ~n2947;
  assign n2949 = ~n310 & n356;
  assign n2950 = ~n355 & n447;
  assign n2951 = ~n2949 & ~n2950;
  assign n2952 = n311 & ~n583;
  assign n2953 = n402 & ~n446;
  assign n2954 = ~n2952 & ~n2953;
  assign n2955 = n2951 & n2954;
  assign n2956 = pi134  & ~n2955;
  assign po48  = n2948 | n2956;
  assign n2958 = n311 & ~n790;
  assign n2959 = n356 & ~n949;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = n402 & ~n998;
  assign n2962 = n447 & ~n1050;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = n2960 & n2963;
  assign n2965 = ~pi134  & ~n2964;
  assign n2966 = n311 & ~n897;
  assign n2967 = n356 & ~n685;
  assign n2968 = ~n2966 & ~n2967;
  assign n2969 = n402 & ~n842;
  assign n2970 = n447 & ~n737;
  assign n2971 = ~n2969 & ~n2970;
  assign n2972 = n2968 & n2971;
  assign n2973 = pi134  & ~n2972;
  assign po49  = n2965 | n2973;
  assign n2975 = n311 & ~n1115;
  assign n2976 = n356 & ~n1178;
  assign n2977 = ~n2975 & ~n2976;
  assign n2978 = n402 & ~n1201;
  assign n2979 = n447 & ~n1221;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = n2977 & n2980;
  assign n2982 = ~pi134  & ~n2981;
  assign n2983 = n311 & ~n1158;
  assign n2984 = n356 & ~n1074;
  assign n2985 = ~n2983 & ~n2984;
  assign n2986 = n402 & ~n1135;
  assign n2987 = n447 & ~n1094;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = n2985 & n2988;
  assign n2990 = pi134  & ~n2989;
  assign po50  = n2982 | n2990;
  assign n2992 = n402 & ~n1442;
  assign n2993 = n447 & ~n1515;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = n311 & ~n1334;
  assign n2996 = n356 & ~n1479;
  assign n2997 = ~n2995 & ~n2996;
  assign n2998 = n2994 & n2997;
  assign n2999 = ~pi134  & ~n2998;
  assign n3000 = n311 & ~n1409;
  assign n3001 = n402 & ~n1261;
  assign n3002 = ~n3000 & ~n3001;
  assign n3003 = n356 & ~n1370;
  assign n3004 = n447 & ~n1297;
  assign n3005 = ~n3003 & ~n3004;
  assign n3006 = n3002 & n3005;
  assign n3007 = pi134  & ~n3006;
  assign po51  = n2999 | n3007;
  assign n3009 = n402 & ~n1563;
  assign n3010 = n311 & ~n1544;
  assign n3011 = ~n3009 & ~n3010;
  assign n3012 = n447 & ~n1580;
  assign n3013 = n356 & ~n1588;
  assign n3014 = ~n3012 & ~n3013;
  assign n3015 = n3011 & n3014;
  assign n3016 = ~pi134  & ~n3015;
  assign n3017 = n356 & ~n1527;
  assign n3018 = n447 & ~n1535;
  assign n3019 = ~n3017 & ~n3018;
  assign n3020 = n402 & ~n1552;
  assign n3021 = n311 & ~n1571;
  assign n3022 = ~n3020 & ~n3021;
  assign n3023 = n3019 & n3022;
  assign n3024 = pi134  & ~n3023;
  assign po52  = n3016 | n3024;
  assign n3026 = n402 & ~n1636;
  assign n3027 = n311 & ~n1617;
  assign n3028 = ~n3026 & ~n3027;
  assign n3029 = n447 & ~n1653;
  assign n3030 = n356 & ~n1661;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = n3028 & n3031;
  assign n3033 = ~pi134  & ~n3032;
  assign n3034 = n356 & ~n1600;
  assign n3035 = n447 & ~n1608;
  assign n3036 = ~n3034 & ~n3035;
  assign n3037 = n402 & ~n1625;
  assign n3038 = n311 & ~n1644;
  assign n3039 = ~n3037 & ~n3038;
  assign n3040 = n3036 & n3039;
  assign n3041 = pi134  & ~n3040;
  assign po53  = n3033 | n3041;
  assign n3043 = n402 & ~n1709;
  assign n3044 = n311 & ~n1690;
  assign n3045 = ~n3043 & ~n3044;
  assign n3046 = n447 & ~n1726;
  assign n3047 = n356 & ~n1734;
  assign n3048 = ~n3046 & ~n3047;
  assign n3049 = n3045 & n3048;
  assign n3050 = ~pi134  & ~n3049;
  assign n3051 = n356 & ~n1673;
  assign n3052 = n447 & ~n1681;
  assign n3053 = ~n3051 & ~n3052;
  assign n3054 = n402 & ~n1698;
  assign n3055 = n311 & ~n1717;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = n3053 & n3056;
  assign n3058 = pi134  & ~n3057;
  assign po54  = n3050 | n3058;
  assign n3060 = n402 & ~n1782;
  assign n3061 = n356 & ~n1807;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = n311 & ~n1763;
  assign n3064 = n447 & ~n1799;
  assign n3065 = ~n3063 & ~n3064;
  assign n3066 = n3062 & n3065;
  assign n3067 = ~pi134  & ~n3066;
  assign n3068 = n311 & ~n1790;
  assign n3069 = n356 & ~n1746;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = n402 & ~n1771;
  assign n3072 = n447 & ~n1754;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = n3070 & n3073;
  assign n3075 = pi134  & ~n3074;
  assign po55  = n3067 | n3075;
  assign n3077 = n402 & ~n1855;
  assign n3078 = n356 & ~n1880;
  assign n3079 = ~n3077 & ~n3078;
  assign n3080 = n311 & ~n1836;
  assign n3081 = n447 & ~n1872;
  assign n3082 = ~n3080 & ~n3081;
  assign n3083 = n3079 & n3082;
  assign n3084 = ~pi134  & ~n3083;
  assign n3085 = n311 & ~n1863;
  assign n3086 = n356 & ~n1819;
  assign n3087 = ~n3085 & ~n3086;
  assign n3088 = n402 & ~n1844;
  assign n3089 = n447 & ~n1827;
  assign n3090 = ~n3088 & ~n3089;
  assign n3091 = n3087 & n3090;
  assign n3092 = pi134  & ~n3091;
  assign po56  = n3084 | n3092;
  assign n3094 = n402 & ~n1928;
  assign n3095 = n356 & ~n1953;
  assign n3096 = ~n3094 & ~n3095;
  assign n3097 = n311 & ~n1909;
  assign n3098 = n447 & ~n1945;
  assign n3099 = ~n3097 & ~n3098;
  assign n3100 = n3096 & n3099;
  assign n3101 = ~pi134  & ~n3100;
  assign n3102 = n311 & ~n1936;
  assign n3103 = n356 & ~n1892;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = n402 & ~n1917;
  assign n3106 = n447 & ~n1900;
  assign n3107 = ~n3105 & ~n3106;
  assign n3108 = n3104 & n3107;
  assign n3109 = pi134  & ~n3108;
  assign po57  = n3101 | n3109;
  assign n3111 = n402 & ~n2001;
  assign n3112 = n311 & ~n1982;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = n447 & ~n2018;
  assign n3115 = n356 & ~n2026;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = n3113 & n3116;
  assign n3118 = ~pi134  & ~n3117;
  assign n3119 = n311 & ~n2009;
  assign n3120 = n356 & ~n1965;
  assign n3121 = ~n3119 & ~n3120;
  assign n3122 = n402 & ~n1990;
  assign n3123 = n447 & ~n1973;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = n3121 & n3124;
  assign n3126 = pi134  & ~n3125;
  assign po58  = n3118 | n3126;
  assign n3128 = n402 & ~n2074;
  assign n3129 = n311 & ~n2055;
  assign n3130 = ~n3128 & ~n3129;
  assign n3131 = n447 & ~n2091;
  assign n3132 = n356 & ~n2099;
  assign n3133 = ~n3131 & ~n3132;
  assign n3134 = n3130 & n3133;
  assign n3135 = ~pi134  & ~n3134;
  assign n3136 = n311 & ~n2082;
  assign n3137 = n356 & ~n2038;
  assign n3138 = ~n3136 & ~n3137;
  assign n3139 = n402 & ~n2063;
  assign n3140 = n447 & ~n2046;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = n3138 & n3141;
  assign n3143 = pi134  & ~n3142;
  assign po59  = n3135 | n3143;
  assign n3145 = n402 & ~n2147;
  assign n3146 = n311 & ~n2128;
  assign n3147 = ~n3145 & ~n3146;
  assign n3148 = n447 & ~n2164;
  assign n3149 = n356 & ~n2172;
  assign n3150 = ~n3148 & ~n3149;
  assign n3151 = n3147 & n3150;
  assign n3152 = ~pi134  & ~n3151;
  assign n3153 = n311 & ~n2155;
  assign n3154 = n356 & ~n2111;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = n402 & ~n2136;
  assign n3157 = n447 & ~n2119;
  assign n3158 = ~n3156 & ~n3157;
  assign n3159 = n3155 & n3158;
  assign n3160 = pi134  & ~n3159;
  assign po60  = n3152 | n3160;
  assign n3162 = n402 & ~n2220;
  assign n3163 = n311 & ~n2201;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = n447 & ~n2237;
  assign n3166 = n356 & ~n2245;
  assign n3167 = ~n3165 & ~n3166;
  assign n3168 = n3164 & n3167;
  assign n3169 = ~pi134  & ~n3168;
  assign n3170 = n311 & ~n2228;
  assign n3171 = n356 & ~n2184;
  assign n3172 = ~n3170 & ~n3171;
  assign n3173 = n402 & ~n2209;
  assign n3174 = n447 & ~n2192;
  assign n3175 = ~n3173 & ~n3174;
  assign n3176 = n3172 & n3175;
  assign n3177 = pi134  & ~n3176;
  assign po61  = n3169 | n3177;
  assign n3179 = n402 & ~n2293;
  assign n3180 = n311 & ~n2274;
  assign n3181 = ~n3179 & ~n3180;
  assign n3182 = n447 & ~n2310;
  assign n3183 = n356 & ~n2318;
  assign n3184 = ~n3182 & ~n3183;
  assign n3185 = n3181 & n3184;
  assign n3186 = ~pi134  & ~n3185;
  assign n3187 = n311 & ~n2301;
  assign n3188 = n356 & ~n2257;
  assign n3189 = ~n3187 & ~n3188;
  assign n3190 = n402 & ~n2282;
  assign n3191 = n447 & ~n2265;
  assign n3192 = ~n3190 & ~n3191;
  assign n3193 = n3189 & n3192;
  assign n3194 = pi134  & ~n3193;
  assign po62  = n3186 | n3194;
  assign n3196 = n402 & ~n2366;
  assign n3197 = n311 & ~n2347;
  assign n3198 = ~n3196 & ~n3197;
  assign n3199 = n447 & ~n2383;
  assign n3200 = n356 & ~n2391;
  assign n3201 = ~n3199 & ~n3200;
  assign n3202 = n3198 & n3201;
  assign n3203 = ~pi134  & ~n3202;
  assign n3204 = n311 & ~n2374;
  assign n3205 = n356 & ~n2330;
  assign n3206 = ~n3204 & ~n3205;
  assign n3207 = n402 & ~n2355;
  assign n3208 = n447 & ~n2338;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = n3206 & n3209;
  assign n3211 = pi134  & ~n3210;
  assign po63  = n3203 | n3211;
  assign n3213 = ~pi134  & ~n632;
  assign n3214 = pi134  & ~n450;
  assign po64  = n3213 | n3214;
  assign n3216 = ~pi134  & ~n1053;
  assign n3217 = pi134  & ~n845;
  assign po65  = n3216 | n3217;
  assign n3219 = ~pi134  & ~n1224;
  assign n3220 = pi134  & ~n1138;
  assign po66  = n3219 | n3220;
  assign n3222 = ~pi134  & ~n1518;
  assign n3223 = pi134  & ~n1373;
  assign po67  = n3222 | n3223;
  assign n3225 = ~pi134  & ~n1591;
  assign n3226 = pi134  & ~n1555;
  assign po68  = n3225 | n3226;
  assign n3228 = ~pi134  & ~n1664;
  assign n3229 = pi134  & ~n1628;
  assign po69  = n3228 | n3229;
  assign n3231 = ~pi134  & ~n1737;
  assign n3232 = pi134  & ~n1701;
  assign po70  = n3231 | n3232;
  assign n3234 = ~pi134  & ~n1810;
  assign n3235 = pi134  & ~n1774;
  assign po71  = n3234 | n3235;
  assign n3237 = ~pi134  & ~n1883;
  assign n3238 = pi134  & ~n1847;
  assign po72  = n3237 | n3238;
  assign n3240 = ~pi134  & ~n1956;
  assign n3241 = pi134  & ~n1920;
  assign po73  = n3240 | n3241;
  assign n3243 = ~pi134  & ~n2029;
  assign n3244 = pi134  & ~n1993;
  assign po74  = n3243 | n3244;
  assign n3246 = ~pi134  & ~n2102;
  assign n3247 = pi134  & ~n2066;
  assign po75  = n3246 | n3247;
  assign n3249 = ~pi134  & ~n2175;
  assign n3250 = pi134  & ~n2139;
  assign po76  = n3249 | n3250;
  assign n3252 = ~pi134  & ~n2248;
  assign n3253 = pi134  & ~n2212;
  assign po77  = n3252 | n3253;
  assign n3255 = ~pi134  & ~n2321;
  assign n3256 = pi134  & ~n2285;
  assign po78  = n3255 | n3256;
  assign n3258 = ~pi134  & ~n2394;
  assign n3259 = pi134  & ~n2358;
  assign po79  = n3258 | n3259;
  assign n3261 = ~pi134  & ~n2411;
  assign n3262 = pi134  & ~n2403;
  assign po80  = n3261 | n3262;
  assign n3264 = ~pi134  & ~n2428;
  assign n3265 = pi134  & ~n2420;
  assign po81  = n3264 | n3265;
  assign n3267 = ~pi134  & ~n2445;
  assign n3268 = pi134  & ~n2437;
  assign po82  = n3267 | n3268;
  assign n3270 = ~pi134  & ~n2462;
  assign n3271 = pi134  & ~n2454;
  assign po83  = n3270 | n3271;
  assign n3273 = ~pi134  & ~n2479;
  assign n3274 = pi134  & ~n2471;
  assign po84  = n3273 | n3274;
  assign n3276 = ~pi134  & ~n2496;
  assign n3277 = pi134  & ~n2488;
  assign po85  = n3276 | n3277;
  assign n3279 = ~pi134  & ~n2513;
  assign n3280 = pi134  & ~n2505;
  assign po86  = n3279 | n3280;
  assign n3282 = ~pi134  & ~n2530;
  assign n3283 = pi134  & ~n2522;
  assign po87  = n3282 | n3283;
  assign n3285 = ~pi134  & ~n2547;
  assign n3286 = pi134  & ~n2539;
  assign po88  = n3285 | n3286;
  assign n3288 = ~pi134  & ~n2564;
  assign n3289 = pi134  & ~n2556;
  assign po89  = n3288 | n3289;
  assign n3291 = ~pi134  & ~n2581;
  assign n3292 = pi134  & ~n2573;
  assign po90  = n3291 | n3292;
  assign n3294 = ~pi134  & ~n2598;
  assign n3295 = pi134  & ~n2590;
  assign po91  = n3294 | n3295;
  assign n3297 = ~pi134  & ~n2615;
  assign n3298 = pi134  & ~n2607;
  assign po92  = n3297 | n3298;
  assign n3300 = ~pi134  & ~n2632;
  assign n3301 = pi134  & ~n2624;
  assign po93  = n3300 | n3301;
  assign n3303 = ~pi134  & ~n2649;
  assign n3304 = pi134  & ~n2641;
  assign po94  = n3303 | n3304;
  assign n3306 = ~pi134  & ~n2666;
  assign n3307 = pi134  & ~n2658;
  assign po95  = n3306 | n3307;
  assign n3309 = ~pi134  & ~n2683;
  assign n3310 = pi134  & ~n2675;
  assign po96  = n3309 | n3310;
  assign n3312 = ~pi134  & ~n2700;
  assign n3313 = pi134  & ~n2692;
  assign po97  = n3312 | n3313;
  assign n3315 = ~pi134  & ~n2717;
  assign n3316 = pi134  & ~n2709;
  assign po98  = n3315 | n3316;
  assign n3318 = ~pi134  & ~n2734;
  assign n3319 = pi134  & ~n2726;
  assign po99  = n3318 | n3319;
  assign n3321 = ~pi134  & ~n2751;
  assign n3322 = pi134  & ~n2743;
  assign po100  = n3321 | n3322;
  assign n3324 = ~pi134  & ~n2768;
  assign n3325 = pi134  & ~n2760;
  assign po101  = n3324 | n3325;
  assign n3327 = ~pi134  & ~n2785;
  assign n3328 = pi134  & ~n2777;
  assign po102  = n3327 | n3328;
  assign n3330 = ~pi134  & ~n2802;
  assign n3331 = pi134  & ~n2794;
  assign po103  = n3330 | n3331;
  assign n3333 = ~pi134  & ~n2819;
  assign n3334 = pi134  & ~n2811;
  assign po104  = n3333 | n3334;
  assign n3336 = ~pi134  & ~n2836;
  assign n3337 = pi134  & ~n2828;
  assign po105  = n3336 | n3337;
  assign n3339 = ~pi134  & ~n2853;
  assign n3340 = pi134  & ~n2845;
  assign po106  = n3339 | n3340;
  assign n3342 = ~pi134  & ~n2870;
  assign n3343 = pi134  & ~n2862;
  assign po107  = n3342 | n3343;
  assign n3345 = ~pi134  & ~n2887;
  assign n3346 = pi134  & ~n2879;
  assign po108  = n3345 | n3346;
  assign n3348 = ~pi134  & ~n2904;
  assign n3349 = pi134  & ~n2896;
  assign po109  = n3348 | n3349;
  assign n3351 = ~pi134  & ~n2921;
  assign n3352 = pi134  & ~n2913;
  assign po110  = n3351 | n3352;
  assign n3354 = ~pi134  & ~n2938;
  assign n3355 = pi134  & ~n2930;
  assign po111  = n3354 | n3355;
  assign n3357 = ~pi134  & ~n2955;
  assign n3358 = pi134  & ~n2947;
  assign po112  = n3357 | n3358;
  assign n3360 = ~pi134  & ~n2972;
  assign n3361 = pi134  & ~n2964;
  assign po113  = n3360 | n3361;
  assign n3363 = ~pi134  & ~n2989;
  assign n3364 = pi134  & ~n2981;
  assign po114  = n3363 | n3364;
  assign n3366 = ~pi134  & ~n3006;
  assign n3367 = pi134  & ~n2998;
  assign po115  = n3366 | n3367;
  assign n3369 = ~pi134  & ~n3023;
  assign n3370 = pi134  & ~n3015;
  assign po116  = n3369 | n3370;
  assign n3372 = ~pi134  & ~n3040;
  assign n3373 = pi134  & ~n3032;
  assign po117  = n3372 | n3373;
  assign n3375 = ~pi134  & ~n3057;
  assign n3376 = pi134  & ~n3049;
  assign po118  = n3375 | n3376;
  assign n3378 = ~pi134  & ~n3074;
  assign n3379 = pi134  & ~n3066;
  assign po119  = n3378 | n3379;
  assign n3381 = ~pi134  & ~n3091;
  assign n3382 = pi134  & ~n3083;
  assign po120  = n3381 | n3382;
  assign n3384 = ~pi134  & ~n3108;
  assign n3385 = pi134  & ~n3100;
  assign po121  = n3384 | n3385;
  assign n3387 = ~pi134  & ~n3125;
  assign n3388 = pi134  & ~n3117;
  assign po122  = n3387 | n3388;
  assign n3390 = ~pi134  & ~n3142;
  assign n3391 = pi134  & ~n3134;
  assign po123  = n3390 | n3391;
  assign n3393 = ~pi134  & ~n3159;
  assign n3394 = pi134  & ~n3151;
  assign po124  = n3393 | n3394;
  assign n3396 = ~pi134  & ~n3176;
  assign n3397 = pi134  & ~n3168;
  assign po125  = n3396 | n3397;
  assign n3399 = ~pi134  & ~n3193;
  assign n3400 = pi134  & ~n3185;
  assign po126  = n3399 | n3400;
  assign n3402 = ~pi134  & ~n3210;
  assign n3403 = pi134  & ~n3202;
  assign po127  = n3402 | n3403;
endmodule
