module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24 ;
  wire n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591,
    n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3626, n3627,
    n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651,
    n3652, n3653, n3654, n3655, n3656, n3657,
    n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681,
    n3682, n3683, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742,
    n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772,
    n3773, n3774, n3775, n3776, n3777, n3778,
    n3779, n3780, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790,
    n3791, n3792, n3793, n3794, n3795, n3796,
    n3797, n3798, n3799, n3800, n3801, n3802,
    n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3819, n3820,
    n3821, n3822, n3823, n3824, n3825, n3826,
    n3827, n3828, n3829, n3830, n3831, n3832,
    n3833, n3834, n3835, n3836, n3837, n3838,
    n3839, n3840, n3841, n3842, n3843, n3844,
    n3845, n3846, n3847, n3848, n3849, n3850,
    n3851, n3852, n3853, n3854, n3855, n3856,
    n3857, n3858, n3859, n3860, n3861, n3862,
    n3863, n3864, n3865, n3866, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881,
    n3882, n3883, n3884, n3885, n3886, n3887,
    n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3901, n3902, n3903, n3904, n3905,
    n3906, n3907, n3908, n3909, n3910, n3911,
    n3912, n3913, n3914, n3915, n3916, n3917,
    n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3934, n3935,
    n3936, n3937, n3938, n3939, n3940, n3941,
    n3942, n3943, n3944, n3945, n3946, n3947,
    n3948, n3949, n3950, n3951, n3952, n3953,
    n3954, n3955, n3956, n3957, n3958, n3959,
    n3960, n3961, n3962, n3963, n3964, n3965,
    n3966, n3967, n3968, n3969, n3970, n3971,
    n3972, n3973, n3974, n3975, n3976, n3977,
    n3978, n3979, n3980, n3981, n3982, n3983,
    n3984, n3985, n3986, n3987, n3989, n3990,
    n3991, n3992, n3993, n3994, n3995, n3996,
    n3997, n3998, n3999, n4000, n4001, n4002,
    n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014,
    n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4023, n4024, n4025, n4026,
    n4027, n4028, n4029, n4030, n4031, n4032,
    n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044,
    n4045, n4046, n4047, n4048, n4049, n4050,
    n4051, n4052, n4053, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4062,
    n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074,
    n4075, n4076, n4077, n4078, n4079, n4080,
    n4081, n4082, n4083, n4084, n4085, n4086,
    n4087, n4088, n4089, n4090, n4091, n4092,
    n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117,
    n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141,
    n4142, n4143, n4144, n4145, n4146, n4147,
    n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171,
    n4172, n4173, n4174, n4175, n4176, n4177,
    n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195,
    n4196, n4197, n4198, n4199, n4200, n4201,
    n4202, n4203, n4204, n4205, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292,
    n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4315, n4316, n4317,
    n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341,
    n4342, n4343, n4344, n4345, n4346, n4347,
    n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4375, n4376, n4377,
    n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395,
    n4396, n4397, n4398, n4399, n4400, n4401,
    n4402, n4403, n4404, n4405, n4406, n4407,
    n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4422, n4423, n4424, n4425, n4426,
    n4427, n4428, n4429, n4430, n4431, n4432,
    n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450,
    n4451, n4452, n4453, n4454, n4455, n4456,
    n4457, n4458, n4459, n4460, n4461, n4462,
    n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4479, n4480,
    n4481, n4482, n4483, n4484, n4485, n4486,
    n4487, n4488, n4489, n4490, n4491, n4492,
    n4493, n4494, n4495, n4496, n4497, n4498,
    n4499, n4500, n4501, n4502, n4503, n4504,
    n4505, n4506, n4507, n4508, n4509, n4510,
    n4511, n4512, n4514, n4515, n4516, n4517,
    n4518, n4519, n4520, n4521, n4522, n4523,
    n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535,
    n4536, n4537, n4538, n4539, n4540, n4541,
    n4542, n4543, n4544, n4545, n4546, n4547,
    n4548, n4549, n4550, n4551, n4552, n4553,
    n4554, n4555, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571,
    n4572, n4573, n4574, n4575, n4576, n4577,
    n4578, n4579, n4580, n4581, n4582, n4583,
    n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601,
    n4602, n4603, n4604, n4605, n4606, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662,
    n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845,
    n4846, n4847, n4848, n4849, n4850, n4851,
    n4852, n4853, n4854, n4855, n4856, n4857,
    n4858, n4859, n4860, n4861, n4862, n4863,
    n4864, n4865, n4866, n4867, n4868, n4869,
    n4870, n4871, n4872, n4873, n4874, n4875,
    n4876, n4877, n4878, n4879, n4880, n4881,
    n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4889, n4890, n4891, n4892, n4894,
    n4895, n4896, n4897, n4898, n4899, n4900,
    n4901, n4902, n4903, n4904, n4905, n4906,
    n4907, n4908, n4909, n4910, n4911, n4912,
    n4913, n4914, n4915, n4916, n4917, n4918,
    n4919, n4920, n4921, n4922, n4923, n4924,
    n4925, n4926, n4927, n4928, n4929, n4930,
    n4931, n4932, n4933, n4934, n4935, n4936,
    n4937, n4938, n4939, n4940, n4941, n4942,
    n4943, n4944, n4945, n4946, n4947, n4948,
    n4949, n4950, n4951, n4952, n4953, n4954,
    n4955, n4956, n4957, n4959, n4960, n4961,
    n4962, n4963, n4964, n4965, n4966, n4967,
    n4968, n4969, n4970, n4971, n4972, n4973,
    n4974, n4975, n4976, n4977, n4978, n4979,
    n4980, n4981, n4982, n4983, n4984, n4985,
    n4986, n4987, n4988, n4989, n4990, n4991,
    n4992, n4993, n4994, n4995, n4996, n4997,
    n4998, n4999, n5000, n5001, n5002, n5003,
    n5004, n5005, n5006, n5007, n5008, n5009,
    n5010, n5011, n5013, n5014, n5015, n5016,
    n5017, n5018, n5019, n5020, n5021, n5022,
    n5023, n5024, n5025, n5026, n5027, n5028,
    n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040,
    n5041, n5042, n5043, n5044, n5045, n5046,
    n5047, n5048, n5049, n5050, n5051, n5052,
    n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5144, n5145, n5146,
    n5147, n5148, n5149, n5150, n5151, n5152,
    n5153, n5154, n5155, n5156, n5157, n5158,
    n5159, n5160, n5161, n5162, n5163, n5164,
    n5165, n5167, n5168, n5169, n5170, n5171,
    n5172, n5173, n5174, n5175, n5176, n5177,
    n5178, n5179, n5180, n5181, n5182, n5183,
    n5184, n5185, n5186, n5188, n5189, n5190,
    n5191, n5192, n5193, n5194, n5195, n5196,
    n5197, n5198, n5199, n5200, n5201, n5202,
    n5203, n5205, n5206, n5207, n5208, n5209,
    n5210, n5211, n5212, n5213, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5225, n5226, n5227, n5228, n5229;
  assign n50 = ~pi1  & ~pi2 ;
  assign n51 = ~pi0  & n50;
  assign n52 = ~pi3  & n51;
  assign n53 = ~pi4  & n52;
  assign n54 = ~pi22  & ~n53;
  assign n55 = pi5  & ~n54;
  assign n56 = ~pi5  & n54;
  assign n57 = ~n55 & ~n56;
  assign n58 = ~pi5  & n53;
  assign n59 = ~pi6  & n58;
  assign n60 = ~pi22  & ~n59;
  assign n61 = pi7  & ~n60;
  assign n62 = ~pi7  & n60;
  assign n63 = ~n61 & ~n62;
  assign n64 = ~pi7  & n59;
  assign n65 = ~pi8  & n64;
  assign n66 = ~pi9  & n65;
  assign n67 = ~pi10  & n66;
  assign n68 = ~pi11  & n67;
  assign n69 = ~pi12  & n68;
  assign n70 = ~pi13  & n69;
  assign n71 = ~pi14  & n70;
  assign n72 = ~pi15  & n71;
  assign n73 = ~pi16  & n72;
  assign n74 = ~pi17  & n73;
  assign n75 = ~pi18  & n74;
  assign n76 = ~pi22  & ~n75;
  assign n77 = pi19  & ~n76;
  assign n78 = ~pi19  & n76;
  assign n79 = ~n77 & ~n78;
  assign n80 = pi18  & pi22 ;
  assign n81 = pi18  & ~n74;
  assign n82 = n76 & ~n81;
  assign n83 = ~n80 & ~n82;
  assign n84 = ~n79 & ~n83;
  assign n85 = ~pi22  & ~n73;
  assign n86 = pi17  & ~n85;
  assign n87 = ~pi17  & n85;
  assign n88 = ~n86 & ~n87;
  assign n89 = ~pi22  & ~n72;
  assign n90 = pi16  & ~n89;
  assign n91 = ~pi16  & n89;
  assign n92 = ~n90 & ~n91;
  assign n93 = ~n88 & ~n92;
  assign n94 = n84 & n93;
  assign n95 = pi15  & pi22 ;
  assign n96 = pi15  & ~n71;
  assign n97 = n89 & ~n96;
  assign n98 = ~n95 & ~n97;
  assign n99 = pi21  & pi22 ;
  assign n100 = ~pi19  & n75;
  assign n101 = ~pi20  & n100;
  assign n102 = ~pi21  & n101;
  assign n103 = pi21  & ~n101;
  assign n104 = ~pi22  & ~n103;
  assign n105 = ~n102 & n104;
  assign n106 = ~n99 & ~n105;
  assign n107 = pi20  & pi22 ;
  assign n108 = pi20  & ~n100;
  assign n109 = ~pi22  & ~n101;
  assign n110 = ~n108 & n109;
  assign n111 = ~n107 & ~n110;
  assign n112 = ~n106 & ~n111;
  assign n113 = n98 & n112;
  assign n114 = n94 & n113;
  assign n115 = ~n98 & n112;
  assign n116 = ~n88 & n92;
  assign n117 = n79 & n83;
  assign n118 = n116 & n117;
  assign n119 = n115 & n118;
  assign n120 = n79 & ~n83;
  assign n121 = n88 & ~n92;
  assign n122 = n120 & n121;
  assign n123 = n113 & n122;
  assign n124 = ~n106 & n111;
  assign n125 = ~n98 & n124;
  assign n126 = n116 & n120;
  assign n127 = n125 & n126;
  assign n128 = n98 & n124;
  assign n129 = n93 & n120;
  assign n130 = n128 & n129;
  assign n131 = ~n127 & ~n130;
  assign n132 = n115 & n122;
  assign n133 = n125 & n129;
  assign n134 = ~n132 & ~n133;
  assign n135 = n131 & n134;
  assign n136 = ~n79 & n83;
  assign n137 = n88 & n92;
  assign n138 = n136 & n137;
  assign n139 = n115 & n138;
  assign n140 = n113 & n138;
  assign n141 = n93 & n136;
  assign n142 = n128 & n141;
  assign n143 = ~n140 & ~n142;
  assign n144 = ~n139 & n143;
  assign n145 = n135 & n144;
  assign n146 = ~n123 & n145;
  assign n147 = n125 & n141;
  assign n148 = n121 & n136;
  assign n149 = n113 & n148;
  assign n150 = n113 & n126;
  assign n151 = ~n149 & ~n150;
  assign n152 = n116 & n136;
  assign n153 = n124 & n152;
  assign n154 = n151 & ~n153;
  assign n155 = ~n147 & n154;
  assign n156 = n146 & n155;
  assign n157 = ~n119 & n156;
  assign n158 = ~n114 & n157;
  assign n159 = n113 & n118;
  assign n160 = n84 & n116;
  assign n161 = n115 & n160;
  assign n162 = n117 & n121;
  assign n163 = n115 & n162;
  assign n164 = ~n161 & ~n163;
  assign n165 = ~n159 & n164;
  assign n166 = n94 & n115;
  assign n167 = n84 & n137;
  assign n168 = n115 & n167;
  assign n169 = n125 & n160;
  assign n170 = ~n168 & ~n169;
  assign n171 = n94 & n128;
  assign n172 = n113 & n167;
  assign n173 = n128 & n160;
  assign n174 = n115 & n141;
  assign n175 = ~n173 & ~n174;
  assign n176 = ~n172 & n175;
  assign n177 = ~n171 & n176;
  assign n178 = n170 & n177;
  assign n179 = ~n166 & n178;
  assign n180 = n165 & n179;
  assign n181 = n84 & n121;
  assign n182 = n113 & n181;
  assign n183 = n113 & n160;
  assign n184 = n117 & n137;
  assign n185 = n115 & n184;
  assign n186 = n94 & n125;
  assign n187 = n113 & n184;
  assign n188 = ~n186 & ~n187;
  assign n189 = ~n185 & n188;
  assign n190 = ~n183 & n189;
  assign n191 = ~n182 & n190;
  assign n192 = n113 & n162;
  assign n193 = n124 & n181;
  assign n194 = n98 & n193;
  assign n195 = n128 & n167;
  assign n196 = n93 & n117;
  assign n197 = n115 & n196;
  assign n198 = n125 & n167;
  assign n199 = n113 & n196;
  assign n200 = ~n198 & ~n199;
  assign n201 = ~n98 & n193;
  assign n202 = n200 & ~n201;
  assign n203 = ~n197 & n202;
  assign n204 = n115 & n152;
  assign n205 = n113 & n152;
  assign n206 = n113 & n141;
  assign n207 = ~n205 & ~n206;
  assign n208 = ~n204 & n207;
  assign n209 = n203 & n208;
  assign n210 = ~n195 & n209;
  assign n211 = ~n194 & n210;
  assign n212 = ~n192 & n211;
  assign n213 = n115 & n181;
  assign n214 = n115 & n148;
  assign n215 = ~n213 & ~n214;
  assign n216 = n212 & n215;
  assign n217 = n128 & n148;
  assign n218 = n115 & n126;
  assign n219 = n113 & n129;
  assign n220 = n120 & n137;
  assign n221 = n113 & n220;
  assign n222 = ~n219 & ~n221;
  assign n223 = ~n218 & n222;
  assign n224 = ~n217 & n223;
  assign n225 = n115 & n220;
  assign n226 = n125 & n138;
  assign n227 = n115 & n129;
  assign n228 = n128 & n138;
  assign n229 = ~n227 & ~n228;
  assign n230 = ~n226 & n229;
  assign n231 = ~n225 & n230;
  assign n232 = n125 & n148;
  assign n233 = n231 & ~n232;
  assign n234 = n224 & n233;
  assign n235 = n216 & n234;
  assign n236 = n191 & n235;
  assign n237 = n180 & n236;
  assign n238 = n158 & n237;
  assign n239 = ~n63 & ~n238;
  assign n240 = n118 & n125;
  assign n241 = n106 & n111;
  assign n242 = n98 & n241;
  assign n243 = n184 & n242;
  assign n244 = ~n232 & ~n243;
  assign n245 = ~n130 & ~n149;
  assign n246 = n106 & ~n111;
  assign n247 = n98 & n246;
  assign n248 = n122 & n247;
  assign n249 = n148 & n247;
  assign n250 = ~n213 & ~n249;
  assign n251 = ~n217 & n250;
  assign n252 = ~n248 & n251;
  assign n253 = n245 & n252;
  assign n254 = n148 & n242;
  assign n255 = n118 & n128;
  assign n256 = n94 & n247;
  assign n257 = ~n98 & n241;
  assign n258 = n138 & n257;
  assign n259 = ~n256 & ~n258;
  assign n260 = ~n255 & n259;
  assign n261 = ~n254 & n260;
  assign n262 = n196 & n257;
  assign n263 = n94 & n257;
  assign n264 = ~n98 & n246;
  assign n265 = n196 & n264;
  assign n266 = ~n263 & ~n265;
  assign n267 = ~n262 & n266;
  assign n268 = ~n197 & n267;
  assign n269 = n261 & n268;
  assign n270 = n94 & n242;
  assign n271 = n196 & n242;
  assign n272 = n230 & ~n271;
  assign n273 = ~n270 & n272;
  assign n274 = n152 & n247;
  assign n275 = ~n204 & ~n274;
  assign n276 = n273 & n275;
  assign n277 = n269 & n276;
  assign n278 = n253 & n277;
  assign n279 = n244 & n278;
  assign n280 = ~n240 & n279;
  assign n281 = n118 & n242;
  assign n282 = n160 & n257;
  assign n283 = n141 & n246;
  assign n284 = n98 & n283;
  assign n285 = ~n166 & ~n284;
  assign n286 = ~n282 & n285;
  assign n287 = n125 & n220;
  assign n288 = ~n147 & ~n218;
  assign n289 = ~n287 & n288;
  assign n290 = n286 & n289;
  assign n291 = ~n281 & n290;
  assign n292 = n280 & n291;
  assign n293 = n162 & n242;
  assign n294 = n220 & n264;
  assign n295 = n162 & n247;
  assign n296 = ~n294 & ~n295;
  assign n297 = n138 & n242;
  assign n298 = ~n225 & ~n297;
  assign n299 = ~n161 & n298;
  assign n300 = n296 & n299;
  assign n301 = ~n293 & n300;
  assign n302 = n162 & n264;
  assign n303 = n94 & n264;
  assign n304 = n138 & n247;
  assign n305 = n196 & n247;
  assign n306 = ~n304 & ~n305;
  assign n307 = ~n303 & n306;
  assign n308 = ~n119 & ~n183;
  assign n309 = ~n127 & n308;
  assign n310 = ~n171 & n309;
  assign n311 = n134 & n310;
  assign n312 = n307 & n311;
  assign n313 = ~n302 & n312;
  assign n314 = ~n198 & n313;
  assign n315 = ~n206 & n314;
  assign n316 = n129 & n257;
  assign n317 = n184 & n257;
  assign n318 = n167 & n242;
  assign n319 = ~n142 & ~n318;
  assign n320 = n98 & n153;
  assign n321 = n319 & ~n320;
  assign n322 = ~n192 & n321;
  assign n323 = ~n317 & n322;
  assign n324 = ~n316 & n323;
  assign n325 = n129 & n264;
  assign n326 = n126 & n264;
  assign n327 = n167 & n247;
  assign n328 = ~n326 & ~n327;
  assign n329 = ~n325 & n328;
  assign n330 = ~n114 & n329;
  assign n331 = n324 & n330;
  assign n332 = n118 & n257;
  assign n333 = n160 & n247;
  assign n334 = ~n182 & ~n333;
  assign n335 = ~n332 & n334;
  assign n336 = n129 & n242;
  assign n337 = n141 & n257;
  assign n338 = n125 & n184;
  assign n339 = n181 & n247;
  assign n340 = ~n338 & ~n339;
  assign n341 = ~n337 & n340;
  assign n342 = ~n336 & n341;
  assign n343 = n335 & n342;
  assign n344 = n331 & n343;
  assign n345 = n315 & n344;
  assign n346 = n167 & n257;
  assign n347 = ~n169 & ~n346;
  assign n348 = ~n98 & n153;
  assign n349 = n128 & n220;
  assign n350 = ~n195 & ~n349;
  assign n351 = n162 & n257;
  assign n352 = ~n185 & ~n351;
  assign n353 = n350 & n352;
  assign n354 = ~n348 & n353;
  assign n355 = n347 & n354;
  assign n356 = n345 & n355;
  assign n357 = ~n186 & n356;
  assign n358 = n301 & n357;
  assign n359 = n292 & n358;
  assign n360 = n220 & n247;
  assign n361 = n129 & n247;
  assign n362 = ~n195 & ~n361;
  assign n363 = ~n161 & n362;
  assign n364 = ~n360 & n363;
  assign n365 = n125 & n196;
  assign n366 = n148 & n264;
  assign n367 = ~n98 & n283;
  assign n368 = ~n366 & ~n367;
  assign n369 = ~n365 & n368;
  assign n370 = ~n320 & n369;
  assign n371 = ~n265 & n370;
  assign n372 = n364 & n371;
  assign n373 = n151 & n372;
  assign n374 = ~n249 & n373;
  assign n375 = ~n217 & n374;
  assign n376 = ~n119 & ~n225;
  assign n377 = ~n316 & n376;
  assign n378 = n122 & n128;
  assign n379 = n184 & n247;
  assign n380 = ~n282 & ~n379;
  assign n381 = n126 & n128;
  assign n382 = ~n174 & ~n381;
  assign n383 = n380 & n382;
  assign n384 = ~n378 & n383;
  assign n385 = n377 & n384;
  assign n386 = n152 & n257;
  assign n387 = ~n263 & ~n386;
  assign n388 = ~n338 & n387;
  assign n389 = n152 & n242;
  assign n390 = ~n169 & ~n228;
  assign n391 = ~n389 & n390;
  assign n392 = ~n130 & ~n305;
  assign n393 = n391 & n392;
  assign n394 = ~n182 & n393;
  assign n395 = n388 & n394;
  assign n396 = n385 & n395;
  assign n397 = n141 & n242;
  assign n398 = ~n284 & ~n326;
  assign n399 = ~n142 & n398;
  assign n400 = ~n287 & n399;
  assign n401 = ~n397 & n400;
  assign n402 = ~n270 & n401;
  assign n403 = n396 & n402;
  assign n404 = ~n140 & ~n168;
  assign n405 = ~n336 & n404;
  assign n406 = ~n173 & ~n339;
  assign n407 = n148 & n257;
  assign n408 = n181 & n264;
  assign n409 = ~n183 & ~n408;
  assign n410 = ~n172 & n409;
  assign n411 = ~n114 & n410;
  assign n412 = ~n159 & n411;
  assign n413 = ~n407 & n412;
  assign n414 = n184 & n264;
  assign n415 = n128 & n162;
  assign n416 = ~n186 & ~n415;
  assign n417 = ~n213 & n416;
  assign n418 = ~n414 & n417;
  assign n419 = n413 & n418;
  assign n420 = n406 & n419;
  assign n421 = ~n139 & ~n166;
  assign n422 = ~n192 & ~n221;
  assign n423 = n421 & n422;
  assign n424 = ~n194 & n423;
  assign n425 = ~n218 & n424;
  assign n426 = n261 & n425;
  assign n427 = n420 & n426;
  assign n428 = n405 & n427;
  assign n429 = ~n297 & n428;
  assign n430 = n403 & n429;
  assign n431 = n375 & n430;
  assign n432 = ~n359 & ~n431;
  assign n433 = ~n192 & ~n389;
  assign n434 = ~n339 & n433;
  assign n435 = ~n187 & n434;
  assign n436 = ~n197 & ~n360;
  assign n437 = ~n317 & n436;
  assign n438 = ~n318 & n437;
  assign n439 = n435 & n438;
  assign n440 = n181 & n242;
  assign n441 = ~n303 & ~n440;
  assign n442 = ~n228 & n441;
  assign n443 = ~n336 & n442;
  assign n444 = ~n333 & n443;
  assign n445 = n138 & n264;
  assign n446 = n126 & n257;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~n254 & n447;
  assign n449 = n122 & n257;
  assign n450 = n220 & n257;
  assign n451 = ~n349 & ~n450;
  assign n452 = ~n449 & n451;
  assign n453 = ~n199 & n452;
  assign n454 = n448 & n453;
  assign n455 = ~n139 & ~n219;
  assign n456 = ~n381 & n455;
  assign n457 = ~n195 & ~n248;
  assign n458 = ~n320 & n457;
  assign n459 = n456 & n458;
  assign n460 = n454 & n459;
  assign n461 = n444 & n460;
  assign n462 = n439 & n461;
  assign n463 = ~n173 & n462;
  assign n464 = ~n169 & n463;
  assign n465 = ~n185 & ~n225;
  assign n466 = ~n326 & n465;
  assign n467 = ~n221 & n466;
  assign n468 = n160 & n242;
  assign n469 = n167 & n264;
  assign n470 = n122 & n125;
  assign n471 = ~n287 & ~n470;
  assign n472 = ~n414 & n471;
  assign n473 = ~n469 & n472;
  assign n474 = ~n149 & n473;
  assign n475 = ~n468 & n474;
  assign n476 = n118 & n264;
  assign n477 = n126 & n247;
  assign n478 = ~n282 & ~n297;
  assign n479 = ~n477 & n478;
  assign n480 = ~n140 & ~n302;
  assign n481 = ~n249 & n480;
  assign n482 = n479 & n481;
  assign n483 = ~n476 & n482;
  assign n484 = ~n325 & ~n332;
  assign n485 = n483 & n484;
  assign n486 = ~n232 & ~n351;
  assign n487 = ~n274 & n486;
  assign n488 = ~n147 & n487;
  assign n489 = n485 & n488;
  assign n490 = n475 & n489;
  assign n491 = ~n227 & ~n305;
  assign n492 = ~n367 & n491;
  assign n493 = ~n133 & ~n397;
  assign n494 = ~n263 & n493;
  assign n495 = n492 & n494;
  assign n496 = n490 & n495;
  assign n497 = ~n262 & n496;
  assign n498 = n467 & n497;
  assign n499 = ~n240 & ~n415;
  assign n500 = ~n201 & n499;
  assign n501 = n498 & n500;
  assign n502 = n464 & n501;
  assign n503 = ~n432 & ~n502;
  assign n504 = n239 & ~n503;
  assign n505 = pi8  & pi22 ;
  assign n506 = ~pi22  & ~n65;
  assign n507 = pi8  & ~n64;
  assign n508 = n506 & ~n507;
  assign n509 = ~n505 & ~n508;
  assign n510 = ~n239 & n503;
  assign n511 = ~n504 & ~n510;
  assign n512 = ~n509 & n511;
  assign n513 = ~n238 & n512;
  assign n514 = ~n504 & ~n513;
  assign n515 = n118 & n247;
  assign n516 = n296 & ~n302;
  assign n517 = ~n305 & n516;
  assign n518 = ~n515 & n517;
  assign n519 = ~n265 & ~n476;
  assign n520 = ~n360 & n519;
  assign n521 = n518 & n520;
  assign n522 = ~n248 & n521;
  assign n523 = ~n349 & ~n378;
  assign n524 = n125 & n162;
  assign n525 = ~n240 & ~n524;
  assign n526 = ~n256 & ~n381;
  assign n527 = n525 & n526;
  assign n528 = ~n338 & n527;
  assign n529 = ~n327 & n528;
  assign n530 = ~n408 & ~n469;
  assign n531 = ~n339 & n530;
  assign n532 = n160 & n264;
  assign n533 = ~n283 & ~n532;
  assign n534 = n531 & n533;
  assign n535 = n128 & n184;
  assign n536 = ~n255 & ~n365;
  assign n537 = ~n535 & n536;
  assign n538 = n534 & n537;
  assign n539 = n128 & n196;
  assign n540 = ~n415 & ~n539;
  assign n541 = n152 & n264;
  assign n542 = ~n303 & ~n333;
  assign n543 = ~n541 & n542;
  assign n544 = n540 & n543;
  assign n545 = n538 & n544;
  assign n546 = n529 & n545;
  assign n547 = n471 & n546;
  assign n548 = n122 & n264;
  assign n549 = ~n361 & ~n548;
  assign n550 = ~n477 & n549;
  assign n551 = ~n249 & ~n445;
  assign n552 = n550 & n551;
  assign n553 = ~n304 & n552;
  assign n554 = ~n274 & ~n325;
  assign n555 = ~n326 & n554;
  assign n556 = ~n366 & n555;
  assign n557 = n553 & n556;
  assign n558 = n547 & n557;
  assign n559 = n523 & n558;
  assign n560 = n522 & n559;
  assign n561 = ~n258 & ~n389;
  assign n562 = n546 & n561;
  assign n563 = ~n254 & n562;
  assign n564 = ~n318 & ~n386;
  assign n565 = n141 & n241;
  assign n566 = ~n468 & n523;
  assign n567 = ~n440 & n566;
  assign n568 = n181 & n257;
  assign n569 = ~n346 & ~n568;
  assign n570 = ~n263 & n380;
  assign n571 = ~n270 & n472;
  assign n572 = n570 & n571;
  assign n573 = n569 & n572;
  assign n574 = n567 & n573;
  assign n575 = ~n565 & n574;
  assign n576 = n564 & n575;
  assign n577 = ~n407 & n576;
  assign n578 = n563 & n577;
  assign n579 = ~n560 & n578;
  assign n580 = n560 & ~n578;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~pi22  & ~n67;
  assign n583 = pi11  & ~n582;
  assign n584 = ~pi11  & n582;
  assign n585 = ~n583 & ~n584;
  assign n586 = ~n238 & ~n585;
  assign n587 = ~n581 & n586;
  assign n588 = pi10  & pi22 ;
  assign n589 = pi10  & ~n66;
  assign n590 = n582 & ~n589;
  assign n591 = ~n588 & ~n590;
  assign n592 = ~n560 & ~n578;
  assign n593 = ~n238 & ~n592;
  assign n594 = n581 & ~n593;
  assign n595 = n591 & n594;
  assign n596 = n238 & ~n581;
  assign n597 = n585 & n596;
  assign n598 = n560 & n578;
  assign n599 = n238 & ~n598;
  assign n600 = n581 & ~n599;
  assign n601 = ~n591 & n600;
  assign n602 = ~n597 & ~n601;
  assign n603 = ~n595 & n602;
  assign n604 = ~n587 & n603;
  assign n605 = ~n514 & n604;
  assign n606 = ~pi22  & ~n69;
  assign n607 = pi13  & ~n606;
  assign n608 = ~pi13  & n606;
  assign n609 = ~n607 & ~n608;
  assign n610 = ~n182 & ~n226;
  assign n611 = ~n201 & ~n217;
  assign n612 = ~n262 & n406;
  assign n613 = ~n568 & n612;
  assign n614 = n611 & n613;
  assign n615 = ~n337 & n614;
  assign n616 = ~n168 & ~n232;
  assign n617 = ~n248 & ~n532;
  assign n618 = ~n293 & n617;
  assign n619 = ~n240 & ~n449;
  assign n620 = ~n389 & n619;
  assign n621 = ~n271 & ~n524;
  assign n622 = n620 & n621;
  assign n623 = n618 & n622;
  assign n624 = ~n469 & n623;
  assign n625 = ~n476 & n624;
  assign n626 = n616 & n625;
  assign n627 = ~n351 & n626;
  assign n628 = ~n414 & n627;
  assign n629 = n615 & n628;
  assign n630 = n610 & n629;
  assign n631 = n164 & ~n199;
  assign n632 = ~n183 & n631;
  assign n633 = ~n361 & n632;
  assign n634 = n207 & ~n470;
  assign n635 = n122 & n242;
  assign n636 = ~n221 & n385;
  assign n637 = ~n635 & n636;
  assign n638 = n634 & n637;
  assign n639 = n554 & n638;
  assign n640 = n633 & n639;
  assign n641 = ~n297 & n640;
  assign n642 = ~n166 & n641;
  assign n643 = ~n114 & ~n294;
  assign n644 = ~n256 & ~n366;
  assign n645 = ~n198 & n644;
  assign n646 = ~n407 & n645;
  assign n647 = ~n194 & n646;
  assign n648 = ~n468 & n647;
  assign n649 = ~n305 & n648;
  assign n650 = ~n172 & ~n303;
  assign n651 = ~n214 & n650;
  assign n652 = ~n197 & n651;
  assign n653 = ~n204 & ~n255;
  assign n654 = ~n159 & n653;
  assign n655 = ~n320 & n654;
  assign n656 = ~n169 & n655;
  assign n657 = n652 & n656;
  assign n658 = ~n213 & ~n318;
  assign n659 = ~n327 & n658;
  assign n660 = n657 & n659;
  assign n661 = n649 & n660;
  assign n662 = n643 & n661;
  assign n663 = ~n515 & n662;
  assign n664 = n642 & n663;
  assign n665 = n630 & n664;
  assign n666 = n502 & ~n665;
  assign n667 = ~n502 & n665;
  assign n668 = ~n666 & ~n667;
  assign n669 = n502 & n665;
  assign n670 = n126 & n242;
  assign n671 = ~n332 & ~n670;
  assign n672 = n112 & n122;
  assign n673 = n671 & ~n672;
  assign n674 = ~n270 & n673;
  assign n675 = ~n381 & n674;
  assign n676 = ~n183 & n675;
  assign n677 = ~n193 & ~n337;
  assign n678 = ~n366 & ~n397;
  assign n679 = ~n142 & n678;
  assign n680 = ~n172 & ~n349;
  assign n681 = ~n213 & n680;
  assign n682 = ~n168 & n681;
  assign n683 = ~n414 & n682;
  assign n684 = n679 & n683;
  assign n685 = n677 & n684;
  assign n686 = ~n166 & ~n204;
  assign n687 = ~n174 & n686;
  assign n688 = ~n281 & n687;
  assign n689 = n685 & n688;
  assign n690 = n267 & n689;
  assign n691 = n676 & n690;
  assign n692 = ~n304 & ~n386;
  assign n693 = n643 & n692;
  assign n694 = ~n249 & n693;
  assign n695 = n691 & n694;
  assign n696 = ~n140 & ~n303;
  assign n697 = ~n365 & n696;
  assign n698 = n289 & ~n318;
  assign n699 = n697 & n698;
  assign n700 = ~n195 & ~n408;
  assign n701 = ~n378 & n700;
  assign n702 = ~n539 & n701;
  assign n703 = n699 & n702;
  assign n704 = ~n173 & ~n297;
  assign n705 = ~n348 & n704;
  assign n706 = ~n274 & n705;
  assign n707 = ~n470 & n706;
  assign n708 = ~n256 & ~n445;
  assign n709 = ~n379 & n708;
  assign n710 = n707 & n709;
  assign n711 = n703 & n710;
  assign n712 = ~n198 & ~n271;
  assign n713 = n151 & ~n227;
  assign n714 = ~n169 & n334;
  assign n715 = n713 & n714;
  assign n716 = ~n214 & n715;
  assign n717 = ~n161 & ~n316;
  assign n718 = n617 & n717;
  assign n719 = n207 & n718;
  assign n720 = ~n219 & n719;
  assign n721 = ~n446 & n720;
  assign n722 = n716 & n721;
  assign n723 = ~n139 & n722;
  assign n724 = ~n360 & n723;
  assign n725 = n712 & n724;
  assign n726 = ~n336 & n725;
  assign n727 = n711 & n726;
  assign n728 = n695 & n727;
  assign n729 = ~n669 & n728;
  assign n730 = n668 & ~n729;
  assign n731 = ~n609 & n730;
  assign n732 = ~n502 & ~n665;
  assign n733 = ~n728 & ~n732;
  assign n734 = n668 & ~n733;
  assign n735 = n609 & n734;
  assign n736 = ~n668 & ~n728;
  assign n737 = pi14  & pi22 ;
  assign n738 = pi14  & ~n70;
  assign n739 = ~pi22  & ~n71;
  assign n740 = ~n738 & n739;
  assign n741 = ~n737 & ~n740;
  assign n742 = n736 & ~n741;
  assign n743 = ~n668 & n728;
  assign n744 = n741 & n743;
  assign n745 = ~n742 & ~n744;
  assign n746 = ~n735 & n745;
  assign n747 = ~n731 & n746;
  assign n748 = n455 & ~n568;
  assign n749 = ~n446 & n654;
  assign n750 = ~n132 & ~n182;
  assign n751 = n416 & n750;
  assign n752 = ~n263 & n751;
  assign n753 = n749 & n752;
  assign n754 = ~n197 & n753;
  assign n755 = ~n524 & n754;
  assign n756 = n680 & n755;
  assign n757 = n748 & n756;
  assign n758 = ~n270 & n757;
  assign n759 = ~n336 & n758;
  assign n760 = ~n365 & ~n548;
  assign n761 = ~n440 & ~n535;
  assign n762 = n220 & n242;
  assign n763 = ~n346 & ~n539;
  assign n764 = ~n218 & ~n445;
  assign n765 = ~n450 & ~n468;
  assign n766 = ~n670 & n765;
  assign n767 = n764 & n766;
  assign n768 = ~n214 & n767;
  assign n769 = n151 & ~n477;
  assign n770 = ~n414 & n769;
  assign n771 = n768 & n770;
  assign n772 = n763 & n771;
  assign n773 = ~n287 & n772;
  assign n774 = ~n762 & n773;
  assign n775 = ~n140 & ~n304;
  assign n776 = ~n192 & n775;
  assign n777 = ~n338 & n776;
  assign n778 = ~n449 & n642;
  assign n779 = n777 & n778;
  assign n780 = ~n123 & ~n185;
  assign n781 = ~n366 & n780;
  assign n782 = ~n227 & n781;
  assign n783 = n779 & n782;
  assign n784 = n774 & n783;
  assign n785 = ~n240 & n250;
  assign n786 = ~n171 & ~n187;
  assign n787 = ~n114 & ~n326;
  assign n788 = n786 & n787;
  assign n789 = ~n168 & n788;
  assign n790 = n785 & n789;
  assign n791 = n784 & n790;
  assign n792 = n761 & n791;
  assign n793 = n760 & n792;
  assign n794 = n759 & n793;
  assign n795 = n728 & ~n794;
  assign n796 = ~n728 & n794;
  assign n797 = ~n795 & ~n796;
  assign n798 = n728 & n794;
  assign n799 = n578 & ~n798;
  assign n800 = n797 & ~n799;
  assign n801 = ~n585 & n800;
  assign n802 = ~n728 & ~n794;
  assign n803 = ~n578 & ~n802;
  assign n804 = n797 & ~n803;
  assign n805 = n585 & n804;
  assign n806 = ~n578 & ~n797;
  assign n807 = pi12  & pi22 ;
  assign n808 = pi12  & ~n68;
  assign n809 = n606 & ~n808;
  assign n810 = ~n807 & ~n809;
  assign n811 = n806 & ~n810;
  assign n812 = n578 & ~n797;
  assign n813 = n810 & n812;
  assign n814 = ~n811 & ~n813;
  assign n815 = ~n805 & n814;
  assign n816 = ~n801 & n815;
  assign n817 = n747 & ~n816;
  assign n818 = ~n747 & n816;
  assign n819 = ~n817 & ~n818;
  assign n820 = ~n238 & ~n591;
  assign n821 = ~n581 & n820;
  assign n822 = pi9  & ~n506;
  assign n823 = ~pi9  & n506;
  assign n824 = ~n822 & ~n823;
  assign n825 = n594 & n824;
  assign n826 = n591 & n596;
  assign n827 = n600 & ~n824;
  assign n828 = ~n826 & ~n827;
  assign n829 = ~n825 & n828;
  assign n830 = ~n821 & n829;
  assign n831 = ~n819 & n830;
  assign n832 = n747 & n816;
  assign n833 = ~n831 & ~n832;
  assign n834 = n514 & ~n604;
  assign n835 = ~n605 & ~n834;
  assign n836 = ~n833 & n835;
  assign n837 = ~n605 & ~n836;
  assign n838 = ~n238 & ~n824;
  assign n839 = ~n733 & n838;
  assign n840 = n733 & ~n838;
  assign n841 = ~n839 & ~n840;
  assign n842 = n820 & n841;
  assign n843 = ~n820 & ~n841;
  assign n844 = ~n842 & ~n843;
  assign n845 = ~n837 & n844;
  assign n846 = n837 & ~n844;
  assign n847 = ~n845 & ~n846;
  assign n848 = n668 & ~n741;
  assign n849 = ~n733 & ~n848;
  assign n850 = ~n729 & n848;
  assign n851 = ~n849 & ~n850;
  assign n852 = ~n838 & n851;
  assign n853 = n838 & ~n851;
  assign n854 = ~n852 & ~n853;
  assign n855 = n800 & ~n810;
  assign n856 = n804 & n810;
  assign n857 = ~n609 & n806;
  assign n858 = n609 & n812;
  assign n859 = ~n857 & ~n858;
  assign n860 = ~n856 & n859;
  assign n861 = ~n855 & n860;
  assign n862 = n854 & n861;
  assign n863 = ~n852 & ~n862;
  assign n864 = ~n609 & n800;
  assign n865 = n609 & n804;
  assign n866 = ~n741 & n806;
  assign n867 = n741 & n812;
  assign n868 = ~n866 & ~n867;
  assign n869 = ~n865 & n868;
  assign n870 = ~n864 & n869;
  assign n871 = ~n238 & ~n810;
  assign n872 = ~n581 & n871;
  assign n873 = n585 & n594;
  assign n874 = n596 & n810;
  assign n875 = ~n585 & n600;
  assign n876 = ~n874 & ~n875;
  assign n877 = ~n873 & n876;
  assign n878 = ~n872 & n877;
  assign n879 = n870 & n878;
  assign n880 = ~n870 & ~n878;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n863 & n881;
  assign n883 = n863 & ~n881;
  assign n884 = ~n882 & ~n883;
  assign n885 = n847 & n884;
  assign n886 = ~n845 & ~n885;
  assign n887 = ~n839 & ~n842;
  assign n888 = ~n879 & ~n882;
  assign n889 = ~n887 & n888;
  assign n890 = n887 & ~n888;
  assign n891 = ~n889 & ~n890;
  assign n892 = ~n741 & n797;
  assign n893 = ~n803 & ~n892;
  assign n894 = ~n799 & n892;
  assign n895 = ~n893 & ~n894;
  assign n896 = ~n586 & n895;
  assign n897 = n586 & ~n895;
  assign n898 = ~n896 & ~n897;
  assign n899 = ~n238 & ~n609;
  assign n900 = ~n581 & n899;
  assign n901 = n594 & n810;
  assign n902 = n596 & n609;
  assign n903 = n600 & ~n810;
  assign n904 = ~n902 & ~n903;
  assign n905 = ~n901 & n904;
  assign n906 = ~n900 & n905;
  assign n907 = n898 & n906;
  assign n908 = ~n898 & ~n906;
  assign n909 = ~n907 & ~n908;
  assign n910 = ~n891 & ~n909;
  assign n911 = n891 & n909;
  assign n912 = ~n910 & ~n911;
  assign n913 = ~n886 & ~n912;
  assign n914 = ~n591 & n800;
  assign n915 = n591 & n804;
  assign n916 = ~n585 & n806;
  assign n917 = n585 & n812;
  assign n918 = ~n916 & ~n917;
  assign n919 = ~n915 & n918;
  assign n920 = ~n914 & n919;
  assign n921 = ~n581 & n838;
  assign n922 = n509 & n594;
  assign n923 = n596 & n824;
  assign n924 = ~n509 & n600;
  assign n925 = ~n923 & ~n924;
  assign n926 = ~n922 & n925;
  assign n927 = ~n921 & n926;
  assign n928 = n920 & n927;
  assign n929 = ~n920 & ~n927;
  assign n930 = ~n928 & ~n929;
  assign n931 = ~n258 & ~n325;
  assign n932 = ~n317 & n536;
  assign n933 = n931 & n932;
  assign n934 = ~n185 & n933;
  assign n935 = ~n195 & ~n515;
  assign n936 = ~n213 & n935;
  assign n937 = n934 & n936;
  assign n938 = n376 & n937;
  assign n939 = ~n476 & n938;
  assign n940 = ~n302 & ~n381;
  assign n941 = ~n295 & n940;
  assign n942 = ~n168 & ~n249;
  assign n943 = ~n539 & n942;
  assign n944 = ~n440 & n943;
  assign n945 = n941 & n944;
  assign n946 = n424 & n945;
  assign n947 = ~n303 & n946;
  assign n948 = ~n114 & n947;
  assign n949 = ~n386 & n617;
  assign n950 = ~n130 & n949;
  assign n951 = ~n173 & ~n338;
  assign n952 = ~n281 & n951;
  assign n953 = n950 & n952;
  assign n954 = n948 & n953;
  assign n955 = n674 & n954;
  assign n956 = ~n336 & n955;
  assign n957 = n939 & n956;
  assign n958 = ~n150 & ~n226;
  assign n959 = ~n287 & n680;
  assign n960 = ~n227 & n959;
  assign n961 = ~n469 & n960;
  assign n962 = ~n217 & n328;
  assign n963 = ~n337 & ~n445;
  assign n964 = n962 & n963;
  assign n965 = n619 & n964;
  assign n966 = n961 & n965;
  assign n967 = n958 & n966;
  assign n968 = ~n199 & n967;
  assign n969 = ~n407 & ~n762;
  assign n970 = ~n153 & ~n294;
  assign n971 = ~n282 & n970;
  assign n972 = ~n283 & n971;
  assign n973 = ~n541 & n972;
  assign n974 = n244 & n973;
  assign n975 = n969 & n974;
  assign n976 = ~n339 & n975;
  assign n977 = ~n169 & n976;
  assign n978 = n968 & n977;
  assign n979 = n957 & n978;
  assign n980 = n359 & n979;
  assign n981 = pi6  & pi22 ;
  assign n982 = pi6  & ~n58;
  assign n983 = n60 & ~n982;
  assign n984 = ~n981 & ~n983;
  assign n985 = ~n238 & ~n984;
  assign n986 = ~n123 & ~n333;
  assign n987 = ~n221 & n986;
  assign n988 = ~n327 & n987;
  assign n989 = n554 & n988;
  assign n990 = ~n197 & n989;
  assign n991 = ~n293 & n471;
  assign n992 = ~n316 & n991;
  assign n993 = ~n336 & ~n381;
  assign n994 = ~n163 & n993;
  assign n995 = ~n217 & n786;
  assign n996 = n352 & n995;
  assign n997 = n319 & n996;
  assign n998 = n994 & n997;
  assign n999 = ~n243 & n998;
  assign n1000 = ~n147 & n999;
  assign n1001 = n992 & n1000;
  assign n1002 = ~n226 & n1001;
  assign n1003 = ~n317 & n677;
  assign n1004 = ~n450 & n1003;
  assign n1005 = n391 & n1004;
  assign n1006 = n1002 & n1005;
  assign n1007 = n531 & n1006;
  assign n1008 = ~n206 & n1007;
  assign n1009 = n990 & n1008;
  assign n1010 = n441 & n1009;
  assign n1011 = ~n535 & n973;
  assign n1012 = ~n114 & n1011;
  assign n1013 = n134 & n748;
  assign n1014 = ~n305 & n1013;
  assign n1015 = ~n183 & n1014;
  assign n1016 = n1012 & n1015;
  assign n1017 = ~n635 & n1016;
  assign n1018 = ~n218 & n616;
  assign n1019 = ~n166 & n969;
  assign n1020 = n525 & n1019;
  assign n1021 = n1018 & n1020;
  assign n1022 = ~n205 & n299;
  assign n1023 = ~n366 & n1022;
  assign n1024 = n1021 & n1023;
  assign n1025 = n1017 & n1024;
  assign n1026 = ~n361 & ~n379;
  assign n1027 = ~n515 & n1026;
  assign n1028 = ~n360 & n760;
  assign n1029 = n1027 & n1028;
  assign n1030 = n151 & n1029;
  assign n1031 = ~n295 & n1030;
  assign n1032 = n1025 & n1031;
  assign n1033 = n1010 & n1032;
  assign n1034 = ~n979 & n1033;
  assign n1035 = ~n359 & n1034;
  assign n1036 = n985 & ~n1035;
  assign n1037 = ~n980 & ~n1036;
  assign n1038 = n930 & ~n1037;
  assign n1039 = ~n928 & ~n1038;
  assign n1040 = n359 & ~n431;
  assign n1041 = ~n359 & n431;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = ~n741 & n1042;
  assign n1044 = ~n503 & ~n1043;
  assign n1045 = n359 & n431;
  assign n1046 = n502 & ~n1045;
  assign n1047 = n1043 & ~n1046;
  assign n1048 = ~n1044 & ~n1047;
  assign n1049 = ~n239 & n1048;
  assign n1050 = n239 & ~n1048;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = n730 & ~n810;
  assign n1053 = n734 & n810;
  assign n1054 = ~n609 & n736;
  assign n1055 = n609 & n743;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = ~n1053 & n1056;
  assign n1058 = ~n1052 & n1057;
  assign n1059 = n1051 & n1058;
  assign n1060 = ~n1049 & ~n1059;
  assign n1061 = ~n1039 & ~n1060;
  assign n1062 = ~n1039 & n1060;
  assign n1063 = n1039 & ~n1060;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = ~n238 & ~n509;
  assign n1066 = ~n511 & ~n1065;
  assign n1067 = ~n513 & ~n1066;
  assign n1068 = ~n1064 & n1067;
  assign n1069 = ~n1061 & ~n1068;
  assign n1070 = ~n854 & ~n861;
  assign n1071 = ~n862 & ~n1070;
  assign n1072 = ~n1069 & n1071;
  assign n1073 = n1069 & ~n1071;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = n833 & ~n835;
  assign n1076 = ~n836 & ~n1075;
  assign n1077 = n1074 & n1076;
  assign n1078 = ~n1072 & ~n1077;
  assign n1079 = ~n847 & ~n884;
  assign n1080 = ~n885 & ~n1079;
  assign n1081 = ~n1078 & n1080;
  assign n1082 = ~n1074 & ~n1076;
  assign n1083 = ~n1077 & ~n1082;
  assign n1084 = n800 & ~n824;
  assign n1085 = n804 & n824;
  assign n1086 = ~n591 & n806;
  assign n1087 = n591 & n812;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = ~n1085 & n1088;
  assign n1090 = ~n1084 & n1089;
  assign n1091 = ~n238 & ~n581;
  assign n1092 = ~n509 & n1091;
  assign n1093 = n63 & n594;
  assign n1094 = n509 & n596;
  assign n1095 = ~n63 & n600;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = ~n1093 & n1096;
  assign n1098 = ~n1092 & n1097;
  assign n1099 = n1090 & ~n1098;
  assign n1100 = ~n1090 & n1098;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = n1042 & ~n1046;
  assign n1103 = ~n609 & n1102;
  assign n1104 = ~n503 & n1042;
  assign n1105 = n609 & n1104;
  assign n1106 = ~n502 & ~n1042;
  assign n1107 = ~n741 & n1106;
  assign n1108 = n502 & ~n1042;
  assign n1109 = n741 & n1108;
  assign n1110 = ~n1107 & ~n1109;
  assign n1111 = ~n1105 & n1110;
  assign n1112 = ~n1103 & n1111;
  assign n1113 = ~n1101 & n1112;
  assign n1114 = n1090 & n1098;
  assign n1115 = ~n1113 & ~n1114;
  assign n1116 = ~n1051 & ~n1058;
  assign n1117 = ~n1059 & ~n1116;
  assign n1118 = ~n1115 & n1117;
  assign n1119 = ~n930 & n1037;
  assign n1120 = ~n1038 & ~n1119;
  assign n1121 = n1115 & ~n1117;
  assign n1122 = ~n1118 & ~n1121;
  assign n1123 = n1120 & n1122;
  assign n1124 = ~n1118 & ~n1123;
  assign n1125 = n819 & n830;
  assign n1126 = ~n819 & ~n830;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = n1124 & n1127;
  assign n1129 = ~n1124 & ~n1127;
  assign n1130 = n1064 & ~n1067;
  assign n1131 = ~n1068 & ~n1130;
  assign n1132 = ~n1129 & ~n1131;
  assign n1133 = ~n1128 & ~n1132;
  assign n1134 = n1083 & n1133;
  assign n1135 = ~n585 & n730;
  assign n1136 = n585 & n734;
  assign n1137 = n736 & ~n810;
  assign n1138 = n743 & n810;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = ~n1136 & n1139;
  assign n1141 = ~n1135 & n1140;
  assign n1142 = ~n980 & ~n1035;
  assign n1143 = n985 & ~n1142;
  assign n1144 = ~n1036 & n1142;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = n1141 & ~n1145;
  assign n1147 = ~n57 & ~n238;
  assign n1148 = ~n979 & n1147;
  assign n1149 = n979 & ~n1147;
  assign n1150 = ~n1148 & ~n1149;
  assign n1151 = ~n979 & ~n1033;
  assign n1152 = ~n359 & ~n1151;
  assign n1153 = n979 & ~n1033;
  assign n1154 = ~n1034 & ~n1153;
  assign n1155 = ~n741 & n1154;
  assign n1156 = ~n1152 & ~n1155;
  assign n1157 = n979 & n1033;
  assign n1158 = n359 & ~n1157;
  assign n1159 = n1155 & ~n1158;
  assign n1160 = ~n1156 & ~n1159;
  assign n1161 = n1150 & n1160;
  assign n1162 = ~n1148 & ~n1161;
  assign n1163 = ~n1141 & n1145;
  assign n1164 = ~n1146 & ~n1163;
  assign n1165 = ~n1162 & n1164;
  assign n1166 = ~n1146 & ~n1165;
  assign n1167 = ~n810 & n1102;
  assign n1168 = n810 & n1104;
  assign n1169 = ~n609 & n1106;
  assign n1170 = n609 & n1108;
  assign n1171 = ~n1169 & ~n1170;
  assign n1172 = ~n1168 & n1171;
  assign n1173 = ~n1167 & n1172;
  assign n1174 = ~n591 & n730;
  assign n1175 = n591 & n734;
  assign n1176 = ~n585 & n736;
  assign n1177 = n585 & n743;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = ~n1175 & n1178;
  assign n1180 = ~n1174 & n1179;
  assign n1181 = n1173 & n1180;
  assign n1182 = n1173 & ~n1180;
  assign n1183 = ~n1173 & n1180;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = ~n509 & n800;
  assign n1186 = n509 & n804;
  assign n1187 = n806 & ~n824;
  assign n1188 = n812 & n824;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1186 & n1189;
  assign n1191 = ~n1185 & n1190;
  assign n1192 = ~n1184 & n1191;
  assign n1193 = ~n1181 & ~n1192;
  assign n1194 = n1101 & ~n1112;
  assign n1195 = ~n1113 & ~n1194;
  assign n1196 = ~n1193 & n1195;
  assign n1197 = pi4  & pi22 ;
  assign n1198 = pi4  & ~n52;
  assign n1199 = n54 & ~n1198;
  assign n1200 = ~n1197 & ~n1199;
  assign n1201 = ~n238 & ~n1200;
  assign n1202 = ~n979 & n1201;
  assign n1203 = n979 & ~n1201;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = n1154 & ~n1158;
  assign n1206 = ~n609 & n1205;
  assign n1207 = ~n1152 & n1154;
  assign n1208 = n609 & n1207;
  assign n1209 = ~n359 & ~n1154;
  assign n1210 = ~n741 & n1209;
  assign n1211 = n359 & ~n1154;
  assign n1212 = n741 & n1211;
  assign n1213 = ~n1210 & ~n1212;
  assign n1214 = ~n1208 & n1213;
  assign n1215 = ~n1206 & n1214;
  assign n1216 = n1204 & n1215;
  assign n1217 = ~n1202 & ~n1216;
  assign n1218 = n239 & ~n581;
  assign n1219 = n594 & n984;
  assign n1220 = n63 & n596;
  assign n1221 = n600 & ~n984;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = ~n1219 & n1222;
  assign n1224 = ~n1218 & n1223;
  assign n1225 = ~n1217 & n1224;
  assign n1226 = n1217 & ~n1224;
  assign n1227 = ~n1225 & ~n1226;
  assign n1228 = n730 & ~n824;
  assign n1229 = n734 & n824;
  assign n1230 = ~n591 & n736;
  assign n1231 = n591 & n743;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = ~n1229 & n1232;
  assign n1234 = ~n1228 & n1233;
  assign n1235 = ~n585 & n1102;
  assign n1236 = n585 & n1104;
  assign n1237 = ~n810 & n1106;
  assign n1238 = n810 & n1108;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = ~n1236 & n1239;
  assign n1241 = ~n1235 & n1240;
  assign n1242 = n1234 & n1241;
  assign n1243 = ~n1234 & n1241;
  assign n1244 = n1234 & ~n1241;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = ~n63 & n800;
  assign n1247 = n63 & n804;
  assign n1248 = ~n509 & n806;
  assign n1249 = n509 & n812;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = ~n1247 & n1250;
  assign n1252 = ~n1246 & n1251;
  assign n1253 = ~n1245 & n1252;
  assign n1254 = ~n1242 & ~n1253;
  assign n1255 = n1227 & ~n1254;
  assign n1256 = ~n1225 & ~n1255;
  assign n1257 = n1193 & ~n1195;
  assign n1258 = ~n1196 & ~n1257;
  assign n1259 = ~n1256 & n1258;
  assign n1260 = ~n1196 & ~n1259;
  assign n1261 = ~n1166 & ~n1260;
  assign n1262 = ~n1166 & n1260;
  assign n1263 = n1166 & ~n1260;
  assign n1264 = ~n1262 & ~n1263;
  assign n1265 = ~n1120 & ~n1122;
  assign n1266 = ~n1123 & ~n1265;
  assign n1267 = ~n1264 & n1266;
  assign n1268 = ~n1261 & ~n1267;
  assign n1269 = ~n1128 & ~n1129;
  assign n1270 = ~n1131 & n1269;
  assign n1271 = n1131 & ~n1269;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = ~n1268 & ~n1272;
  assign n1274 = ~n1264 & ~n1266;
  assign n1275 = n1264 & n1266;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = n1184 & n1191;
  assign n1278 = ~n1184 & ~n1191;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = ~n1150 & ~n1160;
  assign n1281 = ~n1161 & ~n1280;
  assign n1282 = ~n1279 & n1281;
  assign n1283 = n1279 & n1281;
  assign n1284 = ~n1279 & ~n1281;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = ~pi22  & ~n51;
  assign n1287 = pi3  & ~n1286;
  assign n1288 = ~pi3  & n1286;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = ~n238 & ~n1289;
  assign n1291 = ~n365 & ~n379;
  assign n1292 = ~n243 & ~n274;
  assign n1293 = n1291 & n1292;
  assign n1294 = ~n316 & n1293;
  assign n1295 = ~n346 & ~n414;
  assign n1296 = ~n338 & n1295;
  assign n1297 = ~n249 & n1296;
  assign n1298 = n1294 & n1297;
  assign n1299 = ~n548 & n1298;
  assign n1300 = ~n294 & n1299;
  assign n1301 = n209 & n765;
  assign n1302 = ~n762 & n1301;
  assign n1303 = ~n123 & n1302;
  assign n1304 = n1300 & n1303;
  assign n1305 = ~n449 & n1304;
  assign n1306 = ~n265 & n390;
  assign n1307 = ~n140 & n1306;
  assign n1308 = ~n185 & n1307;
  assign n1309 = ~n218 & ~n320;
  assign n1310 = ~n305 & n1309;
  assign n1311 = n164 & n1310;
  assign n1312 = ~n194 & n761;
  assign n1313 = ~n270 & n1312;
  assign n1314 = n1311 & n1313;
  assign n1315 = n702 & n1314;
  assign n1316 = n1308 & n1315;
  assign n1317 = ~n240 & n621;
  assign n1318 = ~n256 & ~n281;
  assign n1319 = n1317 & n1318;
  assign n1320 = ~n142 & n1319;
  assign n1321 = ~n132 & ~n303;
  assign n1322 = ~n232 & n1321;
  assign n1323 = ~n336 & n1322;
  assign n1324 = n1320 & n1323;
  assign n1325 = ~n293 & n1324;
  assign n1326 = ~n172 & n1325;
  assign n1327 = n1316 & n1326;
  assign n1328 = n1305 & n1327;
  assign n1329 = ~n979 & ~n1328;
  assign n1330 = n741 & ~n979;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = n1290 & ~n1331;
  assign n1333 = ~n1290 & n1331;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n810 & n1205;
  assign n1336 = n810 & n1207;
  assign n1337 = ~n609 & n1209;
  assign n1338 = n609 & n1211;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = ~n1336 & n1339;
  assign n1341 = ~n1335 & n1340;
  assign n1342 = n1334 & n1341;
  assign n1343 = ~n1332 & ~n1342;
  assign n1344 = ~n581 & n985;
  assign n1345 = n57 & n594;
  assign n1346 = n596 & n984;
  assign n1347 = ~n57 & n600;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = ~n1345 & n1348;
  assign n1350 = ~n1344 & n1349;
  assign n1351 = ~n1343 & n1350;
  assign n1352 = n1343 & ~n1350;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = ~n509 & n730;
  assign n1355 = n509 & n734;
  assign n1356 = n736 & ~n824;
  assign n1357 = n743 & n824;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = ~n1355 & n1358;
  assign n1360 = ~n1354 & n1359;
  assign n1361 = ~n591 & n1102;
  assign n1362 = n591 & n1104;
  assign n1363 = ~n585 & n1106;
  assign n1364 = n585 & n1108;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = ~n1362 & n1365;
  assign n1367 = ~n1361 & n1366;
  assign n1368 = n1360 & n1367;
  assign n1369 = ~n1360 & n1367;
  assign n1370 = n1360 & ~n1367;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = n800 & ~n984;
  assign n1373 = n804 & n984;
  assign n1374 = ~n63 & n806;
  assign n1375 = n63 & n812;
  assign n1376 = ~n1374 & ~n1375;
  assign n1377 = ~n1373 & n1376;
  assign n1378 = ~n1372 & n1377;
  assign n1379 = ~n1371 & n1378;
  assign n1380 = ~n1368 & ~n1379;
  assign n1381 = n1353 & ~n1380;
  assign n1382 = ~n1351 & ~n1381;
  assign n1383 = ~n1285 & ~n1382;
  assign n1384 = ~n1282 & ~n1383;
  assign n1385 = n1162 & ~n1164;
  assign n1386 = ~n1165 & ~n1385;
  assign n1387 = ~n1384 & n1386;
  assign n1388 = n1384 & ~n1386;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = n1256 & ~n1258;
  assign n1391 = ~n1259 & ~n1390;
  assign n1392 = n1389 & n1391;
  assign n1393 = ~n1387 & ~n1392;
  assign n1394 = ~n1276 & ~n1393;
  assign n1395 = ~n741 & ~n1328;
  assign n1396 = ~n979 & n1395;
  assign n1397 = ~n609 & n1328;
  assign n1398 = n979 & ~n1395;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = ~n1396 & n1399;
  assign n1401 = ~n581 & ~n1289;
  assign n1402 = n593 & ~n1401;
  assign n1403 = n1400 & n1402;
  assign n1404 = ~n581 & n1147;
  assign n1405 = n594 & n1200;
  assign n1406 = n57 & n596;
  assign n1407 = n600 & ~n1200;
  assign n1408 = ~n1406 & ~n1407;
  assign n1409 = ~n1405 & n1408;
  assign n1410 = ~n1404 & n1409;
  assign n1411 = n1403 & n1410;
  assign n1412 = ~n63 & n730;
  assign n1413 = n63 & n734;
  assign n1414 = ~n509 & n736;
  assign n1415 = n509 & n743;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = ~n1413 & n1416;
  assign n1418 = ~n1412 & n1417;
  assign n1419 = ~n57 & n800;
  assign n1420 = n57 & n804;
  assign n1421 = n806 & ~n984;
  assign n1422 = n812 & n984;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = ~n1420 & n1423;
  assign n1425 = ~n1419 & n1424;
  assign n1426 = n1418 & ~n1425;
  assign n1427 = ~n1418 & n1425;
  assign n1428 = ~n1426 & ~n1427;
  assign n1429 = ~n824 & n1102;
  assign n1430 = n824 & n1104;
  assign n1431 = ~n591 & n1106;
  assign n1432 = n591 & n1108;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = ~n1430 & n1433;
  assign n1435 = ~n1429 & n1434;
  assign n1436 = ~n1428 & n1435;
  assign n1437 = n1418 & n1425;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = ~n1403 & ~n1410;
  assign n1440 = ~n1411 & ~n1439;
  assign n1441 = ~n1438 & n1440;
  assign n1442 = ~n1411 & ~n1441;
  assign n1443 = ~n1204 & ~n1215;
  assign n1444 = ~n1216 & ~n1443;
  assign n1445 = ~n1442 & n1444;
  assign n1446 = n1245 & n1252;
  assign n1447 = ~n1245 & ~n1252;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = n1442 & ~n1444;
  assign n1450 = ~n1445 & ~n1449;
  assign n1451 = ~n1448 & n1450;
  assign n1452 = ~n1445 & ~n1451;
  assign n1453 = ~n1227 & n1254;
  assign n1454 = ~n1255 & ~n1453;
  assign n1455 = ~n1452 & n1454;
  assign n1456 = n1285 & ~n1382;
  assign n1457 = ~n1285 & n1382;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = n1452 & ~n1454;
  assign n1460 = ~n1455 & ~n1459;
  assign n1461 = ~n1458 & n1460;
  assign n1462 = ~n1455 & ~n1461;
  assign n1463 = ~n1389 & ~n1391;
  assign n1464 = ~n1392 & ~n1463;
  assign n1465 = ~n1462 & n1464;
  assign n1466 = ~n1353 & n1380;
  assign n1467 = ~n1381 & ~n1466;
  assign n1468 = ~n585 & n1205;
  assign n1469 = n585 & n1207;
  assign n1470 = ~n810 & n1209;
  assign n1471 = n810 & n1211;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = ~n1469 & n1472;
  assign n1474 = ~n1468 & n1473;
  assign n1475 = ~n581 & n1201;
  assign n1476 = n594 & n1289;
  assign n1477 = n596 & n1200;
  assign n1478 = n600 & ~n1289;
  assign n1479 = ~n1477 & ~n1478;
  assign n1480 = ~n1476 & n1479;
  assign n1481 = ~n1475 & n1480;
  assign n1482 = n1474 & n1481;
  assign n1483 = ~n1400 & ~n1402;
  assign n1484 = ~n1403 & ~n1483;
  assign n1485 = ~n1474 & ~n1481;
  assign n1486 = ~n1482 & ~n1485;
  assign n1487 = n1484 & n1486;
  assign n1488 = ~n1482 & ~n1487;
  assign n1489 = ~n1334 & ~n1341;
  assign n1490 = ~n1342 & ~n1489;
  assign n1491 = ~n1488 & n1490;
  assign n1492 = n1488 & ~n1490;
  assign n1493 = n1371 & n1378;
  assign n1494 = ~n1371 & ~n1378;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = ~n1492 & ~n1495;
  assign n1497 = ~n1491 & ~n1496;
  assign n1498 = n1467 & ~n1497;
  assign n1499 = ~n1467 & n1497;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = n1448 & ~n1450;
  assign n1502 = ~n1451 & ~n1501;
  assign n1503 = n1500 & n1502;
  assign n1504 = ~n1498 & ~n1503;
  assign n1505 = n1458 & ~n1460;
  assign n1506 = ~n1461 & ~n1505;
  assign n1507 = ~n1504 & n1506;
  assign n1508 = ~n797 & ~n1289;
  assign n1509 = n803 & ~n1508;
  assign n1510 = ~n810 & ~n1328;
  assign n1511 = ~n979 & n1510;
  assign n1512 = ~n585 & n1328;
  assign n1513 = n979 & ~n1510;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = ~n1511 & n1514;
  assign n1516 = n1509 & n1515;
  assign n1517 = ~n509 & n1102;
  assign n1518 = n509 & n1104;
  assign n1519 = ~n824 & n1106;
  assign n1520 = n824 & n1108;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = ~n1518 & n1521;
  assign n1523 = ~n1517 & n1522;
  assign n1524 = n730 & ~n984;
  assign n1525 = n734 & n984;
  assign n1526 = ~n63 & n736;
  assign n1527 = n63 & n743;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = ~n1525 & n1528;
  assign n1530 = ~n1524 & n1529;
  assign n1531 = n1523 & ~n1530;
  assign n1532 = ~n1523 & n1530;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = n1516 & ~n1533;
  assign n1535 = n1523 & n1530;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = ~n609 & ~n1328;
  assign n1538 = ~n979 & n1537;
  assign n1539 = ~n810 & n1328;
  assign n1540 = n979 & ~n1537;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = ~n1538 & n1541;
  assign n1543 = ~n591 & n1205;
  assign n1544 = n591 & n1207;
  assign n1545 = ~n585 & n1209;
  assign n1546 = n585 & n1211;
  assign n1547 = ~n1545 & ~n1546;
  assign n1548 = ~n1544 & n1547;
  assign n1549 = ~n1543 & n1548;
  assign n1550 = n1542 & ~n1549;
  assign n1551 = ~n1542 & n1549;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = n800 & ~n1200;
  assign n1554 = n804 & n1200;
  assign n1555 = ~n57 & n806;
  assign n1556 = n57 & n812;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = ~n1554 & n1557;
  assign n1559 = ~n1553 & n1558;
  assign n1560 = ~n1552 & n1559;
  assign n1561 = n1542 & n1549;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = ~n1536 & ~n1562;
  assign n1564 = ~n1536 & n1562;
  assign n1565 = n1536 & ~n1562;
  assign n1566 = ~n1564 & ~n1565;
  assign n1567 = n1428 & n1435;
  assign n1568 = ~n1428 & ~n1435;
  assign n1569 = ~n1567 & ~n1568;
  assign n1570 = ~n1566 & ~n1569;
  assign n1571 = ~n1563 & ~n1570;
  assign n1572 = n1438 & ~n1440;
  assign n1573 = ~n1441 & ~n1572;
  assign n1574 = ~n1571 & n1573;
  assign n1575 = n1571 & ~n1573;
  assign n1576 = ~n1574 & ~n1575;
  assign n1577 = ~n1491 & ~n1492;
  assign n1578 = ~n1495 & n1577;
  assign n1579 = n1495 & ~n1577;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = n1576 & n1580;
  assign n1582 = ~n1574 & ~n1581;
  assign n1583 = ~n1500 & ~n1502;
  assign n1584 = ~n1503 & ~n1583;
  assign n1585 = ~n1582 & n1584;
  assign n1586 = n1566 & n1569;
  assign n1587 = ~n1570 & ~n1586;
  assign n1588 = ~n824 & n1205;
  assign n1589 = n824 & n1207;
  assign n1590 = ~n591 & n1209;
  assign n1591 = n591 & n1211;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = ~n1589 & n1592;
  assign n1594 = ~n1588 & n1593;
  assign n1595 = ~n57 & n730;
  assign n1596 = n57 & n734;
  assign n1597 = n736 & ~n984;
  assign n1598 = n743 & n984;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = ~n1596 & n1599;
  assign n1601 = ~n1595 & n1600;
  assign n1602 = n1594 & ~n1601;
  assign n1603 = ~n1594 & n1601;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = ~n63 & n1102;
  assign n1606 = n63 & n1104;
  assign n1607 = ~n509 & n1106;
  assign n1608 = n509 & n1108;
  assign n1609 = ~n1607 & ~n1608;
  assign n1610 = ~n1606 & n1609;
  assign n1611 = ~n1605 & n1610;
  assign n1612 = ~n1604 & n1611;
  assign n1613 = n1594 & n1601;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615 = n1401 & ~n1614;
  assign n1616 = ~n1516 & n1533;
  assign n1617 = ~n1534 & ~n1616;
  assign n1618 = ~n1401 & n1614;
  assign n1619 = ~n1615 & ~n1618;
  assign n1620 = n1617 & n1619;
  assign n1621 = ~n1615 & ~n1620;
  assign n1622 = n1484 & ~n1486;
  assign n1623 = ~n1484 & n1486;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = ~n1621 & ~n1624;
  assign n1626 = n1621 & n1624;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = n1587 & n1627;
  assign n1629 = ~n1625 & ~n1628;
  assign n1630 = ~n1576 & ~n1580;
  assign n1631 = ~n1581 & ~n1630;
  assign n1632 = ~n1629 & n1631;
  assign n1633 = n1629 & ~n1631;
  assign n1634 = ~n1632 & ~n1633;
  assign n1635 = ~n591 & ~n1328;
  assign n1636 = ~n979 & n1635;
  assign n1637 = ~n824 & n1328;
  assign n1638 = n979 & ~n1635;
  assign n1639 = ~n1637 & ~n1638;
  assign n1640 = ~n1636 & n1639;
  assign n1641 = ~n668 & ~n1289;
  assign n1642 = n733 & ~n1641;
  assign n1643 = n1640 & n1642;
  assign n1644 = n730 & ~n1200;
  assign n1645 = n734 & n1200;
  assign n1646 = ~n57 & n736;
  assign n1647 = n57 & n743;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = ~n1645 & n1648;
  assign n1650 = ~n1644 & n1649;
  assign n1651 = n1643 & n1650;
  assign n1652 = n1643 & ~n1650;
  assign n1653 = ~n1643 & n1650;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = n1508 & ~n1654;
  assign n1656 = ~n1651 & ~n1655;
  assign n1657 = n1604 & ~n1611;
  assign n1658 = ~n1612 & ~n1657;
  assign n1659 = ~n1656 & n1658;
  assign n1660 = n1656 & ~n1658;
  assign n1661 = ~n1659 & ~n1660;
  assign n1662 = ~n585 & ~n1328;
  assign n1663 = ~n979 & n1662;
  assign n1664 = ~n591 & n1328;
  assign n1665 = n979 & ~n1662;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = ~n1663 & n1666;
  assign n1668 = ~n509 & n1205;
  assign n1669 = n509 & n1207;
  assign n1670 = ~n824 & n1209;
  assign n1671 = n824 & n1211;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = ~n1669 & n1672;
  assign n1674 = ~n1668 & n1673;
  assign n1675 = n1667 & n1674;
  assign n1676 = n1667 & ~n1674;
  assign n1677 = ~n1667 & n1674;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = ~n984 & n1102;
  assign n1680 = n984 & n1104;
  assign n1681 = ~n63 & n1106;
  assign n1682 = n63 & n1108;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = ~n1680 & n1683;
  assign n1685 = ~n1679 & n1684;
  assign n1686 = ~n1678 & n1685;
  assign n1687 = ~n1675 & ~n1686;
  assign n1688 = ~n1509 & ~n1515;
  assign n1689 = ~n1516 & ~n1688;
  assign n1690 = n800 & ~n1289;
  assign n1691 = n804 & n1289;
  assign n1692 = n806 & ~n1200;
  assign n1693 = n812 & n1200;
  assign n1694 = ~n1692 & ~n1693;
  assign n1695 = ~n1691 & n1694;
  assign n1696 = ~n1690 & n1695;
  assign n1697 = ~n1689 & n1696;
  assign n1698 = n1689 & ~n1696;
  assign n1699 = ~n1697 & ~n1698;
  assign n1700 = ~n1687 & ~n1699;
  assign n1701 = n1687 & n1699;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = n1661 & n1702;
  assign n1704 = ~n1659 & ~n1703;
  assign n1705 = ~n1661 & ~n1702;
  assign n1706 = ~n1703 & ~n1705;
  assign n1707 = ~n63 & n1205;
  assign n1708 = n63 & n1207;
  assign n1709 = ~n509 & n1209;
  assign n1710 = n509 & n1211;
  assign n1711 = ~n1709 & ~n1710;
  assign n1712 = ~n1708 & n1711;
  assign n1713 = ~n1707 & n1712;
  assign n1714 = ~n57 & n1102;
  assign n1715 = n57 & n1104;
  assign n1716 = ~n984 & n1106;
  assign n1717 = n984 & n1108;
  assign n1718 = ~n1716 & ~n1717;
  assign n1719 = ~n1715 & n1718;
  assign n1720 = ~n1714 & n1719;
  assign n1721 = n1713 & ~n1720;
  assign n1722 = ~n1713 & n1720;
  assign n1723 = ~n1721 & ~n1722;
  assign n1724 = n730 & ~n1289;
  assign n1725 = n734 & n1289;
  assign n1726 = n736 & ~n1200;
  assign n1727 = n743 & n1200;
  assign n1728 = ~n1726 & ~n1727;
  assign n1729 = ~n1725 & n1728;
  assign n1730 = ~n1724 & n1729;
  assign n1731 = ~n1723 & n1730;
  assign n1732 = n1713 & n1720;
  assign n1733 = ~n1731 & ~n1732;
  assign n1734 = n1678 & ~n1685;
  assign n1735 = ~n1686 & ~n1734;
  assign n1736 = ~n1733 & n1735;
  assign n1737 = ~n1508 & n1654;
  assign n1738 = ~n1655 & ~n1737;
  assign n1739 = n1733 & ~n1735;
  assign n1740 = ~n1736 & ~n1739;
  assign n1741 = n1738 & n1740;
  assign n1742 = ~n1736 & ~n1741;
  assign n1743 = ~n1640 & ~n1642;
  assign n1744 = ~n1643 & ~n1743;
  assign n1745 = ~n984 & n1205;
  assign n1746 = n984 & n1207;
  assign n1747 = ~n63 & n1209;
  assign n1748 = n63 & n1211;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = ~n1746 & n1749;
  assign n1751 = ~n1745 & n1750;
  assign n1752 = ~n824 & ~n1328;
  assign n1753 = ~n979 & n1752;
  assign n1754 = ~n509 & n1328;
  assign n1755 = n979 & ~n1752;
  assign n1756 = ~n1754 & ~n1755;
  assign n1757 = ~n1753 & n1756;
  assign n1758 = ~n1751 & n1757;
  assign n1759 = n1751 & ~n1757;
  assign n1760 = ~n1758 & ~n1759;
  assign n1761 = n1102 & ~n1200;
  assign n1762 = n1104 & n1200;
  assign n1763 = ~n57 & n1106;
  assign n1764 = n57 & n1108;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = ~n1762 & n1765;
  assign n1767 = ~n1761 & n1766;
  assign n1768 = ~n1760 & n1767;
  assign n1769 = n1751 & n1757;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = n1744 & ~n1770;
  assign n1772 = n1723 & n1730;
  assign n1773 = ~n1723 & ~n1730;
  assign n1774 = ~n1772 & ~n1773;
  assign n1775 = ~n1744 & n1770;
  assign n1776 = ~n1771 & ~n1775;
  assign n1777 = ~n1774 & n1776;
  assign n1778 = ~n1771 & ~n1777;
  assign n1779 = ~n57 & n1205;
  assign n1780 = n57 & n1207;
  assign n1781 = ~n984 & n1209;
  assign n1782 = n984 & n1211;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = ~n1780 & n1783;
  assign n1785 = ~n1779 & n1784;
  assign n1786 = n1102 & ~n1289;
  assign n1787 = n1104 & n1289;
  assign n1788 = n1106 & ~n1200;
  assign n1789 = n1108 & n1200;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~n1787 & n1790;
  assign n1792 = ~n1786 & n1791;
  assign n1793 = n1785 & n1792;
  assign n1794 = ~n1042 & ~n1289;
  assign n1795 = n503 & ~n1794;
  assign n1796 = ~n509 & ~n1328;
  assign n1797 = ~n979 & n1796;
  assign n1798 = ~n63 & n1328;
  assign n1799 = n979 & ~n1796;
  assign n1800 = ~n1798 & ~n1799;
  assign n1801 = ~n1797 & n1800;
  assign n1802 = n1795 & n1801;
  assign n1803 = ~n1795 & ~n1801;
  assign n1804 = ~n1802 & ~n1803;
  assign n1805 = ~n1785 & ~n1792;
  assign n1806 = ~n1793 & ~n1805;
  assign n1807 = n1804 & n1806;
  assign n1808 = ~n1793 & ~n1807;
  assign n1809 = ~n1641 & n1802;
  assign n1810 = n1641 & ~n1802;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = ~n1808 & ~n1811;
  assign n1813 = n1641 & n1802;
  assign n1814 = ~n1812 & ~n1813;
  assign n1815 = n1804 & ~n1806;
  assign n1816 = ~n1804 & n1806;
  assign n1817 = ~n1815 & ~n1816;
  assign n1818 = ~n984 & ~n1328;
  assign n1819 = ~n979 & n1818;
  assign n1820 = ~n57 & n1328;
  assign n1821 = n979 & ~n1818;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = ~n1819 & n1822;
  assign n1824 = ~n1154 & ~n1289;
  assign n1825 = n1152 & ~n1824;
  assign n1826 = n1823 & n1825;
  assign n1827 = ~n63 & ~n1328;
  assign n1828 = ~n979 & n1827;
  assign n1829 = ~n984 & n1328;
  assign n1830 = n979 & ~n1827;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = ~n1828 & n1831;
  assign n1833 = ~n1200 & n1205;
  assign n1834 = n1200 & n1207;
  assign n1835 = ~n57 & n1209;
  assign n1836 = n57 & n1211;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = ~n1834 & n1837;
  assign n1839 = ~n1833 & n1838;
  assign n1840 = n1832 & ~n1839;
  assign n1841 = ~n1832 & n1839;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = n1826 & ~n1842;
  assign n1844 = n1832 & n1839;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = n1817 & n1845;
  assign n1847 = ~n1817 & ~n1845;
  assign n1848 = ~n1823 & ~n1825;
  assign n1849 = ~n1826 & ~n1848;
  assign n1850 = ~n1200 & ~n1328;
  assign n1851 = ~n979 & n1289;
  assign n1852 = ~n1850 & n1851;
  assign n1853 = ~n57 & ~n1328;
  assign n1854 = ~n979 & n1853;
  assign n1855 = ~n1200 & n1328;
  assign n1856 = n979 & ~n1853;
  assign n1857 = ~n1855 & ~n1856;
  assign n1858 = ~n1854 & n1857;
  assign n1859 = n1824 & n1858;
  assign n1860 = ~n1852 & ~n1859;
  assign n1861 = ~n1824 & ~n1858;
  assign n1862 = ~n1860 & ~n1861;
  assign n1863 = ~n1849 & ~n1862;
  assign n1864 = n1849 & n1862;
  assign n1865 = n1207 & n1289;
  assign n1866 = ~n1200 & n1209;
  assign n1867 = n1200 & n1211;
  assign n1868 = n1205 & ~n1289;
  assign n1869 = ~n1867 & ~n1868;
  assign n1870 = ~n1866 & n1869;
  assign n1871 = ~n1865 & n1870;
  assign n1872 = ~n1864 & ~n1871;
  assign n1873 = ~n1863 & ~n1872;
  assign n1874 = ~n1826 & n1842;
  assign n1875 = ~n1843 & ~n1874;
  assign n1876 = n1794 & n1875;
  assign n1877 = ~n1873 & ~n1876;
  assign n1878 = ~n1794 & ~n1875;
  assign n1879 = ~n1877 & ~n1878;
  assign n1880 = ~n1847 & ~n1879;
  assign n1881 = ~n1846 & ~n1880;
  assign n1882 = n1808 & n1811;
  assign n1883 = ~n1812 & ~n1882;
  assign n1884 = n1760 & ~n1767;
  assign n1885 = ~n1768 & ~n1884;
  assign n1886 = n1883 & n1885;
  assign n1887 = ~n1881 & ~n1886;
  assign n1888 = ~n1883 & ~n1885;
  assign n1889 = ~n1887 & ~n1888;
  assign n1890 = ~n1814 & n1889;
  assign n1891 = n1814 & ~n1889;
  assign n1892 = n1774 & ~n1776;
  assign n1893 = ~n1777 & ~n1892;
  assign n1894 = ~n1891 & n1893;
  assign n1895 = ~n1890 & ~n1894;
  assign n1896 = ~n1778 & ~n1895;
  assign n1897 = n1778 & n1895;
  assign n1898 = ~n1738 & ~n1740;
  assign n1899 = ~n1741 & ~n1898;
  assign n1900 = ~n1897 & n1899;
  assign n1901 = ~n1896 & ~n1900;
  assign n1902 = n1742 & n1901;
  assign n1903 = n1706 & ~n1902;
  assign n1904 = ~n1742 & ~n1901;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = ~n1704 & ~n1905;
  assign n1907 = n1704 & n1905;
  assign n1908 = ~n1617 & ~n1619;
  assign n1909 = ~n1620 & ~n1908;
  assign n1910 = n1689 & n1696;
  assign n1911 = ~n1700 & ~n1910;
  assign n1912 = n1552 & n1559;
  assign n1913 = ~n1552 & ~n1559;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = ~n1911 & ~n1914;
  assign n1916 = n1911 & n1914;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = n1909 & n1917;
  assign n1919 = ~n1909 & ~n1917;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = ~n1907 & n1920;
  assign n1922 = ~n1906 & ~n1921;
  assign n1923 = ~n1915 & ~n1918;
  assign n1924 = ~n1587 & ~n1627;
  assign n1925 = ~n1628 & ~n1924;
  assign n1926 = ~n1923 & n1925;
  assign n1927 = n1922 & ~n1926;
  assign n1928 = n1923 & ~n1925;
  assign n1929 = ~n1927 & ~n1928;
  assign n1930 = n1634 & n1929;
  assign n1931 = ~n1632 & ~n1930;
  assign n1932 = n1582 & ~n1584;
  assign n1933 = ~n1585 & ~n1932;
  assign n1934 = ~n1931 & n1933;
  assign n1935 = ~n1585 & ~n1934;
  assign n1936 = n1504 & ~n1506;
  assign n1937 = ~n1507 & ~n1936;
  assign n1938 = ~n1935 & n1937;
  assign n1939 = ~n1507 & ~n1938;
  assign n1940 = n1462 & ~n1464;
  assign n1941 = ~n1465 & ~n1940;
  assign n1942 = ~n1939 & n1941;
  assign n1943 = ~n1465 & ~n1942;
  assign n1944 = n1276 & n1393;
  assign n1945 = ~n1394 & ~n1944;
  assign n1946 = ~n1943 & n1945;
  assign n1947 = ~n1394 & ~n1946;
  assign n1948 = n1268 & n1272;
  assign n1949 = ~n1273 & ~n1948;
  assign n1950 = ~n1947 & n1949;
  assign n1951 = ~n1273 & ~n1950;
  assign n1952 = ~n1083 & ~n1133;
  assign n1953 = ~n1134 & ~n1952;
  assign n1954 = ~n1951 & n1953;
  assign n1955 = ~n1134 & ~n1954;
  assign n1956 = n1078 & ~n1080;
  assign n1957 = ~n1081 & ~n1956;
  assign n1958 = ~n1955 & n1957;
  assign n1959 = ~n1081 & ~n1958;
  assign n1960 = n886 & n912;
  assign n1961 = ~n913 & ~n1960;
  assign n1962 = ~n1959 & n1961;
  assign n1963 = ~n913 & ~n1962;
  assign n1964 = ~n887 & ~n888;
  assign n1965 = ~n891 & n909;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = ~n896 & ~n907;
  assign n1968 = n600 & ~n609;
  assign n1969 = n594 & n609;
  assign n1970 = ~n741 & n1091;
  assign n1971 = n596 & n741;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~n1969 & n1972;
  assign n1974 = ~n1968 & n1973;
  assign n1975 = ~n1967 & n1974;
  assign n1976 = n1967 & ~n1974;
  assign n1977 = ~n1975 & ~n1976;
  assign n1978 = n586 & ~n803;
  assign n1979 = ~n586 & n803;
  assign n1980 = ~n1978 & ~n1979;
  assign n1981 = n871 & n1980;
  assign n1982 = ~n871 & ~n1980;
  assign n1983 = ~n1981 & ~n1982;
  assign n1984 = n1977 & n1983;
  assign n1985 = ~n1977 & ~n1983;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = ~n1966 & n1986;
  assign n1988 = n1966 & ~n1986;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = ~n1963 & n1989;
  assign n1991 = n1963 & ~n1989;
  assign n1992 = ~n1990 & ~n1991;
  assign n1993 = n334 & n659;
  assign n1994 = n380 & n1993;
  assign n1995 = n786 & n1994;
  assign n1996 = ~n515 & n1995;
  assign n1997 = n309 & n954;
  assign n1998 = ~n262 & n1997;
  assign n1999 = n1996 & n1998;
  assign n2000 = n372 & n771;
  assign n2001 = ~n524 & n2000;
  assign n2002 = ~n469 & n488;
  assign n2003 = ~n397 & n2002;
  assign n2004 = n2001 & n2003;
  assign n2005 = n1999 & n2004;
  assign n2006 = ~n1992 & ~n2005;
  assign n2007 = n1959 & ~n1961;
  assign n2008 = ~n1962 & ~n2007;
  assign n2009 = ~n248 & ~n327;
  assign n2010 = ~n415 & n2009;
  assign n2011 = n340 & ~n367;
  assign n2012 = ~n332 & n2011;
  assign n2013 = n2010 & n2012;
  assign n2014 = ~n194 & n2013;
  assign n2015 = ~n174 & n2014;
  assign n2016 = n694 & n782;
  assign n2017 = n486 & n2016;
  assign n2018 = n2015 & n2017;
  assign n2019 = ~n172 & ~n477;
  assign n2020 = ~n263 & n2019;
  assign n2021 = n717 & n2020;
  assign n2022 = n2018 & n2021;
  assign n2023 = ~n226 & n569;
  assign n2024 = ~n119 & n2023;
  assign n2025 = n2022 & n2024;
  assign n2026 = n699 & n2025;
  assign n2027 = ~n214 & ~n258;
  assign n2028 = ~n197 & n2027;
  assign n2029 = ~n201 & n2028;
  assign n2030 = ~n476 & n2029;
  assign n2031 = ~n265 & ~n282;
  assign n2032 = n619 & n2031;
  assign n2033 = n786 & n2032;
  assign n2034 = ~n132 & n2033;
  assign n2035 = ~n186 & ~n378;
  assign n2036 = ~n159 & n2035;
  assign n2037 = ~n333 & n390;
  assign n2038 = ~n548 & n2037;
  assign n2039 = n2036 & n2038;
  assign n2040 = ~n166 & n2039;
  assign n2041 = n2034 & n2040;
  assign n2042 = n707 & n2041;
  assign n2043 = n2030 & n2042;
  assign n2044 = ~n133 & ~n326;
  assign n2045 = ~n254 & n2044;
  assign n2046 = n761 & n2045;
  assign n2047 = ~n670 & n2046;
  assign n2048 = n2043 & n2047;
  assign n2049 = n2026 & n2048;
  assign n2050 = ~n2008 & ~n2049;
  assign n2051 = n1955 & ~n1957;
  assign n2052 = ~n1958 & ~n2051;
  assign n2053 = n143 & ~n295;
  assign n2054 = ~n149 & n531;
  assign n2055 = ~n762 & n2054;
  assign n2056 = n2053 & n2055;
  assign n2057 = ~n270 & n2056;
  assign n2058 = ~n199 & n2020;
  assign n2059 = ~n360 & n2058;
  assign n2060 = ~n183 & n2059;
  assign n2061 = n2057 & n2060;
  assign n2062 = ~n539 & n2061;
  assign n2063 = ~n365 & n2062;
  assign n2064 = ~n147 & n2063;
  assign n2065 = ~n281 & ~n524;
  assign n2066 = n646 & n2065;
  assign n2067 = ~n361 & n2066;
  assign n2068 = ~n150 & ~n217;
  assign n2069 = ~n248 & n2068;
  assign n2070 = n2067 & n2069;
  assign n2071 = n1310 & n2070;
  assign n2072 = ~n133 & n2071;
  assign n2073 = ~n337 & n2043;
  assign n2074 = ~n206 & n2073;
  assign n2075 = ~n450 & n2074;
  assign n2076 = n244 & n2075;
  assign n2077 = n422 & n2076;
  assign n2078 = ~n213 & n2077;
  assign n2079 = n2072 & n2078;
  assign n2080 = ~n262 & ~n336;
  assign n2081 = ~n367 & n2080;
  assign n2082 = n2079 & n2081;
  assign n2083 = n2064 & n2082;
  assign n2084 = ~n2052 & ~n2083;
  assign n2085 = n1951 & ~n1953;
  assign n2086 = ~n1954 & ~n2085;
  assign n2087 = ~n174 & ~n361;
  assign n2088 = ~n232 & ~n274;
  assign n2089 = n2087 & n2088;
  assign n2090 = ~n265 & n2089;
  assign n2091 = ~n219 & ~n414;
  assign n2092 = ~n397 & n2091;
  assign n2093 = n2090 & n2092;
  assign n2094 = ~n159 & n2093;
  assign n2095 = ~n254 & n2094;
  assign n2096 = ~n386 & ~n532;
  assign n2097 = ~n449 & ~n470;
  assign n2098 = ~n139 & n2097;
  assign n2099 = n2096 & n2098;
  assign n2100 = ~n163 & n2099;
  assign n2101 = ~n445 & n2100;
  assign n2102 = n2095 & n2101;
  assign n2103 = n530 & n2102;
  assign n2104 = n345 & ~n635;
  assign n2105 = ~n468 & n2104;
  assign n2106 = ~n204 & ~n389;
  assign n2107 = n151 & ~n367;
  assign n2108 = ~n140 & n2107;
  assign n2109 = n2106 & n2108;
  assign n2110 = ~n524 & n969;
  assign n2111 = ~n256 & n761;
  assign n2112 = n2110 & n2111;
  assign n2113 = n355 & n2112;
  assign n2114 = n2109 & n2113;
  assign n2115 = ~n221 & n2114;
  assign n2116 = ~n197 & n2115;
  assign n2117 = n2105 & n2116;
  assign n2118 = n2103 & n2117;
  assign n2119 = ~n2086 & ~n2118;
  assign n2120 = n1947 & ~n1949;
  assign n2121 = ~n1950 & ~n2120;
  assign n2122 = ~n332 & ~n381;
  assign n2123 = ~n468 & n2122;
  assign n2124 = n164 & n2123;
  assign n2125 = n763 & n2124;
  assign n2126 = n134 & n2125;
  assign n2127 = ~n206 & n2126;
  assign n2128 = n276 & n427;
  assign n2129 = ~n470 & n2128;
  assign n2130 = n2127 & n2129;
  assign n2131 = n971 & n2130;
  assign n2132 = ~n351 & n550;
  assign n2133 = ~n535 & n2132;
  assign n2134 = ~n317 & n2133;
  assign n2135 = ~n219 & ~n532;
  assign n2136 = n245 & n328;
  assign n2137 = ~n366 & n452;
  assign n2138 = ~n635 & n2137;
  assign n2139 = n692 & n2138;
  assign n2140 = n2136 & n2139;
  assign n2141 = n2135 & n2140;
  assign n2142 = ~n302 & n2141;
  assign n2143 = n2134 & n2142;
  assign n2144 = n2131 & n2143;
  assign n2145 = ~n2121 & ~n2144;
  assign n2146 = n1943 & ~n1945;
  assign n2147 = ~n1946 & ~n2146;
  assign n2148 = ~n283 & n447;
  assign n2149 = ~n440 & n2148;
  assign n2150 = ~n114 & n2149;
  assign n2151 = ~n171 & ~n282;
  assign n2152 = n151 & ~n194;
  assign n2153 = ~n133 & ~n281;
  assign n2154 = n2152 & n2153;
  assign n2155 = ~n541 & n2154;
  assign n2156 = n2151 & n2155;
  assign n2157 = ~n532 & n707;
  assign n2158 = ~n169 & n2157;
  assign n2159 = ~n142 & n765;
  assign n2160 = ~n255 & ~n270;
  assign n2161 = n2106 & n2160;
  assign n2162 = ~n407 & n2161;
  assign n2163 = n2159 & n2162;
  assign n2164 = n1029 & n2163;
  assign n2165 = n2158 & n2164;
  assign n2166 = n717 & n2165;
  assign n2167 = ~n320 & n2166;
  assign n2168 = n2156 & n2167;
  assign n2169 = ~n256 & n2168;
  assign n2170 = ~n163 & ~n262;
  assign n2171 = ~n381 & n2170;
  assign n2172 = ~n287 & n2171;
  assign n2173 = ~n199 & n2172;
  assign n2174 = ~n130 & n2035;
  assign n2175 = ~n408 & ~n670;
  assign n2176 = ~n249 & n2175;
  assign n2177 = n2174 & n2176;
  assign n2178 = n343 & n2177;
  assign n2179 = n2173 & n2178;
  assign n2180 = ~n166 & n2179;
  assign n2181 = ~n147 & n2180;
  assign n2182 = n2169 & n2181;
  assign n2183 = ~n132 & n2182;
  assign n2184 = n2150 & n2183;
  assign n2185 = ~n2147 & ~n2184;
  assign n2186 = n1939 & ~n1941;
  assign n2187 = ~n1942 & ~n2186;
  assign n2188 = n523 & ~n541;
  assign n2189 = ~n270 & ~n445;
  assign n2190 = n188 & n2189;
  assign n2191 = ~n294 & n2190;
  assign n2192 = n2188 & n2191;
  assign n2193 = n712 & n2192;
  assign n2194 = ~n197 & n2193;
  assign n2195 = ~n670 & n2194;
  assign n2196 = ~n635 & n687;
  assign n2197 = ~n304 & n2196;
  assign n2198 = n340 & ~n407;
  assign n2199 = ~n365 & n2045;
  assign n2200 = n2198 & n2199;
  assign n2201 = n224 & n2200;
  assign n2202 = n2197 & n2201;
  assign n2203 = n411 & n2202;
  assign n2204 = n490 & n2203;
  assign n2205 = ~n265 & n2204;
  assign n2206 = ~n337 & n2205;
  assign n2207 = n2195 & n2206;
  assign n2208 = ~n139 & n2207;
  assign n2209 = ~n226 & n618;
  assign n2210 = ~n346 & n2209;
  assign n2211 = ~n173 & n2210;
  assign n2212 = n2208 & n2211;
  assign n2213 = ~n2187 & ~n2212;
  assign n2214 = n1935 & ~n1937;
  assign n2215 = ~n1938 & ~n2214;
  assign n2216 = ~n297 & ~n325;
  assign n2217 = n244 & n312;
  assign n2218 = n611 & n2217;
  assign n2219 = n2216 & n2218;
  assign n2220 = ~n228 & n2219;
  assign n2221 = n424 & n722;
  assign n2222 = ~n332 & n2221;
  assign n2223 = n2220 & n2222;
  assign n2224 = n765 & n2081;
  assign n2225 = ~n407 & n2224;
  assign n2226 = ~n337 & ~n408;
  assign n2227 = n261 & n2226;
  assign n2228 = ~n440 & n2227;
  assign n2229 = n2225 & n2228;
  assign n2230 = n387 & n2229;
  assign n2231 = ~n281 & ~n762;
  assign n2232 = ~n295 & ~n327;
  assign n2233 = ~n568 & n2232;
  assign n2234 = n2231 & n2233;
  assign n2235 = ~n360 & n2234;
  assign n2236 = ~n515 & n2235;
  assign n2237 = n2134 & n2236;
  assign n2238 = n2230 & n2237;
  assign n2239 = ~n159 & n2238;
  assign n2240 = ~n185 & n2239;
  assign n2241 = n143 & n2192;
  assign n2242 = ~n365 & n2241;
  assign n2243 = n2240 & n2242;
  assign n2244 = n2223 & n2243;
  assign n2245 = ~n2215 & ~n2244;
  assign n2246 = n1931 & ~n1933;
  assign n2247 = ~n1934 & ~n2246;
  assign n2248 = n416 & n2140;
  assign n2249 = ~n348 & n2248;
  assign n2250 = ~n254 & n2249;
  assign n2251 = n380 & n2226;
  assign n2252 = ~n541 & n2251;
  assign n2253 = ~n140 & n2252;
  assign n2254 = n2250 & n2253;
  assign n2255 = ~n214 & n613;
  assign n2256 = ~n232 & n2255;
  assign n2257 = ~n213 & ~n548;
  assign n2258 = ~n171 & ~n446;
  assign n2259 = ~n255 & n2258;
  assign n2260 = n2257 & n2259;
  assign n2261 = ~n360 & ~n539;
  assign n2262 = n2260 & n2261;
  assign n2263 = ~n316 & n2262;
  assign n2264 = n112 & n141;
  assign n2265 = ~n670 & n958;
  assign n2266 = ~n256 & n2265;
  assign n2267 = ~n2264 & n2266;
  assign n2268 = ~n524 & n2267;
  assign n2269 = ~n336 & n2268;
  assign n2270 = n2263 & n2269;
  assign n2271 = ~n361 & n2270;
  assign n2272 = ~n123 & n2271;
  assign n2273 = n2256 & n2272;
  assign n2274 = n2254 & n2273;
  assign n2275 = ~n2247 & ~n2274;
  assign n2276 = ~n1634 & ~n1929;
  assign n2277 = ~n1930 & ~n2276;
  assign n2278 = ~n187 & n780;
  assign n2279 = ~n379 & n2278;
  assign n2280 = ~n469 & n2279;
  assign n2281 = ~n316 & n2280;
  assign n2282 = n671 & n2038;
  assign n2283 = n472 & n2282;
  assign n2284 = n447 & n941;
  assign n2285 = n2283 & n2284;
  assign n2286 = n411 & n2285;
  assign n2287 = n2281 & n2286;
  assign n2288 = n765 & n2287;
  assign n2289 = ~n515 & n2288;
  assign n2290 = n323 & n500;
  assign n2291 = ~n762 & n2290;
  assign n2292 = n2289 & n2291;
  assign n2293 = ~n194 & n2202;
  assign n2294 = ~n284 & n2293;
  assign n2295 = n488 & n944;
  assign n2296 = ~n348 & n2295;
  assign n2297 = n2294 & n2296;
  assign n2298 = n2292 & n2297;
  assign n2299 = n2277 & n2298;
  assign n2300 = n2247 & n2274;
  assign n2301 = ~n2275 & ~n2300;
  assign n2302 = ~n2299 & n2301;
  assign n2303 = ~n2275 & ~n2302;
  assign n2304 = n2215 & n2244;
  assign n2305 = ~n2245 & ~n2304;
  assign n2306 = ~n2303 & n2305;
  assign n2307 = ~n2245 & ~n2306;
  assign n2308 = n2187 & n2212;
  assign n2309 = ~n2213 & ~n2308;
  assign n2310 = ~n2307 & n2309;
  assign n2311 = ~n2213 & ~n2310;
  assign n2312 = n2147 & n2184;
  assign n2313 = ~n2185 & ~n2312;
  assign n2314 = ~n2311 & n2313;
  assign n2315 = ~n2185 & ~n2314;
  assign n2316 = n2121 & n2144;
  assign n2317 = ~n2145 & ~n2316;
  assign n2318 = ~n2315 & n2317;
  assign n2319 = ~n2145 & ~n2318;
  assign n2320 = n2086 & n2118;
  assign n2321 = ~n2119 & ~n2320;
  assign n2322 = ~n2319 & n2321;
  assign n2323 = ~n2119 & ~n2322;
  assign n2324 = n2052 & n2083;
  assign n2325 = ~n2084 & ~n2324;
  assign n2326 = ~n2323 & n2325;
  assign n2327 = ~n2084 & ~n2326;
  assign n2328 = n2008 & n2049;
  assign n2329 = ~n2050 & ~n2328;
  assign n2330 = ~n2327 & n2329;
  assign n2331 = ~n2050 & ~n2330;
  assign n2332 = n1992 & n2005;
  assign n2333 = ~n2006 & ~n2332;
  assign n2334 = ~n2331 & n2333;
  assign n2335 = ~n2006 & ~n2334;
  assign n2336 = ~n1987 & ~n1990;
  assign n2337 = ~n1975 & ~n1984;
  assign n2338 = ~n1978 & ~n1981;
  assign n2339 = n581 & ~n741;
  assign n2340 = ~n593 & ~n2339;
  assign n2341 = ~n599 & n2339;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = ~n899 & n2342;
  assign n2344 = n899 & ~n2342;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = ~n2338 & n2345;
  assign n2347 = n2338 & ~n2345;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = ~n2337 & n2348;
  assign n2350 = n2337 & ~n2348;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = ~n2336 & n2351;
  assign n2353 = n2336 & ~n2351;
  assign n2354 = ~n2352 & ~n2353;
  assign n2355 = n207 & n495;
  assign n2356 = n131 & n2355;
  assign n2357 = ~n325 & n2356;
  assign n2358 = ~n346 & ~n415;
  assign n2359 = ~n378 & ~n635;
  assign n2360 = ~n515 & n2359;
  assign n2361 = n2358 & n2360;
  assign n2362 = ~n284 & n2361;
  assign n2363 = ~n195 & ~n351;
  assign n2364 = n2362 & n2363;
  assign n2365 = ~n147 & n2364;
  assign n2366 = n441 & ~n476;
  assign n2367 = ~n271 & n2366;
  assign n2368 = ~n173 & n2367;
  assign n2369 = n2365 & n2368;
  assign n2370 = n610 & n2369;
  assign n2371 = ~n159 & n2370;
  assign n2372 = n2357 & n2371;
  assign n2373 = n2070 & n2372;
  assign n2374 = ~n139 & n2287;
  assign n2375 = ~n270 & n2374;
  assign n2376 = n2028 & n2375;
  assign n2377 = n451 & n2376;
  assign n2378 = n2373 & n2377;
  assign n2379 = ~n2354 & ~n2378;
  assign n2380 = n2354 & n2378;
  assign n2381 = ~n2379 & ~n2380;
  assign n2382 = ~n2335 & n2381;
  assign n2383 = n2335 & ~n2381;
  assign n2384 = ~n2382 & ~n2383;
  assign n2385 = n57 & n1200;
  assign n2386 = ~n57 & ~n1200;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = pi2  & pi22 ;
  assign n2389 = ~pi0  & ~pi1 ;
  assign n2390 = pi2  & ~n2389;
  assign n2391 = n1286 & ~n2390;
  assign n2392 = ~n2388 & ~n2391;
  assign n2393 = n1289 & n2392;
  assign n2394 = ~n1289 & ~n2392;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = n1200 & n1289;
  assign n2397 = ~n1200 & ~n1289;
  assign n2398 = ~n2396 & ~n2397;
  assign n2399 = ~n2395 & ~n2398;
  assign n2400 = n2387 & n2399;
  assign n2401 = n2384 & n2400;
  assign n2402 = ~n2395 & n2398;
  assign n2403 = ~n2379 & ~n2382;
  assign n2404 = ~n228 & ~n293;
  assign n2405 = n526 & n2404;
  assign n2406 = n763 & n2405;
  assign n2407 = n966 & n2406;
  assign n2408 = ~n205 & ~n317;
  assign n2409 = ~n397 & ~n635;
  assign n2410 = ~n130 & n2409;
  assign n2411 = n2036 & n2410;
  assign n2412 = n2408 & n2411;
  assign n2413 = n244 & n2412;
  assign n2414 = ~n214 & n2413;
  assign n2415 = n2407 & n2414;
  assign n2416 = ~n123 & n2415;
  assign n2417 = ~n226 & n404;
  assign n2418 = ~n199 & n2417;
  assign n2419 = ~n295 & n2418;
  assign n2420 = n312 & n2167;
  assign n2421 = n2419 & n2420;
  assign n2422 = n2416 & n2421;
  assign n2423 = n609 & n741;
  assign n2424 = ~n609 & ~n741;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = n592 & ~n2425;
  assign n2427 = ~n592 & n2425;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = ~n238 & n2428;
  assign n2430 = ~n2349 & ~n2352;
  assign n2431 = ~n2343 & ~n2346;
  assign n2432 = n2430 & ~n2431;
  assign n2433 = ~n2430 & n2431;
  assign n2434 = ~n2432 & ~n2433;
  assign n2435 = n2429 & n2434;
  assign n2436 = ~n2429 & ~n2434;
  assign n2437 = ~n2435 & ~n2436;
  assign n2438 = ~n2422 & ~n2437;
  assign n2439 = n2422 & n2437;
  assign n2440 = ~n2438 & ~n2439;
  assign n2441 = ~n2403 & n2440;
  assign n2442 = n2403 & ~n2440;
  assign n2443 = ~n2441 & ~n2442;
  assign n2444 = n2402 & n2443;
  assign n2445 = n2387 & n2395;
  assign n2446 = n2384 & n2443;
  assign n2447 = n2331 & ~n2333;
  assign n2448 = ~n2334 & ~n2447;
  assign n2449 = n2384 & n2448;
  assign n2450 = n2327 & ~n2329;
  assign n2451 = ~n2330 & ~n2450;
  assign n2452 = n2448 & n2451;
  assign n2453 = n2323 & ~n2325;
  assign n2454 = ~n2326 & ~n2453;
  assign n2455 = n2451 & n2454;
  assign n2456 = n2319 & ~n2321;
  assign n2457 = ~n2322 & ~n2456;
  assign n2458 = n2454 & n2457;
  assign n2459 = n2315 & ~n2317;
  assign n2460 = ~n2318 & ~n2459;
  assign n2461 = n2457 & n2460;
  assign n2462 = n2311 & ~n2313;
  assign n2463 = ~n2314 & ~n2462;
  assign n2464 = n2460 & n2463;
  assign n2465 = n2307 & ~n2309;
  assign n2466 = ~n2310 & ~n2465;
  assign n2467 = n2463 & n2466;
  assign n2468 = n2303 & ~n2305;
  assign n2469 = ~n2306 & ~n2468;
  assign n2470 = n2466 & n2469;
  assign n2471 = ~n2277 & ~n2298;
  assign n2472 = ~n2299 & ~n2471;
  assign n2473 = ~n2469 & n2472;
  assign n2474 = n2299 & ~n2301;
  assign n2475 = ~n2302 & ~n2474;
  assign n2476 = ~n2473 & n2475;
  assign n2477 = ~n2466 & ~n2469;
  assign n2478 = ~n2470 & ~n2477;
  assign n2479 = n2476 & n2478;
  assign n2480 = ~n2470 & ~n2479;
  assign n2481 = ~n2463 & ~n2466;
  assign n2482 = ~n2467 & ~n2481;
  assign n2483 = ~n2480 & n2482;
  assign n2484 = ~n2467 & ~n2483;
  assign n2485 = ~n2460 & ~n2463;
  assign n2486 = ~n2464 & ~n2485;
  assign n2487 = ~n2484 & n2486;
  assign n2488 = ~n2464 & ~n2487;
  assign n2489 = ~n2457 & ~n2460;
  assign n2490 = ~n2461 & ~n2489;
  assign n2491 = ~n2488 & n2490;
  assign n2492 = ~n2461 & ~n2491;
  assign n2493 = ~n2454 & ~n2457;
  assign n2494 = ~n2458 & ~n2493;
  assign n2495 = ~n2492 & n2494;
  assign n2496 = ~n2458 & ~n2495;
  assign n2497 = ~n2451 & ~n2454;
  assign n2498 = ~n2455 & ~n2497;
  assign n2499 = ~n2496 & n2498;
  assign n2500 = ~n2455 & ~n2499;
  assign n2501 = ~n2448 & ~n2451;
  assign n2502 = ~n2452 & ~n2501;
  assign n2503 = ~n2500 & n2502;
  assign n2504 = ~n2452 & ~n2503;
  assign n2505 = ~n2384 & ~n2448;
  assign n2506 = ~n2449 & ~n2505;
  assign n2507 = ~n2504 & n2506;
  assign n2508 = ~n2449 & ~n2507;
  assign n2509 = ~n2384 & ~n2443;
  assign n2510 = ~n2446 & ~n2509;
  assign n2511 = ~n2508 & n2510;
  assign n2512 = ~n2446 & ~n2511;
  assign n2513 = ~n2438 & ~n2441;
  assign n2514 = ~n217 & n617;
  assign n2515 = ~n407 & n2514;
  assign n2516 = n569 & n2140;
  assign n2517 = n941 & n2516;
  assign n2518 = ~n670 & n2517;
  assign n2519 = ~n174 & ~n221;
  assign n2520 = ~n389 & n2519;
  assign n2521 = ~n142 & ~n199;
  assign n2522 = n651 & n2521;
  assign n2523 = n2520 & n2522;
  assign n2524 = n1316 & n2523;
  assign n2525 = n753 & n2524;
  assign n2526 = ~n336 & n2525;
  assign n2527 = n2518 & n2526;
  assign n2528 = n285 & n2527;
  assign n2529 = n2515 & n2528;
  assign n2530 = n2513 & n2529;
  assign n2531 = ~n2513 & ~n2529;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = n2443 & ~n2532;
  assign n2534 = ~n2443 & n2532;
  assign n2535 = ~n2533 & ~n2534;
  assign n2536 = ~n2512 & n2535;
  assign n2537 = n2512 & ~n2535;
  assign n2538 = ~n2536 & ~n2537;
  assign n2539 = n2445 & n2538;
  assign n2540 = ~n2387 & n2395;
  assign n2541 = ~n2532 & n2540;
  assign n2542 = ~n2539 & ~n2541;
  assign n2543 = ~n2444 & n2542;
  assign n2544 = ~n2401 & n2543;
  assign n2545 = ~n57 & ~n2544;
  assign n2546 = n57 & n2544;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = n509 & n824;
  assign n2549 = ~n509 & ~n824;
  assign n2550 = ~n2548 & ~n2549;
  assign n2551 = n591 & n824;
  assign n2552 = ~n591 & ~n824;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = ~n2550 & n2553;
  assign n2555 = n2466 & n2554;
  assign n2556 = n585 & n591;
  assign n2557 = ~n585 & ~n591;
  assign n2558 = ~n2556 & ~n2557;
  assign n2559 = n2550 & ~n2558;
  assign n2560 = n2463 & n2559;
  assign n2561 = n2550 & n2558;
  assign n2562 = n2480 & ~n2482;
  assign n2563 = ~n2483 & ~n2562;
  assign n2564 = n2561 & n2563;
  assign n2565 = ~n2550 & n2558;
  assign n2566 = ~n2553 & n2565;
  assign n2567 = n2469 & n2566;
  assign n2568 = ~n2564 & ~n2567;
  assign n2569 = ~n2560 & n2568;
  assign n2570 = ~n2555 & n2569;
  assign n2571 = n585 & n2570;
  assign n2572 = ~n585 & ~n2570;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = ~n2472 & ~n2475;
  assign n2575 = ~n2301 & n2472;
  assign n2576 = ~n2574 & ~n2575;
  assign n2577 = n585 & n810;
  assign n2578 = ~n585 & ~n810;
  assign n2579 = ~n2577 & ~n2578;
  assign n2580 = n2425 & n2579;
  assign n2581 = ~n2576 & n2580;
  assign n2582 = ~n2425 & n2579;
  assign n2583 = n2475 & n2582;
  assign n2584 = n609 & n810;
  assign n2585 = ~n609 & ~n810;
  assign n2586 = ~n2584 & ~n2585;
  assign n2587 = ~n2579 & n2586;
  assign n2588 = ~n2472 & n2587;
  assign n2589 = ~n2583 & ~n2588;
  assign n2590 = ~n2581 & n2589;
  assign n2591 = ~n741 & ~n2472;
  assign n2592 = n2579 & n2591;
  assign n2593 = ~n2590 & n2592;
  assign n2594 = n2590 & ~n2592;
  assign n2595 = ~n2593 & ~n2594;
  assign n2596 = n2573 & n2595;
  assign n2597 = ~n2472 & n2579;
  assign n2598 = ~n2472 & n2550;
  assign n2599 = ~n585 & ~n2598;
  assign n2600 = n2561 & ~n2576;
  assign n2601 = n2475 & n2559;
  assign n2602 = ~n2472 & n2554;
  assign n2603 = ~n2601 & ~n2602;
  assign n2604 = ~n2600 & n2603;
  assign n2605 = n2599 & n2604;
  assign n2606 = ~n2472 & n2566;
  assign n2607 = n2475 & n2554;
  assign n2608 = n2469 & ~n2575;
  assign n2609 = ~n2469 & n2575;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = n2561 & ~n2610;
  assign n2612 = n2469 & n2559;
  assign n2613 = ~n2611 & ~n2612;
  assign n2614 = ~n2607 & n2613;
  assign n2615 = ~n2606 & n2614;
  assign n2616 = n2605 & n2615;
  assign n2617 = n2597 & n2616;
  assign n2618 = ~n2597 & n2616;
  assign n2619 = n2597 & ~n2616;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = n2466 & n2559;
  assign n2622 = n2475 & n2566;
  assign n2623 = ~n2476 & ~n2478;
  assign n2624 = ~n2479 & ~n2623;
  assign n2625 = n2561 & n2624;
  assign n2626 = n2469 & n2554;
  assign n2627 = ~n2625 & ~n2626;
  assign n2628 = ~n2622 & n2627;
  assign n2629 = ~n2621 & n2628;
  assign n2630 = ~n585 & ~n2629;
  assign n2631 = n585 & n2629;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = ~n2620 & n2632;
  assign n2634 = ~n2617 & ~n2633;
  assign n2635 = ~n2573 & ~n2595;
  assign n2636 = ~n2596 & ~n2635;
  assign n2637 = ~n2634 & n2636;
  assign n2638 = ~n2596 & ~n2637;
  assign n2639 = n2466 & n2566;
  assign n2640 = n2463 & n2554;
  assign n2641 = n2484 & ~n2486;
  assign n2642 = ~n2487 & ~n2641;
  assign n2643 = n2561 & n2642;
  assign n2644 = n2460 & n2559;
  assign n2645 = ~n2643 & ~n2644;
  assign n2646 = ~n2640 & n2645;
  assign n2647 = ~n2639 & n2646;
  assign n2648 = ~n585 & ~n2647;
  assign n2649 = n585 & n2647;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = n2425 & ~n2579;
  assign n2652 = ~n2586 & n2651;
  assign n2653 = ~n2472 & n2652;
  assign n2654 = n2475 & n2587;
  assign n2655 = n2580 & ~n2610;
  assign n2656 = n2469 & n2582;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = ~n2654 & n2657;
  assign n2659 = ~n2653 & n2658;
  assign n2660 = n2590 & ~n2597;
  assign n2661 = ~n741 & ~n2660;
  assign n2662 = ~n2659 & n2661;
  assign n2663 = n2659 & ~n2661;
  assign n2664 = ~n2662 & ~n2663;
  assign n2665 = n2650 & n2664;
  assign n2666 = ~n2650 & ~n2664;
  assign n2667 = ~n2665 & ~n2666;
  assign n2668 = n2638 & ~n2667;
  assign n2669 = ~n2638 & n2667;
  assign n2670 = ~n2668 & ~n2669;
  assign n2671 = n63 & n509;
  assign n2672 = ~n63 & ~n509;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = n57 & n984;
  assign n2675 = ~n57 & ~n984;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = n63 & n984;
  assign n2678 = ~n63 & ~n984;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = ~n2676 & ~n2679;
  assign n2681 = n2673 & n2680;
  assign n2682 = n2457 & n2681;
  assign n2683 = ~n2676 & n2679;
  assign n2684 = n2454 & n2683;
  assign n2685 = n2496 & ~n2498;
  assign n2686 = ~n2499 & ~n2685;
  assign n2687 = n2673 & n2676;
  assign n2688 = n2686 & n2687;
  assign n2689 = ~n2673 & n2676;
  assign n2690 = n2451 & n2689;
  assign n2691 = ~n2688 & ~n2690;
  assign n2692 = ~n2684 & n2691;
  assign n2693 = ~n2682 & n2692;
  assign n2694 = n509 & n2693;
  assign n2695 = ~n509 & ~n2693;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = n2670 & n2696;
  assign n2698 = ~n2670 & ~n2696;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = n2460 & n2681;
  assign n2701 = n2457 & n2683;
  assign n2702 = n2492 & ~n2494;
  assign n2703 = ~n2495 & ~n2702;
  assign n2704 = n2687 & n2703;
  assign n2705 = n2454 & n2689;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = ~n2701 & n2706;
  assign n2708 = ~n2700 & n2707;
  assign n2709 = n509 & ~n2708;
  assign n2710 = ~n509 & n2708;
  assign n2711 = ~n2709 & ~n2710;
  assign n2712 = n2634 & ~n2636;
  assign n2713 = ~n2637 & ~n2712;
  assign n2714 = n2711 & ~n2713;
  assign n2715 = ~n2711 & n2713;
  assign n2716 = ~n2620 & ~n2632;
  assign n2717 = n2620 & n2632;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = n2463 & n2681;
  assign n2720 = n2460 & n2683;
  assign n2721 = n2488 & ~n2490;
  assign n2722 = ~n2491 & ~n2721;
  assign n2723 = n2687 & n2722;
  assign n2724 = n2457 & n2689;
  assign n2725 = ~n2723 & ~n2724;
  assign n2726 = ~n2720 & n2725;
  assign n2727 = ~n2719 & n2726;
  assign n2728 = n509 & n2727;
  assign n2729 = ~n509 & ~n2727;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = ~n2718 & n2730;
  assign n2732 = ~n2718 & ~n2730;
  assign n2733 = n2718 & n2730;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = n2466 & n2681;
  assign n2736 = n2463 & n2683;
  assign n2737 = n2642 & n2687;
  assign n2738 = n2460 & n2689;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = ~n2736 & n2739;
  assign n2741 = ~n2735 & n2740;
  assign n2742 = n509 & ~n2741;
  assign n2743 = ~n509 & n2741;
  assign n2744 = ~n2742 & ~n2743;
  assign n2745 = ~n585 & ~n2605;
  assign n2746 = ~n2615 & n2745;
  assign n2747 = n2615 & ~n2745;
  assign n2748 = ~n2746 & ~n2747;
  assign n2749 = n2744 & ~n2748;
  assign n2750 = ~n2744 & n2748;
  assign n2751 = n2466 & n2683;
  assign n2752 = n2463 & n2689;
  assign n2753 = n2563 & n2687;
  assign n2754 = n2469 & n2681;
  assign n2755 = ~n2753 & ~n2754;
  assign n2756 = ~n2752 & n2755;
  assign n2757 = ~n2751 & n2756;
  assign n2758 = n509 & n2757;
  assign n2759 = ~n509 & ~n2757;
  assign n2760 = ~n2758 & ~n2759;
  assign n2761 = ~n585 & n2598;
  assign n2762 = ~n2604 & n2761;
  assign n2763 = n2604 & ~n2761;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = n2760 & n2764;
  assign n2766 = ~n2576 & n2687;
  assign n2767 = n2475 & n2689;
  assign n2768 = ~n2472 & n2683;
  assign n2769 = ~n2767 & ~n2768;
  assign n2770 = ~n2766 & n2769;
  assign n2771 = ~n2472 & n2676;
  assign n2772 = ~n509 & ~n2771;
  assign n2773 = n2770 & n2772;
  assign n2774 = ~n2472 & n2681;
  assign n2775 = n2475 & n2683;
  assign n2776 = ~n2610 & n2687;
  assign n2777 = n2469 & n2689;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = ~n2775 & n2778;
  assign n2780 = ~n2774 & n2779;
  assign n2781 = n2773 & n2780;
  assign n2782 = n2598 & n2781;
  assign n2783 = ~n2598 & n2781;
  assign n2784 = n2598 & ~n2781;
  assign n2785 = ~n2783 & ~n2784;
  assign n2786 = n2466 & n2689;
  assign n2787 = n2475 & n2681;
  assign n2788 = n2624 & n2687;
  assign n2789 = n2469 & n2683;
  assign n2790 = ~n2788 & ~n2789;
  assign n2791 = ~n2787 & n2790;
  assign n2792 = ~n2786 & n2791;
  assign n2793 = ~n509 & n2792;
  assign n2794 = n509 & ~n2792;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = ~n2785 & ~n2795;
  assign n2797 = ~n2782 & ~n2796;
  assign n2798 = ~n2760 & ~n2764;
  assign n2799 = ~n2765 & ~n2798;
  assign n2800 = ~n2797 & n2799;
  assign n2801 = ~n2765 & ~n2800;
  assign n2802 = ~n2750 & n2801;
  assign n2803 = ~n2749 & ~n2802;
  assign n2804 = ~n2734 & n2803;
  assign n2805 = ~n2731 & ~n2804;
  assign n2806 = ~n2715 & n2805;
  assign n2807 = ~n2714 & ~n2806;
  assign n2808 = n2699 & n2807;
  assign n2809 = ~n2697 & ~n2808;
  assign n2810 = ~n2665 & ~n2669;
  assign n2811 = n2463 & n2566;
  assign n2812 = n2460 & n2554;
  assign n2813 = n2561 & n2722;
  assign n2814 = n2457 & n2559;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = ~n2812 & n2815;
  assign n2817 = ~n2811 & n2816;
  assign n2818 = ~n585 & ~n2817;
  assign n2819 = n585 & n2817;
  assign n2820 = ~n2818 & ~n2819;
  assign n2821 = n2466 & n2582;
  assign n2822 = n2475 & n2652;
  assign n2823 = n2580 & n2624;
  assign n2824 = n2469 & n2587;
  assign n2825 = ~n2823 & ~n2824;
  assign n2826 = ~n2822 & n2825;
  assign n2827 = ~n2821 & n2826;
  assign n2828 = n741 & ~n2827;
  assign n2829 = ~n741 & n2827;
  assign n2830 = ~n2828 & ~n2829;
  assign n2831 = ~n741 & n2659;
  assign n2832 = n2660 & n2831;
  assign n2833 = ~n2591 & ~n2832;
  assign n2834 = ~n2472 & n2832;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = n2830 & ~n2835;
  assign n2837 = ~n2830 & n2835;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = n2820 & n2838;
  assign n2840 = ~n2820 & ~n2838;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = n2810 & ~n2841;
  assign n2843 = ~n2810 & n2841;
  assign n2844 = ~n2842 & ~n2843;
  assign n2845 = n2454 & n2681;
  assign n2846 = n2451 & n2683;
  assign n2847 = n2500 & ~n2502;
  assign n2848 = ~n2503 & ~n2847;
  assign n2849 = n2687 & n2848;
  assign n2850 = n2448 & n2689;
  assign n2851 = ~n2849 & ~n2850;
  assign n2852 = ~n2846 & n2851;
  assign n2853 = ~n2845 & n2852;
  assign n2854 = n509 & n2853;
  assign n2855 = ~n509 & ~n2853;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857 = n2844 & n2856;
  assign n2858 = ~n2844 & ~n2856;
  assign n2859 = ~n2857 & ~n2858;
  assign n2860 = ~n2809 & n2859;
  assign n2861 = n2809 & ~n2859;
  assign n2862 = ~n2860 & ~n2861;
  assign n2863 = n2547 & n2862;
  assign n2864 = n2400 & n2448;
  assign n2865 = n2384 & n2402;
  assign n2866 = n2508 & ~n2510;
  assign n2867 = ~n2511 & ~n2866;
  assign n2868 = n2445 & n2867;
  assign n2869 = n2443 & n2540;
  assign n2870 = ~n2868 & ~n2869;
  assign n2871 = ~n2865 & n2870;
  assign n2872 = ~n2864 & n2871;
  assign n2873 = ~n57 & ~n2872;
  assign n2874 = n57 & n2872;
  assign n2875 = ~n2873 & ~n2874;
  assign n2876 = ~n2699 & ~n2807;
  assign n2877 = ~n2808 & ~n2876;
  assign n2878 = n2875 & n2877;
  assign n2879 = n2400 & n2451;
  assign n2880 = n2402 & n2448;
  assign n2881 = n2504 & ~n2506;
  assign n2882 = ~n2507 & ~n2881;
  assign n2883 = n2445 & n2882;
  assign n2884 = n2384 & n2540;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = ~n2880 & n2885;
  assign n2887 = ~n2879 & n2886;
  assign n2888 = n57 & n2887;
  assign n2889 = ~n57 & ~n2887;
  assign n2890 = ~n2888 & ~n2889;
  assign n2891 = ~n2714 & ~n2715;
  assign n2892 = n2805 & n2891;
  assign n2893 = ~n2805 & ~n2891;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = n2890 & ~n2894;
  assign n2896 = n2734 & n2803;
  assign n2897 = ~n2734 & ~n2803;
  assign n2898 = ~n2896 & ~n2897;
  assign n2899 = n2400 & n2454;
  assign n2900 = n2402 & n2451;
  assign n2901 = n2445 & n2848;
  assign n2902 = n2448 & n2540;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = ~n2900 & n2903;
  assign n2905 = ~n2899 & n2904;
  assign n2906 = n57 & n2905;
  assign n2907 = ~n57 & ~n2905;
  assign n2908 = ~n2906 & ~n2907;
  assign n2909 = ~n2898 & n2908;
  assign n2910 = n2400 & n2457;
  assign n2911 = n2402 & n2454;
  assign n2912 = n2445 & n2686;
  assign n2913 = n2451 & n2540;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = ~n2911 & n2914;
  assign n2916 = ~n2910 & n2915;
  assign n2917 = n57 & n2916;
  assign n2918 = ~n57 & ~n2916;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = ~n2749 & ~n2750;
  assign n2921 = n2801 & n2920;
  assign n2922 = ~n2801 & ~n2920;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = n2919 & ~n2923;
  assign n2925 = n2400 & n2460;
  assign n2926 = n2402 & n2457;
  assign n2927 = n2445 & n2703;
  assign n2928 = n2454 & n2540;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = ~n2926 & n2929;
  assign n2931 = ~n2925 & n2930;
  assign n2932 = ~n57 & ~n2931;
  assign n2933 = n57 & n2931;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = n2797 & ~n2799;
  assign n2936 = ~n2800 & ~n2935;
  assign n2937 = n2934 & n2936;
  assign n2938 = n2400 & n2463;
  assign n2939 = n2402 & n2460;
  assign n2940 = n2445 & n2722;
  assign n2941 = n2457 & n2540;
  assign n2942 = ~n2940 & ~n2941;
  assign n2943 = ~n2939 & n2942;
  assign n2944 = ~n2938 & n2943;
  assign n2945 = n57 & n2944;
  assign n2946 = ~n57 & ~n2944;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = n2785 & n2795;
  assign n2949 = ~n2796 & ~n2948;
  assign n2950 = n2947 & n2949;
  assign n2951 = n2400 & n2466;
  assign n2952 = n2402 & n2463;
  assign n2953 = n2445 & n2642;
  assign n2954 = n2460 & n2540;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = ~n2952 & n2955;
  assign n2957 = ~n2951 & n2956;
  assign n2958 = ~n57 & ~n2957;
  assign n2959 = n57 & n2957;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = ~n509 & ~n2773;
  assign n2962 = ~n2780 & n2961;
  assign n2963 = n2780 & ~n2961;
  assign n2964 = ~n2962 & ~n2963;
  assign n2965 = n2960 & n2964;
  assign n2966 = n2402 & n2466;
  assign n2967 = n2463 & n2540;
  assign n2968 = n2445 & n2563;
  assign n2969 = n2400 & n2469;
  assign n2970 = ~n2968 & ~n2969;
  assign n2971 = ~n2967 & n2970;
  assign n2972 = ~n2966 & n2971;
  assign n2973 = n57 & n2972;
  assign n2974 = ~n57 & ~n2972;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = ~n509 & n2771;
  assign n2977 = ~n2770 & n2976;
  assign n2978 = n2770 & ~n2976;
  assign n2979 = ~n2977 & ~n2978;
  assign n2980 = n2975 & n2979;
  assign n2981 = n2395 & ~n2472;
  assign n2982 = ~n57 & ~n2981;
  assign n2983 = n2445 & ~n2576;
  assign n2984 = n2475 & n2540;
  assign n2985 = n2402 & ~n2472;
  assign n2986 = ~n2984 & ~n2985;
  assign n2987 = ~n2983 & n2986;
  assign n2988 = n2982 & n2987;
  assign n2989 = n2400 & ~n2472;
  assign n2990 = n2402 & n2475;
  assign n2991 = n2445 & ~n2610;
  assign n2992 = n2469 & n2540;
  assign n2993 = ~n2991 & ~n2992;
  assign n2994 = ~n2990 & n2993;
  assign n2995 = ~n2989 & n2994;
  assign n2996 = n2988 & n2995;
  assign n2997 = n2771 & n2996;
  assign n2998 = ~n2771 & n2996;
  assign n2999 = n2771 & ~n2996;
  assign n3000 = ~n2998 & ~n2999;
  assign n3001 = n2466 & n2540;
  assign n3002 = n2400 & n2475;
  assign n3003 = n2445 & n2624;
  assign n3004 = n2402 & n2469;
  assign n3005 = ~n3003 & ~n3004;
  assign n3006 = ~n3002 & n3005;
  assign n3007 = ~n3001 & n3006;
  assign n3008 = ~n57 & ~n3007;
  assign n3009 = n57 & n3007;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = ~n3000 & n3010;
  assign n3012 = ~n2997 & ~n3011;
  assign n3013 = ~n2975 & ~n2979;
  assign n3014 = ~n2980 & ~n3013;
  assign n3015 = ~n3012 & n3014;
  assign n3016 = ~n2980 & ~n3015;
  assign n3017 = ~n2960 & ~n2964;
  assign n3018 = ~n2965 & ~n3017;
  assign n3019 = ~n3016 & n3018;
  assign n3020 = ~n2965 & ~n3019;
  assign n3021 = ~n2947 & ~n2949;
  assign n3022 = ~n2950 & ~n3021;
  assign n3023 = ~n3020 & n3022;
  assign n3024 = ~n2950 & ~n3023;
  assign n3025 = ~n2934 & ~n2936;
  assign n3026 = ~n2937 & ~n3025;
  assign n3027 = ~n3024 & n3026;
  assign n3028 = ~n2937 & ~n3027;
  assign n3029 = ~n2919 & n2923;
  assign n3030 = ~n2924 & ~n3029;
  assign n3031 = ~n3028 & n3030;
  assign n3032 = ~n2924 & ~n3031;
  assign n3033 = ~n2898 & ~n2908;
  assign n3034 = n2898 & n2908;
  assign n3035 = ~n3033 & ~n3034;
  assign n3036 = ~n3032 & ~n3035;
  assign n3037 = ~n2909 & ~n3036;
  assign n3038 = ~n2890 & n2894;
  assign n3039 = ~n2895 & ~n3038;
  assign n3040 = ~n3037 & n3039;
  assign n3041 = ~n2895 & ~n3040;
  assign n3042 = ~n2875 & ~n2877;
  assign n3043 = ~n2878 & ~n3042;
  assign n3044 = ~n3041 & n3043;
  assign n3045 = ~n2878 & ~n3044;
  assign n3046 = ~n2547 & ~n2862;
  assign n3047 = ~n2863 & ~n3046;
  assign n3048 = ~n3045 & n3047;
  assign n3049 = ~n2863 & ~n3048;
  assign n3050 = n2400 & n2443;
  assign n3051 = n2402 & ~n2532;
  assign n3052 = ~n2533 & ~n2536;
  assign n3053 = ~n295 & n2028;
  assign n3054 = ~n346 & n3053;
  assign n3055 = ~n114 & ~n163;
  assign n3056 = ~n284 & ~n287;
  assign n3057 = ~n348 & n3056;
  assign n3058 = n3055 & n3057;
  assign n3059 = ~n515 & n3058;
  assign n3060 = ~n255 & n3059;
  assign n3061 = n3054 & n3060;
  assign n3062 = n610 & ~n635;
  assign n3063 = ~n240 & n3062;
  assign n3064 = ~n367 & n3063;
  assign n3065 = ~n468 & n3064;
  assign n3066 = ~n173 & ~n187;
  assign n3067 = ~n535 & n3066;
  assign n3068 = ~n304 & n3067;
  assign n3069 = n3065 & n3068;
  assign n3070 = n3061 & n3069;
  assign n3071 = ~n174 & n3070;
  assign n3072 = ~n568 & n3071;
  assign n3073 = ~n338 & n461;
  assign n3074 = ~n213 & n3073;
  assign n3075 = n3072 & n3074;
  assign n3076 = ~n186 & n717;
  assign n3077 = n482 & n3076;
  assign n3078 = ~n198 & n3077;
  assign n3079 = ~n205 & n3078;
  assign n3080 = ~n123 & ~n476;
  assign n3081 = ~n127 & n3080;
  assign n3082 = n2175 & n3081;
  assign n3083 = ~n548 & n3082;
  assign n3084 = ~n218 & n3083;
  assign n3085 = n3079 & n3084;
  assign n3086 = n3075 & n3085;
  assign n3087 = ~n2530 & n3086;
  assign n3088 = n2530 & ~n3086;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090 = ~n2532 & n3089;
  assign n3091 = n2532 & n3086;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = ~n3052 & n3092;
  assign n3094 = n3052 & ~n3092;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = n2445 & n3095;
  assign n3097 = n2540 & n3089;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = ~n3051 & n3098;
  assign n3100 = ~n3050 & n3099;
  assign n3101 = ~n57 & ~n3100;
  assign n3102 = n57 & n3100;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = ~n2857 & ~n2860;
  assign n3105 = n2451 & n2681;
  assign n3106 = n2448 & n2683;
  assign n3107 = n2687 & n2882;
  assign n3108 = n2384 & n2689;
  assign n3109 = ~n3107 & ~n3108;
  assign n3110 = ~n3106 & n3109;
  assign n3111 = ~n3105 & n3110;
  assign n3112 = n509 & n3111;
  assign n3113 = ~n509 & ~n3111;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = ~n2839 & ~n2843;
  assign n3116 = n2460 & n2566;
  assign n3117 = n2457 & n2554;
  assign n3118 = n2561 & n2703;
  assign n3119 = n2454 & n2559;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = ~n3117 & n3120;
  assign n3122 = ~n3116 & n3121;
  assign n3123 = ~n585 & ~n3122;
  assign n3124 = n585 & n3122;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = n2466 & n2587;
  assign n3127 = n2463 & n2582;
  assign n3128 = n2563 & n2580;
  assign n3129 = n2469 & n2652;
  assign n3130 = ~n3128 & ~n3129;
  assign n3131 = ~n3127 & n3130;
  assign n3132 = ~n3126 & n3131;
  assign n3133 = ~n741 & ~n2475;
  assign n3134 = ~n3132 & n3133;
  assign n3135 = n3132 & ~n3133;
  assign n3136 = ~n3134 & ~n3135;
  assign n3137 = n2830 & ~n2834;
  assign n3138 = ~n2833 & ~n3137;
  assign n3139 = n3136 & n3138;
  assign n3140 = ~n3136 & ~n3138;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = n3125 & n3141;
  assign n3143 = ~n3125 & ~n3141;
  assign n3144 = ~n3142 & ~n3143;
  assign n3145 = ~n3115 & n3144;
  assign n3146 = n3115 & ~n3144;
  assign n3147 = ~n3145 & ~n3146;
  assign n3148 = n3114 & n3147;
  assign n3149 = ~n3114 & ~n3147;
  assign n3150 = ~n3148 & ~n3149;
  assign n3151 = ~n3104 & n3150;
  assign n3152 = n3104 & ~n3150;
  assign n3153 = ~n3151 & ~n3152;
  assign n3154 = n3103 & n3153;
  assign n3155 = ~n3103 & ~n3153;
  assign n3156 = ~n3154 & ~n3155;
  assign n3157 = ~n3049 & n3156;
  assign n3158 = n3049 & ~n3156;
  assign n3159 = ~n3157 & ~n3158;
  assign n3160 = n2530 & n3086;
  assign n3161 = n574 & n2231;
  assign n3162 = ~n325 & n3161;
  assign n3163 = n236 & ~n243;
  assign n3164 = n621 & n3163;
  assign n3165 = ~n293 & n3164;
  assign n3166 = ~n303 & n3165;
  assign n3167 = n3162 & n3166;
  assign n3168 = ~n469 & n3167;
  assign n3169 = n398 & n2013;
  assign n3170 = ~n262 & n3169;
  assign n3171 = n2134 & n3170;
  assign n3172 = n3168 & n3171;
  assign n3173 = n3160 & n3172;
  assign n3174 = ~n3160 & ~n3172;
  assign n3175 = ~n3173 & ~n3174;
  assign n3176 = pi2  & n2389;
  assign n3177 = ~n3175 & n3176;
  assign n3178 = pi0  & ~pi22 ;
  assign n3179 = pi1  & ~n3178;
  assign n3180 = ~pi1  & n3178;
  assign n3181 = ~n3179 & ~n3180;
  assign n3182 = ~pi0  & ~n3181;
  assign n3183 = ~n214 & ~n225;
  assign n3184 = n134 & n211;
  assign n3185 = n534 & n3184;
  assign n3186 = n178 & n574;
  assign n3187 = ~n150 & n3186;
  assign n3188 = n3185 & n3187;
  assign n3189 = n3183 & n3188;
  assign n3190 = n526 & n988;
  assign n3191 = n131 & n3190;
  assign n3192 = n521 & n3191;
  assign n3193 = n3189 & n3192;
  assign n3194 = ~n3173 & n3193;
  assign n3195 = n3173 & ~n3193;
  assign n3196 = ~n3194 & ~n3195;
  assign n3197 = n3182 & n3196;
  assign n3198 = n2392 & n3181;
  assign n3199 = ~n2392 & ~n3181;
  assign n3200 = ~n3198 & ~n3199;
  assign n3201 = pi0  & n3200;
  assign n3202 = ~n3175 & n3196;
  assign n3203 = n3089 & ~n3175;
  assign n3204 = ~n3090 & ~n3093;
  assign n3205 = ~n3089 & n3172;
  assign n3206 = ~n3203 & ~n3205;
  assign n3207 = ~n3204 & n3206;
  assign n3208 = ~n3203 & ~n3207;
  assign n3209 = n3175 & n3193;
  assign n3210 = ~n3202 & ~n3209;
  assign n3211 = ~n3208 & n3210;
  assign n3212 = ~n3202 & ~n3211;
  assign n3213 = n3173 & n3193;
  assign n3214 = ~n381 & n522;
  assign n3215 = ~n199 & n3214;
  assign n3216 = ~n197 & n3215;
  assign n3217 = n156 & ~n541;
  assign n3218 = n557 & n574;
  assign n3219 = n3217 & n3218;
  assign n3220 = n234 & n3219;
  assign n3221 = n3216 & n3220;
  assign n3222 = ~n3213 & ~n3221;
  assign n3223 = n3213 & n3221;
  assign n3224 = ~n3222 & ~n3223;
  assign n3225 = n3196 & ~n3224;
  assign n3226 = ~n3196 & n3221;
  assign n3227 = ~n3225 & ~n3226;
  assign n3228 = ~n3212 & n3227;
  assign n3229 = n3212 & ~n3227;
  assign n3230 = ~n3228 & ~n3229;
  assign n3231 = n3201 & n3230;
  assign n3232 = pi0  & ~n3200;
  assign n3233 = ~n3224 & n3232;
  assign n3234 = ~n3231 & ~n3233;
  assign n3235 = ~n3197 & n3234;
  assign n3236 = ~n3177 & n3235;
  assign n3237 = n2392 & n3236;
  assign n3238 = ~n2392 & ~n3236;
  assign n3239 = ~n3237 & ~n3238;
  assign n3240 = n3159 & n3239;
  assign n3241 = n3045 & ~n3047;
  assign n3242 = ~n3048 & ~n3241;
  assign n3243 = n3089 & n3176;
  assign n3244 = ~n3175 & n3182;
  assign n3245 = n3208 & ~n3210;
  assign n3246 = ~n3211 & ~n3245;
  assign n3247 = n3201 & n3246;
  assign n3248 = n3196 & n3232;
  assign n3249 = ~n3247 & ~n3248;
  assign n3250 = ~n3244 & n3249;
  assign n3251 = ~n3243 & n3250;
  assign n3252 = n2392 & n3251;
  assign n3253 = ~n2392 & ~n3251;
  assign n3254 = ~n3252 & ~n3253;
  assign n3255 = n3242 & n3254;
  assign n3256 = n3041 & ~n3043;
  assign n3257 = ~n3044 & ~n3256;
  assign n3258 = ~n2532 & n3176;
  assign n3259 = n3089 & n3182;
  assign n3260 = n3204 & ~n3206;
  assign n3261 = ~n3207 & ~n3260;
  assign n3262 = n3201 & n3261;
  assign n3263 = ~n3175 & n3232;
  assign n3264 = ~n3262 & ~n3263;
  assign n3265 = ~n3259 & n3264;
  assign n3266 = ~n3258 & n3265;
  assign n3267 = n2392 & n3266;
  assign n3268 = ~n2392 & ~n3266;
  assign n3269 = ~n3267 & ~n3268;
  assign n3270 = n3257 & n3269;
  assign n3271 = ~n3257 & ~n3269;
  assign n3272 = ~n3270 & ~n3271;
  assign n3273 = n3037 & ~n3039;
  assign n3274 = ~n3040 & ~n3273;
  assign n3275 = n3032 & n3035;
  assign n3276 = ~n3036 & ~n3275;
  assign n3277 = n3028 & ~n3030;
  assign n3278 = ~n3031 & ~n3277;
  assign n3279 = n3024 & ~n3026;
  assign n3280 = ~n3027 & ~n3279;
  assign n3281 = n3020 & ~n3022;
  assign n3282 = ~n3023 & ~n3281;
  assign n3283 = n3016 & ~n3018;
  assign n3284 = ~n3019 & ~n3283;
  assign n3285 = n3012 & ~n3014;
  assign n3286 = ~n3015 & ~n3285;
  assign n3287 = n2466 & n3176;
  assign n3288 = n2463 & n3182;
  assign n3289 = n2642 & n3201;
  assign n3290 = n2460 & n3232;
  assign n3291 = ~n3289 & ~n3290;
  assign n3292 = ~n3288 & n3291;
  assign n3293 = ~n3287 & n3292;
  assign n3294 = n2392 & ~n3293;
  assign n3295 = ~n2392 & n3293;
  assign n3296 = ~n3294 & ~n3295;
  assign n3297 = ~n57 & n2981;
  assign n3298 = ~n2987 & n3297;
  assign n3299 = n2987 & ~n3297;
  assign n3300 = ~n3298 & ~n3299;
  assign n3301 = n2475 & n3232;
  assign n3302 = ~n2392 & n3201;
  assign n3303 = ~n2610 & n3302;
  assign n3304 = ~n2472 & n3176;
  assign n3305 = n2475 & n3182;
  assign n3306 = n2469 & n3232;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = ~n3304 & n3307;
  assign n3309 = ~n2392 & ~n3308;
  assign n3310 = ~n2576 & n3302;
  assign n3311 = ~n2392 & ~n3310;
  assign n3312 = ~n3309 & n3311;
  assign n3313 = ~n3303 & n3312;
  assign n3314 = ~n2389 & ~n2472;
  assign n3315 = n3313 & ~n3314;
  assign n3316 = ~n3301 & n3315;
  assign n3317 = n2981 & n3316;
  assign n3318 = ~n2981 & ~n3316;
  assign n3319 = n2466 & n3232;
  assign n3320 = n2624 & n3201;
  assign n3321 = n2469 & n3182;
  assign n3322 = ~n3320 & ~n3321;
  assign n3323 = ~n3319 & n3322;
  assign n3324 = n2392 & ~n3323;
  assign n3325 = n2475 & n3176;
  assign n3326 = n3323 & ~n3325;
  assign n3327 = ~n2392 & n3326;
  assign n3328 = ~n3324 & ~n3327;
  assign n3329 = ~n3318 & ~n3328;
  assign n3330 = ~n3317 & ~n3329;
  assign n3331 = ~n3300 & n3330;
  assign n3332 = n3300 & ~n3330;
  assign n3333 = n2563 & n3201;
  assign n3334 = n2466 & n3182;
  assign n3335 = n2463 & n3232;
  assign n3336 = n2469 & n3176;
  assign n3337 = ~n3335 & ~n3336;
  assign n3338 = ~n3334 & n3337;
  assign n3339 = ~n3333 & n3338;
  assign n3340 = n2392 & n3339;
  assign n3341 = ~n2392 & ~n3339;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = ~n3332 & ~n3342;
  assign n3344 = ~n3331 & ~n3343;
  assign n3345 = ~n3296 & n3344;
  assign n3346 = n3296 & ~n3344;
  assign n3347 = ~n57 & ~n2988;
  assign n3348 = ~n2995 & ~n3347;
  assign n3349 = n2995 & n3347;
  assign n3350 = ~n3348 & ~n3349;
  assign n3351 = ~n3346 & ~n3350;
  assign n3352 = ~n3345 & ~n3351;
  assign n3353 = n2722 & n3201;
  assign n3354 = n2463 & n3176;
  assign n3355 = n2460 & n3182;
  assign n3356 = n2457 & n3232;
  assign n3357 = ~n3355 & ~n3356;
  assign n3358 = ~n3354 & n3357;
  assign n3359 = ~n3353 & n3358;
  assign n3360 = n2392 & n3359;
  assign n3361 = ~n2392 & ~n3359;
  assign n3362 = ~n3360 & ~n3361;
  assign n3363 = n3352 & ~n3362;
  assign n3364 = n3000 & ~n3010;
  assign n3365 = ~n3011 & ~n3364;
  assign n3366 = ~n3363 & n3365;
  assign n3367 = ~n3352 & n3362;
  assign n3368 = ~n3366 & ~n3367;
  assign n3369 = ~n3286 & n3368;
  assign n3370 = n3286 & ~n3368;
  assign n3371 = n2460 & n3176;
  assign n3372 = n2457 & n3182;
  assign n3373 = n2703 & n3201;
  assign n3374 = n2454 & n3232;
  assign n3375 = ~n3373 & ~n3374;
  assign n3376 = ~n3372 & n3375;
  assign n3377 = ~n3371 & n3376;
  assign n3378 = n2392 & ~n3377;
  assign n3379 = ~n2392 & n3377;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = ~n3370 & n3380;
  assign n3382 = ~n3369 & ~n3381;
  assign n3383 = ~n3284 & ~n3382;
  assign n3384 = n3284 & n3382;
  assign n3385 = n2686 & n3201;
  assign n3386 = n2457 & n3176;
  assign n3387 = n2454 & n3182;
  assign n3388 = n2451 & n3232;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = ~n3386 & n3389;
  assign n3391 = ~n3385 & n3390;
  assign n3392 = n2392 & n3391;
  assign n3393 = ~n2392 & ~n3391;
  assign n3394 = ~n3392 & ~n3393;
  assign n3395 = ~n3384 & ~n3394;
  assign n3396 = ~n3383 & ~n3395;
  assign n3397 = ~n3282 & ~n3396;
  assign n3398 = n3282 & n3396;
  assign n3399 = n2848 & n3201;
  assign n3400 = n2454 & n3176;
  assign n3401 = n2451 & n3182;
  assign n3402 = n2448 & n3232;
  assign n3403 = ~n3401 & ~n3402;
  assign n3404 = ~n3400 & n3403;
  assign n3405 = ~n3399 & n3404;
  assign n3406 = n2392 & n3405;
  assign n3407 = ~n2392 & ~n3405;
  assign n3408 = ~n3406 & ~n3407;
  assign n3409 = ~n3398 & ~n3408;
  assign n3410 = ~n3397 & ~n3409;
  assign n3411 = ~n3280 & ~n3410;
  assign n3412 = n3280 & n3410;
  assign n3413 = n2882 & n3201;
  assign n3414 = n2451 & n3176;
  assign n3415 = n2448 & n3182;
  assign n3416 = n2384 & n3232;
  assign n3417 = ~n3415 & ~n3416;
  assign n3418 = ~n3414 & n3417;
  assign n3419 = ~n3413 & n3418;
  assign n3420 = n2392 & n3419;
  assign n3421 = ~n2392 & ~n3419;
  assign n3422 = ~n3420 & ~n3421;
  assign n3423 = ~n3412 & ~n3422;
  assign n3424 = ~n3411 & ~n3423;
  assign n3425 = ~n3278 & ~n3424;
  assign n3426 = n3278 & n3424;
  assign n3427 = n2448 & n3176;
  assign n3428 = n2384 & n3182;
  assign n3429 = n2867 & n3201;
  assign n3430 = n2443 & n3232;
  assign n3431 = ~n3429 & ~n3430;
  assign n3432 = ~n3428 & n3431;
  assign n3433 = ~n3427 & n3432;
  assign n3434 = n2392 & ~n3433;
  assign n3435 = ~n2392 & n3433;
  assign n3436 = ~n3434 & ~n3435;
  assign n3437 = ~n3426 & n3436;
  assign n3438 = ~n3425 & ~n3437;
  assign n3439 = n3276 & n3438;
  assign n3440 = ~n3276 & ~n3438;
  assign n3441 = n2384 & n3176;
  assign n3442 = n2443 & n3182;
  assign n3443 = n2538 & n3201;
  assign n3444 = ~n2532 & n3232;
  assign n3445 = ~n3443 & ~n3444;
  assign n3446 = ~n3442 & n3445;
  assign n3447 = ~n3441 & n3446;
  assign n3448 = ~n2392 & ~n3447;
  assign n3449 = n2392 & n3447;
  assign n3450 = ~n3448 & ~n3449;
  assign n3451 = ~n3440 & n3450;
  assign n3452 = ~n3439 & ~n3451;
  assign n3453 = ~n3274 & n3452;
  assign n3454 = n3274 & ~n3452;
  assign n3455 = n2443 & n3176;
  assign n3456 = ~n2532 & n3182;
  assign n3457 = n3095 & n3201;
  assign n3458 = n3089 & n3232;
  assign n3459 = ~n3457 & ~n3458;
  assign n3460 = ~n3456 & n3459;
  assign n3461 = ~n3455 & n3460;
  assign n3462 = n2392 & ~n3461;
  assign n3463 = ~n2392 & n3461;
  assign n3464 = ~n3462 & ~n3463;
  assign n3465 = ~n3454 & n3464;
  assign n3466 = ~n3453 & ~n3465;
  assign n3467 = n3272 & n3466;
  assign n3468 = ~n3270 & ~n3467;
  assign n3469 = ~n3242 & ~n3254;
  assign n3470 = ~n3255 & ~n3469;
  assign n3471 = ~n3468 & n3470;
  assign n3472 = ~n3255 & ~n3471;
  assign n3473 = ~n3159 & ~n3239;
  assign n3474 = ~n3240 & ~n3473;
  assign n3475 = ~n3472 & n3474;
  assign n3476 = ~n3240 & ~n3475;
  assign n3477 = n3176 & n3196;
  assign n3478 = n3182 & ~n3224;
  assign n3479 = ~n3225 & ~n3228;
  assign n3480 = ~n258 & n2411;
  assign n3481 = ~n192 & n3480;
  assign n3482 = ~n446 & n3481;
  assign n3483 = n705 & n2231;
  assign n3484 = ~n449 & n3483;
  assign n3485 = ~n670 & n3484;
  assign n3486 = n3482 & n3485;
  assign n3487 = n350 & n3486;
  assign n3488 = ~n320 & n712;
  assign n3489 = ~n133 & ~n386;
  assign n3490 = n3488 & n3489;
  assign n3491 = ~n127 & n3490;
  assign n3492 = ~n262 & ~n332;
  assign n3493 = ~n232 & n3492;
  assign n3494 = ~n254 & n3493;
  assign n3495 = n3491 & n3494;
  assign n3496 = ~n119 & n3495;
  assign n3497 = ~n407 & n3496;
  assign n3498 = n1006 & n3497;
  assign n3499 = n3487 & n3498;
  assign n3500 = ~n3223 & n3499;
  assign n3501 = n3223 & ~n3499;
  assign n3502 = ~n3500 & ~n3501;
  assign n3503 = ~n3224 & n3502;
  assign n3504 = n3224 & n3499;
  assign n3505 = ~n3503 & ~n3504;
  assign n3506 = ~n3479 & n3505;
  assign n3507 = n3479 & ~n3505;
  assign n3508 = ~n3506 & ~n3507;
  assign n3509 = n3201 & n3508;
  assign n3510 = n3232 & n3502;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = ~n3478 & n3511;
  assign n3513 = ~n3477 & n3512;
  assign n3514 = n2392 & ~n3513;
  assign n3515 = ~n2392 & n3513;
  assign n3516 = ~n3514 & ~n3515;
  assign n3517 = ~n3154 & ~n3157;
  assign n3518 = ~n3148 & ~n3151;
  assign n3519 = n2448 & n2681;
  assign n3520 = n2384 & n2683;
  assign n3521 = n2687 & n2867;
  assign n3522 = n2443 & n2689;
  assign n3523 = ~n3521 & ~n3522;
  assign n3524 = ~n3520 & n3523;
  assign n3525 = ~n3519 & n3524;
  assign n3526 = n509 & ~n3525;
  assign n3527 = ~n509 & n3525;
  assign n3528 = ~n3526 & ~n3527;
  assign n3529 = ~n3142 & ~n3145;
  assign n3530 = ~n741 & ~n2469;
  assign n3531 = n2466 & n2652;
  assign n3532 = n2463 & n2587;
  assign n3533 = n2580 & n2642;
  assign n3534 = n2460 & n2582;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = ~n3532 & n3535;
  assign n3537 = ~n3531 & n3536;
  assign n3538 = n3530 & ~n3537;
  assign n3539 = ~n3530 & n3537;
  assign n3540 = ~n3538 & ~n3539;
  assign n3541 = ~n741 & n2475;
  assign n3542 = n3132 & n3541;
  assign n3543 = ~n3139 & ~n3542;
  assign n3544 = n3540 & ~n3543;
  assign n3545 = ~n3540 & n3543;
  assign n3546 = ~n3544 & ~n3545;
  assign n3547 = n2457 & n2566;
  assign n3548 = n2454 & n2554;
  assign n3549 = n2561 & n2686;
  assign n3550 = n2451 & n2559;
  assign n3551 = ~n3549 & ~n3550;
  assign n3552 = ~n3548 & n3551;
  assign n3553 = ~n3547 & n3552;
  assign n3554 = n585 & n3553;
  assign n3555 = ~n585 & ~n3553;
  assign n3556 = ~n3554 & ~n3555;
  assign n3557 = n3546 & n3556;
  assign n3558 = ~n3546 & ~n3556;
  assign n3559 = ~n3557 & ~n3558;
  assign n3560 = ~n3529 & n3559;
  assign n3561 = n3529 & ~n3559;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = ~n3528 & n3562;
  assign n3564 = n3528 & ~n3562;
  assign n3565 = ~n3563 & ~n3564;
  assign n3566 = n3518 & ~n3565;
  assign n3567 = ~n3518 & n3565;
  assign n3568 = ~n3566 & ~n3567;
  assign n3569 = n2400 & ~n2532;
  assign n3570 = n2402 & n3089;
  assign n3571 = n2445 & n3261;
  assign n3572 = n2540 & ~n3175;
  assign n3573 = ~n3571 & ~n3572;
  assign n3574 = ~n3570 & n3573;
  assign n3575 = ~n3569 & n3574;
  assign n3576 = n57 & n3575;
  assign n3577 = ~n57 & ~n3575;
  assign n3578 = ~n3576 & ~n3577;
  assign n3579 = n3568 & n3578;
  assign n3580 = ~n3568 & ~n3578;
  assign n3581 = ~n3579 & ~n3580;
  assign n3582 = ~n3517 & n3581;
  assign n3583 = n3517 & ~n3581;
  assign n3584 = ~n3582 & ~n3583;
  assign n3585 = ~n3516 & n3584;
  assign n3586 = n3516 & ~n3584;
  assign n3587 = ~n3585 & ~n3586;
  assign n3588 = n3476 & ~n3587;
  assign n3589 = ~n3476 & n3587;
  assign n3590 = ~n3588 & ~n3589;
  assign n3591 = n640 & n952;
  assign n3592 = ~n248 & n3591;
  assign n3593 = ~n186 & n3592;
  assign n3594 = n790 & n3081;
  assign n3595 = n611 & n1310;
  assign n3596 = n3492 & n3595;
  assign n3597 = ~n317 & n3596;
  assign n3598 = n3594 & n3597;
  assign n3599 = n2114 & n3598;
  assign n3600 = n3593 & n3599;
  assign n3601 = ~n3590 & n3600;
  assign n3602 = n3590 & ~n3600;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = n3472 & ~n3474;
  assign n3605 = ~n3475 & ~n3604;
  assign n3606 = n722 & n2404;
  assign n3607 = ~n327 & n3606;
  assign n3608 = ~n303 & ~n449;
  assign n3609 = ~n185 & n3608;
  assign n3610 = ~n218 & n3492;
  assign n3611 = ~n195 & n2031;
  assign n3612 = ~n274 & n3611;
  assign n3613 = n3610 & n3612;
  assign n3614 = ~n132 & n3613;
  assign n3615 = ~n407 & ~n541;
  assign n3616 = ~n201 & n3615;
  assign n3617 = ~n139 & n175;
  assign n3618 = n3616 & n3617;
  assign n3619 = ~n192 & n3618;
  assign n3620 = ~n197 & n3619;
  assign n3621 = ~n450 & n3620;
  assign n3622 = ~n470 & n3621;
  assign n3623 = n3614 & n3622;
  assign n3624 = ~n535 & n3623;
  assign n3625 = n3609 & n3624;
  assign n3626 = n416 & n3625;
  assign n3627 = ~n294 & n3626;
  assign n3628 = ~n204 & n3627;
  assign n3629 = n3607 & n3628;
  assign n3630 = ~n232 & n3081;
  assign n3631 = ~n468 & n3630;
  assign n3632 = ~n339 & n684;
  assign n3633 = ~n147 & n3058;
  assign n3634 = n200 & n3633;
  assign n3635 = n3632 & n3634;
  assign n3636 = ~n304 & n3635;
  assign n3637 = ~n183 & n3636;
  assign n3638 = n3631 & n3637;
  assign n3639 = n3629 & n3638;
  assign n3640 = ~n3605 & n3639;
  assign n3641 = n3605 & ~n3639;
  assign n3642 = n3468 & ~n3470;
  assign n3643 = ~n3471 & ~n3642;
  assign n3644 = ~n130 & n422;
  assign n3645 = ~n346 & n3644;
  assign n3646 = ~n194 & n613;
  assign n3647 = ~n263 & n554;
  assign n3648 = ~n281 & n3647;
  assign n3649 = ~n450 & n3648;
  assign n3650 = ~n302 & n1021;
  assign n3651 = ~n254 & n3650;
  assign n3652 = ~n186 & ~n470;
  assign n3653 = n3651 & n3652;
  assign n3654 = n2161 & n3653;
  assign n3655 = n3649 & n3654;
  assign n3656 = n3646 & n3655;
  assign n3657 = ~n445 & n3656;
  assign n3658 = ~n295 & n3657;
  assign n3659 = ~n532 & n3658;
  assign n3660 = n3645 & n3659;
  assign n3661 = ~n149 & ~n198;
  assign n3662 = ~n333 & n3661;
  assign n3663 = ~n468 & n3662;
  assign n3664 = ~n133 & n611;
  assign n3665 = ~n360 & n3664;
  assign n3666 = ~n169 & ~n205;
  assign n3667 = n3665 & n3666;
  assign n3668 = ~n304 & ~n477;
  assign n3669 = ~n316 & ~n337;
  assign n3670 = ~n351 & n3669;
  assign n3671 = n3668 & n3670;
  assign n3672 = n3667 & n3671;
  assign n3673 = n3663 & n3672;
  assign n3674 = ~n469 & n3673;
  assign n3675 = ~n227 & n3674;
  assign n3676 = ~n338 & n2267;
  assign n3677 = ~n415 & n3676;
  assign n3678 = ~n318 & n3677;
  assign n3679 = n3675 & n3678;
  assign n3680 = n3660 & n3679;
  assign n3681 = ~n3643 & n3680;
  assign n3682 = n3643 & ~n3680;
  assign n3683 = ~n3272 & ~n3466;
  assign n3684 = ~n3467 & ~n3683;
  assign n3685 = n2156 & n2216;
  assign n3686 = ~n326 & n3685;
  assign n3687 = n763 & n2226;
  assign n3688 = n536 & n3687;
  assign n3689 = ~n119 & n3688;
  assign n3690 = ~n142 & n3689;
  assign n3691 = n3686 & n3690;
  assign n3692 = ~n182 & n2081;
  assign n3693 = ~n379 & n3692;
  assign n3694 = ~n249 & ~n568;
  assign n3695 = n131 & n3694;
  assign n3696 = n2093 & n3695;
  assign n3697 = n3693 & n3696;
  assign n3698 = ~n187 & n3697;
  assign n3699 = ~n205 & n3698;
  assign n3700 = ~n161 & n2419;
  assign n3701 = ~n227 & n3700;
  assign n3702 = n623 & n3701;
  assign n3703 = ~n197 & n3702;
  assign n3704 = ~n195 & n3703;
  assign n3705 = n3699 & n3704;
  assign n3706 = n3691 & n3705;
  assign n3707 = n3684 & ~n3706;
  assign n3708 = ~n3682 & ~n3707;
  assign n3709 = ~n3681 & ~n3708;
  assign n3710 = ~n3641 & ~n3709;
  assign n3711 = ~n3640 & ~n3710;
  assign n3712 = n3603 & n3711;
  assign n3713 = ~n3603 & ~n3711;
  assign n3714 = ~n3712 & ~n3713;
  assign n3715 = ~n3640 & ~n3641;
  assign n3716 = n3709 & ~n3715;
  assign n3717 = ~n3709 & n3715;
  assign n3718 = ~n3716 & ~n3717;
  assign n3719 = n3714 & n3718;
  assign n3720 = ~n3714 & ~n3718;
  assign po0  = n3719 | n3720;
  assign n3722 = ~n3602 & ~n3712;
  assign n3723 = ~n3585 & ~n3589;
  assign n3724 = n3176 & ~n3224;
  assign n3725 = n3182 & n3502;
  assign n3726 = ~n3503 & ~n3506;
  assign n3727 = n671 & n1298;
  assign n3728 = n306 & n3727;
  assign n3729 = ~n635 & n3728;
  assign n3730 = n398 & n625;
  assign n3731 = ~n318 & n3730;
  assign n3732 = n3729 & n3731;
  assign n3733 = ~n270 & n3732;
  assign n3734 = ~n339 & n447;
  assign n3735 = ~n294 & n3734;
  assign n3736 = n544 & n2031;
  assign n3737 = n678 & n3736;
  assign n3738 = n2216 & n3737;
  assign n3739 = n3735 & n3738;
  assign n3740 = ~n302 & n2238;
  assign n3741 = n3739 & n3740;
  assign n3742 = n3733 & n3741;
  assign n3743 = ~n3502 & ~n3742;
  assign n3744 = n3223 & n3499;
  assign n3745 = n3742 & ~n3744;
  assign n3746 = ~n3742 & n3744;
  assign n3747 = ~n3745 & ~n3746;
  assign n3748 = n3502 & ~n3747;
  assign n3749 = ~n3743 & ~n3748;
  assign n3750 = ~n3726 & ~n3749;
  assign n3751 = n3726 & n3749;
  assign n3752 = ~n3750 & ~n3751;
  assign n3753 = n3201 & n3752;
  assign n3754 = n3232 & n3747;
  assign n3755 = ~n3753 & ~n3754;
  assign n3756 = ~n3725 & n3755;
  assign n3757 = ~n3724 & n3756;
  assign n3758 = n2392 & ~n3757;
  assign n3759 = ~n2392 & n3757;
  assign n3760 = ~n3758 & ~n3759;
  assign n3761 = ~n3579 & ~n3582;
  assign n3762 = ~n3563 & ~n3567;
  assign n3763 = n2384 & n2681;
  assign n3764 = n2443 & n2683;
  assign n3765 = n2538 & n2687;
  assign n3766 = ~n2532 & n2689;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = ~n3764 & n3767;
  assign n3769 = ~n3763 & n3768;
  assign n3770 = n509 & ~n3769;
  assign n3771 = ~n509 & n3769;
  assign n3772 = ~n3770 & ~n3771;
  assign n3773 = ~n3557 & ~n3560;
  assign n3774 = ~n741 & ~n2466;
  assign n3775 = n2463 & n2652;
  assign n3776 = n2460 & n2587;
  assign n3777 = n2580 & n2722;
  assign n3778 = n2457 & n2582;
  assign n3779 = ~n3777 & ~n3778;
  assign n3780 = ~n3776 & n3779;
  assign n3781 = ~n3775 & n3780;
  assign n3782 = n3774 & ~n3781;
  assign n3783 = ~n3774 & n3781;
  assign n3784 = ~n3782 & ~n3783;
  assign n3785 = ~n741 & n3537;
  assign n3786 = n2469 & n3785;
  assign n3787 = ~n3544 & ~n3786;
  assign n3788 = ~n3784 & ~n3787;
  assign n3789 = n3784 & n3787;
  assign n3790 = ~n3788 & ~n3789;
  assign n3791 = n2454 & n2566;
  assign n3792 = n2451 & n2554;
  assign n3793 = n2561 & n2848;
  assign n3794 = n2448 & n2559;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = ~n3792 & n3795;
  assign n3797 = ~n3791 & n3796;
  assign n3798 = n585 & n3797;
  assign n3799 = ~n585 & ~n3797;
  assign n3800 = ~n3798 & ~n3799;
  assign n3801 = ~n3790 & ~n3800;
  assign n3802 = n3790 & n3800;
  assign n3803 = ~n3801 & ~n3802;
  assign n3804 = ~n3773 & n3803;
  assign n3805 = n3773 & ~n3803;
  assign n3806 = ~n3804 & ~n3805;
  assign n3807 = ~n3772 & ~n3806;
  assign n3808 = n3772 & n3806;
  assign n3809 = ~n3807 & ~n3808;
  assign n3810 = n3762 & ~n3809;
  assign n3811 = ~n3762 & n3809;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = n2400 & n3089;
  assign n3814 = n2402 & ~n3175;
  assign n3815 = n2445 & n3246;
  assign n3816 = n2540 & n3196;
  assign n3817 = ~n3815 & ~n3816;
  assign n3818 = ~n3814 & n3817;
  assign n3819 = ~n3813 & n3818;
  assign n3820 = n57 & n3819;
  assign n3821 = ~n57 & ~n3819;
  assign n3822 = ~n3820 & ~n3821;
  assign n3823 = n3812 & n3822;
  assign n3824 = ~n3812 & ~n3822;
  assign n3825 = ~n3823 & ~n3824;
  assign n3826 = ~n3761 & n3825;
  assign n3827 = n3761 & ~n3825;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = ~n3760 & n3828;
  assign n3830 = n3760 & ~n3828;
  assign n3831 = ~n3829 & ~n3830;
  assign n3832 = n3723 & ~n3831;
  assign n3833 = ~n3723 & n3831;
  assign n3834 = ~n3832 & ~n3833;
  assign n3835 = n2061 & n3081;
  assign n3836 = ~n254 & n3835;
  assign n3837 = ~n150 & ~n225;
  assign n3838 = ~n548 & n3837;
  assign n3839 = ~n293 & n3838;
  assign n3840 = n786 & n3839;
  assign n3841 = ~n168 & n3840;
  assign n3842 = ~n287 & n3841;
  assign n3843 = n3836 & n3842;
  assign n3844 = n2135 & n3063;
  assign n3845 = ~n161 & n3844;
  assign n3846 = n447 & n3623;
  assign n3847 = ~n130 & n3846;
  assign n3848 = ~n294 & n3847;
  assign n3849 = n3845 & n3848;
  assign n3850 = n3843 & n3849;
  assign n3851 = ~n3834 & n3850;
  assign n3852 = n3834 & ~n3850;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = ~n3722 & n3853;
  assign n3855 = n3722 & ~n3853;
  assign n3856 = ~n3854 & ~n3855;
  assign n3857 = pi22  & ~pi23 ;
  assign n3858 = ~pi22  & pi23 ;
  assign n3859 = ~n3857 & ~n3858;
  assign n3860 = po0  & ~n3859;
  assign n3861 = ~n3856 & n3860;
  assign n3862 = n3714 & ~n3718;
  assign n3863 = n3856 & n3862;
  assign n3864 = ~n3856 & ~n3862;
  assign n3865 = ~n3863 & ~n3864;
  assign n3866 = ~n3860 & n3865;
  assign po1  = n3861 | n3866;
  assign n3868 = ~n3852 & ~n3854;
  assign n3869 = ~n3829 & ~n3833;
  assign n3870 = ~n3747 & n3750;
  assign n3871 = ~n3502 & ~n3506;
  assign n3872 = n3747 & n3871;
  assign n3873 = ~n3870 & ~n3872;
  assign n3874 = n3201 & ~n3873;
  assign n3875 = n3182 & n3747;
  assign n3876 = n3176 & n3502;
  assign n3877 = ~n3875 & ~n3876;
  assign n3878 = ~n3874 & n3877;
  assign n3879 = n2392 & ~n3878;
  assign n3880 = ~n2392 & n3878;
  assign n3881 = ~n3879 & ~n3880;
  assign n3882 = ~n3823 & ~n3826;
  assign n3883 = ~n3807 & ~n3811;
  assign n3884 = n2443 & n2681;
  assign n3885 = ~n2532 & n2683;
  assign n3886 = n2687 & n3095;
  assign n3887 = n2689 & n3089;
  assign n3888 = ~n3886 & ~n3887;
  assign n3889 = ~n3885 & n3888;
  assign n3890 = ~n3884 & n3889;
  assign n3891 = n509 & ~n3890;
  assign n3892 = ~n509 & n3890;
  assign n3893 = ~n3891 & ~n3892;
  assign n3894 = ~n3790 & n3800;
  assign n3895 = ~n3773 & ~n3803;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = ~n741 & ~n2463;
  assign n3898 = n2460 & n2652;
  assign n3899 = n2457 & n2587;
  assign n3900 = n2580 & n2703;
  assign n3901 = n2454 & n2582;
  assign n3902 = ~n3900 & ~n3901;
  assign n3903 = ~n3899 & n3902;
  assign n3904 = ~n3898 & n3903;
  assign n3905 = n3897 & ~n3904;
  assign n3906 = ~n3897 & n3904;
  assign n3907 = ~n3905 & ~n3906;
  assign n3908 = n3784 & ~n3787;
  assign n3909 = ~n741 & n3781;
  assign n3910 = n2466 & n3909;
  assign n3911 = ~n3908 & ~n3910;
  assign n3912 = ~n3907 & ~n3911;
  assign n3913 = n3907 & n3911;
  assign n3914 = ~n3912 & ~n3913;
  assign n3915 = n2451 & n2566;
  assign n3916 = n2448 & n2554;
  assign n3917 = n2561 & n2882;
  assign n3918 = n2384 & n2559;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~n3916 & n3919;
  assign n3921 = ~n3915 & n3920;
  assign n3922 = n585 & n3921;
  assign n3923 = ~n585 & ~n3921;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = ~n3914 & ~n3924;
  assign n3926 = n3914 & n3924;
  assign n3927 = ~n3925 & ~n3926;
  assign n3928 = ~n3896 & n3927;
  assign n3929 = n3896 & ~n3927;
  assign n3930 = ~n3928 & ~n3929;
  assign n3931 = ~n3893 & ~n3930;
  assign n3932 = n3893 & n3930;
  assign n3933 = ~n3931 & ~n3932;
  assign n3934 = n3883 & ~n3933;
  assign n3935 = ~n3883 & n3933;
  assign n3936 = ~n3934 & ~n3935;
  assign n3937 = n2400 & ~n3175;
  assign n3938 = n2402 & n3196;
  assign n3939 = n2445 & n3230;
  assign n3940 = n2540 & ~n3224;
  assign n3941 = ~n3939 & ~n3940;
  assign n3942 = ~n3938 & n3941;
  assign n3943 = ~n3937 & n3942;
  assign n3944 = n57 & n3943;
  assign n3945 = ~n57 & ~n3943;
  assign n3946 = ~n3944 & ~n3945;
  assign n3947 = n3936 & n3946;
  assign n3948 = ~n3936 & ~n3946;
  assign n3949 = ~n3947 & ~n3948;
  assign n3950 = ~n3882 & n3949;
  assign n3951 = n3882 & ~n3949;
  assign n3952 = ~n3950 & ~n3951;
  assign n3953 = ~n3881 & n3952;
  assign n3954 = n3881 & ~n3952;
  assign n3955 = ~n3953 & ~n3954;
  assign n3956 = ~n3869 & n3955;
  assign n3957 = n3869 & ~n3955;
  assign n3958 = ~n3956 & ~n3957;
  assign n3959 = n188 & n776;
  assign n3960 = ~n477 & n3959;
  assign n3961 = ~n183 & ~n446;
  assign n3962 = ~n139 & n3961;
  assign n3963 = ~n221 & n2408;
  assign n3964 = ~n333 & n3963;
  assign n3965 = n3962 & n3964;
  assign n3966 = ~n524 & n3965;
  assign n3967 = ~n133 & n3966;
  assign n3968 = ~n532 & n3967;
  assign n3969 = n3960 & n3968;
  assign n3970 = ~n635 & n3969;
  assign n3971 = ~n325 & n661;
  assign n3972 = ~n445 & n3971;
  assign n3973 = n3697 & n3972;
  assign n3974 = n3970 & n3973;
  assign n3975 = n3958 & ~n3974;
  assign n3976 = ~n3958 & n3974;
  assign n3977 = ~n3975 & ~n3976;
  assign n3978 = n3868 & n3977;
  assign n3979 = ~n3868 & ~n3977;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = ~n3863 & n3980;
  assign n3982 = n3863 & ~n3980;
  assign n3983 = ~n3981 & ~n3982;
  assign n3984 = ~po0  & ~n3865;
  assign n3985 = ~n3859 & ~n3984;
  assign n3986 = n3983 & ~n3985;
  assign n3987 = ~n3983 & n3985;
  assign po2  = n3986 | n3987;
  assign n3989 = ~n3983 & n3984;
  assign n3990 = ~n3859 & ~n3989;
  assign n3991 = ~n3953 & ~n3956;
  assign n3992 = ~n3947 & ~n3950;
  assign n3993 = n3201 & ~n3871;
  assign n3994 = ~n3176 & ~n3993;
  assign n3995 = n3747 & ~n3994;
  assign n3996 = n2392 & n3995;
  assign n3997 = ~n2392 & ~n3995;
  assign n3998 = ~n3996 & ~n3997;
  assign n3999 = ~n3931 & ~n3935;
  assign n4000 = ~n2532 & n2681;
  assign n4001 = n2683 & n3089;
  assign n4002 = n2687 & n3261;
  assign n4003 = n2689 & ~n3175;
  assign n4004 = ~n4002 & ~n4003;
  assign n4005 = ~n4001 & n4004;
  assign n4006 = ~n4000 & n4005;
  assign n4007 = n509 & ~n4006;
  assign n4008 = ~n509 & n4006;
  assign n4009 = ~n4007 & ~n4008;
  assign n4010 = ~n3914 & n3924;
  assign n4011 = ~n3896 & ~n3927;
  assign n4012 = ~n4010 & ~n4011;
  assign n4013 = ~n741 & ~n2460;
  assign n4014 = n2457 & n2652;
  assign n4015 = n2454 & n2587;
  assign n4016 = n2580 & n2686;
  assign n4017 = n2451 & n2582;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = ~n4015 & n4018;
  assign n4020 = ~n4014 & n4019;
  assign n4021 = n4013 & ~n4020;
  assign n4022 = ~n4013 & n4020;
  assign n4023 = ~n4021 & ~n4022;
  assign n4024 = n3907 & ~n3911;
  assign n4025 = ~n741 & n3904;
  assign n4026 = n2463 & n4025;
  assign n4027 = ~n4024 & ~n4026;
  assign n4028 = ~n4023 & ~n4027;
  assign n4029 = n4023 & n4027;
  assign n4030 = ~n4028 & ~n4029;
  assign n4031 = n2448 & n2566;
  assign n4032 = n2384 & n2554;
  assign n4033 = n2561 & n2867;
  assign n4034 = n2443 & n2559;
  assign n4035 = ~n4033 & ~n4034;
  assign n4036 = ~n4032 & n4035;
  assign n4037 = ~n4031 & n4036;
  assign n4038 = n585 & n4037;
  assign n4039 = ~n585 & ~n4037;
  assign n4040 = ~n4038 & ~n4039;
  assign n4041 = ~n4030 & n4040;
  assign n4042 = n4030 & ~n4040;
  assign n4043 = ~n4041 & ~n4042;
  assign n4044 = ~n4012 & n4043;
  assign n4045 = n4012 & ~n4043;
  assign n4046 = ~n4044 & ~n4045;
  assign n4047 = ~n4009 & n4046;
  assign n4048 = n4009 & ~n4046;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = n3999 & ~n4049;
  assign n4051 = ~n3999 & n4049;
  assign n4052 = ~n4050 & ~n4051;
  assign n4053 = n2400 & n3196;
  assign n4054 = n2402 & ~n3224;
  assign n4055 = n2445 & n3508;
  assign n4056 = n2540 & n3502;
  assign n4057 = ~n4055 & ~n4056;
  assign n4058 = ~n4054 & n4057;
  assign n4059 = ~n4053 & n4058;
  assign n4060 = n57 & n4059;
  assign n4061 = ~n57 & ~n4059;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = n4052 & n4062;
  assign n4064 = ~n4052 & ~n4062;
  assign n4065 = ~n4063 & ~n4064;
  assign n4066 = ~n3998 & n4065;
  assign n4067 = n3998 & ~n4065;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = ~n3992 & n4068;
  assign n4070 = n3992 & ~n4068;
  assign n4071 = ~n4069 & ~n4070;
  assign n4072 = ~n3991 & n4071;
  assign n4073 = n3991 & ~n4071;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = n439 & n2135;
  assign n4076 = ~n332 & n4075;
  assign n4077 = n131 & n3671;
  assign n4078 = n286 & n4077;
  assign n4079 = ~n119 & n4078;
  assign n4080 = ~n168 & n4079;
  assign n4081 = n4076 & n4080;
  assign n4082 = ~n255 & n2070;
  assign n4083 = ~n293 & n4082;
  assign n4084 = n707 & n1316;
  assign n4085 = ~n327 & n4084;
  assign n4086 = n4083 & n4085;
  assign n4087 = n4081 & n4086;
  assign n4088 = ~n4074 & ~n4087;
  assign n4089 = n4074 & n4087;
  assign n4090 = ~n4088 & ~n4089;
  assign n4091 = n3868 & ~n3975;
  assign n4092 = ~n3976 & ~n4091;
  assign n4093 = ~n4090 & n4092;
  assign n4094 = n4090 & ~n4092;
  assign n4095 = ~n4093 & ~n4094;
  assign n4096 = n3982 & n4095;
  assign n4097 = ~n3982 & ~n4095;
  assign n4098 = ~n4096 & ~n4097;
  assign n4099 = n3990 & n4098;
  assign n4100 = ~n3990 & ~n4098;
  assign po3  = ~n4099 & ~n4100;
  assign n4102 = n4074 & ~n4087;
  assign n4103 = ~n4093 & ~n4102;
  assign n4104 = ~n4069 & ~n4072;
  assign n4105 = ~n4063 & ~n4066;
  assign n4106 = ~n4047 & ~n4051;
  assign n4107 = ~n4041 & ~n4044;
  assign n4108 = n2454 & n2652;
  assign n4109 = n2451 & n2587;
  assign n4110 = n2580 & n2848;
  assign n4111 = n2448 & n2582;
  assign n4112 = ~n4110 & ~n4111;
  assign n4113 = ~n4109 & n4112;
  assign n4114 = ~n4108 & n4113;
  assign n4115 = n741 & ~n4114;
  assign n4116 = ~n741 & n4114;
  assign n4117 = ~n4115 & ~n4116;
  assign n4118 = ~n741 & n2457;
  assign n4119 = ~n2392 & n4118;
  assign n4120 = n2392 & ~n4118;
  assign n4121 = ~n4119 & ~n4120;
  assign n4122 = ~n4117 & n4121;
  assign n4123 = n4117 & ~n4121;
  assign n4124 = ~n4122 & ~n4123;
  assign n4125 = n4023 & ~n4027;
  assign n4126 = ~n741 & n4020;
  assign n4127 = n2460 & n4126;
  assign n4128 = ~n4125 & ~n4127;
  assign n4129 = ~n4124 & ~n4128;
  assign n4130 = n4124 & n4128;
  assign n4131 = ~n4129 & ~n4130;
  assign n4132 = n2384 & n2566;
  assign n4133 = n2443 & n2554;
  assign n4134 = n2538 & n2561;
  assign n4135 = ~n2532 & n2559;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = ~n4133 & n4136;
  assign n4138 = ~n4132 & n4137;
  assign n4139 = ~n585 & ~n4138;
  assign n4140 = n585 & n4138;
  assign n4141 = ~n4139 & ~n4140;
  assign n4142 = ~n4131 & ~n4141;
  assign n4143 = n4131 & n4141;
  assign n4144 = ~n4142 & ~n4143;
  assign n4145 = ~n4107 & n4144;
  assign n4146 = n4107 & ~n4144;
  assign n4147 = ~n4145 & ~n4146;
  assign n4148 = n2681 & n3089;
  assign n4149 = n2683 & ~n3175;
  assign n4150 = n2687 & n3246;
  assign n4151 = n2689 & n3196;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = ~n4149 & n4152;
  assign n4154 = ~n4148 & n4153;
  assign n4155 = ~n509 & n4154;
  assign n4156 = n509 & ~n4154;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~n4147 & ~n4157;
  assign n4159 = n4147 & n4157;
  assign n4160 = ~n4158 & ~n4159;
  assign n4161 = ~n4106 & n4160;
  assign n4162 = n4106 & ~n4160;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = n2400 & ~n3224;
  assign n4165 = n2402 & n3502;
  assign n4166 = n2445 & n3752;
  assign n4167 = n2540 & n3747;
  assign n4168 = ~n4166 & ~n4167;
  assign n4169 = ~n4165 & n4168;
  assign n4170 = ~n4164 & n4169;
  assign n4171 = ~n57 & ~n4170;
  assign n4172 = n57 & n4170;
  assign n4173 = ~n4171 & ~n4172;
  assign n4174 = n4163 & n4173;
  assign n4175 = ~n4163 & ~n4173;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = ~n4105 & n4176;
  assign n4178 = n4105 & ~n4176;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180 = n4104 & ~n4179;
  assign n4181 = ~n4104 & n4179;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = ~n163 & n761;
  assign n4184 = ~n172 & n4183;
  assign n4185 = n395 & n4184;
  assign n4186 = n2231 & n2270;
  assign n4187 = n619 & n2408;
  assign n4188 = n296 & n4187;
  assign n4189 = ~n271 & n4188;
  assign n4190 = n4186 & n4189;
  assign n4191 = n490 & n4190;
  assign n4192 = n4185 & n4191;
  assign n4193 = ~n4182 & n4192;
  assign n4194 = n4182 & ~n4192;
  assign n4195 = ~n4193 & ~n4194;
  assign n4196 = ~n4103 & n4195;
  assign n4197 = n4103 & ~n4195;
  assign n4198 = ~n4196 & ~n4197;
  assign n4199 = ~n4096 & ~n4198;
  assign n4200 = n4096 & n4198;
  assign n4201 = ~n4199 & ~n4200;
  assign n4202 = n3989 & ~n4098;
  assign n4203 = ~n3859 & ~n4202;
  assign n4204 = n4201 & ~n4203;
  assign n4205 = ~n4201 & n4203;
  assign po4  = n4204 | n4205;
  assign n4207 = ~n4194 & ~n4196;
  assign n4208 = ~n4177 & ~n4181;
  assign n4209 = ~n4161 & ~n4174;
  assign n4210 = n2445 & ~n3873;
  assign n4211 = n2402 & n3747;
  assign n4212 = n2400 & n3502;
  assign n4213 = ~n4211 & ~n4212;
  assign n4214 = ~n4210 & n4213;
  assign n4215 = ~n57 & ~n4214;
  assign n4216 = n57 & n4214;
  assign n4217 = ~n4215 & ~n4216;
  assign n4218 = ~n4107 & ~n4144;
  assign n4219 = ~n4158 & ~n4218;
  assign n4220 = n2681 & ~n3175;
  assign n4221 = n2683 & n3196;
  assign n4222 = n2687 & n3230;
  assign n4223 = n2689 & ~n3224;
  assign n4224 = ~n4222 & ~n4223;
  assign n4225 = ~n4221 & n4224;
  assign n4226 = ~n4220 & n4225;
  assign n4227 = n509 & ~n4226;
  assign n4228 = ~n509 & n4226;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = ~n4131 & n4141;
  assign n4231 = n4124 & ~n4128;
  assign n4232 = ~n4230 & ~n4231;
  assign n4233 = ~n4119 & ~n4122;
  assign n4234 = ~n741 & ~n2392;
  assign n4235 = n2454 & n4234;
  assign n4236 = ~n2392 & ~n4235;
  assign n4237 = ~n741 & ~n4234;
  assign n4238 = n2454 & n4237;
  assign n4239 = ~n4236 & ~n4238;
  assign n4240 = ~n4233 & n4239;
  assign n4241 = n4233 & ~n4239;
  assign n4242 = ~n4240 & ~n4241;
  assign n4243 = n2451 & n2652;
  assign n4244 = n2448 & n2587;
  assign n4245 = n2580 & n2882;
  assign n4246 = n2384 & n2582;
  assign n4247 = ~n4245 & ~n4246;
  assign n4248 = ~n4244 & n4247;
  assign n4249 = ~n4243 & n4248;
  assign n4250 = n741 & n4249;
  assign n4251 = ~n741 & ~n4249;
  assign n4252 = ~n4250 & ~n4251;
  assign n4253 = ~n4242 & ~n4252;
  assign n4254 = n4242 & n4252;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = n2443 & n2566;
  assign n4257 = ~n2532 & n2554;
  assign n4258 = n2561 & n3095;
  assign n4259 = n2559 & n3089;
  assign n4260 = ~n4258 & ~n4259;
  assign n4261 = ~n4257 & n4260;
  assign n4262 = ~n4256 & n4261;
  assign n4263 = ~n585 & ~n4262;
  assign n4264 = n585 & n4262;
  assign n4265 = ~n4263 & ~n4264;
  assign n4266 = ~n4255 & n4265;
  assign n4267 = n4255 & ~n4265;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = ~n4232 & ~n4268;
  assign n4270 = n4232 & n4268;
  assign n4271 = ~n4269 & ~n4270;
  assign n4272 = ~n4229 & ~n4271;
  assign n4273 = n4229 & n4271;
  assign n4274 = ~n4272 & ~n4273;
  assign n4275 = ~n4219 & n4274;
  assign n4276 = n4219 & ~n4274;
  assign n4277 = ~n4275 & ~n4276;
  assign n4278 = n4217 & n4277;
  assign n4279 = ~n4217 & ~n4277;
  assign n4280 = ~n4278 & ~n4279;
  assign n4281 = ~n4209 & n4280;
  assign n4282 = n4209 & ~n4280;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = ~n4208 & n4283;
  assign n4285 = n4208 & ~n4283;
  assign n4286 = ~n4284 & ~n4285;
  assign n4287 = n134 & n3839;
  assign n4288 = n2099 & n4287;
  assign n4289 = ~n194 & n616;
  assign n4290 = ~n262 & n4289;
  assign n4291 = n4288 & n4290;
  assign n4292 = n3070 & n3739;
  assign n4293 = ~n217 & n4292;
  assign n4294 = ~n360 & ~n440;
  assign n4295 = ~n119 & n4294;
  assign n4296 = n200 & n4295;
  assign n4297 = n2106 & n4296;
  assign n4298 = ~n172 & n4297;
  assign n4299 = n4293 & n4298;
  assign n4300 = n4291 & n4299;
  assign n4301 = ~n4286 & n4300;
  assign n4302 = n4286 & ~n4300;
  assign n4303 = ~n4301 & ~n4302;
  assign n4304 = ~n4207 & n4303;
  assign n4305 = n4207 & ~n4303;
  assign n4306 = ~n4304 & ~n4305;
  assign n4307 = ~n4200 & ~n4306;
  assign n4308 = n4200 & n4306;
  assign n4309 = ~n4307 & ~n4308;
  assign n4310 = ~n4201 & n4202;
  assign n4311 = ~n3859 & ~n4310;
  assign n4312 = n4309 & ~n4311;
  assign n4313 = ~n4309 & n4311;
  assign po5  = n4312 | n4313;
  assign n4315 = ~n4302 & ~n4304;
  assign n4316 = ~n4281 & ~n4284;
  assign n4317 = ~n4275 & ~n4278;
  assign n4318 = ~n4232 & n4268;
  assign n4319 = ~n4272 & ~n4318;
  assign n4320 = n2445 & ~n3871;
  assign n4321 = ~n2400 & ~n4320;
  assign n4322 = n3747 & ~n4321;
  assign n4323 = n57 & n4322;
  assign n4324 = ~n57 & ~n4322;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = ~n4319 & ~n4325;
  assign n4327 = n4319 & n4325;
  assign n4328 = ~n4326 & ~n4327;
  assign n4329 = n2681 & n3196;
  assign n4330 = n2683 & ~n3224;
  assign n4331 = n2687 & n3508;
  assign n4332 = n2689 & n3502;
  assign n4333 = ~n4331 & ~n4332;
  assign n4334 = ~n4330 & n4333;
  assign n4335 = ~n4329 & n4334;
  assign n4336 = n509 & ~n4335;
  assign n4337 = ~n509 & n4335;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = ~n4242 & n4252;
  assign n4340 = ~n4266 & ~n4339;
  assign n4341 = ~n2532 & n2566;
  assign n4342 = n2554 & n3089;
  assign n4343 = n2561 & n3261;
  assign n4344 = n2559 & ~n3175;
  assign n4345 = ~n4343 & ~n4344;
  assign n4346 = ~n4342 & n4345;
  assign n4347 = ~n4341 & n4346;
  assign n4348 = ~n585 & ~n4347;
  assign n4349 = n585 & n4347;
  assign n4350 = ~n4348 & ~n4349;
  assign n4351 = n2448 & n2652;
  assign n4352 = n2384 & n2587;
  assign n4353 = n2580 & n2867;
  assign n4354 = n2443 & n2582;
  assign n4355 = ~n4353 & ~n4354;
  assign n4356 = ~n4352 & n4355;
  assign n4357 = ~n4351 & n4356;
  assign n4358 = n741 & n4357;
  assign n4359 = ~n741 & ~n4357;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = ~n4233 & ~n4239;
  assign n4362 = ~n4235 & ~n4361;
  assign n4363 = ~n741 & n2451;
  assign n4364 = ~n2392 & n4363;
  assign n4365 = n2392 & ~n4363;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = ~n4362 & n4366;
  assign n4368 = n4362 & ~n4366;
  assign n4369 = ~n4367 & ~n4368;
  assign n4370 = n4360 & n4369;
  assign n4371 = ~n4360 & ~n4369;
  assign n4372 = ~n4370 & ~n4371;
  assign n4373 = n4350 & n4372;
  assign n4374 = ~n4350 & ~n4372;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = ~n4340 & n4375;
  assign n4377 = n4340 & ~n4375;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = ~n4338 & n4378;
  assign n4380 = n4338 & ~n4378;
  assign n4381 = ~n4379 & ~n4380;
  assign n4382 = n4328 & n4381;
  assign n4383 = ~n4328 & ~n4381;
  assign n4384 = ~n4382 & ~n4383;
  assign n4385 = ~n4317 & n4384;
  assign n4386 = n4317 & ~n4384;
  assign n4387 = ~n4385 & ~n4386;
  assign n4388 = ~n4316 & n4387;
  assign n4389 = n4316 & ~n4387;
  assign n4390 = ~n4388 & ~n4389;
  assign n4391 = n387 & n3183;
  assign n4392 = ~n140 & n4391;
  assign n4393 = n368 & n4392;
  assign n4394 = n709 & n717;
  assign n4395 = ~n361 & n4394;
  assign n4396 = n2106 & n4395;
  assign n4397 = n306 & n2234;
  assign n4398 = n398 & n958;
  assign n4399 = n4397 & n4398;
  assign n4400 = n2135 & n4399;
  assign n4401 = n4396 & n4400;
  assign n4402 = ~n248 & n4401;
  assign n4403 = ~n205 & n3625;
  assign n4404 = ~n414 & n4403;
  assign n4405 = n4402 & n4404;
  assign n4406 = n2260 & n4405;
  assign n4407 = n4393 & n4406;
  assign n4408 = ~n4390 & n4407;
  assign n4409 = n4390 & ~n4407;
  assign n4410 = ~n4408 & ~n4409;
  assign n4411 = ~n4315 & n4410;
  assign n4412 = n4315 & ~n4410;
  assign n4413 = ~n4411 & ~n4412;
  assign n4414 = ~n4308 & ~n4413;
  assign n4415 = n4308 & n4413;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = ~n4309 & n4310;
  assign n4418 = ~n3859 & ~n4417;
  assign n4419 = n4416 & ~n4418;
  assign n4420 = ~n4416 & n4418;
  assign po6  = n4419 | n4420;
  assign n4422 = ~n4409 & ~n4411;
  assign n4423 = ~n4385 & ~n4388;
  assign n4424 = ~n4326 & ~n4382;
  assign n4425 = ~n4376 & ~n4379;
  assign n4426 = n2681 & ~n3224;
  assign n4427 = n2683 & n3502;
  assign n4428 = n2687 & n3752;
  assign n4429 = n2689 & n3747;
  assign n4430 = ~n4428 & ~n4429;
  assign n4431 = ~n4427 & n4430;
  assign n4432 = ~n4426 & n4431;
  assign n4433 = n509 & n4432;
  assign n4434 = ~n509 & ~n4432;
  assign n4435 = ~n4433 & ~n4434;
  assign n4436 = ~n4425 & n4435;
  assign n4437 = n4425 & ~n4435;
  assign n4438 = ~n4436 & ~n4437;
  assign n4439 = ~n4370 & ~n4373;
  assign n4440 = n2566 & n3089;
  assign n4441 = n2554 & ~n3175;
  assign n4442 = n2561 & n3246;
  assign n4443 = n2559 & n3196;
  assign n4444 = ~n4442 & ~n4443;
  assign n4445 = ~n4441 & n4444;
  assign n4446 = ~n4440 & n4445;
  assign n4447 = n585 & n4446;
  assign n4448 = ~n585 & ~n4446;
  assign n4449 = ~n4447 & ~n4448;
  assign n4450 = ~n4364 & ~n4367;
  assign n4451 = n2384 & n2652;
  assign n4452 = n2443 & n2587;
  assign n4453 = n2538 & n2580;
  assign n4454 = ~n2532 & n2582;
  assign n4455 = ~n4453 & ~n4454;
  assign n4456 = ~n4452 & n4455;
  assign n4457 = ~n4451 & n4456;
  assign n4458 = n741 & ~n4457;
  assign n4459 = ~n741 & n4457;
  assign n4460 = ~n4458 & ~n4459;
  assign n4461 = ~n741 & n2448;
  assign n4462 = n57 & n2392;
  assign n4463 = ~n57 & ~n2392;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = n4461 & n4464;
  assign n4466 = ~n4461 & ~n4464;
  assign n4467 = ~n4465 & ~n4466;
  assign n4468 = ~n4460 & ~n4467;
  assign n4469 = n4460 & n4467;
  assign n4470 = ~n4468 & ~n4469;
  assign n4471 = ~n4450 & ~n4470;
  assign n4472 = n4450 & n4470;
  assign n4473 = ~n4471 & ~n4472;
  assign n4474 = n4449 & n4473;
  assign n4475 = ~n4449 & ~n4473;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = ~n4439 & n4476;
  assign n4478 = n4439 & ~n4476;
  assign n4479 = ~n4477 & ~n4478;
  assign n4480 = n4438 & n4479;
  assign n4481 = ~n4438 & ~n4479;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = ~n4424 & n4482;
  assign n4484 = n4424 & ~n4482;
  assign n4485 = ~n4483 & ~n4484;
  assign n4486 = n4423 & ~n4485;
  assign n4487 = ~n4423 & n4485;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = ~n227 & n4401;
  assign n4490 = ~n397 & n4489;
  assign n4491 = n940 & n4490;
  assign n4492 = ~n163 & n4295;
  assign n4493 = ~n254 & n4492;
  assign n4494 = n245 & n621;
  assign n4495 = ~n183 & n4494;
  assign n4496 = ~n195 & n4495;
  assign n4497 = n4493 & n4496;
  assign n4498 = n2075 & n4497;
  assign n4499 = n4491 & n4498;
  assign n4500 = n4488 & ~n4499;
  assign n4501 = ~n4488 & n4499;
  assign n4502 = ~n4500 & ~n4501;
  assign n4503 = ~n4422 & n4502;
  assign n4504 = n4422 & ~n4502;
  assign n4505 = ~n4503 & ~n4504;
  assign n4506 = n4415 & n4505;
  assign n4507 = ~n4415 & ~n4505;
  assign n4508 = ~n4506 & ~n4507;
  assign n4509 = ~n4416 & n4417;
  assign n4510 = ~n3859 & ~n4509;
  assign n4511 = n4508 & ~n4510;
  assign n4512 = ~n4508 & n4510;
  assign po7  = n4511 | n4512;
  assign n4514 = ~n4500 & ~n4503;
  assign n4515 = ~n4483 & ~n4487;
  assign n4516 = ~n4436 & ~n4480;
  assign n4517 = n2687 & ~n3873;
  assign n4518 = n2683 & n3747;
  assign n4519 = n2681 & n3502;
  assign n4520 = ~n4518 & ~n4519;
  assign n4521 = ~n4517 & n4520;
  assign n4522 = n509 & ~n4521;
  assign n4523 = ~n509 & n4521;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = ~n4474 & ~n4477;
  assign n4526 = n2566 & ~n3175;
  assign n4527 = n2554 & n3196;
  assign n4528 = n2561 & n3230;
  assign n4529 = n2559 & ~n3224;
  assign n4530 = ~n4528 & ~n4529;
  assign n4531 = ~n4527 & n4530;
  assign n4532 = ~n4526 & n4531;
  assign n4533 = ~n585 & ~n4532;
  assign n4534 = n585 & n4532;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = ~n4460 & n4467;
  assign n4537 = ~n4471 & ~n4536;
  assign n4538 = ~n741 & n2384;
  assign n4539 = ~n4462 & ~n4465;
  assign n4540 = ~n4538 & n4539;
  assign n4541 = n4538 & ~n4539;
  assign n4542 = ~n4540 & ~n4541;
  assign n4543 = n2443 & n2652;
  assign n4544 = ~n2532 & n2587;
  assign n4545 = n2580 & n3095;
  assign n4546 = n2582 & n3089;
  assign n4547 = ~n4545 & ~n4546;
  assign n4548 = ~n4544 & n4547;
  assign n4549 = ~n4543 & n4548;
  assign n4550 = n741 & n4549;
  assign n4551 = ~n741 & ~n4549;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = ~n4542 & n4552;
  assign n4554 = n4542 & ~n4552;
  assign n4555 = ~n4553 & ~n4554;
  assign n4556 = ~n4537 & n4555;
  assign n4557 = n4537 & ~n4555;
  assign n4558 = ~n4556 & ~n4557;
  assign n4559 = n4535 & n4558;
  assign n4560 = ~n4535 & ~n4558;
  assign n4561 = ~n4559 & ~n4560;
  assign n4562 = ~n4525 & n4561;
  assign n4563 = n4525 & ~n4561;
  assign n4564 = ~n4562 & ~n4563;
  assign n4565 = ~n4524 & n4564;
  assign n4566 = n4524 & ~n4564;
  assign n4567 = ~n4565 & ~n4566;
  assign n4568 = ~n4516 & n4567;
  assign n4569 = n4516 & ~n4567;
  assign n4570 = ~n4568 & ~n4569;
  assign n4571 = ~n4515 & n4570;
  assign n4572 = n4515 & ~n4570;
  assign n4573 = ~n4571 & ~n4572;
  assign n4574 = n369 & n401;
  assign n4575 = ~n127 & n4574;
  assign n4576 = ~n221 & n3657;
  assign n4577 = ~n635 & n4576;
  assign n4578 = ~n548 & n4577;
  assign n4579 = n4575 & n4578;
  assign n4580 = ~n541 & n4579;
  assign n4581 = ~n449 & n722;
  assign n4582 = ~n338 & n376;
  assign n4583 = ~n197 & n4582;
  assign n4584 = n4581 & n4583;
  assign n4585 = ~n132 & n4584;
  assign n4586 = ~n201 & n2280;
  assign n4587 = ~n327 & n4586;
  assign n4588 = ~n147 & n4587;
  assign n4589 = n4585 & n4588;
  assign n4590 = ~n228 & n2123;
  assign n4591 = ~n386 & n4590;
  assign n4592 = n4589 & n4591;
  assign n4593 = n4580 & n4592;
  assign n4594 = ~n4573 & n4593;
  assign n4595 = n4573 & ~n4593;
  assign n4596 = ~n4594 & ~n4595;
  assign n4597 = ~n4514 & n4596;
  assign n4598 = n4514 & ~n4596;
  assign n4599 = ~n4597 & ~n4598;
  assign n4600 = ~n4506 & ~n4599;
  assign n4601 = n4506 & n4599;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = ~n4508 & n4509;
  assign n4604 = ~n3859 & ~n4603;
  assign n4605 = n4602 & ~n4604;
  assign n4606 = ~n4602 & n4604;
  assign po8  = n4605 | n4606;
  assign n4608 = ~n4595 & ~n4597;
  assign n4609 = ~n4568 & ~n4571;
  assign n4610 = ~n4562 & ~n4565;
  assign n4611 = ~n4556 & ~n4559;
  assign n4612 = n2687 & ~n3871;
  assign n4613 = ~n2681 & ~n4612;
  assign n4614 = n3747 & ~n4613;
  assign n4615 = ~n509 & ~n4614;
  assign n4616 = n509 & n4614;
  assign n4617 = ~n4615 & ~n4616;
  assign n4618 = ~n4611 & ~n4617;
  assign n4619 = n4611 & n4617;
  assign n4620 = ~n4618 & ~n4619;
  assign n4621 = n2566 & n3196;
  assign n4622 = n2554 & ~n3224;
  assign n4623 = n2561 & n3508;
  assign n4624 = n2559 & n3502;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = ~n4622 & n4625;
  assign n4627 = ~n4621 & n4626;
  assign n4628 = ~n585 & ~n4627;
  assign n4629 = n585 & n4627;
  assign n4630 = ~n4628 & ~n4629;
  assign n4631 = ~n4538 & ~n4539;
  assign n4632 = ~n4553 & ~n4631;
  assign n4633 = ~n2532 & n2652;
  assign n4634 = n2587 & n3089;
  assign n4635 = n2580 & n3261;
  assign n4636 = n2582 & ~n3175;
  assign n4637 = ~n4635 & ~n4636;
  assign n4638 = ~n4634 & n4637;
  assign n4639 = ~n4633 & n4638;
  assign n4640 = n741 & ~n4639;
  assign n4641 = ~n741 & n4639;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = ~n741 & n2510;
  assign n4644 = ~n4642 & ~n4643;
  assign n4645 = n4642 & n4643;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = ~n4632 & n4646;
  assign n4648 = n4632 & ~n4646;
  assign n4649 = ~n4647 & ~n4648;
  assign n4650 = n4630 & n4649;
  assign n4651 = ~n4630 & ~n4649;
  assign n4652 = ~n4650 & ~n4651;
  assign n4653 = n4620 & n4652;
  assign n4654 = ~n4620 & ~n4652;
  assign n4655 = ~n4653 & ~n4654;
  assign n4656 = ~n4610 & n4655;
  assign n4657 = n4610 & ~n4655;
  assign n4658 = ~n4656 & ~n4657;
  assign n4659 = n4609 & ~n4658;
  assign n4660 = ~n4609 & n4658;
  assign n4661 = ~n4659 & ~n4660;
  assign n4662 = n1317 & n3062;
  assign n4663 = ~n265 & n4662;
  assign n4664 = n3183 & n3635;
  assign n4665 = ~n130 & n4664;
  assign n4666 = ~n274 & n4665;
  assign n4667 = n4663 & n4666;
  assign n4668 = ~n201 & n459;
  assign n4669 = ~n169 & n4668;
  assign n4670 = ~n379 & n2238;
  assign n4671 = ~n140 & n4670;
  assign n4672 = n4669 & n4671;
  assign n4673 = n4667 & n4672;
  assign n4674 = ~n4661 & n4673;
  assign n4675 = n4661 & ~n4673;
  assign n4676 = ~n4674 & ~n4675;
  assign n4677 = ~n4608 & n4676;
  assign n4678 = n4608 & ~n4676;
  assign n4679 = ~n4677 & ~n4678;
  assign n4680 = ~n4601 & ~n4679;
  assign n4681 = n4601 & n4679;
  assign n4682 = ~n4680 & ~n4681;
  assign n4683 = ~n4602 & n4603;
  assign n4684 = ~n3859 & ~n4683;
  assign n4685 = n4682 & ~n4684;
  assign n4686 = ~n4682 & n4684;
  assign po9  = n4685 | n4686;
  assign n4688 = ~n4675 & ~n4677;
  assign n4689 = ~n4656 & ~n4660;
  assign n4690 = ~n4618 & ~n4653;
  assign n4691 = ~n4647 & ~n4650;
  assign n4692 = n2566 & ~n3224;
  assign n4693 = n2554 & n3502;
  assign n4694 = n2561 & n3752;
  assign n4695 = n2559 & n3747;
  assign n4696 = ~n4694 & ~n4695;
  assign n4697 = ~n4693 & n4696;
  assign n4698 = ~n4692 & n4697;
  assign n4699 = n585 & n4698;
  assign n4700 = ~n585 & ~n4698;
  assign n4701 = ~n4699 & ~n4700;
  assign n4702 = ~n4691 & n4701;
  assign n4703 = n4691 & ~n4701;
  assign n4704 = ~n4702 & ~n4703;
  assign n4705 = n2652 & n3089;
  assign n4706 = n2587 & ~n3175;
  assign n4707 = n2580 & n3246;
  assign n4708 = n2582 & n3196;
  assign n4709 = ~n4707 & ~n4708;
  assign n4710 = ~n4706 & n4709;
  assign n4711 = ~n4705 & n4710;
  assign n4712 = ~n741 & n4711;
  assign n4713 = n741 & ~n4711;
  assign n4714 = ~n4712 & ~n4713;
  assign n4715 = ~n741 & ~n2532;
  assign n4716 = ~n509 & ~n4715;
  assign n4717 = n509 & n4715;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = n4538 & ~n4718;
  assign n4720 = ~n4538 & n4718;
  assign n4721 = ~n4719 & ~n4720;
  assign n4722 = ~n741 & ~n2384;
  assign n4723 = n2443 & n4722;
  assign n4724 = ~n4644 & ~n4723;
  assign n4725 = ~n4721 & ~n4724;
  assign n4726 = n4721 & n4724;
  assign n4727 = ~n4725 & ~n4726;
  assign n4728 = n4714 & ~n4727;
  assign n4729 = ~n4714 & n4727;
  assign n4730 = ~n4728 & ~n4729;
  assign n4731 = n4704 & n4730;
  assign n4732 = ~n4704 & ~n4730;
  assign n4733 = ~n4731 & ~n4732;
  assign n4734 = ~n4690 & n4733;
  assign n4735 = n4690 & ~n4733;
  assign n4736 = ~n4734 & ~n4735;
  assign n4737 = ~n4689 & n4736;
  assign n4738 = n4689 & ~n4736;
  assign n4739 = ~n4737 & ~n4738;
  assign n4740 = n755 & n3081;
  assign n4741 = ~n348 & n4740;
  assign n4742 = n472 & n2404;
  assign n4743 = n554 & n4742;
  assign n4744 = n3183 & n4743;
  assign n4745 = ~n171 & n4744;
  assign n4746 = n4741 & n4745;
  assign n4747 = ~n305 & n4746;
  assign n4748 = n399 & n954;
  assign n4749 = n3673 & n4748;
  assign n4750 = n4747 & n4749;
  assign n4751 = ~n4739 & n4750;
  assign n4752 = n4739 & ~n4750;
  assign n4753 = ~n4751 & ~n4752;
  assign n4754 = ~n4688 & n4753;
  assign n4755 = n4688 & ~n4753;
  assign n4756 = ~n4754 & ~n4755;
  assign n4757 = ~n4681 & ~n4756;
  assign n4758 = n4681 & n4756;
  assign n4759 = ~n4757 & ~n4758;
  assign n4760 = ~n4682 & n4683;
  assign n4761 = ~n3859 & ~n4760;
  assign n4762 = n4759 & ~n4761;
  assign n4763 = ~n4759 & n4761;
  assign po10  = n4762 | n4763;
  assign n4765 = ~n4752 & ~n4754;
  assign n4766 = ~n4734 & ~n4737;
  assign n4767 = ~n4702 & ~n4731;
  assign n4768 = n2561 & ~n3873;
  assign n4769 = n2554 & n3747;
  assign n4770 = n2566 & n3502;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = ~n4768 & n4771;
  assign n4773 = ~n585 & ~n4772;
  assign n4774 = n585 & n4772;
  assign n4775 = ~n4773 & ~n4774;
  assign n4776 = n2652 & ~n3175;
  assign n4777 = n2587 & n3196;
  assign n4778 = n2580 & n3230;
  assign n4779 = n2582 & ~n3224;
  assign n4780 = ~n4778 & ~n4779;
  assign n4781 = ~n4777 & n4780;
  assign n4782 = ~n4776 & n4781;
  assign n4783 = n741 & n4782;
  assign n4784 = ~n741 & ~n4782;
  assign n4785 = ~n4783 & ~n4784;
  assign n4786 = ~n741 & n3089;
  assign n4787 = ~n4538 & ~n4717;
  assign n4788 = ~n4716 & ~n4787;
  assign n4789 = ~n4786 & n4788;
  assign n4790 = n4786 & ~n4788;
  assign n4791 = ~n4789 & ~n4790;
  assign n4792 = n4785 & n4791;
  assign n4793 = ~n4785 & ~n4791;
  assign n4794 = ~n4792 & ~n4793;
  assign n4795 = n4714 & ~n4725;
  assign n4796 = ~n4726 & ~n4795;
  assign n4797 = n4794 & n4796;
  assign n4798 = ~n4794 & ~n4796;
  assign n4799 = ~n4797 & ~n4798;
  assign n4800 = n4775 & n4799;
  assign n4801 = ~n4775 & ~n4799;
  assign n4802 = ~n4800 & ~n4801;
  assign n4803 = ~n4767 & n4802;
  assign n4804 = n4767 & ~n4802;
  assign n4805 = ~n4803 & ~n4804;
  assign n4806 = ~n4766 & n4805;
  assign n4807 = n4766 & ~n4805;
  assign n4808 = ~n4806 & ~n4807;
  assign n4809 = n319 & n3495;
  assign n4810 = n391 & n534;
  assign n4811 = n4809 & n4810;
  assign n4812 = ~n226 & n4811;
  assign n4813 = n518 & n784;
  assign n4814 = n4812 & n4813;
  assign n4815 = ~n4808 & n4814;
  assign n4816 = n4808 & ~n4814;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = ~n4765 & n4817;
  assign n4819 = n4765 & ~n4817;
  assign n4820 = ~n4818 & ~n4819;
  assign n4821 = ~n4758 & ~n4820;
  assign n4822 = n4758 & n4820;
  assign n4823 = ~n4821 & ~n4822;
  assign n4824 = ~n4759 & n4760;
  assign n4825 = ~n3859 & ~n4824;
  assign n4826 = n4823 & ~n4825;
  assign n4827 = ~n4823 & n4825;
  assign po11  = n4826 | n4827;
  assign n4829 = ~n4816 & ~n4818;
  assign n4830 = ~n4803 & ~n4806;
  assign n4831 = ~n4797 & ~n4800;
  assign n4832 = n2652 & n3196;
  assign n4833 = n2587 & ~n3224;
  assign n4834 = n2580 & n3508;
  assign n4835 = n2582 & n3502;
  assign n4836 = ~n4834 & ~n4835;
  assign n4837 = ~n4833 & n4836;
  assign n4838 = ~n4832 & n4837;
  assign n4839 = ~n741 & n4838;
  assign n4840 = n741 & ~n4838;
  assign n4841 = ~n4839 & ~n4840;
  assign n4842 = n2561 & ~n3871;
  assign n4843 = ~n2566 & ~n4842;
  assign n4844 = n3747 & ~n4843;
  assign n4845 = n585 & n4844;
  assign n4846 = ~n585 & ~n4844;
  assign n4847 = ~n4845 & ~n4846;
  assign n4848 = ~n4841 & ~n4847;
  assign n4849 = n4841 & n4847;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4789 & ~n4792;
  assign n4852 = ~n741 & ~n3175;
  assign n4853 = ~n3089 & n4852;
  assign n4854 = n3175 & n4786;
  assign n4855 = ~n4853 & ~n4854;
  assign n4856 = n4851 & ~n4855;
  assign n4857 = ~n4851 & n4855;
  assign n4858 = ~n4856 & ~n4857;
  assign n4859 = n4850 & n4858;
  assign n4860 = ~n4850 & ~n4858;
  assign n4861 = ~n4859 & ~n4860;
  assign n4862 = ~n4831 & n4861;
  assign n4863 = n4831 & ~n4861;
  assign n4864 = ~n4862 & ~n4863;
  assign n4865 = ~n4830 & n4864;
  assign n4866 = n4830 & ~n4864;
  assign n4867 = ~n4865 & ~n4866;
  assign n4868 = ~n214 & n2018;
  assign n4869 = ~n149 & n4868;
  assign n4870 = n2165 & n2170;
  assign n4871 = ~n127 & ~n198;
  assign n4872 = ~n295 & n4871;
  assign n4873 = ~n265 & ~n349;
  assign n4874 = n4872 & n4873;
  assign n4875 = n286 & n4874;
  assign n4876 = ~n449 & n4875;
  assign n4877 = n4870 & n4876;
  assign n4878 = n3965 & n4877;
  assign n4879 = n4869 & n4878;
  assign n4880 = ~n4867 & n4879;
  assign n4881 = n4867 & ~n4879;
  assign n4882 = ~n4880 & ~n4881;
  assign n4883 = ~n4829 & n4882;
  assign n4884 = n4829 & ~n4882;
  assign n4885 = ~n4883 & ~n4884;
  assign n4886 = ~n4822 & ~n4885;
  assign n4887 = n4822 & n4885;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = ~n4823 & n4824;
  assign n4890 = ~n3859 & ~n4889;
  assign n4891 = n4888 & ~n4890;
  assign n4892 = ~n4888 & n4890;
  assign po12  = n4891 | n4892;
  assign n4894 = ~n4881 & ~n4883;
  assign n4895 = ~n4862 & ~n4865;
  assign n4896 = ~n4848 & ~n4859;
  assign n4897 = n2652 & ~n3224;
  assign n4898 = n2587 & n3502;
  assign n4899 = n2580 & n3752;
  assign n4900 = n2582 & n3747;
  assign n4901 = ~n4899 & ~n4900;
  assign n4902 = ~n4898 & n4901;
  assign n4903 = ~n4897 & n4902;
  assign n4904 = n741 & ~n4903;
  assign n4905 = ~n741 & n4903;
  assign n4906 = ~n4904 & ~n4905;
  assign n4907 = n585 & n4852;
  assign n4908 = ~n585 & ~n4852;
  assign n4909 = ~n4907 & ~n4908;
  assign n4910 = ~n741 & n3196;
  assign n4911 = n4909 & n4910;
  assign n4912 = ~n4909 & ~n4910;
  assign n4913 = ~n4911 & ~n4912;
  assign n4914 = ~n4906 & ~n4913;
  assign n4915 = n4906 & n4913;
  assign n4916 = ~n4914 & ~n4915;
  assign n4917 = ~n4851 & ~n4853;
  assign n4918 = ~n4854 & ~n4917;
  assign n4919 = ~n4916 & ~n4918;
  assign n4920 = n4916 & n4918;
  assign n4921 = ~n4919 & ~n4920;
  assign n4922 = ~n4896 & n4921;
  assign n4923 = n4896 & ~n4921;
  assign n4924 = ~n4922 & ~n4923;
  assign n4925 = ~n4895 & n4924;
  assign n4926 = n4895 & ~n4924;
  assign n4927 = ~n4925 & ~n4926;
  assign n4928 = n966 & n3697;
  assign n4929 = ~n366 & n4928;
  assign n4930 = ~n166 & ~n365;
  assign n4931 = ~n186 & ~n294;
  assign n4932 = ~n163 & n4931;
  assign n4933 = n4930 & n4932;
  assign n4934 = n717 & n4933;
  assign n4935 = ~n228 & n4934;
  assign n4936 = ~n297 & n4935;
  assign n4937 = n4929 & n4936;
  assign n4938 = ~n114 & n3839;
  assign n4939 = ~n333 & n4938;
  assign n4940 = n422 & n2369;
  assign n4941 = ~n539 & n4940;
  assign n4942 = ~n318 & n4941;
  assign n4943 = n4939 & n4942;
  assign n4944 = n4937 & n4943;
  assign n4945 = n4927 & ~n4944;
  assign n4946 = ~n4927 & n4944;
  assign n4947 = ~n4945 & ~n4946;
  assign n4948 = n4894 & n4947;
  assign n4949 = ~n4894 & ~n4947;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = ~n4887 & n4950;
  assign n4952 = n4887 & ~n4950;
  assign n4953 = ~n4951 & ~n4952;
  assign n4954 = ~n4888 & n4889;
  assign n4955 = ~n3859 & ~n4954;
  assign n4956 = n4953 & ~n4955;
  assign n4957 = ~n4953 & n4955;
  assign po13  = n4956 | n4957;
  assign n4959 = ~n4922 & ~n4925;
  assign n4960 = ~n4906 & n4913;
  assign n4961 = ~n4919 & ~n4960;
  assign n4962 = ~n741 & ~n3224;
  assign n4963 = ~n4907 & ~n4911;
  assign n4964 = ~n4962 & n4963;
  assign n4965 = n4962 & ~n4963;
  assign n4966 = ~n4964 & ~n4965;
  assign n4967 = n2580 & ~n3873;
  assign n4968 = n2587 & n3747;
  assign n4969 = n2652 & n3502;
  assign n4970 = ~n4968 & ~n4969;
  assign n4971 = ~n4967 & n4970;
  assign n4972 = n741 & n4971;
  assign n4973 = ~n741 & ~n4971;
  assign n4974 = ~n4972 & ~n4973;
  assign n4975 = ~n4966 & n4974;
  assign n4976 = n4966 & ~n4974;
  assign n4977 = ~n4975 & ~n4976;
  assign n4978 = ~n4961 & n4977;
  assign n4979 = n4961 & ~n4977;
  assign n4980 = ~n4978 & ~n4979;
  assign n4981 = ~n4959 & n4980;
  assign n4982 = n4959 & ~n4980;
  assign n4983 = ~n4981 & ~n4982;
  assign n4984 = n372 & n523;
  assign n4985 = n2170 & n4984;
  assign n4986 = ~n213 & n4985;
  assign n4987 = ~n477 & n4986;
  assign n4988 = n424 & n2216;
  assign n4989 = ~n226 & n4988;
  assign n4990 = ~n539 & n4989;
  assign n4991 = n4987 & n4990;
  assign n4992 = n653 & n4991;
  assign n4993 = n1324 & n3183;
  assign n4994 = ~n219 & n4993;
  assign n4995 = n2287 & n4994;
  assign n4996 = n4992 & n4995;
  assign n4997 = ~n4983 & n4996;
  assign n4998 = n4983 & ~n4996;
  assign n4999 = ~n4997 & ~n4998;
  assign n5000 = n4894 & ~n4945;
  assign n5001 = ~n4946 & ~n5000;
  assign n5002 = n4999 & n5001;
  assign n5003 = ~n4999 & ~n5001;
  assign n5004 = ~n5002 & ~n5003;
  assign n5005 = ~n4952 & ~n5004;
  assign n5006 = n4952 & n5004;
  assign n5007 = ~n5005 & ~n5006;
  assign n5008 = ~n4953 & n4954;
  assign n5009 = ~n3859 & ~n5008;
  assign n5010 = n5007 & ~n5009;
  assign n5011 = ~n5007 & n5009;
  assign po14  = n5010 | n5011;
  assign n5013 = ~n4998 & ~n5002;
  assign n5014 = n2580 & ~n3871;
  assign n5015 = ~n2652 & ~n5014;
  assign n5016 = n3747 & ~n5015;
  assign n5017 = n741 & n5016;
  assign n5018 = ~n741 & ~n5016;
  assign n5019 = ~n5017 & ~n5018;
  assign n5020 = ~n741 & n3505;
  assign n5021 = n5019 & ~n5020;
  assign n5022 = n3505 & n5018;
  assign n5023 = ~n5021 & ~n5022;
  assign n5024 = ~n4962 & ~n4963;
  assign n5025 = ~n4975 & ~n5024;
  assign n5026 = n5023 & n5025;
  assign n5027 = ~n5023 & ~n5025;
  assign n5028 = ~n5026 & ~n5027;
  assign n5029 = ~n4978 & ~n4981;
  assign n5030 = ~n5028 & n5029;
  assign n5031 = n5028 & ~n5029;
  assign n5032 = ~n5030 & ~n5031;
  assign n5033 = n387 & n937;
  assign n5034 = ~n204 & n5033;
  assign n5035 = ~n140 & n1025;
  assign n5036 = ~n415 & n5035;
  assign n5037 = ~n159 & n5036;
  assign n5038 = n763 & n5037;
  assign n5039 = ~n477 & n5038;
  assign n5040 = ~n470 & n5039;
  assign n5041 = n5034 & n5040;
  assign n5042 = ~n351 & n5041;
  assign n5043 = ~n379 & n2179;
  assign n5044 = ~n173 & n5043;
  assign n5045 = n4874 & n5044;
  assign n5046 = n5042 & n5045;
  assign n5047 = n5032 & ~n5046;
  assign n5048 = ~n5032 & n5046;
  assign n5049 = ~n5047 & ~n5048;
  assign n5050 = n5013 & n5049;
  assign n5051 = ~n5013 & ~n5049;
  assign n5052 = ~n5050 & ~n5051;
  assign n5053 = ~n5006 & n5052;
  assign n5054 = n5006 & ~n5052;
  assign n5055 = ~n5053 & ~n5054;
  assign n5056 = ~n5007 & n5008;
  assign n5057 = ~n3859 & ~n5056;
  assign n5058 = n5055 & ~n5057;
  assign n5059 = ~n5055 & n5057;
  assign po15  = n5058 | n5059;
  assign n5061 = ~n367 & n471;
  assign n5062 = ~n123 & n5061;
  assign n5063 = n3618 & n5062;
  assign n5064 = n2020 & n2105;
  assign n5065 = n250 & n3702;
  assign n5066 = ~n568 & n5065;
  assign n5067 = n5064 & n5066;
  assign n5068 = n4933 & n5067;
  assign n5069 = n5063 & n5068;
  assign n5070 = ~n5019 & ~n5020;
  assign n5071 = ~n741 & n3224;
  assign n5072 = n3502 & n5071;
  assign n5073 = ~n5070 & ~n5072;
  assign n5074 = ~n5027 & ~n5031;
  assign n5075 = ~n3747 & n4962;
  assign n5076 = n3747 & ~n4962;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = ~n741 & n5077;
  assign n5079 = n5074 & ~n5078;
  assign n5080 = ~n5074 & n5078;
  assign n5081 = ~n5079 & ~n5080;
  assign n5082 = n5073 & n5081;
  assign n5083 = ~n5073 & ~n5081;
  assign n5084 = ~n5082 & ~n5083;
  assign n5085 = ~n5069 & n5084;
  assign n5086 = n5069 & ~n5084;
  assign n5087 = ~n5085 & ~n5086;
  assign n5088 = n5013 & ~n5047;
  assign n5089 = ~n5048 & ~n5088;
  assign n5090 = n5087 & ~n5089;
  assign n5091 = ~n5087 & n5089;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = ~n5054 & n5092;
  assign n5094 = n5054 & ~n5092;
  assign n5095 = ~n5093 & ~n5094;
  assign n5096 = ~n5055 & n5056;
  assign n5097 = ~n3859 & ~n5096;
  assign n5098 = n5095 & ~n5097;
  assign n5099 = ~n5095 & n5097;
  assign po16  = n5098 | n5099;
  assign n5101 = ~n5095 & n5096;
  assign n5102 = ~n3859 & ~n5101;
  assign n5103 = ~n5085 & ~n5089;
  assign n5104 = ~n5086 & ~n5103;
  assign n5105 = n691 & n2404;
  assign n5106 = ~n389 & n5105;
  assign n5107 = n340 & n719;
  assign n5108 = ~n127 & n5107;
  assign n5109 = ~n149 & n5108;
  assign n5110 = n5106 & n5109;
  assign n5111 = ~n469 & n5110;
  assign n5112 = n422 & n3070;
  assign n5113 = ~n450 & n5112;
  assign n5114 = n466 & n5113;
  assign n5115 = n5111 & n5114;
  assign n5116 = n5104 & ~n5115;
  assign n5117 = ~n5104 & n5115;
  assign n5118 = ~n5116 & ~n5117;
  assign n5119 = n5094 & n5118;
  assign n5120 = ~n5094 & ~n5118;
  assign n5121 = ~n5119 & ~n5120;
  assign n5122 = n5102 & n5121;
  assign n5123 = ~n5102 & ~n5121;
  assign po17  = ~n5122 & ~n5123;
  assign n5125 = n5101 & ~n5121;
  assign n5126 = ~n3859 & ~n5125;
  assign n5127 = ~n5116 & ~n5119;
  assign n5128 = n973 & n998;
  assign n5129 = ~n213 & n5128;
  assign n5130 = n411 & n5129;
  assign n5131 = n776 & n2361;
  assign n5132 = ~n127 & n5131;
  assign n5133 = n724 & n3655;
  assign n5134 = ~n332 & n5133;
  assign n5135 = n5132 & n5134;
  assign n5136 = n2087 & n5135;
  assign n5137 = n5130 & n5136;
  assign n5138 = ~n5127 & n5137;
  assign n5139 = n5127 & ~n5137;
  assign n5140 = ~n5138 & ~n5139;
  assign n5141 = n5126 & n5140;
  assign n5142 = ~n5126 & ~n5140;
  assign po18  = n5141 | n5142;
  assign n5144 = n5116 & ~n5137;
  assign n5145 = n278 & n765;
  assign n5146 = ~n338 & n5037;
  assign n5147 = n5145 & n5146;
  assign n5148 = ~n206 & n2523;
  assign n5149 = ~n150 & n5148;
  assign n5150 = ~n182 & n4295;
  assign n5151 = ~n445 & n5150;
  assign n5152 = n5149 & n5151;
  assign n5153 = n5147 & n5152;
  assign n5154 = n3080 & n5153;
  assign n5155 = ~n5144 & n5154;
  assign n5156 = n5144 & ~n5154;
  assign n5157 = ~n5155 & ~n5156;
  assign n5158 = n5119 & ~n5137;
  assign n5159 = ~n5157 & ~n5158;
  assign n5160 = n5157 & n5158;
  assign n5161 = ~n5159 & ~n5160;
  assign n5162 = n5125 & n5140;
  assign n5163 = ~n3859 & ~n5162;
  assign n5164 = n5161 & ~n5163;
  assign n5165 = ~n5161 & n5163;
  assign po19  = n5164 | n5165;
  assign n5167 = ~n5161 & n5162;
  assign n5168 = ~n3859 & ~n5167;
  assign n5169 = n200 & n2106;
  assign n5170 = ~n535 & n5169;
  assign n5171 = n429 & n525;
  assign n5172 = ~n171 & n5171;
  assign n5173 = ~n670 & n5172;
  assign n5174 = n5170 & n5173;
  assign n5175 = ~n174 & n521;
  assign n5176 = ~n163 & n5175;
  assign n5177 = ~n195 & n4589;
  assign n5178 = ~n303 & n5177;
  assign n5179 = n5176 & n5178;
  assign n5180 = n5174 & n5179;
  assign n5181 = ~n5156 & ~n5160;
  assign n5182 = n5180 & ~n5181;
  assign n5183 = ~n5180 & n5181;
  assign n5184 = ~n5182 & ~n5183;
  assign n5185 = n5168 & n5184;
  assign n5186 = ~n5168 & ~n5184;
  assign po20  = n5185 | n5186;
  assign n5188 = n5156 & ~n5180;
  assign n5189 = n238 & ~n539;
  assign n5190 = ~n365 & n3214;
  assign n5191 = n576 & n5190;
  assign n5192 = n5189 & n5191;
  assign n5193 = ~n5188 & n5192;
  assign n5194 = n5188 & ~n5192;
  assign n5195 = ~n5193 & ~n5194;
  assign n5196 = n5160 & ~n5180;
  assign n5197 = ~n5195 & ~n5196;
  assign n5198 = n5195 & n5196;
  assign n5199 = ~n5197 & ~n5198;
  assign n5200 = n5167 & n5184;
  assign n5201 = ~n3859 & ~n5200;
  assign n5202 = n5199 & ~n5201;
  assign n5203 = ~n5199 & n5201;
  assign po21  = n5202 | n5203;
  assign n5205 = ~n5199 & n5200;
  assign n5206 = ~n3859 & ~n5205;
  assign n5207 = n238 & n559;
  assign n5208 = ~n5194 & ~n5198;
  assign n5209 = n5207 & ~n5208;
  assign n5210 = ~n5207 & n5208;
  assign n5211 = ~n5209 & ~n5210;
  assign n5212 = n5206 & n5211;
  assign n5213 = ~n5206 & ~n5211;
  assign po22  = n5212 | n5213;
  assign n5215 = ~pi22  & n102;
  assign n5216 = n5205 & n5211;
  assign n5217 = ~n3859 & ~n5216;
  assign n5218 = ~n5207 & ~n5208;
  assign n5219 = n5194 & n5198;
  assign n5220 = n5218 & ~n5219;
  assign n5221 = n5217 & ~n5220;
  assign n5222 = ~n5217 & n5220;
  assign n5223 = ~n5221 & ~n5222;
  assign po23  = n5215 | ~n5223;
  assign n5225 = ~n5207 & n5219;
  assign n5226 = ~n5216 & ~n5225;
  assign n5227 = n5205 & n5218;
  assign n5228 = ~n5215 & ~n5227;
  assign n5229 = ~n5226 & n5228;
  assign po24  = ~n3859 & ~n5229;
endmodule
