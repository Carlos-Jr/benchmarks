module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7;
  wire n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n655, n657, n658, n660, n661,
    n662, n663, n664, n665;
  assign n137 = ~pi124  & ~pi125 ;
  assign n138 = ~pi126  & ~pi127 ;
  assign n139 = n137 & n138;
  assign n140 = ~pi122  & ~pi123 ;
  assign n141 = ~pi120  & ~pi121 ;
  assign n142 = n140 & n141;
  assign n143 = n139 & n142;
  assign n144 = pi123  & n139;
  assign n145 = pi125  & ~pi126 ;
  assign n146 = ~pi127  & ~n145;
  assign n147 = ~n144 & n146;
  assign n148 = pi121  & ~pi122 ;
  assign n149 = n139 & n148;
  assign n150 = n147 & ~n149;
  assign n151 = ~n143 & n150;
  assign n152 = ~pi118  & ~n151;
  assign n153 = ~pi116  & n152;
  assign n154 = ~pi114  & n153;
  assign n155 = pi117  & n152;
  assign n156 = pi119  & n143;
  assign n157 = pi115  & n153;
  assign n158 = n150 & ~n157;
  assign n159 = ~n156 & n158;
  assign n160 = ~n155 & n159;
  assign n161 = ~n154 & n160;
  assign n162 = ~pi112  & ~n161;
  assign n163 = ~pi110  & n162;
  assign n164 = pi111  & ~pi112 ;
  assign n165 = ~pi113  & ~n164;
  assign n166 = n154 & ~n165;
  assign n167 = n160 & ~n166;
  assign n168 = ~n163 & n167;
  assign n169 = ~pi108  & ~n168;
  assign n170 = ~pi106  & n169;
  assign n171 = ~pi104  & n170;
  assign n172 = pi107  & n169;
  assign n173 = pi109  & n163;
  assign n174 = pi105  & n170;
  assign n175 = n167 & ~n174;
  assign n176 = ~n173 & n175;
  assign n177 = ~n172 & n176;
  assign n178 = ~n171 & n177;
  assign n179 = ~pi102  & ~n178;
  assign n180 = ~pi100  & n179;
  assign n181 = pi101  & ~pi102 ;
  assign n182 = ~pi103  & ~n181;
  assign n183 = n171 & ~n182;
  assign n184 = n177 & ~n183;
  assign n185 = ~n180 & n184;
  assign n186 = ~pi98  & ~n185;
  assign n187 = ~pi96  & n186;
  assign n188 = ~pi94  & n187;
  assign n189 = pi97  & n186;
  assign n190 = pi99  & n180;
  assign n191 = pi95  & n187;
  assign n192 = n184 & ~n191;
  assign n193 = ~n190 & n192;
  assign n194 = ~n189 & n193;
  assign n195 = ~n188 & n194;
  assign n196 = ~pi92  & ~n195;
  assign n197 = ~pi90  & n196;
  assign n198 = pi91  & ~pi92 ;
  assign n199 = ~pi93  & ~n198;
  assign n200 = n188 & ~n199;
  assign n201 = n194 & ~n200;
  assign n202 = ~n197 & n201;
  assign n203 = ~pi88  & ~n202;
  assign n204 = ~pi86  & n203;
  assign n205 = ~pi84  & n204;
  assign n206 = pi87  & n203;
  assign n207 = pi89  & n197;
  assign n208 = pi85  & n204;
  assign n209 = n201 & ~n208;
  assign n210 = ~n207 & n209;
  assign n211 = ~n206 & n210;
  assign n212 = ~n205 & n211;
  assign n213 = ~pi82  & ~n212;
  assign n214 = ~pi80  & n213;
  assign n215 = pi81  & ~pi82 ;
  assign n216 = ~pi83  & ~n215;
  assign n217 = n205 & ~n216;
  assign n218 = n211 & ~n217;
  assign n219 = ~n214 & n218;
  assign n220 = ~pi78  & ~n219;
  assign n221 = ~pi76  & n220;
  assign n222 = ~pi74  & n221;
  assign n223 = pi77  & n220;
  assign n224 = pi79  & n214;
  assign n225 = pi75  & n221;
  assign n226 = n218 & ~n225;
  assign n227 = ~n224 & n226;
  assign n228 = ~n223 & n227;
  assign n229 = ~n222 & n228;
  assign n230 = ~pi72  & ~n229;
  assign n231 = ~pi70  & n230;
  assign n232 = pi71  & ~pi72 ;
  assign n233 = ~pi73  & ~n232;
  assign n234 = n222 & ~n233;
  assign n235 = n228 & ~n234;
  assign n236 = ~n231 & n235;
  assign n237 = ~pi68  & ~n236;
  assign n238 = ~pi66  & n237;
  assign n239 = ~pi64  & n238;
  assign n240 = pi67  & n237;
  assign n241 = pi69  & n231;
  assign n242 = pi65  & n238;
  assign n243 = n235 & ~n242;
  assign n244 = ~n241 & n243;
  assign n245 = ~n240 & n244;
  assign n246 = ~n239 & n245;
  assign n247 = ~pi62  & ~n246;
  assign n248 = ~pi60  & n247;
  assign n249 = pi61  & ~pi62 ;
  assign n250 = ~pi63  & ~n249;
  assign n251 = n239 & ~n250;
  assign n252 = n245 & ~n251;
  assign n253 = ~n248 & n252;
  assign n254 = ~pi58  & ~n253;
  assign n255 = ~pi56  & n254;
  assign n256 = ~pi54  & n255;
  assign n257 = pi57  & n254;
  assign n258 = pi59  & n248;
  assign n259 = pi55  & n255;
  assign n260 = n252 & ~n259;
  assign n261 = ~n258 & n260;
  assign n262 = ~n257 & n261;
  assign n263 = ~n256 & n262;
  assign n264 = ~pi52  & ~n263;
  assign n265 = ~pi50  & n264;
  assign n266 = pi51  & ~pi52 ;
  assign n267 = ~pi53  & ~n266;
  assign n268 = n256 & ~n267;
  assign n269 = n262 & ~n268;
  assign n270 = ~n265 & n269;
  assign n271 = ~pi48  & ~n270;
  assign n272 = ~pi46  & n271;
  assign n273 = ~pi44  & n272;
  assign n274 = pi47  & n271;
  assign n275 = pi49  & n265;
  assign n276 = pi45  & n272;
  assign n277 = n269 & ~n276;
  assign n278 = ~n275 & n277;
  assign n279 = ~n274 & n278;
  assign n280 = ~n273 & n279;
  assign n281 = ~pi42  & ~n280;
  assign n282 = ~pi40  & n281;
  assign n283 = pi41  & ~pi42 ;
  assign n284 = ~pi43  & ~n283;
  assign n285 = n273 & ~n284;
  assign n286 = n279 & ~n285;
  assign n287 = ~n282 & n286;
  assign n288 = ~pi38  & ~n287;
  assign n289 = ~pi36  & n288;
  assign n290 = ~pi34  & n289;
  assign n291 = pi37  & n288;
  assign n292 = pi39  & n282;
  assign n293 = pi35  & n289;
  assign n294 = n286 & ~n293;
  assign n295 = ~n292 & n294;
  assign n296 = ~n291 & n295;
  assign n297 = ~n290 & n296;
  assign n298 = ~pi32  & ~n297;
  assign n299 = ~pi30  & n298;
  assign n300 = pi31  & ~pi32 ;
  assign n301 = ~pi33  & ~n300;
  assign n302 = n290 & ~n301;
  assign n303 = n296 & ~n302;
  assign n304 = ~n299 & n303;
  assign n305 = ~pi28  & ~n304;
  assign n306 = ~pi26  & n305;
  assign n307 = ~pi24  & n306;
  assign n308 = pi27  & n305;
  assign n309 = pi29  & n299;
  assign n310 = pi25  & n306;
  assign n311 = n303 & ~n310;
  assign n312 = ~n309 & n311;
  assign n313 = ~n308 & n312;
  assign n314 = ~n307 & n313;
  assign n315 = ~pi22  & ~n314;
  assign n316 = ~pi20  & n315;
  assign n317 = pi21  & ~pi22 ;
  assign n318 = ~pi23  & ~n317;
  assign n319 = n307 & ~n318;
  assign n320 = n313 & ~n319;
  assign n321 = ~n316 & n320;
  assign n322 = ~pi18  & ~n321;
  assign n323 = ~pi16  & n322;
  assign n324 = ~pi14  & n323;
  assign n325 = pi17  & n322;
  assign n326 = pi19  & n316;
  assign n327 = pi15  & n323;
  assign n328 = n320 & ~n327;
  assign n329 = ~n326 & n328;
  assign n330 = ~n325 & n329;
  assign n331 = ~n324 & n330;
  assign n332 = ~pi12  & ~n331;
  assign n333 = ~pi10  & n332;
  assign n334 = pi11  & ~pi12 ;
  assign n335 = ~pi13  & ~n334;
  assign n336 = n324 & ~n335;
  assign n337 = n330 & ~n336;
  assign n338 = ~n333 & n337;
  assign n339 = ~pi8  & ~n338;
  assign n340 = pi7  & n339;
  assign n341 = pi9  & n333;
  assign n342 = ~pi6  & n339;
  assign n343 = pi5  & n342;
  assign n344 = n337 & ~n343;
  assign n345 = ~n341 & n344;
  assign n346 = ~n340 & n345;
  assign n347 = pi1  & ~pi2 ;
  assign n348 = ~pi3  & ~n347;
  assign n349 = ~pi4  & ~n348;
  assign n350 = n342 & n349;
  assign po0  = ~n346 | n350;
  assign n352 = ~pi74  & ~pi75 ;
  assign n353 = ~pi90  & ~pi91 ;
  assign n354 = n137 & ~n140;
  assign n355 = n138 & ~n143;
  assign n356 = ~n354 & n355;
  assign n357 = ~pi118  & ~pi119 ;
  assign n358 = ~pi116  & ~pi117 ;
  assign n359 = ~pi114  & ~pi115 ;
  assign n360 = n358 & ~n359;
  assign n361 = n357 & ~n360;
  assign n362 = n143 & n361;
  assign n363 = ~n356 & ~n362;
  assign n364 = ~pi112  & n359;
  assign n365 = n357 & n358;
  assign n366 = ~pi113  & n365;
  assign n367 = n364 & n366;
  assign n368 = n143 & n367;
  assign n369 = ~pi110  & ~pi111 ;
  assign n370 = ~pi106  & ~pi107 ;
  assign n371 = ~pi108  & ~pi109 ;
  assign n372 = ~n370 & n371;
  assign n373 = n369 & ~n372;
  assign n374 = n368 & ~n373;
  assign n375 = ~n363 & ~n374;
  assign n376 = ~pi102  & ~pi103 ;
  assign n377 = ~pi98  & ~pi99 ;
  assign n378 = n376 & n377;
  assign n379 = ~pi94  & ~pi95 ;
  assign n380 = n378 & n379;
  assign n381 = n375 & n380;
  assign n382 = n353 & n381;
  assign n383 = ~pi86  & ~pi87 ;
  assign n384 = n382 & n383;
  assign n385 = ~pi82  & ~pi83 ;
  assign n386 = n384 & n385;
  assign n387 = ~pi78  & n386;
  assign n388 = ~pi79  & n387;
  assign n389 = n352 & n388;
  assign n390 = ~pi70  & ~pi71 ;
  assign n391 = n389 & n390;
  assign n392 = ~pi66  & ~pi67 ;
  assign n393 = n391 & n392;
  assign n394 = ~pi62  & ~pi63 ;
  assign n395 = n393 & n394;
  assign n396 = ~pi58  & ~pi59 ;
  assign n397 = n395 & n396;
  assign n398 = ~pi54  & ~pi55 ;
  assign n399 = n397 & n398;
  assign n400 = ~pi50  & ~pi51 ;
  assign n401 = n399 & n400;
  assign n402 = ~pi46  & ~pi47 ;
  assign n403 = n401 & n402;
  assign n404 = ~pi42  & ~pi43 ;
  assign n405 = n403 & n404;
  assign n406 = ~pi38  & ~pi39 ;
  assign n407 = n405 & n406;
  assign n408 = ~pi34  & ~pi35 ;
  assign n409 = n407 & n408;
  assign n410 = ~pi30  & ~pi31 ;
  assign n411 = n409 & n410;
  assign n412 = ~pi26  & ~pi27 ;
  assign n413 = n411 & n412;
  assign n414 = ~pi22  & ~pi23 ;
  assign n415 = n413 & n414;
  assign n416 = ~pi18  & ~pi19 ;
  assign n417 = n415 & n416;
  assign n418 = ~pi14  & ~pi15 ;
  assign n419 = n417 & n418;
  assign n420 = ~pi100  & ~pi101 ;
  assign n421 = n369 & n371;
  assign n422 = n368 & n421;
  assign n423 = ~pi105  & n370;
  assign n424 = ~pi104  & n423;
  assign n425 = n422 & n424;
  assign n426 = n420 & n425;
  assign n427 = ~pi96  & ~pi97 ;
  assign n428 = n426 & n427;
  assign n429 = ~pi92  & ~pi93 ;
  assign n430 = n428 & n429;
  assign n431 = ~pi88  & ~pi89 ;
  assign n432 = n430 & n431;
  assign n433 = ~pi84  & ~pi85 ;
  assign n434 = n432 & n433;
  assign n435 = ~pi80  & ~pi81 ;
  assign n436 = n434 & n435;
  assign n437 = ~pi76  & ~pi77 ;
  assign n438 = n436 & n437;
  assign n439 = ~pi72  & ~pi73 ;
  assign n440 = n438 & n439;
  assign n441 = ~pi68  & ~pi69 ;
  assign n442 = n440 & n441;
  assign n443 = ~pi64  & ~pi65 ;
  assign n444 = n442 & n443;
  assign n445 = ~pi60  & ~pi61 ;
  assign n446 = n444 & n445;
  assign n447 = ~pi56  & ~pi57 ;
  assign n448 = n446 & n447;
  assign n449 = ~pi52  & ~pi53 ;
  assign n450 = n448 & n449;
  assign n451 = ~pi48  & ~pi49 ;
  assign n452 = n450 & n451;
  assign n453 = ~pi44  & ~pi45 ;
  assign n454 = n452 & n453;
  assign n455 = ~pi40  & ~pi41 ;
  assign n456 = n454 & n455;
  assign n457 = ~pi36  & ~pi37 ;
  assign n458 = n456 & n457;
  assign n459 = ~pi32  & ~pi33 ;
  assign n460 = n458 & n459;
  assign n461 = ~pi28  & ~pi29 ;
  assign n462 = n460 & n461;
  assign n463 = ~pi24  & ~pi25 ;
  assign n464 = n462 & n463;
  assign n465 = ~pi20  & ~pi21 ;
  assign n466 = n464 & n465;
  assign n467 = ~pi16  & ~pi17 ;
  assign n468 = n466 & n467;
  assign n469 = n376 & ~n420;
  assign n470 = ~n378 & ~n469;
  assign n471 = n425 & n470;
  assign n472 = ~n428 & ~n471;
  assign n473 = ~n380 & ~n472;
  assign n474 = ~n430 & ~n473;
  assign n475 = n375 & n474;
  assign n476 = ~n382 & ~n475;
  assign n477 = ~n432 & ~n476;
  assign n478 = ~n384 & ~n477;
  assign n479 = ~n434 & ~n478;
  assign n480 = ~n386 & ~n479;
  assign n481 = ~n436 & ~n480;
  assign n482 = ~n388 & ~n481;
  assign n483 = ~n438 & ~n482;
  assign n484 = ~n389 & ~n483;
  assign n485 = ~n440 & ~n484;
  assign n486 = ~n391 & ~n485;
  assign n487 = ~n442 & ~n486;
  assign n488 = ~n393 & ~n487;
  assign n489 = ~n444 & ~n488;
  assign n490 = ~n395 & ~n489;
  assign n491 = ~n446 & ~n490;
  assign n492 = ~n397 & ~n491;
  assign n493 = ~n448 & ~n492;
  assign n494 = ~n399 & ~n493;
  assign n495 = ~n450 & ~n494;
  assign n496 = ~n401 & ~n495;
  assign n497 = ~n452 & ~n496;
  assign n498 = ~n403 & ~n497;
  assign n499 = ~n454 & ~n498;
  assign n500 = ~n405 & ~n499;
  assign n501 = ~n456 & ~n500;
  assign n502 = ~n407 & ~n501;
  assign n503 = ~n458 & ~n502;
  assign n504 = ~n409 & ~n503;
  assign n505 = ~n460 & ~n504;
  assign n506 = ~n411 & ~n505;
  assign n507 = ~n462 & ~n506;
  assign n508 = ~n413 & ~n507;
  assign n509 = ~n464 & ~n508;
  assign n510 = ~n415 & ~n509;
  assign n511 = ~n466 & ~n510;
  assign n512 = ~n417 & ~n511;
  assign n513 = ~n468 & ~n512;
  assign n514 = ~n419 & ~n513;
  assign n515 = ~pi12  & ~pi13 ;
  assign n516 = ~pi10  & ~pi11 ;
  assign n517 = n419 & n516;
  assign n518 = ~pi8  & ~pi9 ;
  assign n519 = n517 & ~n518;
  assign n520 = n515 & ~n519;
  assign n521 = n468 & n520;
  assign n522 = ~n514 & ~n521;
  assign n523 = ~pi6  & ~pi7 ;
  assign n524 = ~pi4  & ~pi5 ;
  assign n525 = ~pi2  & ~pi3 ;
  assign n526 = n524 & ~n525;
  assign n527 = n517 & ~n526;
  assign n528 = n523 & n527;
  assign po1  = ~n522 & ~n528;
  assign n530 = n377 & n427;
  assign n531 = n376 & n426;
  assign n532 = ~n530 & n531;
  assign n533 = n352 & n439;
  assign n534 = n379 & n429;
  assign n535 = n531 & n534;
  assign n536 = n383 & n433;
  assign n537 = n535 & n536;
  assign n538 = n385 & n435;
  assign n539 = ~pi78  & n437;
  assign n540 = ~pi79  & n539;
  assign n541 = n538 & ~n540;
  assign n542 = n537 & ~n541;
  assign n543 = ~n533 & n542;
  assign n544 = n142 & ~n365;
  assign n545 = ~n368 & ~n544;
  assign n546 = n139 & n545;
  assign n547 = ~n422 & ~n546;
  assign n548 = ~n425 & ~n547;
  assign n549 = n353 & n431;
  assign n550 = n535 & ~n549;
  assign n551 = ~n548 & ~n550;
  assign n552 = ~n543 & n551;
  assign n553 = ~n532 & n552;
  assign n554 = n533 & ~n538;
  assign n555 = n537 & n554;
  assign n556 = n553 & ~n555;
  assign n557 = n390 & n441;
  assign n558 = n542 & n557;
  assign n559 = n394 & n445;
  assign n560 = n392 & n443;
  assign n561 = ~n559 & n560;
  assign n562 = n558 & ~n561;
  assign n563 = n556 & ~n562;
  assign n564 = n398 & n449;
  assign n565 = n558 & ~n560;
  assign n566 = n396 & n447;
  assign n567 = n556 & n566;
  assign n568 = ~n565 & n567;
  assign n569 = ~n564 & n568;
  assign n570 = n402 & n453;
  assign n571 = n400 & n451;
  assign n572 = n568 & n571;
  assign n573 = ~n570 & n572;
  assign n574 = ~n569 & ~n573;
  assign n575 = ~n563 & n574;
  assign n576 = n404 & n455;
  assign n577 = n572 & n576;
  assign n578 = n408 & n459;
  assign n579 = n406 & n457;
  assign n580 = ~n578 & n579;
  assign n581 = n577 & ~n580;
  assign n582 = n575 & ~n581;
  assign n583 = n577 & ~n579;
  assign n584 = n410 & n461;
  assign n585 = ~n583 & n584;
  assign n586 = n575 & n585;
  assign n587 = ~n582 & ~n586;
  assign n588 = n414 & n465;
  assign n589 = n412 & n463;
  assign n590 = ~n582 & n589;
  assign n591 = ~n588 & n590;
  assign n592 = ~n587 & ~n591;
  assign n593 = n416 & n467;
  assign n594 = n418 & n515;
  assign n595 = n516 & n518;
  assign n596 = n523 & n524;
  assign n597 = n595 & ~n596;
  assign n598 = n594 & ~n597;
  assign n599 = ~n587 & ~n590;
  assign n600 = ~n598 & ~n599;
  assign n601 = n593 & n600;
  assign po2  = ~n592 | n601;
  assign n603 = n421 & n424;
  assign n604 = ~pi102  & n530;
  assign n605 = n420 & n604;
  assign n606 = ~n603 & ~n605;
  assign n607 = n367 & n606;
  assign n608 = n143 & ~n607;
  assign n609 = pi103  & n603;
  assign n610 = n367 & ~n609;
  assign n611 = n605 & n610;
  assign n612 = n608 & ~n611;
  assign n613 = n536 & n538;
  assign n614 = n534 & n549;
  assign n615 = n425 & n614;
  assign n616 = ~n613 & n615;
  assign n617 = n564 & n571;
  assign n618 = n533 & n540;
  assign n619 = n615 & n618;
  assign n620 = n559 & n566;
  assign n621 = n557 & n560;
  assign n622 = ~n620 & n621;
  assign n623 = n619 & ~n622;
  assign n624 = ~n617 & n623;
  assign n625 = ~n616 & ~n624;
  assign n626 = ~n612 & n625;
  assign n627 = n617 & ~n621;
  assign n628 = n619 & n627;
  assign n629 = n626 & ~n628;
  assign n630 = n570 & n576;
  assign n631 = n623 & n630;
  assign n632 = n584 & n589;
  assign n633 = n588 & n593;
  assign n634 = n594 & n595;
  assign n635 = n633 & ~n634;
  assign n636 = n632 & ~n635;
  assign n637 = n578 & n579;
  assign n638 = ~n636 & n637;
  assign n639 = n631 & ~n638;
  assign po3  = n629 & ~n639;
  assign n641 = n613 & n614;
  assign n642 = n603 & n605;
  assign n643 = ~pi103  & n642;
  assign n644 = ~n641 & n643;
  assign n645 = n368 & ~n644;
  assign n646 = n617 & n620;
  assign n647 = n632 & n633;
  assign n648 = n630 & n637;
  assign n649 = ~n647 & n648;
  assign n650 = n646 & ~n649;
  assign n651 = n368 & n643;
  assign n652 = n618 & n621;
  assign n653 = n641 & n652;
  assign po6  = ~n651 | ~n653;
  assign n655 = ~n650 & ~po6 ;
  assign po4  = ~n645 | n655;
  assign n657 = n646 & n648;
  assign n658 = n653 & ~n657;
  assign po5  = ~n651 | n658;
  assign n660 = n596 & n647;
  assign n661 = ~pi1  & n660;
  assign n662 = n634 & n661;
  assign n663 = ~pi0  & n525;
  assign n664 = ~po6  & n663;
  assign n665 = n657 & n664;
  assign po7 = ~n662 | ~n665;
endmodule
