module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 , pi132 ,
    pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 , pi140 ,
    pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 , pi148 ,
    pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 , pi156 ,
    pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 , pi164 ,
    pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 , pi172 ,
    pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 , pi188 ,
    pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 , pi196 ,
    pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 , pi204 ,
    pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 , pi212 ,
    pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 , pi220 ,
    pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 ,
    po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 ,
    po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 , po30 , po31 , po32 ,
    po33 , po34 , po35 , po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 , po46 , po47 , po48 ,
    po49 , po50 , po51 , po52 , po53 , po54 , po55 , po56 ,
    po57 , po58 , po59 , po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 , po70 , po71 , po72 ,
    po73 , po74 , po75 , po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 , po86 , po87 , po88 ,
    po89 , po90 , po91 , po92 , po93 , po94 , po95 , po96 ,
    po97 , po98 , po99 , po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 , po116 , po117 ,
    po118 , po119 , po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127 , po128  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 ,
    pi140 , pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 ,
    pi148 , pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 ,
    pi156 , pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 ,
    pi164 , pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 ,
    pi172 , pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 ,
    pi180 , pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 ,
    pi196 , pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 ,
    pi204 , pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 ,
    pi212 , pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 ,
    pi220 , pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 , po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 , po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 , po101 , po102 ,
    po103 , po104 , po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 , po115 , po116 ,
    po117 , po118 , po119 , po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 , po128;
  wire n386, n387, n389, n390, n391, n392, n393,
    n395, n396, n397, n398, n399, n400, n401,
    n403, n404, n405, n406, n407, n408, n410,
    n411, n412, n413, n414, n415, n417, n418,
    n419, n420, n421, n422, n424, n425, n426,
    n427, n428, n429, n431, n432, n433, n434,
    n435, n436, n438, n439, n440, n441, n442,
    n443, n445, n446, n447, n448, n449, n450,
    n452, n453, n454, n455, n456, n457, n459,
    n460, n461, n462, n463, n464, n466, n467,
    n468, n469, n470, n471, n473, n474, n475,
    n476, n477, n478, n480, n481, n482, n483,
    n484, n485, n487, n488, n489, n490, n491,
    n492, n494, n495, n496, n497, n498, n499,
    n501, n502, n503, n504, n505, n506, n508,
    n509, n510, n511, n512, n513, n515, n516,
    n517, n518, n519, n520, n522, n523, n524,
    n525, n526, n527, n529, n530, n531, n532,
    n533, n534, n536, n537, n538, n539, n540,
    n541, n543, n544, n545, n546, n547, n548,
    n550, n551, n552, n553, n554, n555, n557,
    n558, n559, n560, n561, n562, n564, n565,
    n566, n567, n568, n569, n571, n572, n573,
    n574, n575, n576, n578, n579, n580, n581,
    n582, n583, n585, n586, n587, n588, n589,
    n590, n592, n593, n594, n595, n596, n597,
    n599, n600, n601, n602, n603, n604, n606,
    n607, n608, n609, n610, n611, n613, n614,
    n615, n616, n617, n618, n620, n621, n622,
    n623, n624, n625, n627, n628, n629, n630,
    n631, n632, n634, n635, n636, n637, n638,
    n639, n641, n642, n643, n644, n645, n646,
    n648, n649, n650, n651, n652, n653, n655,
    n656, n657, n658, n659, n660, n662, n663,
    n664, n665, n666, n667, n669, n670, n671,
    n672, n673, n674, n676, n677, n678, n679,
    n680, n681, n683, n684, n685, n686, n687,
    n688, n690, n691, n692, n693, n694, n695,
    n697, n698, n699, n700, n701, n702, n704,
    n705, n706, n707, n708, n709, n711, n712,
    n713, n714, n715, n716, n718, n719, n720,
    n721, n722, n723, n725, n726, n727, n728,
    n729, n730, n732, n733, n734, n735, n736,
    n737, n739, n740, n741, n742, n743, n744,
    n746, n747, n748, n749, n750, n751, n753,
    n754, n755, n756, n757, n758, n760, n761,
    n762, n763, n764, n765, n767, n768, n769,
    n770, n771, n772, n774, n775, n776, n777,
    n778, n779, n781, n782, n783, n784, n785,
    n786, n788, n789, n790, n791, n792, n793,
    n795, n796, n797, n798, n799, n800, n802,
    n803, n804, n805, n806, n807, n809, n810,
    n811, n812, n813, n814, n816, n817, n818,
    n819, n820, n821, n823, n824, n825, n826,
    n827, n828, n830, n831, n832, n833, n834,
    n835, n837, n838, n839, n840, n841, n842,
    n844, n845, n846, n847, n848, n849, n851,
    n852, n853, n854, n855, n856, n858, n859,
    n860, n861, n862, n863, n865, n866, n867,
    n868, n869, n870, n872, n873, n874, n875,
    n876, n877, n879, n880, n881, n882, n883,
    n884, n886, n887, n888, n889, n890, n891,
    n893, n894, n895, n896, n897, n898, n900,
    n901, n902, n903, n904, n905, n907, n908,
    n909, n910, n911, n912, n914, n915, n916,
    n917, n918, n919, n921, n922, n923, n924,
    n925, n926, n928, n929, n930, n931, n932,
    n933, n935, n936, n937, n938, n939, n940,
    n942, n943, n944, n945, n946, n947, n949,
    n950, n951, n952, n953, n954, n956, n957,
    n958, n959, n960, n961, n963, n964, n965,
    n966, n967, n968, n970, n971, n972, n973,
    n974, n975, n977, n978, n979, n980, n981,
    n982, n984, n985, n986, n987, n988, n989,
    n991, n992, n993, n994, n995, n996, n998,
    n999, n1000, n1001, n1002, n1003, n1005,
    n1006, n1007, n1008, n1009, n1010, n1012,
    n1013, n1014, n1015, n1016, n1017, n1019,
    n1020, n1021, n1022, n1023, n1024, n1026,
    n1027, n1028, n1029, n1030, n1031, n1033,
    n1034, n1035, n1036, n1037, n1038, n1040,
    n1041, n1042, n1043, n1044, n1045, n1047,
    n1048, n1049, n1050, n1051, n1052, n1054,
    n1055, n1056, n1057, n1058, n1059, n1061,
    n1062, n1063, n1064, n1065, n1066, n1068,
    n1069, n1070, n1071, n1072, n1073, n1075,
    n1076, n1077, n1078, n1079, n1080, n1082,
    n1083, n1084, n1085, n1086, n1087, n1089,
    n1090, n1091, n1092, n1093, n1094, n1096,
    n1097, n1098, n1099, n1100, n1101, n1103,
    n1104, n1105, n1106, n1107, n1108, n1110,
    n1111, n1112, n1113, n1114, n1115, n1117,
    n1118, n1119, n1120, n1121, n1122, n1124,
    n1125, n1126, n1127, n1128, n1129, n1131,
    n1132, n1133, n1134, n1135, n1136, n1138,
    n1139, n1140, n1141, n1142, n1143, n1145,
    n1146, n1147, n1148, n1149, n1150, n1152,
    n1153, n1154, n1155, n1156, n1157, n1159,
    n1160, n1161, n1162, n1163, n1164, n1166,
    n1167, n1168, n1169, n1170, n1171, n1173,
    n1174, n1175, n1176, n1177, n1178, n1180,
    n1181, n1182, n1183, n1184, n1185, n1187,
    n1188, n1189, n1190, n1191, n1192, n1194,
    n1195, n1196, n1197, n1198, n1199, n1201,
    n1202, n1203, n1204, n1205, n1206, n1208,
    n1209, n1210, n1211, n1212, n1213, n1215,
    n1216, n1217, n1218, n1219, n1220, n1222,
    n1223, n1224, n1225, n1226, n1227, n1229,
    n1230, n1231, n1232, n1233, n1234, n1236,
    n1237, n1238, n1239, n1240, n1241, n1243,
    n1244, n1245, n1246, n1247, n1248, n1250,
    n1251, n1252, n1253, n1254, n1255, n1257,
    n1258, n1259, n1260, n1261, n1262, n1264,
    n1265, n1266, n1267, n1268, n1269, n1271,
    n1272, n1273, n1274, n1275, n1276;
  assign n386 = pi0  & pi128 ;
  assign n387 = ~pi0  & ~pi128 ;
  assign po0  = ~n386 & ~n387;
  assign n389 = ~pi1  & ~pi129 ;
  assign n390 = pi1  & pi129 ;
  assign n391 = ~n389 & ~n390;
  assign n392 = n386 & ~n391;
  assign n393 = ~n386 & n391;
  assign po1  = n392 | n393;
  assign n395 = ~pi2  & ~pi130 ;
  assign n396 = pi2  & pi130 ;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~n386 & ~n390;
  assign n399 = ~n389 & ~n398;
  assign n400 = ~n397 & ~n399;
  assign n401 = n397 & n399;
  assign po2  = ~n400 & ~n401;
  assign n403 = ~pi3  & ~pi131 ;
  assign n404 = pi3  & pi131 ;
  assign n405 = ~n403 & ~n404;
  assign n406 = ~n396 & ~n401;
  assign n407 = ~n405 & n406;
  assign n408 = n405 & ~n406;
  assign po3  = ~n407 & ~n408;
  assign n410 = ~pi4  & ~pi132 ;
  assign n411 = pi4  & pi132 ;
  assign n412 = ~n410 & ~n411;
  assign n413 = ~n404 & ~n408;
  assign n414 = ~n412 & n413;
  assign n415 = n412 & ~n413;
  assign po4  = ~n414 & ~n415;
  assign n417 = ~pi5  & ~pi133 ;
  assign n418 = pi5  & pi133 ;
  assign n419 = ~n417 & ~n418;
  assign n420 = ~n411 & ~n415;
  assign n421 = ~n419 & n420;
  assign n422 = n419 & ~n420;
  assign po5  = ~n421 & ~n422;
  assign n424 = ~pi6  & ~pi134 ;
  assign n425 = pi6  & pi134 ;
  assign n426 = ~n424 & ~n425;
  assign n427 = ~n418 & ~n422;
  assign n428 = ~n426 & n427;
  assign n429 = n426 & ~n427;
  assign po6  = ~n428 & ~n429;
  assign n431 = ~pi7  & ~pi135 ;
  assign n432 = pi7  & pi135 ;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~n425 & ~n429;
  assign n435 = ~n433 & n434;
  assign n436 = n433 & ~n434;
  assign po7  = ~n435 & ~n436;
  assign n438 = ~pi8  & ~pi136 ;
  assign n439 = pi8  & pi136 ;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~n432 & ~n436;
  assign n442 = ~n440 & n441;
  assign n443 = n440 & ~n441;
  assign po8  = ~n442 & ~n443;
  assign n445 = ~pi9  & ~pi137 ;
  assign n446 = pi9  & pi137 ;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~n439 & ~n443;
  assign n449 = ~n447 & n448;
  assign n450 = n447 & ~n448;
  assign po9  = ~n449 & ~n450;
  assign n452 = ~pi10  & ~pi138 ;
  assign n453 = pi10  & pi138 ;
  assign n454 = ~n452 & ~n453;
  assign n455 = ~n446 & ~n450;
  assign n456 = ~n454 & n455;
  assign n457 = n454 & ~n455;
  assign po10  = ~n456 & ~n457;
  assign n459 = ~pi11  & ~pi139 ;
  assign n460 = pi11  & pi139 ;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n453 & ~n457;
  assign n463 = ~n461 & n462;
  assign n464 = n461 & ~n462;
  assign po11  = ~n463 & ~n464;
  assign n466 = ~pi12  & ~pi140 ;
  assign n467 = pi12  & pi140 ;
  assign n468 = ~n466 & ~n467;
  assign n469 = ~n460 & ~n464;
  assign n470 = ~n468 & n469;
  assign n471 = n468 & ~n469;
  assign po12  = ~n470 & ~n471;
  assign n473 = ~pi13  & ~pi141 ;
  assign n474 = pi13  & pi141 ;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~n467 & ~n471;
  assign n477 = ~n475 & n476;
  assign n478 = n475 & ~n476;
  assign po13  = ~n477 & ~n478;
  assign n480 = ~pi14  & ~pi142 ;
  assign n481 = pi14  & pi142 ;
  assign n482 = ~n480 & ~n481;
  assign n483 = ~n474 & ~n478;
  assign n484 = ~n482 & n483;
  assign n485 = n482 & ~n483;
  assign po14  = ~n484 & ~n485;
  assign n487 = ~pi15  & ~pi143 ;
  assign n488 = pi15  & pi143 ;
  assign n489 = ~n487 & ~n488;
  assign n490 = ~n481 & ~n485;
  assign n491 = ~n489 & n490;
  assign n492 = n489 & ~n490;
  assign po15  = ~n491 & ~n492;
  assign n494 = ~pi16  & ~pi144 ;
  assign n495 = pi16  & pi144 ;
  assign n496 = ~n494 & ~n495;
  assign n497 = ~n488 & ~n492;
  assign n498 = ~n496 & n497;
  assign n499 = n496 & ~n497;
  assign po16  = ~n498 & ~n499;
  assign n501 = ~pi17  & ~pi145 ;
  assign n502 = pi17  & pi145 ;
  assign n503 = ~n501 & ~n502;
  assign n504 = ~n495 & ~n499;
  assign n505 = ~n503 & n504;
  assign n506 = n503 & ~n504;
  assign po17  = ~n505 & ~n506;
  assign n508 = ~pi18  & ~pi146 ;
  assign n509 = pi18  & pi146 ;
  assign n510 = ~n508 & ~n509;
  assign n511 = ~n502 & ~n506;
  assign n512 = ~n510 & n511;
  assign n513 = n510 & ~n511;
  assign po18  = ~n512 & ~n513;
  assign n515 = ~pi19  & ~pi147 ;
  assign n516 = pi19  & pi147 ;
  assign n517 = ~n515 & ~n516;
  assign n518 = ~n509 & ~n513;
  assign n519 = ~n517 & n518;
  assign n520 = n517 & ~n518;
  assign po19  = ~n519 & ~n520;
  assign n522 = ~pi20  & ~pi148 ;
  assign n523 = pi20  & pi148 ;
  assign n524 = ~n522 & ~n523;
  assign n525 = ~n516 & ~n520;
  assign n526 = ~n524 & n525;
  assign n527 = n524 & ~n525;
  assign po20  = ~n526 & ~n527;
  assign n529 = ~pi21  & ~pi149 ;
  assign n530 = pi21  & pi149 ;
  assign n531 = ~n529 & ~n530;
  assign n532 = ~n523 & ~n527;
  assign n533 = ~n531 & n532;
  assign n534 = n531 & ~n532;
  assign po21  = ~n533 & ~n534;
  assign n536 = ~pi22  & ~pi150 ;
  assign n537 = pi22  & pi150 ;
  assign n538 = ~n536 & ~n537;
  assign n539 = ~n530 & ~n534;
  assign n540 = ~n538 & n539;
  assign n541 = n538 & ~n539;
  assign po22  = ~n540 & ~n541;
  assign n543 = ~pi23  & ~pi151 ;
  assign n544 = pi23  & pi151 ;
  assign n545 = ~n543 & ~n544;
  assign n546 = ~n537 & ~n541;
  assign n547 = ~n545 & n546;
  assign n548 = n545 & ~n546;
  assign po23  = ~n547 & ~n548;
  assign n550 = ~pi24  & ~pi152 ;
  assign n551 = pi24  & pi152 ;
  assign n552 = ~n550 & ~n551;
  assign n553 = ~n544 & ~n548;
  assign n554 = ~n552 & n553;
  assign n555 = n552 & ~n553;
  assign po24  = ~n554 & ~n555;
  assign n557 = ~pi25  & ~pi153 ;
  assign n558 = pi25  & pi153 ;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~n551 & ~n555;
  assign n561 = ~n559 & n560;
  assign n562 = n559 & ~n560;
  assign po25  = ~n561 & ~n562;
  assign n564 = ~pi26  & ~pi154 ;
  assign n565 = pi26  & pi154 ;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~n558 & ~n562;
  assign n568 = ~n566 & n567;
  assign n569 = n566 & ~n567;
  assign po26  = ~n568 & ~n569;
  assign n571 = ~pi27  & ~pi155 ;
  assign n572 = pi27  & pi155 ;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~n565 & ~n569;
  assign n575 = ~n573 & n574;
  assign n576 = n573 & ~n574;
  assign po27  = ~n575 & ~n576;
  assign n578 = ~pi28  & ~pi156 ;
  assign n579 = pi28  & pi156 ;
  assign n580 = ~n578 & ~n579;
  assign n581 = ~n572 & ~n576;
  assign n582 = ~n580 & n581;
  assign n583 = n580 & ~n581;
  assign po28  = ~n582 & ~n583;
  assign n585 = ~pi29  & ~pi157 ;
  assign n586 = pi29  & pi157 ;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~n579 & ~n583;
  assign n589 = ~n587 & n588;
  assign n590 = n587 & ~n588;
  assign po29  = ~n589 & ~n590;
  assign n592 = ~pi30  & ~pi158 ;
  assign n593 = pi30  & pi158 ;
  assign n594 = ~n592 & ~n593;
  assign n595 = ~n586 & ~n590;
  assign n596 = ~n594 & n595;
  assign n597 = n594 & ~n595;
  assign po30  = ~n596 & ~n597;
  assign n599 = ~pi31  & ~pi159 ;
  assign n600 = pi31  & pi159 ;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n593 & ~n597;
  assign n603 = ~n601 & n602;
  assign n604 = n601 & ~n602;
  assign po31  = ~n603 & ~n604;
  assign n606 = ~pi32  & ~pi160 ;
  assign n607 = pi32  & pi160 ;
  assign n608 = ~n606 & ~n607;
  assign n609 = ~n600 & ~n604;
  assign n610 = ~n608 & n609;
  assign n611 = n608 & ~n609;
  assign po32  = ~n610 & ~n611;
  assign n613 = ~pi33  & ~pi161 ;
  assign n614 = pi33  & pi161 ;
  assign n615 = ~n613 & ~n614;
  assign n616 = ~n607 & ~n611;
  assign n617 = ~n615 & n616;
  assign n618 = n615 & ~n616;
  assign po33  = ~n617 & ~n618;
  assign n620 = ~pi34  & ~pi162 ;
  assign n621 = pi34  & pi162 ;
  assign n622 = ~n620 & ~n621;
  assign n623 = ~n614 & ~n618;
  assign n624 = ~n622 & n623;
  assign n625 = n622 & ~n623;
  assign po34  = ~n624 & ~n625;
  assign n627 = ~pi35  & ~pi163 ;
  assign n628 = pi35  & pi163 ;
  assign n629 = ~n627 & ~n628;
  assign n630 = ~n621 & ~n625;
  assign n631 = ~n629 & n630;
  assign n632 = n629 & ~n630;
  assign po35  = ~n631 & ~n632;
  assign n634 = ~pi36  & ~pi164 ;
  assign n635 = pi36  & pi164 ;
  assign n636 = ~n634 & ~n635;
  assign n637 = ~n628 & ~n632;
  assign n638 = ~n636 & n637;
  assign n639 = n636 & ~n637;
  assign po36  = ~n638 & ~n639;
  assign n641 = ~pi37  & ~pi165 ;
  assign n642 = pi37  & pi165 ;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~n635 & ~n639;
  assign n645 = ~n643 & n644;
  assign n646 = n643 & ~n644;
  assign po37  = ~n645 & ~n646;
  assign n648 = ~pi38  & ~pi166 ;
  assign n649 = pi38  & pi166 ;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~n642 & ~n646;
  assign n652 = ~n650 & n651;
  assign n653 = n650 & ~n651;
  assign po38  = ~n652 & ~n653;
  assign n655 = ~pi39  & ~pi167 ;
  assign n656 = pi39  & pi167 ;
  assign n657 = ~n655 & ~n656;
  assign n658 = ~n649 & ~n653;
  assign n659 = ~n657 & n658;
  assign n660 = n657 & ~n658;
  assign po39  = ~n659 & ~n660;
  assign n662 = ~pi40  & ~pi168 ;
  assign n663 = pi40  & pi168 ;
  assign n664 = ~n662 & ~n663;
  assign n665 = ~n656 & ~n660;
  assign n666 = ~n664 & n665;
  assign n667 = n664 & ~n665;
  assign po40  = ~n666 & ~n667;
  assign n669 = ~pi41  & ~pi169 ;
  assign n670 = pi41  & pi169 ;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~n663 & ~n667;
  assign n673 = ~n671 & n672;
  assign n674 = n671 & ~n672;
  assign po41  = ~n673 & ~n674;
  assign n676 = ~pi42  & ~pi170 ;
  assign n677 = pi42  & pi170 ;
  assign n678 = ~n676 & ~n677;
  assign n679 = ~n670 & ~n674;
  assign n680 = ~n678 & n679;
  assign n681 = n678 & ~n679;
  assign po42  = ~n680 & ~n681;
  assign n683 = ~pi43  & ~pi171 ;
  assign n684 = pi43  & pi171 ;
  assign n685 = ~n683 & ~n684;
  assign n686 = ~n677 & ~n681;
  assign n687 = ~n685 & n686;
  assign n688 = n685 & ~n686;
  assign po43  = ~n687 & ~n688;
  assign n690 = ~pi44  & ~pi172 ;
  assign n691 = pi44  & pi172 ;
  assign n692 = ~n690 & ~n691;
  assign n693 = ~n684 & ~n688;
  assign n694 = ~n692 & n693;
  assign n695 = n692 & ~n693;
  assign po44  = ~n694 & ~n695;
  assign n697 = ~pi45  & ~pi173 ;
  assign n698 = pi45  & pi173 ;
  assign n699 = ~n697 & ~n698;
  assign n700 = ~n691 & ~n695;
  assign n701 = ~n699 & n700;
  assign n702 = n699 & ~n700;
  assign po45  = ~n701 & ~n702;
  assign n704 = ~pi46  & ~pi174 ;
  assign n705 = pi46  & pi174 ;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n698 & ~n702;
  assign n708 = ~n706 & n707;
  assign n709 = n706 & ~n707;
  assign po46  = ~n708 & ~n709;
  assign n711 = ~pi47  & ~pi175 ;
  assign n712 = pi47  & pi175 ;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n705 & ~n709;
  assign n715 = ~n713 & n714;
  assign n716 = n713 & ~n714;
  assign po47  = ~n715 & ~n716;
  assign n718 = ~pi48  & ~pi176 ;
  assign n719 = pi48  & pi176 ;
  assign n720 = ~n718 & ~n719;
  assign n721 = ~n712 & ~n716;
  assign n722 = ~n720 & n721;
  assign n723 = n720 & ~n721;
  assign po48  = ~n722 & ~n723;
  assign n725 = ~pi49  & ~pi177 ;
  assign n726 = pi49  & pi177 ;
  assign n727 = ~n725 & ~n726;
  assign n728 = ~n719 & ~n723;
  assign n729 = ~n727 & n728;
  assign n730 = n727 & ~n728;
  assign po49  = ~n729 & ~n730;
  assign n732 = ~pi50  & ~pi178 ;
  assign n733 = pi50  & pi178 ;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n726 & ~n730;
  assign n736 = ~n734 & n735;
  assign n737 = n734 & ~n735;
  assign po50  = ~n736 & ~n737;
  assign n739 = ~pi51  & ~pi179 ;
  assign n740 = pi51  & pi179 ;
  assign n741 = ~n739 & ~n740;
  assign n742 = ~n733 & ~n737;
  assign n743 = ~n741 & n742;
  assign n744 = n741 & ~n742;
  assign po51  = ~n743 & ~n744;
  assign n746 = ~pi52  & ~pi180 ;
  assign n747 = pi52  & pi180 ;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~n740 & ~n744;
  assign n750 = ~n748 & n749;
  assign n751 = n748 & ~n749;
  assign po52  = ~n750 & ~n751;
  assign n753 = ~pi53  & ~pi181 ;
  assign n754 = pi53  & pi181 ;
  assign n755 = ~n753 & ~n754;
  assign n756 = ~n747 & ~n751;
  assign n757 = ~n755 & n756;
  assign n758 = n755 & ~n756;
  assign po53  = ~n757 & ~n758;
  assign n760 = ~pi54  & ~pi182 ;
  assign n761 = pi54  & pi182 ;
  assign n762 = ~n760 & ~n761;
  assign n763 = ~n754 & ~n758;
  assign n764 = ~n762 & n763;
  assign n765 = n762 & ~n763;
  assign po54  = ~n764 & ~n765;
  assign n767 = ~pi55  & ~pi183 ;
  assign n768 = pi55  & pi183 ;
  assign n769 = ~n767 & ~n768;
  assign n770 = ~n761 & ~n765;
  assign n771 = ~n769 & n770;
  assign n772 = n769 & ~n770;
  assign po55  = ~n771 & ~n772;
  assign n774 = ~pi56  & ~pi184 ;
  assign n775 = pi56  & pi184 ;
  assign n776 = ~n774 & ~n775;
  assign n777 = ~n768 & ~n772;
  assign n778 = ~n776 & n777;
  assign n779 = n776 & ~n777;
  assign po56  = ~n778 & ~n779;
  assign n781 = ~pi57  & ~pi185 ;
  assign n782 = pi57  & pi185 ;
  assign n783 = ~n781 & ~n782;
  assign n784 = ~n775 & ~n779;
  assign n785 = ~n783 & n784;
  assign n786 = n783 & ~n784;
  assign po57  = ~n785 & ~n786;
  assign n788 = ~pi58  & ~pi186 ;
  assign n789 = pi58  & pi186 ;
  assign n790 = ~n788 & ~n789;
  assign n791 = ~n782 & ~n786;
  assign n792 = ~n790 & n791;
  assign n793 = n790 & ~n791;
  assign po58  = ~n792 & ~n793;
  assign n795 = ~pi59  & ~pi187 ;
  assign n796 = pi59  & pi187 ;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~n789 & ~n793;
  assign n799 = ~n797 & n798;
  assign n800 = n797 & ~n798;
  assign po59  = ~n799 & ~n800;
  assign n802 = ~pi60  & ~pi188 ;
  assign n803 = pi60  & pi188 ;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~n796 & ~n800;
  assign n806 = ~n804 & n805;
  assign n807 = n804 & ~n805;
  assign po60  = ~n806 & ~n807;
  assign n809 = ~pi61  & ~pi189 ;
  assign n810 = pi61  & pi189 ;
  assign n811 = ~n809 & ~n810;
  assign n812 = ~n803 & ~n807;
  assign n813 = ~n811 & n812;
  assign n814 = n811 & ~n812;
  assign po61  = ~n813 & ~n814;
  assign n816 = ~pi62  & ~pi190 ;
  assign n817 = pi62  & pi190 ;
  assign n818 = ~n816 & ~n817;
  assign n819 = ~n810 & ~n814;
  assign n820 = ~n818 & n819;
  assign n821 = n818 & ~n819;
  assign po62  = ~n820 & ~n821;
  assign n823 = ~pi63  & ~pi191 ;
  assign n824 = pi63  & pi191 ;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~n817 & ~n821;
  assign n827 = ~n825 & n826;
  assign n828 = n825 & ~n826;
  assign po63  = ~n827 & ~n828;
  assign n830 = ~pi64  & ~pi192 ;
  assign n831 = pi64  & pi192 ;
  assign n832 = ~n830 & ~n831;
  assign n833 = ~n824 & ~n828;
  assign n834 = ~n832 & n833;
  assign n835 = n832 & ~n833;
  assign po64  = ~n834 & ~n835;
  assign n837 = ~pi65  & ~pi193 ;
  assign n838 = pi65  & pi193 ;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~n831 & ~n835;
  assign n841 = ~n839 & n840;
  assign n842 = n839 & ~n840;
  assign po65  = ~n841 & ~n842;
  assign n844 = ~pi66  & ~pi194 ;
  assign n845 = pi66  & pi194 ;
  assign n846 = ~n844 & ~n845;
  assign n847 = ~n838 & ~n842;
  assign n848 = ~n846 & n847;
  assign n849 = n846 & ~n847;
  assign po66  = ~n848 & ~n849;
  assign n851 = ~pi67  & ~pi195 ;
  assign n852 = pi67  & pi195 ;
  assign n853 = ~n851 & ~n852;
  assign n854 = ~n845 & ~n849;
  assign n855 = ~n853 & n854;
  assign n856 = n853 & ~n854;
  assign po67  = ~n855 & ~n856;
  assign n858 = ~pi68  & ~pi196 ;
  assign n859 = pi68  & pi196 ;
  assign n860 = ~n858 & ~n859;
  assign n861 = ~n852 & ~n856;
  assign n862 = ~n860 & n861;
  assign n863 = n860 & ~n861;
  assign po68  = ~n862 & ~n863;
  assign n865 = ~pi69  & ~pi197 ;
  assign n866 = pi69  & pi197 ;
  assign n867 = ~n865 & ~n866;
  assign n868 = ~n859 & ~n863;
  assign n869 = ~n867 & n868;
  assign n870 = n867 & ~n868;
  assign po69  = ~n869 & ~n870;
  assign n872 = ~pi70  & ~pi198 ;
  assign n873 = pi70  & pi198 ;
  assign n874 = ~n872 & ~n873;
  assign n875 = ~n866 & ~n870;
  assign n876 = ~n874 & n875;
  assign n877 = n874 & ~n875;
  assign po70  = ~n876 & ~n877;
  assign n879 = ~pi71  & ~pi199 ;
  assign n880 = pi71  & pi199 ;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n873 & ~n877;
  assign n883 = ~n881 & n882;
  assign n884 = n881 & ~n882;
  assign po71  = ~n883 & ~n884;
  assign n886 = ~pi72  & ~pi200 ;
  assign n887 = pi72  & pi200 ;
  assign n888 = ~n886 & ~n887;
  assign n889 = ~n880 & ~n884;
  assign n890 = ~n888 & n889;
  assign n891 = n888 & ~n889;
  assign po72  = ~n890 & ~n891;
  assign n893 = ~pi73  & ~pi201 ;
  assign n894 = pi73  & pi201 ;
  assign n895 = ~n893 & ~n894;
  assign n896 = ~n887 & ~n891;
  assign n897 = ~n895 & n896;
  assign n898 = n895 & ~n896;
  assign po73  = ~n897 & ~n898;
  assign n900 = ~pi74  & ~pi202 ;
  assign n901 = pi74  & pi202 ;
  assign n902 = ~n900 & ~n901;
  assign n903 = ~n894 & ~n898;
  assign n904 = ~n902 & n903;
  assign n905 = n902 & ~n903;
  assign po74  = ~n904 & ~n905;
  assign n907 = ~pi75  & ~pi203 ;
  assign n908 = pi75  & pi203 ;
  assign n909 = ~n907 & ~n908;
  assign n910 = ~n901 & ~n905;
  assign n911 = ~n909 & n910;
  assign n912 = n909 & ~n910;
  assign po75  = ~n911 & ~n912;
  assign n914 = ~pi76  & ~pi204 ;
  assign n915 = pi76  & pi204 ;
  assign n916 = ~n914 & ~n915;
  assign n917 = ~n908 & ~n912;
  assign n918 = ~n916 & n917;
  assign n919 = n916 & ~n917;
  assign po76  = ~n918 & ~n919;
  assign n921 = ~pi77  & ~pi205 ;
  assign n922 = pi77  & pi205 ;
  assign n923 = ~n921 & ~n922;
  assign n924 = ~n915 & ~n919;
  assign n925 = ~n923 & n924;
  assign n926 = n923 & ~n924;
  assign po77  = ~n925 & ~n926;
  assign n928 = ~pi78  & ~pi206 ;
  assign n929 = pi78  & pi206 ;
  assign n930 = ~n928 & ~n929;
  assign n931 = ~n922 & ~n926;
  assign n932 = ~n930 & n931;
  assign n933 = n930 & ~n931;
  assign po78  = ~n932 & ~n933;
  assign n935 = ~pi79  & ~pi207 ;
  assign n936 = pi79  & pi207 ;
  assign n937 = ~n935 & ~n936;
  assign n938 = ~n929 & ~n933;
  assign n939 = ~n937 & n938;
  assign n940 = n937 & ~n938;
  assign po79  = ~n939 & ~n940;
  assign n942 = ~pi80  & ~pi208 ;
  assign n943 = pi80  & pi208 ;
  assign n944 = ~n942 & ~n943;
  assign n945 = ~n936 & ~n940;
  assign n946 = ~n944 & n945;
  assign n947 = n944 & ~n945;
  assign po80  = ~n946 & ~n947;
  assign n949 = ~pi81  & ~pi209 ;
  assign n950 = pi81  & pi209 ;
  assign n951 = ~n949 & ~n950;
  assign n952 = ~n943 & ~n947;
  assign n953 = ~n951 & n952;
  assign n954 = n951 & ~n952;
  assign po81  = ~n953 & ~n954;
  assign n956 = ~pi82  & ~pi210 ;
  assign n957 = pi82  & pi210 ;
  assign n958 = ~n956 & ~n957;
  assign n959 = ~n950 & ~n954;
  assign n960 = ~n958 & n959;
  assign n961 = n958 & ~n959;
  assign po82  = ~n960 & ~n961;
  assign n963 = ~pi83  & ~pi211 ;
  assign n964 = pi83  & pi211 ;
  assign n965 = ~n963 & ~n964;
  assign n966 = ~n957 & ~n961;
  assign n967 = ~n965 & n966;
  assign n968 = n965 & ~n966;
  assign po83  = ~n967 & ~n968;
  assign n970 = ~pi84  & ~pi212 ;
  assign n971 = pi84  & pi212 ;
  assign n972 = ~n970 & ~n971;
  assign n973 = ~n964 & ~n968;
  assign n974 = ~n972 & n973;
  assign n975 = n972 & ~n973;
  assign po84  = ~n974 & ~n975;
  assign n977 = ~pi85  & ~pi213 ;
  assign n978 = pi85  & pi213 ;
  assign n979 = ~n977 & ~n978;
  assign n980 = ~n971 & ~n975;
  assign n981 = ~n979 & n980;
  assign n982 = n979 & ~n980;
  assign po85  = ~n981 & ~n982;
  assign n984 = ~pi86  & ~pi214 ;
  assign n985 = pi86  & pi214 ;
  assign n986 = ~n984 & ~n985;
  assign n987 = ~n978 & ~n982;
  assign n988 = ~n986 & n987;
  assign n989 = n986 & ~n987;
  assign po86  = ~n988 & ~n989;
  assign n991 = ~pi87  & ~pi215 ;
  assign n992 = pi87  & pi215 ;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~n985 & ~n989;
  assign n995 = ~n993 & n994;
  assign n996 = n993 & ~n994;
  assign po87  = ~n995 & ~n996;
  assign n998 = ~pi88  & ~pi216 ;
  assign n999 = pi88  & pi216 ;
  assign n1000 = ~n998 & ~n999;
  assign n1001 = ~n992 & ~n996;
  assign n1002 = ~n1000 & n1001;
  assign n1003 = n1000 & ~n1001;
  assign po88  = ~n1002 & ~n1003;
  assign n1005 = ~pi89  & ~pi217 ;
  assign n1006 = pi89  & pi217 ;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = ~n999 & ~n1003;
  assign n1009 = ~n1007 & n1008;
  assign n1010 = n1007 & ~n1008;
  assign po89  = ~n1009 & ~n1010;
  assign n1012 = ~pi90  & ~pi218 ;
  assign n1013 = pi90  & pi218 ;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = ~n1006 & ~n1010;
  assign n1016 = ~n1014 & n1015;
  assign n1017 = n1014 & ~n1015;
  assign po90  = ~n1016 & ~n1017;
  assign n1019 = ~pi91  & ~pi219 ;
  assign n1020 = pi91  & pi219 ;
  assign n1021 = ~n1019 & ~n1020;
  assign n1022 = ~n1013 & ~n1017;
  assign n1023 = ~n1021 & n1022;
  assign n1024 = n1021 & ~n1022;
  assign po91  = ~n1023 & ~n1024;
  assign n1026 = ~pi92  & ~pi220 ;
  assign n1027 = pi92  & pi220 ;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = ~n1020 & ~n1024;
  assign n1030 = ~n1028 & n1029;
  assign n1031 = n1028 & ~n1029;
  assign po92  = ~n1030 & ~n1031;
  assign n1033 = ~pi93  & ~pi221 ;
  assign n1034 = pi93  & pi221 ;
  assign n1035 = ~n1033 & ~n1034;
  assign n1036 = ~n1027 & ~n1031;
  assign n1037 = ~n1035 & n1036;
  assign n1038 = n1035 & ~n1036;
  assign po93  = ~n1037 & ~n1038;
  assign n1040 = ~pi94  & ~pi222 ;
  assign n1041 = pi94  & pi222 ;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = ~n1034 & ~n1038;
  assign n1044 = ~n1042 & n1043;
  assign n1045 = n1042 & ~n1043;
  assign po94  = ~n1044 & ~n1045;
  assign n1047 = ~pi95  & ~pi223 ;
  assign n1048 = pi95  & pi223 ;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = ~n1041 & ~n1045;
  assign n1051 = ~n1049 & n1050;
  assign n1052 = n1049 & ~n1050;
  assign po95  = ~n1051 & ~n1052;
  assign n1054 = ~pi96  & ~pi224 ;
  assign n1055 = pi96  & pi224 ;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = ~n1048 & ~n1052;
  assign n1058 = ~n1056 & n1057;
  assign n1059 = n1056 & ~n1057;
  assign po96  = ~n1058 & ~n1059;
  assign n1061 = ~pi97  & ~pi225 ;
  assign n1062 = pi97  & pi225 ;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = ~n1055 & ~n1059;
  assign n1065 = ~n1063 & n1064;
  assign n1066 = n1063 & ~n1064;
  assign po97  = ~n1065 & ~n1066;
  assign n1068 = ~pi98  & ~pi226 ;
  assign n1069 = pi98  & pi226 ;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = ~n1062 & ~n1066;
  assign n1072 = ~n1070 & n1071;
  assign n1073 = n1070 & ~n1071;
  assign po98  = ~n1072 & ~n1073;
  assign n1075 = ~pi99  & ~pi227 ;
  assign n1076 = pi99  & pi227 ;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~n1069 & ~n1073;
  assign n1079 = ~n1077 & n1078;
  assign n1080 = n1077 & ~n1078;
  assign po99  = ~n1079 & ~n1080;
  assign n1082 = ~pi100  & ~pi228 ;
  assign n1083 = pi100  & pi228 ;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = ~n1076 & ~n1080;
  assign n1086 = ~n1084 & n1085;
  assign n1087 = n1084 & ~n1085;
  assign po100  = ~n1086 & ~n1087;
  assign n1089 = ~pi101  & ~pi229 ;
  assign n1090 = pi101  & pi229 ;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = ~n1083 & ~n1087;
  assign n1093 = ~n1091 & n1092;
  assign n1094 = n1091 & ~n1092;
  assign po101  = ~n1093 & ~n1094;
  assign n1096 = ~pi102  & ~pi230 ;
  assign n1097 = pi102  & pi230 ;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~n1090 & ~n1094;
  assign n1100 = ~n1098 & n1099;
  assign n1101 = n1098 & ~n1099;
  assign po102  = ~n1100 & ~n1101;
  assign n1103 = ~pi103  & ~pi231 ;
  assign n1104 = pi103  & pi231 ;
  assign n1105 = ~n1103 & ~n1104;
  assign n1106 = ~n1097 & ~n1101;
  assign n1107 = ~n1105 & n1106;
  assign n1108 = n1105 & ~n1106;
  assign po103  = ~n1107 & ~n1108;
  assign n1110 = ~pi104  & ~pi232 ;
  assign n1111 = pi104  & pi232 ;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = ~n1104 & ~n1108;
  assign n1114 = ~n1112 & n1113;
  assign n1115 = n1112 & ~n1113;
  assign po104  = ~n1114 & ~n1115;
  assign n1117 = ~pi105  & ~pi233 ;
  assign n1118 = pi105  & pi233 ;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~n1111 & ~n1115;
  assign n1121 = ~n1119 & n1120;
  assign n1122 = n1119 & ~n1120;
  assign po105  = ~n1121 & ~n1122;
  assign n1124 = ~pi106  & ~pi234 ;
  assign n1125 = pi106  & pi234 ;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = ~n1118 & ~n1122;
  assign n1128 = ~n1126 & n1127;
  assign n1129 = n1126 & ~n1127;
  assign po106  = ~n1128 & ~n1129;
  assign n1131 = ~pi107  & ~pi235 ;
  assign n1132 = pi107  & pi235 ;
  assign n1133 = ~n1131 & ~n1132;
  assign n1134 = ~n1125 & ~n1129;
  assign n1135 = ~n1133 & n1134;
  assign n1136 = n1133 & ~n1134;
  assign po107  = ~n1135 & ~n1136;
  assign n1138 = ~pi108  & ~pi236 ;
  assign n1139 = pi108  & pi236 ;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = ~n1132 & ~n1136;
  assign n1142 = ~n1140 & n1141;
  assign n1143 = n1140 & ~n1141;
  assign po108  = ~n1142 & ~n1143;
  assign n1145 = ~pi109  & ~pi237 ;
  assign n1146 = pi109  & pi237 ;
  assign n1147 = ~n1145 & ~n1146;
  assign n1148 = ~n1139 & ~n1143;
  assign n1149 = ~n1147 & n1148;
  assign n1150 = n1147 & ~n1148;
  assign po109  = ~n1149 & ~n1150;
  assign n1152 = ~pi110  & ~pi238 ;
  assign n1153 = pi110  & pi238 ;
  assign n1154 = ~n1152 & ~n1153;
  assign n1155 = ~n1146 & ~n1150;
  assign n1156 = ~n1154 & n1155;
  assign n1157 = n1154 & ~n1155;
  assign po110  = ~n1156 & ~n1157;
  assign n1159 = ~pi111  & ~pi239 ;
  assign n1160 = pi111  & pi239 ;
  assign n1161 = ~n1159 & ~n1160;
  assign n1162 = ~n1153 & ~n1157;
  assign n1163 = ~n1161 & n1162;
  assign n1164 = n1161 & ~n1162;
  assign po111  = ~n1163 & ~n1164;
  assign n1166 = ~pi112  & ~pi240 ;
  assign n1167 = pi112  & pi240 ;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = ~n1160 & ~n1164;
  assign n1170 = ~n1168 & n1169;
  assign n1171 = n1168 & ~n1169;
  assign po112  = ~n1170 & ~n1171;
  assign n1173 = ~pi113  & ~pi241 ;
  assign n1174 = pi113  & pi241 ;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = ~n1167 & ~n1171;
  assign n1177 = ~n1175 & n1176;
  assign n1178 = n1175 & ~n1176;
  assign po113  = ~n1177 & ~n1178;
  assign n1180 = ~pi114  & ~pi242 ;
  assign n1181 = pi114  & pi242 ;
  assign n1182 = ~n1180 & ~n1181;
  assign n1183 = ~n1174 & ~n1178;
  assign n1184 = ~n1182 & n1183;
  assign n1185 = n1182 & ~n1183;
  assign po114  = ~n1184 & ~n1185;
  assign n1187 = ~pi115  & ~pi243 ;
  assign n1188 = pi115  & pi243 ;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1181 & ~n1185;
  assign n1191 = ~n1189 & n1190;
  assign n1192 = n1189 & ~n1190;
  assign po115  = ~n1191 & ~n1192;
  assign n1194 = ~pi116  & ~pi244 ;
  assign n1195 = pi116  & pi244 ;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = ~n1188 & ~n1192;
  assign n1198 = ~n1196 & n1197;
  assign n1199 = n1196 & ~n1197;
  assign po116  = ~n1198 & ~n1199;
  assign n1201 = ~pi117  & ~pi245 ;
  assign n1202 = pi117  & pi245 ;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = ~n1195 & ~n1199;
  assign n1205 = ~n1203 & n1204;
  assign n1206 = n1203 & ~n1204;
  assign po117  = ~n1205 & ~n1206;
  assign n1208 = ~pi118  & ~pi246 ;
  assign n1209 = pi118  & pi246 ;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = ~n1202 & ~n1206;
  assign n1212 = ~n1210 & n1211;
  assign n1213 = n1210 & ~n1211;
  assign po118  = ~n1212 & ~n1213;
  assign n1215 = ~pi119  & ~pi247 ;
  assign n1216 = pi119  & pi247 ;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = ~n1209 & ~n1213;
  assign n1219 = ~n1217 & n1218;
  assign n1220 = n1217 & ~n1218;
  assign po119  = ~n1219 & ~n1220;
  assign n1222 = ~pi120  & ~pi248 ;
  assign n1223 = pi120  & pi248 ;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = ~n1216 & ~n1220;
  assign n1226 = ~n1224 & n1225;
  assign n1227 = n1224 & ~n1225;
  assign po120  = ~n1226 & ~n1227;
  assign n1229 = ~pi121  & ~pi249 ;
  assign n1230 = pi121  & pi249 ;
  assign n1231 = ~n1229 & ~n1230;
  assign n1232 = ~n1223 & ~n1227;
  assign n1233 = ~n1231 & n1232;
  assign n1234 = n1231 & ~n1232;
  assign po121  = ~n1233 & ~n1234;
  assign n1236 = ~pi122  & ~pi250 ;
  assign n1237 = pi122  & pi250 ;
  assign n1238 = ~n1236 & ~n1237;
  assign n1239 = ~n1230 & ~n1234;
  assign n1240 = ~n1238 & n1239;
  assign n1241 = n1238 & ~n1239;
  assign po122  = ~n1240 & ~n1241;
  assign n1243 = ~pi123  & ~pi251 ;
  assign n1244 = pi123  & pi251 ;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = ~n1237 & ~n1241;
  assign n1247 = ~n1245 & n1246;
  assign n1248 = n1245 & ~n1246;
  assign po123  = ~n1247 & ~n1248;
  assign n1250 = ~pi124  & ~pi252 ;
  assign n1251 = pi124  & pi252 ;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = ~n1244 & ~n1248;
  assign n1254 = ~n1252 & n1253;
  assign n1255 = n1252 & ~n1253;
  assign po124  = ~n1254 & ~n1255;
  assign n1257 = ~pi125  & ~pi253 ;
  assign n1258 = pi125  & pi253 ;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = ~n1251 & ~n1255;
  assign n1261 = ~n1259 & n1260;
  assign n1262 = n1259 & ~n1260;
  assign po125  = ~n1261 & ~n1262;
  assign n1264 = ~pi126  & ~pi254 ;
  assign n1265 = pi126  & pi254 ;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = ~n1258 & ~n1262;
  assign n1268 = ~n1266 & n1267;
  assign n1269 = n1266 & ~n1267;
  assign po126  = ~n1268 & ~n1269;
  assign n1271 = ~pi127  & ~pi255 ;
  assign n1272 = pi127  & pi255 ;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = ~n1265 & ~n1269;
  assign n1275 = ~n1273 & n1274;
  assign n1276 = n1273 & ~n1274;
  assign po127  = ~n1275 & ~n1276;
  assign po128 = n1272 | n1276;
endmodule
