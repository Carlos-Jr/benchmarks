module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n414, n415, n416, n417, n418,
    n419, n420, n422, n423, n424, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504,
    n505, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589,
    n590, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646,
    n647, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682,
    n684, n685, n686, n687, n688, n689;
  assign n22 = ~pi0  & pi9 ;
  assign n23 = pi1  & ~n22;
  assign n24 = ~pi3  & ~pi5 ;
  assign n25 = ~pi1  & pi9 ;
  assign n26 = n24 & ~n25;
  assign n27 = ~n23 & n26;
  assign n28 = pi0  & ~pi9 ;
  assign n29 = ~pi1  & ~n28;
  assign n30 = pi1  & ~pi9 ;
  assign n31 = ~pi7  & ~n30;
  assign n32 = ~n29 & n31;
  assign n33 = ~n27 & ~n32;
  assign n34 = ~pi2  & ~n33;
  assign n35 = ~pi2  & ~pi3 ;
  assign n36 = pi9  & ~n35;
  assign n37 = pi0  & pi3 ;
  assign n38 = ~n36 & ~n37;
  assign n39 = ~pi1  & ~n38;
  assign n40 = ~pi0  & pi5 ;
  assign n41 = ~pi0  & pi2 ;
  assign n42 = pi1  & pi2 ;
  assign n43 = ~n40 & ~n41;
  assign n44 = ~n42 & n43;
  assign n45 = ~pi9  & ~n44;
  assign n46 = pi1  & ~pi3 ;
  assign n47 = ~n39 & ~n46;
  assign n48 = ~n45 & n47;
  assign n49 = ~pi7  & ~n48;
  assign n50 = ~n34 & ~n49;
  assign n51 = ~pi8  & ~n50;
  assign n52 = pi7  & pi8 ;
  assign n53 = ~pi5  & n52;
  assign n54 = ~pi7  & pi9 ;
  assign n55 = ~n53 & ~n54;
  assign n56 = pi1  & ~n55;
  assign n57 = pi1  & ~pi7 ;
  assign n58 = ~pi5  & ~pi9 ;
  assign n59 = ~n57 & n58;
  assign n60 = ~n56 & ~n59;
  assign n61 = pi0  & ~pi2 ;
  assign n62 = ~n60 & n61;
  assign n63 = pi2  & ~pi9 ;
  assign n64 = ~pi0  & ~pi1 ;
  assign n65 = n63 & n64;
  assign n66 = n53 & n65;
  assign n67 = ~n62 & ~n66;
  assign n68 = ~pi3  & ~n67;
  assign n69 = ~n51 & ~n68;
  assign n70 = ~pi6  & ~n69;
  assign n71 = ~pi2  & ~n28;
  assign n72 = pi6  & ~n71;
  assign n73 = ~pi0  & ~pi9 ;
  assign n74 = pi0  & pi9 ;
  assign n75 = ~n73 & ~n74;
  assign n76 = pi1  & ~n75;
  assign n77 = n35 & n76;
  assign n78 = ~n72 & ~n77;
  assign n79 = pi5  & ~n78;
  assign n80 = pi2  & pi9 ;
  assign n81 = ~pi2  & n30;
  assign n82 = ~n80 & ~n81;
  assign n83 = ~pi0  & ~pi3 ;
  assign n84 = pi6  & n83;
  assign n85 = ~n82 & n84;
  assign n86 = ~n79 & ~n85;
  assign n87 = pi8  & ~n86;
  assign n88 = ~pi0  & ~pi2 ;
  assign n89 = n25 & n88;
  assign n90 = ~pi5  & ~n89;
  assign n91 = pi6  & ~n90;
  assign n92 = pi2  & pi5 ;
  assign n93 = n76 & n92;
  assign n94 = ~n91 & ~n93;
  assign n95 = pi8  & ~n94;
  assign n96 = ~pi1  & ~n22;
  assign n97 = ~pi8  & ~n96;
  assign n98 = ~pi1  & pi2 ;
  assign n99 = n28 & n98;
  assign n100 = ~n97 & ~n99;
  assign n101 = ~pi5  & ~n100;
  assign n102 = ~n95 & ~n101;
  assign n103 = pi3  & ~n102;
  assign n104 = pi2  & ~pi3 ;
  assign n105 = n25 & n104;
  assign n106 = pi1  & ~pi8 ;
  assign n107 = ~n105 & ~n106;
  assign n108 = ~pi0  & ~n107;
  assign n109 = pi3  & ~pi6 ;
  assign n110 = pi2  & pi3 ;
  assign n111 = ~pi1  & ~pi9 ;
  assign n112 = ~n109 & ~n110;
  assign n113 = n111 & n112;
  assign n114 = ~n80 & ~n113;
  assign n115 = ~pi8  & ~n114;
  assign n116 = ~n108 & ~n115;
  assign n117 = ~pi5  & ~n116;
  assign n118 = ~pi1  & ~pi3 ;
  assign n119 = ~pi2  & ~pi8 ;
  assign n120 = n73 & n119;
  assign n121 = n118 & n120;
  assign n122 = ~n117 & ~n121;
  assign n123 = ~n87 & n122;
  assign n124 = ~n103 & n123;
  assign n125 = ~pi7  & ~n124;
  assign n126 = ~n70 & ~n125;
  assign n127 = ~pi4  & ~n126;
  assign n128 = ~pi8  & ~pi9 ;
  assign n129 = ~pi6  & n128;
  assign n130 = pi4  & pi8 ;
  assign n131 = pi6  & n130;
  assign n132 = ~n129 & ~n131;
  assign n133 = pi5  & ~n132;
  assign n134 = pi6  & ~pi9 ;
  assign n135 = pi4  & pi9 ;
  assign n136 = ~n134 & ~n135;
  assign n137 = pi5  & pi6 ;
  assign n138 = ~pi8  & ~n137;
  assign n139 = ~n136 & n138;
  assign n140 = ~n133 & ~n139;
  assign n141 = ~pi2  & n118;
  assign n142 = ~pi0  & ~pi7 ;
  assign n143 = n141 & n142;
  assign n144 = ~n140 & n143;
  assign po0  = n127 | n144;
  assign n146 = pi0  & pi8 ;
  assign n147 = n80 & n146;
  assign n148 = ~n120 & ~n147;
  assign n149 = pi5  & ~n148;
  assign n150 = ~pi5  & pi8 ;
  assign n151 = pi6  & pi9 ;
  assign n152 = ~n150 & ~n151;
  assign n153 = ~pi0  & ~n152;
  assign n154 = pi8  & n151;
  assign n155 = ~pi8  & n58;
  assign n156 = ~n154 & ~n155;
  assign n157 = ~n153 & n156;
  assign n158 = pi2  & ~n157;
  assign n159 = ~n149 & ~n158;
  assign n160 = ~pi4  & ~n159;
  assign n161 = pi5  & ~pi8 ;
  assign n162 = ~n130 & ~n161;
  assign n163 = ~pi6  & ~n162;
  assign n164 = ~n135 & ~n163;
  assign n165 = ~pi6  & pi9 ;
  assign n166 = n88 & ~n165;
  assign n167 = ~n164 & n166;
  assign n168 = ~n160 & ~n167;
  assign n169 = ~pi1  & ~n168;
  assign n170 = pi6  & pi8 ;
  assign n171 = pi0  & ~n170;
  assign n172 = ~n152 & n171;
  assign n173 = ~pi8  & pi9 ;
  assign n174 = n40 & n173;
  assign n175 = ~n172 & ~n174;
  assign n176 = ~pi2  & ~n175;
  assign n177 = ~pi6  & ~pi8 ;
  assign n178 = ~pi0  & pi6 ;
  assign n179 = ~pi2  & ~n178;
  assign n180 = n150 & ~n179;
  assign n181 = ~n177 & ~n180;
  assign n182 = ~pi9  & ~n181;
  assign n183 = ~n176 & ~n182;
  assign n184 = pi1  & ~n183;
  assign n185 = ~pi6  & pi8 ;
  assign n186 = n63 & n185;
  assign n187 = ~n184 & ~n186;
  assign n188 = ~pi4  & ~n187;
  assign n189 = ~n169 & ~n188;
  assign n190 = ~pi3  & ~n189;
  assign n191 = pi5  & n119;
  assign n192 = ~pi3  & ~pi8 ;
  assign n193 = ~n150 & ~n192;
  assign n194 = pi0  & n193;
  assign n195 = ~n191 & ~n194;
  assign n196 = ~pi1  & ~n195;
  assign n197 = ~n35 & ~n119;
  assign n198 = ~pi0  & n197;
  assign n199 = ~pi2  & pi8 ;
  assign n200 = pi0  & n199;
  assign n201 = pi0  & ~pi5 ;
  assign n202 = ~n40 & ~n201;
  assign n203 = ~n200 & n202;
  assign n204 = pi1  & ~n203;
  assign n205 = ~n198 & ~n204;
  assign n206 = ~n196 & n205;
  assign n207 = ~pi6  & ~n206;
  assign n208 = ~pi1  & pi6 ;
  assign n209 = pi2  & ~n208;
  assign n210 = ~pi1  & ~pi8 ;
  assign n211 = pi3  & ~n210;
  assign n212 = ~n209 & n211;
  assign n213 = ~pi0  & pi8 ;
  assign n214 = ~pi1  & ~pi6 ;
  assign n215 = pi0  & pi1 ;
  assign n216 = ~pi2  & ~n213;
  assign n217 = ~n214 & ~n215;
  assign n218 = n216 & n217;
  assign n219 = ~n212 & ~n218;
  assign n220 = ~pi5  & ~n219;
  assign n221 = ~n207 & ~n220;
  assign n222 = ~pi9  & ~n221;
  assign n223 = pi1  & pi5 ;
  assign n224 = pi3  & ~pi8 ;
  assign n225 = ~pi1  & ~pi2 ;
  assign n226 = n224 & n225;
  assign n227 = ~n223 & ~n226;
  assign n228 = pi0  & ~n227;
  assign n229 = pi5  & ~n35;
  assign n230 = pi3  & n42;
  assign n231 = ~n229 & ~n230;
  assign n232 = ~n228 & n231;
  assign n233 = pi6  & ~n232;
  assign n234 = n161 & n230;
  assign n235 = ~n233 & ~n234;
  assign n236 = pi9  & ~n235;
  assign n237 = ~n222 & ~n236;
  assign n238 = ~pi4  & ~n237;
  assign n239 = ~n190 & ~n238;
  assign n240 = ~pi7  & ~n239;
  assign n241 = n71 & ~n215;
  assign n242 = pi2  & ~n64;
  assign n243 = ~pi8  & ~n242;
  assign n244 = ~n241 & n243;
  assign n245 = n30 & n199;
  assign n246 = ~n244 & ~n245;
  assign n247 = pi7  & ~n246;
  assign n248 = ~n65 & ~n247;
  assign n249 = ~pi6  & n24;
  assign n250 = ~pi4  & n249;
  assign n251 = ~n248 & n250;
  assign po1  = n240 | n251;
  assign n253 = pi3  & ~n199;
  assign n254 = pi5  & ~n253;
  assign n255 = pi2  & ~pi5 ;
  assign n256 = pi3  & ~n255;
  assign n257 = pi8  & ~n256;
  assign n258 = ~n254 & ~n257;
  assign n259 = pi1  & ~n258;
  assign n260 = ~pi5  & pi6 ;
  assign n261 = ~pi8  & n260;
  assign n262 = n118 & n261;
  assign n263 = ~n259 & ~n262;
  assign n264 = ~pi9  & ~n263;
  assign n265 = pi6  & ~pi8 ;
  assign n266 = ~pi9  & ~n208;
  assign n267 = ~n265 & n266;
  assign n268 = ~pi2  & ~n267;
  assign n269 = ~pi1  & n173;
  assign n270 = ~n268 & ~n269;
  assign n271 = pi3  & ~n270;
  assign n272 = ~pi1  & n197;
  assign n273 = pi2  & ~n185;
  assign n274 = ~n272 & ~n273;
  assign n275 = pi5  & ~n274;
  assign n276 = ~n46 & ~n173;
  assign n277 = ~pi3  & pi9 ;
  assign n278 = ~pi6  & ~n277;
  assign n279 = ~n276 & n278;
  assign n280 = pi1  & n277;
  assign n281 = n265 & n280;
  assign n282 = ~n279 & ~n281;
  assign n283 = ~n275 & n282;
  assign n284 = ~n271 & n283;
  assign n285 = ~n264 & n284;
  assign n286 = ~pi4  & ~n285;
  assign n287 = pi8  & ~pi9 ;
  assign n288 = ~pi5  & ~n177;
  assign n289 = ~n287 & n288;
  assign n290 = ~pi3  & pi4 ;
  assign n291 = n225 & n290;
  assign n292 = ~n289 & n291;
  assign n293 = ~n286 & ~n292;
  assign n294 = ~pi0  & ~n293;
  assign n295 = pi8  & n74;
  assign n296 = ~n128 & ~n295;
  assign n297 = pi5  & ~n296;
  assign n298 = ~pi5  & n80;
  assign n299 = ~n297 & ~n298;
  assign n300 = pi1  & ~n299;
  assign n301 = pi8  & pi9 ;
  assign n302 = ~n128 & ~n301;
  assign n303 = ~n111 & ~n302;
  assign n304 = pi2  & ~n303;
  assign n305 = ~n300 & ~n304;
  assign n306 = ~pi3  & ~n305;
  assign n307 = ~pi1  & pi3 ;
  assign n308 = pi5  & ~n307;
  assign n309 = ~pi2  & n128;
  assign n310 = ~n308 & n309;
  assign n311 = ~pi1  & pi8 ;
  assign n312 = n36 & n311;
  assign n313 = ~n310 & ~n312;
  assign n314 = pi0  & ~n313;
  assign n315 = ~n306 & ~n314;
  assign n316 = ~pi6  & ~n315;
  assign n317 = pi1  & pi9 ;
  assign n318 = pi2  & n317;
  assign n319 = ~n311 & ~n318;
  assign n320 = pi6  & ~n319;
  assign n321 = pi8  & ~n63;
  assign n322 = pi2  & n128;
  assign n323 = ~n321 & ~n322;
  assign n324 = ~n320 & n323;
  assign n325 = pi3  & ~n324;
  assign n326 = pi6  & ~n25;
  assign n327 = ~n30 & ~n326;
  assign n328 = pi8  & ~n327;
  assign n329 = ~n111 & ~n317;
  assign n330 = n192 & ~n329;
  assign n331 = ~n328 & ~n330;
  assign n332 = ~pi2  & ~n331;
  assign n333 = ~n325 & ~n332;
  assign n334 = n201 & ~n333;
  assign n335 = ~n316 & ~n334;
  assign n336 = ~pi4  & ~n335;
  assign n337 = ~n294 & ~n336;
  assign n338 = ~pi7  & ~n337;
  assign n339 = n52 & n74;
  assign n340 = ~n73 & ~n339;
  assign n341 = pi1  & ~n340;
  assign n342 = n28 & n210;
  assign n343 = ~n341 & ~n342;
  assign n344 = ~pi2  & n250;
  assign n345 = ~n343 & n344;
  assign po2  = n338 | n345;
  assign n347 = pi3  & ~n165;
  assign n348 = pi2  & pi6 ;
  assign n349 = ~n347 & ~n348;
  assign n350 = ~pi4  & ~n349;
  assign n351 = ~pi5  & ~pi6 ;
  assign n352 = n301 & n351;
  assign n353 = ~n137 & ~n352;
  assign n354 = ~pi2  & n290;
  assign n355 = ~n353 & n354;
  assign n356 = ~n350 & ~n355;
  assign n357 = ~pi1  & ~n356;
  assign n358 = pi5  & pi8 ;
  assign n359 = n165 & n358;
  assign n360 = ~n155 & ~n359;
  assign n361 = pi2  & ~n360;
  assign n362 = ~pi6  & ~n224;
  assign n363 = pi3  & ~pi5 ;
  assign n364 = ~n362 & ~n363;
  assign n365 = pi3  & ~n364;
  assign n366 = ~n261 & ~n361;
  assign n367 = ~n365 & n366;
  assign n368 = pi1  & ~n367;
  assign n369 = pi2  & n260;
  assign n370 = ~n368 & ~n369;
  assign n371 = ~pi4  & ~n370;
  assign n372 = ~n357 & ~n371;
  assign n373 = ~pi0  & ~n372;
  assign n374 = pi2  & ~n193;
  assign n375 = ~pi2  & n358;
  assign n376 = ~n374 & ~n375;
  assign n377 = ~pi9  & ~n376;
  assign n378 = pi5  & pi9 ;
  assign n379 = ~pi8  & n378;
  assign n380 = ~pi3  & ~n379;
  assign n381 = ~pi2  & ~n380;
  assign n382 = ~n364 & ~n381;
  assign n383 = ~n377 & n382;
  assign n384 = pi1  & ~n383;
  assign n385 = ~pi3  & n260;
  assign n386 = n191 & n214;
  assign n387 = ~n385 & ~n386;
  assign n388 = ~pi9  & ~n387;
  assign n389 = ~n384 & ~n388;
  assign n390 = pi0  & ~n389;
  assign n391 = ~n35 & n260;
  assign n392 = pi2  & n109;
  assign n393 = ~n391 & ~n392;
  assign n394 = pi9  & ~n393;
  assign n395 = ~pi9  & n260;
  assign n396 = ~n109 & ~n395;
  assign n397 = ~pi8  & ~n396;
  assign n398 = ~n394 & ~n397;
  assign n399 = ~pi1  & ~n398;
  assign n400 = ~n58 & ~n177;
  assign n401 = ~pi2  & ~n400;
  assign n402 = ~pi6  & ~n378;
  assign n403 = ~n317 & ~n358;
  assign n404 = n402 & ~n403;
  assign n405 = ~n401 & ~n404;
  assign n406 = pi3  & ~n405;
  assign n407 = n260 & n267;
  assign n408 = ~n406 & ~n407;
  assign n409 = ~n399 & n408;
  assign n410 = ~n390 & n409;
  assign n411 = ~pi4  & ~n410;
  assign n412 = ~n373 & ~n411;
  assign po3  = ~pi7  & ~n412;
  assign n414 = ~pi4  & n242;
  assign n415 = pi3  & ~pi4 ;
  assign n416 = ~n290 & ~n415;
  assign n417 = ~pi0  & n225;
  assign n418 = ~n416 & n417;
  assign n419 = ~n414 & ~n418;
  assign n420 = ~pi7  & n137;
  assign po4  = ~n419 & n420;
  assign n422 = n415 & ~n417;
  assign n423 = pi4  & n418;
  assign n424 = ~n422 & ~n423;
  assign po5  = n420 & ~n424;
  assign n426 = ~pi1  & ~pi5 ;
  assign n427 = pi2  & ~n426;
  assign n428 = ~pi6  & ~pi9 ;
  assign n429 = ~n427 & n428;
  assign n430 = pi5  & n317;
  assign n431 = ~n429 & ~n430;
  assign n432 = pi0  & ~n431;
  assign n433 = n41 & ~n58;
  assign n434 = ~n432 & ~n433;
  assign n435 = pi8  & ~n434;
  assign n436 = ~pi8  & n111;
  assign n437 = pi2  & n22;
  assign n438 = ~n436 & ~n437;
  assign n439 = pi5  & ~n438;
  assign n440 = pi6  & ~n302;
  assign n441 = ~pi2  & pi9 ;
  assign n442 = ~n63 & ~n441;
  assign n443 = n440 & n442;
  assign n444 = ~n439 & ~n443;
  assign n445 = ~n435 & n444;
  assign n446 = ~pi7  & ~n445;
  assign n447 = ~pi9  & n52;
  assign n448 = pi8  & ~n447;
  assign n449 = n98 & ~n448;
  assign n450 = ~n81 & ~n449;
  assign n451 = ~pi0  & ~n450;
  assign n452 = ~pi2  & pi7 ;
  assign n453 = ~n311 & n452;
  assign n454 = ~n296 & n453;
  assign n455 = ~n451 & ~n454;
  assign n456 = n351 & ~n455;
  assign n457 = ~n446 & ~n456;
  assign n458 = ~pi3  & ~n457;
  assign n459 = ~pi8  & n215;
  assign n460 = pi0  & n170;
  assign n461 = ~n106 & ~n460;
  assign n462 = ~pi2  & ~n461;
  assign n463 = ~n459 & ~n462;
  assign n464 = pi9  & ~n463;
  assign n465 = ~n317 & ~n436;
  assign n466 = pi0  & ~n465;
  assign n467 = pi2  & n30;
  assign n468 = ~pi0  & ~pi6 ;
  assign n469 = ~n210 & n468;
  assign n470 = n329 & n469;
  assign n471 = ~n467 & ~n470;
  assign n472 = ~n466 & n471;
  assign n473 = ~pi5  & ~n472;
  assign n474 = ~pi0  & ~pi8 ;
  assign n475 = n30 & ~n201;
  assign n476 = ~n474 & n475;
  assign n477 = ~n464 & ~n476;
  assign n478 = ~n473 & n477;
  assign n479 = pi3  & ~n478;
  assign n480 = ~pi2  & pi5 ;
  assign n481 = ~n75 & n480;
  assign n482 = ~pi6  & ~n255;
  assign n483 = n22 & ~n482;
  assign n484 = ~n481 & ~n483;
  assign n485 = ~pi8  & ~n484;
  assign n486 = pi2  & ~n128;
  assign n487 = ~n295 & ~n486;
  assign n488 = pi6  & ~n487;
  assign n489 = ~n485 & ~n488;
  assign n490 = pi1  & ~n489;
  assign n491 = ~pi8  & ~n468;
  assign n492 = ~n201 & ~n491;
  assign n493 = ~pi2  & ~pi9 ;
  assign n494 = ~n492 & n493;
  assign n495 = pi2  & pi8 ;
  assign n496 = n22 & n495;
  assign n497 = ~n494 & ~n496;
  assign n498 = ~pi1  & ~n497;
  assign n499 = ~n490 & ~n498;
  assign n500 = ~n479 & n499;
  assign n501 = ~pi7  & ~n500;
  assign n502 = ~n458 & ~n501;
  assign n503 = ~pi4  & ~n502;
  assign n504 = ~n137 & ~n423;
  assign n505 = ~pi7  & ~n504;
  assign po6  = ~n503 & ~n505;
  assign n507 = ~pi3  & n301;
  assign n508 = pi3  & ~n301;
  assign n509 = ~n146 & ~n508;
  assign n510 = ~pi6  & ~n509;
  assign n511 = ~n507 & ~n510;
  assign n512 = pi2  & ~n511;
  assign n513 = n109 & n213;
  assign n514 = ~n265 & ~n513;
  assign n515 = pi9  & ~n514;
  assign n516 = ~pi3  & pi8 ;
  assign n517 = ~n151 & ~n516;
  assign n518 = pi0  & ~n517;
  assign n519 = ~pi9  & n170;
  assign n520 = ~n518 & ~n519;
  assign n521 = ~n515 & n520;
  assign n522 = ~pi2  & ~n521;
  assign n523 = ~pi3  & n129;
  assign n524 = ~n512 & ~n523;
  assign n525 = ~n522 & n524;
  assign n526 = pi1  & ~n525;
  assign n527 = ~n73 & ~n173;
  assign n528 = ~pi2  & ~pi6 ;
  assign n529 = ~n527 & n528;
  assign n530 = ~pi0  & n440;
  assign n531 = ~n529 & ~n530;
  assign n532 = pi3  & ~n531;
  assign n533 = ~pi0  & n119;
  assign n534 = ~n460 & ~n533;
  assign n535 = ~pi9  & ~n534;
  assign n536 = ~pi6  & ~n192;
  assign n537 = n486 & ~n536;
  assign n538 = ~n535 & ~n537;
  assign n539 = ~n532 & n538;
  assign n540 = ~pi1  & ~n539;
  assign n541 = ~pi2  & pi3 ;
  assign n542 = n443 & n541;
  assign n543 = ~n540 & ~n542;
  assign n544 = ~n526 & n543;
  assign n545 = ~pi5  & ~n544;
  assign n546 = pi0  & ~n442;
  assign n547 = pi5  & ~pi9 ;
  assign n548 = ~pi0  & n547;
  assign n549 = ~n546 & ~n548;
  assign n550 = pi8  & ~n549;
  assign n551 = n80 & n161;
  assign n552 = ~n550 & ~n551;
  assign n553 = ~pi3  & ~n552;
  assign n554 = pi3  & pi5 ;
  assign n555 = ~n63 & ~n554;
  assign n556 = ~pi0  & ~n555;
  assign n557 = pi3  & n480;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~pi8  & ~n558;
  assign n560 = n541 & n547;
  assign n561 = ~n559 & ~n560;
  assign n562 = ~n553 & n561;
  assign n563 = pi1  & ~n562;
  assign n564 = ~pi2  & ~n37;
  assign n565 = ~n302 & ~n564;
  assign n566 = ~n110 & ~n565;
  assign n567 = pi5  & ~n566;
  assign n568 = n37 & n322;
  assign n569 = ~n567 & ~n568;
  assign n570 = ~pi1  & ~n569;
  assign n571 = pi8  & n378;
  assign n572 = n110 & n571;
  assign n573 = ~n570 & ~n572;
  assign n574 = ~n563 & n573;
  assign n575 = ~pi6  & ~n574;
  assign n576 = ~n545 & ~n575;
  assign n577 = ~pi7  & ~n576;
  assign n578 = n41 & n302;
  assign n579 = n61 & n447;
  assign n580 = ~n578 & ~n579;
  assign n581 = n24 & n214;
  assign n582 = ~n580 & n581;
  assign n583 = ~n577 & ~n582;
  assign n584 = ~pi4  & ~n583;
  assign n585 = pi4  & ~pi7 ;
  assign n586 = n24 & n585;
  assign n587 = n417 & n586;
  assign n588 = pi4  & ~n351;
  assign n589 = ~pi3  & ~n588;
  assign n590 = n587 & n589;
  assign po7  = ~n584 & ~n590;
  assign n592 = ~n223 & ~n363;
  assign n593 = ~pi2  & ~n83;
  assign n594 = n592 & n593;
  assign n595 = n118 & n201;
  assign n596 = ~n594 & ~n595;
  assign n597 = pi8  & ~n596;
  assign n598 = ~pi5  & ~n213;
  assign n599 = n42 & ~n554;
  assign n600 = ~n598 & n599;
  assign n601 = ~n597 & ~n600;
  assign n602 = ~pi9  & ~n601;
  assign n603 = n225 & n547;
  assign n604 = ~n280 & ~n603;
  assign n605 = ~pi0  & ~n604;
  assign n606 = ~pi2  & ~n111;
  assign n607 = ~n277 & n606;
  assign n608 = n592 & n607;
  assign n609 = n329 & ~n426;
  assign n610 = n104 & ~n609;
  assign n611 = ~n605 & ~n608;
  assign n612 = ~n610 & n611;
  assign n613 = ~pi8  & ~n612;
  assign n614 = ~n255 & ~n554;
  assign n615 = pi1  & ~n253;
  assign n616 = ~n614 & n615;
  assign n617 = ~n40 & n199;
  assign n618 = n307 & n617;
  assign n619 = ~n616 & ~n618;
  assign n620 = pi9  & ~n619;
  assign n621 = ~n602 & ~n620;
  assign n622 = ~n613 & n621;
  assign n623 = ~pi6  & ~n622;
  assign n624 = ~pi1  & ~n128;
  assign n625 = pi2  & ~n624;
  assign n626 = ~n326 & ~n625;
  assign n627 = pi0  & ~n626;
  assign n628 = pi8  & ~n30;
  assign n629 = n326 & ~n628;
  assign n630 = ~n214 & n273;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n627 & n631;
  assign n633 = n363 & ~n632;
  assign n634 = ~n623 & ~n633;
  assign n635 = ~pi7  & ~n634;
  assign n636 = ~n119 & ~n495;
  assign n637 = ~pi0  & ~n636;
  assign n638 = ~n200 & ~n637;
  assign n639 = ~pi9  & ~n638;
  assign n640 = n80 & n474;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~pi1  & ~n641;
  assign n643 = n317 & n533;
  assign n644 = ~n642 & ~n643;
  assign n645 = n249 & ~n644;
  assign n646 = ~n635 & ~n645;
  assign n647 = ~pi4  & ~n646;
  assign po8  = ~n587 & ~n647;
  assign n649 = n213 & ~n402;
  assign n650 = ~n151 & ~n649;
  assign n651 = pi3  & ~n650;
  assign n652 = ~n589 & ~n651;
  assign n653 = ~pi2  & ~n652;
  assign n654 = ~pi3  & ~n58;
  assign n655 = ~n495 & ~n551;
  assign n656 = n654 & ~n655;
  assign n657 = ~n653 & ~n656;
  assign n658 = ~pi1  & ~n657;
  assign n659 = n213 & ~n517;
  assign n660 = ~n654 & ~n659;
  assign n661 = ~pi2  & ~n660;
  assign n662 = ~pi5  & ~n301;
  assign n663 = n392 & n662;
  assign n664 = ~pi6  & ~n571;
  assign n665 = ~pi3  & ~n664;
  assign n666 = ~n663 & ~n665;
  assign n667 = ~n661 & n666;
  assign n668 = pi1  & ~n667;
  assign n669 = n201 & n392;
  assign n670 = ~pi7  & ~n669;
  assign n671 = ~n624 & ~n670;
  assign n672 = ~pi7  & ~n141;
  assign n673 = pi0  & ~n672;
  assign n674 = ~pi5  & ~n104;
  assign n675 = pi6  & ~n674;
  assign n676 = pi4  & ~n141;
  assign n677 = pi7  & ~n104;
  assign n678 = ~n675 & ~n677;
  assign n679 = ~n676 & n678;
  assign n680 = ~n673 & n679;
  assign n681 = ~n671 & n680;
  assign n682 = ~n668 & n681;
  assign po9  = ~n658 & n682;
  assign n684 = ~pi8  & ~n29;
  assign n685 = ~n23 & ~n684;
  assign n686 = pi2  & n415;
  assign n687 = ~n685 & n686;
  assign n688 = ~n423 & ~n687;
  assign n689 = ~pi7  & n351;
  assign po10  = ~n688 & n689;
endmodule
