module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n403, n404,
    n405, n406, n407, n408, n410, n411, n412,
    n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647,
    n648, n650, n651, n652, n653, n654, n655;
  assign n22 = pi1  & ~pi9 ;
  assign n23 = pi0  & ~pi9 ;
  assign n24 = ~pi1  & ~n23;
  assign n25 = ~pi7  & ~n22;
  assign n26 = ~n24 & n25;
  assign n27 = ~pi3  & ~pi5 ;
  assign n28 = ~pi0  & pi9 ;
  assign n29 = pi1  & ~n28;
  assign n30 = ~pi1  & pi9 ;
  assign n31 = n27 & ~n30;
  assign n32 = ~n29 & n31;
  assign n33 = ~n26 & ~n32;
  assign n34 = ~pi2  & ~n33;
  assign n35 = ~pi2  & ~pi3 ;
  assign n36 = pi9  & ~n35;
  assign n37 = pi0  & pi3 ;
  assign n38 = ~n36 & ~n37;
  assign n39 = ~pi1  & ~n38;
  assign n40 = pi1  & ~pi3 ;
  assign n41 = pi0  & ~n22;
  assign n42 = pi2  & ~pi9 ;
  assign n43 = ~n23 & ~n28;
  assign n44 = ~pi2  & pi5 ;
  assign n45 = n43 & n44;
  assign n46 = ~n42 & ~n45;
  assign n47 = ~n41 & ~n46;
  assign n48 = ~n40 & ~n47;
  assign n49 = ~n39 & n48;
  assign n50 = ~pi7  & ~n49;
  assign n51 = ~n34 & ~n50;
  assign n52 = ~pi8  & ~n51;
  assign n53 = pi7  & pi8 ;
  assign n54 = ~pi5  & n53;
  assign n55 = ~pi7  & pi9 ;
  assign n56 = ~n54 & ~n55;
  assign n57 = pi1  & ~n56;
  assign n58 = pi1  & ~pi7 ;
  assign n59 = ~pi5  & ~pi9 ;
  assign n60 = ~n58 & n59;
  assign n61 = ~n57 & ~n60;
  assign n62 = pi0  & ~pi2 ;
  assign n63 = ~n61 & n62;
  assign n64 = ~pi0  & ~pi1 ;
  assign n65 = n42 & n64;
  assign n66 = n54 & n65;
  assign n67 = ~n63 & ~n66;
  assign n68 = ~pi3  & ~n67;
  assign n69 = ~n52 & ~n68;
  assign n70 = ~pi6  & ~n69;
  assign n71 = ~pi3  & ~pi8 ;
  assign n72 = ~pi1  & ~pi9 ;
  assign n73 = pi1  & pi9 ;
  assign n74 = ~n72 & ~n73;
  assign n75 = n71 & ~n74;
  assign n76 = ~pi1  & ~pi2 ;
  assign n77 = ~pi0  & n76;
  assign n78 = n75 & n77;
  assign n79 = ~pi2  & ~n23;
  assign n80 = pi6  & ~n79;
  assign n81 = pi1  & n43;
  assign n82 = n35 & n81;
  assign n83 = ~n80 & ~n82;
  assign n84 = pi5  & ~n83;
  assign n85 = pi2  & pi9 ;
  assign n86 = ~pi2  & n22;
  assign n87 = ~n85 & ~n86;
  assign n88 = ~pi0  & ~pi3 ;
  assign n89 = pi6  & n88;
  assign n90 = ~n87 & n89;
  assign n91 = ~n84 & ~n90;
  assign n92 = pi8  & ~n91;
  assign n93 = pi1  & ~pi8 ;
  assign n94 = pi2  & ~pi3 ;
  assign n95 = n30 & n94;
  assign n96 = ~n93 & ~n95;
  assign n97 = ~pi0  & ~n96;
  assign n98 = pi3  & ~pi6 ;
  assign n99 = pi2  & pi3 ;
  assign n100 = n72 & ~n98;
  assign n101 = ~n99 & n100;
  assign n102 = ~n85 & ~n101;
  assign n103 = ~pi8  & ~n102;
  assign n104 = ~n97 & ~n103;
  assign n105 = ~pi5  & ~n104;
  assign n106 = ~pi1  & ~n28;
  assign n107 = ~pi8  & ~n106;
  assign n108 = ~pi1  & pi2 ;
  assign n109 = n23 & n108;
  assign n110 = ~n107 & ~n109;
  assign n111 = ~pi5  & ~n110;
  assign n112 = ~pi0  & ~pi2 ;
  assign n113 = ~pi6  & pi9 ;
  assign n114 = n112 & ~n113;
  assign n115 = n30 & n114;
  assign n116 = pi5  & pi6 ;
  assign n117 = pi2  & pi5 ;
  assign n118 = n81 & n117;
  assign n119 = ~n115 & ~n116;
  assign n120 = ~n118 & n119;
  assign n121 = pi8  & ~n120;
  assign n122 = ~n111 & ~n121;
  assign n123 = pi3  & ~n122;
  assign n124 = ~n78 & ~n105;
  assign n125 = ~n92 & n124;
  assign n126 = ~n123 & n125;
  assign n127 = ~pi7  & ~n126;
  assign n128 = ~n70 & ~n127;
  assign n129 = ~pi4  & ~n128;
  assign n130 = ~pi1  & ~pi3 ;
  assign n131 = pi6  & ~pi9 ;
  assign n132 = pi4  & pi9 ;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~pi8  & ~n116;
  assign n135 = ~n133 & n134;
  assign n136 = pi4  & pi8 ;
  assign n137 = ~pi6  & ~pi9 ;
  assign n138 = ~n136 & ~n137;
  assign n139 = ~pi6  & pi8 ;
  assign n140 = pi5  & ~n139;
  assign n141 = ~n138 & n140;
  assign n142 = ~n135 & ~n141;
  assign n143 = ~pi7  & n112;
  assign n144 = n130 & n143;
  assign n145 = ~n142 & n144;
  assign po0  = n129 | n145;
  assign n147 = pi2  & ~n64;
  assign n148 = pi0  & pi1 ;
  assign n149 = n79 & ~n148;
  assign n150 = ~pi8  & ~n147;
  assign n151 = ~n149 & n150;
  assign n152 = ~pi2  & pi8 ;
  assign n153 = n22 & n152;
  assign n154 = ~n151 & ~n153;
  assign n155 = pi7  & ~n154;
  assign n156 = ~n65 & ~n155;
  assign n157 = ~pi6  & n27;
  assign n158 = ~pi4  & n157;
  assign n159 = ~n156 & n158;
  assign n160 = pi1  & pi2 ;
  assign n161 = pi5  & ~pi8 ;
  assign n162 = ~pi6  & ~n161;
  assign n163 = pi3  & n160;
  assign n164 = ~n162 & n163;
  assign n165 = pi1  & pi5 ;
  assign n166 = pi3  & ~pi8 ;
  assign n167 = n76 & n166;
  assign n168 = ~n165 & ~n167;
  assign n169 = pi0  & ~n168;
  assign n170 = pi5  & ~n35;
  assign n171 = ~n169 & ~n170;
  assign n172 = pi6  & ~n171;
  assign n173 = ~n164 & ~n172;
  assign n174 = pi9  & ~n173;
  assign n175 = ~pi2  & ~pi8 ;
  assign n176 = pi5  & n175;
  assign n177 = ~pi5  & pi8 ;
  assign n178 = ~n71 & ~n177;
  assign n179 = pi0  & n178;
  assign n180 = ~n176 & ~n179;
  assign n181 = ~pi1  & ~n180;
  assign n182 = ~pi0  & pi5 ;
  assign n183 = pi0  & n152;
  assign n184 = pi0  & ~pi5 ;
  assign n185 = ~n182 & ~n184;
  assign n186 = ~n183 & n185;
  assign n187 = pi1  & ~n186;
  assign n188 = ~pi0  & ~n35;
  assign n189 = ~n175 & n188;
  assign n190 = ~n187 & ~n189;
  assign n191 = ~n181 & n190;
  assign n192 = ~pi6  & ~n191;
  assign n193 = ~pi1  & pi6 ;
  assign n194 = pi2  & ~n193;
  assign n195 = ~pi1  & ~pi8 ;
  assign n196 = pi3  & ~n195;
  assign n197 = ~n194 & n196;
  assign n198 = ~pi0  & pi8 ;
  assign n199 = ~pi1  & ~pi6 ;
  assign n200 = ~pi2  & ~n148;
  assign n201 = ~n198 & ~n199;
  assign n202 = n200 & n201;
  assign n203 = ~n197 & ~n202;
  assign n204 = ~pi5  & ~n203;
  assign n205 = ~n192 & ~n204;
  assign n206 = ~pi9  & ~n205;
  assign n207 = n42 & n139;
  assign n208 = ~pi8  & ~pi9 ;
  assign n209 = pi8  & pi9 ;
  assign n210 = pi0  & n209;
  assign n211 = ~n208 & ~n210;
  assign n212 = pi5  & ~n211;
  assign n213 = ~n42 & ~n62;
  assign n214 = n212 & n213;
  assign n215 = ~pi8  & n59;
  assign n216 = pi6  & pi9 ;
  assign n217 = ~n177 & ~n216;
  assign n218 = pi6  & pi8 ;
  assign n219 = pi0  & ~n218;
  assign n220 = ~n23 & ~n217;
  assign n221 = ~n219 & n220;
  assign n222 = ~n215 & ~n221;
  assign n223 = pi2  & ~n222;
  assign n224 = ~n214 & ~n223;
  assign n225 = ~pi1  & ~n224;
  assign n226 = ~n217 & n219;
  assign n227 = ~pi8  & pi9 ;
  assign n228 = n182 & n227;
  assign n229 = ~n226 & ~n228;
  assign n230 = ~pi2  & ~n229;
  assign n231 = ~pi6  & ~pi8 ;
  assign n232 = pi2  & ~pi5 ;
  assign n233 = ~pi6  & ~n232;
  assign n234 = ~n62 & n177;
  assign n235 = ~n233 & n234;
  assign n236 = ~n231 & ~n235;
  assign n237 = ~pi9  & ~n236;
  assign n238 = ~n230 & ~n237;
  assign n239 = pi1  & ~n238;
  assign n240 = ~n207 & ~n239;
  assign n241 = ~n225 & n240;
  assign n242 = ~pi3  & ~n241;
  assign n243 = ~n174 & ~n206;
  assign n244 = ~n242 & n243;
  assign n245 = ~pi4  & ~n244;
  assign n246 = ~n136 & ~n161;
  assign n247 = ~pi6  & ~n246;
  assign n248 = ~n132 & ~n247;
  assign n249 = n114 & n130;
  assign n250 = ~n248 & n249;
  assign n251 = ~n245 & ~n250;
  assign n252 = ~pi7  & ~n251;
  assign po1  = n159 | n252;
  assign n254 = ~pi5  & n85;
  assign n255 = ~n212 & ~n254;
  assign n256 = pi1  & ~n255;
  assign n257 = ~n208 & ~n209;
  assign n258 = ~n72 & ~n257;
  assign n259 = pi2  & ~n258;
  assign n260 = ~n256 & ~n259;
  assign n261 = ~pi3  & ~n260;
  assign n262 = ~pi1  & pi8 ;
  assign n263 = n36 & n262;
  assign n264 = ~pi2  & ~pi5 ;
  assign n265 = ~n167 & ~n264;
  assign n266 = n208 & ~n265;
  assign n267 = ~n263 & ~n266;
  assign n268 = pi0  & ~n267;
  assign n269 = ~n261 & ~n268;
  assign n270 = ~pi6  & ~n269;
  assign n271 = pi6  & ~n30;
  assign n272 = ~n22 & ~n271;
  assign n273 = pi8  & ~n272;
  assign n274 = ~n75 & ~n273;
  assign n275 = ~pi2  & ~n274;
  assign n276 = pi8  & ~n42;
  assign n277 = pi2  & n73;
  assign n278 = ~n262 & ~n277;
  assign n279 = pi6  & ~n278;
  assign n280 = pi2  & n208;
  assign n281 = ~n276 & ~n280;
  assign n282 = ~n279 & n281;
  assign n283 = pi3  & ~n282;
  assign n284 = ~n275 & ~n283;
  assign n285 = n184 & ~n284;
  assign n286 = ~n270 & ~n285;
  assign n287 = ~pi4  & ~n286;
  assign n288 = ~pi3  & pi9 ;
  assign n289 = ~pi1  & ~n208;
  assign n290 = pi6  & ~n209;
  assign n291 = ~n289 & n290;
  assign n292 = n288 & n291;
  assign n293 = pi3  & ~n152;
  assign n294 = pi5  & ~n293;
  assign n295 = pi3  & ~n232;
  assign n296 = pi8  & ~n295;
  assign n297 = ~n294 & ~n296;
  assign n298 = pi1  & ~n297;
  assign n299 = ~pi5  & pi6 ;
  assign n300 = ~pi3  & n299;
  assign n301 = n195 & n300;
  assign n302 = ~n298 & ~n301;
  assign n303 = ~pi9  & ~n302;
  assign n304 = pi6  & ~pi8 ;
  assign n305 = ~pi9  & ~n193;
  assign n306 = ~n304 & n305;
  assign n307 = ~pi2  & ~n306;
  assign n308 = ~pi8  & n30;
  assign n309 = ~n307 & ~n308;
  assign n310 = pi3  & ~n309;
  assign n311 = pi2  & ~n139;
  assign n312 = ~n262 & ~n311;
  assign n313 = n170 & ~n312;
  assign n314 = ~n40 & ~n227;
  assign n315 = ~pi6  & ~n288;
  assign n316 = ~n314 & n315;
  assign n317 = ~n292 & ~n316;
  assign n318 = ~n313 & n317;
  assign n319 = ~n310 & n318;
  assign n320 = ~n303 & n319;
  assign n321 = ~pi4  & ~n320;
  assign n322 = ~n209 & ~n304;
  assign n323 = ~pi5  & ~n322;
  assign n324 = ~pi3  & pi4 ;
  assign n325 = n76 & n324;
  assign n326 = ~n323 & n325;
  assign n327 = ~n321 & ~n326;
  assign n328 = ~pi0  & ~n327;
  assign n329 = ~n287 & ~n328;
  assign n330 = ~pi7  & ~n329;
  assign n331 = n23 & n195;
  assign n332 = pi0  & ~n53;
  assign n333 = n81 & ~n332;
  assign n334 = ~n331 & ~n333;
  assign n335 = ~pi2  & n158;
  assign n336 = ~n334 & n335;
  assign po2  = n330 | n336;
  assign n338 = n299 & n306;
  assign n339 = n176 & n199;
  assign n340 = ~n300 & ~n339;
  assign n341 = ~pi9  & ~n340;
  assign n342 = pi2  & ~n178;
  assign n343 = pi8  & n44;
  assign n344 = ~n342 & ~n343;
  assign n345 = ~pi9  & ~n344;
  assign n346 = ~pi6  & ~n166;
  assign n347 = pi3  & ~pi5 ;
  assign n348 = ~n346 & ~n347;
  assign n349 = ~pi2  & pi3 ;
  assign n350 = pi9  & n176;
  assign n351 = ~n348 & ~n349;
  assign n352 = ~n350 & n351;
  assign n353 = ~n345 & n352;
  assign n354 = pi1  & ~n353;
  assign n355 = ~n341 & ~n354;
  assign n356 = pi0  & ~n355;
  assign n357 = ~pi8  & n299;
  assign n358 = pi5  & pi8 ;
  assign n359 = n113 & n358;
  assign n360 = ~n215 & ~n359;
  assign n361 = pi2  & ~n360;
  assign n362 = pi3  & ~n348;
  assign n363 = ~n357 & ~n361;
  assign n364 = ~n362 & n363;
  assign n365 = pi1  & ~n364;
  assign n366 = pi2  & n299;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~pi0  & ~n367;
  assign n369 = ~n59 & ~n231;
  assign n370 = ~pi2  & ~n369;
  assign n371 = pi5  & pi9 ;
  assign n372 = ~pi6  & ~n371;
  assign n373 = ~n73 & ~n358;
  assign n374 = n372 & ~n373;
  assign n375 = ~n370 & ~n374;
  assign n376 = pi3  & ~n375;
  assign n377 = pi2  & n98;
  assign n378 = ~n299 & ~n377;
  assign n379 = n36 & ~n378;
  assign n380 = ~pi5  & ~pi6 ;
  assign n381 = ~n116 & ~n380;
  assign n382 = ~pi6  & ~n209;
  assign n383 = ~n381 & ~n382;
  assign n384 = n217 & ~n346;
  assign n385 = ~n383 & n384;
  assign n386 = ~n379 & ~n385;
  assign n387 = ~pi1  & ~n386;
  assign n388 = ~n338 & ~n376;
  assign n389 = ~n387 & n388;
  assign n390 = ~n356 & n389;
  assign n391 = ~n368 & n390;
  assign n392 = ~pi4  & ~n391;
  assign n393 = pi3  & ~n113;
  assign n394 = pi2  & pi6 ;
  assign n395 = ~n393 & ~n394;
  assign n396 = ~pi4  & ~n395;
  assign n397 = ~pi2  & n324;
  assign n398 = n383 & n397;
  assign n399 = ~n396 & ~n398;
  assign n400 = n64 & ~n399;
  assign n401 = ~n392 & ~n400;
  assign po3  = ~pi7  & ~n401;
  assign n403 = ~pi4  & n147;
  assign n404 = pi3  & ~pi4 ;
  assign n405 = ~n324 & ~n404;
  assign n406 = n77 & ~n405;
  assign n407 = ~n403 & ~n406;
  assign n408 = ~pi7  & n116;
  assign po4  = ~n407 & n408;
  assign n410 = ~n77 & n404;
  assign n411 = n64 & n397;
  assign n412 = ~n410 & ~n411;
  assign po5  = n408 & ~n412;
  assign n414 = pi7  & ~pi9 ;
  assign n415 = pi8  & ~n414;
  assign n416 = n108 & ~n415;
  assign n417 = ~n86 & ~n416;
  assign n418 = ~pi0  & ~n417;
  assign n419 = ~pi2  & pi7 ;
  assign n420 = ~n262 & n419;
  assign n421 = ~n211 & n420;
  assign n422 = ~n418 & ~n421;
  assign n423 = n380 & ~n422;
  assign n424 = ~pi8  & n72;
  assign n425 = pi2  & n28;
  assign n426 = ~n424 & ~n425;
  assign n427 = pi5  & ~n426;
  assign n428 = ~pi1  & ~pi5 ;
  assign n429 = pi2  & ~n428;
  assign n430 = n137 & ~n429;
  assign n431 = pi5  & n73;
  assign n432 = ~n430 & ~n431;
  assign n433 = pi0  & ~n432;
  assign n434 = ~pi0  & pi2 ;
  assign n435 = ~n59 & n434;
  assign n436 = ~n433 & ~n435;
  assign n437 = pi8  & ~n436;
  assign n438 = pi6  & ~n257;
  assign n439 = pi2  & pi8 ;
  assign n440 = ~n175 & ~n439;
  assign n441 = n438 & ~n440;
  assign n442 = ~n427 & ~n441;
  assign n443 = ~n437 & n442;
  assign n444 = ~pi7  & ~n443;
  assign n445 = ~n423 & ~n444;
  assign n446 = ~pi3  & ~n445;
  assign n447 = ~pi0  & ~pi6 ;
  assign n448 = pi8  & ~n184;
  assign n449 = ~pi2  & ~pi9 ;
  assign n450 = ~n447 & n449;
  assign n451 = ~n448 & n450;
  assign n452 = pi8  & n425;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~pi1  & ~n453;
  assign n455 = n41 & ~n289;
  assign n456 = ~n195 & n447;
  assign n457 = ~n160 & ~n456;
  assign n458 = n74 & ~n457;
  assign n459 = ~n455 & ~n458;
  assign n460 = ~pi5  & ~n459;
  assign n461 = pi0  & n218;
  assign n462 = ~n93 & ~n461;
  assign n463 = ~pi2  & ~n462;
  assign n464 = ~pi8  & n148;
  assign n465 = ~n463 & ~n464;
  assign n466 = pi9  & ~n465;
  assign n467 = ~pi0  & ~pi8 ;
  assign n468 = n22 & ~n184;
  assign n469 = ~n467 & n468;
  assign n470 = ~n460 & ~n469;
  assign n471 = ~n466 & n470;
  assign n472 = pi3  & ~n471;
  assign n473 = n28 & ~n233;
  assign n474 = ~n45 & ~n473;
  assign n475 = ~pi8  & ~n474;
  assign n476 = pi2  & ~n208;
  assign n477 = ~n210 & ~n476;
  assign n478 = pi6  & ~n477;
  assign n479 = ~n475 & ~n478;
  assign n480 = pi1  & ~n479;
  assign n481 = ~n454 & ~n480;
  assign n482 = ~n472 & n481;
  assign n483 = ~pi7  & ~n482;
  assign n484 = ~n446 & ~n483;
  assign n485 = ~pi4  & ~n484;
  assign n486 = ~n116 & ~n411;
  assign n487 = ~pi7  & ~n486;
  assign po6  = ~n485 & ~n487;
  assign n489 = n349 & n441;
  assign n490 = ~pi6  & ~n71;
  assign n491 = n476 & ~n490;
  assign n492 = ~pi0  & n438;
  assign n493 = n79 & n382;
  assign n494 = ~n492 & ~n493;
  assign n495 = pi3  & ~n494;
  assign n496 = ~pi0  & n175;
  assign n497 = ~n461 & ~n496;
  assign n498 = ~pi9  & ~n497;
  assign n499 = ~pi1  & ~n491;
  assign n500 = ~n498 & n499;
  assign n501 = ~n495 & n500;
  assign n502 = n71 & n137;
  assign n503 = n98 & n198;
  assign n504 = ~n304 & ~n503;
  assign n505 = pi9  & ~n504;
  assign n506 = ~n88 & n490;
  assign n507 = ~n505 & n506;
  assign n508 = ~pi3  & n209;
  assign n509 = pi2  & ~n508;
  assign n510 = ~n507 & n509;
  assign n511 = ~pi3  & pi8 ;
  assign n512 = ~n216 & ~n511;
  assign n513 = pi0  & ~n512;
  assign n514 = pi8  & n131;
  assign n515 = ~pi2  & ~n514;
  assign n516 = ~n513 & n515;
  assign n517 = ~n505 & n516;
  assign n518 = ~n510 & ~n517;
  assign n519 = pi1  & ~n502;
  assign n520 = ~n518 & n519;
  assign n521 = ~n501 & ~n520;
  assign n522 = ~n489 & ~n521;
  assign n523 = ~pi5  & ~n522;
  assign n524 = pi8  & n371;
  assign n525 = n99 & n524;
  assign n526 = n85 & n161;
  assign n527 = ~pi0  & ~n440;
  assign n528 = ~n183 & ~n527;
  assign n529 = ~pi9  & ~n528;
  assign n530 = pi8  & ~n213;
  assign n531 = ~n529 & n530;
  assign n532 = ~n526 & ~n531;
  assign n533 = ~pi3  & ~n532;
  assign n534 = pi3  & pi5 ;
  assign n535 = ~n42 & ~n534;
  assign n536 = n467 & ~n535;
  assign n537 = pi8  & n88;
  assign n538 = ~n349 & ~n537;
  assign n539 = pi5  & ~n209;
  assign n540 = ~n538 & n539;
  assign n541 = pi1  & ~n536;
  assign n542 = ~n540 & n541;
  assign n543 = ~n533 & n542;
  assign n544 = ~n112 & ~n257;
  assign n545 = ~n99 & ~n544;
  assign n546 = n170 & ~n545;
  assign n547 = n37 & n280;
  assign n548 = ~pi1  & ~n547;
  assign n549 = ~n546 & n548;
  assign n550 = ~n543 & ~n549;
  assign n551 = ~n525 & ~n550;
  assign n552 = ~pi6  & ~n551;
  assign n553 = ~n523 & ~n552;
  assign n554 = ~pi7  & ~n553;
  assign n555 = ~pi8  & n425;
  assign n556 = ~n529 & ~n555;
  assign n557 = ~pi2  & ~n53;
  assign n558 = n130 & n380;
  assign n559 = ~n557 & n558;
  assign n560 = ~n556 & n559;
  assign n561 = ~n554 & ~n560;
  assign n562 = ~pi4  & ~n561;
  assign n563 = ~pi5  & ~pi7 ;
  assign n564 = n411 & n563;
  assign n565 = ~pi6  & n564;
  assign po7  = ~n562 & ~n565;
  assign n567 = n74 & ~n428;
  assign n568 = n94 & ~n567;
  assign n569 = ~n165 & ~n347;
  assign n570 = ~pi2  & ~n72;
  assign n571 = ~n288 & n570;
  assign n572 = n569 & n571;
  assign n573 = ~n29 & ~n108;
  assign n574 = ~n48 & n573;
  assign n575 = ~n568 & ~n572;
  assign n576 = ~n574 & n575;
  assign n577 = ~pi8  & ~n576;
  assign n578 = n130 & n184;
  assign n579 = ~pi2  & ~n88;
  assign n580 = n569 & n579;
  assign n581 = ~n578 & ~n580;
  assign n582 = pi8  & ~n581;
  assign n583 = pi2  & ~n184;
  assign n584 = n298 & n583;
  assign n585 = ~n582 & ~n584;
  assign n586 = ~pi9  & ~n585;
  assign n587 = ~n232 & ~n534;
  assign n588 = pi1  & ~n293;
  assign n589 = ~n587 & n588;
  assign n590 = n76 & ~n182;
  assign n591 = n196 & n590;
  assign n592 = ~n589 & ~n591;
  assign n593 = pi9  & ~n592;
  assign n594 = ~n586 & ~n593;
  assign n595 = ~n577 & n594;
  assign n596 = ~pi6  & ~n595;
  assign n597 = pi2  & ~n289;
  assign n598 = ~n271 & ~n597;
  assign n599 = pi0  & ~n598;
  assign n600 = ~n199 & n311;
  assign n601 = ~n291 & ~n600;
  assign n602 = ~n599 & n601;
  assign n603 = n347 & ~n602;
  assign n604 = ~n596 & ~n603;
  assign n605 = ~pi7  & ~n604;
  assign n606 = ~pi1  & ~n556;
  assign n607 = n73 & n496;
  assign n608 = ~n606 & ~n607;
  assign n609 = n157 & ~n608;
  assign n610 = ~n605 & ~n609;
  assign n611 = ~pi4  & ~n610;
  assign po8  = ~n564 & ~n611;
  assign n613 = ~pi2  & n130;
  assign n614 = pi4  & ~n613;
  assign n615 = ~pi3  & ~n59;
  assign n616 = n198 & ~n512;
  assign n617 = ~n615 & ~n616;
  assign n618 = ~pi2  & ~n617;
  assign n619 = ~pi6  & ~n524;
  assign n620 = ~pi3  & ~n619;
  assign n621 = ~pi5  & ~n209;
  assign n622 = n377 & n621;
  assign n623 = ~n620 & ~n622;
  assign n624 = ~n618 & n623;
  assign n625 = pi1  & ~n624;
  assign n626 = n324 & ~n380;
  assign n627 = n198 & ~n372;
  assign n628 = pi3  & ~n216;
  assign n629 = ~n627 & n628;
  assign n630 = ~pi2  & ~n626;
  assign n631 = ~n629 & n630;
  assign n632 = n476 & n615;
  assign n633 = ~n297 & n632;
  assign n634 = ~n631 & ~n633;
  assign n635 = ~pi1  & ~n634;
  assign n636 = n184 & n377;
  assign n637 = ~pi7  & ~n636;
  assign n638 = ~n289 & ~n637;
  assign n639 = pi7  & ~n94;
  assign n640 = ~pi7  & ~n613;
  assign n641 = pi0  & ~n640;
  assign n642 = ~pi5  & ~n94;
  assign n643 = pi6  & ~n642;
  assign n644 = ~n614 & ~n639;
  assign n645 = ~n643 & n644;
  assign n646 = ~n641 & n645;
  assign n647 = ~n638 & n646;
  assign n648 = ~n625 & n647;
  assign po9  = ~n635 & n648;
  assign n650 = pi8  & ~n29;
  assign n651 = pi2  & n404;
  assign n652 = ~n24 & n651;
  assign n653 = ~n650 & n652;
  assign n654 = ~n411 & ~n653;
  assign n655 = ~pi7  & n380;
  assign po10  = ~n654 & n655;
endmodule
