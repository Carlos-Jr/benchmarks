module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 ,
    po6 , po7 , po8 , po9 , po10 ,
    po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 ,
    po21 , po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 , po30 ,
    po31 , po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 ,
    po46 , po47 , po48 , po49 , po50 ,
    po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 ,
    po61 , po62 , po63   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 ;
  wire n194, n195, n196, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244,
    n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330,
    n331, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n713, n714,
    n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925,
    n926, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474,
    n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492,
    n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552,
    n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582,
    n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612,
    n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661,
    n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721,
    n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751,
    n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781,
    n1782, n1783, n1784, n1785, n1786, n1787,
    n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962,
    n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101,
    n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131,
    n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554,
    n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566,
    n2567, n2568, n2569, n2570, n2571, n2572,
    n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596,
    n2597, n2598, n2599, n2600, n2601, n2602,
    n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614,
    n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2688, n2689, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716,
    n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734,
    n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752,
    n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771,
    n2772, n2773, n2774, n2775, n2776, n2777,
    n2778, n2779, n2780, n2781, n2782, n2783,
    n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801,
    n2802, n2803, n2804, n2805, n2806, n2807,
    n2808, n2809, n2810, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831,
    n2832, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861,
    n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885,
    n2886, n2887, n2888, n2889, n2890, n2891,
    n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915,
    n2916, n2917, n2918, n2919, n2920, n2921,
    n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933,
    n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211,
    n3212, n3213, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241,
    n3242, n3243, n3244, n3245, n3246, n3247,
    n3248, n3249, n3250, n3251, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271,
    n3272, n3273, n3274, n3275, n3276, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3441, n3442, n3443, n3444, n3445, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476,
    n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927,
    n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156,
    n4157, n4158, n4159, n4160, n4161, n4162,
    n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174,
    n4175, n4176, n4177, n4178, n4179, n4180,
    n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192,
    n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204,
    n4205, n4206, n4207, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277,
    n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307,
    n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367,
    n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385,
    n4386, n4387, n4388, n4389, n4390, n4391,
    n4392, n4393, n4394, n4395, n4396, n4397,
    n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4421,
    n4422, n4423, n4424, n4425, n4426, n4427,
    n4428, n4429, n4430, n4431, n4432, n4433,
    n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451,
    n4452, n4453, n4454, n4455, n4456, n4457,
    n4458, n4459, n4460, n4461, n4462, n4463,
    n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596,
    n4597, n4598, n4599, n4600, n4601, n4602,
    n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662,
    n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686,
    n4687, n4688, n4689, n4690, n4691, n4692,
    n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710,
    n4711, n4712, n4713, n4714, n4715, n4716,
    n4717, n4718, n4719, n4720, n4721, n4722,
    n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734,
    n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752,
    n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764,
    n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843,
    n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861,
    n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873,
    n4874, n4875, n4876, n4877, n4878, n4879,
    n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891,
    n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072,
    n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5359, n5360, n5361,
    n5362, n5363, n5364, n5365, n5366, n5367,
    n5368, n5369, n5370, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391,
    n5392, n5393, n5394, n5395, n5396, n5397,
    n5398, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409,
    n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421,
    n5422, n5423, n5424, n5425, n5426, n5427,
    n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451,
    n5452, n5453, n5454, n5455, n5456, n5457,
    n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481,
    n5482, n5483, n5484, n5485, n5486, n5487,
    n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499,
    n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511,
    n5512, n5513, n5514, n5515, n5516, n5517,
    n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541,
    n5542, n5543, n5544, n5545, n5546, n5547,
    n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571,
    n5572, n5573, n5574, n5575, n5576, n5577,
    n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601,
    n5602, n5603, n5604, n5605, n5606, n5607,
    n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619,
    n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631,
    n5632, n5633, n5634, n5635, n5636, n5637,
    n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649,
    n5650, n5651, n5652, n5653, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661,
    n5662, n5663, n5664, n5665, n5666, n5667,
    n5669, n5670, n5671, n5672, n5673, n5674,
    n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5684, n5685, n5686,
    n5687, n5688, n5689, n5690, n5691, n5692,
    n5693, n5694, n5695, n5696, n5697, n5698,
    n5699, n5700, n5701, n5702, n5703, n5704,
    n5705, n5706, n5707, n5708, n5709, n5710,
    n5711, n5712, n5713, n5714, n5715, n5716,
    n5717, n5718, n5719, n5720, n5721, n5722,
    n5723, n5724, n5725, n5726, n5727, n5728,
    n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740,
    n5741, n5742, n5743, n5744, n5745, n5746,
    n5747, n5748, n5749, n5750, n5751, n5752,
    n5753, n5754, n5755, n5756, n5757, n5758,
    n5759, n5760, n5761, n5762, n5763, n5764,
    n5765, n5766, n5767, n5768, n5769, n5770,
    n5771, n5772, n5773, n5774, n5775, n5776,
    n5777, n5778, n5779, n5780, n5781, n5782,
    n5783, n5784, n5785, n5786, n5787, n5788,
    n5789, n5790, n5791, n5792, n5793, n5794,
    n5795, n5796, n5797, n5798, n5799, n5800,
    n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5812,
    n5813, n5814, n5815, n5816, n5817, n5818,
    n5819, n5820, n5821, n5822, n5823, n5824,
    n5825, n5826, n5827, n5828, n5829, n5830,
    n5831, n5832, n5833, n5834, n5835, n5836,
    n5837, n5838, n5839, n5840, n5841, n5842,
    n5843, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854,
    n5855, n5856, n5857, n5858, n5859, n5860,
    n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872,
    n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884,
    n5885, n5886, n5887, n5888, n5889, n5890,
    n5891, n5892, n5893, n5894, n5895, n5896,
    n5897, n5898, n5899, n5900, n5901, n5902,
    n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914,
    n5915, n5916, n5917, n5918, n5919, n5920,
    n5921, n5922, n5923, n5924, n5925, n5926,
    n5927, n5928, n5929, n5930, n5931, n5932,
    n5933, n5934, n5935, n5936, n5937, n5938,
    n5939, n5940, n5941, n5942, n5943, n5944,
    n5945, n5946, n5947, n5948, n5949, n5950,
    n5951, n5952, n5953, n5954, n5955, n5956,
    n5957, n5958, n5959, n5960, n5961, n5962,
    n5963, n5964, n5965, n5966, n5967, n5968,
    n5969, n5970, n5971, n5972, n5973, n5974,
    n5975, n5976, n5977, n5978, n5979, n5980,
    n5981, n5982, n5983, n5984, n5985, n5986,
    n5988, n5989, n5990, n5991, n5992, n5993,
    n5994, n5995, n5996, n5997, n5998, n5999,
    n6000, n6001, n6002, n6003, n6004, n6005,
    n6006, n6007, n6008, n6009, n6010, n6011,
    n6012, n6013, n6014, n6015, n6016, n6017,
    n6018, n6019, n6020, n6021, n6022, n6023,
    n6024, n6025, n6026, n6027, n6028, n6029,
    n6030, n6031, n6032, n6033, n6034, n6035,
    n6036, n6037, n6038, n6039, n6040, n6041,
    n6042, n6043, n6044, n6045, n6046, n6047,
    n6048, n6049, n6050, n6051, n6052, n6053,
    n6054, n6055, n6056, n6057, n6058, n6059,
    n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071,
    n6072, n6073, n6074, n6075, n6076, n6077,
    n6078, n6079, n6080, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087, n6088, n6089,
    n6090, n6091, n6092, n6093, n6094, n6095,
    n6096, n6097, n6098, n6099, n6100, n6101,
    n6102, n6103, n6104, n6105, n6106, n6107,
    n6108, n6109, n6110, n6111, n6112, n6113,
    n6114, n6115, n6116, n6117, n6118, n6119,
    n6120, n6121, n6122, n6123, n6124, n6125,
    n6126, n6127, n6128, n6129, n6130, n6131,
    n6132, n6133, n6134, n6135, n6136, n6137,
    n6138, n6139, n6140, n6141, n6142, n6143,
    n6144, n6145, n6146, n6147, n6148, n6149,
    n6150, n6151, n6152, n6153, n6154, n6155,
    n6156, n6157, n6158, n6159, n6160, n6161,
    n6162, n6163, n6164, n6165, n6166, n6167,
    n6168, n6169, n6170, n6171, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6179,
    n6180, n6181, n6182, n6183, n6184, n6185,
    n6186, n6187, n6188, n6189, n6190, n6191,
    n6192, n6193, n6194, n6195, n6196, n6197,
    n6198, n6199, n6200, n6201, n6202, n6203,
    n6204, n6205, n6206, n6207, n6208, n6209,
    n6210, n6211, n6212, n6213, n6214, n6215,
    n6216, n6217, n6218, n6219, n6220, n6221,
    n6222, n6223, n6224, n6225, n6226, n6227,
    n6228, n6229, n6230, n6231, n6232, n6233,
    n6234, n6235, n6236, n6237, n6238, n6239,
    n6240, n6241, n6242, n6243, n6244, n6245,
    n6246, n6247, n6248, n6249, n6250, n6251,
    n6252, n6253, n6254, n6255, n6256, n6257,
    n6258, n6259, n6260, n6261, n6262, n6263,
    n6264, n6265, n6266, n6267, n6268, n6269,
    n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6277, n6278, n6279, n6280, n6281,
    n6282, n6283, n6284, n6285, n6286, n6287,
    n6288, n6289, n6290, n6291, n6292, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311,
    n6312, n6313, n6314, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546,
    n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570,
    n6571, n6572, n6573, n6574, n6575, n6576,
    n6577, n6578, n6579, n6580, n6581, n6582,
    n6583, n6584, n6585, n6586, n6587, n6588,
    n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600,
    n6601, n6602, n6603, n6604, n6605, n6606,
    n6607, n6608, n6609, n6610, n6611, n6612,
    n6613, n6614, n6615, n6616, n6617, n6618,
    n6619, n6620, n6621, n6622, n6623, n6624,
    n6625, n6626, n6627, n6628, n6629, n6630,
    n6631, n6632, n6633, n6634, n6635, n6636,
    n6637, n6638, n6639, n6640, n6641, n6642,
    n6643, n6644, n6645, n6646, n6647, n6648,
    n6649, n6650, n6651, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661,
    n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691,
    n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721,
    n6722, n6723, n6724, n6725, n6726, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751,
    n6752, n6753, n6754, n6755, n6756, n6757,
    n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781,
    n6782, n6783, n6784, n6785, n6786, n6787,
    n6788, n6789, n6790, n6791, n6792, n6793,
    n6794, n6795, n6796, n6797, n6798, n6799,
    n6800, n6801, n6802, n6803, n6804, n6805,
    n6806, n6807, n6808, n6809, n6810, n6811,
    n6812, n6813, n6814, n6815, n6816, n6817,
    n6818, n6819, n6820, n6821, n6822, n6823,
    n6824, n6825, n6826, n6827, n6828, n6829,
    n6830, n6831, n6832, n6833, n6834, n6835,
    n6836, n6837, n6838, n6839, n6840, n6841,
    n6842, n6843, n6844, n6845, n6846, n6847,
    n6848, n6849, n6850, n6851, n6852, n6853,
    n6854, n6855, n6856, n6857, n6858, n6859,
    n6860, n6861, n6862, n6863, n6864, n6865,
    n6866, n6867, n6868, n6869, n6870, n6871,
    n6872, n6873, n6874, n6875, n6876, n6877,
    n6878, n6879, n6880, n6881, n6882, n6883,
    n6884, n6885, n6886, n6887, n6888, n6889,
    n6890, n6891, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901,
    n6902, n6903, n6904, n6905, n6906, n6907,
    n6908, n6909, n6910, n6911, n6912, n6913,
    n6914, n6915, n6916, n6917, n6918, n6919,
    n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931,
    n6932, n6933, n6934, n6935, n6936, n6937,
    n6938, n6939, n6940, n6941, n6942, n6943,
    n6944, n6945, n6946, n6947, n6948, n6949,
    n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961,
    n6962, n6963, n6964, n6965, n6966, n6967,
    n6968, n6969, n6970, n6971, n6972, n6973,
    n6974, n6975, n6976, n6977, n6978, n6979,
    n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991,
    n6992, n6993, n6994, n6995, n6996, n6997,
    n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112,
    n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136,
    n7137, n7138, n7139, n7140, n7141, n7142,
    n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154,
    n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172,
    n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214,
    n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352,
    n7354, n7355, n7356, n7357, n7358, n7359,
    n7360, n7361, n7362, n7363, n7364, n7365,
    n7366, n7367, n7368, n7369, n7370, n7371,
    n7372, n7373, n7374, n7375, n7376, n7377,
    n7378, n7379, n7380, n7381, n7382, n7383,
    n7384, n7385, n7386, n7387, n7388, n7389,
    n7390, n7391, n7392, n7393, n7394, n7395,
    n7396, n7397, n7398, n7399, n7400, n7401,
    n7402, n7403, n7404, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431,
    n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443,
    n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461,
    n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479,
    n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491,
    n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503,
    n7504, n7505, n7506, n7507, n7508, n7509,
    n7510, n7511, n7512, n7513, n7514, n7515,
    n7516, n7517, n7518, n7519, n7520, n7521,
    n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551,
    n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581,
    n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7716, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726,
    n7727, n7728, n7729, n7730, n7731, n7732,
    n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744,
    n7745, n7746, n7747, n7748, n7749, n7750,
    n7751, n7752, n7753, n7754, n7755, n7756,
    n7757, n7758, n7759, n7760, n7761, n7762,
    n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7786,
    n7787, n7788, n7789, n7790, n7791, n7792,
    n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7813, n7814, n7815, n7816,
    n7817, n7818, n7819, n7820, n7821, n7822,
    n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062,
    n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8091, n8092, n8093,
    n8094, n8095, n8096, n8097, n8098, n8099,
    n8100, n8101, n8102, n8103, n8104, n8105,
    n8106, n8107, n8108, n8109, n8110, n8111,
    n8112, n8113, n8114, n8115, n8116, n8117,
    n8118, n8119, n8120, n8121, n8122, n8123,
    n8124, n8125, n8126, n8127, n8128, n8129,
    n8130, n8131, n8132, n8133, n8134, n8135,
    n8136, n8137, n8138, n8139, n8140, n8141,
    n8142, n8143, n8144, n8145, n8146, n8147,
    n8148, n8149, n8150, n8151, n8152, n8153,
    n8154, n8155, n8156, n8157, n8158, n8159,
    n8160, n8161, n8162, n8163, n8164, n8165,
    n8166, n8167, n8168, n8169, n8170, n8171,
    n8172, n8173, n8174, n8175, n8176, n8177,
    n8178, n8179, n8180, n8181, n8182, n8183,
    n8184, n8185, n8186, n8187, n8188, n8189,
    n8190, n8191, n8192, n8193, n8194, n8195,
    n8196, n8197, n8198, n8199, n8200, n8201,
    n8202, n8203, n8204, n8205, n8206, n8207,
    n8208, n8209, n8210, n8211, n8212, n8213,
    n8214, n8215, n8216, n8217, n8218, n8219,
    n8220, n8221, n8222, n8223, n8224, n8225,
    n8226, n8227, n8228, n8229, n8230, n8231,
    n8232, n8233, n8234, n8235, n8236, n8237,
    n8238, n8239, n8240, n8241, n8242, n8243,
    n8244, n8245, n8246, n8247, n8248, n8249,
    n8250, n8251, n8252, n8253, n8254, n8255,
    n8256, n8257, n8258, n8259, n8260, n8261,
    n8262, n8263, n8264, n8265, n8266, n8267,
    n8268, n8269, n8270, n8271, n8272, n8273,
    n8274, n8275, n8276, n8277, n8278, n8279,
    n8280, n8281, n8282, n8283, n8284, n8285,
    n8286, n8287, n8288, n8289, n8290, n8291,
    n8292, n8293, n8294, n8295, n8296, n8297,
    n8298, n8299, n8300, n8301, n8302, n8303,
    n8304, n8305, n8306, n8307, n8308, n8309,
    n8310, n8311, n8312, n8313, n8314, n8315,
    n8316, n8317, n8318, n8319, n8320, n8321,
    n8322, n8323, n8324, n8325, n8326, n8327,
    n8328, n8329, n8330, n8331, n8332, n8333,
    n8334, n8335, n8336, n8337, n8338, n8339,
    n8340, n8341, n8342, n8343, n8344, n8345,
    n8346, n8347, n8348, n8349, n8350, n8351,
    n8352, n8353, n8354, n8355, n8356, n8357,
    n8358, n8359, n8360, n8361, n8362, n8363,
    n8364, n8365, n8366, n8367, n8368, n8369,
    n8370, n8371, n8372, n8373, n8374, n8375,
    n8376, n8377, n8378, n8379, n8380, n8381,
    n8382, n8383, n8384, n8385, n8386, n8387,
    n8388, n8389, n8390, n8391, n8392, n8393,
    n8394, n8395, n8396, n8397, n8398, n8399,
    n8400, n8401, n8402, n8403, n8404, n8405,
    n8406, n8407, n8408, n8409, n8410, n8411,
    n8412, n8413, n8414, n8415, n8416, n8417,
    n8418, n8419, n8420, n8421, n8422, n8423,
    n8424, n8425, n8426, n8427, n8428, n8429,
    n8430, n8431, n8432, n8433, n8434, n8435,
    n8436, n8437, n8438, n8439, n8440, n8441,
    n8442, n8443, n8444, n8445, n8446, n8447,
    n8448, n8449, n8450, n8451, n8452, n8453,
    n8454, n8455, n8456, n8457, n8458, n8459,
    n8460, n8461, n8462, n8463, n8464, n8465,
    n8466, n8467, n8468, n8469, n8470, n8471,
    n8473, n8474, n8475, n8476, n8477, n8478,
    n8479, n8480, n8481, n8482, n8483, n8484,
    n8485, n8486, n8487, n8488, n8489, n8490,
    n8491, n8492, n8493, n8494, n8495, n8496,
    n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508,
    n8509, n8510, n8511, n8512, n8513, n8514,
    n8515, n8516, n8517, n8518, n8519, n8520,
    n8521, n8522, n8523, n8524, n8525, n8526,
    n8527, n8528, n8529, n8530, n8531, n8532,
    n8533, n8534, n8535, n8536, n8537, n8538,
    n8539, n8540, n8541, n8542, n8543, n8544,
    n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556,
    n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568,
    n8569, n8570, n8571, n8572, n8573, n8574,
    n8575, n8576, n8577, n8578, n8579, n8580,
    n8581, n8582, n8583, n8584, n8585, n8586,
    n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8601, n8602, n8603, n8604,
    n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616,
    n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658,
    n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8678, n8679, n8680, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688,
    n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706,
    n8707, n8708, n8709, n8710, n8711, n8712,
    n8713, n8714, n8715, n8716, n8717, n8718,
    n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736,
    n8737, n8738, n8739, n8740, n8741, n8742,
    n8743, n8744, n8745, n8746, n8747, n8748,
    n8749, n8750, n8751, n8752, n8753, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766,
    n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778,
    n8779, n8780, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796,
    n8797, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826,
    n8827, n8828, n8829, n8830, n8831, n8832,
    n8833, n8834, n8835, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844,
    n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856,
    n8857, n8858, n8859, n8860, n8861, n8862,
    n8864, n8865, n8866, n8867, n8868, n8869,
    n8870, n8871, n8872, n8873, n8874, n8875,
    n8876, n8877, n8878, n8879, n8880, n8881,
    n8882, n8883, n8884, n8885, n8886, n8887,
    n8888, n8889, n8890, n8891, n8892, n8893,
    n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8908, n8909, n8910, n8911,
    n8912, n8913, n8914, n8915, n8916, n8917,
    n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8929,
    n8930, n8931, n8932, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941,
    n8942, n8943, n8944, n8945, n8946, n8947,
    n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959,
    n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971,
    n8972, n8973, n8974, n8975, n8976, n8977,
    n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001,
    n9002, n9003, n9004, n9005, n9006, n9007,
    n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019,
    n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031,
    n9032, n9033, n9034, n9035, n9036, n9037,
    n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121,
    n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151,
    n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9262, n9264, n9265, n9266,
    n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296,
    n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326,
    n9327, n9328, n9329, n9330, n9331, n9332,
    n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386,
    n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416,
    n9417, n9418, n9419, n9420, n9421, n9422,
    n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446,
    n9447, n9448, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9673, n9674, n9675,
    n9676, n9677, n9678, n9679, n9680, n9681,
    n9682, n9683, n9684, n9685, n9686, n9687,
    n9688, n9689, n9690, n9691, n9692, n9693,
    n9694, n9695, n9696, n9697, n9698, n9699,
    n9700, n9701, n9702, n9703, n9704, n9705,
    n9706, n9707, n9708, n9709, n9710, n9711,
    n9712, n9713, n9714, n9715, n9716, n9717,
    n9718, n9719, n9720, n9721, n9722, n9723,
    n9724, n9725, n9726, n9727, n9728, n9729,
    n9730, n9731, n9732, n9733, n9734, n9735,
    n9736, n9737, n9738, n9739, n9740, n9741,
    n9742, n9743, n9744, n9745, n9746, n9747,
    n9748, n9749, n9750, n9751, n9752, n9753,
    n9754, n9755, n9756, n9757, n9758, n9759,
    n9760, n9761, n9762, n9763, n9764, n9765,
    n9766, n9767, n9768, n9769, n9770, n9771,
    n9772, n9773, n9774, n9775, n9776, n9777,
    n9778, n9779, n9780, n9781, n9782, n9783,
    n9784, n9785, n9786, n9787, n9788, n9789,
    n9790, n9791, n9792, n9793, n9794, n9795,
    n9796, n9797, n9798, n9799, n9800, n9801,
    n9802, n9803, n9804, n9805, n9806, n9807,
    n9808, n9809, n9810, n9811, n9812, n9813,
    n9814, n9815, n9816, n9817, n9818, n9819,
    n9820, n9821, n9822, n9823, n9824, n9825,
    n9826, n9827, n9828, n9829, n9830, n9831,
    n9832, n9833, n9834, n9835, n9836, n9837,
    n9838, n9839, n9840, n9841, n9842, n9843,
    n9844, n9845, n9846, n9847, n9848, n9849,
    n9850, n9851, n9852, n9853, n9854, n9855,
    n9856, n9857, n9858, n9859, n9860, n9861,
    n9862, n9863, n9864, n9865, n9866, n9867,
    n9868, n9869, n9870, n9871, n9872, n9873,
    n9874, n9875, n9876, n9877, n9878, n9879,
    n9880, n9881, n9882, n9883, n9884, n9885,
    n9886, n9887, n9888, n9889, n9890, n9891,
    n9892, n9893, n9894, n9895, n9896, n9897,
    n9898, n9899, n9900, n9901, n9902, n9903,
    n9904, n9905, n9906, n9907, n9908, n9909,
    n9910, n9911, n9912, n9913, n9914, n9915,
    n9916, n9917, n9918, n9919, n9920, n9921,
    n9922, n9923, n9924, n9925, n9926, n9927,
    n9928, n9929, n9930, n9931, n9932, n9933,
    n9934, n9935, n9936, n9937, n9938, n9939,
    n9940, n9941, n9942, n9943, n9944, n9945,
    n9946, n9947, n9948, n9949, n9950, n9951,
    n9952, n9953, n9954, n9955, n9956, n9957,
    n9958, n9959, n9960, n9961, n9962, n9963,
    n9964, n9965, n9966, n9967, n9968, n9969,
    n9970, n9971, n9972, n9973, n9974, n9975,
    n9976, n9977, n9978, n9979, n9980, n9981,
    n9982, n9983, n9984, n9985, n9986, n9987,
    n9988, n9989, n9990, n9991, n9992, n9993,
    n9994, n9995, n9996, n9997, n9998, n9999,
    n10000, n10001, n10002, n10003, n10004, n10005,
    n10006, n10007, n10008, n10009, n10010, n10011,
    n10012, n10013, n10014, n10015, n10016, n10017,
    n10018, n10019, n10020, n10021, n10022, n10023,
    n10024, n10025, n10026, n10027, n10028, n10029,
    n10030, n10031, n10032, n10033, n10034, n10035,
    n10036, n10037, n10038, n10039, n10040, n10041,
    n10042, n10043, n10044, n10045, n10046, n10047,
    n10048, n10049, n10050, n10051, n10052, n10053,
    n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065,
    n10066, n10067, n10068, n10069, n10070, n10071,
    n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083,
    n10084, n10085, n10086, n10087, n10088, n10089,
    n10091, n10092, n10093, n10094, n10095, n10096,
    n10097, n10098, n10099, n10100, n10101, n10102,
    n10103, n10104, n10105, n10106, n10107, n10108,
    n10109, n10110, n10111, n10112, n10113, n10114,
    n10115, n10116, n10117, n10118, n10119, n10120,
    n10121, n10122, n10123, n10124, n10125, n10126,
    n10127, n10128, n10129, n10130, n10131, n10132,
    n10133, n10134, n10135, n10136, n10137, n10138,
    n10139, n10140, n10141, n10142, n10143, n10144,
    n10145, n10146, n10147, n10148, n10149, n10150,
    n10151, n10152, n10153, n10154, n10155, n10156,
    n10157, n10158, n10159, n10160, n10161, n10162,
    n10163, n10164, n10165, n10166, n10167, n10168,
    n10169, n10170, n10171, n10172, n10173, n10174,
    n10175, n10176, n10177, n10178, n10179, n10180,
    n10181, n10182, n10183, n10184, n10185, n10186,
    n10187, n10188, n10189, n10190, n10191, n10192,
    n10193, n10194, n10195, n10196, n10197, n10198,
    n10199, n10200, n10201, n10202, n10203, n10204,
    n10205, n10206, n10207, n10208, n10209, n10210,
    n10211, n10212, n10213, n10214, n10215, n10216,
    n10217, n10218, n10219, n10220, n10221, n10222,
    n10223, n10224, n10225, n10226, n10227, n10228,
    n10229, n10230, n10231, n10232, n10233, n10234,
    n10235, n10236, n10237, n10238, n10239, n10240,
    n10241, n10242, n10243, n10244, n10245, n10246,
    n10247, n10248, n10249, n10250, n10251, n10252,
    n10253, n10254, n10255, n10256, n10257, n10258,
    n10259, n10260, n10261, n10262, n10263, n10264,
    n10265, n10266, n10267, n10268, n10269, n10270,
    n10271, n10272, n10273, n10274, n10275, n10276,
    n10277, n10278, n10279, n10280, n10281, n10282,
    n10283, n10284, n10285, n10286, n10287, n10288,
    n10289, n10290, n10291, n10292, n10293, n10294,
    n10295, n10296, n10297, n10298, n10299, n10300,
    n10301, n10302, n10303, n10304, n10305, n10306,
    n10307, n10308, n10309, n10310, n10311, n10312,
    n10313, n10314, n10315, n10316, n10317, n10318,
    n10319, n10320, n10321, n10322, n10323, n10324,
    n10325, n10326, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10335, n10336,
    n10337, n10338, n10339, n10340, n10341, n10342,
    n10343, n10344, n10345, n10346, n10347, n10348,
    n10349, n10350, n10351, n10352, n10353, n10354,
    n10355, n10356, n10357, n10358, n10359, n10360,
    n10361, n10362, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10371, n10372,
    n10373, n10374, n10375, n10376, n10377, n10378,
    n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10387, n10388, n10389, n10390,
    n10391, n10392, n10393, n10394, n10395, n10396,
    n10397, n10398, n10399, n10400, n10401, n10402,
    n10403, n10404, n10405, n10406, n10407, n10408,
    n10409, n10410, n10411, n10412, n10413, n10414,
    n10415, n10416, n10417, n10418, n10419, n10420,
    n10421, n10422, n10423, n10424, n10425, n10426,
    n10427, n10428, n10429, n10430, n10431, n10432,
    n10433, n10434, n10435, n10436, n10437, n10438,
    n10439, n10440, n10441, n10442, n10443, n10444,
    n10445, n10446, n10447, n10448, n10449, n10450,
    n10451, n10452, n10453, n10454, n10455, n10456,
    n10457, n10458, n10459, n10460, n10461, n10462,
    n10463, n10464, n10465, n10466, n10467, n10468,
    n10469, n10470, n10471, n10472, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10480,
    n10481, n10482, n10483, n10484, n10485, n10486,
    n10487, n10488, n10489, n10490, n10491, n10492,
    n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504,
    n10505, n10506, n10507, n10508, n10509, n10510,
    n10511, n10512, n10513, n10514, n10515, n10516,
    n10518, n10519, n10520, n10521, n10522, n10523,
    n10524, n10525, n10526, n10527, n10528, n10529,
    n10530, n10531, n10532, n10533, n10534, n10535,
    n10536, n10537, n10538, n10539, n10540, n10541,
    n10542, n10543, n10544, n10545, n10546, n10547,
    n10548, n10549, n10550, n10551, n10552, n10553,
    n10554, n10555, n10556, n10557, n10558, n10559,
    n10560, n10561, n10562, n10563, n10564, n10565,
    n10566, n10567, n10568, n10569, n10570, n10571,
    n10572, n10573, n10574, n10575, n10576, n10577,
    n10578, n10579, n10580, n10581, n10582, n10583,
    n10584, n10585, n10586, n10587, n10588, n10589,
    n10590, n10591, n10592, n10593, n10594, n10595,
    n10596, n10597, n10598, n10599, n10600, n10601,
    n10602, n10603, n10604, n10605, n10606, n10607,
    n10608, n10609, n10610, n10611, n10612, n10613,
    n10614, n10615, n10616, n10617, n10618, n10619,
    n10620, n10621, n10622, n10623, n10624, n10625,
    n10626, n10627, n10628, n10629, n10630, n10631,
    n10632, n10633, n10634, n10635, n10636, n10637,
    n10638, n10639, n10640, n10641, n10642, n10643,
    n10644, n10645, n10646, n10647, n10648, n10649,
    n10650, n10651, n10652, n10653, n10654, n10655,
    n10656, n10657, n10658, n10659, n10660, n10661,
    n10662, n10663, n10664, n10665, n10666, n10667,
    n10668, n10669, n10670, n10671, n10672, n10673,
    n10674, n10675, n10676, n10677, n10678, n10679,
    n10680, n10681, n10682, n10683, n10684, n10685,
    n10686, n10687, n10688, n10689, n10690, n10691,
    n10692, n10693, n10694, n10695, n10696, n10697,
    n10698, n10699, n10700, n10701, n10702, n10703,
    n10704, n10705, n10706, n10707, n10708, n10709,
    n10710, n10711, n10712, n10713, n10714, n10715,
    n10716, n10717, n10718, n10719, n10720, n10721,
    n10722, n10723, n10724, n10725, n10726, n10727,
    n10728, n10729, n10730, n10731, n10732, n10733,
    n10734, n10735, n10736, n10737, n10738, n10739,
    n10740, n10741, n10742, n10743, n10744, n10745,
    n10746, n10747, n10748, n10749, n10750, n10751,
    n10752, n10753, n10754, n10755, n10756, n10757,
    n10758, n10759, n10760, n10761, n10762, n10763,
    n10764, n10765, n10766, n10767, n10768, n10769,
    n10770, n10771, n10772, n10773, n10774, n10775,
    n10776, n10777, n10778, n10779, n10780, n10781,
    n10782, n10783, n10784, n10785, n10786, n10787,
    n10788, n10789, n10790, n10791, n10792, n10793,
    n10794, n10795, n10796, n10797, n10798, n10799,
    n10800, n10801, n10802, n10803, n10804, n10805,
    n10806, n10807, n10808, n10809, n10810, n10811,
    n10812, n10813, n10814, n10815, n10816, n10817,
    n10818, n10819, n10820, n10821, n10822, n10823,
    n10824, n10825, n10826, n10827, n10828, n10829,
    n10830, n10831, n10832, n10833, n10834, n10835,
    n10836, n10837, n10838, n10839, n10840, n10841,
    n10842, n10843, n10844, n10845, n10846, n10847,
    n10848, n10849, n10850, n10851, n10852, n10853,
    n10854, n10855, n10856, n10857, n10858, n10859,
    n10860, n10861, n10862, n10863, n10864, n10865,
    n10866, n10867, n10868, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877,
    n10878, n10879, n10880, n10881, n10882, n10883,
    n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895,
    n10896, n10897, n10898, n10899, n10900, n10901,
    n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913,
    n10914, n10915, n10916, n10917, n10918, n10919,
    n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931,
    n10932, n10933, n10934, n10935, n10936, n10937,
    n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949,
    n10950, n10951, n10952, n10954, n10955, n10956,
    n10957, n10958, n10959, n10960, n10961, n10962,
    n10963, n10964, n10965, n10966, n10967, n10968,
    n10969, n10970, n10971, n10972, n10973, n10974,
    n10975, n10976, n10977, n10978, n10979, n10980,
    n10981, n10982, n10983, n10984, n10985, n10986,
    n10987, n10988, n10989, n10990, n10991, n10992,
    n10993, n10994, n10995, n10996, n10997, n10998,
    n10999, n11000, n11001, n11002, n11003, n11004,
    n11005, n11006, n11007, n11008, n11009, n11010,
    n11011, n11012, n11013, n11014, n11015, n11016,
    n11017, n11018, n11019, n11020, n11021, n11022,
    n11023, n11024, n11025, n11026, n11027, n11028,
    n11029, n11030, n11031, n11032, n11033, n11034,
    n11035, n11036, n11037, n11038, n11039, n11040,
    n11041, n11042, n11043, n11044, n11045, n11046,
    n11047, n11048, n11049, n11050, n11051, n11052,
    n11053, n11054, n11055, n11056, n11057, n11058,
    n11059, n11060, n11061, n11062, n11063, n11064,
    n11065, n11066, n11067, n11068, n11069, n11070,
    n11071, n11072, n11073, n11074, n11075, n11076,
    n11077, n11078, n11079, n11080, n11081, n11082,
    n11083, n11084, n11085, n11086, n11087, n11088,
    n11089, n11090, n11091, n11092, n11093, n11094,
    n11095, n11096, n11097, n11098, n11099, n11100,
    n11101, n11102, n11103, n11104, n11105, n11106,
    n11107, n11108, n11109, n11110, n11111, n11112,
    n11113, n11114, n11115, n11116, n11117, n11118,
    n11119, n11120, n11121, n11122, n11123, n11124,
    n11125, n11126, n11127, n11128, n11129, n11130,
    n11131, n11132, n11133, n11134, n11135, n11136,
    n11137, n11138, n11139, n11140, n11141, n11142,
    n11143, n11144, n11145, n11146, n11147, n11148,
    n11149, n11150, n11151, n11152, n11153, n11154,
    n11155, n11156, n11157, n11158, n11159, n11160,
    n11161, n11162, n11163, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172,
    n11173, n11174, n11175, n11176, n11177, n11178,
    n11179, n11180, n11181, n11182, n11183, n11184,
    n11185, n11186, n11187, n11188, n11189, n11190,
    n11191, n11192, n11193, n11194, n11195, n11196,
    n11197, n11198, n11199, n11200, n11201, n11202,
    n11203, n11204, n11205, n11206, n11207, n11208,
    n11209, n11210, n11211, n11212, n11213, n11214,
    n11215, n11216, n11217, n11218, n11219, n11220,
    n11221, n11222, n11223, n11224, n11225, n11226,
    n11227, n11228, n11229, n11230, n11231, n11232,
    n11233, n11234, n11235, n11236, n11237, n11238,
    n11239, n11240, n11241, n11242, n11243, n11244,
    n11245, n11246, n11247, n11248, n11249, n11250,
    n11251, n11252, n11253, n11254, n11255, n11256,
    n11257, n11258, n11259, n11260, n11261, n11262,
    n11263, n11264, n11265, n11266, n11267, n11268,
    n11269, n11270, n11271, n11272, n11273, n11274,
    n11275, n11276, n11277, n11278, n11279, n11280,
    n11281, n11282, n11283, n11284, n11285, n11286,
    n11287, n11288, n11289, n11290, n11291, n11292,
    n11293, n11294, n11295, n11296, n11297, n11298,
    n11299, n11300, n11301, n11302, n11303, n11304,
    n11305, n11306, n11307, n11308, n11309, n11310,
    n11311, n11312, n11313, n11314, n11315, n11316,
    n11317, n11318, n11319, n11320, n11321, n11322,
    n11323, n11324, n11325, n11326, n11327, n11328,
    n11329, n11330, n11331, n11332, n11333, n11334,
    n11335, n11336, n11337, n11338, n11339, n11340,
    n11341, n11342, n11343, n11344, n11345, n11346,
    n11347, n11348, n11349, n11350, n11351, n11352,
    n11353, n11354, n11355, n11356, n11357, n11358,
    n11359, n11360, n11361, n11362, n11363, n11364,
    n11365, n11366, n11367, n11368, n11369, n11370,
    n11371, n11372, n11373, n11374, n11375, n11376,
    n11377, n11378, n11379, n11380, n11381, n11382,
    n11383, n11384, n11385, n11386, n11387, n11388,
    n11389, n11390, n11391, n11392, n11393, n11394,
    n11395, n11396, n11397, n11399, n11400, n11401,
    n11402, n11403, n11404, n11405, n11406, n11407,
    n11408, n11409, n11410, n11411, n11412, n11413,
    n11414, n11415, n11416, n11417, n11418, n11419,
    n11420, n11421, n11422, n11423, n11424, n11425,
    n11426, n11427, n11428, n11429, n11430, n11431,
    n11432, n11433, n11434, n11435, n11436, n11437,
    n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449,
    n11450, n11451, n11452, n11453, n11454, n11455,
    n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473,
    n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497,
    n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515,
    n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527,
    n11528, n11529, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545,
    n11546, n11547, n11548, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575,
    n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11590, n11591, n11592, n11593,
    n11594, n11595, n11596, n11597, n11598, n11599,
    n11600, n11601, n11602, n11603, n11604, n11605,
    n11606, n11607, n11608, n11609, n11610, n11611,
    n11612, n11613, n11614, n11615, n11616, n11617,
    n11618, n11619, n11620, n11621, n11622, n11623,
    n11624, n11625, n11626, n11627, n11628, n11629,
    n11630, n11631, n11632, n11633, n11634, n11635,
    n11636, n11637, n11638, n11639, n11640, n11641,
    n11642, n11643, n11644, n11645, n11646, n11647,
    n11648, n11649, n11650, n11651, n11652, n11653,
    n11654, n11655, n11656, n11657, n11658, n11659,
    n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671,
    n11672, n11673, n11674, n11675, n11676, n11677,
    n11678, n11679, n11680, n11681, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11693, n11694, n11695,
    n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11706, n11707,
    n11708, n11709, n11710, n11711, n11712, n11713,
    n11714, n11715, n11716, n11717, n11718, n11719,
    n11720, n11721, n11722, n11723, n11724, n11725,
    n11726, n11727, n11728, n11729, n11730, n11731,
    n11732, n11733, n11734, n11735, n11736, n11737,
    n11738, n11739, n11740, n11741, n11742, n11743,
    n11744, n11745, n11746, n11747, n11748, n11749,
    n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761,
    n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779,
    n11780, n11781, n11782, n11783, n11784, n11785,
    n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797,
    n11798, n11799, n11800, n11801, n11802, n11803,
    n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815,
    n11816, n11817, n11818, n11819, n11820, n11821,
    n11822, n11823, n11824, n11825, n11826, n11827,
    n11828, n11829, n11830, n11831, n11832, n11833,
    n11834, n11835, n11836, n11837, n11838, n11839,
    n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11849, n11850, n11851,
    n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218,
    n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236,
    n12237, n12238, n12239, n12240, n12241, n12242,
    n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254,
    n12255, n12256, n12257, n12258, n12259, n12260,
    n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272,
    n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290,
    n12291, n12292, n12293, n12294, n12295, n12296,
    n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314,
    n12316, n12317, n12318, n12319, n12320, n12321,
    n12322, n12323, n12324, n12325, n12326, n12327,
    n12328, n12329, n12330, n12331, n12332, n12333,
    n12334, n12335, n12336, n12337, n12338, n12339,
    n12340, n12341, n12342, n12343, n12344, n12345,
    n12346, n12347, n12348, n12349, n12350, n12351,
    n12352, n12353, n12354, n12355, n12356, n12357,
    n12358, n12359, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369,
    n12370, n12371, n12372, n12373, n12374, n12375,
    n12376, n12377, n12378, n12379, n12380, n12381,
    n12382, n12383, n12384, n12385, n12386, n12387,
    n12388, n12389, n12390, n12391, n12392, n12393,
    n12394, n12395, n12396, n12397, n12398, n12399,
    n12400, n12401, n12402, n12403, n12404, n12405,
    n12406, n12407, n12408, n12409, n12410, n12411,
    n12412, n12413, n12414, n12415, n12416, n12417,
    n12418, n12419, n12420, n12421, n12422, n12423,
    n12424, n12425, n12426, n12427, n12428, n12429,
    n12430, n12431, n12432, n12433, n12434, n12435,
    n12436, n12437, n12438, n12439, n12440, n12441,
    n12442, n12443, n12444, n12445, n12446, n12447,
    n12448, n12449, n12450, n12451, n12452, n12453,
    n12454, n12455, n12456, n12457, n12458, n12459,
    n12460, n12461, n12462, n12463, n12464, n12465,
    n12466, n12467, n12468, n12469, n12470, n12471,
    n12472, n12473, n12474, n12475, n12476, n12477,
    n12478, n12479, n12480, n12481, n12482, n12483,
    n12484, n12485, n12486, n12487, n12488, n12489,
    n12490, n12491, n12492, n12493, n12494, n12495,
    n12496, n12497, n12498, n12499, n12500, n12501,
    n12502, n12503, n12504, n12505, n12506, n12507,
    n12508, n12509, n12510, n12511, n12512, n12513,
    n12514, n12515, n12516, n12517, n12518, n12519,
    n12520, n12521, n12522, n12523, n12524, n12525,
    n12526, n12527, n12528, n12529, n12530, n12531,
    n12532, n12533, n12534, n12535, n12536, n12537,
    n12538, n12539, n12540, n12541, n12542, n12543,
    n12544, n12545, n12546, n12547, n12548, n12549,
    n12550, n12551, n12552, n12553, n12554, n12555,
    n12556, n12557, n12558, n12559, n12560, n12561,
    n12562, n12563, n12564, n12565, n12566, n12567,
    n12568, n12569, n12570, n12571, n12572, n12573,
    n12574, n12575, n12576, n12577, n12578, n12579,
    n12580, n12581, n12582, n12583, n12584, n12585,
    n12586, n12587, n12588, n12589, n12590, n12591,
    n12592, n12593, n12594, n12595, n12596, n12597,
    n12598, n12599, n12600, n12601, n12602, n12603,
    n12604, n12605, n12606, n12607, n12608, n12609,
    n12610, n12611, n12612, n12613, n12614, n12615,
    n12616, n12617, n12618, n12619, n12620, n12621,
    n12622, n12623, n12624, n12625, n12626, n12627,
    n12628, n12629, n12630, n12631, n12632, n12633,
    n12634, n12635, n12636, n12637, n12638, n12639,
    n12640, n12641, n12642, n12643, n12644, n12645,
    n12646, n12647, n12648, n12649, n12650, n12651,
    n12652, n12653, n12654, n12655, n12656, n12657,
    n12658, n12659, n12660, n12661, n12662, n12663,
    n12664, n12665, n12666, n12667, n12668, n12669,
    n12670, n12671, n12672, n12673, n12674, n12675,
    n12676, n12677, n12678, n12679, n12680, n12681,
    n12682, n12683, n12684, n12685, n12686, n12687,
    n12688, n12689, n12690, n12691, n12692, n12693,
    n12694, n12695, n12696, n12697, n12698, n12699,
    n12700, n12701, n12702, n12703, n12704, n12705,
    n12706, n12707, n12708, n12709, n12710, n12711,
    n12712, n12713, n12714, n12715, n12716, n12717,
    n12718, n12719, n12720, n12721, n12722, n12723,
    n12724, n12725, n12726, n12727, n12728, n12729,
    n12730, n12731, n12732, n12733, n12734, n12735,
    n12736, n12737, n12738, n12739, n12740, n12741,
    n12742, n12743, n12744, n12745, n12746, n12747,
    n12748, n12749, n12750, n12751, n12752, n12753,
    n12754, n12755, n12756, n12757, n12758, n12759,
    n12760, n12761, n12762, n12763, n12764, n12765,
    n12766, n12767, n12768, n12769, n12770, n12771,
    n12772, n12773, n12774, n12775, n12776, n12777,
    n12778, n12779, n12780, n12781, n12782, n12783,
    n12784, n12785, n12786, n12788, n12789, n12790,
    n12791, n12792, n12793, n12794, n12795, n12796,
    n12797, n12798, n12799, n12800, n12801, n12802,
    n12803, n12804, n12805, n12806, n12807, n12808,
    n12809, n12810, n12811, n12812, n12813, n12814,
    n12815, n12816, n12817, n12818, n12819, n12820,
    n12821, n12822, n12823, n12824, n12825, n12826,
    n12827, n12828, n12829, n12830, n12831, n12832,
    n12833, n12834, n12835, n12836, n12837, n12838,
    n12839, n12840, n12841, n12842, n12843, n12844,
    n12845, n12846, n12847, n12848, n12849, n12850,
    n12851, n12852, n12853, n12854, n12855, n12856,
    n12857, n12858, n12859, n12860, n12861, n12862,
    n12863, n12864, n12865, n12866, n12867, n12868,
    n12869, n12870, n12871, n12872, n12873, n12874,
    n12875, n12876, n12877, n12878, n12879, n12880,
    n12881, n12882, n12883, n12884, n12885, n12886,
    n12887, n12888, n12889, n12890, n12891, n12892,
    n12893, n12894, n12895, n12896, n12897, n12898,
    n12899, n12900, n12901, n12902, n12903, n12904,
    n12905, n12906, n12907, n12908, n12909, n12910,
    n12911, n12912, n12913, n12914, n12915, n12916,
    n12917, n12918, n12919, n12920, n12921, n12922,
    n12923, n12924, n12925, n12926, n12927, n12928,
    n12929, n12930, n12931, n12932, n12933, n12934,
    n12935, n12936, n12937, n12938, n12939, n12940,
    n12941, n12942, n12943, n12944, n12945, n12946,
    n12947, n12948, n12949, n12950, n12951, n12952,
    n12953, n12954, n12955, n12956, n12957, n12958,
    n12959, n12960, n12961, n12962, n12963, n12964,
    n12965, n12966, n12967, n12968, n12969, n12970,
    n12971, n12972, n12973, n12974, n12975, n12976,
    n12977, n12978, n12979, n12980, n12981, n12982,
    n12983, n12984, n12985, n12986, n12987, n12988,
    n12989, n12990, n12991, n12992, n12993, n12994,
    n12995, n12996, n12997, n12998, n12999, n13000,
    n13001, n13002, n13003, n13004, n13005, n13006,
    n13007, n13008, n13009, n13010, n13011, n13012,
    n13013, n13014, n13015, n13016, n13017, n13018,
    n13019, n13020, n13021, n13022, n13023, n13024,
    n13025, n13026, n13027, n13028, n13029, n13030,
    n13031, n13032, n13033, n13034, n13035, n13036,
    n13037, n13038, n13039, n13040, n13041, n13042,
    n13043, n13044, n13045, n13046, n13047, n13048,
    n13049, n13050, n13051, n13052, n13053, n13054,
    n13055, n13056, n13057, n13058, n13059, n13060,
    n13061, n13062, n13063, n13064, n13065, n13066,
    n13067, n13068, n13069, n13070, n13071, n13072,
    n13073, n13074, n13075, n13076, n13077, n13078,
    n13079, n13080, n13081, n13082, n13083, n13084,
    n13085, n13086, n13087, n13088, n13089, n13090,
    n13091, n13092, n13093, n13094, n13095, n13096,
    n13097, n13098, n13099, n13100, n13101, n13102,
    n13103, n13104, n13105, n13106, n13107, n13108,
    n13109, n13110, n13111, n13112, n13113, n13114,
    n13115, n13116, n13117, n13118, n13119, n13120,
    n13121, n13122, n13123, n13124, n13125, n13126,
    n13127, n13128, n13129, n13130, n13131, n13132,
    n13133, n13134, n13135, n13136, n13137, n13138,
    n13139, n13140, n13141, n13142, n13143, n13144,
    n13145, n13146, n13147, n13148, n13149, n13150,
    n13151, n13152, n13153, n13154, n13155, n13156,
    n13157, n13158, n13159, n13160, n13161, n13162,
    n13163, n13164, n13165, n13166, n13167, n13168,
    n13169, n13170, n13171, n13172, n13173, n13174,
    n13175, n13176, n13177, n13178, n13179, n13180,
    n13181, n13182, n13183, n13184, n13185, n13186,
    n13187, n13188, n13189, n13190, n13191, n13192,
    n13193, n13194, n13195, n13196, n13197, n13198,
    n13199, n13200, n13201, n13202, n13203, n13204,
    n13205, n13206, n13207, n13208, n13209, n13210,
    n13211, n13212, n13213, n13214, n13215, n13216,
    n13217, n13218, n13219, n13220, n13221, n13222,
    n13223, n13224, n13225, n13226, n13227, n13228,
    n13229, n13230, n13231, n13232, n13233, n13234,
    n13235, n13236, n13237, n13238, n13239, n13240,
    n13241, n13242, n13243, n13244, n13245, n13246,
    n13247, n13248, n13249, n13250, n13251, n13252,
    n13253, n13254, n13255, n13256, n13257, n13258,
    n13259, n13260, n13261, n13262, n13263, n13264,
    n13265, n13266, n13267, n13269, n13270, n13271,
    n13272, n13273, n13274, n13275, n13276, n13277,
    n13278, n13279, n13280, n13281, n13282, n13283,
    n13284, n13285, n13286, n13287, n13288, n13289,
    n13290, n13291, n13292, n13293, n13294, n13295,
    n13296, n13297, n13298, n13299, n13300, n13301,
    n13302, n13303, n13304, n13305, n13306, n13307,
    n13308, n13309, n13310, n13311, n13312, n13313,
    n13314, n13315, n13316, n13317, n13318, n13319,
    n13320, n13321, n13322, n13323, n13324, n13325,
    n13326, n13327, n13328, n13329, n13330, n13331,
    n13332, n13333, n13334, n13335, n13336, n13337,
    n13338, n13339, n13340, n13341, n13342, n13343,
    n13344, n13345, n13346, n13347, n13348, n13349,
    n13350, n13351, n13352, n13353, n13354, n13355,
    n13356, n13357, n13358, n13359, n13360, n13361,
    n13362, n13363, n13364, n13365, n13366, n13367,
    n13368, n13369, n13370, n13371, n13372, n13373,
    n13374, n13375, n13376, n13377, n13378, n13379,
    n13380, n13381, n13382, n13383, n13384, n13385,
    n13386, n13387, n13388, n13389, n13390, n13391,
    n13392, n13393, n13394, n13395, n13396, n13397,
    n13398, n13399, n13400, n13401, n13402, n13403,
    n13404, n13405, n13406, n13407, n13408, n13409,
    n13410, n13411, n13412, n13413, n13414, n13415,
    n13416, n13417, n13418, n13419, n13420, n13421,
    n13422, n13423, n13424, n13425, n13426, n13427,
    n13428, n13429, n13430, n13431, n13432, n13433,
    n13434, n13435, n13436, n13437, n13438, n13439,
    n13440, n13441, n13442, n13443, n13444, n13445,
    n13446, n13447, n13448, n13449, n13450, n13451,
    n13452, n13453, n13454, n13455, n13456, n13457,
    n13458, n13459, n13460, n13461, n13462, n13463,
    n13464, n13465, n13466, n13467, n13468, n13469,
    n13470, n13471, n13472, n13473, n13474, n13475,
    n13476, n13477, n13478, n13479, n13480, n13481,
    n13482, n13483, n13484, n13485, n13486, n13487,
    n13488, n13489, n13490, n13491, n13492, n13493,
    n13494, n13495, n13496, n13497, n13498, n13499,
    n13500, n13501, n13502, n13503, n13504, n13505,
    n13506, n13507, n13508, n13509, n13510, n13511,
    n13512, n13513, n13514, n13515, n13516, n13517,
    n13518, n13519, n13520, n13521, n13522, n13523,
    n13524, n13525, n13526, n13527, n13528, n13529,
    n13530, n13531, n13532, n13533, n13534, n13535,
    n13536, n13537, n13538, n13539, n13540, n13541,
    n13542, n13543, n13544, n13545, n13546, n13547,
    n13548, n13549, n13550, n13551, n13552, n13553,
    n13554, n13555, n13556, n13557, n13558, n13559,
    n13560, n13561, n13562, n13563, n13564, n13565,
    n13566, n13567, n13568, n13569, n13570, n13571,
    n13572, n13573, n13574, n13575, n13576, n13577,
    n13578, n13579, n13580, n13581, n13582, n13583,
    n13584, n13585, n13586, n13587, n13588, n13589,
    n13590, n13591, n13592, n13593, n13594, n13595,
    n13596, n13597, n13598, n13599, n13600, n13601,
    n13602, n13603, n13604, n13605, n13606, n13607,
    n13608, n13609, n13610, n13611, n13612, n13613,
    n13614, n13615, n13616, n13617, n13618, n13619,
    n13620, n13621, n13622, n13623, n13624, n13625,
    n13626, n13627, n13628, n13629, n13630, n13631,
    n13632, n13633, n13634, n13635, n13636, n13637,
    n13638, n13639, n13640, n13641, n13642, n13643,
    n13644, n13645, n13646, n13647, n13648, n13649,
    n13650, n13651, n13652, n13653, n13654, n13655,
    n13656, n13657, n13658, n13659, n13660, n13661,
    n13662, n13663, n13664, n13665, n13666, n13667,
    n13668, n13669, n13670, n13671, n13672, n13673,
    n13674, n13675, n13676, n13677, n13678, n13679,
    n13680, n13681, n13682, n13683, n13684, n13685,
    n13686, n13687, n13688, n13689, n13690, n13691,
    n13692, n13693, n13694, n13695, n13696, n13697,
    n13698, n13699, n13700, n13701, n13702, n13703,
    n13704, n13705, n13706, n13707, n13708, n13709,
    n13710, n13711, n13712, n13713, n13714, n13715,
    n13716, n13717, n13718, n13719, n13720, n13721,
    n13722, n13723, n13724, n13725, n13726, n13727,
    n13728, n13729, n13730, n13731, n13732, n13733,
    n13734, n13735, n13736, n13737, n13738, n13739,
    n13740, n13741, n13742, n13743, n13744, n13745,
    n13746, n13747, n13748, n13749, n13750, n13751,
    n13752, n13753, n13754, n13755, n13756, n13757,
    n13759, n13760, n13761, n13762, n13763, n13764,
    n13765, n13766, n13767, n13768, n13769, n13770,
    n13771, n13772, n13773, n13774, n13775, n13776,
    n13777, n13778, n13779, n13780, n13781, n13782,
    n13783, n13784, n13785, n13786, n13787, n13788,
    n13789, n13790, n13791, n13792, n13793, n13794,
    n13795, n13796, n13797, n13798, n13799, n13800,
    n13801, n13802, n13803, n13804, n13805, n13806,
    n13807, n13808, n13809, n13810, n13811, n13812,
    n13813, n13814, n13815, n13816, n13817, n13818,
    n13819, n13820, n13821, n13822, n13823, n13824,
    n13825, n13826, n13827, n13828, n13829, n13830,
    n13831, n13832, n13833, n13834, n13835, n13836,
    n13837, n13838, n13839, n13840, n13841, n13842,
    n13843, n13844, n13845, n13846, n13847, n13848,
    n13849, n13850, n13851, n13852, n13853, n13854,
    n13855, n13856, n13857, n13858, n13859, n13860,
    n13861, n13862, n13863, n13864, n13865, n13866,
    n13867, n13868, n13869, n13870, n13871, n13872,
    n13873, n13874, n13875, n13876, n13877, n13878,
    n13879, n13880, n13881, n13882, n13883, n13884,
    n13885, n13886, n13887, n13888, n13889, n13890,
    n13891, n13892, n13893, n13894, n13895, n13896,
    n13897, n13898, n13899, n13900, n13901, n13902,
    n13903, n13904, n13905, n13906, n13907, n13908,
    n13909, n13910, n13911, n13912, n13913, n13914,
    n13915, n13916, n13917, n13918, n13919, n13920,
    n13921, n13922, n13923, n13924, n13925, n13926,
    n13927, n13928, n13929, n13930, n13931, n13932,
    n13933, n13934, n13935, n13936, n13937, n13938,
    n13939, n13940, n13941, n13942, n13943, n13944,
    n13945, n13946, n13947, n13948, n13949, n13950,
    n13951, n13952, n13953, n13954, n13955, n13956,
    n13957, n13958, n13959, n13960, n13961, n13962,
    n13963, n13964, n13965, n13966, n13967, n13968,
    n13969, n13970, n13971, n13972, n13973, n13974,
    n13975, n13976, n13977, n13978, n13979, n13980,
    n13981, n13982, n13983, n13984, n13985, n13986,
    n13987, n13988, n13989, n13990, n13991, n13992,
    n13993, n13994, n13995, n13996, n13997, n13998,
    n13999, n14000, n14001, n14002, n14003, n14004,
    n14005, n14006, n14007, n14008, n14009, n14010,
    n14011, n14012, n14013, n14014, n14015, n14016,
    n14017, n14018, n14019, n14020, n14021, n14022,
    n14023, n14024, n14025, n14026, n14027, n14028,
    n14029, n14030, n14031, n14032, n14033, n14034,
    n14035, n14036, n14037, n14038, n14039, n14040,
    n14041, n14042, n14043, n14044, n14045, n14046,
    n14047, n14048, n14049, n14050, n14051, n14052,
    n14053, n14054, n14055, n14056, n14057, n14058,
    n14059, n14060, n14061, n14062, n14063, n14064,
    n14065, n14066, n14067, n14068, n14069, n14070,
    n14071, n14072, n14073, n14074, n14075, n14076,
    n14077, n14078, n14079, n14080, n14081, n14082,
    n14083, n14084, n14085, n14086, n14087, n14088,
    n14089, n14090, n14091, n14092, n14093, n14094,
    n14095, n14096, n14097, n14098, n14099, n14100,
    n14101, n14102, n14103, n14104, n14105, n14106,
    n14107, n14108, n14109, n14110, n14111, n14112,
    n14113, n14114, n14115, n14116, n14117, n14118,
    n14119, n14120, n14121, n14122, n14123, n14124,
    n14125, n14126, n14127, n14128, n14129, n14130,
    n14131, n14132, n14133, n14134, n14135, n14136,
    n14137, n14138, n14139, n14140, n14141, n14142,
    n14143, n14144, n14145, n14146, n14147, n14148,
    n14149, n14150, n14151, n14152, n14153, n14154,
    n14155, n14156, n14157, n14158, n14159, n14160,
    n14161, n14162, n14163, n14164, n14165, n14166,
    n14167, n14168, n14169, n14170, n14171, n14172,
    n14173, n14174, n14175, n14176, n14177, n14178,
    n14179, n14180, n14181, n14182, n14183, n14184,
    n14185, n14186, n14187, n14188, n14189, n14190,
    n14191, n14192, n14193, n14194, n14195, n14196,
    n14197, n14198, n14199, n14200, n14201, n14202,
    n14203, n14204, n14205, n14206, n14207, n14208,
    n14209, n14210, n14211, n14212, n14213, n14214,
    n14215, n14216, n14217, n14218, n14219, n14220,
    n14221, n14222, n14223, n14224, n14225, n14226,
    n14227, n14228, n14229, n14230, n14231, n14232,
    n14233, n14234, n14235, n14236, n14237, n14238,
    n14239, n14240, n14241, n14242, n14243, n14244,
    n14245, n14246, n14247, n14248, n14249, n14250,
    n14251, n14252, n14253, n14254, n14255, n14256,
    n14258, n14259, n14260, n14261, n14262, n14263,
    n14264, n14265, n14266, n14267, n14268, n14269,
    n14270, n14271, n14272, n14273, n14274, n14275,
    n14276, n14277, n14278, n14279, n14280, n14281,
    n14282, n14283, n14284, n14285, n14286, n14287,
    n14288, n14289, n14290, n14291, n14292, n14293,
    n14294, n14295, n14296, n14297, n14298, n14299,
    n14300, n14301, n14302, n14303, n14304, n14305,
    n14306, n14307, n14308, n14309, n14310, n14311,
    n14312, n14313, n14314, n14315, n14316, n14317,
    n14318, n14319, n14320, n14321, n14322, n14323,
    n14324, n14325, n14326, n14327, n14328, n14329,
    n14330, n14331, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14340, n14341,
    n14342, n14343, n14344, n14345, n14346, n14347,
    n14348, n14349, n14350, n14351, n14352, n14353,
    n14354, n14355, n14356, n14357, n14358, n14359,
    n14360, n14361, n14362, n14363, n14364, n14365,
    n14366, n14367, n14368, n14369, n14370, n14371,
    n14372, n14373, n14374, n14375, n14376, n14377,
    n14378, n14379, n14380, n14381, n14382, n14383,
    n14384, n14385, n14386, n14387, n14388, n14389,
    n14390, n14391, n14392, n14393, n14394, n14395,
    n14396, n14397, n14398, n14399, n14400, n14401,
    n14402, n14403, n14404, n14405, n14406, n14407,
    n14408, n14409, n14410, n14411, n14412, n14413,
    n14414, n14415, n14416, n14417, n14418, n14419,
    n14420, n14421, n14422, n14423, n14424, n14425,
    n14426, n14427, n14428, n14429, n14430, n14431,
    n14432, n14433, n14434, n14435, n14436, n14437,
    n14438, n14439, n14440, n14441, n14442, n14443,
    n14444, n14445, n14446, n14447, n14448, n14449,
    n14450, n14451, n14452, n14453, n14454, n14455,
    n14456, n14457, n14458, n14459, n14460, n14461,
    n14462, n14463, n14464, n14465, n14466, n14467,
    n14468, n14469, n14470, n14471, n14472, n14473,
    n14474, n14475, n14476, n14477, n14478, n14479,
    n14480, n14481, n14482, n14483, n14484, n14485,
    n14486, n14487, n14488, n14489, n14490, n14491,
    n14492, n14493, n14494, n14495, n14496, n14497,
    n14498, n14499, n14500, n14501, n14502, n14503,
    n14504, n14505, n14506, n14507, n14508, n14509,
    n14510, n14511, n14512, n14513, n14514, n14515,
    n14516, n14517, n14518, n14519, n14520, n14521,
    n14522, n14523, n14524, n14525, n14526, n14527,
    n14528, n14529, n14530, n14531, n14532, n14533,
    n14534, n14535, n14536, n14537, n14538, n14539,
    n14540, n14541, n14542, n14543, n14544, n14545,
    n14546, n14547, n14548, n14549, n14550, n14551,
    n14552, n14553, n14554, n14555, n14556, n14557,
    n14558, n14559, n14560, n14561, n14562, n14563,
    n14564, n14565, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14573, n14574, n14575,
    n14576, n14577, n14578, n14579, n14580, n14581,
    n14582, n14583, n14584, n14585, n14586, n14587,
    n14588, n14589, n14590, n14591, n14592, n14593,
    n14594, n14595, n14596, n14597, n14598, n14599,
    n14600, n14601, n14602, n14603, n14604, n14605,
    n14606, n14607, n14608, n14609, n14610, n14611,
    n14612, n14613, n14614, n14615, n14616, n14617,
    n14618, n14619, n14620, n14621, n14622, n14623,
    n14624, n14625, n14626, n14627, n14628, n14629,
    n14630, n14631, n14632, n14633, n14634, n14635,
    n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647,
    n14648, n14649, n14650, n14651, n14652, n14653,
    n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665,
    n14666, n14667, n14668, n14669, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683,
    n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701,
    n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719,
    n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731,
    n14732, n14733, n14734, n14735, n14736, n14737,
    n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749,
    n14750, n14751, n14752, n14753, n14754, n14755,
    n14756, n14757, n14758, n14759, n14760, n14761,
    n14762, n14763, n14764, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816,
    n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834,
    n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846,
    n14847, n14848, n14849, n14850, n14851, n14852,
    n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864,
    n14865, n14866, n14867, n14868, n14869, n14870,
    n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882,
    n14883, n14884, n14885, n14886, n14887, n14888,
    n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906,
    n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924,
    n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942,
    n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978,
    n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996,
    n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014,
    n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032,
    n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050,
    n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068,
    n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086,
    n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122,
    n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194,
    n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230,
    n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248,
    n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15281, n15283, n15284, n15285,
    n15286, n15287, n15288, n15289, n15290, n15291,
    n15292, n15293, n15294, n15295, n15296, n15297,
    n15298, n15299, n15300, n15301, n15302, n15303,
    n15304, n15305, n15306, n15307, n15308, n15309,
    n15310, n15311, n15312, n15313, n15314, n15315,
    n15316, n15317, n15318, n15319, n15320, n15321,
    n15322, n15323, n15324, n15325, n15326, n15327,
    n15328, n15329, n15330, n15331, n15332, n15333,
    n15334, n15335, n15336, n15337, n15338, n15339,
    n15340, n15341, n15342, n15343, n15344, n15345,
    n15346, n15347, n15348, n15349, n15350, n15351,
    n15352, n15353, n15354, n15355, n15356, n15357,
    n15358, n15359, n15360, n15361, n15362, n15363,
    n15364, n15365, n15366, n15367, n15368, n15369,
    n15370, n15371, n15372, n15373, n15374, n15375,
    n15376, n15377, n15378, n15379, n15380, n15381,
    n15382, n15383, n15384, n15385, n15386, n15387,
    n15388, n15389, n15390, n15391, n15392, n15393,
    n15394, n15395, n15396, n15397, n15398, n15399,
    n15400, n15401, n15402, n15403, n15404, n15405,
    n15406, n15407, n15408, n15409, n15410, n15411,
    n15412, n15413, n15414, n15415, n15416, n15417,
    n15418, n15419, n15420, n15421, n15422, n15423,
    n15424, n15425, n15426, n15427, n15428, n15429,
    n15430, n15431, n15432, n15433, n15434, n15435,
    n15436, n15437, n15438, n15439, n15440, n15441,
    n15442, n15443, n15444, n15445, n15446, n15447,
    n15448, n15449, n15450, n15451, n15452, n15453,
    n15454, n15455, n15456, n15457, n15458, n15459,
    n15460, n15461, n15462, n15463, n15464, n15465,
    n15466, n15467, n15468, n15469, n15470, n15471,
    n15472, n15473, n15474, n15475, n15476, n15477,
    n15478, n15479, n15480, n15481, n15482, n15483,
    n15484, n15485, n15486, n15487, n15488, n15489,
    n15490, n15491, n15492, n15493, n15494, n15495,
    n15496, n15497, n15498, n15499, n15500, n15501,
    n15502, n15503, n15504, n15505, n15506, n15507,
    n15508, n15509, n15510, n15511, n15512, n15513,
    n15514, n15515, n15516, n15517, n15518, n15519,
    n15520, n15521, n15522, n15523, n15524, n15525,
    n15526, n15527, n15528, n15529, n15530, n15531,
    n15532, n15533, n15534, n15535, n15536, n15537,
    n15538, n15539, n15540, n15541, n15542, n15543,
    n15544, n15545, n15546, n15547, n15548, n15549,
    n15550, n15551, n15552, n15553, n15554, n15555,
    n15556, n15557, n15558, n15559, n15560, n15561,
    n15562, n15563, n15564, n15565, n15566, n15567,
    n15568, n15569, n15570, n15571, n15572, n15573,
    n15574, n15575, n15576, n15577, n15578, n15579,
    n15580, n15581, n15582, n15583, n15584, n15585,
    n15586, n15587, n15588, n15589, n15590, n15591,
    n15592, n15593, n15594, n15595, n15596, n15597,
    n15598, n15599, n15600, n15601, n15602, n15603,
    n15604, n15605, n15606, n15607, n15608, n15609,
    n15610, n15611, n15612, n15613, n15614, n15615,
    n15616, n15617, n15618, n15619, n15620, n15621,
    n15622, n15623, n15624, n15625, n15626, n15627,
    n15628, n15629, n15630, n15631, n15632, n15633,
    n15634, n15635, n15636, n15637, n15638, n15639,
    n15640, n15641, n15642, n15643, n15644, n15645,
    n15646, n15647, n15648, n15649, n15650, n15651,
    n15652, n15653, n15654, n15655, n15656, n15657,
    n15658, n15659, n15660, n15661, n15662, n15663,
    n15664, n15665, n15666, n15667, n15668, n15669,
    n15670, n15671, n15672, n15673, n15674, n15675,
    n15676, n15677, n15678, n15679, n15680, n15681,
    n15682, n15683, n15684, n15685, n15686, n15687,
    n15688, n15689, n15690, n15691, n15692, n15693,
    n15694, n15695, n15696, n15697, n15698, n15699,
    n15700, n15701, n15702, n15703, n15704, n15705,
    n15706, n15707, n15708, n15709, n15710, n15711,
    n15712, n15713, n15714, n15715, n15716, n15717,
    n15718, n15719, n15720, n15721, n15722, n15723,
    n15724, n15725, n15726, n15727, n15728, n15729,
    n15730, n15731, n15732, n15733, n15734, n15735,
    n15736, n15737, n15738, n15739, n15740, n15741,
    n15742, n15743, n15744, n15745, n15746, n15747,
    n15748, n15749, n15750, n15751, n15752, n15753,
    n15754, n15755, n15756, n15757, n15758, n15759,
    n15760, n15761, n15762, n15763, n15764, n15765,
    n15766, n15767, n15768, n15769, n15770, n15771,
    n15772, n15773, n15774, n15775, n15776, n15777,
    n15778, n15779, n15780, n15781, n15782, n15783,
    n15784, n15785, n15786, n15787, n15788, n15789,
    n15790, n15791, n15792, n15793, n15794, n15795,
    n15796, n15797, n15798, n15799, n15800, n15801,
    n15802, n15803, n15804, n15805, n15807, n15808,
    n15809, n15810, n15811, n15812, n15813, n15814,
    n15815, n15816, n15817, n15818, n15819, n15820,
    n15821, n15822, n15823, n15824, n15825, n15826,
    n15827, n15828, n15829, n15830, n15831, n15832,
    n15833, n15834, n15835, n15836, n15837, n15838,
    n15839, n15840, n15841, n15842, n15843, n15844,
    n15845, n15846, n15847, n15848, n15849, n15850,
    n15851, n15852, n15853, n15854, n15855, n15856,
    n15857, n15858, n15859, n15860, n15861, n15862,
    n15863, n15864, n15865, n15866, n15867, n15868,
    n15869, n15870, n15871, n15872, n15873, n15874,
    n15875, n15876, n15877, n15878, n15879, n15880,
    n15881, n15882, n15883, n15884, n15885, n15886,
    n15887, n15888, n15889, n15890, n15891, n15892,
    n15893, n15894, n15895, n15896, n15897, n15898,
    n15899, n15900, n15901, n15902, n15903, n15904,
    n15905, n15906, n15907, n15908, n15909, n15910,
    n15911, n15912, n15913, n15914, n15915, n15916,
    n15917, n15918, n15919, n15920, n15921, n15922,
    n15923, n15924, n15925, n15926, n15927, n15928,
    n15929, n15930, n15931, n15932, n15933, n15934,
    n15935, n15936, n15937, n15938, n15939, n15940,
    n15941, n15942, n15943, n15944, n15945, n15946,
    n15947, n15948, n15949, n15950, n15951, n15952,
    n15953, n15954, n15955, n15956, n15957, n15958,
    n15959, n15960, n15961, n15962, n15963, n15964,
    n15965, n15966, n15967, n15968, n15969, n15970,
    n15971, n15972, n15973, n15974, n15975, n15976,
    n15977, n15978, n15979, n15980, n15981, n15982,
    n15983, n15984, n15985, n15986, n15987, n15988,
    n15989, n15990, n15991, n15992, n15993, n15994,
    n15995, n15996, n15997, n15998, n15999, n16000,
    n16001, n16002, n16003, n16004, n16005, n16006,
    n16007, n16008, n16009, n16010, n16011, n16012,
    n16013, n16014, n16015, n16016, n16017, n16018,
    n16019, n16020, n16021, n16022, n16023, n16024,
    n16025, n16026, n16027, n16028, n16029, n16030,
    n16031, n16032, n16033, n16034, n16035, n16036,
    n16037, n16038, n16039, n16040, n16041, n16042,
    n16043, n16044, n16045, n16046, n16047, n16048,
    n16049, n16050, n16051, n16052, n16053, n16054,
    n16055, n16056, n16057, n16058, n16059, n16060,
    n16061, n16062, n16063, n16064, n16065, n16066,
    n16067, n16068, n16069, n16070, n16071, n16072,
    n16073, n16074, n16075, n16076, n16077, n16078,
    n16079, n16080, n16081, n16082, n16083, n16084,
    n16085, n16086, n16087, n16088, n16089, n16090,
    n16091, n16092, n16093, n16094, n16095, n16096,
    n16097, n16098, n16099, n16100, n16101, n16102,
    n16103, n16104, n16105, n16106, n16107, n16108,
    n16109, n16110, n16111, n16112, n16113, n16114,
    n16115, n16116, n16117, n16118, n16119, n16120,
    n16121, n16122, n16123, n16124, n16125, n16126,
    n16127, n16128, n16129, n16130, n16131, n16132,
    n16133, n16134, n16135, n16136, n16137, n16138,
    n16139, n16140, n16141, n16142, n16143, n16144,
    n16145, n16146, n16147, n16148, n16149, n16150,
    n16151, n16152, n16153, n16154, n16155, n16156,
    n16157, n16158, n16159, n16160, n16161, n16162,
    n16163, n16164, n16165, n16166, n16167, n16168,
    n16169, n16170, n16171, n16172, n16173, n16174,
    n16175, n16176, n16177, n16178, n16179, n16180,
    n16181, n16182, n16183, n16184, n16185, n16186,
    n16187, n16188, n16189, n16190, n16191, n16192,
    n16193, n16194, n16195, n16196, n16197, n16198,
    n16199, n16200, n16201, n16202, n16203, n16204,
    n16205, n16206, n16207, n16208, n16209, n16210,
    n16211, n16212, n16213, n16214, n16215, n16216,
    n16217, n16218, n16219, n16220, n16221, n16222,
    n16223, n16224, n16225, n16226, n16227, n16228,
    n16229, n16230, n16231, n16232, n16233, n16234,
    n16235, n16236, n16237, n16238, n16239, n16240,
    n16241, n16242, n16243, n16244, n16245, n16246,
    n16247, n16248, n16249, n16250, n16251, n16252,
    n16253, n16254, n16255, n16256, n16257, n16258,
    n16259, n16260, n16261, n16262, n16263, n16264,
    n16265, n16266, n16267, n16268, n16269, n16270,
    n16271, n16272, n16273, n16274, n16275, n16276,
    n16277, n16278, n16279, n16280, n16281, n16282,
    n16283, n16284, n16285, n16286, n16287, n16288,
    n16289, n16290, n16291, n16292, n16293, n16294,
    n16295, n16296, n16297, n16298, n16299, n16300,
    n16301, n16302, n16303, n16304, n16305, n16306,
    n16307, n16308, n16309, n16310, n16311, n16312,
    n16313, n16314, n16315, n16316, n16317, n16318,
    n16319, n16320, n16321, n16322, n16323, n16324,
    n16325, n16326, n16327, n16328, n16329, n16330,
    n16331, n16332, n16333, n16334, n16335, n16336,
    n16337, n16338, n16340, n16341, n16342, n16343,
    n16344, n16345, n16346, n16347, n16348, n16349,
    n16350, n16351, n16352, n16353, n16354, n16355,
    n16356, n16357, n16358, n16359, n16360, n16361,
    n16362, n16363, n16364, n16365, n16366, n16367,
    n16368, n16369, n16370, n16371, n16372, n16373,
    n16374, n16375, n16376, n16377, n16378, n16379,
    n16380, n16381, n16382, n16383, n16384, n16385,
    n16386, n16387, n16388, n16389, n16390, n16391,
    n16392, n16393, n16394, n16395, n16396, n16397,
    n16398, n16399, n16400, n16401, n16402, n16403,
    n16404, n16405, n16406, n16407, n16408, n16409,
    n16410, n16411, n16412, n16413, n16414, n16415,
    n16416, n16417, n16418, n16419, n16420, n16421,
    n16422, n16423, n16424, n16425, n16426, n16427,
    n16428, n16429, n16430, n16431, n16432, n16433,
    n16434, n16435, n16436, n16437, n16438, n16439,
    n16440, n16441, n16442, n16443, n16444, n16445,
    n16446, n16447, n16448, n16449, n16450, n16451,
    n16452, n16453, n16454, n16455, n16456, n16457,
    n16458, n16459, n16460, n16461, n16462, n16463,
    n16464, n16465, n16466, n16467, n16468, n16469,
    n16470, n16471, n16472, n16473, n16474, n16475,
    n16476, n16477, n16478, n16479, n16480, n16481,
    n16482, n16483, n16484, n16485, n16486, n16487,
    n16488, n16489, n16490, n16491, n16492, n16493,
    n16494, n16495, n16496, n16497, n16498, n16499,
    n16500, n16501, n16502, n16503, n16504, n16505,
    n16506, n16507, n16508, n16509, n16510, n16511,
    n16512, n16513, n16514, n16515, n16516, n16517,
    n16518, n16519, n16520, n16521, n16522, n16523,
    n16524, n16525, n16526, n16527, n16528, n16529,
    n16530, n16531, n16532, n16533, n16534, n16535,
    n16536, n16537, n16538, n16539, n16540, n16541,
    n16542, n16543, n16544, n16545, n16546, n16547,
    n16548, n16549, n16550, n16551, n16552, n16553,
    n16554, n16555, n16556, n16557, n16558, n16559,
    n16560, n16561, n16562, n16563, n16564, n16565,
    n16566, n16567, n16568, n16569, n16570, n16571,
    n16572, n16573, n16574, n16575, n16576, n16577,
    n16578, n16579, n16580, n16581, n16582, n16583,
    n16584, n16585, n16586, n16587, n16588, n16589,
    n16590, n16591, n16592, n16593, n16594, n16595,
    n16596, n16597, n16598, n16599, n16600, n16601,
    n16602, n16603, n16604, n16605, n16606, n16607,
    n16608, n16609, n16610, n16611, n16612, n16613,
    n16614, n16615, n16616, n16617, n16618, n16619,
    n16620, n16621, n16622, n16623, n16624, n16625,
    n16626, n16627, n16628, n16629, n16630, n16631,
    n16632, n16633, n16634, n16635, n16636, n16637,
    n16638, n16639, n16640, n16641, n16642, n16643,
    n16644, n16645, n16646, n16647, n16648, n16649,
    n16650, n16651, n16652, n16653, n16654, n16655,
    n16656, n16657, n16658, n16659, n16660, n16661,
    n16662, n16663, n16664, n16665, n16666, n16667,
    n16668, n16669, n16670, n16671, n16672, n16673,
    n16674, n16675, n16676, n16677, n16678, n16679,
    n16680, n16681, n16682, n16683, n16684, n16685,
    n16686, n16687, n16688, n16689, n16690, n16691,
    n16692, n16693, n16694, n16695, n16696, n16697,
    n16698, n16699, n16700, n16701, n16702, n16703,
    n16704, n16705, n16706, n16707, n16708, n16709,
    n16710, n16711, n16712, n16713, n16714, n16715,
    n16716, n16717, n16718, n16719, n16720, n16721,
    n16722, n16723, n16724, n16725, n16726, n16727,
    n16728, n16729, n16730, n16731, n16732, n16733,
    n16734, n16735, n16736, n16737, n16738, n16739,
    n16740, n16741, n16742, n16743, n16744, n16745,
    n16746, n16747, n16748, n16749, n16750, n16751,
    n16752, n16753, n16754, n16755, n16756, n16757,
    n16758, n16759, n16760, n16761, n16762, n16763,
    n16764, n16765, n16766, n16767, n16768, n16769,
    n16770, n16771, n16772, n16773, n16774, n16775,
    n16776, n16777, n16778, n16779, n16780, n16781,
    n16782, n16783, n16784, n16785, n16786, n16787,
    n16788, n16789, n16790, n16791, n16792, n16793,
    n16794, n16795, n16796, n16797, n16798, n16799,
    n16800, n16801, n16802, n16803, n16804, n16805,
    n16806, n16807, n16808, n16809, n16810, n16811,
    n16812, n16813, n16814, n16815, n16816, n16817,
    n16818, n16819, n16820, n16821, n16822, n16823,
    n16824, n16825, n16826, n16827, n16828, n16829,
    n16830, n16831, n16832, n16833, n16834, n16835,
    n16836, n16837, n16838, n16839, n16840, n16841,
    n16842, n16843, n16844, n16845, n16846, n16847,
    n16848, n16849, n16850, n16851, n16852, n16853,
    n16854, n16855, n16856, n16857, n16858, n16859,
    n16860, n16861, n16862, n16863, n16864, n16865,
    n16866, n16867, n16868, n16869, n16870, n16871,
    n16872, n16873, n16874, n16875, n16876, n16877,
    n16878, n16879, n16880, n16882, n16883, n16884,
    n16885, n16886, n16887, n16888, n16889, n16890,
    n16891, n16892, n16893, n16894, n16895, n16896,
    n16897, n16898, n16899, n16900, n16901, n16902,
    n16903, n16904, n16905, n16906, n16907, n16908,
    n16909, n16910, n16911, n16912, n16913, n16914,
    n16915, n16916, n16917, n16918, n16919, n16920,
    n16921, n16922, n16923, n16924, n16925, n16926,
    n16927, n16928, n16929, n16930, n16931, n16932,
    n16933, n16934, n16935, n16936, n16937, n16938,
    n16939, n16940, n16941, n16942, n16943, n16944,
    n16945, n16946, n16947, n16948, n16949, n16950,
    n16951, n16952, n16953, n16954, n16955, n16956,
    n16957, n16958, n16959, n16960, n16961, n16962,
    n16963, n16964, n16965, n16966, n16967, n16968,
    n16969, n16970, n16971, n16972, n16973, n16974,
    n16975, n16976, n16977, n16978, n16979, n16980,
    n16981, n16982, n16983, n16984, n16985, n16986,
    n16987, n16988, n16989, n16990, n16991, n16992,
    n16993, n16994, n16995, n16996, n16997, n16998,
    n16999, n17000, n17001, n17002, n17003, n17004,
    n17005, n17006, n17007, n17008, n17009, n17010,
    n17011, n17012, n17013, n17014, n17015, n17016,
    n17017, n17018, n17019, n17020, n17021, n17022,
    n17023, n17024, n17025, n17026, n17027, n17028,
    n17029, n17030, n17031, n17032, n17033, n17034,
    n17035, n17036, n17037, n17038, n17039, n17040,
    n17041, n17042, n17043, n17044, n17045, n17046,
    n17047, n17048, n17049, n17050, n17051, n17052,
    n17053, n17054, n17055, n17056, n17057, n17058,
    n17059, n17060, n17061, n17062, n17063, n17064,
    n17065, n17066, n17067, n17068, n17069, n17070,
    n17071, n17072, n17073, n17074, n17075, n17076,
    n17077, n17078, n17079, n17080, n17081, n17082,
    n17083, n17084, n17085, n17086, n17087, n17088,
    n17089, n17090, n17091, n17092, n17093, n17094,
    n17095, n17096, n17097, n17098, n17099, n17100,
    n17101, n17102, n17103, n17104, n17105, n17106,
    n17107, n17108, n17109, n17110, n17111, n17112,
    n17113, n17114, n17115, n17116, n17117, n17118,
    n17119, n17120, n17121, n17122, n17123, n17124,
    n17125, n17126, n17127, n17128, n17129, n17130,
    n17131, n17132, n17133, n17134, n17135, n17136,
    n17137, n17138, n17139, n17140, n17141, n17142,
    n17143, n17144, n17145, n17146, n17147, n17148,
    n17149, n17150, n17151, n17152, n17153, n17154,
    n17155, n17156, n17157, n17158, n17159, n17160,
    n17161, n17162, n17163, n17164, n17165, n17166,
    n17167, n17168, n17169, n17170, n17171, n17172,
    n17173, n17174, n17175, n17176, n17177, n17178,
    n17179, n17180, n17181, n17182, n17183, n17184,
    n17185, n17186, n17187, n17188, n17189, n17190,
    n17191, n17192, n17193, n17194, n17195, n17196,
    n17197, n17198, n17199, n17200, n17201, n17202,
    n17203, n17204, n17205, n17206, n17207, n17208,
    n17209, n17210, n17211, n17212, n17213, n17214,
    n17215, n17216, n17217, n17218, n17219, n17220,
    n17221, n17222, n17223, n17224, n17225, n17226,
    n17227, n17228, n17229, n17230, n17231, n17232,
    n17233, n17234, n17235, n17236, n17237, n17238,
    n17239, n17240, n17241, n17242, n17243, n17244,
    n17245, n17246, n17247, n17248, n17249, n17250,
    n17251, n17252, n17253, n17254, n17255, n17256,
    n17257, n17258, n17259, n17260, n17261, n17262,
    n17263, n17264, n17265, n17266, n17267, n17268,
    n17269, n17270, n17271, n17272, n17273, n17274,
    n17275, n17276, n17277, n17278, n17279, n17280,
    n17281, n17282, n17283, n17284, n17285, n17286,
    n17287, n17288, n17289, n17290, n17291, n17292,
    n17293, n17294, n17295, n17296, n17297, n17298,
    n17299, n17300, n17301, n17302, n17303, n17304,
    n17305, n17306, n17307, n17308, n17309, n17310,
    n17311, n17312, n17313, n17314, n17315, n17316,
    n17317, n17318, n17319, n17320, n17321, n17322,
    n17323, n17324, n17325, n17326, n17327, n17328,
    n17329, n17330, n17331, n17332, n17333, n17334,
    n17335, n17336, n17337, n17338, n17339, n17340,
    n17341, n17342, n17343, n17344, n17345, n17346,
    n17347, n17348, n17349, n17350, n17351, n17352,
    n17353, n17354, n17355, n17356, n17357, n17358,
    n17359, n17360, n17361, n17362, n17363, n17364,
    n17365, n17366, n17367, n17368, n17369, n17370,
    n17371, n17372, n17373, n17374, n17375, n17376,
    n17377, n17378, n17379, n17380, n17381, n17382,
    n17383, n17384, n17385, n17386, n17387, n17388,
    n17389, n17390, n17391, n17392, n17393, n17394,
    n17395, n17396, n17397, n17398, n17399, n17400,
    n17401, n17402, n17403, n17404, n17405, n17406,
    n17407, n17408, n17409, n17410, n17411, n17412,
    n17413, n17414, n17415, n17416, n17417, n17418,
    n17419, n17420, n17421, n17422, n17423, n17424,
    n17425, n17426, n17427, n17428, n17429, n17430,
    n17431, n17433, n17434, n17435, n17436, n17437,
    n17438, n17439, n17440, n17441, n17442, n17443,
    n17444, n17445, n17446, n17447, n17448, n17449,
    n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461,
    n17462, n17463, n17464, n17465, n17466, n17467,
    n17468, n17469, n17470, n17471, n17472, n17473,
    n17474, n17475, n17476, n17477, n17478, n17479,
    n17480, n17481, n17482, n17483, n17484, n17485,
    n17486, n17487, n17488, n17489, n17490, n17491,
    n17492, n17493, n17494, n17495, n17496, n17497,
    n17498, n17499, n17500, n17501, n17502, n17503,
    n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515,
    n17516, n17517, n17518, n17519, n17520, n17521,
    n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533,
    n17534, n17535, n17536, n17537, n17538, n17539,
    n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551,
    n17552, n17553, n17554, n17555, n17556, n17557,
    n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569,
    n17570, n17571, n17572, n17573, n17574, n17575,
    n17576, n17577, n17578, n17579, n17580, n17581,
    n17582, n17583, n17584, n17585, n17586, n17587,
    n17588, n17589, n17590, n17591, n17592, n17593,
    n17594, n17595, n17596, n17597, n17598, n17599,
    n17600, n17601, n17602, n17603, n17604, n17605,
    n17606, n17607, n17608, n17609, n17610, n17611,
    n17612, n17613, n17614, n17615, n17616, n17617,
    n17618, n17619, n17620, n17621, n17622, n17623,
    n17624, n17625, n17626, n17627, n17628, n17629,
    n17630, n17631, n17632, n17633, n17634, n17635,
    n17636, n17637, n17638, n17639, n17640, n17641,
    n17642, n17643, n17644, n17645, n17646, n17647,
    n17648, n17649, n17650, n17651, n17652, n17653,
    n17654, n17655, n17656, n17657, n17658, n17659,
    n17660, n17661, n17662, n17663, n17664, n17665,
    n17666, n17667, n17668, n17669, n17670, n17671,
    n17672, n17673, n17674, n17675, n17676, n17677,
    n17678, n17679, n17680, n17681, n17682, n17683,
    n17684, n17685, n17686, n17687, n17688, n17689,
    n17690, n17691, n17692, n17693, n17694, n17695,
    n17696, n17697, n17698, n17699, n17700, n17701,
    n17702, n17703, n17704, n17705, n17706, n17707,
    n17708, n17709, n17710, n17711, n17712, n17713,
    n17714, n17715, n17716, n17717, n17718, n17719,
    n17720, n17721, n17722, n17723, n17724, n17725,
    n17726, n17727, n17728, n17729, n17730, n17731,
    n17732, n17733, n17734, n17735, n17736, n17737,
    n17738, n17739, n17740, n17741, n17742, n17743,
    n17744, n17745, n17746, n17747, n17748, n17749,
    n17750, n17751, n17752, n17753, n17754, n17755,
    n17756, n17757, n17758, n17759, n17760, n17761,
    n17762, n17763, n17764, n17765, n17766, n17767,
    n17768, n17769, n17770, n17771, n17772, n17773,
    n17774, n17775, n17776, n17777, n17778, n17779,
    n17780, n17781, n17782, n17783, n17784, n17785,
    n17786, n17787, n17788, n17789, n17790, n17791,
    n17792, n17793, n17794, n17795, n17796, n17797,
    n17798, n17799, n17800, n17801, n17802, n17803,
    n17804, n17805, n17806, n17807, n17808, n17809,
    n17810, n17811, n17812, n17813, n17814, n17815,
    n17816, n17817, n17818, n17819, n17820, n17821,
    n17822, n17823, n17824, n17825, n17826, n17827,
    n17828, n17829, n17830, n17831, n17832, n17833,
    n17834, n17835, n17836, n17837, n17838, n17839,
    n17840, n17841, n17842, n17843, n17844, n17845,
    n17846, n17847, n17848, n17849, n17850, n17851,
    n17852, n17853, n17854, n17855, n17856, n17857,
    n17858, n17859, n17860, n17861, n17862, n17863,
    n17864, n17865, n17866, n17867, n17868, n17869,
    n17870, n17871, n17872, n17873, n17874, n17875,
    n17876, n17877, n17878, n17879, n17880, n17881,
    n17882, n17883, n17884, n17885, n17886, n17887,
    n17888, n17889, n17890, n17891, n17892, n17893,
    n17894, n17895, n17896, n17897, n17898, n17899,
    n17900, n17901, n17902, n17903, n17904, n17905,
    n17906, n17907, n17908, n17909, n17910, n17911,
    n17912, n17913, n17914, n17915, n17916, n17917,
    n17918, n17919, n17920, n17921, n17922, n17923,
    n17924, n17925, n17926, n17927, n17928, n17929,
    n17930, n17931, n17932, n17933, n17934, n17935,
    n17936, n17937, n17938, n17939, n17940, n17941,
    n17942, n17943, n17944, n17945, n17946, n17947,
    n17948, n17949, n17950, n17951, n17952, n17953,
    n17954, n17955, n17956, n17957, n17958, n17959,
    n17960, n17961, n17962, n17963, n17964, n17965,
    n17966, n17967, n17968, n17969, n17970, n17971,
    n17972, n17973, n17974, n17975, n17976, n17977,
    n17978, n17979, n17980, n17981, n17982, n17983,
    n17984, n17985, n17986, n17987, n17988, n17989,
    n17990, n17991, n17992, n17993, n17994, n17995,
    n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014,
    n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032,
    n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050,
    n18051, n18052, n18053, n18054, n18055, n18056,
    n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068,
    n18069, n18070, n18071, n18072, n18073, n18074,
    n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086,
    n18087, n18088, n18089, n18090, n18091, n18092,
    n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104,
    n18105, n18106, n18107, n18108, n18109, n18110,
    n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122,
    n18123, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140,
    n18141, n18142, n18143, n18144, n18145, n18146,
    n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158,
    n18159, n18160, n18161, n18162, n18163, n18164,
    n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176,
    n18177, n18178, n18179, n18180, n18181, n18182,
    n18183, n18184, n18185, n18186, n18187, n18188,
    n18189, n18190, n18191, n18192, n18193, n18194,
    n18195, n18196, n18197, n18198, n18199, n18200,
    n18201, n18202, n18203, n18204, n18205, n18206,
    n18207, n18208, n18209, n18210, n18211, n18212,
    n18213, n18214, n18215, n18216, n18217, n18218,
    n18219, n18220, n18221, n18222, n18223, n18224,
    n18225, n18226, n18227, n18228, n18229, n18230,
    n18231, n18232, n18233, n18234, n18235, n18236,
    n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18248,
    n18249, n18250, n18251, n18252, n18253, n18254,
    n18255, n18256, n18257, n18258, n18259, n18260,
    n18261, n18262, n18263, n18264, n18265, n18266,
    n18267, n18268, n18269, n18270, n18271, n18272,
    n18273, n18274, n18275, n18276, n18277, n18278,
    n18279, n18280, n18281, n18282, n18283, n18284,
    n18285, n18286, n18287, n18288, n18289, n18290,
    n18291, n18292, n18293, n18294, n18295, n18296,
    n18297, n18298, n18299, n18300, n18301, n18302,
    n18303, n18304, n18305, n18306, n18307, n18308,
    n18309, n18310, n18311, n18312, n18313, n18314,
    n18315, n18316, n18317, n18318, n18319, n18320,
    n18321, n18322, n18323, n18324, n18325, n18326,
    n18327, n18328, n18329, n18330, n18331, n18332,
    n18333, n18334, n18335, n18336, n18337, n18338,
    n18339, n18340, n18341, n18342, n18343, n18344,
    n18345, n18346, n18347, n18348, n18349, n18350,
    n18351, n18352, n18353, n18354, n18355, n18356,
    n18357, n18358, n18359, n18360, n18361, n18362,
    n18363, n18364, n18365, n18366, n18367, n18368,
    n18369, n18370, n18371, n18372, n18373, n18374,
    n18375, n18376, n18377, n18378, n18379, n18380,
    n18381, n18382, n18383, n18384, n18385, n18386,
    n18387, n18388, n18389, n18390, n18391, n18392,
    n18393, n18394, n18395, n18396, n18397, n18398,
    n18399, n18400, n18401, n18402, n18403, n18404,
    n18405, n18406, n18407, n18408, n18409, n18410,
    n18411, n18412, n18413, n18414, n18415, n18416,
    n18417, n18418, n18419, n18420, n18421, n18422,
    n18423, n18424, n18425, n18426, n18427, n18428,
    n18429, n18430, n18431, n18432, n18433, n18434,
    n18435, n18436, n18437, n18438, n18439, n18440,
    n18441, n18442, n18443, n18444, n18445, n18446,
    n18447, n18448, n18449, n18450, n18451, n18452,
    n18453, n18454, n18455, n18456, n18457, n18458,
    n18459, n18460, n18461, n18462, n18463, n18464,
    n18465, n18466, n18467, n18468, n18469, n18470,
    n18471, n18472, n18473, n18474, n18475, n18476,
    n18477, n18478, n18479, n18480, n18481, n18482,
    n18483, n18484, n18485, n18486, n18487, n18488,
    n18489, n18490, n18491, n18492, n18493, n18494,
    n18495, n18496, n18497, n18498, n18499, n18500,
    n18501, n18502, n18503, n18504, n18505, n18506,
    n18507, n18508, n18509, n18510, n18511, n18512,
    n18513, n18514, n18515, n18516, n18517, n18518,
    n18519, n18520, n18521, n18522, n18523, n18524,
    n18525, n18526, n18527, n18528, n18529, n18530,
    n18531, n18532, n18533, n18534, n18535, n18536,
    n18537, n18538, n18539, n18540, n18541, n18542,
    n18543, n18544, n18545, n18546, n18547, n18548,
    n18549, n18550, n18551, n18552, n18553, n18554,
    n18555, n18556, n18557, n18558, n18559, n18560;
  assign po63  = pi126  | pi127 ;
  assign n194 = pi126  & pi127 ;
  assign n195 = ~pi124  & ~pi125 ;
  assign n196 = ~pi126  & ~n195;
  assign po62  = n194 | n196;
  assign n198 = ~pi124  & po62 ;
  assign n199 = pi125  & ~n198;
  assign n200 = n194 & n195;
  assign n201 = ~n199 & ~n200;
  assign n202 = pi124  & po62 ;
  assign n203 = ~pi122  & ~pi123 ;
  assign n204 = ~pi124  & n203;
  assign n205 = ~n202 & ~n204;
  assign n206 = n201 & ~n205;
  assign n207 = ~po63  & ~n206;
  assign n208 = ~n201 & n205;
  assign n209 = pi126  & n195;
  assign n210 = ~n196 & ~n209;
  assign n211 = pi127  & n210;
  assign n212 = ~n208 & ~n211;
  assign po61  = n207 | ~n212;
  assign n214 = n201 & ~n212;
  assign n215 = n205 & ~n214;
  assign n216 = po63  & ~n215;
  assign n217 = ~n206 & n216;
  assign n218 = po62  & ~po61 ;
  assign n219 = n203 & po61 ;
  assign n220 = ~n218 & ~n219;
  assign n221 = pi124  & ~n220;
  assign n222 = ~pi124  & n220;
  assign n223 = ~n221 & ~n222;
  assign n224 = ~pi120  & ~pi121 ;
  assign n225 = ~pi122  & ~n224;
  assign n226 = pi122  & ~po61 ;
  assign n227 = ~n225 & ~n226;
  assign n228 = ~po62  & ~n227;
  assign n229 = po62  & n227;
  assign n230 = ~pi122  & po61 ;
  assign n231 = pi123  & ~n230;
  assign n232 = ~n219 & ~n231;
  assign n233 = ~n229 & ~n232;
  assign n234 = ~n228 & ~n233;
  assign n235 = n223 & ~n234;
  assign n236 = ~n223 & n234;
  assign n237 = n206 & ~n212;
  assign n238 = ~n208 & ~n237;
  assign n239 = n236 & n238;
  assign n240 = ~po63  & ~n239;
  assign n241 = ~n235 & ~n240;
  assign n242 = ~n217 & n241;
  assign n243 = po61  & n242;
  assign n244 = ~n201 & ~po61 ;
  assign po60  = ~n242 | n244;
  assign n246 = n224 & po60 ;
  assign n247 = ~n243 & ~n246;
  assign n248 = pi122  & ~n247;
  assign n249 = ~pi122  & n247;
  assign n250 = ~n248 & ~n249;
  assign n251 = ~n223 & ~po60 ;
  assign n252 = po63  & ~n236;
  assign n253 = ~n235 & n252;
  assign n254 = po60  & ~n253;
  assign n255 = ~n251 & ~n254;
  assign n256 = pi120  & po60 ;
  assign n257 = ~pi118  & ~pi119 ;
  assign n258 = ~pi120  & n257;
  assign n259 = ~n256 & ~n258;
  assign n260 = po61  & ~n259;
  assign n261 = ~po61  & n259;
  assign n262 = ~pi120  & po60 ;
  assign n263 = pi121  & ~n262;
  assign n264 = ~n246 & ~n263;
  assign n265 = ~n261 & n264;
  assign n266 = ~n260 & ~n265;
  assign n267 = po62  & ~n266;
  assign n268 = ~po62  & n266;
  assign n269 = ~n250 & ~n268;
  assign n270 = ~n267 & ~n269;
  assign n271 = ~n228 & ~n229;
  assign n272 = po60  & n271;
  assign n273 = n232 & ~n272;
  assign n274 = ~n232 & n272;
  assign n275 = ~n273 & ~n274;
  assign n276 = n270 & n275;
  assign n277 = ~n270 & ~n275;
  assign n278 = n236 & po60 ;
  assign n279 = ~n235 & ~n278;
  assign n280 = n277 & n279;
  assign n281 = ~po63  & ~n280;
  assign n282 = ~n276 & ~n281;
  assign po59  = n255 | ~n282;
  assign n284 = ~n267 & ~n268;
  assign n285 = po59  & n284;
  assign n286 = ~n250 & ~n285;
  assign n287 = n250 & n285;
  assign n288 = ~n286 & ~n287;
  assign n289 = n275 & ~po59 ;
  assign n290 = ~n275 & ~po59 ;
  assign n291 = po63  & ~n290;
  assign n292 = ~n276 & n291;
  assign n293 = ~n277 & n292;
  assign n294 = pi118  & po59 ;
  assign n295 = ~pi116  & ~pi117 ;
  assign n296 = ~pi118  & n295;
  assign n297 = ~n294 & ~n296;
  assign n298 = po60  & ~n297;
  assign n299 = ~po60  & n297;
  assign n300 = ~pi118  & po59 ;
  assign n301 = pi119  & ~n300;
  assign n302 = n257 & po59 ;
  assign n303 = ~n301 & ~n302;
  assign n304 = ~n299 & n303;
  assign n305 = ~n298 & ~n304;
  assign n306 = po61  & ~n305;
  assign n307 = n254 & n282;
  assign n308 = ~n302 & ~n307;
  assign n309 = pi120  & ~n308;
  assign n310 = ~pi120  & n308;
  assign n311 = ~n309 & ~n310;
  assign n312 = ~po61  & n305;
  assign n313 = ~n311 & ~n312;
  assign n314 = ~n306 & ~n313;
  assign n315 = po62  & ~n314;
  assign n316 = ~po62  & n314;
  assign n317 = ~n260 & ~n261;
  assign n318 = po59  & n317;
  assign n319 = n264 & ~n318;
  assign n320 = ~n264 & n318;
  assign n321 = ~n319 & ~n320;
  assign n322 = ~n316 & ~n321;
  assign n323 = ~n315 & ~n322;
  assign n324 = n288 & n323;
  assign n325 = ~n288 & ~n323;
  assign n326 = n277 & po59 ;
  assign n327 = ~n276 & ~n326;
  assign n328 = n325 & n327;
  assign n329 = ~po63  & ~n328;
  assign n330 = ~n324 & ~n329;
  assign n331 = ~n293 & n330;
  assign po58  = n289 | ~n331;
  assign n333 = n288 & ~po58 ;
  assign n334 = ~n288 & po58 ;
  assign n335 = n323 & ~n334;
  assign n336 = po63  & ~n335;
  assign n337 = ~n325 & n336;
  assign n338 = pi116  & po58 ;
  assign n339 = ~pi114  & ~pi115 ;
  assign n340 = ~pi116  & n339;
  assign n341 = ~n338 & ~n340;
  assign n342 = po59  & ~n341;
  assign n343 = ~po59  & n341;
  assign n344 = ~pi116  & po58 ;
  assign n345 = pi117  & ~n344;
  assign n346 = n295 & po58 ;
  assign n347 = ~n345 & ~n346;
  assign n348 = ~n343 & n347;
  assign n349 = ~n342 & ~n348;
  assign n350 = po60  & ~n349;
  assign n351 = ~po60  & n349;
  assign n352 = po59  & n331;
  assign n353 = ~n346 & ~n352;
  assign n354 = pi118  & ~n353;
  assign n355 = ~pi118  & n353;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n351 & ~n356;
  assign n358 = ~n350 & ~n357;
  assign n359 = po61  & ~n358;
  assign n360 = ~po61  & n358;
  assign n361 = ~n298 & ~n299;
  assign n362 = po58  & n361;
  assign n363 = n303 & ~n362;
  assign n364 = ~n303 & n362;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~n360 & ~n365;
  assign n367 = ~n359 & ~n366;
  assign n368 = po62  & ~n367;
  assign n369 = ~n306 & ~n312;
  assign n370 = po58  & n369;
  assign n371 = ~n311 & ~n370;
  assign n372 = n311 & n370;
  assign n373 = ~n371 & ~n372;
  assign n374 = ~po62  & n367;
  assign n375 = ~n373 & ~n374;
  assign n376 = ~n368 & ~n375;
  assign n377 = ~n315 & ~n316;
  assign n378 = po58  & n377;
  assign n379 = n321 & n378;
  assign n380 = ~n321 & ~n378;
  assign n381 = ~n379 & ~n380;
  assign n382 = n376 & n381;
  assign n383 = ~n376 & ~n381;
  assign n384 = n325 & po58 ;
  assign n385 = ~n324 & ~n384;
  assign n386 = n383 & n385;
  assign n387 = ~po63  & ~n386;
  assign n388 = ~n382 & ~n387;
  assign n389 = ~n337 & n388;
  assign po57  = n333 | ~n389;
  assign n391 = n381 & ~po57 ;
  assign n392 = ~n381 & po57 ;
  assign n393 = n376 & ~n392;
  assign n394 = po63  & ~n393;
  assign n395 = ~n383 & n394;
  assign n396 = ~n368 & ~n374;
  assign n397 = po57  & n396;
  assign n398 = ~n373 & ~n397;
  assign n399 = n373 & n397;
  assign n400 = ~n398 & ~n399;
  assign n401 = pi114  & po57 ;
  assign n402 = ~pi112  & ~pi113 ;
  assign n403 = ~pi114  & n402;
  assign n404 = ~n401 & ~n403;
  assign n405 = po58  & ~n404;
  assign n406 = ~po58  & n404;
  assign n407 = ~pi114  & po57 ;
  assign n408 = pi115  & ~n407;
  assign n409 = n339 & po57 ;
  assign n410 = ~n408 & ~n409;
  assign n411 = ~n406 & n410;
  assign n412 = ~n405 & ~n411;
  assign n413 = po59  & ~n412;
  assign n414 = ~po59  & n412;
  assign n415 = po58  & n389;
  assign n416 = ~n409 & ~n415;
  assign n417 = pi116  & ~n416;
  assign n418 = ~pi116  & n416;
  assign n419 = ~n417 & ~n418;
  assign n420 = ~n414 & ~n419;
  assign n421 = ~n413 & ~n420;
  assign n422 = po60  & ~n421;
  assign n423 = ~po60  & n421;
  assign n424 = ~n342 & ~n343;
  assign n425 = po57  & n424;
  assign n426 = n347 & ~n425;
  assign n427 = ~n347 & n425;
  assign n428 = ~n426 & ~n427;
  assign n429 = ~n423 & ~n428;
  assign n430 = ~n422 & ~n429;
  assign n431 = po61  & ~n430;
  assign n432 = ~po61  & n430;
  assign n433 = ~n350 & ~n351;
  assign n434 = po57  & n433;
  assign n435 = ~n356 & ~n434;
  assign n436 = n356 & n434;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~n432 & ~n437;
  assign n439 = ~n431 & ~n438;
  assign n440 = po62  & ~n439;
  assign n441 = ~po62  & n439;
  assign n442 = ~n359 & ~n360;
  assign n443 = po57  & n442;
  assign n444 = n365 & n443;
  assign n445 = ~n365 & ~n443;
  assign n446 = ~n444 & ~n445;
  assign n447 = ~n441 & ~n446;
  assign n448 = ~n440 & ~n447;
  assign n449 = n400 & n448;
  assign n450 = ~n400 & ~n448;
  assign n451 = n383 & po57 ;
  assign n452 = ~n382 & ~n451;
  assign n453 = n450 & n452;
  assign n454 = ~po63  & ~n453;
  assign n455 = ~n449 & ~n454;
  assign n456 = ~n395 & n455;
  assign po56  = n391 | ~n456;
  assign n458 = ~pi112  & po56 ;
  assign n459 = pi113  & ~n458;
  assign n460 = n402 & po56 ;
  assign n461 = ~n459 & ~n460;
  assign n462 = n400 & ~po56 ;
  assign n463 = ~n400 & po56 ;
  assign n464 = n448 & ~n463;
  assign n465 = po63  & ~n464;
  assign n466 = ~n450 & n465;
  assign n467 = ~n440 & ~n441;
  assign n468 = po56  & n467;
  assign n469 = ~n446 & ~n468;
  assign n470 = n446 & n468;
  assign n471 = ~n469 & ~n470;
  assign n472 = pi112  & po56 ;
  assign n473 = ~pi110  & ~pi111 ;
  assign n474 = ~pi112  & n473;
  assign n475 = ~n472 & ~n474;
  assign n476 = po57  & ~n475;
  assign n477 = ~po57  & n475;
  assign n478 = n461 & ~n477;
  assign n479 = ~n476 & ~n478;
  assign n480 = po58  & ~n479;
  assign n481 = ~po58  & n479;
  assign n482 = po57  & n456;
  assign n483 = ~n460 & ~n482;
  assign n484 = pi114  & ~n483;
  assign n485 = ~pi114  & n483;
  assign n486 = ~n484 & ~n485;
  assign n487 = ~n481 & ~n486;
  assign n488 = ~n480 & ~n487;
  assign n489 = po59  & ~n488;
  assign n490 = ~po59  & n488;
  assign n491 = ~n405 & ~n406;
  assign n492 = po56  & n491;
  assign n493 = n410 & ~n492;
  assign n494 = ~n410 & n492;
  assign n495 = ~n493 & ~n494;
  assign n496 = ~n490 & ~n495;
  assign n497 = ~n489 & ~n496;
  assign n498 = po60  & ~n497;
  assign n499 = ~po60  & n497;
  assign n500 = ~n413 & ~n414;
  assign n501 = po56  & n500;
  assign n502 = ~n419 & ~n501;
  assign n503 = n419 & n501;
  assign n504 = ~n502 & ~n503;
  assign n505 = ~n499 & ~n504;
  assign n506 = ~n498 & ~n505;
  assign n507 = po61  & ~n506;
  assign n508 = ~po61  & n506;
  assign n509 = ~n422 & ~n423;
  assign n510 = po56  & n509;
  assign n511 = n428 & n510;
  assign n512 = ~n428 & ~n510;
  assign n513 = ~n511 & ~n512;
  assign n514 = ~n508 & ~n513;
  assign n515 = ~n507 & ~n514;
  assign n516 = po62  & ~n515;
  assign n517 = ~po62  & n515;
  assign n518 = ~n431 & ~n432;
  assign n519 = po56  & n518;
  assign n520 = ~n437 & ~n519;
  assign n521 = n437 & n519;
  assign n522 = ~n520 & ~n521;
  assign n523 = ~n517 & ~n522;
  assign n524 = ~n516 & ~n523;
  assign n525 = n471 & n524;
  assign n526 = ~n471 & ~n524;
  assign n527 = n450 & po56 ;
  assign n528 = ~n449 & ~n527;
  assign n529 = n526 & n528;
  assign n530 = ~po63  & ~n529;
  assign n531 = ~n525 & ~n530;
  assign n532 = ~n466 & n531;
  assign po55  = n462 | ~n532;
  assign n534 = ~n476 & ~n477;
  assign n535 = po55  & n534;
  assign n536 = n461 & ~n535;
  assign n537 = ~n461 & n535;
  assign n538 = ~n536 & ~n537;
  assign n539 = n471 & ~po55 ;
  assign n540 = ~n471 & po55 ;
  assign n541 = n524 & ~n540;
  assign n542 = po63  & ~n541;
  assign n543 = ~n526 & n542;
  assign n544 = ~n516 & ~n517;
  assign n545 = po55  & n544;
  assign n546 = ~n522 & ~n545;
  assign n547 = n522 & n545;
  assign n548 = ~n546 & ~n547;
  assign n549 = pi110  & po55 ;
  assign n550 = ~pi108  & ~pi109 ;
  assign n551 = ~pi110  & n550;
  assign n552 = ~n549 & ~n551;
  assign n553 = po56  & ~n552;
  assign n554 = ~po56  & n552;
  assign n555 = ~pi110  & po55 ;
  assign n556 = pi111  & ~n555;
  assign n557 = n473 & po55 ;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~n554 & n558;
  assign n560 = ~n553 & ~n559;
  assign n561 = po57  & ~n560;
  assign n562 = po56  & n532;
  assign n563 = ~n557 & ~n562;
  assign n564 = pi112  & ~n563;
  assign n565 = ~pi112  & n563;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~po57  & n560;
  assign n568 = ~n566 & ~n567;
  assign n569 = ~n561 & ~n568;
  assign n570 = po58  & ~n569;
  assign n571 = ~po58  & n569;
  assign n572 = ~n538 & ~n571;
  assign n573 = ~n570 & ~n572;
  assign n574 = po59  & ~n573;
  assign n575 = ~po59  & n573;
  assign n576 = ~n480 & ~n481;
  assign n577 = po55  & n576;
  assign n578 = ~n486 & ~n577;
  assign n579 = n486 & n577;
  assign n580 = ~n578 & ~n579;
  assign n581 = ~n575 & ~n580;
  assign n582 = ~n574 & ~n581;
  assign n583 = po60  & ~n582;
  assign n584 = ~po60  & n582;
  assign n585 = ~n489 & ~n490;
  assign n586 = po55  & n585;
  assign n587 = n495 & n586;
  assign n588 = ~n495 & ~n586;
  assign n589 = ~n587 & ~n588;
  assign n590 = ~n584 & ~n589;
  assign n591 = ~n583 & ~n590;
  assign n592 = po61  & ~n591;
  assign n593 = ~po61  & n591;
  assign n594 = ~n498 & ~n499;
  assign n595 = po55  & n594;
  assign n596 = ~n504 & ~n595;
  assign n597 = n504 & n595;
  assign n598 = ~n596 & ~n597;
  assign n599 = ~n593 & ~n598;
  assign n600 = ~n592 & ~n599;
  assign n601 = po62  & ~n600;
  assign n602 = ~po62  & n600;
  assign n603 = ~n507 & ~n508;
  assign n604 = po55  & n603;
  assign n605 = ~n513 & ~n604;
  assign n606 = n513 & n604;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~n602 & ~n607;
  assign n609 = ~n601 & ~n608;
  assign n610 = n548 & n609;
  assign n611 = ~n548 & ~n609;
  assign n612 = n526 & po55 ;
  assign n613 = ~n525 & ~n612;
  assign n614 = n611 & n613;
  assign n615 = ~po63  & ~n614;
  assign n616 = ~n610 & ~n615;
  assign n617 = ~n543 & n616;
  assign po54  = n539 | ~n617;
  assign n619 = ~n570 & ~n571;
  assign n620 = po54  & n619;
  assign n621 = n538 & n620;
  assign n622 = ~n538 & ~n620;
  assign n623 = ~n621 & ~n622;
  assign n624 = n548 & ~po54 ;
  assign n625 = ~n548 & po54 ;
  assign n626 = n609 & ~n625;
  assign n627 = po63  & ~n626;
  assign n628 = ~n611 & n627;
  assign n629 = ~n601 & ~n602;
  assign n630 = po54  & n629;
  assign n631 = ~n607 & ~n630;
  assign n632 = n607 & n630;
  assign n633 = ~n631 & ~n632;
  assign n634 = pi108  & po54 ;
  assign n635 = ~pi106  & ~pi107 ;
  assign n636 = ~pi108  & n635;
  assign n637 = ~n634 & ~n636;
  assign n638 = po55  & ~n637;
  assign n639 = ~po55  & n637;
  assign n640 = ~pi108  & po54 ;
  assign n641 = pi109  & ~n640;
  assign n642 = n550 & po54 ;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~n639 & n643;
  assign n645 = ~n638 & ~n644;
  assign n646 = po56  & ~n645;
  assign n647 = ~po56  & n645;
  assign n648 = po55  & n617;
  assign n649 = ~n642 & ~n648;
  assign n650 = pi110  & ~n649;
  assign n651 = ~pi110  & n649;
  assign n652 = ~n650 & ~n651;
  assign n653 = ~n647 & ~n652;
  assign n654 = ~n646 & ~n653;
  assign n655 = po57  & ~n654;
  assign n656 = ~po57  & n654;
  assign n657 = ~n553 & ~n554;
  assign n658 = po54  & n657;
  assign n659 = n558 & ~n658;
  assign n660 = ~n558 & n658;
  assign n661 = ~n659 & ~n660;
  assign n662 = ~n656 & ~n661;
  assign n663 = ~n655 & ~n662;
  assign n664 = po58  & ~n663;
  assign n665 = ~n561 & ~n567;
  assign n666 = po54  & n665;
  assign n667 = ~n566 & ~n666;
  assign n668 = n566 & n666;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~po58  & n663;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~n664 & ~n671;
  assign n673 = po59  & ~n672;
  assign n674 = ~po59  & n672;
  assign n675 = ~n623 & ~n674;
  assign n676 = ~n673 & ~n675;
  assign n677 = po60  & ~n676;
  assign n678 = ~po60  & n676;
  assign n679 = ~n574 & ~n575;
  assign n680 = po54  & n679;
  assign n681 = ~n580 & ~n680;
  assign n682 = n580 & n680;
  assign n683 = ~n681 & ~n682;
  assign n684 = ~n678 & ~n683;
  assign n685 = ~n677 & ~n684;
  assign n686 = po61  & ~n685;
  assign n687 = ~po61  & n685;
  assign n688 = ~n583 & ~n584;
  assign n689 = po54  & n688;
  assign n690 = ~n589 & ~n689;
  assign n691 = n589 & n689;
  assign n692 = ~n690 & ~n691;
  assign n693 = ~n687 & ~n692;
  assign n694 = ~n686 & ~n693;
  assign n695 = po62  & ~n694;
  assign n696 = ~po62  & n694;
  assign n697 = ~n592 & ~n593;
  assign n698 = po54  & n697;
  assign n699 = ~n598 & ~n698;
  assign n700 = n598 & n698;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n696 & ~n701;
  assign n703 = ~n695 & ~n702;
  assign n704 = n633 & n703;
  assign n705 = ~n633 & ~n703;
  assign n706 = n611 & po54 ;
  assign n707 = ~n610 & ~n706;
  assign n708 = n705 & n707;
  assign n709 = ~po63  & ~n708;
  assign n710 = ~n704 & ~n709;
  assign n711 = ~n628 & n710;
  assign po53  = n624 | ~n711;
  assign n713 = ~n673 & ~n674;
  assign n714 = po53  & n713;
  assign n715 = ~n623 & ~n714;
  assign n716 = n623 & n714;
  assign n717 = ~n715 & ~n716;
  assign n718 = n633 & ~po53 ;
  assign n719 = ~n633 & po53 ;
  assign n720 = n703 & ~n719;
  assign n721 = po63  & ~n720;
  assign n722 = ~n705 & n721;
  assign n723 = ~n695 & ~n696;
  assign n724 = po53  & n723;
  assign n725 = ~n701 & ~n724;
  assign n726 = n701 & n724;
  assign n727 = ~n725 & ~n726;
  assign n728 = pi106  & po53 ;
  assign n729 = ~pi104  & ~pi105 ;
  assign n730 = ~pi106  & n729;
  assign n731 = ~n728 & ~n730;
  assign n732 = po54  & ~n731;
  assign n733 = ~po54  & n731;
  assign n734 = ~pi106  & po53 ;
  assign n735 = pi107  & ~n734;
  assign n736 = n635 & po53 ;
  assign n737 = ~n735 & ~n736;
  assign n738 = ~n733 & n737;
  assign n739 = ~n732 & ~n738;
  assign n740 = po55  & ~n739;
  assign n741 = ~po55  & n739;
  assign n742 = po54  & n711;
  assign n743 = ~n736 & ~n742;
  assign n744 = pi108  & ~n743;
  assign n745 = ~pi108  & n743;
  assign n746 = ~n744 & ~n745;
  assign n747 = ~n741 & ~n746;
  assign n748 = ~n740 & ~n747;
  assign n749 = po56  & ~n748;
  assign n750 = ~po56  & n748;
  assign n751 = ~n638 & ~n639;
  assign n752 = po53  & n751;
  assign n753 = n643 & ~n752;
  assign n754 = ~n643 & n752;
  assign n755 = ~n753 & ~n754;
  assign n756 = ~n750 & ~n755;
  assign n757 = ~n749 & ~n756;
  assign n758 = po57  & ~n757;
  assign n759 = ~po57  & n757;
  assign n760 = ~n646 & ~n647;
  assign n761 = po53  & n760;
  assign n762 = ~n652 & ~n761;
  assign n763 = n652 & n761;
  assign n764 = ~n762 & ~n763;
  assign n765 = ~n759 & ~n764;
  assign n766 = ~n758 & ~n765;
  assign n767 = po58  & ~n766;
  assign n768 = ~po58  & n766;
  assign n769 = ~n655 & ~n656;
  assign n770 = po53  & n769;
  assign n771 = n661 & n770;
  assign n772 = ~n661 & ~n770;
  assign n773 = ~n771 & ~n772;
  assign n774 = ~n768 & ~n773;
  assign n775 = ~n767 & ~n774;
  assign n776 = po59  & ~n775;
  assign n777 = ~n664 & ~n670;
  assign n778 = po53  & n777;
  assign n779 = ~n669 & ~n778;
  assign n780 = n669 & n778;
  assign n781 = ~n779 & ~n780;
  assign n782 = ~po59  & n775;
  assign n783 = ~n781 & ~n782;
  assign n784 = ~n776 & ~n783;
  assign n785 = po60  & ~n784;
  assign n786 = ~po60  & n784;
  assign n787 = ~n717 & ~n786;
  assign n788 = ~n785 & ~n787;
  assign n789 = po61  & ~n788;
  assign n790 = ~po61  & n788;
  assign n791 = ~n677 & ~n678;
  assign n792 = po53  & n791;
  assign n793 = ~n683 & ~n792;
  assign n794 = n683 & n792;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~n790 & ~n795;
  assign n797 = ~n789 & ~n796;
  assign n798 = po62  & ~n797;
  assign n799 = ~po62  & n797;
  assign n800 = ~n686 & ~n687;
  assign n801 = po53  & n800;
  assign n802 = ~n692 & ~n801;
  assign n803 = n692 & n801;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~n799 & ~n804;
  assign n806 = ~n798 & ~n805;
  assign n807 = n727 & n806;
  assign n808 = ~n727 & ~n806;
  assign n809 = n705 & po53 ;
  assign n810 = ~n704 & ~n809;
  assign n811 = n808 & n810;
  assign n812 = ~po63  & ~n811;
  assign n813 = ~n807 & ~n812;
  assign n814 = ~n722 & n813;
  assign po52  = n718 | ~n814;
  assign n816 = ~n785 & ~n786;
  assign n817 = po52  & n816;
  assign n818 = ~n717 & ~n817;
  assign n819 = n717 & n817;
  assign n820 = ~n818 & ~n819;
  assign n821 = n727 & ~po52 ;
  assign n822 = ~n727 & po52 ;
  assign n823 = n806 & ~n822;
  assign n824 = po63  & ~n823;
  assign n825 = ~n808 & n824;
  assign n826 = ~n798 & ~n799;
  assign n827 = po52  & n826;
  assign n828 = ~n804 & ~n827;
  assign n829 = n804 & n827;
  assign n830 = ~n828 & ~n829;
  assign n831 = pi104  & po52 ;
  assign n832 = ~pi102  & ~pi103 ;
  assign n833 = ~pi104  & n832;
  assign n834 = ~n831 & ~n833;
  assign n835 = po53  & ~n834;
  assign n836 = ~po53  & n834;
  assign n837 = ~pi104  & po52 ;
  assign n838 = pi105  & ~n837;
  assign n839 = n729 & po52 ;
  assign n840 = ~n838 & ~n839;
  assign n841 = ~n836 & n840;
  assign n842 = ~n835 & ~n841;
  assign n843 = po54  & ~n842;
  assign n844 = ~po54  & n842;
  assign n845 = po53  & n814;
  assign n846 = ~n839 & ~n845;
  assign n847 = pi106  & ~n846;
  assign n848 = ~pi106  & n846;
  assign n849 = ~n847 & ~n848;
  assign n850 = ~n844 & ~n849;
  assign n851 = ~n843 & ~n850;
  assign n852 = po55  & ~n851;
  assign n853 = ~po55  & n851;
  assign n854 = ~n732 & ~n733;
  assign n855 = po52  & n854;
  assign n856 = n737 & ~n855;
  assign n857 = ~n737 & n855;
  assign n858 = ~n856 & ~n857;
  assign n859 = ~n853 & ~n858;
  assign n860 = ~n852 & ~n859;
  assign n861 = po56  & ~n860;
  assign n862 = ~po56  & n860;
  assign n863 = ~n740 & ~n741;
  assign n864 = po52  & n863;
  assign n865 = ~n746 & ~n864;
  assign n866 = n746 & n864;
  assign n867 = ~n865 & ~n866;
  assign n868 = ~n862 & ~n867;
  assign n869 = ~n861 & ~n868;
  assign n870 = po57  & ~n869;
  assign n871 = ~po57  & n869;
  assign n872 = ~n749 & ~n750;
  assign n873 = po52  & n872;
  assign n874 = n755 & n873;
  assign n875 = ~n755 & ~n873;
  assign n876 = ~n874 & ~n875;
  assign n877 = ~n871 & ~n876;
  assign n878 = ~n870 & ~n877;
  assign n879 = po58  & ~n878;
  assign n880 = ~po58  & n878;
  assign n881 = ~n758 & ~n759;
  assign n882 = po52  & n881;
  assign n883 = ~n764 & ~n882;
  assign n884 = n764 & n882;
  assign n885 = ~n883 & ~n884;
  assign n886 = ~n880 & ~n885;
  assign n887 = ~n879 & ~n886;
  assign n888 = po59  & ~n887;
  assign n889 = ~po59  & n887;
  assign n890 = ~n767 & ~n768;
  assign n891 = po52  & n890;
  assign n892 = ~n773 & ~n891;
  assign n893 = n773 & n891;
  assign n894 = ~n892 & ~n893;
  assign n895 = ~n889 & ~n894;
  assign n896 = ~n888 & ~n895;
  assign n897 = po60  & ~n896;
  assign n898 = ~n776 & ~n782;
  assign n899 = po52  & n898;
  assign n900 = ~n781 & ~n899;
  assign n901 = n781 & n899;
  assign n902 = ~n900 & ~n901;
  assign n903 = ~po60  & n896;
  assign n904 = ~n902 & ~n903;
  assign n905 = ~n897 & ~n904;
  assign n906 = po61  & ~n905;
  assign n907 = ~po61  & n905;
  assign n908 = ~n820 & ~n907;
  assign n909 = ~n906 & ~n908;
  assign n910 = po62  & ~n909;
  assign n911 = ~po62  & n909;
  assign n912 = ~n789 & ~n790;
  assign n913 = po52  & n912;
  assign n914 = ~n795 & ~n913;
  assign n915 = n795 & n913;
  assign n916 = ~n914 & ~n915;
  assign n917 = ~n911 & ~n916;
  assign n918 = ~n910 & ~n917;
  assign n919 = n830 & n918;
  assign n920 = ~n830 & ~n918;
  assign n921 = n808 & po52 ;
  assign n922 = ~n807 & ~n921;
  assign n923 = n920 & n922;
  assign n924 = ~po63  & ~n923;
  assign n925 = ~n919 & ~n924;
  assign n926 = ~n825 & n925;
  assign po51  = n821 | ~n926;
  assign n928 = ~n906 & ~n907;
  assign n929 = po51  & n928;
  assign n930 = ~n820 & ~n929;
  assign n931 = n820 & n929;
  assign n932 = ~n930 & ~n931;
  assign n933 = n830 & ~po51 ;
  assign n934 = ~n830 & po51 ;
  assign n935 = n918 & ~n934;
  assign n936 = po63  & ~n935;
  assign n937 = ~n920 & n936;
  assign n938 = ~n910 & ~n911;
  assign n939 = po51  & n938;
  assign n940 = ~n916 & ~n939;
  assign n941 = n916 & n939;
  assign n942 = ~n940 & ~n941;
  assign n943 = pi102  & po51 ;
  assign n944 = ~pi100  & ~pi101 ;
  assign n945 = ~pi102  & n944;
  assign n946 = ~n943 & ~n945;
  assign n947 = po52  & ~n946;
  assign n948 = ~po52  & n946;
  assign n949 = ~pi102  & po51 ;
  assign n950 = pi103  & ~n949;
  assign n951 = n832 & po51 ;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~n948 & n952;
  assign n954 = ~n947 & ~n953;
  assign n955 = po53  & ~n954;
  assign n956 = ~po53  & n954;
  assign n957 = po52  & n926;
  assign n958 = ~n951 & ~n957;
  assign n959 = pi104  & ~n958;
  assign n960 = ~pi104  & n958;
  assign n961 = ~n959 & ~n960;
  assign n962 = ~n956 & ~n961;
  assign n963 = ~n955 & ~n962;
  assign n964 = po54  & ~n963;
  assign n965 = ~po54  & n963;
  assign n966 = ~n835 & ~n836;
  assign n967 = po51  & n966;
  assign n968 = n840 & ~n967;
  assign n969 = ~n840 & n967;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~n965 & ~n970;
  assign n972 = ~n964 & ~n971;
  assign n973 = po55  & ~n972;
  assign n974 = ~po55  & n972;
  assign n975 = ~n843 & ~n844;
  assign n976 = po51  & n975;
  assign n977 = ~n849 & ~n976;
  assign n978 = n849 & n976;
  assign n979 = ~n977 & ~n978;
  assign n980 = ~n974 & ~n979;
  assign n981 = ~n973 & ~n980;
  assign n982 = po56  & ~n981;
  assign n983 = ~po56  & n981;
  assign n984 = ~n852 & ~n853;
  assign n985 = po51  & n984;
  assign n986 = n858 & n985;
  assign n987 = ~n858 & ~n985;
  assign n988 = ~n986 & ~n987;
  assign n989 = ~n983 & ~n988;
  assign n990 = ~n982 & ~n989;
  assign n991 = po57  & ~n990;
  assign n992 = ~po57  & n990;
  assign n993 = ~n861 & ~n862;
  assign n994 = po51  & n993;
  assign n995 = ~n867 & ~n994;
  assign n996 = n867 & n994;
  assign n997 = ~n995 & ~n996;
  assign n998 = ~n992 & ~n997;
  assign n999 = ~n991 & ~n998;
  assign n1000 = po58  & ~n999;
  assign n1001 = ~po58  & n999;
  assign n1002 = ~n870 & ~n871;
  assign n1003 = po51  & n1002;
  assign n1004 = ~n876 & ~n1003;
  assign n1005 = n876 & n1003;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~n1001 & ~n1006;
  assign n1008 = ~n1000 & ~n1007;
  assign n1009 = po59  & ~n1008;
  assign n1010 = ~po59  & n1008;
  assign n1011 = ~n879 & ~n880;
  assign n1012 = po51  & n1011;
  assign n1013 = ~n885 & ~n1012;
  assign n1014 = n885 & n1012;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = ~n1010 & ~n1015;
  assign n1017 = ~n1009 & ~n1016;
  assign n1018 = po60  & ~n1017;
  assign n1019 = ~po60  & n1017;
  assign n1020 = ~n888 & ~n889;
  assign n1021 = po51  & n1020;
  assign n1022 = ~n894 & ~n1021;
  assign n1023 = n894 & n1021;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = ~n1019 & ~n1024;
  assign n1026 = ~n1018 & ~n1025;
  assign n1027 = po61  & ~n1026;
  assign n1028 = ~n897 & ~n903;
  assign n1029 = po51  & n1028;
  assign n1030 = ~n902 & ~n1029;
  assign n1031 = n902 & n1029;
  assign n1032 = ~n1030 & ~n1031;
  assign n1033 = ~po61  & n1026;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = ~n1027 & ~n1034;
  assign n1036 = po62  & ~n1035;
  assign n1037 = ~po62  & n1035;
  assign n1038 = ~n932 & ~n1037;
  assign n1039 = ~n1036 & ~n1038;
  assign n1040 = n942 & n1039;
  assign n1041 = ~n942 & ~n1039;
  assign n1042 = n920 & po51 ;
  assign n1043 = ~n919 & ~n1042;
  assign n1044 = n1041 & n1043;
  assign n1045 = ~po63  & ~n1044;
  assign n1046 = ~n1040 & ~n1045;
  assign n1047 = ~n937 & n1046;
  assign po50  = n933 | ~n1047;
  assign n1049 = ~n1036 & ~n1037;
  assign n1050 = po50  & n1049;
  assign n1051 = ~n932 & ~n1050;
  assign n1052 = n932 & n1050;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = n942 & ~po50 ;
  assign n1055 = ~n942 & po50 ;
  assign n1056 = n1039 & ~n1055;
  assign n1057 = po63  & ~n1056;
  assign n1058 = ~n1041 & n1057;
  assign n1059 = pi100  & po50 ;
  assign n1060 = ~pi98  & ~pi99 ;
  assign n1061 = ~pi100  & n1060;
  assign n1062 = ~n1059 & ~n1061;
  assign n1063 = po51  & ~n1062;
  assign n1064 = ~po51  & n1062;
  assign n1065 = ~pi100  & po50 ;
  assign n1066 = pi101  & ~n1065;
  assign n1067 = n944 & po50 ;
  assign n1068 = ~n1066 & ~n1067;
  assign n1069 = ~n1064 & n1068;
  assign n1070 = ~n1063 & ~n1069;
  assign n1071 = po52  & ~n1070;
  assign n1072 = ~po52  & n1070;
  assign n1073 = po51  & n1047;
  assign n1074 = ~n1067 & ~n1073;
  assign n1075 = pi102  & ~n1074;
  assign n1076 = ~pi102  & n1074;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~n1072 & ~n1077;
  assign n1079 = ~n1071 & ~n1078;
  assign n1080 = po53  & ~n1079;
  assign n1081 = ~po53  & n1079;
  assign n1082 = ~n947 & ~n948;
  assign n1083 = po50  & n1082;
  assign n1084 = n952 & ~n1083;
  assign n1085 = ~n952 & n1083;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = ~n1081 & ~n1086;
  assign n1088 = ~n1080 & ~n1087;
  assign n1089 = po54  & ~n1088;
  assign n1090 = ~po54  & n1088;
  assign n1091 = ~n955 & ~n956;
  assign n1092 = po50  & n1091;
  assign n1093 = ~n961 & ~n1092;
  assign n1094 = n961 & n1092;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = ~n1090 & ~n1095;
  assign n1097 = ~n1089 & ~n1096;
  assign n1098 = po55  & ~n1097;
  assign n1099 = ~po55  & n1097;
  assign n1100 = ~n964 & ~n965;
  assign n1101 = po50  & n1100;
  assign n1102 = n970 & n1101;
  assign n1103 = ~n970 & ~n1101;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~n1099 & ~n1104;
  assign n1106 = ~n1098 & ~n1105;
  assign n1107 = po56  & ~n1106;
  assign n1108 = ~po56  & n1106;
  assign n1109 = ~n973 & ~n974;
  assign n1110 = po50  & n1109;
  assign n1111 = ~n979 & ~n1110;
  assign n1112 = n979 & n1110;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = ~n1108 & ~n1113;
  assign n1115 = ~n1107 & ~n1114;
  assign n1116 = po57  & ~n1115;
  assign n1117 = ~po57  & n1115;
  assign n1118 = ~n982 & ~n983;
  assign n1119 = po50  & n1118;
  assign n1120 = ~n988 & ~n1119;
  assign n1121 = n988 & n1119;
  assign n1122 = ~n1120 & ~n1121;
  assign n1123 = ~n1117 & ~n1122;
  assign n1124 = ~n1116 & ~n1123;
  assign n1125 = po58  & ~n1124;
  assign n1126 = ~po58  & n1124;
  assign n1127 = ~n991 & ~n992;
  assign n1128 = po50  & n1127;
  assign n1129 = ~n997 & ~n1128;
  assign n1130 = n997 & n1128;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = ~n1126 & ~n1131;
  assign n1133 = ~n1125 & ~n1132;
  assign n1134 = po59  & ~n1133;
  assign n1135 = ~po59  & n1133;
  assign n1136 = ~n1000 & ~n1001;
  assign n1137 = po50  & n1136;
  assign n1138 = ~n1006 & ~n1137;
  assign n1139 = n1006 & n1137;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = ~n1135 & ~n1140;
  assign n1142 = ~n1134 & ~n1141;
  assign n1143 = po60  & ~n1142;
  assign n1144 = ~po60  & n1142;
  assign n1145 = ~n1009 & ~n1010;
  assign n1146 = po50  & n1145;
  assign n1147 = ~n1015 & ~n1146;
  assign n1148 = n1015 & n1146;
  assign n1149 = ~n1147 & ~n1148;
  assign n1150 = ~n1144 & ~n1149;
  assign n1151 = ~n1143 & ~n1150;
  assign n1152 = po61  & ~n1151;
  assign n1153 = ~po61  & n1151;
  assign n1154 = ~n1018 & ~n1019;
  assign n1155 = po50  & n1154;
  assign n1156 = ~n1024 & ~n1155;
  assign n1157 = n1024 & n1155;
  assign n1158 = ~n1156 & ~n1157;
  assign n1159 = ~n1153 & ~n1158;
  assign n1160 = ~n1152 & ~n1159;
  assign n1161 = po62  & ~n1160;
  assign n1162 = ~n1027 & ~n1033;
  assign n1163 = po50  & n1162;
  assign n1164 = ~n1032 & ~n1163;
  assign n1165 = n1032 & n1163;
  assign n1166 = ~n1164 & ~n1165;
  assign n1167 = ~po62  & n1160;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = ~n1161 & ~n1168;
  assign n1170 = n1053 & n1169;
  assign n1171 = ~n1053 & ~n1169;
  assign n1172 = n1041 & po50 ;
  assign n1173 = ~n1040 & ~n1172;
  assign n1174 = n1171 & n1173;
  assign n1175 = ~po63  & ~n1174;
  assign n1176 = ~n1170 & ~n1175;
  assign n1177 = ~n1058 & n1176;
  assign po49  = n1054 | ~n1177;
  assign n1179 = n1053 & ~po49 ;
  assign n1180 = ~n1053 & po49 ;
  assign n1181 = n1169 & ~n1180;
  assign n1182 = po63  & ~n1181;
  assign n1183 = ~n1171 & n1182;
  assign n1184 = ~n1161 & ~n1167;
  assign n1185 = po49  & n1184;
  assign n1186 = ~n1166 & ~n1185;
  assign n1187 = n1166 & n1185;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = pi98  & po49 ;
  assign n1190 = ~pi96  & ~pi97 ;
  assign n1191 = ~pi98  & n1190;
  assign n1192 = ~n1189 & ~n1191;
  assign n1193 = po50  & ~n1192;
  assign n1194 = ~po50  & n1192;
  assign n1195 = ~pi98  & po49 ;
  assign n1196 = pi99  & ~n1195;
  assign n1197 = n1060 & po49 ;
  assign n1198 = ~n1196 & ~n1197;
  assign n1199 = ~n1194 & n1198;
  assign n1200 = ~n1193 & ~n1199;
  assign n1201 = po51  & ~n1200;
  assign n1202 = ~po51  & n1200;
  assign n1203 = po50  & n1177;
  assign n1204 = ~n1197 & ~n1203;
  assign n1205 = pi100  & ~n1204;
  assign n1206 = ~pi100  & n1204;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = ~n1202 & ~n1207;
  assign n1209 = ~n1201 & ~n1208;
  assign n1210 = po52  & ~n1209;
  assign n1211 = ~po52  & n1209;
  assign n1212 = ~n1063 & ~n1064;
  assign n1213 = po49  & n1212;
  assign n1214 = n1068 & ~n1213;
  assign n1215 = ~n1068 & n1213;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1211 & ~n1216;
  assign n1218 = ~n1210 & ~n1217;
  assign n1219 = po53  & ~n1218;
  assign n1220 = ~po53  & n1218;
  assign n1221 = ~n1071 & ~n1072;
  assign n1222 = po49  & n1221;
  assign n1223 = ~n1077 & ~n1222;
  assign n1224 = n1077 & n1222;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = ~n1220 & ~n1225;
  assign n1227 = ~n1219 & ~n1226;
  assign n1228 = po54  & ~n1227;
  assign n1229 = ~po54  & n1227;
  assign n1230 = ~n1080 & ~n1081;
  assign n1231 = po49  & n1230;
  assign n1232 = n1086 & n1231;
  assign n1233 = ~n1086 & ~n1231;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = ~n1229 & ~n1234;
  assign n1236 = ~n1228 & ~n1235;
  assign n1237 = po55  & ~n1236;
  assign n1238 = ~po55  & n1236;
  assign n1239 = ~n1089 & ~n1090;
  assign n1240 = po49  & n1239;
  assign n1241 = ~n1095 & ~n1240;
  assign n1242 = n1095 & n1240;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = ~n1238 & ~n1243;
  assign n1245 = ~n1237 & ~n1244;
  assign n1246 = po56  & ~n1245;
  assign n1247 = ~po56  & n1245;
  assign n1248 = ~n1098 & ~n1099;
  assign n1249 = po49  & n1248;
  assign n1250 = ~n1104 & ~n1249;
  assign n1251 = n1104 & n1249;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = ~n1247 & ~n1252;
  assign n1254 = ~n1246 & ~n1253;
  assign n1255 = po57  & ~n1254;
  assign n1256 = ~po57  & n1254;
  assign n1257 = ~n1107 & ~n1108;
  assign n1258 = po49  & n1257;
  assign n1259 = ~n1113 & ~n1258;
  assign n1260 = n1113 & n1258;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = ~n1256 & ~n1261;
  assign n1263 = ~n1255 & ~n1262;
  assign n1264 = po58  & ~n1263;
  assign n1265 = ~po58  & n1263;
  assign n1266 = ~n1116 & ~n1117;
  assign n1267 = po49  & n1266;
  assign n1268 = ~n1122 & ~n1267;
  assign n1269 = n1122 & n1267;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = ~n1265 & ~n1270;
  assign n1272 = ~n1264 & ~n1271;
  assign n1273 = po59  & ~n1272;
  assign n1274 = ~po59  & n1272;
  assign n1275 = ~n1125 & ~n1126;
  assign n1276 = po49  & n1275;
  assign n1277 = ~n1131 & ~n1276;
  assign n1278 = n1131 & n1276;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = ~n1274 & ~n1279;
  assign n1281 = ~n1273 & ~n1280;
  assign n1282 = po60  & ~n1281;
  assign n1283 = ~po60  & n1281;
  assign n1284 = ~n1134 & ~n1135;
  assign n1285 = po49  & n1284;
  assign n1286 = ~n1140 & ~n1285;
  assign n1287 = n1140 & n1285;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = ~n1283 & ~n1288;
  assign n1290 = ~n1282 & ~n1289;
  assign n1291 = po61  & ~n1290;
  assign n1292 = ~po61  & n1290;
  assign n1293 = ~n1143 & ~n1144;
  assign n1294 = po49  & n1293;
  assign n1295 = ~n1149 & ~n1294;
  assign n1296 = n1149 & n1294;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = ~n1292 & ~n1297;
  assign n1299 = ~n1291 & ~n1298;
  assign n1300 = po62  & ~n1299;
  assign n1301 = ~po62  & n1299;
  assign n1302 = ~n1152 & ~n1153;
  assign n1303 = po49  & n1302;
  assign n1304 = ~n1158 & ~n1303;
  assign n1305 = n1158 & n1303;
  assign n1306 = ~n1304 & ~n1305;
  assign n1307 = ~n1301 & ~n1306;
  assign n1308 = ~n1300 & ~n1307;
  assign n1309 = n1188 & n1308;
  assign n1310 = ~n1188 & ~n1308;
  assign n1311 = n1171 & po49 ;
  assign n1312 = ~n1170 & ~n1311;
  assign n1313 = n1310 & n1312;
  assign n1314 = ~po63  & ~n1313;
  assign n1315 = ~n1309 & ~n1314;
  assign n1316 = ~n1183 & n1315;
  assign po48  = n1179 | ~n1316;
  assign n1318 = ~pi96  & po48 ;
  assign n1319 = pi97  & ~n1318;
  assign n1320 = n1190 & po48 ;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = n1188 & ~po48 ;
  assign n1323 = ~n1188 & po48 ;
  assign n1324 = n1308 & ~n1323;
  assign n1325 = po63  & ~n1324;
  assign n1326 = ~n1310 & n1325;
  assign n1327 = ~n1300 & ~n1301;
  assign n1328 = po48  & n1327;
  assign n1329 = ~n1306 & ~n1328;
  assign n1330 = n1306 & n1328;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = pi96  & po48 ;
  assign n1333 = ~pi94  & ~pi95 ;
  assign n1334 = ~pi96  & n1333;
  assign n1335 = ~n1332 & ~n1334;
  assign n1336 = po49  & ~n1335;
  assign n1337 = ~po49  & n1335;
  assign n1338 = n1321 & ~n1337;
  assign n1339 = ~n1336 & ~n1338;
  assign n1340 = po50  & ~n1339;
  assign n1341 = ~po50  & n1339;
  assign n1342 = po49  & n1316;
  assign n1343 = ~n1320 & ~n1342;
  assign n1344 = pi98  & ~n1343;
  assign n1345 = ~pi98  & n1343;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = ~n1341 & ~n1346;
  assign n1348 = ~n1340 & ~n1347;
  assign n1349 = po51  & ~n1348;
  assign n1350 = ~po51  & n1348;
  assign n1351 = ~n1193 & ~n1194;
  assign n1352 = po48  & n1351;
  assign n1353 = n1198 & ~n1352;
  assign n1354 = ~n1198 & n1352;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = ~n1350 & ~n1355;
  assign n1357 = ~n1349 & ~n1356;
  assign n1358 = po52  & ~n1357;
  assign n1359 = ~po52  & n1357;
  assign n1360 = ~n1201 & ~n1202;
  assign n1361 = po48  & n1360;
  assign n1362 = ~n1207 & ~n1361;
  assign n1363 = n1207 & n1361;
  assign n1364 = ~n1362 & ~n1363;
  assign n1365 = ~n1359 & ~n1364;
  assign n1366 = ~n1358 & ~n1365;
  assign n1367 = po53  & ~n1366;
  assign n1368 = ~po53  & n1366;
  assign n1369 = ~n1210 & ~n1211;
  assign n1370 = po48  & n1369;
  assign n1371 = n1216 & n1370;
  assign n1372 = ~n1216 & ~n1370;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = ~n1368 & ~n1373;
  assign n1375 = ~n1367 & ~n1374;
  assign n1376 = po54  & ~n1375;
  assign n1377 = ~po54  & n1375;
  assign n1378 = ~n1219 & ~n1220;
  assign n1379 = po48  & n1378;
  assign n1380 = ~n1225 & ~n1379;
  assign n1381 = n1225 & n1379;
  assign n1382 = ~n1380 & ~n1381;
  assign n1383 = ~n1377 & ~n1382;
  assign n1384 = ~n1376 & ~n1383;
  assign n1385 = po55  & ~n1384;
  assign n1386 = ~po55  & n1384;
  assign n1387 = ~n1228 & ~n1229;
  assign n1388 = po48  & n1387;
  assign n1389 = ~n1234 & ~n1388;
  assign n1390 = n1234 & n1388;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = ~n1386 & ~n1391;
  assign n1393 = ~n1385 & ~n1392;
  assign n1394 = po56  & ~n1393;
  assign n1395 = ~po56  & n1393;
  assign n1396 = ~n1237 & ~n1238;
  assign n1397 = po48  & n1396;
  assign n1398 = ~n1243 & ~n1397;
  assign n1399 = n1243 & n1397;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = ~n1395 & ~n1400;
  assign n1402 = ~n1394 & ~n1401;
  assign n1403 = po57  & ~n1402;
  assign n1404 = ~po57  & n1402;
  assign n1405 = ~n1246 & ~n1247;
  assign n1406 = po48  & n1405;
  assign n1407 = ~n1252 & ~n1406;
  assign n1408 = n1252 & n1406;
  assign n1409 = ~n1407 & ~n1408;
  assign n1410 = ~n1404 & ~n1409;
  assign n1411 = ~n1403 & ~n1410;
  assign n1412 = po58  & ~n1411;
  assign n1413 = ~po58  & n1411;
  assign n1414 = ~n1255 & ~n1256;
  assign n1415 = po48  & n1414;
  assign n1416 = ~n1261 & ~n1415;
  assign n1417 = n1261 & n1415;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = ~n1413 & ~n1418;
  assign n1420 = ~n1412 & ~n1419;
  assign n1421 = po59  & ~n1420;
  assign n1422 = ~po59  & n1420;
  assign n1423 = ~n1264 & ~n1265;
  assign n1424 = po48  & n1423;
  assign n1425 = ~n1270 & ~n1424;
  assign n1426 = n1270 & n1424;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~n1422 & ~n1427;
  assign n1429 = ~n1421 & ~n1428;
  assign n1430 = po60  & ~n1429;
  assign n1431 = ~po60  & n1429;
  assign n1432 = ~n1273 & ~n1274;
  assign n1433 = po48  & n1432;
  assign n1434 = ~n1279 & ~n1433;
  assign n1435 = n1279 & n1433;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = ~n1431 & ~n1436;
  assign n1438 = ~n1430 & ~n1437;
  assign n1439 = po61  & ~n1438;
  assign n1440 = ~po61  & n1438;
  assign n1441 = ~n1282 & ~n1283;
  assign n1442 = po48  & n1441;
  assign n1443 = ~n1288 & ~n1442;
  assign n1444 = n1288 & n1442;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = ~n1440 & ~n1445;
  assign n1447 = ~n1439 & ~n1446;
  assign n1448 = po62  & ~n1447;
  assign n1449 = ~po62  & n1447;
  assign n1450 = ~n1291 & ~n1292;
  assign n1451 = po48  & n1450;
  assign n1452 = ~n1297 & ~n1451;
  assign n1453 = n1297 & n1451;
  assign n1454 = ~n1452 & ~n1453;
  assign n1455 = ~n1449 & ~n1454;
  assign n1456 = ~n1448 & ~n1455;
  assign n1457 = n1331 & n1456;
  assign n1458 = ~n1331 & ~n1456;
  assign n1459 = n1310 & po48 ;
  assign n1460 = ~n1309 & ~n1459;
  assign n1461 = n1458 & n1460;
  assign n1462 = ~po63  & ~n1461;
  assign n1463 = ~n1457 & ~n1462;
  assign n1464 = ~n1326 & n1463;
  assign po47  = n1322 | ~n1464;
  assign n1466 = ~n1336 & ~n1337;
  assign n1467 = po47  & n1466;
  assign n1468 = n1321 & ~n1467;
  assign n1469 = ~n1321 & n1467;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = n1331 & ~po47 ;
  assign n1472 = ~n1331 & po47 ;
  assign n1473 = n1456 & ~n1472;
  assign n1474 = po63  & ~n1473;
  assign n1475 = ~n1458 & n1474;
  assign n1476 = ~n1448 & ~n1449;
  assign n1477 = po47  & n1476;
  assign n1478 = ~n1454 & ~n1477;
  assign n1479 = n1454 & n1477;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = pi94  & po47 ;
  assign n1482 = ~pi92  & ~pi93 ;
  assign n1483 = ~pi94  & n1482;
  assign n1484 = ~n1481 & ~n1483;
  assign n1485 = po48  & ~n1484;
  assign n1486 = ~po48  & n1484;
  assign n1487 = ~pi94  & po47 ;
  assign n1488 = pi95  & ~n1487;
  assign n1489 = n1333 & po47 ;
  assign n1490 = ~n1488 & ~n1489;
  assign n1491 = ~n1486 & n1490;
  assign n1492 = ~n1485 & ~n1491;
  assign n1493 = po49  & ~n1492;
  assign n1494 = po48  & n1464;
  assign n1495 = ~n1489 & ~n1494;
  assign n1496 = pi96  & ~n1495;
  assign n1497 = ~pi96  & n1495;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = ~po49  & n1492;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = ~n1493 & ~n1500;
  assign n1502 = po50  & ~n1501;
  assign n1503 = ~po50  & n1501;
  assign n1504 = ~n1470 & ~n1503;
  assign n1505 = ~n1502 & ~n1504;
  assign n1506 = po51  & ~n1505;
  assign n1507 = ~po51  & n1505;
  assign n1508 = ~n1340 & ~n1341;
  assign n1509 = po47  & n1508;
  assign n1510 = ~n1346 & ~n1509;
  assign n1511 = n1346 & n1509;
  assign n1512 = ~n1510 & ~n1511;
  assign n1513 = ~n1507 & ~n1512;
  assign n1514 = ~n1506 & ~n1513;
  assign n1515 = po52  & ~n1514;
  assign n1516 = ~po52  & n1514;
  assign n1517 = ~n1349 & ~n1350;
  assign n1518 = po47  & n1517;
  assign n1519 = n1355 & n1518;
  assign n1520 = ~n1355 & ~n1518;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = ~n1516 & ~n1521;
  assign n1523 = ~n1515 & ~n1522;
  assign n1524 = po53  & ~n1523;
  assign n1525 = ~po53  & n1523;
  assign n1526 = ~n1358 & ~n1359;
  assign n1527 = po47  & n1526;
  assign n1528 = ~n1364 & ~n1527;
  assign n1529 = n1364 & n1527;
  assign n1530 = ~n1528 & ~n1529;
  assign n1531 = ~n1525 & ~n1530;
  assign n1532 = ~n1524 & ~n1531;
  assign n1533 = po54  & ~n1532;
  assign n1534 = ~po54  & n1532;
  assign n1535 = ~n1367 & ~n1368;
  assign n1536 = po47  & n1535;
  assign n1537 = ~n1373 & ~n1536;
  assign n1538 = n1373 & n1536;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = ~n1534 & ~n1539;
  assign n1541 = ~n1533 & ~n1540;
  assign n1542 = po55  & ~n1541;
  assign n1543 = ~po55  & n1541;
  assign n1544 = ~n1376 & ~n1377;
  assign n1545 = po47  & n1544;
  assign n1546 = ~n1382 & ~n1545;
  assign n1547 = n1382 & n1545;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = ~n1543 & ~n1548;
  assign n1550 = ~n1542 & ~n1549;
  assign n1551 = po56  & ~n1550;
  assign n1552 = ~po56  & n1550;
  assign n1553 = ~n1385 & ~n1386;
  assign n1554 = po47  & n1553;
  assign n1555 = ~n1391 & ~n1554;
  assign n1556 = n1391 & n1554;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = ~n1552 & ~n1557;
  assign n1559 = ~n1551 & ~n1558;
  assign n1560 = po57  & ~n1559;
  assign n1561 = ~po57  & n1559;
  assign n1562 = ~n1394 & ~n1395;
  assign n1563 = po47  & n1562;
  assign n1564 = ~n1400 & ~n1563;
  assign n1565 = n1400 & n1563;
  assign n1566 = ~n1564 & ~n1565;
  assign n1567 = ~n1561 & ~n1566;
  assign n1568 = ~n1560 & ~n1567;
  assign n1569 = po58  & ~n1568;
  assign n1570 = ~po58  & n1568;
  assign n1571 = ~n1403 & ~n1404;
  assign n1572 = po47  & n1571;
  assign n1573 = ~n1409 & ~n1572;
  assign n1574 = n1409 & n1572;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = ~n1570 & ~n1575;
  assign n1577 = ~n1569 & ~n1576;
  assign n1578 = po59  & ~n1577;
  assign n1579 = ~po59  & n1577;
  assign n1580 = ~n1412 & ~n1413;
  assign n1581 = po47  & n1580;
  assign n1582 = ~n1418 & ~n1581;
  assign n1583 = n1418 & n1581;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = ~n1579 & ~n1584;
  assign n1586 = ~n1578 & ~n1585;
  assign n1587 = po60  & ~n1586;
  assign n1588 = ~po60  & n1586;
  assign n1589 = ~n1421 & ~n1422;
  assign n1590 = po47  & n1589;
  assign n1591 = ~n1427 & ~n1590;
  assign n1592 = n1427 & n1590;
  assign n1593 = ~n1591 & ~n1592;
  assign n1594 = ~n1588 & ~n1593;
  assign n1595 = ~n1587 & ~n1594;
  assign n1596 = po61  & ~n1595;
  assign n1597 = ~po61  & n1595;
  assign n1598 = ~n1430 & ~n1431;
  assign n1599 = po47  & n1598;
  assign n1600 = ~n1436 & ~n1599;
  assign n1601 = n1436 & n1599;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = ~n1597 & ~n1602;
  assign n1604 = ~n1596 & ~n1603;
  assign n1605 = po62  & ~n1604;
  assign n1606 = ~po62  & n1604;
  assign n1607 = ~n1439 & ~n1440;
  assign n1608 = po47  & n1607;
  assign n1609 = ~n1445 & ~n1608;
  assign n1610 = n1445 & n1608;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = ~n1606 & ~n1611;
  assign n1613 = ~n1605 & ~n1612;
  assign n1614 = n1480 & n1613;
  assign n1615 = ~n1480 & ~n1613;
  assign n1616 = n1458 & po47 ;
  assign n1617 = ~n1457 & ~n1616;
  assign n1618 = n1615 & n1617;
  assign n1619 = ~po63  & ~n1618;
  assign n1620 = ~n1614 & ~n1619;
  assign n1621 = ~n1475 & n1620;
  assign po46  = n1471 | ~n1621;
  assign n1623 = ~n1502 & ~n1503;
  assign n1624 = po46  & n1623;
  assign n1625 = n1470 & n1624;
  assign n1626 = ~n1470 & ~n1624;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = n1480 & ~po46 ;
  assign n1629 = ~n1480 & po46 ;
  assign n1630 = n1613 & ~n1629;
  assign n1631 = po63  & ~n1630;
  assign n1632 = ~n1615 & n1631;
  assign n1633 = ~n1605 & ~n1606;
  assign n1634 = po46  & n1633;
  assign n1635 = ~n1611 & ~n1634;
  assign n1636 = n1611 & n1634;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = pi92  & po46 ;
  assign n1639 = ~pi90  & ~pi91 ;
  assign n1640 = ~pi92  & n1639;
  assign n1641 = ~n1638 & ~n1640;
  assign n1642 = po47  & ~n1641;
  assign n1643 = ~po47  & n1641;
  assign n1644 = ~pi92  & po46 ;
  assign n1645 = pi93  & ~n1644;
  assign n1646 = n1482 & po46 ;
  assign n1647 = ~n1645 & ~n1646;
  assign n1648 = ~n1643 & n1647;
  assign n1649 = ~n1642 & ~n1648;
  assign n1650 = po48  & ~n1649;
  assign n1651 = ~po48  & n1649;
  assign n1652 = po47  & n1621;
  assign n1653 = ~n1646 & ~n1652;
  assign n1654 = pi94  & ~n1653;
  assign n1655 = ~pi94  & n1653;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = ~n1651 & ~n1656;
  assign n1658 = ~n1650 & ~n1657;
  assign n1659 = po49  & ~n1658;
  assign n1660 = ~po49  & n1658;
  assign n1661 = ~n1485 & ~n1486;
  assign n1662 = po46  & n1661;
  assign n1663 = n1490 & ~n1662;
  assign n1664 = ~n1490 & n1662;
  assign n1665 = ~n1663 & ~n1664;
  assign n1666 = ~n1660 & ~n1665;
  assign n1667 = ~n1659 & ~n1666;
  assign n1668 = po50  & ~n1667;
  assign n1669 = ~n1493 & ~n1499;
  assign n1670 = po46  & n1669;
  assign n1671 = ~n1498 & ~n1670;
  assign n1672 = n1498 & n1670;
  assign n1673 = ~n1671 & ~n1672;
  assign n1674 = ~po50  & n1667;
  assign n1675 = ~n1673 & ~n1674;
  assign n1676 = ~n1668 & ~n1675;
  assign n1677 = po51  & ~n1676;
  assign n1678 = ~po51  & n1676;
  assign n1679 = ~n1627 & ~n1678;
  assign n1680 = ~n1677 & ~n1679;
  assign n1681 = po52  & ~n1680;
  assign n1682 = ~po52  & n1680;
  assign n1683 = ~n1506 & ~n1507;
  assign n1684 = po46  & n1683;
  assign n1685 = ~n1512 & ~n1684;
  assign n1686 = n1512 & n1684;
  assign n1687 = ~n1685 & ~n1686;
  assign n1688 = ~n1682 & ~n1687;
  assign n1689 = ~n1681 & ~n1688;
  assign n1690 = po53  & ~n1689;
  assign n1691 = ~po53  & n1689;
  assign n1692 = ~n1515 & ~n1516;
  assign n1693 = po46  & n1692;
  assign n1694 = ~n1521 & ~n1693;
  assign n1695 = n1521 & n1693;
  assign n1696 = ~n1694 & ~n1695;
  assign n1697 = ~n1691 & ~n1696;
  assign n1698 = ~n1690 & ~n1697;
  assign n1699 = po54  & ~n1698;
  assign n1700 = ~po54  & n1698;
  assign n1701 = ~n1524 & ~n1525;
  assign n1702 = po46  & n1701;
  assign n1703 = ~n1530 & ~n1702;
  assign n1704 = n1530 & n1702;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = ~n1700 & ~n1705;
  assign n1707 = ~n1699 & ~n1706;
  assign n1708 = po55  & ~n1707;
  assign n1709 = ~po55  & n1707;
  assign n1710 = ~n1533 & ~n1534;
  assign n1711 = po46  & n1710;
  assign n1712 = ~n1539 & ~n1711;
  assign n1713 = n1539 & n1711;
  assign n1714 = ~n1712 & ~n1713;
  assign n1715 = ~n1709 & ~n1714;
  assign n1716 = ~n1708 & ~n1715;
  assign n1717 = po56  & ~n1716;
  assign n1718 = ~po56  & n1716;
  assign n1719 = ~n1542 & ~n1543;
  assign n1720 = po46  & n1719;
  assign n1721 = ~n1548 & ~n1720;
  assign n1722 = n1548 & n1720;
  assign n1723 = ~n1721 & ~n1722;
  assign n1724 = ~n1718 & ~n1723;
  assign n1725 = ~n1717 & ~n1724;
  assign n1726 = po57  & ~n1725;
  assign n1727 = ~po57  & n1725;
  assign n1728 = ~n1551 & ~n1552;
  assign n1729 = po46  & n1728;
  assign n1730 = ~n1557 & ~n1729;
  assign n1731 = n1557 & n1729;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = ~n1727 & ~n1732;
  assign n1734 = ~n1726 & ~n1733;
  assign n1735 = po58  & ~n1734;
  assign n1736 = ~po58  & n1734;
  assign n1737 = ~n1560 & ~n1561;
  assign n1738 = po46  & n1737;
  assign n1739 = ~n1566 & ~n1738;
  assign n1740 = n1566 & n1738;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = ~n1736 & ~n1741;
  assign n1743 = ~n1735 & ~n1742;
  assign n1744 = po59  & ~n1743;
  assign n1745 = ~po59  & n1743;
  assign n1746 = ~n1569 & ~n1570;
  assign n1747 = po46  & n1746;
  assign n1748 = ~n1575 & ~n1747;
  assign n1749 = n1575 & n1747;
  assign n1750 = ~n1748 & ~n1749;
  assign n1751 = ~n1745 & ~n1750;
  assign n1752 = ~n1744 & ~n1751;
  assign n1753 = po60  & ~n1752;
  assign n1754 = ~po60  & n1752;
  assign n1755 = ~n1578 & ~n1579;
  assign n1756 = po46  & n1755;
  assign n1757 = ~n1584 & ~n1756;
  assign n1758 = n1584 & n1756;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = ~n1754 & ~n1759;
  assign n1761 = ~n1753 & ~n1760;
  assign n1762 = po61  & ~n1761;
  assign n1763 = ~po61  & n1761;
  assign n1764 = ~n1587 & ~n1588;
  assign n1765 = po46  & n1764;
  assign n1766 = ~n1593 & ~n1765;
  assign n1767 = n1593 & n1765;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = ~n1763 & ~n1768;
  assign n1770 = ~n1762 & ~n1769;
  assign n1771 = po62  & ~n1770;
  assign n1772 = ~po62  & n1770;
  assign n1773 = ~n1596 & ~n1597;
  assign n1774 = po46  & n1773;
  assign n1775 = ~n1602 & ~n1774;
  assign n1776 = n1602 & n1774;
  assign n1777 = ~n1775 & ~n1776;
  assign n1778 = ~n1772 & ~n1777;
  assign n1779 = ~n1771 & ~n1778;
  assign n1780 = n1637 & n1779;
  assign n1781 = ~n1637 & ~n1779;
  assign n1782 = n1615 & po46 ;
  assign n1783 = ~n1614 & ~n1782;
  assign n1784 = n1781 & n1783;
  assign n1785 = ~po63  & ~n1784;
  assign n1786 = ~n1780 & ~n1785;
  assign n1787 = ~n1632 & n1786;
  assign po45  = n1628 | ~n1787;
  assign n1789 = ~n1677 & ~n1678;
  assign n1790 = po45  & n1789;
  assign n1791 = ~n1627 & ~n1790;
  assign n1792 = n1627 & n1790;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = n1637 & ~po45 ;
  assign n1795 = ~n1637 & po45 ;
  assign n1796 = n1779 & ~n1795;
  assign n1797 = po63  & ~n1796;
  assign n1798 = ~n1781 & n1797;
  assign n1799 = ~n1771 & ~n1772;
  assign n1800 = po45  & n1799;
  assign n1801 = ~n1777 & ~n1800;
  assign n1802 = n1777 & n1800;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = pi90  & po45 ;
  assign n1805 = ~pi88  & ~pi89 ;
  assign n1806 = ~pi90  & n1805;
  assign n1807 = ~n1804 & ~n1806;
  assign n1808 = po46  & ~n1807;
  assign n1809 = ~po46  & n1807;
  assign n1810 = ~pi90  & po45 ;
  assign n1811 = pi91  & ~n1810;
  assign n1812 = n1639 & po45 ;
  assign n1813 = ~n1811 & ~n1812;
  assign n1814 = ~n1809 & n1813;
  assign n1815 = ~n1808 & ~n1814;
  assign n1816 = po47  & ~n1815;
  assign n1817 = ~po47  & n1815;
  assign n1818 = po46  & n1787;
  assign n1819 = ~n1812 & ~n1818;
  assign n1820 = pi92  & ~n1819;
  assign n1821 = ~pi92  & n1819;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = ~n1817 & ~n1822;
  assign n1824 = ~n1816 & ~n1823;
  assign n1825 = po48  & ~n1824;
  assign n1826 = ~po48  & n1824;
  assign n1827 = ~n1642 & ~n1643;
  assign n1828 = po45  & n1827;
  assign n1829 = n1647 & ~n1828;
  assign n1830 = ~n1647 & n1828;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = ~n1826 & ~n1831;
  assign n1833 = ~n1825 & ~n1832;
  assign n1834 = po49  & ~n1833;
  assign n1835 = ~po49  & n1833;
  assign n1836 = ~n1650 & ~n1651;
  assign n1837 = po45  & n1836;
  assign n1838 = ~n1656 & ~n1837;
  assign n1839 = n1656 & n1837;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = ~n1835 & ~n1840;
  assign n1842 = ~n1834 & ~n1841;
  assign n1843 = po50  & ~n1842;
  assign n1844 = ~po50  & n1842;
  assign n1845 = ~n1659 & ~n1660;
  assign n1846 = po45  & n1845;
  assign n1847 = n1665 & n1846;
  assign n1848 = ~n1665 & ~n1846;
  assign n1849 = ~n1847 & ~n1848;
  assign n1850 = ~n1844 & ~n1849;
  assign n1851 = ~n1843 & ~n1850;
  assign n1852 = po51  & ~n1851;
  assign n1853 = ~n1668 & ~n1674;
  assign n1854 = po45  & n1853;
  assign n1855 = ~n1673 & ~n1854;
  assign n1856 = n1673 & n1854;
  assign n1857 = ~n1855 & ~n1856;
  assign n1858 = ~po51  & n1851;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = ~n1852 & ~n1859;
  assign n1861 = po52  & ~n1860;
  assign n1862 = ~po52  & n1860;
  assign n1863 = ~n1793 & ~n1862;
  assign n1864 = ~n1861 & ~n1863;
  assign n1865 = po53  & ~n1864;
  assign n1866 = ~po53  & n1864;
  assign n1867 = ~n1681 & ~n1682;
  assign n1868 = po45  & n1867;
  assign n1869 = ~n1687 & ~n1868;
  assign n1870 = n1687 & n1868;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = ~n1866 & ~n1871;
  assign n1873 = ~n1865 & ~n1872;
  assign n1874 = po54  & ~n1873;
  assign n1875 = ~po54  & n1873;
  assign n1876 = ~n1690 & ~n1691;
  assign n1877 = po45  & n1876;
  assign n1878 = ~n1696 & ~n1877;
  assign n1879 = n1696 & n1877;
  assign n1880 = ~n1878 & ~n1879;
  assign n1881 = ~n1875 & ~n1880;
  assign n1882 = ~n1874 & ~n1881;
  assign n1883 = po55  & ~n1882;
  assign n1884 = ~po55  & n1882;
  assign n1885 = ~n1699 & ~n1700;
  assign n1886 = po45  & n1885;
  assign n1887 = ~n1705 & ~n1886;
  assign n1888 = n1705 & n1886;
  assign n1889 = ~n1887 & ~n1888;
  assign n1890 = ~n1884 & ~n1889;
  assign n1891 = ~n1883 & ~n1890;
  assign n1892 = po56  & ~n1891;
  assign n1893 = ~po56  & n1891;
  assign n1894 = ~n1708 & ~n1709;
  assign n1895 = po45  & n1894;
  assign n1896 = ~n1714 & ~n1895;
  assign n1897 = n1714 & n1895;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = ~n1893 & ~n1898;
  assign n1900 = ~n1892 & ~n1899;
  assign n1901 = po57  & ~n1900;
  assign n1902 = ~po57  & n1900;
  assign n1903 = ~n1717 & ~n1718;
  assign n1904 = po45  & n1903;
  assign n1905 = ~n1723 & ~n1904;
  assign n1906 = n1723 & n1904;
  assign n1907 = ~n1905 & ~n1906;
  assign n1908 = ~n1902 & ~n1907;
  assign n1909 = ~n1901 & ~n1908;
  assign n1910 = po58  & ~n1909;
  assign n1911 = ~po58  & n1909;
  assign n1912 = ~n1726 & ~n1727;
  assign n1913 = po45  & n1912;
  assign n1914 = ~n1732 & ~n1913;
  assign n1915 = n1732 & n1913;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = ~n1911 & ~n1916;
  assign n1918 = ~n1910 & ~n1917;
  assign n1919 = po59  & ~n1918;
  assign n1920 = ~po59  & n1918;
  assign n1921 = ~n1735 & ~n1736;
  assign n1922 = po45  & n1921;
  assign n1923 = ~n1741 & ~n1922;
  assign n1924 = n1741 & n1922;
  assign n1925 = ~n1923 & ~n1924;
  assign n1926 = ~n1920 & ~n1925;
  assign n1927 = ~n1919 & ~n1926;
  assign n1928 = po60  & ~n1927;
  assign n1929 = ~po60  & n1927;
  assign n1930 = ~n1744 & ~n1745;
  assign n1931 = po45  & n1930;
  assign n1932 = ~n1750 & ~n1931;
  assign n1933 = n1750 & n1931;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = ~n1929 & ~n1934;
  assign n1936 = ~n1928 & ~n1935;
  assign n1937 = po61  & ~n1936;
  assign n1938 = ~po61  & n1936;
  assign n1939 = ~n1753 & ~n1754;
  assign n1940 = po45  & n1939;
  assign n1941 = ~n1759 & ~n1940;
  assign n1942 = n1759 & n1940;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = ~n1938 & ~n1943;
  assign n1945 = ~n1937 & ~n1944;
  assign n1946 = po62  & ~n1945;
  assign n1947 = ~po62  & n1945;
  assign n1948 = ~n1762 & ~n1763;
  assign n1949 = po45  & n1948;
  assign n1950 = ~n1768 & ~n1949;
  assign n1951 = n1768 & n1949;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = ~n1947 & ~n1952;
  assign n1954 = ~n1946 & ~n1953;
  assign n1955 = n1803 & n1954;
  assign n1956 = ~n1803 & ~n1954;
  assign n1957 = n1781 & po45 ;
  assign n1958 = ~n1780 & ~n1957;
  assign n1959 = n1956 & n1958;
  assign n1960 = ~po63  & ~n1959;
  assign n1961 = ~n1955 & ~n1960;
  assign n1962 = ~n1798 & n1961;
  assign po44  = n1794 | ~n1962;
  assign n1964 = ~n1861 & ~n1862;
  assign n1965 = po44  & n1964;
  assign n1966 = ~n1793 & ~n1965;
  assign n1967 = n1793 & n1965;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = n1803 & ~po44 ;
  assign n1970 = ~n1803 & po44 ;
  assign n1971 = n1954 & ~n1970;
  assign n1972 = po63  & ~n1971;
  assign n1973 = ~n1956 & n1972;
  assign n1974 = ~n1946 & ~n1947;
  assign n1975 = po44  & n1974;
  assign n1976 = ~n1952 & ~n1975;
  assign n1977 = n1952 & n1975;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = pi88  & po44 ;
  assign n1980 = ~pi86  & ~pi87 ;
  assign n1981 = ~pi88  & n1980;
  assign n1982 = ~n1979 & ~n1981;
  assign n1983 = po45  & ~n1982;
  assign n1984 = ~po45  & n1982;
  assign n1985 = ~pi88  & po44 ;
  assign n1986 = pi89  & ~n1985;
  assign n1987 = n1805 & po44 ;
  assign n1988 = ~n1986 & ~n1987;
  assign n1989 = ~n1984 & n1988;
  assign n1990 = ~n1983 & ~n1989;
  assign n1991 = po46  & ~n1990;
  assign n1992 = ~po46  & n1990;
  assign n1993 = po45  & n1962;
  assign n1994 = ~n1987 & ~n1993;
  assign n1995 = pi90  & ~n1994;
  assign n1996 = ~pi90  & n1994;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = ~n1992 & ~n1997;
  assign n1999 = ~n1991 & ~n1998;
  assign n2000 = po47  & ~n1999;
  assign n2001 = ~po47  & n1999;
  assign n2002 = ~n1808 & ~n1809;
  assign n2003 = po44  & n2002;
  assign n2004 = n1813 & ~n2003;
  assign n2005 = ~n1813 & n2003;
  assign n2006 = ~n2004 & ~n2005;
  assign n2007 = ~n2001 & ~n2006;
  assign n2008 = ~n2000 & ~n2007;
  assign n2009 = po48  & ~n2008;
  assign n2010 = ~po48  & n2008;
  assign n2011 = ~n1816 & ~n1817;
  assign n2012 = po44  & n2011;
  assign n2013 = ~n1822 & ~n2012;
  assign n2014 = n1822 & n2012;
  assign n2015 = ~n2013 & ~n2014;
  assign n2016 = ~n2010 & ~n2015;
  assign n2017 = ~n2009 & ~n2016;
  assign n2018 = po49  & ~n2017;
  assign n2019 = ~po49  & n2017;
  assign n2020 = ~n1825 & ~n1826;
  assign n2021 = po44  & n2020;
  assign n2022 = n1831 & n2021;
  assign n2023 = ~n1831 & ~n2021;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = ~n2019 & ~n2024;
  assign n2026 = ~n2018 & ~n2025;
  assign n2027 = po50  & ~n2026;
  assign n2028 = ~po50  & n2026;
  assign n2029 = ~n1834 & ~n1835;
  assign n2030 = po44  & n2029;
  assign n2031 = ~n1840 & ~n2030;
  assign n2032 = n1840 & n2030;
  assign n2033 = ~n2031 & ~n2032;
  assign n2034 = ~n2028 & ~n2033;
  assign n2035 = ~n2027 & ~n2034;
  assign n2036 = po51  & ~n2035;
  assign n2037 = ~po51  & n2035;
  assign n2038 = ~n1843 & ~n1844;
  assign n2039 = po44  & n2038;
  assign n2040 = ~n1849 & ~n2039;
  assign n2041 = n1849 & n2039;
  assign n2042 = ~n2040 & ~n2041;
  assign n2043 = ~n2037 & ~n2042;
  assign n2044 = ~n2036 & ~n2043;
  assign n2045 = po52  & ~n2044;
  assign n2046 = ~n1852 & ~n1858;
  assign n2047 = po44  & n2046;
  assign n2048 = ~n1857 & ~n2047;
  assign n2049 = n1857 & n2047;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = ~po52  & n2044;
  assign n2052 = ~n2050 & ~n2051;
  assign n2053 = ~n2045 & ~n2052;
  assign n2054 = po53  & ~n2053;
  assign n2055 = ~po53  & n2053;
  assign n2056 = ~n1968 & ~n2055;
  assign n2057 = ~n2054 & ~n2056;
  assign n2058 = po54  & ~n2057;
  assign n2059 = ~po54  & n2057;
  assign n2060 = ~n1865 & ~n1866;
  assign n2061 = po44  & n2060;
  assign n2062 = ~n1871 & ~n2061;
  assign n2063 = n1871 & n2061;
  assign n2064 = ~n2062 & ~n2063;
  assign n2065 = ~n2059 & ~n2064;
  assign n2066 = ~n2058 & ~n2065;
  assign n2067 = po55  & ~n2066;
  assign n2068 = ~po55  & n2066;
  assign n2069 = ~n1874 & ~n1875;
  assign n2070 = po44  & n2069;
  assign n2071 = ~n1880 & ~n2070;
  assign n2072 = n1880 & n2070;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = ~n2068 & ~n2073;
  assign n2075 = ~n2067 & ~n2074;
  assign n2076 = po56  & ~n2075;
  assign n2077 = ~po56  & n2075;
  assign n2078 = ~n1883 & ~n1884;
  assign n2079 = po44  & n2078;
  assign n2080 = ~n1889 & ~n2079;
  assign n2081 = n1889 & n2079;
  assign n2082 = ~n2080 & ~n2081;
  assign n2083 = ~n2077 & ~n2082;
  assign n2084 = ~n2076 & ~n2083;
  assign n2085 = po57  & ~n2084;
  assign n2086 = ~po57  & n2084;
  assign n2087 = ~n1892 & ~n1893;
  assign n2088 = po44  & n2087;
  assign n2089 = ~n1898 & ~n2088;
  assign n2090 = n1898 & n2088;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = ~n2086 & ~n2091;
  assign n2093 = ~n2085 & ~n2092;
  assign n2094 = po58  & ~n2093;
  assign n2095 = ~po58  & n2093;
  assign n2096 = ~n1901 & ~n1902;
  assign n2097 = po44  & n2096;
  assign n2098 = ~n1907 & ~n2097;
  assign n2099 = n1907 & n2097;
  assign n2100 = ~n2098 & ~n2099;
  assign n2101 = ~n2095 & ~n2100;
  assign n2102 = ~n2094 & ~n2101;
  assign n2103 = po59  & ~n2102;
  assign n2104 = ~po59  & n2102;
  assign n2105 = ~n1910 & ~n1911;
  assign n2106 = po44  & n2105;
  assign n2107 = ~n1916 & ~n2106;
  assign n2108 = n1916 & n2106;
  assign n2109 = ~n2107 & ~n2108;
  assign n2110 = ~n2104 & ~n2109;
  assign n2111 = ~n2103 & ~n2110;
  assign n2112 = po60  & ~n2111;
  assign n2113 = ~po60  & n2111;
  assign n2114 = ~n1919 & ~n1920;
  assign n2115 = po44  & n2114;
  assign n2116 = ~n1925 & ~n2115;
  assign n2117 = n1925 & n2115;
  assign n2118 = ~n2116 & ~n2117;
  assign n2119 = ~n2113 & ~n2118;
  assign n2120 = ~n2112 & ~n2119;
  assign n2121 = po61  & ~n2120;
  assign n2122 = ~po61  & n2120;
  assign n2123 = ~n1928 & ~n1929;
  assign n2124 = po44  & n2123;
  assign n2125 = ~n1934 & ~n2124;
  assign n2126 = n1934 & n2124;
  assign n2127 = ~n2125 & ~n2126;
  assign n2128 = ~n2122 & ~n2127;
  assign n2129 = ~n2121 & ~n2128;
  assign n2130 = po62  & ~n2129;
  assign n2131 = ~po62  & n2129;
  assign n2132 = ~n1937 & ~n1938;
  assign n2133 = po44  & n2132;
  assign n2134 = ~n1943 & ~n2133;
  assign n2135 = n1943 & n2133;
  assign n2136 = ~n2134 & ~n2135;
  assign n2137 = ~n2131 & ~n2136;
  assign n2138 = ~n2130 & ~n2137;
  assign n2139 = n1978 & n2138;
  assign n2140 = ~n1978 & ~n2138;
  assign n2141 = n1956 & po44 ;
  assign n2142 = ~n1955 & ~n2141;
  assign n2143 = n2140 & n2142;
  assign n2144 = ~po63  & ~n2143;
  assign n2145 = ~n2139 & ~n2144;
  assign n2146 = ~n1973 & n2145;
  assign po43  = n1969 | ~n2146;
  assign n2148 = ~n2054 & ~n2055;
  assign n2149 = po43  & n2148;
  assign n2150 = ~n1968 & ~n2149;
  assign n2151 = n1968 & n2149;
  assign n2152 = ~n2150 & ~n2151;
  assign n2153 = n1978 & ~po43 ;
  assign n2154 = ~n1978 & po43 ;
  assign n2155 = n2138 & ~n2154;
  assign n2156 = po63  & ~n2155;
  assign n2157 = ~n2140 & n2156;
  assign n2158 = ~n2130 & ~n2131;
  assign n2159 = po43  & n2158;
  assign n2160 = ~n2136 & ~n2159;
  assign n2161 = n2136 & n2159;
  assign n2162 = ~n2160 & ~n2161;
  assign n2163 = pi86  & po43 ;
  assign n2164 = ~pi84  & ~pi85 ;
  assign n2165 = ~pi86  & n2164;
  assign n2166 = ~n2163 & ~n2165;
  assign n2167 = po44  & ~n2166;
  assign n2168 = ~po44  & n2166;
  assign n2169 = ~pi86  & po43 ;
  assign n2170 = pi87  & ~n2169;
  assign n2171 = n1980 & po43 ;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = ~n2168 & n2172;
  assign n2174 = ~n2167 & ~n2173;
  assign n2175 = po45  & ~n2174;
  assign n2176 = ~po45  & n2174;
  assign n2177 = po44  & n2146;
  assign n2178 = ~n2171 & ~n2177;
  assign n2179 = pi88  & ~n2178;
  assign n2180 = ~pi88  & n2178;
  assign n2181 = ~n2179 & ~n2180;
  assign n2182 = ~n2176 & ~n2181;
  assign n2183 = ~n2175 & ~n2182;
  assign n2184 = po46  & ~n2183;
  assign n2185 = ~po46  & n2183;
  assign n2186 = ~n1983 & ~n1984;
  assign n2187 = po43  & n2186;
  assign n2188 = n1988 & ~n2187;
  assign n2189 = ~n1988 & n2187;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = ~n2185 & ~n2190;
  assign n2192 = ~n2184 & ~n2191;
  assign n2193 = po47  & ~n2192;
  assign n2194 = ~po47  & n2192;
  assign n2195 = ~n1991 & ~n1992;
  assign n2196 = po43  & n2195;
  assign n2197 = ~n1997 & ~n2196;
  assign n2198 = n1997 & n2196;
  assign n2199 = ~n2197 & ~n2198;
  assign n2200 = ~n2194 & ~n2199;
  assign n2201 = ~n2193 & ~n2200;
  assign n2202 = po48  & ~n2201;
  assign n2203 = ~po48  & n2201;
  assign n2204 = ~n2000 & ~n2001;
  assign n2205 = po43  & n2204;
  assign n2206 = n2006 & n2205;
  assign n2207 = ~n2006 & ~n2205;
  assign n2208 = ~n2206 & ~n2207;
  assign n2209 = ~n2203 & ~n2208;
  assign n2210 = ~n2202 & ~n2209;
  assign n2211 = po49  & ~n2210;
  assign n2212 = ~po49  & n2210;
  assign n2213 = ~n2009 & ~n2010;
  assign n2214 = po43  & n2213;
  assign n2215 = ~n2015 & ~n2214;
  assign n2216 = n2015 & n2214;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~n2212 & ~n2217;
  assign n2219 = ~n2211 & ~n2218;
  assign n2220 = po50  & ~n2219;
  assign n2221 = ~po50  & n2219;
  assign n2222 = ~n2018 & ~n2019;
  assign n2223 = po43  & n2222;
  assign n2224 = ~n2024 & ~n2223;
  assign n2225 = n2024 & n2223;
  assign n2226 = ~n2224 & ~n2225;
  assign n2227 = ~n2221 & ~n2226;
  assign n2228 = ~n2220 & ~n2227;
  assign n2229 = po51  & ~n2228;
  assign n2230 = ~po51  & n2228;
  assign n2231 = ~n2027 & ~n2028;
  assign n2232 = po43  & n2231;
  assign n2233 = ~n2033 & ~n2232;
  assign n2234 = n2033 & n2232;
  assign n2235 = ~n2233 & ~n2234;
  assign n2236 = ~n2230 & ~n2235;
  assign n2237 = ~n2229 & ~n2236;
  assign n2238 = po52  & ~n2237;
  assign n2239 = ~po52  & n2237;
  assign n2240 = ~n2036 & ~n2037;
  assign n2241 = po43  & n2240;
  assign n2242 = ~n2042 & ~n2241;
  assign n2243 = n2042 & n2241;
  assign n2244 = ~n2242 & ~n2243;
  assign n2245 = ~n2239 & ~n2244;
  assign n2246 = ~n2238 & ~n2245;
  assign n2247 = po53  & ~n2246;
  assign n2248 = ~n2045 & ~n2051;
  assign n2249 = po43  & n2248;
  assign n2250 = ~n2050 & ~n2249;
  assign n2251 = n2050 & n2249;
  assign n2252 = ~n2250 & ~n2251;
  assign n2253 = ~po53  & n2246;
  assign n2254 = ~n2252 & ~n2253;
  assign n2255 = ~n2247 & ~n2254;
  assign n2256 = po54  & ~n2255;
  assign n2257 = ~po54  & n2255;
  assign n2258 = ~n2152 & ~n2257;
  assign n2259 = ~n2256 & ~n2258;
  assign n2260 = po55  & ~n2259;
  assign n2261 = ~po55  & n2259;
  assign n2262 = ~n2058 & ~n2059;
  assign n2263 = po43  & n2262;
  assign n2264 = ~n2064 & ~n2263;
  assign n2265 = n2064 & n2263;
  assign n2266 = ~n2264 & ~n2265;
  assign n2267 = ~n2261 & ~n2266;
  assign n2268 = ~n2260 & ~n2267;
  assign n2269 = po56  & ~n2268;
  assign n2270 = ~po56  & n2268;
  assign n2271 = ~n2067 & ~n2068;
  assign n2272 = po43  & n2271;
  assign n2273 = ~n2073 & ~n2272;
  assign n2274 = n2073 & n2272;
  assign n2275 = ~n2273 & ~n2274;
  assign n2276 = ~n2270 & ~n2275;
  assign n2277 = ~n2269 & ~n2276;
  assign n2278 = po57  & ~n2277;
  assign n2279 = ~po57  & n2277;
  assign n2280 = ~n2076 & ~n2077;
  assign n2281 = po43  & n2280;
  assign n2282 = ~n2082 & ~n2281;
  assign n2283 = n2082 & n2281;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = ~n2279 & ~n2284;
  assign n2286 = ~n2278 & ~n2285;
  assign n2287 = po58  & ~n2286;
  assign n2288 = ~po58  & n2286;
  assign n2289 = ~n2085 & ~n2086;
  assign n2290 = po43  & n2289;
  assign n2291 = ~n2091 & ~n2290;
  assign n2292 = n2091 & n2290;
  assign n2293 = ~n2291 & ~n2292;
  assign n2294 = ~n2288 & ~n2293;
  assign n2295 = ~n2287 & ~n2294;
  assign n2296 = po59  & ~n2295;
  assign n2297 = ~po59  & n2295;
  assign n2298 = ~n2094 & ~n2095;
  assign n2299 = po43  & n2298;
  assign n2300 = ~n2100 & ~n2299;
  assign n2301 = n2100 & n2299;
  assign n2302 = ~n2300 & ~n2301;
  assign n2303 = ~n2297 & ~n2302;
  assign n2304 = ~n2296 & ~n2303;
  assign n2305 = po60  & ~n2304;
  assign n2306 = ~po60  & n2304;
  assign n2307 = ~n2103 & ~n2104;
  assign n2308 = po43  & n2307;
  assign n2309 = ~n2109 & ~n2308;
  assign n2310 = n2109 & n2308;
  assign n2311 = ~n2309 & ~n2310;
  assign n2312 = ~n2306 & ~n2311;
  assign n2313 = ~n2305 & ~n2312;
  assign n2314 = po61  & ~n2313;
  assign n2315 = ~po61  & n2313;
  assign n2316 = ~n2112 & ~n2113;
  assign n2317 = po43  & n2316;
  assign n2318 = ~n2118 & ~n2317;
  assign n2319 = n2118 & n2317;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = ~n2315 & ~n2320;
  assign n2322 = ~n2314 & ~n2321;
  assign n2323 = po62  & ~n2322;
  assign n2324 = ~po62  & n2322;
  assign n2325 = ~n2121 & ~n2122;
  assign n2326 = po43  & n2325;
  assign n2327 = ~n2127 & ~n2326;
  assign n2328 = n2127 & n2326;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = ~n2324 & ~n2329;
  assign n2331 = ~n2323 & ~n2330;
  assign n2332 = n2162 & n2331;
  assign n2333 = ~n2162 & ~n2331;
  assign n2334 = n2140 & po43 ;
  assign n2335 = ~n2139 & ~n2334;
  assign n2336 = n2333 & n2335;
  assign n2337 = ~po63  & ~n2336;
  assign n2338 = ~n2332 & ~n2337;
  assign n2339 = ~n2157 & n2338;
  assign po42  = n2153 | ~n2339;
  assign n2341 = ~n2256 & ~n2257;
  assign n2342 = po42  & n2341;
  assign n2343 = ~n2152 & ~n2342;
  assign n2344 = n2152 & n2342;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = n2162 & ~po42 ;
  assign n2347 = ~n2162 & po42 ;
  assign n2348 = n2331 & ~n2347;
  assign n2349 = po63  & ~n2348;
  assign n2350 = ~n2333 & n2349;
  assign n2351 = ~n2323 & ~n2324;
  assign n2352 = po42  & n2351;
  assign n2353 = ~n2329 & ~n2352;
  assign n2354 = n2329 & n2352;
  assign n2355 = ~n2353 & ~n2354;
  assign n2356 = pi84  & po42 ;
  assign n2357 = ~pi82  & ~pi83 ;
  assign n2358 = ~pi84  & n2357;
  assign n2359 = ~n2356 & ~n2358;
  assign n2360 = po43  & ~n2359;
  assign n2361 = ~po43  & n2359;
  assign n2362 = ~pi84  & po42 ;
  assign n2363 = pi85  & ~n2362;
  assign n2364 = n2164 & po42 ;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = ~n2361 & n2365;
  assign n2367 = ~n2360 & ~n2366;
  assign n2368 = po44  & ~n2367;
  assign n2369 = ~po44  & n2367;
  assign n2370 = po43  & n2339;
  assign n2371 = ~n2364 & ~n2370;
  assign n2372 = pi86  & ~n2371;
  assign n2373 = ~pi86  & n2371;
  assign n2374 = ~n2372 & ~n2373;
  assign n2375 = ~n2369 & ~n2374;
  assign n2376 = ~n2368 & ~n2375;
  assign n2377 = po45  & ~n2376;
  assign n2378 = ~po45  & n2376;
  assign n2379 = ~n2167 & ~n2168;
  assign n2380 = po42  & n2379;
  assign n2381 = n2172 & ~n2380;
  assign n2382 = ~n2172 & n2380;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = ~n2378 & ~n2383;
  assign n2385 = ~n2377 & ~n2384;
  assign n2386 = po46  & ~n2385;
  assign n2387 = ~po46  & n2385;
  assign n2388 = ~n2175 & ~n2176;
  assign n2389 = po42  & n2388;
  assign n2390 = ~n2181 & ~n2389;
  assign n2391 = n2181 & n2389;
  assign n2392 = ~n2390 & ~n2391;
  assign n2393 = ~n2387 & ~n2392;
  assign n2394 = ~n2386 & ~n2393;
  assign n2395 = po47  & ~n2394;
  assign n2396 = ~po47  & n2394;
  assign n2397 = ~n2184 & ~n2185;
  assign n2398 = po42  & n2397;
  assign n2399 = n2190 & n2398;
  assign n2400 = ~n2190 & ~n2398;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = ~n2396 & ~n2401;
  assign n2403 = ~n2395 & ~n2402;
  assign n2404 = po48  & ~n2403;
  assign n2405 = ~po48  & n2403;
  assign n2406 = ~n2193 & ~n2194;
  assign n2407 = po42  & n2406;
  assign n2408 = ~n2199 & ~n2407;
  assign n2409 = n2199 & n2407;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = ~n2405 & ~n2410;
  assign n2412 = ~n2404 & ~n2411;
  assign n2413 = po49  & ~n2412;
  assign n2414 = ~po49  & n2412;
  assign n2415 = ~n2202 & ~n2203;
  assign n2416 = po42  & n2415;
  assign n2417 = ~n2208 & ~n2416;
  assign n2418 = n2208 & n2416;
  assign n2419 = ~n2417 & ~n2418;
  assign n2420 = ~n2414 & ~n2419;
  assign n2421 = ~n2413 & ~n2420;
  assign n2422 = po50  & ~n2421;
  assign n2423 = ~po50  & n2421;
  assign n2424 = ~n2211 & ~n2212;
  assign n2425 = po42  & n2424;
  assign n2426 = ~n2217 & ~n2425;
  assign n2427 = n2217 & n2425;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = ~n2423 & ~n2428;
  assign n2430 = ~n2422 & ~n2429;
  assign n2431 = po51  & ~n2430;
  assign n2432 = ~po51  & n2430;
  assign n2433 = ~n2220 & ~n2221;
  assign n2434 = po42  & n2433;
  assign n2435 = ~n2226 & ~n2434;
  assign n2436 = n2226 & n2434;
  assign n2437 = ~n2435 & ~n2436;
  assign n2438 = ~n2432 & ~n2437;
  assign n2439 = ~n2431 & ~n2438;
  assign n2440 = po52  & ~n2439;
  assign n2441 = ~po52  & n2439;
  assign n2442 = ~n2229 & ~n2230;
  assign n2443 = po42  & n2442;
  assign n2444 = ~n2235 & ~n2443;
  assign n2445 = n2235 & n2443;
  assign n2446 = ~n2444 & ~n2445;
  assign n2447 = ~n2441 & ~n2446;
  assign n2448 = ~n2440 & ~n2447;
  assign n2449 = po53  & ~n2448;
  assign n2450 = ~po53  & n2448;
  assign n2451 = ~n2238 & ~n2239;
  assign n2452 = po42  & n2451;
  assign n2453 = ~n2244 & ~n2452;
  assign n2454 = n2244 & n2452;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = ~n2450 & ~n2455;
  assign n2457 = ~n2449 & ~n2456;
  assign n2458 = po54  & ~n2457;
  assign n2459 = ~n2247 & ~n2253;
  assign n2460 = po42  & n2459;
  assign n2461 = ~n2252 & ~n2460;
  assign n2462 = n2252 & n2460;
  assign n2463 = ~n2461 & ~n2462;
  assign n2464 = ~po54  & n2457;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = ~n2458 & ~n2465;
  assign n2467 = po55  & ~n2466;
  assign n2468 = ~po55  & n2466;
  assign n2469 = ~n2345 & ~n2468;
  assign n2470 = ~n2467 & ~n2469;
  assign n2471 = po56  & ~n2470;
  assign n2472 = ~po56  & n2470;
  assign n2473 = ~n2260 & ~n2261;
  assign n2474 = po42  & n2473;
  assign n2475 = ~n2266 & ~n2474;
  assign n2476 = n2266 & n2474;
  assign n2477 = ~n2475 & ~n2476;
  assign n2478 = ~n2472 & ~n2477;
  assign n2479 = ~n2471 & ~n2478;
  assign n2480 = po57  & ~n2479;
  assign n2481 = ~po57  & n2479;
  assign n2482 = ~n2269 & ~n2270;
  assign n2483 = po42  & n2482;
  assign n2484 = ~n2275 & ~n2483;
  assign n2485 = n2275 & n2483;
  assign n2486 = ~n2484 & ~n2485;
  assign n2487 = ~n2481 & ~n2486;
  assign n2488 = ~n2480 & ~n2487;
  assign n2489 = po58  & ~n2488;
  assign n2490 = ~po58  & n2488;
  assign n2491 = ~n2278 & ~n2279;
  assign n2492 = po42  & n2491;
  assign n2493 = ~n2284 & ~n2492;
  assign n2494 = n2284 & n2492;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = ~n2490 & ~n2495;
  assign n2497 = ~n2489 & ~n2496;
  assign n2498 = po59  & ~n2497;
  assign n2499 = ~po59  & n2497;
  assign n2500 = ~n2287 & ~n2288;
  assign n2501 = po42  & n2500;
  assign n2502 = ~n2293 & ~n2501;
  assign n2503 = n2293 & n2501;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = ~n2499 & ~n2504;
  assign n2506 = ~n2498 & ~n2505;
  assign n2507 = po60  & ~n2506;
  assign n2508 = ~po60  & n2506;
  assign n2509 = ~n2296 & ~n2297;
  assign n2510 = po42  & n2509;
  assign n2511 = ~n2302 & ~n2510;
  assign n2512 = n2302 & n2510;
  assign n2513 = ~n2511 & ~n2512;
  assign n2514 = ~n2508 & ~n2513;
  assign n2515 = ~n2507 & ~n2514;
  assign n2516 = po61  & ~n2515;
  assign n2517 = ~po61  & n2515;
  assign n2518 = ~n2305 & ~n2306;
  assign n2519 = po42  & n2518;
  assign n2520 = ~n2311 & ~n2519;
  assign n2521 = n2311 & n2519;
  assign n2522 = ~n2520 & ~n2521;
  assign n2523 = ~n2517 & ~n2522;
  assign n2524 = ~n2516 & ~n2523;
  assign n2525 = po62  & ~n2524;
  assign n2526 = ~po62  & n2524;
  assign n2527 = ~n2314 & ~n2315;
  assign n2528 = po42  & n2527;
  assign n2529 = ~n2320 & ~n2528;
  assign n2530 = n2320 & n2528;
  assign n2531 = ~n2529 & ~n2530;
  assign n2532 = ~n2526 & ~n2531;
  assign n2533 = ~n2525 & ~n2532;
  assign n2534 = n2355 & n2533;
  assign n2535 = ~n2355 & ~n2533;
  assign n2536 = n2333 & po42 ;
  assign n2537 = ~n2332 & ~n2536;
  assign n2538 = n2535 & n2537;
  assign n2539 = ~po63  & ~n2538;
  assign n2540 = ~n2534 & ~n2539;
  assign n2541 = ~n2350 & n2540;
  assign po41  = n2346 | ~n2541;
  assign n2543 = ~n2467 & ~n2468;
  assign n2544 = po41  & n2543;
  assign n2545 = ~n2345 & ~n2544;
  assign n2546 = n2345 & n2544;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = n2355 & ~po41 ;
  assign n2549 = ~n2355 & po41 ;
  assign n2550 = n2533 & ~n2549;
  assign n2551 = po63  & ~n2550;
  assign n2552 = ~n2535 & n2551;
  assign n2553 = ~n2525 & ~n2526;
  assign n2554 = po41  & n2553;
  assign n2555 = ~n2531 & ~n2554;
  assign n2556 = n2531 & n2554;
  assign n2557 = ~n2555 & ~n2556;
  assign n2558 = pi82  & po41 ;
  assign n2559 = ~pi80  & ~pi81 ;
  assign n2560 = ~pi82  & n2559;
  assign n2561 = ~n2558 & ~n2560;
  assign n2562 = po42  & ~n2561;
  assign n2563 = ~po42  & n2561;
  assign n2564 = ~pi82  & po41 ;
  assign n2565 = pi83  & ~n2564;
  assign n2566 = n2357 & po41 ;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = ~n2563 & n2567;
  assign n2569 = ~n2562 & ~n2568;
  assign n2570 = po43  & ~n2569;
  assign n2571 = ~po43  & n2569;
  assign n2572 = po42  & n2541;
  assign n2573 = ~n2566 & ~n2572;
  assign n2574 = pi84  & ~n2573;
  assign n2575 = ~pi84  & n2573;
  assign n2576 = ~n2574 & ~n2575;
  assign n2577 = ~n2571 & ~n2576;
  assign n2578 = ~n2570 & ~n2577;
  assign n2579 = po44  & ~n2578;
  assign n2580 = ~po44  & n2578;
  assign n2581 = ~n2360 & ~n2361;
  assign n2582 = po41  & n2581;
  assign n2583 = n2365 & ~n2582;
  assign n2584 = ~n2365 & n2582;
  assign n2585 = ~n2583 & ~n2584;
  assign n2586 = ~n2580 & ~n2585;
  assign n2587 = ~n2579 & ~n2586;
  assign n2588 = po45  & ~n2587;
  assign n2589 = ~po45  & n2587;
  assign n2590 = ~n2368 & ~n2369;
  assign n2591 = po41  & n2590;
  assign n2592 = ~n2374 & ~n2591;
  assign n2593 = n2374 & n2591;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = ~n2589 & ~n2594;
  assign n2596 = ~n2588 & ~n2595;
  assign n2597 = po46  & ~n2596;
  assign n2598 = ~po46  & n2596;
  assign n2599 = ~n2377 & ~n2378;
  assign n2600 = po41  & n2599;
  assign n2601 = n2383 & n2600;
  assign n2602 = ~n2383 & ~n2600;
  assign n2603 = ~n2601 & ~n2602;
  assign n2604 = ~n2598 & ~n2603;
  assign n2605 = ~n2597 & ~n2604;
  assign n2606 = po47  & ~n2605;
  assign n2607 = ~po47  & n2605;
  assign n2608 = ~n2386 & ~n2387;
  assign n2609 = po41  & n2608;
  assign n2610 = ~n2392 & ~n2609;
  assign n2611 = n2392 & n2609;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = ~n2607 & ~n2612;
  assign n2614 = ~n2606 & ~n2613;
  assign n2615 = po48  & ~n2614;
  assign n2616 = ~po48  & n2614;
  assign n2617 = ~n2395 & ~n2396;
  assign n2618 = po41  & n2617;
  assign n2619 = ~n2401 & ~n2618;
  assign n2620 = n2401 & n2618;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = ~n2616 & ~n2621;
  assign n2623 = ~n2615 & ~n2622;
  assign n2624 = po49  & ~n2623;
  assign n2625 = ~po49  & n2623;
  assign n2626 = ~n2404 & ~n2405;
  assign n2627 = po41  & n2626;
  assign n2628 = ~n2410 & ~n2627;
  assign n2629 = n2410 & n2627;
  assign n2630 = ~n2628 & ~n2629;
  assign n2631 = ~n2625 & ~n2630;
  assign n2632 = ~n2624 & ~n2631;
  assign n2633 = po50  & ~n2632;
  assign n2634 = ~po50  & n2632;
  assign n2635 = ~n2413 & ~n2414;
  assign n2636 = po41  & n2635;
  assign n2637 = ~n2419 & ~n2636;
  assign n2638 = n2419 & n2636;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = ~n2634 & ~n2639;
  assign n2641 = ~n2633 & ~n2640;
  assign n2642 = po51  & ~n2641;
  assign n2643 = ~po51  & n2641;
  assign n2644 = ~n2422 & ~n2423;
  assign n2645 = po41  & n2644;
  assign n2646 = ~n2428 & ~n2645;
  assign n2647 = n2428 & n2645;
  assign n2648 = ~n2646 & ~n2647;
  assign n2649 = ~n2643 & ~n2648;
  assign n2650 = ~n2642 & ~n2649;
  assign n2651 = po52  & ~n2650;
  assign n2652 = ~po52  & n2650;
  assign n2653 = ~n2431 & ~n2432;
  assign n2654 = po41  & n2653;
  assign n2655 = ~n2437 & ~n2654;
  assign n2656 = n2437 & n2654;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = ~n2652 & ~n2657;
  assign n2659 = ~n2651 & ~n2658;
  assign n2660 = po53  & ~n2659;
  assign n2661 = ~po53  & n2659;
  assign n2662 = ~n2440 & ~n2441;
  assign n2663 = po41  & n2662;
  assign n2664 = ~n2446 & ~n2663;
  assign n2665 = n2446 & n2663;
  assign n2666 = ~n2664 & ~n2665;
  assign n2667 = ~n2661 & ~n2666;
  assign n2668 = ~n2660 & ~n2667;
  assign n2669 = po54  & ~n2668;
  assign n2670 = ~po54  & n2668;
  assign n2671 = ~n2449 & ~n2450;
  assign n2672 = po41  & n2671;
  assign n2673 = ~n2455 & ~n2672;
  assign n2674 = n2455 & n2672;
  assign n2675 = ~n2673 & ~n2674;
  assign n2676 = ~n2670 & ~n2675;
  assign n2677 = ~n2669 & ~n2676;
  assign n2678 = po55  & ~n2677;
  assign n2679 = ~n2458 & ~n2464;
  assign n2680 = po41  & n2679;
  assign n2681 = ~n2463 & ~n2680;
  assign n2682 = n2463 & n2680;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = ~po55  & n2677;
  assign n2685 = ~n2683 & ~n2684;
  assign n2686 = ~n2678 & ~n2685;
  assign n2687 = po56  & ~n2686;
  assign n2688 = ~po56  & n2686;
  assign n2689 = ~n2547 & ~n2688;
  assign n2690 = ~n2687 & ~n2689;
  assign n2691 = po57  & ~n2690;
  assign n2692 = ~po57  & n2690;
  assign n2693 = ~n2471 & ~n2472;
  assign n2694 = po41  & n2693;
  assign n2695 = ~n2477 & ~n2694;
  assign n2696 = n2477 & n2694;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = ~n2692 & ~n2697;
  assign n2699 = ~n2691 & ~n2698;
  assign n2700 = po58  & ~n2699;
  assign n2701 = ~po58  & n2699;
  assign n2702 = ~n2480 & ~n2481;
  assign n2703 = po41  & n2702;
  assign n2704 = ~n2486 & ~n2703;
  assign n2705 = n2486 & n2703;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = ~n2701 & ~n2706;
  assign n2708 = ~n2700 & ~n2707;
  assign n2709 = po59  & ~n2708;
  assign n2710 = ~po59  & n2708;
  assign n2711 = ~n2489 & ~n2490;
  assign n2712 = po41  & n2711;
  assign n2713 = ~n2495 & ~n2712;
  assign n2714 = n2495 & n2712;
  assign n2715 = ~n2713 & ~n2714;
  assign n2716 = ~n2710 & ~n2715;
  assign n2717 = ~n2709 & ~n2716;
  assign n2718 = po60  & ~n2717;
  assign n2719 = ~po60  & n2717;
  assign n2720 = ~n2498 & ~n2499;
  assign n2721 = po41  & n2720;
  assign n2722 = ~n2504 & ~n2721;
  assign n2723 = n2504 & n2721;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = ~n2719 & ~n2724;
  assign n2726 = ~n2718 & ~n2725;
  assign n2727 = po61  & ~n2726;
  assign n2728 = ~po61  & n2726;
  assign n2729 = ~n2507 & ~n2508;
  assign n2730 = po41  & n2729;
  assign n2731 = ~n2513 & ~n2730;
  assign n2732 = n2513 & n2730;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = ~n2728 & ~n2733;
  assign n2735 = ~n2727 & ~n2734;
  assign n2736 = po62  & ~n2735;
  assign n2737 = ~po62  & n2735;
  assign n2738 = ~n2516 & ~n2517;
  assign n2739 = po41  & n2738;
  assign n2740 = ~n2522 & ~n2739;
  assign n2741 = n2522 & n2739;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = ~n2737 & ~n2742;
  assign n2744 = ~n2736 & ~n2743;
  assign n2745 = n2557 & n2744;
  assign n2746 = ~n2557 & ~n2744;
  assign n2747 = n2535 & po41 ;
  assign n2748 = ~n2534 & ~n2747;
  assign n2749 = n2746 & n2748;
  assign n2750 = ~po63  & ~n2749;
  assign n2751 = ~n2745 & ~n2750;
  assign n2752 = ~n2552 & n2751;
  assign po40  = n2548 | ~n2752;
  assign n2754 = ~n2687 & ~n2688;
  assign n2755 = po40  & n2754;
  assign n2756 = ~n2547 & ~n2755;
  assign n2757 = n2547 & n2755;
  assign n2758 = ~n2756 & ~n2757;
  assign n2759 = n2557 & ~po40 ;
  assign n2760 = ~n2557 & po40 ;
  assign n2761 = n2744 & ~n2760;
  assign n2762 = po63  & ~n2761;
  assign n2763 = ~n2746 & n2762;
  assign n2764 = ~n2736 & ~n2737;
  assign n2765 = po40  & n2764;
  assign n2766 = ~n2742 & ~n2765;
  assign n2767 = n2742 & n2765;
  assign n2768 = ~n2766 & ~n2767;
  assign n2769 = pi80  & po40 ;
  assign n2770 = ~pi78  & ~pi79 ;
  assign n2771 = ~pi80  & n2770;
  assign n2772 = ~n2769 & ~n2771;
  assign n2773 = po41  & ~n2772;
  assign n2774 = ~po41  & n2772;
  assign n2775 = ~pi80  & po40 ;
  assign n2776 = pi81  & ~n2775;
  assign n2777 = n2559 & po40 ;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = ~n2774 & n2778;
  assign n2780 = ~n2773 & ~n2779;
  assign n2781 = po42  & ~n2780;
  assign n2782 = ~po42  & n2780;
  assign n2783 = po41  & n2752;
  assign n2784 = ~n2777 & ~n2783;
  assign n2785 = pi82  & ~n2784;
  assign n2786 = ~pi82  & n2784;
  assign n2787 = ~n2785 & ~n2786;
  assign n2788 = ~n2782 & ~n2787;
  assign n2789 = ~n2781 & ~n2788;
  assign n2790 = po43  & ~n2789;
  assign n2791 = ~po43  & n2789;
  assign n2792 = ~n2562 & ~n2563;
  assign n2793 = po40  & n2792;
  assign n2794 = n2567 & ~n2793;
  assign n2795 = ~n2567 & n2793;
  assign n2796 = ~n2794 & ~n2795;
  assign n2797 = ~n2791 & ~n2796;
  assign n2798 = ~n2790 & ~n2797;
  assign n2799 = po44  & ~n2798;
  assign n2800 = ~po44  & n2798;
  assign n2801 = ~n2570 & ~n2571;
  assign n2802 = po40  & n2801;
  assign n2803 = ~n2576 & ~n2802;
  assign n2804 = n2576 & n2802;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = ~n2800 & ~n2805;
  assign n2807 = ~n2799 & ~n2806;
  assign n2808 = po45  & ~n2807;
  assign n2809 = ~po45  & n2807;
  assign n2810 = ~n2579 & ~n2580;
  assign n2811 = po40  & n2810;
  assign n2812 = n2585 & n2811;
  assign n2813 = ~n2585 & ~n2811;
  assign n2814 = ~n2812 & ~n2813;
  assign n2815 = ~n2809 & ~n2814;
  assign n2816 = ~n2808 & ~n2815;
  assign n2817 = po46  & ~n2816;
  assign n2818 = ~po46  & n2816;
  assign n2819 = ~n2588 & ~n2589;
  assign n2820 = po40  & n2819;
  assign n2821 = ~n2594 & ~n2820;
  assign n2822 = n2594 & n2820;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = ~n2818 & ~n2823;
  assign n2825 = ~n2817 & ~n2824;
  assign n2826 = po47  & ~n2825;
  assign n2827 = ~po47  & n2825;
  assign n2828 = ~n2597 & ~n2598;
  assign n2829 = po40  & n2828;
  assign n2830 = ~n2603 & ~n2829;
  assign n2831 = n2603 & n2829;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = ~n2827 & ~n2832;
  assign n2834 = ~n2826 & ~n2833;
  assign n2835 = po48  & ~n2834;
  assign n2836 = ~po48  & n2834;
  assign n2837 = ~n2606 & ~n2607;
  assign n2838 = po40  & n2837;
  assign n2839 = ~n2612 & ~n2838;
  assign n2840 = n2612 & n2838;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = ~n2836 & ~n2841;
  assign n2843 = ~n2835 & ~n2842;
  assign n2844 = po49  & ~n2843;
  assign n2845 = ~po49  & n2843;
  assign n2846 = ~n2615 & ~n2616;
  assign n2847 = po40  & n2846;
  assign n2848 = ~n2621 & ~n2847;
  assign n2849 = n2621 & n2847;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = ~n2845 & ~n2850;
  assign n2852 = ~n2844 & ~n2851;
  assign n2853 = po50  & ~n2852;
  assign n2854 = ~po50  & n2852;
  assign n2855 = ~n2624 & ~n2625;
  assign n2856 = po40  & n2855;
  assign n2857 = ~n2630 & ~n2856;
  assign n2858 = n2630 & n2856;
  assign n2859 = ~n2857 & ~n2858;
  assign n2860 = ~n2854 & ~n2859;
  assign n2861 = ~n2853 & ~n2860;
  assign n2862 = po51  & ~n2861;
  assign n2863 = ~po51  & n2861;
  assign n2864 = ~n2633 & ~n2634;
  assign n2865 = po40  & n2864;
  assign n2866 = ~n2639 & ~n2865;
  assign n2867 = n2639 & n2865;
  assign n2868 = ~n2866 & ~n2867;
  assign n2869 = ~n2863 & ~n2868;
  assign n2870 = ~n2862 & ~n2869;
  assign n2871 = po52  & ~n2870;
  assign n2872 = ~po52  & n2870;
  assign n2873 = ~n2642 & ~n2643;
  assign n2874 = po40  & n2873;
  assign n2875 = ~n2648 & ~n2874;
  assign n2876 = n2648 & n2874;
  assign n2877 = ~n2875 & ~n2876;
  assign n2878 = ~n2872 & ~n2877;
  assign n2879 = ~n2871 & ~n2878;
  assign n2880 = po53  & ~n2879;
  assign n2881 = ~po53  & n2879;
  assign n2882 = ~n2651 & ~n2652;
  assign n2883 = po40  & n2882;
  assign n2884 = ~n2657 & ~n2883;
  assign n2885 = n2657 & n2883;
  assign n2886 = ~n2884 & ~n2885;
  assign n2887 = ~n2881 & ~n2886;
  assign n2888 = ~n2880 & ~n2887;
  assign n2889 = po54  & ~n2888;
  assign n2890 = ~po54  & n2888;
  assign n2891 = ~n2660 & ~n2661;
  assign n2892 = po40  & n2891;
  assign n2893 = ~n2666 & ~n2892;
  assign n2894 = n2666 & n2892;
  assign n2895 = ~n2893 & ~n2894;
  assign n2896 = ~n2890 & ~n2895;
  assign n2897 = ~n2889 & ~n2896;
  assign n2898 = po55  & ~n2897;
  assign n2899 = ~po55  & n2897;
  assign n2900 = ~n2669 & ~n2670;
  assign n2901 = po40  & n2900;
  assign n2902 = ~n2675 & ~n2901;
  assign n2903 = n2675 & n2901;
  assign n2904 = ~n2902 & ~n2903;
  assign n2905 = ~n2899 & ~n2904;
  assign n2906 = ~n2898 & ~n2905;
  assign n2907 = po56  & ~n2906;
  assign n2908 = ~n2678 & ~n2684;
  assign n2909 = po40  & n2908;
  assign n2910 = ~n2683 & ~n2909;
  assign n2911 = n2683 & n2909;
  assign n2912 = ~n2910 & ~n2911;
  assign n2913 = ~po56  & n2906;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = ~n2907 & ~n2914;
  assign n2916 = po57  & ~n2915;
  assign n2917 = ~po57  & n2915;
  assign n2918 = ~n2758 & ~n2917;
  assign n2919 = ~n2916 & ~n2918;
  assign n2920 = po58  & ~n2919;
  assign n2921 = ~po58  & n2919;
  assign n2922 = ~n2691 & ~n2692;
  assign n2923 = po40  & n2922;
  assign n2924 = ~n2697 & ~n2923;
  assign n2925 = n2697 & n2923;
  assign n2926 = ~n2924 & ~n2925;
  assign n2927 = ~n2921 & ~n2926;
  assign n2928 = ~n2920 & ~n2927;
  assign n2929 = po59  & ~n2928;
  assign n2930 = ~po59  & n2928;
  assign n2931 = ~n2700 & ~n2701;
  assign n2932 = po40  & n2931;
  assign n2933 = ~n2706 & ~n2932;
  assign n2934 = n2706 & n2932;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = ~n2930 & ~n2935;
  assign n2937 = ~n2929 & ~n2936;
  assign n2938 = po60  & ~n2937;
  assign n2939 = ~po60  & n2937;
  assign n2940 = ~n2709 & ~n2710;
  assign n2941 = po40  & n2940;
  assign n2942 = ~n2715 & ~n2941;
  assign n2943 = n2715 & n2941;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = ~n2939 & ~n2944;
  assign n2946 = ~n2938 & ~n2945;
  assign n2947 = po61  & ~n2946;
  assign n2948 = ~po61  & n2946;
  assign n2949 = ~n2718 & ~n2719;
  assign n2950 = po40  & n2949;
  assign n2951 = ~n2724 & ~n2950;
  assign n2952 = n2724 & n2950;
  assign n2953 = ~n2951 & ~n2952;
  assign n2954 = ~n2948 & ~n2953;
  assign n2955 = ~n2947 & ~n2954;
  assign n2956 = po62  & ~n2955;
  assign n2957 = ~po62  & n2955;
  assign n2958 = ~n2727 & ~n2728;
  assign n2959 = po40  & n2958;
  assign n2960 = ~n2733 & ~n2959;
  assign n2961 = n2733 & n2959;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = ~n2957 & ~n2962;
  assign n2964 = ~n2956 & ~n2963;
  assign n2965 = n2768 & n2964;
  assign n2966 = ~n2768 & ~n2964;
  assign n2967 = n2746 & po40 ;
  assign n2968 = ~n2745 & ~n2967;
  assign n2969 = n2966 & n2968;
  assign n2970 = ~po63  & ~n2969;
  assign n2971 = ~n2965 & ~n2970;
  assign n2972 = ~n2763 & n2971;
  assign po39  = n2759 | ~n2972;
  assign n2974 = ~n2916 & ~n2917;
  assign n2975 = po39  & n2974;
  assign n2976 = ~n2758 & ~n2975;
  assign n2977 = n2758 & n2975;
  assign n2978 = ~n2976 & ~n2977;
  assign n2979 = n2768 & ~po39 ;
  assign n2980 = ~n2768 & po39 ;
  assign n2981 = n2964 & ~n2980;
  assign n2982 = po63  & ~n2981;
  assign n2983 = ~n2966 & n2982;
  assign n2984 = ~n2956 & ~n2957;
  assign n2985 = po39  & n2984;
  assign n2986 = ~n2962 & ~n2985;
  assign n2987 = n2962 & n2985;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = pi78  & po39 ;
  assign n2990 = ~pi76  & ~pi77 ;
  assign n2991 = ~pi78  & n2990;
  assign n2992 = ~n2989 & ~n2991;
  assign n2993 = po40  & ~n2992;
  assign n2994 = ~po40  & n2992;
  assign n2995 = ~pi78  & po39 ;
  assign n2996 = pi79  & ~n2995;
  assign n2997 = n2770 & po39 ;
  assign n2998 = ~n2996 & ~n2997;
  assign n2999 = ~n2994 & n2998;
  assign n3000 = ~n2993 & ~n2999;
  assign n3001 = po41  & ~n3000;
  assign n3002 = ~po41  & n3000;
  assign n3003 = po40  & n2972;
  assign n3004 = ~n2997 & ~n3003;
  assign n3005 = pi80  & ~n3004;
  assign n3006 = ~pi80  & n3004;
  assign n3007 = ~n3005 & ~n3006;
  assign n3008 = ~n3002 & ~n3007;
  assign n3009 = ~n3001 & ~n3008;
  assign n3010 = po42  & ~n3009;
  assign n3011 = ~po42  & n3009;
  assign n3012 = ~n2773 & ~n2774;
  assign n3013 = po39  & n3012;
  assign n3014 = n2778 & ~n3013;
  assign n3015 = ~n2778 & n3013;
  assign n3016 = ~n3014 & ~n3015;
  assign n3017 = ~n3011 & ~n3016;
  assign n3018 = ~n3010 & ~n3017;
  assign n3019 = po43  & ~n3018;
  assign n3020 = ~po43  & n3018;
  assign n3021 = ~n2781 & ~n2782;
  assign n3022 = po39  & n3021;
  assign n3023 = ~n2787 & ~n3022;
  assign n3024 = n2787 & n3022;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = ~n3020 & ~n3025;
  assign n3027 = ~n3019 & ~n3026;
  assign n3028 = po44  & ~n3027;
  assign n3029 = ~po44  & n3027;
  assign n3030 = ~n2790 & ~n2791;
  assign n3031 = po39  & n3030;
  assign n3032 = n2796 & n3031;
  assign n3033 = ~n2796 & ~n3031;
  assign n3034 = ~n3032 & ~n3033;
  assign n3035 = ~n3029 & ~n3034;
  assign n3036 = ~n3028 & ~n3035;
  assign n3037 = po45  & ~n3036;
  assign n3038 = ~po45  & n3036;
  assign n3039 = ~n2799 & ~n2800;
  assign n3040 = po39  & n3039;
  assign n3041 = ~n2805 & ~n3040;
  assign n3042 = n2805 & n3040;
  assign n3043 = ~n3041 & ~n3042;
  assign n3044 = ~n3038 & ~n3043;
  assign n3045 = ~n3037 & ~n3044;
  assign n3046 = po46  & ~n3045;
  assign n3047 = ~po46  & n3045;
  assign n3048 = ~n2808 & ~n2809;
  assign n3049 = po39  & n3048;
  assign n3050 = ~n2814 & ~n3049;
  assign n3051 = n2814 & n3049;
  assign n3052 = ~n3050 & ~n3051;
  assign n3053 = ~n3047 & ~n3052;
  assign n3054 = ~n3046 & ~n3053;
  assign n3055 = po47  & ~n3054;
  assign n3056 = ~po47  & n3054;
  assign n3057 = ~n2817 & ~n2818;
  assign n3058 = po39  & n3057;
  assign n3059 = ~n2823 & ~n3058;
  assign n3060 = n2823 & n3058;
  assign n3061 = ~n3059 & ~n3060;
  assign n3062 = ~n3056 & ~n3061;
  assign n3063 = ~n3055 & ~n3062;
  assign n3064 = po48  & ~n3063;
  assign n3065 = ~po48  & n3063;
  assign n3066 = ~n2826 & ~n2827;
  assign n3067 = po39  & n3066;
  assign n3068 = ~n2832 & ~n3067;
  assign n3069 = n2832 & n3067;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = ~n3065 & ~n3070;
  assign n3072 = ~n3064 & ~n3071;
  assign n3073 = po49  & ~n3072;
  assign n3074 = ~po49  & n3072;
  assign n3075 = ~n2835 & ~n2836;
  assign n3076 = po39  & n3075;
  assign n3077 = ~n2841 & ~n3076;
  assign n3078 = n2841 & n3076;
  assign n3079 = ~n3077 & ~n3078;
  assign n3080 = ~n3074 & ~n3079;
  assign n3081 = ~n3073 & ~n3080;
  assign n3082 = po50  & ~n3081;
  assign n3083 = ~po50  & n3081;
  assign n3084 = ~n2844 & ~n2845;
  assign n3085 = po39  & n3084;
  assign n3086 = ~n2850 & ~n3085;
  assign n3087 = n2850 & n3085;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = ~n3083 & ~n3088;
  assign n3090 = ~n3082 & ~n3089;
  assign n3091 = po51  & ~n3090;
  assign n3092 = ~po51  & n3090;
  assign n3093 = ~n2853 & ~n2854;
  assign n3094 = po39  & n3093;
  assign n3095 = ~n2859 & ~n3094;
  assign n3096 = n2859 & n3094;
  assign n3097 = ~n3095 & ~n3096;
  assign n3098 = ~n3092 & ~n3097;
  assign n3099 = ~n3091 & ~n3098;
  assign n3100 = po52  & ~n3099;
  assign n3101 = ~po52  & n3099;
  assign n3102 = ~n2862 & ~n2863;
  assign n3103 = po39  & n3102;
  assign n3104 = ~n2868 & ~n3103;
  assign n3105 = n2868 & n3103;
  assign n3106 = ~n3104 & ~n3105;
  assign n3107 = ~n3101 & ~n3106;
  assign n3108 = ~n3100 & ~n3107;
  assign n3109 = po53  & ~n3108;
  assign n3110 = ~po53  & n3108;
  assign n3111 = ~n2871 & ~n2872;
  assign n3112 = po39  & n3111;
  assign n3113 = ~n2877 & ~n3112;
  assign n3114 = n2877 & n3112;
  assign n3115 = ~n3113 & ~n3114;
  assign n3116 = ~n3110 & ~n3115;
  assign n3117 = ~n3109 & ~n3116;
  assign n3118 = po54  & ~n3117;
  assign n3119 = ~po54  & n3117;
  assign n3120 = ~n2880 & ~n2881;
  assign n3121 = po39  & n3120;
  assign n3122 = ~n2886 & ~n3121;
  assign n3123 = n2886 & n3121;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = ~n3119 & ~n3124;
  assign n3126 = ~n3118 & ~n3125;
  assign n3127 = po55  & ~n3126;
  assign n3128 = ~po55  & n3126;
  assign n3129 = ~n2889 & ~n2890;
  assign n3130 = po39  & n3129;
  assign n3131 = ~n2895 & ~n3130;
  assign n3132 = n2895 & n3130;
  assign n3133 = ~n3131 & ~n3132;
  assign n3134 = ~n3128 & ~n3133;
  assign n3135 = ~n3127 & ~n3134;
  assign n3136 = po56  & ~n3135;
  assign n3137 = ~po56  & n3135;
  assign n3138 = ~n2898 & ~n2899;
  assign n3139 = po39  & n3138;
  assign n3140 = ~n2904 & ~n3139;
  assign n3141 = n2904 & n3139;
  assign n3142 = ~n3140 & ~n3141;
  assign n3143 = ~n3137 & ~n3142;
  assign n3144 = ~n3136 & ~n3143;
  assign n3145 = po57  & ~n3144;
  assign n3146 = ~n2907 & ~n2913;
  assign n3147 = po39  & n3146;
  assign n3148 = ~n2912 & ~n3147;
  assign n3149 = n2912 & n3147;
  assign n3150 = ~n3148 & ~n3149;
  assign n3151 = ~po57  & n3144;
  assign n3152 = ~n3150 & ~n3151;
  assign n3153 = ~n3145 & ~n3152;
  assign n3154 = po58  & ~n3153;
  assign n3155 = ~po58  & n3153;
  assign n3156 = ~n2978 & ~n3155;
  assign n3157 = ~n3154 & ~n3156;
  assign n3158 = po59  & ~n3157;
  assign n3159 = ~po59  & n3157;
  assign n3160 = ~n2920 & ~n2921;
  assign n3161 = po39  & n3160;
  assign n3162 = ~n2926 & ~n3161;
  assign n3163 = n2926 & n3161;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = ~n3159 & ~n3164;
  assign n3166 = ~n3158 & ~n3165;
  assign n3167 = po60  & ~n3166;
  assign n3168 = ~po60  & n3166;
  assign n3169 = ~n2929 & ~n2930;
  assign n3170 = po39  & n3169;
  assign n3171 = ~n2935 & ~n3170;
  assign n3172 = n2935 & n3170;
  assign n3173 = ~n3171 & ~n3172;
  assign n3174 = ~n3168 & ~n3173;
  assign n3175 = ~n3167 & ~n3174;
  assign n3176 = po61  & ~n3175;
  assign n3177 = ~po61  & n3175;
  assign n3178 = ~n2938 & ~n2939;
  assign n3179 = po39  & n3178;
  assign n3180 = ~n2944 & ~n3179;
  assign n3181 = n2944 & n3179;
  assign n3182 = ~n3180 & ~n3181;
  assign n3183 = ~n3177 & ~n3182;
  assign n3184 = ~n3176 & ~n3183;
  assign n3185 = po62  & ~n3184;
  assign n3186 = ~po62  & n3184;
  assign n3187 = ~n2947 & ~n2948;
  assign n3188 = po39  & n3187;
  assign n3189 = ~n2953 & ~n3188;
  assign n3190 = n2953 & n3188;
  assign n3191 = ~n3189 & ~n3190;
  assign n3192 = ~n3186 & ~n3191;
  assign n3193 = ~n3185 & ~n3192;
  assign n3194 = n2988 & n3193;
  assign n3195 = ~n2988 & ~n3193;
  assign n3196 = n2966 & po39 ;
  assign n3197 = ~n2965 & ~n3196;
  assign n3198 = n3195 & n3197;
  assign n3199 = ~po63  & ~n3198;
  assign n3200 = ~n3194 & ~n3199;
  assign n3201 = ~n2983 & n3200;
  assign po38  = n2979 | ~n3201;
  assign n3203 = ~n3154 & ~n3155;
  assign n3204 = po38  & n3203;
  assign n3205 = ~n2978 & ~n3204;
  assign n3206 = n2978 & n3204;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = n2988 & ~po38 ;
  assign n3209 = ~n2988 & po38 ;
  assign n3210 = n3193 & ~n3209;
  assign n3211 = po63  & ~n3210;
  assign n3212 = ~n3195 & n3211;
  assign n3213 = ~n3185 & ~n3186;
  assign n3214 = po38  & n3213;
  assign n3215 = ~n3191 & ~n3214;
  assign n3216 = n3191 & n3214;
  assign n3217 = ~n3215 & ~n3216;
  assign n3218 = pi76  & po38 ;
  assign n3219 = ~pi74  & ~pi75 ;
  assign n3220 = ~pi76  & n3219;
  assign n3221 = ~n3218 & ~n3220;
  assign n3222 = po39  & ~n3221;
  assign n3223 = ~po39  & n3221;
  assign n3224 = ~pi76  & po38 ;
  assign n3225 = pi77  & ~n3224;
  assign n3226 = n2990 & po38 ;
  assign n3227 = ~n3225 & ~n3226;
  assign n3228 = ~n3223 & n3227;
  assign n3229 = ~n3222 & ~n3228;
  assign n3230 = po40  & ~n3229;
  assign n3231 = ~po40  & n3229;
  assign n3232 = po39  & n3201;
  assign n3233 = ~n3226 & ~n3232;
  assign n3234 = pi78  & ~n3233;
  assign n3235 = ~pi78  & n3233;
  assign n3236 = ~n3234 & ~n3235;
  assign n3237 = ~n3231 & ~n3236;
  assign n3238 = ~n3230 & ~n3237;
  assign n3239 = po41  & ~n3238;
  assign n3240 = ~po41  & n3238;
  assign n3241 = ~n2993 & ~n2994;
  assign n3242 = po38  & n3241;
  assign n3243 = n2998 & ~n3242;
  assign n3244 = ~n2998 & n3242;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = ~n3240 & ~n3245;
  assign n3247 = ~n3239 & ~n3246;
  assign n3248 = po42  & ~n3247;
  assign n3249 = ~po42  & n3247;
  assign n3250 = ~n3001 & ~n3002;
  assign n3251 = po38  & n3250;
  assign n3252 = ~n3007 & ~n3251;
  assign n3253 = n3007 & n3251;
  assign n3254 = ~n3252 & ~n3253;
  assign n3255 = ~n3249 & ~n3254;
  assign n3256 = ~n3248 & ~n3255;
  assign n3257 = po43  & ~n3256;
  assign n3258 = ~po43  & n3256;
  assign n3259 = ~n3010 & ~n3011;
  assign n3260 = po38  & n3259;
  assign n3261 = n3016 & n3260;
  assign n3262 = ~n3016 & ~n3260;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = ~n3258 & ~n3263;
  assign n3265 = ~n3257 & ~n3264;
  assign n3266 = po44  & ~n3265;
  assign n3267 = ~po44  & n3265;
  assign n3268 = ~n3019 & ~n3020;
  assign n3269 = po38  & n3268;
  assign n3270 = ~n3025 & ~n3269;
  assign n3271 = n3025 & n3269;
  assign n3272 = ~n3270 & ~n3271;
  assign n3273 = ~n3267 & ~n3272;
  assign n3274 = ~n3266 & ~n3273;
  assign n3275 = po45  & ~n3274;
  assign n3276 = ~po45  & n3274;
  assign n3277 = ~n3028 & ~n3029;
  assign n3278 = po38  & n3277;
  assign n3279 = ~n3034 & ~n3278;
  assign n3280 = n3034 & n3278;
  assign n3281 = ~n3279 & ~n3280;
  assign n3282 = ~n3276 & ~n3281;
  assign n3283 = ~n3275 & ~n3282;
  assign n3284 = po46  & ~n3283;
  assign n3285 = ~po46  & n3283;
  assign n3286 = ~n3037 & ~n3038;
  assign n3287 = po38  & n3286;
  assign n3288 = ~n3043 & ~n3287;
  assign n3289 = n3043 & n3287;
  assign n3290 = ~n3288 & ~n3289;
  assign n3291 = ~n3285 & ~n3290;
  assign n3292 = ~n3284 & ~n3291;
  assign n3293 = po47  & ~n3292;
  assign n3294 = ~po47  & n3292;
  assign n3295 = ~n3046 & ~n3047;
  assign n3296 = po38  & n3295;
  assign n3297 = ~n3052 & ~n3296;
  assign n3298 = n3052 & n3296;
  assign n3299 = ~n3297 & ~n3298;
  assign n3300 = ~n3294 & ~n3299;
  assign n3301 = ~n3293 & ~n3300;
  assign n3302 = po48  & ~n3301;
  assign n3303 = ~po48  & n3301;
  assign n3304 = ~n3055 & ~n3056;
  assign n3305 = po38  & n3304;
  assign n3306 = ~n3061 & ~n3305;
  assign n3307 = n3061 & n3305;
  assign n3308 = ~n3306 & ~n3307;
  assign n3309 = ~n3303 & ~n3308;
  assign n3310 = ~n3302 & ~n3309;
  assign n3311 = po49  & ~n3310;
  assign n3312 = ~po49  & n3310;
  assign n3313 = ~n3064 & ~n3065;
  assign n3314 = po38  & n3313;
  assign n3315 = ~n3070 & ~n3314;
  assign n3316 = n3070 & n3314;
  assign n3317 = ~n3315 & ~n3316;
  assign n3318 = ~n3312 & ~n3317;
  assign n3319 = ~n3311 & ~n3318;
  assign n3320 = po50  & ~n3319;
  assign n3321 = ~po50  & n3319;
  assign n3322 = ~n3073 & ~n3074;
  assign n3323 = po38  & n3322;
  assign n3324 = ~n3079 & ~n3323;
  assign n3325 = n3079 & n3323;
  assign n3326 = ~n3324 & ~n3325;
  assign n3327 = ~n3321 & ~n3326;
  assign n3328 = ~n3320 & ~n3327;
  assign n3329 = po51  & ~n3328;
  assign n3330 = ~po51  & n3328;
  assign n3331 = ~n3082 & ~n3083;
  assign n3332 = po38  & n3331;
  assign n3333 = ~n3088 & ~n3332;
  assign n3334 = n3088 & n3332;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = ~n3330 & ~n3335;
  assign n3337 = ~n3329 & ~n3336;
  assign n3338 = po52  & ~n3337;
  assign n3339 = ~po52  & n3337;
  assign n3340 = ~n3091 & ~n3092;
  assign n3341 = po38  & n3340;
  assign n3342 = ~n3097 & ~n3341;
  assign n3343 = n3097 & n3341;
  assign n3344 = ~n3342 & ~n3343;
  assign n3345 = ~n3339 & ~n3344;
  assign n3346 = ~n3338 & ~n3345;
  assign n3347 = po53  & ~n3346;
  assign n3348 = ~po53  & n3346;
  assign n3349 = ~n3100 & ~n3101;
  assign n3350 = po38  & n3349;
  assign n3351 = ~n3106 & ~n3350;
  assign n3352 = n3106 & n3350;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = ~n3348 & ~n3353;
  assign n3355 = ~n3347 & ~n3354;
  assign n3356 = po54  & ~n3355;
  assign n3357 = ~po54  & n3355;
  assign n3358 = ~n3109 & ~n3110;
  assign n3359 = po38  & n3358;
  assign n3360 = ~n3115 & ~n3359;
  assign n3361 = n3115 & n3359;
  assign n3362 = ~n3360 & ~n3361;
  assign n3363 = ~n3357 & ~n3362;
  assign n3364 = ~n3356 & ~n3363;
  assign n3365 = po55  & ~n3364;
  assign n3366 = ~po55  & n3364;
  assign n3367 = ~n3118 & ~n3119;
  assign n3368 = po38  & n3367;
  assign n3369 = ~n3124 & ~n3368;
  assign n3370 = n3124 & n3368;
  assign n3371 = ~n3369 & ~n3370;
  assign n3372 = ~n3366 & ~n3371;
  assign n3373 = ~n3365 & ~n3372;
  assign n3374 = po56  & ~n3373;
  assign n3375 = ~po56  & n3373;
  assign n3376 = ~n3127 & ~n3128;
  assign n3377 = po38  & n3376;
  assign n3378 = ~n3133 & ~n3377;
  assign n3379 = n3133 & n3377;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = ~n3375 & ~n3380;
  assign n3382 = ~n3374 & ~n3381;
  assign n3383 = po57  & ~n3382;
  assign n3384 = ~po57  & n3382;
  assign n3385 = ~n3136 & ~n3137;
  assign n3386 = po38  & n3385;
  assign n3387 = ~n3142 & ~n3386;
  assign n3388 = n3142 & n3386;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = ~n3384 & ~n3389;
  assign n3391 = ~n3383 & ~n3390;
  assign n3392 = po58  & ~n3391;
  assign n3393 = ~n3145 & ~n3151;
  assign n3394 = po38  & n3393;
  assign n3395 = ~n3150 & ~n3394;
  assign n3396 = n3150 & n3394;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = ~po58  & n3391;
  assign n3399 = ~n3397 & ~n3398;
  assign n3400 = ~n3392 & ~n3399;
  assign n3401 = po59  & ~n3400;
  assign n3402 = ~po59  & n3400;
  assign n3403 = ~n3207 & ~n3402;
  assign n3404 = ~n3401 & ~n3403;
  assign n3405 = po60  & ~n3404;
  assign n3406 = ~po60  & n3404;
  assign n3407 = ~n3158 & ~n3159;
  assign n3408 = po38  & n3407;
  assign n3409 = ~n3164 & ~n3408;
  assign n3410 = n3164 & n3408;
  assign n3411 = ~n3409 & ~n3410;
  assign n3412 = ~n3406 & ~n3411;
  assign n3413 = ~n3405 & ~n3412;
  assign n3414 = po61  & ~n3413;
  assign n3415 = ~po61  & n3413;
  assign n3416 = ~n3167 & ~n3168;
  assign n3417 = po38  & n3416;
  assign n3418 = ~n3173 & ~n3417;
  assign n3419 = n3173 & n3417;
  assign n3420 = ~n3418 & ~n3419;
  assign n3421 = ~n3415 & ~n3420;
  assign n3422 = ~n3414 & ~n3421;
  assign n3423 = po62  & ~n3422;
  assign n3424 = ~po62  & n3422;
  assign n3425 = ~n3176 & ~n3177;
  assign n3426 = po38  & n3425;
  assign n3427 = ~n3182 & ~n3426;
  assign n3428 = n3182 & n3426;
  assign n3429 = ~n3427 & ~n3428;
  assign n3430 = ~n3424 & ~n3429;
  assign n3431 = ~n3423 & ~n3430;
  assign n3432 = n3217 & n3431;
  assign n3433 = ~n3217 & ~n3431;
  assign n3434 = n3195 & po38 ;
  assign n3435 = ~n3194 & ~n3434;
  assign n3436 = n3433 & n3435;
  assign n3437 = ~po63  & ~n3436;
  assign n3438 = ~n3432 & ~n3437;
  assign n3439 = ~n3212 & n3438;
  assign po37  = n3208 | ~n3439;
  assign n3441 = ~n3401 & ~n3402;
  assign n3442 = po37  & n3441;
  assign n3443 = ~n3207 & ~n3442;
  assign n3444 = n3207 & n3442;
  assign n3445 = ~n3443 & ~n3444;
  assign n3446 = n3217 & ~po37 ;
  assign n3447 = ~n3217 & po37 ;
  assign n3448 = n3431 & ~n3447;
  assign n3449 = po63  & ~n3448;
  assign n3450 = ~n3433 & n3449;
  assign n3451 = ~n3423 & ~n3424;
  assign n3452 = po37  & n3451;
  assign n3453 = ~n3429 & ~n3452;
  assign n3454 = n3429 & n3452;
  assign n3455 = ~n3453 & ~n3454;
  assign n3456 = pi74  & po37 ;
  assign n3457 = ~pi72  & ~pi73 ;
  assign n3458 = ~pi74  & n3457;
  assign n3459 = ~n3456 & ~n3458;
  assign n3460 = po38  & ~n3459;
  assign n3461 = ~po38  & n3459;
  assign n3462 = ~pi74  & po37 ;
  assign n3463 = pi75  & ~n3462;
  assign n3464 = n3219 & po37 ;
  assign n3465 = ~n3463 & ~n3464;
  assign n3466 = ~n3461 & n3465;
  assign n3467 = ~n3460 & ~n3466;
  assign n3468 = po39  & ~n3467;
  assign n3469 = ~po39  & n3467;
  assign n3470 = po38  & n3439;
  assign n3471 = ~n3464 & ~n3470;
  assign n3472 = pi76  & ~n3471;
  assign n3473 = ~pi76  & n3471;
  assign n3474 = ~n3472 & ~n3473;
  assign n3475 = ~n3469 & ~n3474;
  assign n3476 = ~n3468 & ~n3475;
  assign n3477 = po40  & ~n3476;
  assign n3478 = ~po40  & n3476;
  assign n3479 = ~n3222 & ~n3223;
  assign n3480 = po37  & n3479;
  assign n3481 = n3227 & ~n3480;
  assign n3482 = ~n3227 & n3480;
  assign n3483 = ~n3481 & ~n3482;
  assign n3484 = ~n3478 & ~n3483;
  assign n3485 = ~n3477 & ~n3484;
  assign n3486 = po41  & ~n3485;
  assign n3487 = ~po41  & n3485;
  assign n3488 = ~n3230 & ~n3231;
  assign n3489 = po37  & n3488;
  assign n3490 = ~n3236 & ~n3489;
  assign n3491 = n3236 & n3489;
  assign n3492 = ~n3490 & ~n3491;
  assign n3493 = ~n3487 & ~n3492;
  assign n3494 = ~n3486 & ~n3493;
  assign n3495 = po42  & ~n3494;
  assign n3496 = ~po42  & n3494;
  assign n3497 = ~n3239 & ~n3240;
  assign n3498 = po37  & n3497;
  assign n3499 = n3245 & n3498;
  assign n3500 = ~n3245 & ~n3498;
  assign n3501 = ~n3499 & ~n3500;
  assign n3502 = ~n3496 & ~n3501;
  assign n3503 = ~n3495 & ~n3502;
  assign n3504 = po43  & ~n3503;
  assign n3505 = ~po43  & n3503;
  assign n3506 = ~n3248 & ~n3249;
  assign n3507 = po37  & n3506;
  assign n3508 = ~n3254 & ~n3507;
  assign n3509 = n3254 & n3507;
  assign n3510 = ~n3508 & ~n3509;
  assign n3511 = ~n3505 & ~n3510;
  assign n3512 = ~n3504 & ~n3511;
  assign n3513 = po44  & ~n3512;
  assign n3514 = ~po44  & n3512;
  assign n3515 = ~n3257 & ~n3258;
  assign n3516 = po37  & n3515;
  assign n3517 = ~n3263 & ~n3516;
  assign n3518 = n3263 & n3516;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520 = ~n3514 & ~n3519;
  assign n3521 = ~n3513 & ~n3520;
  assign n3522 = po45  & ~n3521;
  assign n3523 = ~po45  & n3521;
  assign n3524 = ~n3266 & ~n3267;
  assign n3525 = po37  & n3524;
  assign n3526 = ~n3272 & ~n3525;
  assign n3527 = n3272 & n3525;
  assign n3528 = ~n3526 & ~n3527;
  assign n3529 = ~n3523 & ~n3528;
  assign n3530 = ~n3522 & ~n3529;
  assign n3531 = po46  & ~n3530;
  assign n3532 = ~po46  & n3530;
  assign n3533 = ~n3275 & ~n3276;
  assign n3534 = po37  & n3533;
  assign n3535 = ~n3281 & ~n3534;
  assign n3536 = n3281 & n3534;
  assign n3537 = ~n3535 & ~n3536;
  assign n3538 = ~n3532 & ~n3537;
  assign n3539 = ~n3531 & ~n3538;
  assign n3540 = po47  & ~n3539;
  assign n3541 = ~po47  & n3539;
  assign n3542 = ~n3284 & ~n3285;
  assign n3543 = po37  & n3542;
  assign n3544 = ~n3290 & ~n3543;
  assign n3545 = n3290 & n3543;
  assign n3546 = ~n3544 & ~n3545;
  assign n3547 = ~n3541 & ~n3546;
  assign n3548 = ~n3540 & ~n3547;
  assign n3549 = po48  & ~n3548;
  assign n3550 = ~po48  & n3548;
  assign n3551 = ~n3293 & ~n3294;
  assign n3552 = po37  & n3551;
  assign n3553 = ~n3299 & ~n3552;
  assign n3554 = n3299 & n3552;
  assign n3555 = ~n3553 & ~n3554;
  assign n3556 = ~n3550 & ~n3555;
  assign n3557 = ~n3549 & ~n3556;
  assign n3558 = po49  & ~n3557;
  assign n3559 = ~po49  & n3557;
  assign n3560 = ~n3302 & ~n3303;
  assign n3561 = po37  & n3560;
  assign n3562 = ~n3308 & ~n3561;
  assign n3563 = n3308 & n3561;
  assign n3564 = ~n3562 & ~n3563;
  assign n3565 = ~n3559 & ~n3564;
  assign n3566 = ~n3558 & ~n3565;
  assign n3567 = po50  & ~n3566;
  assign n3568 = ~po50  & n3566;
  assign n3569 = ~n3311 & ~n3312;
  assign n3570 = po37  & n3569;
  assign n3571 = ~n3317 & ~n3570;
  assign n3572 = n3317 & n3570;
  assign n3573 = ~n3571 & ~n3572;
  assign n3574 = ~n3568 & ~n3573;
  assign n3575 = ~n3567 & ~n3574;
  assign n3576 = po51  & ~n3575;
  assign n3577 = ~po51  & n3575;
  assign n3578 = ~n3320 & ~n3321;
  assign n3579 = po37  & n3578;
  assign n3580 = ~n3326 & ~n3579;
  assign n3581 = n3326 & n3579;
  assign n3582 = ~n3580 & ~n3581;
  assign n3583 = ~n3577 & ~n3582;
  assign n3584 = ~n3576 & ~n3583;
  assign n3585 = po52  & ~n3584;
  assign n3586 = ~po52  & n3584;
  assign n3587 = ~n3329 & ~n3330;
  assign n3588 = po37  & n3587;
  assign n3589 = ~n3335 & ~n3588;
  assign n3590 = n3335 & n3588;
  assign n3591 = ~n3589 & ~n3590;
  assign n3592 = ~n3586 & ~n3591;
  assign n3593 = ~n3585 & ~n3592;
  assign n3594 = po53  & ~n3593;
  assign n3595 = ~po53  & n3593;
  assign n3596 = ~n3338 & ~n3339;
  assign n3597 = po37  & n3596;
  assign n3598 = ~n3344 & ~n3597;
  assign n3599 = n3344 & n3597;
  assign n3600 = ~n3598 & ~n3599;
  assign n3601 = ~n3595 & ~n3600;
  assign n3602 = ~n3594 & ~n3601;
  assign n3603 = po54  & ~n3602;
  assign n3604 = ~po54  & n3602;
  assign n3605 = ~n3347 & ~n3348;
  assign n3606 = po37  & n3605;
  assign n3607 = ~n3353 & ~n3606;
  assign n3608 = n3353 & n3606;
  assign n3609 = ~n3607 & ~n3608;
  assign n3610 = ~n3604 & ~n3609;
  assign n3611 = ~n3603 & ~n3610;
  assign n3612 = po55  & ~n3611;
  assign n3613 = ~po55  & n3611;
  assign n3614 = ~n3356 & ~n3357;
  assign n3615 = po37  & n3614;
  assign n3616 = ~n3362 & ~n3615;
  assign n3617 = n3362 & n3615;
  assign n3618 = ~n3616 & ~n3617;
  assign n3619 = ~n3613 & ~n3618;
  assign n3620 = ~n3612 & ~n3619;
  assign n3621 = po56  & ~n3620;
  assign n3622 = ~po56  & n3620;
  assign n3623 = ~n3365 & ~n3366;
  assign n3624 = po37  & n3623;
  assign n3625 = ~n3371 & ~n3624;
  assign n3626 = n3371 & n3624;
  assign n3627 = ~n3625 & ~n3626;
  assign n3628 = ~n3622 & ~n3627;
  assign n3629 = ~n3621 & ~n3628;
  assign n3630 = po57  & ~n3629;
  assign n3631 = ~po57  & n3629;
  assign n3632 = ~n3374 & ~n3375;
  assign n3633 = po37  & n3632;
  assign n3634 = ~n3380 & ~n3633;
  assign n3635 = n3380 & n3633;
  assign n3636 = ~n3634 & ~n3635;
  assign n3637 = ~n3631 & ~n3636;
  assign n3638 = ~n3630 & ~n3637;
  assign n3639 = po58  & ~n3638;
  assign n3640 = ~po58  & n3638;
  assign n3641 = ~n3383 & ~n3384;
  assign n3642 = po37  & n3641;
  assign n3643 = ~n3389 & ~n3642;
  assign n3644 = n3389 & n3642;
  assign n3645 = ~n3643 & ~n3644;
  assign n3646 = ~n3640 & ~n3645;
  assign n3647 = ~n3639 & ~n3646;
  assign n3648 = po59  & ~n3647;
  assign n3649 = ~n3392 & ~n3398;
  assign n3650 = po37  & n3649;
  assign n3651 = ~n3397 & ~n3650;
  assign n3652 = n3397 & n3650;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = ~po59  & n3647;
  assign n3655 = ~n3653 & ~n3654;
  assign n3656 = ~n3648 & ~n3655;
  assign n3657 = po60  & ~n3656;
  assign n3658 = ~po60  & n3656;
  assign n3659 = ~n3445 & ~n3658;
  assign n3660 = ~n3657 & ~n3659;
  assign n3661 = po61  & ~n3660;
  assign n3662 = ~po61  & n3660;
  assign n3663 = ~n3405 & ~n3406;
  assign n3664 = po37  & n3663;
  assign n3665 = ~n3411 & ~n3664;
  assign n3666 = n3411 & n3664;
  assign n3667 = ~n3665 & ~n3666;
  assign n3668 = ~n3662 & ~n3667;
  assign n3669 = ~n3661 & ~n3668;
  assign n3670 = po62  & ~n3669;
  assign n3671 = ~po62  & n3669;
  assign n3672 = ~n3414 & ~n3415;
  assign n3673 = po37  & n3672;
  assign n3674 = ~n3420 & ~n3673;
  assign n3675 = n3420 & n3673;
  assign n3676 = ~n3674 & ~n3675;
  assign n3677 = ~n3671 & ~n3676;
  assign n3678 = ~n3670 & ~n3677;
  assign n3679 = n3455 & n3678;
  assign n3680 = ~n3455 & ~n3678;
  assign n3681 = n3433 & po37 ;
  assign n3682 = ~n3432 & ~n3681;
  assign n3683 = n3680 & n3682;
  assign n3684 = ~po63  & ~n3683;
  assign n3685 = ~n3679 & ~n3684;
  assign n3686 = ~n3450 & n3685;
  assign po36  = n3446 | ~n3686;
  assign n3688 = ~n3657 & ~n3658;
  assign n3689 = po36  & n3688;
  assign n3690 = ~n3445 & ~n3689;
  assign n3691 = n3445 & n3689;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = n3455 & ~po36 ;
  assign n3694 = ~n3455 & po36 ;
  assign n3695 = n3678 & ~n3694;
  assign n3696 = po63  & ~n3695;
  assign n3697 = ~n3680 & n3696;
  assign n3698 = ~n3670 & ~n3671;
  assign n3699 = po36  & n3698;
  assign n3700 = ~n3676 & ~n3699;
  assign n3701 = n3676 & n3699;
  assign n3702 = ~n3700 & ~n3701;
  assign n3703 = pi72  & po36 ;
  assign n3704 = ~pi70  & ~pi71 ;
  assign n3705 = ~pi72  & n3704;
  assign n3706 = ~n3703 & ~n3705;
  assign n3707 = po37  & ~n3706;
  assign n3708 = ~po37  & n3706;
  assign n3709 = ~pi72  & po36 ;
  assign n3710 = pi73  & ~n3709;
  assign n3711 = n3457 & po36 ;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = ~n3708 & n3712;
  assign n3714 = ~n3707 & ~n3713;
  assign n3715 = po38  & ~n3714;
  assign n3716 = ~po38  & n3714;
  assign n3717 = po37  & n3686;
  assign n3718 = ~n3711 & ~n3717;
  assign n3719 = pi74  & ~n3718;
  assign n3720 = ~pi74  & n3718;
  assign n3721 = ~n3719 & ~n3720;
  assign n3722 = ~n3716 & ~n3721;
  assign n3723 = ~n3715 & ~n3722;
  assign n3724 = po39  & ~n3723;
  assign n3725 = ~po39  & n3723;
  assign n3726 = ~n3460 & ~n3461;
  assign n3727 = po36  & n3726;
  assign n3728 = n3465 & ~n3727;
  assign n3729 = ~n3465 & n3727;
  assign n3730 = ~n3728 & ~n3729;
  assign n3731 = ~n3725 & ~n3730;
  assign n3732 = ~n3724 & ~n3731;
  assign n3733 = po40  & ~n3732;
  assign n3734 = ~po40  & n3732;
  assign n3735 = ~n3468 & ~n3469;
  assign n3736 = po36  & n3735;
  assign n3737 = ~n3474 & ~n3736;
  assign n3738 = n3474 & n3736;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = ~n3734 & ~n3739;
  assign n3741 = ~n3733 & ~n3740;
  assign n3742 = po41  & ~n3741;
  assign n3743 = ~po41  & n3741;
  assign n3744 = ~n3477 & ~n3478;
  assign n3745 = po36  & n3744;
  assign n3746 = n3483 & n3745;
  assign n3747 = ~n3483 & ~n3745;
  assign n3748 = ~n3746 & ~n3747;
  assign n3749 = ~n3743 & ~n3748;
  assign n3750 = ~n3742 & ~n3749;
  assign n3751 = po42  & ~n3750;
  assign n3752 = ~po42  & n3750;
  assign n3753 = ~n3486 & ~n3487;
  assign n3754 = po36  & n3753;
  assign n3755 = ~n3492 & ~n3754;
  assign n3756 = n3492 & n3754;
  assign n3757 = ~n3755 & ~n3756;
  assign n3758 = ~n3752 & ~n3757;
  assign n3759 = ~n3751 & ~n3758;
  assign n3760 = po43  & ~n3759;
  assign n3761 = ~po43  & n3759;
  assign n3762 = ~n3495 & ~n3496;
  assign n3763 = po36  & n3762;
  assign n3764 = ~n3501 & ~n3763;
  assign n3765 = n3501 & n3763;
  assign n3766 = ~n3764 & ~n3765;
  assign n3767 = ~n3761 & ~n3766;
  assign n3768 = ~n3760 & ~n3767;
  assign n3769 = po44  & ~n3768;
  assign n3770 = ~po44  & n3768;
  assign n3771 = ~n3504 & ~n3505;
  assign n3772 = po36  & n3771;
  assign n3773 = ~n3510 & ~n3772;
  assign n3774 = n3510 & n3772;
  assign n3775 = ~n3773 & ~n3774;
  assign n3776 = ~n3770 & ~n3775;
  assign n3777 = ~n3769 & ~n3776;
  assign n3778 = po45  & ~n3777;
  assign n3779 = ~po45  & n3777;
  assign n3780 = ~n3513 & ~n3514;
  assign n3781 = po36  & n3780;
  assign n3782 = ~n3519 & ~n3781;
  assign n3783 = n3519 & n3781;
  assign n3784 = ~n3782 & ~n3783;
  assign n3785 = ~n3779 & ~n3784;
  assign n3786 = ~n3778 & ~n3785;
  assign n3787 = po46  & ~n3786;
  assign n3788 = ~po46  & n3786;
  assign n3789 = ~n3522 & ~n3523;
  assign n3790 = po36  & n3789;
  assign n3791 = ~n3528 & ~n3790;
  assign n3792 = n3528 & n3790;
  assign n3793 = ~n3791 & ~n3792;
  assign n3794 = ~n3788 & ~n3793;
  assign n3795 = ~n3787 & ~n3794;
  assign n3796 = po47  & ~n3795;
  assign n3797 = ~po47  & n3795;
  assign n3798 = ~n3531 & ~n3532;
  assign n3799 = po36  & n3798;
  assign n3800 = ~n3537 & ~n3799;
  assign n3801 = n3537 & n3799;
  assign n3802 = ~n3800 & ~n3801;
  assign n3803 = ~n3797 & ~n3802;
  assign n3804 = ~n3796 & ~n3803;
  assign n3805 = po48  & ~n3804;
  assign n3806 = ~po48  & n3804;
  assign n3807 = ~n3540 & ~n3541;
  assign n3808 = po36  & n3807;
  assign n3809 = ~n3546 & ~n3808;
  assign n3810 = n3546 & n3808;
  assign n3811 = ~n3809 & ~n3810;
  assign n3812 = ~n3806 & ~n3811;
  assign n3813 = ~n3805 & ~n3812;
  assign n3814 = po49  & ~n3813;
  assign n3815 = ~po49  & n3813;
  assign n3816 = ~n3549 & ~n3550;
  assign n3817 = po36  & n3816;
  assign n3818 = ~n3555 & ~n3817;
  assign n3819 = n3555 & n3817;
  assign n3820 = ~n3818 & ~n3819;
  assign n3821 = ~n3815 & ~n3820;
  assign n3822 = ~n3814 & ~n3821;
  assign n3823 = po50  & ~n3822;
  assign n3824 = ~po50  & n3822;
  assign n3825 = ~n3558 & ~n3559;
  assign n3826 = po36  & n3825;
  assign n3827 = ~n3564 & ~n3826;
  assign n3828 = n3564 & n3826;
  assign n3829 = ~n3827 & ~n3828;
  assign n3830 = ~n3824 & ~n3829;
  assign n3831 = ~n3823 & ~n3830;
  assign n3832 = po51  & ~n3831;
  assign n3833 = ~po51  & n3831;
  assign n3834 = ~n3567 & ~n3568;
  assign n3835 = po36  & n3834;
  assign n3836 = ~n3573 & ~n3835;
  assign n3837 = n3573 & n3835;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = ~n3833 & ~n3838;
  assign n3840 = ~n3832 & ~n3839;
  assign n3841 = po52  & ~n3840;
  assign n3842 = ~po52  & n3840;
  assign n3843 = ~n3576 & ~n3577;
  assign n3844 = po36  & n3843;
  assign n3845 = ~n3582 & ~n3844;
  assign n3846 = n3582 & n3844;
  assign n3847 = ~n3845 & ~n3846;
  assign n3848 = ~n3842 & ~n3847;
  assign n3849 = ~n3841 & ~n3848;
  assign n3850 = po53  & ~n3849;
  assign n3851 = ~po53  & n3849;
  assign n3852 = ~n3585 & ~n3586;
  assign n3853 = po36  & n3852;
  assign n3854 = ~n3591 & ~n3853;
  assign n3855 = n3591 & n3853;
  assign n3856 = ~n3854 & ~n3855;
  assign n3857 = ~n3851 & ~n3856;
  assign n3858 = ~n3850 & ~n3857;
  assign n3859 = po54  & ~n3858;
  assign n3860 = ~po54  & n3858;
  assign n3861 = ~n3594 & ~n3595;
  assign n3862 = po36  & n3861;
  assign n3863 = ~n3600 & ~n3862;
  assign n3864 = n3600 & n3862;
  assign n3865 = ~n3863 & ~n3864;
  assign n3866 = ~n3860 & ~n3865;
  assign n3867 = ~n3859 & ~n3866;
  assign n3868 = po55  & ~n3867;
  assign n3869 = ~po55  & n3867;
  assign n3870 = ~n3603 & ~n3604;
  assign n3871 = po36  & n3870;
  assign n3872 = ~n3609 & ~n3871;
  assign n3873 = n3609 & n3871;
  assign n3874 = ~n3872 & ~n3873;
  assign n3875 = ~n3869 & ~n3874;
  assign n3876 = ~n3868 & ~n3875;
  assign n3877 = po56  & ~n3876;
  assign n3878 = ~po56  & n3876;
  assign n3879 = ~n3612 & ~n3613;
  assign n3880 = po36  & n3879;
  assign n3881 = ~n3618 & ~n3880;
  assign n3882 = n3618 & n3880;
  assign n3883 = ~n3881 & ~n3882;
  assign n3884 = ~n3878 & ~n3883;
  assign n3885 = ~n3877 & ~n3884;
  assign n3886 = po57  & ~n3885;
  assign n3887 = ~po57  & n3885;
  assign n3888 = ~n3621 & ~n3622;
  assign n3889 = po36  & n3888;
  assign n3890 = ~n3627 & ~n3889;
  assign n3891 = n3627 & n3889;
  assign n3892 = ~n3890 & ~n3891;
  assign n3893 = ~n3887 & ~n3892;
  assign n3894 = ~n3886 & ~n3893;
  assign n3895 = po58  & ~n3894;
  assign n3896 = ~po58  & n3894;
  assign n3897 = ~n3630 & ~n3631;
  assign n3898 = po36  & n3897;
  assign n3899 = ~n3636 & ~n3898;
  assign n3900 = n3636 & n3898;
  assign n3901 = ~n3899 & ~n3900;
  assign n3902 = ~n3896 & ~n3901;
  assign n3903 = ~n3895 & ~n3902;
  assign n3904 = po59  & ~n3903;
  assign n3905 = ~po59  & n3903;
  assign n3906 = ~n3639 & ~n3640;
  assign n3907 = po36  & n3906;
  assign n3908 = ~n3645 & ~n3907;
  assign n3909 = n3645 & n3907;
  assign n3910 = ~n3908 & ~n3909;
  assign n3911 = ~n3905 & ~n3910;
  assign n3912 = ~n3904 & ~n3911;
  assign n3913 = po60  & ~n3912;
  assign n3914 = ~n3648 & ~n3654;
  assign n3915 = po36  & n3914;
  assign n3916 = ~n3653 & ~n3915;
  assign n3917 = n3653 & n3915;
  assign n3918 = ~n3916 & ~n3917;
  assign n3919 = ~po60  & n3912;
  assign n3920 = ~n3918 & ~n3919;
  assign n3921 = ~n3913 & ~n3920;
  assign n3922 = po61  & ~n3921;
  assign n3923 = ~po61  & n3921;
  assign n3924 = ~n3692 & ~n3923;
  assign n3925 = ~n3922 & ~n3924;
  assign n3926 = po62  & ~n3925;
  assign n3927 = ~po62  & n3925;
  assign n3928 = ~n3661 & ~n3662;
  assign n3929 = po36  & n3928;
  assign n3930 = ~n3667 & ~n3929;
  assign n3931 = n3667 & n3929;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = ~n3927 & ~n3932;
  assign n3934 = ~n3926 & ~n3933;
  assign n3935 = n3702 & n3934;
  assign n3936 = ~n3702 & ~n3934;
  assign n3937 = n3680 & po36 ;
  assign n3938 = ~n3679 & ~n3937;
  assign n3939 = n3936 & n3938;
  assign n3940 = ~po63  & ~n3939;
  assign n3941 = ~n3935 & ~n3940;
  assign n3942 = ~n3697 & n3941;
  assign po35  = n3693 | ~n3942;
  assign n3944 = ~n3922 & ~n3923;
  assign n3945 = po35  & n3944;
  assign n3946 = ~n3692 & ~n3945;
  assign n3947 = n3692 & n3945;
  assign n3948 = ~n3946 & ~n3947;
  assign n3949 = n3702 & ~po35 ;
  assign n3950 = ~n3702 & po35 ;
  assign n3951 = n3934 & ~n3950;
  assign n3952 = po63  & ~n3951;
  assign n3953 = ~n3936 & n3952;
  assign n3954 = ~n3926 & ~n3927;
  assign n3955 = po35  & n3954;
  assign n3956 = ~n3932 & ~n3955;
  assign n3957 = n3932 & n3955;
  assign n3958 = ~n3956 & ~n3957;
  assign n3959 = pi70  & po35 ;
  assign n3960 = ~pi68  & ~pi69 ;
  assign n3961 = ~pi70  & n3960;
  assign n3962 = ~n3959 & ~n3961;
  assign n3963 = po36  & ~n3962;
  assign n3964 = ~po36  & n3962;
  assign n3965 = ~pi70  & po35 ;
  assign n3966 = pi71  & ~n3965;
  assign n3967 = n3704 & po35 ;
  assign n3968 = ~n3966 & ~n3967;
  assign n3969 = ~n3964 & n3968;
  assign n3970 = ~n3963 & ~n3969;
  assign n3971 = po37  & ~n3970;
  assign n3972 = ~po37  & n3970;
  assign n3973 = po36  & n3942;
  assign n3974 = ~n3967 & ~n3973;
  assign n3975 = pi72  & ~n3974;
  assign n3976 = ~pi72  & n3974;
  assign n3977 = ~n3975 & ~n3976;
  assign n3978 = ~n3972 & ~n3977;
  assign n3979 = ~n3971 & ~n3978;
  assign n3980 = po38  & ~n3979;
  assign n3981 = ~po38  & n3979;
  assign n3982 = ~n3707 & ~n3708;
  assign n3983 = po35  & n3982;
  assign n3984 = n3712 & ~n3983;
  assign n3985 = ~n3712 & n3983;
  assign n3986 = ~n3984 & ~n3985;
  assign n3987 = ~n3981 & ~n3986;
  assign n3988 = ~n3980 & ~n3987;
  assign n3989 = po39  & ~n3988;
  assign n3990 = ~po39  & n3988;
  assign n3991 = ~n3715 & ~n3716;
  assign n3992 = po35  & n3991;
  assign n3993 = ~n3721 & ~n3992;
  assign n3994 = n3721 & n3992;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = ~n3990 & ~n3995;
  assign n3997 = ~n3989 & ~n3996;
  assign n3998 = po40  & ~n3997;
  assign n3999 = ~po40  & n3997;
  assign n4000 = ~n3724 & ~n3725;
  assign n4001 = po35  & n4000;
  assign n4002 = n3730 & n4001;
  assign n4003 = ~n3730 & ~n4001;
  assign n4004 = ~n4002 & ~n4003;
  assign n4005 = ~n3999 & ~n4004;
  assign n4006 = ~n3998 & ~n4005;
  assign n4007 = po41  & ~n4006;
  assign n4008 = ~po41  & n4006;
  assign n4009 = ~n3733 & ~n3734;
  assign n4010 = po35  & n4009;
  assign n4011 = ~n3739 & ~n4010;
  assign n4012 = n3739 & n4010;
  assign n4013 = ~n4011 & ~n4012;
  assign n4014 = ~n4008 & ~n4013;
  assign n4015 = ~n4007 & ~n4014;
  assign n4016 = po42  & ~n4015;
  assign n4017 = ~po42  & n4015;
  assign n4018 = ~n3742 & ~n3743;
  assign n4019 = po35  & n4018;
  assign n4020 = ~n3748 & ~n4019;
  assign n4021 = n3748 & n4019;
  assign n4022 = ~n4020 & ~n4021;
  assign n4023 = ~n4017 & ~n4022;
  assign n4024 = ~n4016 & ~n4023;
  assign n4025 = po43  & ~n4024;
  assign n4026 = ~po43  & n4024;
  assign n4027 = ~n3751 & ~n3752;
  assign n4028 = po35  & n4027;
  assign n4029 = ~n3757 & ~n4028;
  assign n4030 = n3757 & n4028;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = ~n4026 & ~n4031;
  assign n4033 = ~n4025 & ~n4032;
  assign n4034 = po44  & ~n4033;
  assign n4035 = ~po44  & n4033;
  assign n4036 = ~n3760 & ~n3761;
  assign n4037 = po35  & n4036;
  assign n4038 = ~n3766 & ~n4037;
  assign n4039 = n3766 & n4037;
  assign n4040 = ~n4038 & ~n4039;
  assign n4041 = ~n4035 & ~n4040;
  assign n4042 = ~n4034 & ~n4041;
  assign n4043 = po45  & ~n4042;
  assign n4044 = ~po45  & n4042;
  assign n4045 = ~n3769 & ~n3770;
  assign n4046 = po35  & n4045;
  assign n4047 = ~n3775 & ~n4046;
  assign n4048 = n3775 & n4046;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = ~n4044 & ~n4049;
  assign n4051 = ~n4043 & ~n4050;
  assign n4052 = po46  & ~n4051;
  assign n4053 = ~po46  & n4051;
  assign n4054 = ~n3778 & ~n3779;
  assign n4055 = po35  & n4054;
  assign n4056 = ~n3784 & ~n4055;
  assign n4057 = n3784 & n4055;
  assign n4058 = ~n4056 & ~n4057;
  assign n4059 = ~n4053 & ~n4058;
  assign n4060 = ~n4052 & ~n4059;
  assign n4061 = po47  & ~n4060;
  assign n4062 = ~po47  & n4060;
  assign n4063 = ~n3787 & ~n3788;
  assign n4064 = po35  & n4063;
  assign n4065 = ~n3793 & ~n4064;
  assign n4066 = n3793 & n4064;
  assign n4067 = ~n4065 & ~n4066;
  assign n4068 = ~n4062 & ~n4067;
  assign n4069 = ~n4061 & ~n4068;
  assign n4070 = po48  & ~n4069;
  assign n4071 = ~po48  & n4069;
  assign n4072 = ~n3796 & ~n3797;
  assign n4073 = po35  & n4072;
  assign n4074 = ~n3802 & ~n4073;
  assign n4075 = n3802 & n4073;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = ~n4071 & ~n4076;
  assign n4078 = ~n4070 & ~n4077;
  assign n4079 = po49  & ~n4078;
  assign n4080 = ~po49  & n4078;
  assign n4081 = ~n3805 & ~n3806;
  assign n4082 = po35  & n4081;
  assign n4083 = ~n3811 & ~n4082;
  assign n4084 = n3811 & n4082;
  assign n4085 = ~n4083 & ~n4084;
  assign n4086 = ~n4080 & ~n4085;
  assign n4087 = ~n4079 & ~n4086;
  assign n4088 = po50  & ~n4087;
  assign n4089 = ~po50  & n4087;
  assign n4090 = ~n3814 & ~n3815;
  assign n4091 = po35  & n4090;
  assign n4092 = ~n3820 & ~n4091;
  assign n4093 = n3820 & n4091;
  assign n4094 = ~n4092 & ~n4093;
  assign n4095 = ~n4089 & ~n4094;
  assign n4096 = ~n4088 & ~n4095;
  assign n4097 = po51  & ~n4096;
  assign n4098 = ~po51  & n4096;
  assign n4099 = ~n3823 & ~n3824;
  assign n4100 = po35  & n4099;
  assign n4101 = ~n3829 & ~n4100;
  assign n4102 = n3829 & n4100;
  assign n4103 = ~n4101 & ~n4102;
  assign n4104 = ~n4098 & ~n4103;
  assign n4105 = ~n4097 & ~n4104;
  assign n4106 = po52  & ~n4105;
  assign n4107 = ~po52  & n4105;
  assign n4108 = ~n3832 & ~n3833;
  assign n4109 = po35  & n4108;
  assign n4110 = ~n3838 & ~n4109;
  assign n4111 = n3838 & n4109;
  assign n4112 = ~n4110 & ~n4111;
  assign n4113 = ~n4107 & ~n4112;
  assign n4114 = ~n4106 & ~n4113;
  assign n4115 = po53  & ~n4114;
  assign n4116 = ~po53  & n4114;
  assign n4117 = ~n3841 & ~n3842;
  assign n4118 = po35  & n4117;
  assign n4119 = ~n3847 & ~n4118;
  assign n4120 = n3847 & n4118;
  assign n4121 = ~n4119 & ~n4120;
  assign n4122 = ~n4116 & ~n4121;
  assign n4123 = ~n4115 & ~n4122;
  assign n4124 = po54  & ~n4123;
  assign n4125 = ~po54  & n4123;
  assign n4126 = ~n3850 & ~n3851;
  assign n4127 = po35  & n4126;
  assign n4128 = ~n3856 & ~n4127;
  assign n4129 = n3856 & n4127;
  assign n4130 = ~n4128 & ~n4129;
  assign n4131 = ~n4125 & ~n4130;
  assign n4132 = ~n4124 & ~n4131;
  assign n4133 = po55  & ~n4132;
  assign n4134 = ~po55  & n4132;
  assign n4135 = ~n3859 & ~n3860;
  assign n4136 = po35  & n4135;
  assign n4137 = ~n3865 & ~n4136;
  assign n4138 = n3865 & n4136;
  assign n4139 = ~n4137 & ~n4138;
  assign n4140 = ~n4134 & ~n4139;
  assign n4141 = ~n4133 & ~n4140;
  assign n4142 = po56  & ~n4141;
  assign n4143 = ~po56  & n4141;
  assign n4144 = ~n3868 & ~n3869;
  assign n4145 = po35  & n4144;
  assign n4146 = ~n3874 & ~n4145;
  assign n4147 = n3874 & n4145;
  assign n4148 = ~n4146 & ~n4147;
  assign n4149 = ~n4143 & ~n4148;
  assign n4150 = ~n4142 & ~n4149;
  assign n4151 = po57  & ~n4150;
  assign n4152 = ~po57  & n4150;
  assign n4153 = ~n3877 & ~n3878;
  assign n4154 = po35  & n4153;
  assign n4155 = ~n3883 & ~n4154;
  assign n4156 = n3883 & n4154;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~n4152 & ~n4157;
  assign n4159 = ~n4151 & ~n4158;
  assign n4160 = po58  & ~n4159;
  assign n4161 = ~po58  & n4159;
  assign n4162 = ~n3886 & ~n3887;
  assign n4163 = po35  & n4162;
  assign n4164 = ~n3892 & ~n4163;
  assign n4165 = n3892 & n4163;
  assign n4166 = ~n4164 & ~n4165;
  assign n4167 = ~n4161 & ~n4166;
  assign n4168 = ~n4160 & ~n4167;
  assign n4169 = po59  & ~n4168;
  assign n4170 = ~po59  & n4168;
  assign n4171 = ~n3895 & ~n3896;
  assign n4172 = po35  & n4171;
  assign n4173 = ~n3901 & ~n4172;
  assign n4174 = n3901 & n4172;
  assign n4175 = ~n4173 & ~n4174;
  assign n4176 = ~n4170 & ~n4175;
  assign n4177 = ~n4169 & ~n4176;
  assign n4178 = po60  & ~n4177;
  assign n4179 = ~po60  & n4177;
  assign n4180 = ~n3904 & ~n3905;
  assign n4181 = po35  & n4180;
  assign n4182 = ~n3910 & ~n4181;
  assign n4183 = n3910 & n4181;
  assign n4184 = ~n4182 & ~n4183;
  assign n4185 = ~n4179 & ~n4184;
  assign n4186 = ~n4178 & ~n4185;
  assign n4187 = po61  & ~n4186;
  assign n4188 = ~n3913 & ~n3919;
  assign n4189 = po35  & n4188;
  assign n4190 = ~n3918 & ~n4189;
  assign n4191 = n3918 & n4189;
  assign n4192 = ~n4190 & ~n4191;
  assign n4193 = ~po61  & n4186;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = ~n4187 & ~n4194;
  assign n4196 = po62  & ~n4195;
  assign n4197 = ~po62  & n4195;
  assign n4198 = ~n3948 & ~n4197;
  assign n4199 = ~n4196 & ~n4198;
  assign n4200 = n3958 & n4199;
  assign n4201 = ~n3958 & ~n4199;
  assign n4202 = n3936 & po35 ;
  assign n4203 = ~n3935 & ~n4202;
  assign n4204 = n4201 & n4203;
  assign n4205 = ~po63  & ~n4204;
  assign n4206 = ~n4200 & ~n4205;
  assign n4207 = ~n3953 & n4206;
  assign po34  = n3949 | ~n4207;
  assign n4209 = ~n4196 & ~n4197;
  assign n4210 = po34  & n4209;
  assign n4211 = ~n3948 & ~n4210;
  assign n4212 = n3948 & n4210;
  assign n4213 = ~n4211 & ~n4212;
  assign n4214 = n3958 & ~po34 ;
  assign n4215 = ~n3958 & po34 ;
  assign n4216 = n4199 & ~n4215;
  assign n4217 = po63  & ~n4216;
  assign n4218 = ~n4201 & n4217;
  assign n4219 = pi68  & po34 ;
  assign n4220 = ~pi66  & ~pi67 ;
  assign n4221 = ~pi68  & n4220;
  assign n4222 = ~n4219 & ~n4221;
  assign n4223 = po35  & ~n4222;
  assign n4224 = ~po35  & n4222;
  assign n4225 = ~pi68  & po34 ;
  assign n4226 = pi69  & ~n4225;
  assign n4227 = n3960 & po34 ;
  assign n4228 = ~n4226 & ~n4227;
  assign n4229 = ~n4224 & n4228;
  assign n4230 = ~n4223 & ~n4229;
  assign n4231 = po36  & ~n4230;
  assign n4232 = ~po36  & n4230;
  assign n4233 = po35  & n4207;
  assign n4234 = ~n4227 & ~n4233;
  assign n4235 = pi70  & ~n4234;
  assign n4236 = ~pi70  & n4234;
  assign n4237 = ~n4235 & ~n4236;
  assign n4238 = ~n4232 & ~n4237;
  assign n4239 = ~n4231 & ~n4238;
  assign n4240 = po37  & ~n4239;
  assign n4241 = ~po37  & n4239;
  assign n4242 = ~n3963 & ~n3964;
  assign n4243 = po34  & n4242;
  assign n4244 = n3968 & ~n4243;
  assign n4245 = ~n3968 & n4243;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = ~n4241 & ~n4246;
  assign n4248 = ~n4240 & ~n4247;
  assign n4249 = po38  & ~n4248;
  assign n4250 = ~po38  & n4248;
  assign n4251 = ~n3971 & ~n3972;
  assign n4252 = po34  & n4251;
  assign n4253 = ~n3977 & ~n4252;
  assign n4254 = n3977 & n4252;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = ~n4250 & ~n4255;
  assign n4257 = ~n4249 & ~n4256;
  assign n4258 = po39  & ~n4257;
  assign n4259 = ~po39  & n4257;
  assign n4260 = ~n3980 & ~n3981;
  assign n4261 = po34  & n4260;
  assign n4262 = n3986 & n4261;
  assign n4263 = ~n3986 & ~n4261;
  assign n4264 = ~n4262 & ~n4263;
  assign n4265 = ~n4259 & ~n4264;
  assign n4266 = ~n4258 & ~n4265;
  assign n4267 = po40  & ~n4266;
  assign n4268 = ~po40  & n4266;
  assign n4269 = ~n3989 & ~n3990;
  assign n4270 = po34  & n4269;
  assign n4271 = ~n3995 & ~n4270;
  assign n4272 = n3995 & n4270;
  assign n4273 = ~n4271 & ~n4272;
  assign n4274 = ~n4268 & ~n4273;
  assign n4275 = ~n4267 & ~n4274;
  assign n4276 = po41  & ~n4275;
  assign n4277 = ~po41  & n4275;
  assign n4278 = ~n3998 & ~n3999;
  assign n4279 = po34  & n4278;
  assign n4280 = ~n4004 & ~n4279;
  assign n4281 = n4004 & n4279;
  assign n4282 = ~n4280 & ~n4281;
  assign n4283 = ~n4277 & ~n4282;
  assign n4284 = ~n4276 & ~n4283;
  assign n4285 = po42  & ~n4284;
  assign n4286 = ~po42  & n4284;
  assign n4287 = ~n4007 & ~n4008;
  assign n4288 = po34  & n4287;
  assign n4289 = ~n4013 & ~n4288;
  assign n4290 = n4013 & n4288;
  assign n4291 = ~n4289 & ~n4290;
  assign n4292 = ~n4286 & ~n4291;
  assign n4293 = ~n4285 & ~n4292;
  assign n4294 = po43  & ~n4293;
  assign n4295 = ~po43  & n4293;
  assign n4296 = ~n4016 & ~n4017;
  assign n4297 = po34  & n4296;
  assign n4298 = ~n4022 & ~n4297;
  assign n4299 = n4022 & n4297;
  assign n4300 = ~n4298 & ~n4299;
  assign n4301 = ~n4295 & ~n4300;
  assign n4302 = ~n4294 & ~n4301;
  assign n4303 = po44  & ~n4302;
  assign n4304 = ~po44  & n4302;
  assign n4305 = ~n4025 & ~n4026;
  assign n4306 = po34  & n4305;
  assign n4307 = ~n4031 & ~n4306;
  assign n4308 = n4031 & n4306;
  assign n4309 = ~n4307 & ~n4308;
  assign n4310 = ~n4304 & ~n4309;
  assign n4311 = ~n4303 & ~n4310;
  assign n4312 = po45  & ~n4311;
  assign n4313 = ~po45  & n4311;
  assign n4314 = ~n4034 & ~n4035;
  assign n4315 = po34  & n4314;
  assign n4316 = ~n4040 & ~n4315;
  assign n4317 = n4040 & n4315;
  assign n4318 = ~n4316 & ~n4317;
  assign n4319 = ~n4313 & ~n4318;
  assign n4320 = ~n4312 & ~n4319;
  assign n4321 = po46  & ~n4320;
  assign n4322 = ~po46  & n4320;
  assign n4323 = ~n4043 & ~n4044;
  assign n4324 = po34  & n4323;
  assign n4325 = ~n4049 & ~n4324;
  assign n4326 = n4049 & n4324;
  assign n4327 = ~n4325 & ~n4326;
  assign n4328 = ~n4322 & ~n4327;
  assign n4329 = ~n4321 & ~n4328;
  assign n4330 = po47  & ~n4329;
  assign n4331 = ~po47  & n4329;
  assign n4332 = ~n4052 & ~n4053;
  assign n4333 = po34  & n4332;
  assign n4334 = ~n4058 & ~n4333;
  assign n4335 = n4058 & n4333;
  assign n4336 = ~n4334 & ~n4335;
  assign n4337 = ~n4331 & ~n4336;
  assign n4338 = ~n4330 & ~n4337;
  assign n4339 = po48  & ~n4338;
  assign n4340 = ~po48  & n4338;
  assign n4341 = ~n4061 & ~n4062;
  assign n4342 = po34  & n4341;
  assign n4343 = ~n4067 & ~n4342;
  assign n4344 = n4067 & n4342;
  assign n4345 = ~n4343 & ~n4344;
  assign n4346 = ~n4340 & ~n4345;
  assign n4347 = ~n4339 & ~n4346;
  assign n4348 = po49  & ~n4347;
  assign n4349 = ~po49  & n4347;
  assign n4350 = ~n4070 & ~n4071;
  assign n4351 = po34  & n4350;
  assign n4352 = ~n4076 & ~n4351;
  assign n4353 = n4076 & n4351;
  assign n4354 = ~n4352 & ~n4353;
  assign n4355 = ~n4349 & ~n4354;
  assign n4356 = ~n4348 & ~n4355;
  assign n4357 = po50  & ~n4356;
  assign n4358 = ~po50  & n4356;
  assign n4359 = ~n4079 & ~n4080;
  assign n4360 = po34  & n4359;
  assign n4361 = ~n4085 & ~n4360;
  assign n4362 = n4085 & n4360;
  assign n4363 = ~n4361 & ~n4362;
  assign n4364 = ~n4358 & ~n4363;
  assign n4365 = ~n4357 & ~n4364;
  assign n4366 = po51  & ~n4365;
  assign n4367 = ~po51  & n4365;
  assign n4368 = ~n4088 & ~n4089;
  assign n4369 = po34  & n4368;
  assign n4370 = ~n4094 & ~n4369;
  assign n4371 = n4094 & n4369;
  assign n4372 = ~n4370 & ~n4371;
  assign n4373 = ~n4367 & ~n4372;
  assign n4374 = ~n4366 & ~n4373;
  assign n4375 = po52  & ~n4374;
  assign n4376 = ~po52  & n4374;
  assign n4377 = ~n4097 & ~n4098;
  assign n4378 = po34  & n4377;
  assign n4379 = ~n4103 & ~n4378;
  assign n4380 = n4103 & n4378;
  assign n4381 = ~n4379 & ~n4380;
  assign n4382 = ~n4376 & ~n4381;
  assign n4383 = ~n4375 & ~n4382;
  assign n4384 = po53  & ~n4383;
  assign n4385 = ~po53  & n4383;
  assign n4386 = ~n4106 & ~n4107;
  assign n4387 = po34  & n4386;
  assign n4388 = ~n4112 & ~n4387;
  assign n4389 = n4112 & n4387;
  assign n4390 = ~n4388 & ~n4389;
  assign n4391 = ~n4385 & ~n4390;
  assign n4392 = ~n4384 & ~n4391;
  assign n4393 = po54  & ~n4392;
  assign n4394 = ~po54  & n4392;
  assign n4395 = ~n4115 & ~n4116;
  assign n4396 = po34  & n4395;
  assign n4397 = ~n4121 & ~n4396;
  assign n4398 = n4121 & n4396;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n4394 & ~n4399;
  assign n4401 = ~n4393 & ~n4400;
  assign n4402 = po55  & ~n4401;
  assign n4403 = ~po55  & n4401;
  assign n4404 = ~n4124 & ~n4125;
  assign n4405 = po34  & n4404;
  assign n4406 = ~n4130 & ~n4405;
  assign n4407 = n4130 & n4405;
  assign n4408 = ~n4406 & ~n4407;
  assign n4409 = ~n4403 & ~n4408;
  assign n4410 = ~n4402 & ~n4409;
  assign n4411 = po56  & ~n4410;
  assign n4412 = ~po56  & n4410;
  assign n4413 = ~n4133 & ~n4134;
  assign n4414 = po34  & n4413;
  assign n4415 = ~n4139 & ~n4414;
  assign n4416 = n4139 & n4414;
  assign n4417 = ~n4415 & ~n4416;
  assign n4418 = ~n4412 & ~n4417;
  assign n4419 = ~n4411 & ~n4418;
  assign n4420 = po57  & ~n4419;
  assign n4421 = ~po57  & n4419;
  assign n4422 = ~n4142 & ~n4143;
  assign n4423 = po34  & n4422;
  assign n4424 = ~n4148 & ~n4423;
  assign n4425 = n4148 & n4423;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = ~n4421 & ~n4426;
  assign n4428 = ~n4420 & ~n4427;
  assign n4429 = po58  & ~n4428;
  assign n4430 = ~po58  & n4428;
  assign n4431 = ~n4151 & ~n4152;
  assign n4432 = po34  & n4431;
  assign n4433 = ~n4157 & ~n4432;
  assign n4434 = n4157 & n4432;
  assign n4435 = ~n4433 & ~n4434;
  assign n4436 = ~n4430 & ~n4435;
  assign n4437 = ~n4429 & ~n4436;
  assign n4438 = po59  & ~n4437;
  assign n4439 = ~po59  & n4437;
  assign n4440 = ~n4160 & ~n4161;
  assign n4441 = po34  & n4440;
  assign n4442 = ~n4166 & ~n4441;
  assign n4443 = n4166 & n4441;
  assign n4444 = ~n4442 & ~n4443;
  assign n4445 = ~n4439 & ~n4444;
  assign n4446 = ~n4438 & ~n4445;
  assign n4447 = po60  & ~n4446;
  assign n4448 = ~po60  & n4446;
  assign n4449 = ~n4169 & ~n4170;
  assign n4450 = po34  & n4449;
  assign n4451 = ~n4175 & ~n4450;
  assign n4452 = n4175 & n4450;
  assign n4453 = ~n4451 & ~n4452;
  assign n4454 = ~n4448 & ~n4453;
  assign n4455 = ~n4447 & ~n4454;
  assign n4456 = po61  & ~n4455;
  assign n4457 = ~po61  & n4455;
  assign n4458 = ~n4178 & ~n4179;
  assign n4459 = po34  & n4458;
  assign n4460 = ~n4184 & ~n4459;
  assign n4461 = n4184 & n4459;
  assign n4462 = ~n4460 & ~n4461;
  assign n4463 = ~n4457 & ~n4462;
  assign n4464 = ~n4456 & ~n4463;
  assign n4465 = po62  & ~n4464;
  assign n4466 = ~n4187 & ~n4193;
  assign n4467 = po34  & n4466;
  assign n4468 = ~n4192 & ~n4467;
  assign n4469 = n4192 & n4467;
  assign n4470 = ~n4468 & ~n4469;
  assign n4471 = ~po62  & n4464;
  assign n4472 = ~n4470 & ~n4471;
  assign n4473 = ~n4465 & ~n4472;
  assign n4474 = n4213 & n4473;
  assign n4475 = ~n4213 & ~n4473;
  assign n4476 = n4201 & po34 ;
  assign n4477 = ~n4200 & ~n4476;
  assign n4478 = n4475 & n4477;
  assign n4479 = ~po63  & ~n4478;
  assign n4480 = ~n4474 & ~n4479;
  assign n4481 = ~n4218 & n4480;
  assign po33  = n4214 | ~n4481;
  assign n4483 = n4213 & ~po33 ;
  assign n4484 = ~n4213 & po33 ;
  assign n4485 = n4473 & ~n4484;
  assign n4486 = po63  & ~n4485;
  assign n4487 = ~n4475 & n4486;
  assign n4488 = ~n4465 & ~n4471;
  assign n4489 = po33  & n4488;
  assign n4490 = ~n4470 & ~n4489;
  assign n4491 = n4470 & n4489;
  assign n4492 = ~n4490 & ~n4491;
  assign n4493 = pi66  & po33 ;
  assign n4494 = ~pi64  & ~pi65 ;
  assign n4495 = ~pi66  & n4494;
  assign n4496 = ~n4493 & ~n4495;
  assign n4497 = po34  & ~n4496;
  assign n4498 = ~po34  & n4496;
  assign n4499 = ~pi66  & po33 ;
  assign n4500 = pi67  & ~n4499;
  assign n4501 = n4220 & po33 ;
  assign n4502 = ~n4500 & ~n4501;
  assign n4503 = ~n4498 & n4502;
  assign n4504 = ~n4497 & ~n4503;
  assign n4505 = po35  & ~n4504;
  assign n4506 = ~po35  & n4504;
  assign n4507 = po34  & n4481;
  assign n4508 = ~n4501 & ~n4507;
  assign n4509 = pi68  & ~n4508;
  assign n4510 = ~pi68  & n4508;
  assign n4511 = ~n4509 & ~n4510;
  assign n4512 = ~n4506 & ~n4511;
  assign n4513 = ~n4505 & ~n4512;
  assign n4514 = po36  & ~n4513;
  assign n4515 = ~po36  & n4513;
  assign n4516 = ~n4223 & ~n4224;
  assign n4517 = po33  & n4516;
  assign n4518 = n4228 & ~n4517;
  assign n4519 = ~n4228 & n4517;
  assign n4520 = ~n4518 & ~n4519;
  assign n4521 = ~n4515 & ~n4520;
  assign n4522 = ~n4514 & ~n4521;
  assign n4523 = po37  & ~n4522;
  assign n4524 = ~po37  & n4522;
  assign n4525 = ~n4231 & ~n4232;
  assign n4526 = po33  & n4525;
  assign n4527 = ~n4237 & ~n4526;
  assign n4528 = n4237 & n4526;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = ~n4524 & ~n4529;
  assign n4531 = ~n4523 & ~n4530;
  assign n4532 = po38  & ~n4531;
  assign n4533 = ~po38  & n4531;
  assign n4534 = ~n4240 & ~n4241;
  assign n4535 = po33  & n4534;
  assign n4536 = n4246 & n4535;
  assign n4537 = ~n4246 & ~n4535;
  assign n4538 = ~n4536 & ~n4537;
  assign n4539 = ~n4533 & ~n4538;
  assign n4540 = ~n4532 & ~n4539;
  assign n4541 = po39  & ~n4540;
  assign n4542 = ~po39  & n4540;
  assign n4543 = ~n4249 & ~n4250;
  assign n4544 = po33  & n4543;
  assign n4545 = ~n4255 & ~n4544;
  assign n4546 = n4255 & n4544;
  assign n4547 = ~n4545 & ~n4546;
  assign n4548 = ~n4542 & ~n4547;
  assign n4549 = ~n4541 & ~n4548;
  assign n4550 = po40  & ~n4549;
  assign n4551 = ~po40  & n4549;
  assign n4552 = ~n4258 & ~n4259;
  assign n4553 = po33  & n4552;
  assign n4554 = ~n4264 & ~n4553;
  assign n4555 = n4264 & n4553;
  assign n4556 = ~n4554 & ~n4555;
  assign n4557 = ~n4551 & ~n4556;
  assign n4558 = ~n4550 & ~n4557;
  assign n4559 = po41  & ~n4558;
  assign n4560 = ~po41  & n4558;
  assign n4561 = ~n4267 & ~n4268;
  assign n4562 = po33  & n4561;
  assign n4563 = ~n4273 & ~n4562;
  assign n4564 = n4273 & n4562;
  assign n4565 = ~n4563 & ~n4564;
  assign n4566 = ~n4560 & ~n4565;
  assign n4567 = ~n4559 & ~n4566;
  assign n4568 = po42  & ~n4567;
  assign n4569 = ~po42  & n4567;
  assign n4570 = ~n4276 & ~n4277;
  assign n4571 = po33  & n4570;
  assign n4572 = ~n4282 & ~n4571;
  assign n4573 = n4282 & n4571;
  assign n4574 = ~n4572 & ~n4573;
  assign n4575 = ~n4569 & ~n4574;
  assign n4576 = ~n4568 & ~n4575;
  assign n4577 = po43  & ~n4576;
  assign n4578 = ~po43  & n4576;
  assign n4579 = ~n4285 & ~n4286;
  assign n4580 = po33  & n4579;
  assign n4581 = ~n4291 & ~n4580;
  assign n4582 = n4291 & n4580;
  assign n4583 = ~n4581 & ~n4582;
  assign n4584 = ~n4578 & ~n4583;
  assign n4585 = ~n4577 & ~n4584;
  assign n4586 = po44  & ~n4585;
  assign n4587 = ~po44  & n4585;
  assign n4588 = ~n4294 & ~n4295;
  assign n4589 = po33  & n4588;
  assign n4590 = ~n4300 & ~n4589;
  assign n4591 = n4300 & n4589;
  assign n4592 = ~n4590 & ~n4591;
  assign n4593 = ~n4587 & ~n4592;
  assign n4594 = ~n4586 & ~n4593;
  assign n4595 = po45  & ~n4594;
  assign n4596 = ~po45  & n4594;
  assign n4597 = ~n4303 & ~n4304;
  assign n4598 = po33  & n4597;
  assign n4599 = ~n4309 & ~n4598;
  assign n4600 = n4309 & n4598;
  assign n4601 = ~n4599 & ~n4600;
  assign n4602 = ~n4596 & ~n4601;
  assign n4603 = ~n4595 & ~n4602;
  assign n4604 = po46  & ~n4603;
  assign n4605 = ~po46  & n4603;
  assign n4606 = ~n4312 & ~n4313;
  assign n4607 = po33  & n4606;
  assign n4608 = ~n4318 & ~n4607;
  assign n4609 = n4318 & n4607;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = ~n4605 & ~n4610;
  assign n4612 = ~n4604 & ~n4611;
  assign n4613 = po47  & ~n4612;
  assign n4614 = ~po47  & n4612;
  assign n4615 = ~n4321 & ~n4322;
  assign n4616 = po33  & n4615;
  assign n4617 = ~n4327 & ~n4616;
  assign n4618 = n4327 & n4616;
  assign n4619 = ~n4617 & ~n4618;
  assign n4620 = ~n4614 & ~n4619;
  assign n4621 = ~n4613 & ~n4620;
  assign n4622 = po48  & ~n4621;
  assign n4623 = ~po48  & n4621;
  assign n4624 = ~n4330 & ~n4331;
  assign n4625 = po33  & n4624;
  assign n4626 = ~n4336 & ~n4625;
  assign n4627 = n4336 & n4625;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = ~n4623 & ~n4628;
  assign n4630 = ~n4622 & ~n4629;
  assign n4631 = po49  & ~n4630;
  assign n4632 = ~po49  & n4630;
  assign n4633 = ~n4339 & ~n4340;
  assign n4634 = po33  & n4633;
  assign n4635 = ~n4345 & ~n4634;
  assign n4636 = n4345 & n4634;
  assign n4637 = ~n4635 & ~n4636;
  assign n4638 = ~n4632 & ~n4637;
  assign n4639 = ~n4631 & ~n4638;
  assign n4640 = po50  & ~n4639;
  assign n4641 = ~po50  & n4639;
  assign n4642 = ~n4348 & ~n4349;
  assign n4643 = po33  & n4642;
  assign n4644 = ~n4354 & ~n4643;
  assign n4645 = n4354 & n4643;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = ~n4641 & ~n4646;
  assign n4648 = ~n4640 & ~n4647;
  assign n4649 = po51  & ~n4648;
  assign n4650 = ~po51  & n4648;
  assign n4651 = ~n4357 & ~n4358;
  assign n4652 = po33  & n4651;
  assign n4653 = ~n4363 & ~n4652;
  assign n4654 = n4363 & n4652;
  assign n4655 = ~n4653 & ~n4654;
  assign n4656 = ~n4650 & ~n4655;
  assign n4657 = ~n4649 & ~n4656;
  assign n4658 = po52  & ~n4657;
  assign n4659 = ~po52  & n4657;
  assign n4660 = ~n4366 & ~n4367;
  assign n4661 = po33  & n4660;
  assign n4662 = ~n4372 & ~n4661;
  assign n4663 = n4372 & n4661;
  assign n4664 = ~n4662 & ~n4663;
  assign n4665 = ~n4659 & ~n4664;
  assign n4666 = ~n4658 & ~n4665;
  assign n4667 = po53  & ~n4666;
  assign n4668 = ~po53  & n4666;
  assign n4669 = ~n4375 & ~n4376;
  assign n4670 = po33  & n4669;
  assign n4671 = ~n4381 & ~n4670;
  assign n4672 = n4381 & n4670;
  assign n4673 = ~n4671 & ~n4672;
  assign n4674 = ~n4668 & ~n4673;
  assign n4675 = ~n4667 & ~n4674;
  assign n4676 = po54  & ~n4675;
  assign n4677 = ~po54  & n4675;
  assign n4678 = ~n4384 & ~n4385;
  assign n4679 = po33  & n4678;
  assign n4680 = ~n4390 & ~n4679;
  assign n4681 = n4390 & n4679;
  assign n4682 = ~n4680 & ~n4681;
  assign n4683 = ~n4677 & ~n4682;
  assign n4684 = ~n4676 & ~n4683;
  assign n4685 = po55  & ~n4684;
  assign n4686 = ~po55  & n4684;
  assign n4687 = ~n4393 & ~n4394;
  assign n4688 = po33  & n4687;
  assign n4689 = ~n4399 & ~n4688;
  assign n4690 = n4399 & n4688;
  assign n4691 = ~n4689 & ~n4690;
  assign n4692 = ~n4686 & ~n4691;
  assign n4693 = ~n4685 & ~n4692;
  assign n4694 = po56  & ~n4693;
  assign n4695 = ~po56  & n4693;
  assign n4696 = ~n4402 & ~n4403;
  assign n4697 = po33  & n4696;
  assign n4698 = ~n4408 & ~n4697;
  assign n4699 = n4408 & n4697;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = ~n4695 & ~n4700;
  assign n4702 = ~n4694 & ~n4701;
  assign n4703 = po57  & ~n4702;
  assign n4704 = ~po57  & n4702;
  assign n4705 = ~n4411 & ~n4412;
  assign n4706 = po33  & n4705;
  assign n4707 = ~n4417 & ~n4706;
  assign n4708 = n4417 & n4706;
  assign n4709 = ~n4707 & ~n4708;
  assign n4710 = ~n4704 & ~n4709;
  assign n4711 = ~n4703 & ~n4710;
  assign n4712 = po58  & ~n4711;
  assign n4713 = ~po58  & n4711;
  assign n4714 = ~n4420 & ~n4421;
  assign n4715 = po33  & n4714;
  assign n4716 = ~n4426 & ~n4715;
  assign n4717 = n4426 & n4715;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = ~n4713 & ~n4718;
  assign n4720 = ~n4712 & ~n4719;
  assign n4721 = po59  & ~n4720;
  assign n4722 = ~po59  & n4720;
  assign n4723 = ~n4429 & ~n4430;
  assign n4724 = po33  & n4723;
  assign n4725 = ~n4435 & ~n4724;
  assign n4726 = n4435 & n4724;
  assign n4727 = ~n4725 & ~n4726;
  assign n4728 = ~n4722 & ~n4727;
  assign n4729 = ~n4721 & ~n4728;
  assign n4730 = po60  & ~n4729;
  assign n4731 = ~po60  & n4729;
  assign n4732 = ~n4438 & ~n4439;
  assign n4733 = po33  & n4732;
  assign n4734 = ~n4444 & ~n4733;
  assign n4735 = n4444 & n4733;
  assign n4736 = ~n4734 & ~n4735;
  assign n4737 = ~n4731 & ~n4736;
  assign n4738 = ~n4730 & ~n4737;
  assign n4739 = po61  & ~n4738;
  assign n4740 = ~po61  & n4738;
  assign n4741 = ~n4447 & ~n4448;
  assign n4742 = po33  & n4741;
  assign n4743 = ~n4453 & ~n4742;
  assign n4744 = n4453 & n4742;
  assign n4745 = ~n4743 & ~n4744;
  assign n4746 = ~n4740 & ~n4745;
  assign n4747 = ~n4739 & ~n4746;
  assign n4748 = po62  & ~n4747;
  assign n4749 = ~po62  & n4747;
  assign n4750 = ~n4456 & ~n4457;
  assign n4751 = po33  & n4750;
  assign n4752 = ~n4462 & ~n4751;
  assign n4753 = n4462 & n4751;
  assign n4754 = ~n4752 & ~n4753;
  assign n4755 = ~n4749 & ~n4754;
  assign n4756 = ~n4748 & ~n4755;
  assign n4757 = n4492 & n4756;
  assign n4758 = ~n4492 & ~n4756;
  assign n4759 = n4475 & po33 ;
  assign n4760 = ~n4474 & ~n4759;
  assign n4761 = n4758 & n4760;
  assign n4762 = ~po63  & ~n4761;
  assign n4763 = ~n4757 & ~n4762;
  assign n4764 = ~n4487 & n4763;
  assign po32  = n4483 | ~n4764;
  assign n4766 = ~pi64  & po32 ;
  assign n4767 = pi65  & ~n4766;
  assign n4768 = n4494 & po32 ;
  assign n4769 = ~n4767 & ~n4768;
  assign n4770 = n4492 & ~po32 ;
  assign n4771 = ~n4492 & po32 ;
  assign n4772 = n4756 & ~n4771;
  assign n4773 = po63  & ~n4772;
  assign n4774 = ~n4758 & n4773;
  assign n4775 = ~n4748 & ~n4749;
  assign n4776 = po32  & n4775;
  assign n4777 = ~n4754 & ~n4776;
  assign n4778 = n4754 & n4776;
  assign n4779 = ~n4777 & ~n4778;
  assign n4780 = pi64  & po32 ;
  assign n4781 = ~pi62  & ~pi63 ;
  assign n4782 = ~pi64  & n4781;
  assign n4783 = ~n4780 & ~n4782;
  assign n4784 = po33  & ~n4783;
  assign n4785 = ~po33  & n4783;
  assign n4786 = n4769 & ~n4785;
  assign n4787 = ~n4784 & ~n4786;
  assign n4788 = po34  & ~n4787;
  assign n4789 = ~po34  & n4787;
  assign n4790 = po33  & n4764;
  assign n4791 = ~n4768 & ~n4790;
  assign n4792 = pi66  & ~n4791;
  assign n4793 = ~pi66  & n4791;
  assign n4794 = ~n4792 & ~n4793;
  assign n4795 = ~n4789 & ~n4794;
  assign n4796 = ~n4788 & ~n4795;
  assign n4797 = po35  & ~n4796;
  assign n4798 = ~po35  & n4796;
  assign n4799 = ~n4497 & ~n4498;
  assign n4800 = po32  & n4799;
  assign n4801 = n4502 & ~n4800;
  assign n4802 = ~n4502 & n4800;
  assign n4803 = ~n4801 & ~n4802;
  assign n4804 = ~n4798 & ~n4803;
  assign n4805 = ~n4797 & ~n4804;
  assign n4806 = po36  & ~n4805;
  assign n4807 = ~po36  & n4805;
  assign n4808 = ~n4505 & ~n4506;
  assign n4809 = po32  & n4808;
  assign n4810 = ~n4511 & ~n4809;
  assign n4811 = n4511 & n4809;
  assign n4812 = ~n4810 & ~n4811;
  assign n4813 = ~n4807 & ~n4812;
  assign n4814 = ~n4806 & ~n4813;
  assign n4815 = po37  & ~n4814;
  assign n4816 = ~po37  & n4814;
  assign n4817 = ~n4514 & ~n4515;
  assign n4818 = po32  & n4817;
  assign n4819 = n4520 & n4818;
  assign n4820 = ~n4520 & ~n4818;
  assign n4821 = ~n4819 & ~n4820;
  assign n4822 = ~n4816 & ~n4821;
  assign n4823 = ~n4815 & ~n4822;
  assign n4824 = po38  & ~n4823;
  assign n4825 = ~po38  & n4823;
  assign n4826 = ~n4523 & ~n4524;
  assign n4827 = po32  & n4826;
  assign n4828 = ~n4529 & ~n4827;
  assign n4829 = n4529 & n4827;
  assign n4830 = ~n4828 & ~n4829;
  assign n4831 = ~n4825 & ~n4830;
  assign n4832 = ~n4824 & ~n4831;
  assign n4833 = po39  & ~n4832;
  assign n4834 = ~po39  & n4832;
  assign n4835 = ~n4532 & ~n4533;
  assign n4836 = po32  & n4835;
  assign n4837 = ~n4538 & ~n4836;
  assign n4838 = n4538 & n4836;
  assign n4839 = ~n4837 & ~n4838;
  assign n4840 = ~n4834 & ~n4839;
  assign n4841 = ~n4833 & ~n4840;
  assign n4842 = po40  & ~n4841;
  assign n4843 = ~po40  & n4841;
  assign n4844 = ~n4541 & ~n4542;
  assign n4845 = po32  & n4844;
  assign n4846 = ~n4547 & ~n4845;
  assign n4847 = n4547 & n4845;
  assign n4848 = ~n4846 & ~n4847;
  assign n4849 = ~n4843 & ~n4848;
  assign n4850 = ~n4842 & ~n4849;
  assign n4851 = po41  & ~n4850;
  assign n4852 = ~po41  & n4850;
  assign n4853 = ~n4550 & ~n4551;
  assign n4854 = po32  & n4853;
  assign n4855 = ~n4556 & ~n4854;
  assign n4856 = n4556 & n4854;
  assign n4857 = ~n4855 & ~n4856;
  assign n4858 = ~n4852 & ~n4857;
  assign n4859 = ~n4851 & ~n4858;
  assign n4860 = po42  & ~n4859;
  assign n4861 = ~po42  & n4859;
  assign n4862 = ~n4559 & ~n4560;
  assign n4863 = po32  & n4862;
  assign n4864 = ~n4565 & ~n4863;
  assign n4865 = n4565 & n4863;
  assign n4866 = ~n4864 & ~n4865;
  assign n4867 = ~n4861 & ~n4866;
  assign n4868 = ~n4860 & ~n4867;
  assign n4869 = po43  & ~n4868;
  assign n4870 = ~po43  & n4868;
  assign n4871 = ~n4568 & ~n4569;
  assign n4872 = po32  & n4871;
  assign n4873 = ~n4574 & ~n4872;
  assign n4874 = n4574 & n4872;
  assign n4875 = ~n4873 & ~n4874;
  assign n4876 = ~n4870 & ~n4875;
  assign n4877 = ~n4869 & ~n4876;
  assign n4878 = po44  & ~n4877;
  assign n4879 = ~po44  & n4877;
  assign n4880 = ~n4577 & ~n4578;
  assign n4881 = po32  & n4880;
  assign n4882 = ~n4583 & ~n4881;
  assign n4883 = n4583 & n4881;
  assign n4884 = ~n4882 & ~n4883;
  assign n4885 = ~n4879 & ~n4884;
  assign n4886 = ~n4878 & ~n4885;
  assign n4887 = po45  & ~n4886;
  assign n4888 = ~po45  & n4886;
  assign n4889 = ~n4586 & ~n4587;
  assign n4890 = po32  & n4889;
  assign n4891 = ~n4592 & ~n4890;
  assign n4892 = n4592 & n4890;
  assign n4893 = ~n4891 & ~n4892;
  assign n4894 = ~n4888 & ~n4893;
  assign n4895 = ~n4887 & ~n4894;
  assign n4896 = po46  & ~n4895;
  assign n4897 = ~po46  & n4895;
  assign n4898 = ~n4595 & ~n4596;
  assign n4899 = po32  & n4898;
  assign n4900 = ~n4601 & ~n4899;
  assign n4901 = n4601 & n4899;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = ~n4897 & ~n4902;
  assign n4904 = ~n4896 & ~n4903;
  assign n4905 = po47  & ~n4904;
  assign n4906 = ~po47  & n4904;
  assign n4907 = ~n4604 & ~n4605;
  assign n4908 = po32  & n4907;
  assign n4909 = ~n4610 & ~n4908;
  assign n4910 = n4610 & n4908;
  assign n4911 = ~n4909 & ~n4910;
  assign n4912 = ~n4906 & ~n4911;
  assign n4913 = ~n4905 & ~n4912;
  assign n4914 = po48  & ~n4913;
  assign n4915 = ~po48  & n4913;
  assign n4916 = ~n4613 & ~n4614;
  assign n4917 = po32  & n4916;
  assign n4918 = ~n4619 & ~n4917;
  assign n4919 = n4619 & n4917;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = ~n4915 & ~n4920;
  assign n4922 = ~n4914 & ~n4921;
  assign n4923 = po49  & ~n4922;
  assign n4924 = ~po49  & n4922;
  assign n4925 = ~n4622 & ~n4623;
  assign n4926 = po32  & n4925;
  assign n4927 = ~n4628 & ~n4926;
  assign n4928 = n4628 & n4926;
  assign n4929 = ~n4927 & ~n4928;
  assign n4930 = ~n4924 & ~n4929;
  assign n4931 = ~n4923 & ~n4930;
  assign n4932 = po50  & ~n4931;
  assign n4933 = ~po50  & n4931;
  assign n4934 = ~n4631 & ~n4632;
  assign n4935 = po32  & n4934;
  assign n4936 = ~n4637 & ~n4935;
  assign n4937 = n4637 & n4935;
  assign n4938 = ~n4936 & ~n4937;
  assign n4939 = ~n4933 & ~n4938;
  assign n4940 = ~n4932 & ~n4939;
  assign n4941 = po51  & ~n4940;
  assign n4942 = ~po51  & n4940;
  assign n4943 = ~n4640 & ~n4641;
  assign n4944 = po32  & n4943;
  assign n4945 = ~n4646 & ~n4944;
  assign n4946 = n4646 & n4944;
  assign n4947 = ~n4945 & ~n4946;
  assign n4948 = ~n4942 & ~n4947;
  assign n4949 = ~n4941 & ~n4948;
  assign n4950 = po52  & ~n4949;
  assign n4951 = ~po52  & n4949;
  assign n4952 = ~n4649 & ~n4650;
  assign n4953 = po32  & n4952;
  assign n4954 = ~n4655 & ~n4953;
  assign n4955 = n4655 & n4953;
  assign n4956 = ~n4954 & ~n4955;
  assign n4957 = ~n4951 & ~n4956;
  assign n4958 = ~n4950 & ~n4957;
  assign n4959 = po53  & ~n4958;
  assign n4960 = ~po53  & n4958;
  assign n4961 = ~n4658 & ~n4659;
  assign n4962 = po32  & n4961;
  assign n4963 = ~n4664 & ~n4962;
  assign n4964 = n4664 & n4962;
  assign n4965 = ~n4963 & ~n4964;
  assign n4966 = ~n4960 & ~n4965;
  assign n4967 = ~n4959 & ~n4966;
  assign n4968 = po54  & ~n4967;
  assign n4969 = ~po54  & n4967;
  assign n4970 = ~n4667 & ~n4668;
  assign n4971 = po32  & n4970;
  assign n4972 = ~n4673 & ~n4971;
  assign n4973 = n4673 & n4971;
  assign n4974 = ~n4972 & ~n4973;
  assign n4975 = ~n4969 & ~n4974;
  assign n4976 = ~n4968 & ~n4975;
  assign n4977 = po55  & ~n4976;
  assign n4978 = ~po55  & n4976;
  assign n4979 = ~n4676 & ~n4677;
  assign n4980 = po32  & n4979;
  assign n4981 = ~n4682 & ~n4980;
  assign n4982 = n4682 & n4980;
  assign n4983 = ~n4981 & ~n4982;
  assign n4984 = ~n4978 & ~n4983;
  assign n4985 = ~n4977 & ~n4984;
  assign n4986 = po56  & ~n4985;
  assign n4987 = ~po56  & n4985;
  assign n4988 = ~n4685 & ~n4686;
  assign n4989 = po32  & n4988;
  assign n4990 = ~n4691 & ~n4989;
  assign n4991 = n4691 & n4989;
  assign n4992 = ~n4990 & ~n4991;
  assign n4993 = ~n4987 & ~n4992;
  assign n4994 = ~n4986 & ~n4993;
  assign n4995 = po57  & ~n4994;
  assign n4996 = ~po57  & n4994;
  assign n4997 = ~n4694 & ~n4695;
  assign n4998 = po32  & n4997;
  assign n4999 = ~n4700 & ~n4998;
  assign n5000 = n4700 & n4998;
  assign n5001 = ~n4999 & ~n5000;
  assign n5002 = ~n4996 & ~n5001;
  assign n5003 = ~n4995 & ~n5002;
  assign n5004 = po58  & ~n5003;
  assign n5005 = ~po58  & n5003;
  assign n5006 = ~n4703 & ~n4704;
  assign n5007 = po32  & n5006;
  assign n5008 = ~n4709 & ~n5007;
  assign n5009 = n4709 & n5007;
  assign n5010 = ~n5008 & ~n5009;
  assign n5011 = ~n5005 & ~n5010;
  assign n5012 = ~n5004 & ~n5011;
  assign n5013 = po59  & ~n5012;
  assign n5014 = ~po59  & n5012;
  assign n5015 = ~n4712 & ~n4713;
  assign n5016 = po32  & n5015;
  assign n5017 = ~n4718 & ~n5016;
  assign n5018 = n4718 & n5016;
  assign n5019 = ~n5017 & ~n5018;
  assign n5020 = ~n5014 & ~n5019;
  assign n5021 = ~n5013 & ~n5020;
  assign n5022 = po60  & ~n5021;
  assign n5023 = ~po60  & n5021;
  assign n5024 = ~n4721 & ~n4722;
  assign n5025 = po32  & n5024;
  assign n5026 = ~n4727 & ~n5025;
  assign n5027 = n4727 & n5025;
  assign n5028 = ~n5026 & ~n5027;
  assign n5029 = ~n5023 & ~n5028;
  assign n5030 = ~n5022 & ~n5029;
  assign n5031 = po61  & ~n5030;
  assign n5032 = ~po61  & n5030;
  assign n5033 = ~n4730 & ~n4731;
  assign n5034 = po32  & n5033;
  assign n5035 = ~n4736 & ~n5034;
  assign n5036 = n4736 & n5034;
  assign n5037 = ~n5035 & ~n5036;
  assign n5038 = ~n5032 & ~n5037;
  assign n5039 = ~n5031 & ~n5038;
  assign n5040 = po62  & ~n5039;
  assign n5041 = ~po62  & n5039;
  assign n5042 = ~n4739 & ~n4740;
  assign n5043 = po32  & n5042;
  assign n5044 = ~n4745 & ~n5043;
  assign n5045 = n4745 & n5043;
  assign n5046 = ~n5044 & ~n5045;
  assign n5047 = ~n5041 & ~n5046;
  assign n5048 = ~n5040 & ~n5047;
  assign n5049 = n4779 & n5048;
  assign n5050 = ~n4779 & ~n5048;
  assign n5051 = n4758 & po32 ;
  assign n5052 = ~n4757 & ~n5051;
  assign n5053 = n5050 & n5052;
  assign n5054 = ~po63  & ~n5053;
  assign n5055 = ~n5049 & ~n5054;
  assign n5056 = ~n4774 & n5055;
  assign po31  = n4770 | ~n5056;
  assign n5058 = ~n4784 & ~n4785;
  assign n5059 = po31  & n5058;
  assign n5060 = n4769 & ~n5059;
  assign n5061 = ~n4769 & n5059;
  assign n5062 = ~n5060 & ~n5061;
  assign n5063 = n4779 & ~po31 ;
  assign n5064 = ~n4779 & po31 ;
  assign n5065 = n5048 & ~n5064;
  assign n5066 = po63  & ~n5065;
  assign n5067 = ~n5050 & n5066;
  assign n5068 = ~n5040 & ~n5041;
  assign n5069 = po31  & n5068;
  assign n5070 = ~n5046 & ~n5069;
  assign n5071 = n5046 & n5069;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = pi62  & po31 ;
  assign n5074 = ~pi60  & ~pi61 ;
  assign n5075 = ~pi62  & n5074;
  assign n5076 = ~n5073 & ~n5075;
  assign n5077 = po32  & ~n5076;
  assign n5078 = ~po32  & n5076;
  assign n5079 = ~pi62  & po31 ;
  assign n5080 = pi63  & ~n5079;
  assign n5081 = n4781 & po31 ;
  assign n5082 = ~n5080 & ~n5081;
  assign n5083 = ~n5078 & n5082;
  assign n5084 = ~n5077 & ~n5083;
  assign n5085 = po33  & ~n5084;
  assign n5086 = po32  & n5056;
  assign n5087 = ~n5081 & ~n5086;
  assign n5088 = pi64  & ~n5087;
  assign n5089 = ~pi64  & n5087;
  assign n5090 = ~n5088 & ~n5089;
  assign n5091 = ~po33  & n5084;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = ~n5085 & ~n5092;
  assign n5094 = po34  & ~n5093;
  assign n5095 = ~po34  & n5093;
  assign n5096 = ~n5062 & ~n5095;
  assign n5097 = ~n5094 & ~n5096;
  assign n5098 = po35  & ~n5097;
  assign n5099 = ~po35  & n5097;
  assign n5100 = ~n4788 & ~n4789;
  assign n5101 = po31  & n5100;
  assign n5102 = ~n4794 & ~n5101;
  assign n5103 = n4794 & n5101;
  assign n5104 = ~n5102 & ~n5103;
  assign n5105 = ~n5099 & ~n5104;
  assign n5106 = ~n5098 & ~n5105;
  assign n5107 = po36  & ~n5106;
  assign n5108 = ~po36  & n5106;
  assign n5109 = ~n4797 & ~n4798;
  assign n5110 = po31  & n5109;
  assign n5111 = n4803 & n5110;
  assign n5112 = ~n4803 & ~n5110;
  assign n5113 = ~n5111 & ~n5112;
  assign n5114 = ~n5108 & ~n5113;
  assign n5115 = ~n5107 & ~n5114;
  assign n5116 = po37  & ~n5115;
  assign n5117 = ~po37  & n5115;
  assign n5118 = ~n4806 & ~n4807;
  assign n5119 = po31  & n5118;
  assign n5120 = ~n4812 & ~n5119;
  assign n5121 = n4812 & n5119;
  assign n5122 = ~n5120 & ~n5121;
  assign n5123 = ~n5117 & ~n5122;
  assign n5124 = ~n5116 & ~n5123;
  assign n5125 = po38  & ~n5124;
  assign n5126 = ~po38  & n5124;
  assign n5127 = ~n4815 & ~n4816;
  assign n5128 = po31  & n5127;
  assign n5129 = ~n4821 & ~n5128;
  assign n5130 = n4821 & n5128;
  assign n5131 = ~n5129 & ~n5130;
  assign n5132 = ~n5126 & ~n5131;
  assign n5133 = ~n5125 & ~n5132;
  assign n5134 = po39  & ~n5133;
  assign n5135 = ~po39  & n5133;
  assign n5136 = ~n4824 & ~n4825;
  assign n5137 = po31  & n5136;
  assign n5138 = ~n4830 & ~n5137;
  assign n5139 = n4830 & n5137;
  assign n5140 = ~n5138 & ~n5139;
  assign n5141 = ~n5135 & ~n5140;
  assign n5142 = ~n5134 & ~n5141;
  assign n5143 = po40  & ~n5142;
  assign n5144 = ~po40  & n5142;
  assign n5145 = ~n4833 & ~n4834;
  assign n5146 = po31  & n5145;
  assign n5147 = ~n4839 & ~n5146;
  assign n5148 = n4839 & n5146;
  assign n5149 = ~n5147 & ~n5148;
  assign n5150 = ~n5144 & ~n5149;
  assign n5151 = ~n5143 & ~n5150;
  assign n5152 = po41  & ~n5151;
  assign n5153 = ~po41  & n5151;
  assign n5154 = ~n4842 & ~n4843;
  assign n5155 = po31  & n5154;
  assign n5156 = ~n4848 & ~n5155;
  assign n5157 = n4848 & n5155;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = ~n5153 & ~n5158;
  assign n5160 = ~n5152 & ~n5159;
  assign n5161 = po42  & ~n5160;
  assign n5162 = ~po42  & n5160;
  assign n5163 = ~n4851 & ~n4852;
  assign n5164 = po31  & n5163;
  assign n5165 = ~n4857 & ~n5164;
  assign n5166 = n4857 & n5164;
  assign n5167 = ~n5165 & ~n5166;
  assign n5168 = ~n5162 & ~n5167;
  assign n5169 = ~n5161 & ~n5168;
  assign n5170 = po43  & ~n5169;
  assign n5171 = ~po43  & n5169;
  assign n5172 = ~n4860 & ~n4861;
  assign n5173 = po31  & n5172;
  assign n5174 = ~n4866 & ~n5173;
  assign n5175 = n4866 & n5173;
  assign n5176 = ~n5174 & ~n5175;
  assign n5177 = ~n5171 & ~n5176;
  assign n5178 = ~n5170 & ~n5177;
  assign n5179 = po44  & ~n5178;
  assign n5180 = ~po44  & n5178;
  assign n5181 = ~n4869 & ~n4870;
  assign n5182 = po31  & n5181;
  assign n5183 = ~n4875 & ~n5182;
  assign n5184 = n4875 & n5182;
  assign n5185 = ~n5183 & ~n5184;
  assign n5186 = ~n5180 & ~n5185;
  assign n5187 = ~n5179 & ~n5186;
  assign n5188 = po45  & ~n5187;
  assign n5189 = ~po45  & n5187;
  assign n5190 = ~n4878 & ~n4879;
  assign n5191 = po31  & n5190;
  assign n5192 = ~n4884 & ~n5191;
  assign n5193 = n4884 & n5191;
  assign n5194 = ~n5192 & ~n5193;
  assign n5195 = ~n5189 & ~n5194;
  assign n5196 = ~n5188 & ~n5195;
  assign n5197 = po46  & ~n5196;
  assign n5198 = ~po46  & n5196;
  assign n5199 = ~n4887 & ~n4888;
  assign n5200 = po31  & n5199;
  assign n5201 = ~n4893 & ~n5200;
  assign n5202 = n4893 & n5200;
  assign n5203 = ~n5201 & ~n5202;
  assign n5204 = ~n5198 & ~n5203;
  assign n5205 = ~n5197 & ~n5204;
  assign n5206 = po47  & ~n5205;
  assign n5207 = ~po47  & n5205;
  assign n5208 = ~n4896 & ~n4897;
  assign n5209 = po31  & n5208;
  assign n5210 = ~n4902 & ~n5209;
  assign n5211 = n4902 & n5209;
  assign n5212 = ~n5210 & ~n5211;
  assign n5213 = ~n5207 & ~n5212;
  assign n5214 = ~n5206 & ~n5213;
  assign n5215 = po48  & ~n5214;
  assign n5216 = ~po48  & n5214;
  assign n5217 = ~n4905 & ~n4906;
  assign n5218 = po31  & n5217;
  assign n5219 = ~n4911 & ~n5218;
  assign n5220 = n4911 & n5218;
  assign n5221 = ~n5219 & ~n5220;
  assign n5222 = ~n5216 & ~n5221;
  assign n5223 = ~n5215 & ~n5222;
  assign n5224 = po49  & ~n5223;
  assign n5225 = ~po49  & n5223;
  assign n5226 = ~n4914 & ~n4915;
  assign n5227 = po31  & n5226;
  assign n5228 = ~n4920 & ~n5227;
  assign n5229 = n4920 & n5227;
  assign n5230 = ~n5228 & ~n5229;
  assign n5231 = ~n5225 & ~n5230;
  assign n5232 = ~n5224 & ~n5231;
  assign n5233 = po50  & ~n5232;
  assign n5234 = ~po50  & n5232;
  assign n5235 = ~n4923 & ~n4924;
  assign n5236 = po31  & n5235;
  assign n5237 = ~n4929 & ~n5236;
  assign n5238 = n4929 & n5236;
  assign n5239 = ~n5237 & ~n5238;
  assign n5240 = ~n5234 & ~n5239;
  assign n5241 = ~n5233 & ~n5240;
  assign n5242 = po51  & ~n5241;
  assign n5243 = ~po51  & n5241;
  assign n5244 = ~n4932 & ~n4933;
  assign n5245 = po31  & n5244;
  assign n5246 = ~n4938 & ~n5245;
  assign n5247 = n4938 & n5245;
  assign n5248 = ~n5246 & ~n5247;
  assign n5249 = ~n5243 & ~n5248;
  assign n5250 = ~n5242 & ~n5249;
  assign n5251 = po52  & ~n5250;
  assign n5252 = ~po52  & n5250;
  assign n5253 = ~n4941 & ~n4942;
  assign n5254 = po31  & n5253;
  assign n5255 = ~n4947 & ~n5254;
  assign n5256 = n4947 & n5254;
  assign n5257 = ~n5255 & ~n5256;
  assign n5258 = ~n5252 & ~n5257;
  assign n5259 = ~n5251 & ~n5258;
  assign n5260 = po53  & ~n5259;
  assign n5261 = ~po53  & n5259;
  assign n5262 = ~n4950 & ~n4951;
  assign n5263 = po31  & n5262;
  assign n5264 = ~n4956 & ~n5263;
  assign n5265 = n4956 & n5263;
  assign n5266 = ~n5264 & ~n5265;
  assign n5267 = ~n5261 & ~n5266;
  assign n5268 = ~n5260 & ~n5267;
  assign n5269 = po54  & ~n5268;
  assign n5270 = ~po54  & n5268;
  assign n5271 = ~n4959 & ~n4960;
  assign n5272 = po31  & n5271;
  assign n5273 = ~n4965 & ~n5272;
  assign n5274 = n4965 & n5272;
  assign n5275 = ~n5273 & ~n5274;
  assign n5276 = ~n5270 & ~n5275;
  assign n5277 = ~n5269 & ~n5276;
  assign n5278 = po55  & ~n5277;
  assign n5279 = ~po55  & n5277;
  assign n5280 = ~n4968 & ~n4969;
  assign n5281 = po31  & n5280;
  assign n5282 = ~n4974 & ~n5281;
  assign n5283 = n4974 & n5281;
  assign n5284 = ~n5282 & ~n5283;
  assign n5285 = ~n5279 & ~n5284;
  assign n5286 = ~n5278 & ~n5285;
  assign n5287 = po56  & ~n5286;
  assign n5288 = ~po56  & n5286;
  assign n5289 = ~n4977 & ~n4978;
  assign n5290 = po31  & n5289;
  assign n5291 = ~n4983 & ~n5290;
  assign n5292 = n4983 & n5290;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~n5288 & ~n5293;
  assign n5295 = ~n5287 & ~n5294;
  assign n5296 = po57  & ~n5295;
  assign n5297 = ~po57  & n5295;
  assign n5298 = ~n4986 & ~n4987;
  assign n5299 = po31  & n5298;
  assign n5300 = ~n4992 & ~n5299;
  assign n5301 = n4992 & n5299;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = ~n5297 & ~n5302;
  assign n5304 = ~n5296 & ~n5303;
  assign n5305 = po58  & ~n5304;
  assign n5306 = ~po58  & n5304;
  assign n5307 = ~n4995 & ~n4996;
  assign n5308 = po31  & n5307;
  assign n5309 = ~n5001 & ~n5308;
  assign n5310 = n5001 & n5308;
  assign n5311 = ~n5309 & ~n5310;
  assign n5312 = ~n5306 & ~n5311;
  assign n5313 = ~n5305 & ~n5312;
  assign n5314 = po59  & ~n5313;
  assign n5315 = ~po59  & n5313;
  assign n5316 = ~n5004 & ~n5005;
  assign n5317 = po31  & n5316;
  assign n5318 = ~n5010 & ~n5317;
  assign n5319 = n5010 & n5317;
  assign n5320 = ~n5318 & ~n5319;
  assign n5321 = ~n5315 & ~n5320;
  assign n5322 = ~n5314 & ~n5321;
  assign n5323 = po60  & ~n5322;
  assign n5324 = ~po60  & n5322;
  assign n5325 = ~n5013 & ~n5014;
  assign n5326 = po31  & n5325;
  assign n5327 = ~n5019 & ~n5326;
  assign n5328 = n5019 & n5326;
  assign n5329 = ~n5327 & ~n5328;
  assign n5330 = ~n5324 & ~n5329;
  assign n5331 = ~n5323 & ~n5330;
  assign n5332 = po61  & ~n5331;
  assign n5333 = ~po61  & n5331;
  assign n5334 = ~n5022 & ~n5023;
  assign n5335 = po31  & n5334;
  assign n5336 = ~n5028 & ~n5335;
  assign n5337 = n5028 & n5335;
  assign n5338 = ~n5336 & ~n5337;
  assign n5339 = ~n5333 & ~n5338;
  assign n5340 = ~n5332 & ~n5339;
  assign n5341 = po62  & ~n5340;
  assign n5342 = ~po62  & n5340;
  assign n5343 = ~n5031 & ~n5032;
  assign n5344 = po31  & n5343;
  assign n5345 = ~n5037 & ~n5344;
  assign n5346 = n5037 & n5344;
  assign n5347 = ~n5345 & ~n5346;
  assign n5348 = ~n5342 & ~n5347;
  assign n5349 = ~n5341 & ~n5348;
  assign n5350 = n5072 & n5349;
  assign n5351 = ~n5072 & ~n5349;
  assign n5352 = n5050 & po31 ;
  assign n5353 = ~n5049 & ~n5352;
  assign n5354 = n5351 & n5353;
  assign n5355 = ~po63  & ~n5354;
  assign n5356 = ~n5350 & ~n5355;
  assign n5357 = ~n5067 & n5356;
  assign po30  = n5063 | ~n5357;
  assign n5359 = ~n5094 & ~n5095;
  assign n5360 = po30  & n5359;
  assign n5361 = n5062 & n5360;
  assign n5362 = ~n5062 & ~n5360;
  assign n5363 = ~n5361 & ~n5362;
  assign n5364 = n5072 & ~po30 ;
  assign n5365 = ~n5072 & po30 ;
  assign n5366 = n5349 & ~n5365;
  assign n5367 = po63  & ~n5366;
  assign n5368 = ~n5351 & n5367;
  assign n5369 = ~n5341 & ~n5342;
  assign n5370 = po30  & n5369;
  assign n5371 = ~n5347 & ~n5370;
  assign n5372 = n5347 & n5370;
  assign n5373 = ~n5371 & ~n5372;
  assign n5374 = pi60  & po30 ;
  assign n5375 = ~pi58  & ~pi59 ;
  assign n5376 = ~pi60  & n5375;
  assign n5377 = ~n5374 & ~n5376;
  assign n5378 = po31  & ~n5377;
  assign n5379 = ~po31  & n5377;
  assign n5380 = ~pi60  & po30 ;
  assign n5381 = pi61  & ~n5380;
  assign n5382 = n5074 & po30 ;
  assign n5383 = ~n5381 & ~n5382;
  assign n5384 = ~n5379 & n5383;
  assign n5385 = ~n5378 & ~n5384;
  assign n5386 = po32  & ~n5385;
  assign n5387 = ~po32  & n5385;
  assign n5388 = po31  & n5357;
  assign n5389 = ~n5382 & ~n5388;
  assign n5390 = pi62  & ~n5389;
  assign n5391 = ~pi62  & n5389;
  assign n5392 = ~n5390 & ~n5391;
  assign n5393 = ~n5387 & ~n5392;
  assign n5394 = ~n5386 & ~n5393;
  assign n5395 = po33  & ~n5394;
  assign n5396 = ~po33  & n5394;
  assign n5397 = ~n5077 & ~n5078;
  assign n5398 = po30  & n5397;
  assign n5399 = n5082 & ~n5398;
  assign n5400 = ~n5082 & n5398;
  assign n5401 = ~n5399 & ~n5400;
  assign n5402 = ~n5396 & ~n5401;
  assign n5403 = ~n5395 & ~n5402;
  assign n5404 = po34  & ~n5403;
  assign n5405 = ~n5085 & ~n5091;
  assign n5406 = po30  & n5405;
  assign n5407 = ~n5090 & ~n5406;
  assign n5408 = n5090 & n5406;
  assign n5409 = ~n5407 & ~n5408;
  assign n5410 = ~po34  & n5403;
  assign n5411 = ~n5409 & ~n5410;
  assign n5412 = ~n5404 & ~n5411;
  assign n5413 = po35  & ~n5412;
  assign n5414 = ~po35  & n5412;
  assign n5415 = ~n5363 & ~n5414;
  assign n5416 = ~n5413 & ~n5415;
  assign n5417 = po36  & ~n5416;
  assign n5418 = ~po36  & n5416;
  assign n5419 = ~n5098 & ~n5099;
  assign n5420 = po30  & n5419;
  assign n5421 = ~n5104 & ~n5420;
  assign n5422 = n5104 & n5420;
  assign n5423 = ~n5421 & ~n5422;
  assign n5424 = ~n5418 & ~n5423;
  assign n5425 = ~n5417 & ~n5424;
  assign n5426 = po37  & ~n5425;
  assign n5427 = ~po37  & n5425;
  assign n5428 = ~n5107 & ~n5108;
  assign n5429 = po30  & n5428;
  assign n5430 = ~n5113 & ~n5429;
  assign n5431 = n5113 & n5429;
  assign n5432 = ~n5430 & ~n5431;
  assign n5433 = ~n5427 & ~n5432;
  assign n5434 = ~n5426 & ~n5433;
  assign n5435 = po38  & ~n5434;
  assign n5436 = ~po38  & n5434;
  assign n5437 = ~n5116 & ~n5117;
  assign n5438 = po30  & n5437;
  assign n5439 = ~n5122 & ~n5438;
  assign n5440 = n5122 & n5438;
  assign n5441 = ~n5439 & ~n5440;
  assign n5442 = ~n5436 & ~n5441;
  assign n5443 = ~n5435 & ~n5442;
  assign n5444 = po39  & ~n5443;
  assign n5445 = ~po39  & n5443;
  assign n5446 = ~n5125 & ~n5126;
  assign n5447 = po30  & n5446;
  assign n5448 = ~n5131 & ~n5447;
  assign n5449 = n5131 & n5447;
  assign n5450 = ~n5448 & ~n5449;
  assign n5451 = ~n5445 & ~n5450;
  assign n5452 = ~n5444 & ~n5451;
  assign n5453 = po40  & ~n5452;
  assign n5454 = ~po40  & n5452;
  assign n5455 = ~n5134 & ~n5135;
  assign n5456 = po30  & n5455;
  assign n5457 = ~n5140 & ~n5456;
  assign n5458 = n5140 & n5456;
  assign n5459 = ~n5457 & ~n5458;
  assign n5460 = ~n5454 & ~n5459;
  assign n5461 = ~n5453 & ~n5460;
  assign n5462 = po41  & ~n5461;
  assign n5463 = ~po41  & n5461;
  assign n5464 = ~n5143 & ~n5144;
  assign n5465 = po30  & n5464;
  assign n5466 = ~n5149 & ~n5465;
  assign n5467 = n5149 & n5465;
  assign n5468 = ~n5466 & ~n5467;
  assign n5469 = ~n5463 & ~n5468;
  assign n5470 = ~n5462 & ~n5469;
  assign n5471 = po42  & ~n5470;
  assign n5472 = ~po42  & n5470;
  assign n5473 = ~n5152 & ~n5153;
  assign n5474 = po30  & n5473;
  assign n5475 = ~n5158 & ~n5474;
  assign n5476 = n5158 & n5474;
  assign n5477 = ~n5475 & ~n5476;
  assign n5478 = ~n5472 & ~n5477;
  assign n5479 = ~n5471 & ~n5478;
  assign n5480 = po43  & ~n5479;
  assign n5481 = ~po43  & n5479;
  assign n5482 = ~n5161 & ~n5162;
  assign n5483 = po30  & n5482;
  assign n5484 = ~n5167 & ~n5483;
  assign n5485 = n5167 & n5483;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = ~n5481 & ~n5486;
  assign n5488 = ~n5480 & ~n5487;
  assign n5489 = po44  & ~n5488;
  assign n5490 = ~po44  & n5488;
  assign n5491 = ~n5170 & ~n5171;
  assign n5492 = po30  & n5491;
  assign n5493 = ~n5176 & ~n5492;
  assign n5494 = n5176 & n5492;
  assign n5495 = ~n5493 & ~n5494;
  assign n5496 = ~n5490 & ~n5495;
  assign n5497 = ~n5489 & ~n5496;
  assign n5498 = po45  & ~n5497;
  assign n5499 = ~po45  & n5497;
  assign n5500 = ~n5179 & ~n5180;
  assign n5501 = po30  & n5500;
  assign n5502 = ~n5185 & ~n5501;
  assign n5503 = n5185 & n5501;
  assign n5504 = ~n5502 & ~n5503;
  assign n5505 = ~n5499 & ~n5504;
  assign n5506 = ~n5498 & ~n5505;
  assign n5507 = po46  & ~n5506;
  assign n5508 = ~po46  & n5506;
  assign n5509 = ~n5188 & ~n5189;
  assign n5510 = po30  & n5509;
  assign n5511 = ~n5194 & ~n5510;
  assign n5512 = n5194 & n5510;
  assign n5513 = ~n5511 & ~n5512;
  assign n5514 = ~n5508 & ~n5513;
  assign n5515 = ~n5507 & ~n5514;
  assign n5516 = po47  & ~n5515;
  assign n5517 = ~po47  & n5515;
  assign n5518 = ~n5197 & ~n5198;
  assign n5519 = po30  & n5518;
  assign n5520 = ~n5203 & ~n5519;
  assign n5521 = n5203 & n5519;
  assign n5522 = ~n5520 & ~n5521;
  assign n5523 = ~n5517 & ~n5522;
  assign n5524 = ~n5516 & ~n5523;
  assign n5525 = po48  & ~n5524;
  assign n5526 = ~po48  & n5524;
  assign n5527 = ~n5206 & ~n5207;
  assign n5528 = po30  & n5527;
  assign n5529 = ~n5212 & ~n5528;
  assign n5530 = n5212 & n5528;
  assign n5531 = ~n5529 & ~n5530;
  assign n5532 = ~n5526 & ~n5531;
  assign n5533 = ~n5525 & ~n5532;
  assign n5534 = po49  & ~n5533;
  assign n5535 = ~po49  & n5533;
  assign n5536 = ~n5215 & ~n5216;
  assign n5537 = po30  & n5536;
  assign n5538 = ~n5221 & ~n5537;
  assign n5539 = n5221 & n5537;
  assign n5540 = ~n5538 & ~n5539;
  assign n5541 = ~n5535 & ~n5540;
  assign n5542 = ~n5534 & ~n5541;
  assign n5543 = po50  & ~n5542;
  assign n5544 = ~po50  & n5542;
  assign n5545 = ~n5224 & ~n5225;
  assign n5546 = po30  & n5545;
  assign n5547 = ~n5230 & ~n5546;
  assign n5548 = n5230 & n5546;
  assign n5549 = ~n5547 & ~n5548;
  assign n5550 = ~n5544 & ~n5549;
  assign n5551 = ~n5543 & ~n5550;
  assign n5552 = po51  & ~n5551;
  assign n5553 = ~po51  & n5551;
  assign n5554 = ~n5233 & ~n5234;
  assign n5555 = po30  & n5554;
  assign n5556 = ~n5239 & ~n5555;
  assign n5557 = n5239 & n5555;
  assign n5558 = ~n5556 & ~n5557;
  assign n5559 = ~n5553 & ~n5558;
  assign n5560 = ~n5552 & ~n5559;
  assign n5561 = po52  & ~n5560;
  assign n5562 = ~po52  & n5560;
  assign n5563 = ~n5242 & ~n5243;
  assign n5564 = po30  & n5563;
  assign n5565 = ~n5248 & ~n5564;
  assign n5566 = n5248 & n5564;
  assign n5567 = ~n5565 & ~n5566;
  assign n5568 = ~n5562 & ~n5567;
  assign n5569 = ~n5561 & ~n5568;
  assign n5570 = po53  & ~n5569;
  assign n5571 = ~po53  & n5569;
  assign n5572 = ~n5251 & ~n5252;
  assign n5573 = po30  & n5572;
  assign n5574 = ~n5257 & ~n5573;
  assign n5575 = n5257 & n5573;
  assign n5576 = ~n5574 & ~n5575;
  assign n5577 = ~n5571 & ~n5576;
  assign n5578 = ~n5570 & ~n5577;
  assign n5579 = po54  & ~n5578;
  assign n5580 = ~po54  & n5578;
  assign n5581 = ~n5260 & ~n5261;
  assign n5582 = po30  & n5581;
  assign n5583 = ~n5266 & ~n5582;
  assign n5584 = n5266 & n5582;
  assign n5585 = ~n5583 & ~n5584;
  assign n5586 = ~n5580 & ~n5585;
  assign n5587 = ~n5579 & ~n5586;
  assign n5588 = po55  & ~n5587;
  assign n5589 = ~po55  & n5587;
  assign n5590 = ~n5269 & ~n5270;
  assign n5591 = po30  & n5590;
  assign n5592 = ~n5275 & ~n5591;
  assign n5593 = n5275 & n5591;
  assign n5594 = ~n5592 & ~n5593;
  assign n5595 = ~n5589 & ~n5594;
  assign n5596 = ~n5588 & ~n5595;
  assign n5597 = po56  & ~n5596;
  assign n5598 = ~po56  & n5596;
  assign n5599 = ~n5278 & ~n5279;
  assign n5600 = po30  & n5599;
  assign n5601 = ~n5284 & ~n5600;
  assign n5602 = n5284 & n5600;
  assign n5603 = ~n5601 & ~n5602;
  assign n5604 = ~n5598 & ~n5603;
  assign n5605 = ~n5597 & ~n5604;
  assign n5606 = po57  & ~n5605;
  assign n5607 = ~po57  & n5605;
  assign n5608 = ~n5287 & ~n5288;
  assign n5609 = po30  & n5608;
  assign n5610 = ~n5293 & ~n5609;
  assign n5611 = n5293 & n5609;
  assign n5612 = ~n5610 & ~n5611;
  assign n5613 = ~n5607 & ~n5612;
  assign n5614 = ~n5606 & ~n5613;
  assign n5615 = po58  & ~n5614;
  assign n5616 = ~po58  & n5614;
  assign n5617 = ~n5296 & ~n5297;
  assign n5618 = po30  & n5617;
  assign n5619 = ~n5302 & ~n5618;
  assign n5620 = n5302 & n5618;
  assign n5621 = ~n5619 & ~n5620;
  assign n5622 = ~n5616 & ~n5621;
  assign n5623 = ~n5615 & ~n5622;
  assign n5624 = po59  & ~n5623;
  assign n5625 = ~po59  & n5623;
  assign n5626 = ~n5305 & ~n5306;
  assign n5627 = po30  & n5626;
  assign n5628 = ~n5311 & ~n5627;
  assign n5629 = n5311 & n5627;
  assign n5630 = ~n5628 & ~n5629;
  assign n5631 = ~n5625 & ~n5630;
  assign n5632 = ~n5624 & ~n5631;
  assign n5633 = po60  & ~n5632;
  assign n5634 = ~po60  & n5632;
  assign n5635 = ~n5314 & ~n5315;
  assign n5636 = po30  & n5635;
  assign n5637 = ~n5320 & ~n5636;
  assign n5638 = n5320 & n5636;
  assign n5639 = ~n5637 & ~n5638;
  assign n5640 = ~n5634 & ~n5639;
  assign n5641 = ~n5633 & ~n5640;
  assign n5642 = po61  & ~n5641;
  assign n5643 = ~po61  & n5641;
  assign n5644 = ~n5323 & ~n5324;
  assign n5645 = po30  & n5644;
  assign n5646 = ~n5329 & ~n5645;
  assign n5647 = n5329 & n5645;
  assign n5648 = ~n5646 & ~n5647;
  assign n5649 = ~n5643 & ~n5648;
  assign n5650 = ~n5642 & ~n5649;
  assign n5651 = po62  & ~n5650;
  assign n5652 = ~po62  & n5650;
  assign n5653 = ~n5332 & ~n5333;
  assign n5654 = po30  & n5653;
  assign n5655 = ~n5338 & ~n5654;
  assign n5656 = n5338 & n5654;
  assign n5657 = ~n5655 & ~n5656;
  assign n5658 = ~n5652 & ~n5657;
  assign n5659 = ~n5651 & ~n5658;
  assign n5660 = n5373 & n5659;
  assign n5661 = ~n5373 & ~n5659;
  assign n5662 = n5351 & po30 ;
  assign n5663 = ~n5350 & ~n5662;
  assign n5664 = n5661 & n5663;
  assign n5665 = ~po63  & ~n5664;
  assign n5666 = ~n5660 & ~n5665;
  assign n5667 = ~n5368 & n5666;
  assign po29  = n5364 | ~n5667;
  assign n5669 = ~n5413 & ~n5414;
  assign n5670 = po29  & n5669;
  assign n5671 = ~n5363 & ~n5670;
  assign n5672 = n5363 & n5670;
  assign n5673 = ~n5671 & ~n5672;
  assign n5674 = n5373 & ~po29 ;
  assign n5675 = ~n5373 & po29 ;
  assign n5676 = n5659 & ~n5675;
  assign n5677 = po63  & ~n5676;
  assign n5678 = ~n5661 & n5677;
  assign n5679 = ~n5651 & ~n5652;
  assign n5680 = po29  & n5679;
  assign n5681 = ~n5657 & ~n5680;
  assign n5682 = n5657 & n5680;
  assign n5683 = ~n5681 & ~n5682;
  assign n5684 = pi58  & po29 ;
  assign n5685 = ~pi56  & ~pi57 ;
  assign n5686 = ~pi58  & n5685;
  assign n5687 = ~n5684 & ~n5686;
  assign n5688 = po30  & ~n5687;
  assign n5689 = ~po30  & n5687;
  assign n5690 = ~pi58  & po29 ;
  assign n5691 = pi59  & ~n5690;
  assign n5692 = n5375 & po29 ;
  assign n5693 = ~n5691 & ~n5692;
  assign n5694 = ~n5689 & n5693;
  assign n5695 = ~n5688 & ~n5694;
  assign n5696 = po31  & ~n5695;
  assign n5697 = ~po31  & n5695;
  assign n5698 = po30  & n5667;
  assign n5699 = ~n5692 & ~n5698;
  assign n5700 = pi60  & ~n5699;
  assign n5701 = ~pi60  & n5699;
  assign n5702 = ~n5700 & ~n5701;
  assign n5703 = ~n5697 & ~n5702;
  assign n5704 = ~n5696 & ~n5703;
  assign n5705 = po32  & ~n5704;
  assign n5706 = ~po32  & n5704;
  assign n5707 = ~n5378 & ~n5379;
  assign n5708 = po29  & n5707;
  assign n5709 = n5383 & ~n5708;
  assign n5710 = ~n5383 & n5708;
  assign n5711 = ~n5709 & ~n5710;
  assign n5712 = ~n5706 & ~n5711;
  assign n5713 = ~n5705 & ~n5712;
  assign n5714 = po33  & ~n5713;
  assign n5715 = ~po33  & n5713;
  assign n5716 = ~n5386 & ~n5387;
  assign n5717 = po29  & n5716;
  assign n5718 = ~n5392 & ~n5717;
  assign n5719 = n5392 & n5717;
  assign n5720 = ~n5718 & ~n5719;
  assign n5721 = ~n5715 & ~n5720;
  assign n5722 = ~n5714 & ~n5721;
  assign n5723 = po34  & ~n5722;
  assign n5724 = ~po34  & n5722;
  assign n5725 = ~n5395 & ~n5396;
  assign n5726 = po29  & n5725;
  assign n5727 = n5401 & n5726;
  assign n5728 = ~n5401 & ~n5726;
  assign n5729 = ~n5727 & ~n5728;
  assign n5730 = ~n5724 & ~n5729;
  assign n5731 = ~n5723 & ~n5730;
  assign n5732 = po35  & ~n5731;
  assign n5733 = ~n5404 & ~n5410;
  assign n5734 = po29  & n5733;
  assign n5735 = ~n5409 & ~n5734;
  assign n5736 = n5409 & n5734;
  assign n5737 = ~n5735 & ~n5736;
  assign n5738 = ~po35  & n5731;
  assign n5739 = ~n5737 & ~n5738;
  assign n5740 = ~n5732 & ~n5739;
  assign n5741 = po36  & ~n5740;
  assign n5742 = ~po36  & n5740;
  assign n5743 = ~n5673 & ~n5742;
  assign n5744 = ~n5741 & ~n5743;
  assign n5745 = po37  & ~n5744;
  assign n5746 = ~po37  & n5744;
  assign n5747 = ~n5417 & ~n5418;
  assign n5748 = po29  & n5747;
  assign n5749 = ~n5423 & ~n5748;
  assign n5750 = n5423 & n5748;
  assign n5751 = ~n5749 & ~n5750;
  assign n5752 = ~n5746 & ~n5751;
  assign n5753 = ~n5745 & ~n5752;
  assign n5754 = po38  & ~n5753;
  assign n5755 = ~po38  & n5753;
  assign n5756 = ~n5426 & ~n5427;
  assign n5757 = po29  & n5756;
  assign n5758 = ~n5432 & ~n5757;
  assign n5759 = n5432 & n5757;
  assign n5760 = ~n5758 & ~n5759;
  assign n5761 = ~n5755 & ~n5760;
  assign n5762 = ~n5754 & ~n5761;
  assign n5763 = po39  & ~n5762;
  assign n5764 = ~po39  & n5762;
  assign n5765 = ~n5435 & ~n5436;
  assign n5766 = po29  & n5765;
  assign n5767 = ~n5441 & ~n5766;
  assign n5768 = n5441 & n5766;
  assign n5769 = ~n5767 & ~n5768;
  assign n5770 = ~n5764 & ~n5769;
  assign n5771 = ~n5763 & ~n5770;
  assign n5772 = po40  & ~n5771;
  assign n5773 = ~po40  & n5771;
  assign n5774 = ~n5444 & ~n5445;
  assign n5775 = po29  & n5774;
  assign n5776 = ~n5450 & ~n5775;
  assign n5777 = n5450 & n5775;
  assign n5778 = ~n5776 & ~n5777;
  assign n5779 = ~n5773 & ~n5778;
  assign n5780 = ~n5772 & ~n5779;
  assign n5781 = po41  & ~n5780;
  assign n5782 = ~po41  & n5780;
  assign n5783 = ~n5453 & ~n5454;
  assign n5784 = po29  & n5783;
  assign n5785 = ~n5459 & ~n5784;
  assign n5786 = n5459 & n5784;
  assign n5787 = ~n5785 & ~n5786;
  assign n5788 = ~n5782 & ~n5787;
  assign n5789 = ~n5781 & ~n5788;
  assign n5790 = po42  & ~n5789;
  assign n5791 = ~po42  & n5789;
  assign n5792 = ~n5462 & ~n5463;
  assign n5793 = po29  & n5792;
  assign n5794 = ~n5468 & ~n5793;
  assign n5795 = n5468 & n5793;
  assign n5796 = ~n5794 & ~n5795;
  assign n5797 = ~n5791 & ~n5796;
  assign n5798 = ~n5790 & ~n5797;
  assign n5799 = po43  & ~n5798;
  assign n5800 = ~po43  & n5798;
  assign n5801 = ~n5471 & ~n5472;
  assign n5802 = po29  & n5801;
  assign n5803 = ~n5477 & ~n5802;
  assign n5804 = n5477 & n5802;
  assign n5805 = ~n5803 & ~n5804;
  assign n5806 = ~n5800 & ~n5805;
  assign n5807 = ~n5799 & ~n5806;
  assign n5808 = po44  & ~n5807;
  assign n5809 = ~po44  & n5807;
  assign n5810 = ~n5480 & ~n5481;
  assign n5811 = po29  & n5810;
  assign n5812 = ~n5486 & ~n5811;
  assign n5813 = n5486 & n5811;
  assign n5814 = ~n5812 & ~n5813;
  assign n5815 = ~n5809 & ~n5814;
  assign n5816 = ~n5808 & ~n5815;
  assign n5817 = po45  & ~n5816;
  assign n5818 = ~po45  & n5816;
  assign n5819 = ~n5489 & ~n5490;
  assign n5820 = po29  & n5819;
  assign n5821 = ~n5495 & ~n5820;
  assign n5822 = n5495 & n5820;
  assign n5823 = ~n5821 & ~n5822;
  assign n5824 = ~n5818 & ~n5823;
  assign n5825 = ~n5817 & ~n5824;
  assign n5826 = po46  & ~n5825;
  assign n5827 = ~po46  & n5825;
  assign n5828 = ~n5498 & ~n5499;
  assign n5829 = po29  & n5828;
  assign n5830 = ~n5504 & ~n5829;
  assign n5831 = n5504 & n5829;
  assign n5832 = ~n5830 & ~n5831;
  assign n5833 = ~n5827 & ~n5832;
  assign n5834 = ~n5826 & ~n5833;
  assign n5835 = po47  & ~n5834;
  assign n5836 = ~po47  & n5834;
  assign n5837 = ~n5507 & ~n5508;
  assign n5838 = po29  & n5837;
  assign n5839 = ~n5513 & ~n5838;
  assign n5840 = n5513 & n5838;
  assign n5841 = ~n5839 & ~n5840;
  assign n5842 = ~n5836 & ~n5841;
  assign n5843 = ~n5835 & ~n5842;
  assign n5844 = po48  & ~n5843;
  assign n5845 = ~po48  & n5843;
  assign n5846 = ~n5516 & ~n5517;
  assign n5847 = po29  & n5846;
  assign n5848 = ~n5522 & ~n5847;
  assign n5849 = n5522 & n5847;
  assign n5850 = ~n5848 & ~n5849;
  assign n5851 = ~n5845 & ~n5850;
  assign n5852 = ~n5844 & ~n5851;
  assign n5853 = po49  & ~n5852;
  assign n5854 = ~po49  & n5852;
  assign n5855 = ~n5525 & ~n5526;
  assign n5856 = po29  & n5855;
  assign n5857 = ~n5531 & ~n5856;
  assign n5858 = n5531 & n5856;
  assign n5859 = ~n5857 & ~n5858;
  assign n5860 = ~n5854 & ~n5859;
  assign n5861 = ~n5853 & ~n5860;
  assign n5862 = po50  & ~n5861;
  assign n5863 = ~po50  & n5861;
  assign n5864 = ~n5534 & ~n5535;
  assign n5865 = po29  & n5864;
  assign n5866 = ~n5540 & ~n5865;
  assign n5867 = n5540 & n5865;
  assign n5868 = ~n5866 & ~n5867;
  assign n5869 = ~n5863 & ~n5868;
  assign n5870 = ~n5862 & ~n5869;
  assign n5871 = po51  & ~n5870;
  assign n5872 = ~po51  & n5870;
  assign n5873 = ~n5543 & ~n5544;
  assign n5874 = po29  & n5873;
  assign n5875 = ~n5549 & ~n5874;
  assign n5876 = n5549 & n5874;
  assign n5877 = ~n5875 & ~n5876;
  assign n5878 = ~n5872 & ~n5877;
  assign n5879 = ~n5871 & ~n5878;
  assign n5880 = po52  & ~n5879;
  assign n5881 = ~po52  & n5879;
  assign n5882 = ~n5552 & ~n5553;
  assign n5883 = po29  & n5882;
  assign n5884 = ~n5558 & ~n5883;
  assign n5885 = n5558 & n5883;
  assign n5886 = ~n5884 & ~n5885;
  assign n5887 = ~n5881 & ~n5886;
  assign n5888 = ~n5880 & ~n5887;
  assign n5889 = po53  & ~n5888;
  assign n5890 = ~po53  & n5888;
  assign n5891 = ~n5561 & ~n5562;
  assign n5892 = po29  & n5891;
  assign n5893 = ~n5567 & ~n5892;
  assign n5894 = n5567 & n5892;
  assign n5895 = ~n5893 & ~n5894;
  assign n5896 = ~n5890 & ~n5895;
  assign n5897 = ~n5889 & ~n5896;
  assign n5898 = po54  & ~n5897;
  assign n5899 = ~po54  & n5897;
  assign n5900 = ~n5570 & ~n5571;
  assign n5901 = po29  & n5900;
  assign n5902 = ~n5576 & ~n5901;
  assign n5903 = n5576 & n5901;
  assign n5904 = ~n5902 & ~n5903;
  assign n5905 = ~n5899 & ~n5904;
  assign n5906 = ~n5898 & ~n5905;
  assign n5907 = po55  & ~n5906;
  assign n5908 = ~po55  & n5906;
  assign n5909 = ~n5579 & ~n5580;
  assign n5910 = po29  & n5909;
  assign n5911 = ~n5585 & ~n5910;
  assign n5912 = n5585 & n5910;
  assign n5913 = ~n5911 & ~n5912;
  assign n5914 = ~n5908 & ~n5913;
  assign n5915 = ~n5907 & ~n5914;
  assign n5916 = po56  & ~n5915;
  assign n5917 = ~po56  & n5915;
  assign n5918 = ~n5588 & ~n5589;
  assign n5919 = po29  & n5918;
  assign n5920 = ~n5594 & ~n5919;
  assign n5921 = n5594 & n5919;
  assign n5922 = ~n5920 & ~n5921;
  assign n5923 = ~n5917 & ~n5922;
  assign n5924 = ~n5916 & ~n5923;
  assign n5925 = po57  & ~n5924;
  assign n5926 = ~po57  & n5924;
  assign n5927 = ~n5597 & ~n5598;
  assign n5928 = po29  & n5927;
  assign n5929 = ~n5603 & ~n5928;
  assign n5930 = n5603 & n5928;
  assign n5931 = ~n5929 & ~n5930;
  assign n5932 = ~n5926 & ~n5931;
  assign n5933 = ~n5925 & ~n5932;
  assign n5934 = po58  & ~n5933;
  assign n5935 = ~po58  & n5933;
  assign n5936 = ~n5606 & ~n5607;
  assign n5937 = po29  & n5936;
  assign n5938 = ~n5612 & ~n5937;
  assign n5939 = n5612 & n5937;
  assign n5940 = ~n5938 & ~n5939;
  assign n5941 = ~n5935 & ~n5940;
  assign n5942 = ~n5934 & ~n5941;
  assign n5943 = po59  & ~n5942;
  assign n5944 = ~po59  & n5942;
  assign n5945 = ~n5615 & ~n5616;
  assign n5946 = po29  & n5945;
  assign n5947 = ~n5621 & ~n5946;
  assign n5948 = n5621 & n5946;
  assign n5949 = ~n5947 & ~n5948;
  assign n5950 = ~n5944 & ~n5949;
  assign n5951 = ~n5943 & ~n5950;
  assign n5952 = po60  & ~n5951;
  assign n5953 = ~po60  & n5951;
  assign n5954 = ~n5624 & ~n5625;
  assign n5955 = po29  & n5954;
  assign n5956 = ~n5630 & ~n5955;
  assign n5957 = n5630 & n5955;
  assign n5958 = ~n5956 & ~n5957;
  assign n5959 = ~n5953 & ~n5958;
  assign n5960 = ~n5952 & ~n5959;
  assign n5961 = po61  & ~n5960;
  assign n5962 = ~po61  & n5960;
  assign n5963 = ~n5633 & ~n5634;
  assign n5964 = po29  & n5963;
  assign n5965 = ~n5639 & ~n5964;
  assign n5966 = n5639 & n5964;
  assign n5967 = ~n5965 & ~n5966;
  assign n5968 = ~n5962 & ~n5967;
  assign n5969 = ~n5961 & ~n5968;
  assign n5970 = po62  & ~n5969;
  assign n5971 = ~po62  & n5969;
  assign n5972 = ~n5642 & ~n5643;
  assign n5973 = po29  & n5972;
  assign n5974 = ~n5648 & ~n5973;
  assign n5975 = n5648 & n5973;
  assign n5976 = ~n5974 & ~n5975;
  assign n5977 = ~n5971 & ~n5976;
  assign n5978 = ~n5970 & ~n5977;
  assign n5979 = n5683 & n5978;
  assign n5980 = ~n5683 & ~n5978;
  assign n5981 = n5661 & po29 ;
  assign n5982 = ~n5660 & ~n5981;
  assign n5983 = n5980 & n5982;
  assign n5984 = ~po63  & ~n5983;
  assign n5985 = ~n5979 & ~n5984;
  assign n5986 = ~n5678 & n5985;
  assign po28  = n5674 | ~n5986;
  assign n5988 = ~n5741 & ~n5742;
  assign n5989 = po28  & n5988;
  assign n5990 = ~n5673 & ~n5989;
  assign n5991 = n5673 & n5989;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = n5683 & ~po28 ;
  assign n5994 = ~n5683 & po28 ;
  assign n5995 = n5978 & ~n5994;
  assign n5996 = po63  & ~n5995;
  assign n5997 = ~n5980 & n5996;
  assign n5998 = ~n5970 & ~n5971;
  assign n5999 = po28  & n5998;
  assign n6000 = ~n5976 & ~n5999;
  assign n6001 = n5976 & n5999;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = pi56  & po28 ;
  assign n6004 = ~pi54  & ~pi55 ;
  assign n6005 = ~pi56  & n6004;
  assign n6006 = ~n6003 & ~n6005;
  assign n6007 = po29  & ~n6006;
  assign n6008 = ~po29  & n6006;
  assign n6009 = ~pi56  & po28 ;
  assign n6010 = pi57  & ~n6009;
  assign n6011 = n5685 & po28 ;
  assign n6012 = ~n6010 & ~n6011;
  assign n6013 = ~n6008 & n6012;
  assign n6014 = ~n6007 & ~n6013;
  assign n6015 = po30  & ~n6014;
  assign n6016 = ~po30  & n6014;
  assign n6017 = po29  & n5986;
  assign n6018 = ~n6011 & ~n6017;
  assign n6019 = pi58  & ~n6018;
  assign n6020 = ~pi58  & n6018;
  assign n6021 = ~n6019 & ~n6020;
  assign n6022 = ~n6016 & ~n6021;
  assign n6023 = ~n6015 & ~n6022;
  assign n6024 = po31  & ~n6023;
  assign n6025 = ~po31  & n6023;
  assign n6026 = ~n5688 & ~n5689;
  assign n6027 = po28  & n6026;
  assign n6028 = n5693 & ~n6027;
  assign n6029 = ~n5693 & n6027;
  assign n6030 = ~n6028 & ~n6029;
  assign n6031 = ~n6025 & ~n6030;
  assign n6032 = ~n6024 & ~n6031;
  assign n6033 = po32  & ~n6032;
  assign n6034 = ~po32  & n6032;
  assign n6035 = ~n5696 & ~n5697;
  assign n6036 = po28  & n6035;
  assign n6037 = ~n5702 & ~n6036;
  assign n6038 = n5702 & n6036;
  assign n6039 = ~n6037 & ~n6038;
  assign n6040 = ~n6034 & ~n6039;
  assign n6041 = ~n6033 & ~n6040;
  assign n6042 = po33  & ~n6041;
  assign n6043 = ~po33  & n6041;
  assign n6044 = ~n5705 & ~n5706;
  assign n6045 = po28  & n6044;
  assign n6046 = n5711 & n6045;
  assign n6047 = ~n5711 & ~n6045;
  assign n6048 = ~n6046 & ~n6047;
  assign n6049 = ~n6043 & ~n6048;
  assign n6050 = ~n6042 & ~n6049;
  assign n6051 = po34  & ~n6050;
  assign n6052 = ~po34  & n6050;
  assign n6053 = ~n5714 & ~n5715;
  assign n6054 = po28  & n6053;
  assign n6055 = ~n5720 & ~n6054;
  assign n6056 = n5720 & n6054;
  assign n6057 = ~n6055 & ~n6056;
  assign n6058 = ~n6052 & ~n6057;
  assign n6059 = ~n6051 & ~n6058;
  assign n6060 = po35  & ~n6059;
  assign n6061 = ~po35  & n6059;
  assign n6062 = ~n5723 & ~n5724;
  assign n6063 = po28  & n6062;
  assign n6064 = ~n5729 & ~n6063;
  assign n6065 = n5729 & n6063;
  assign n6066 = ~n6064 & ~n6065;
  assign n6067 = ~n6061 & ~n6066;
  assign n6068 = ~n6060 & ~n6067;
  assign n6069 = po36  & ~n6068;
  assign n6070 = ~n5732 & ~n5738;
  assign n6071 = po28  & n6070;
  assign n6072 = ~n5737 & ~n6071;
  assign n6073 = n5737 & n6071;
  assign n6074 = ~n6072 & ~n6073;
  assign n6075 = ~po36  & n6068;
  assign n6076 = ~n6074 & ~n6075;
  assign n6077 = ~n6069 & ~n6076;
  assign n6078 = po37  & ~n6077;
  assign n6079 = ~po37  & n6077;
  assign n6080 = ~n5992 & ~n6079;
  assign n6081 = ~n6078 & ~n6080;
  assign n6082 = po38  & ~n6081;
  assign n6083 = ~po38  & n6081;
  assign n6084 = ~n5745 & ~n5746;
  assign n6085 = po28  & n6084;
  assign n6086 = ~n5751 & ~n6085;
  assign n6087 = n5751 & n6085;
  assign n6088 = ~n6086 & ~n6087;
  assign n6089 = ~n6083 & ~n6088;
  assign n6090 = ~n6082 & ~n6089;
  assign n6091 = po39  & ~n6090;
  assign n6092 = ~po39  & n6090;
  assign n6093 = ~n5754 & ~n5755;
  assign n6094 = po28  & n6093;
  assign n6095 = ~n5760 & ~n6094;
  assign n6096 = n5760 & n6094;
  assign n6097 = ~n6095 & ~n6096;
  assign n6098 = ~n6092 & ~n6097;
  assign n6099 = ~n6091 & ~n6098;
  assign n6100 = po40  & ~n6099;
  assign n6101 = ~po40  & n6099;
  assign n6102 = ~n5763 & ~n5764;
  assign n6103 = po28  & n6102;
  assign n6104 = ~n5769 & ~n6103;
  assign n6105 = n5769 & n6103;
  assign n6106 = ~n6104 & ~n6105;
  assign n6107 = ~n6101 & ~n6106;
  assign n6108 = ~n6100 & ~n6107;
  assign n6109 = po41  & ~n6108;
  assign n6110 = ~po41  & n6108;
  assign n6111 = ~n5772 & ~n5773;
  assign n6112 = po28  & n6111;
  assign n6113 = ~n5778 & ~n6112;
  assign n6114 = n5778 & n6112;
  assign n6115 = ~n6113 & ~n6114;
  assign n6116 = ~n6110 & ~n6115;
  assign n6117 = ~n6109 & ~n6116;
  assign n6118 = po42  & ~n6117;
  assign n6119 = ~po42  & n6117;
  assign n6120 = ~n5781 & ~n5782;
  assign n6121 = po28  & n6120;
  assign n6122 = ~n5787 & ~n6121;
  assign n6123 = n5787 & n6121;
  assign n6124 = ~n6122 & ~n6123;
  assign n6125 = ~n6119 & ~n6124;
  assign n6126 = ~n6118 & ~n6125;
  assign n6127 = po43  & ~n6126;
  assign n6128 = ~po43  & n6126;
  assign n6129 = ~n5790 & ~n5791;
  assign n6130 = po28  & n6129;
  assign n6131 = ~n5796 & ~n6130;
  assign n6132 = n5796 & n6130;
  assign n6133 = ~n6131 & ~n6132;
  assign n6134 = ~n6128 & ~n6133;
  assign n6135 = ~n6127 & ~n6134;
  assign n6136 = po44  & ~n6135;
  assign n6137 = ~po44  & n6135;
  assign n6138 = ~n5799 & ~n5800;
  assign n6139 = po28  & n6138;
  assign n6140 = ~n5805 & ~n6139;
  assign n6141 = n5805 & n6139;
  assign n6142 = ~n6140 & ~n6141;
  assign n6143 = ~n6137 & ~n6142;
  assign n6144 = ~n6136 & ~n6143;
  assign n6145 = po45  & ~n6144;
  assign n6146 = ~po45  & n6144;
  assign n6147 = ~n5808 & ~n5809;
  assign n6148 = po28  & n6147;
  assign n6149 = ~n5814 & ~n6148;
  assign n6150 = n5814 & n6148;
  assign n6151 = ~n6149 & ~n6150;
  assign n6152 = ~n6146 & ~n6151;
  assign n6153 = ~n6145 & ~n6152;
  assign n6154 = po46  & ~n6153;
  assign n6155 = ~po46  & n6153;
  assign n6156 = ~n5817 & ~n5818;
  assign n6157 = po28  & n6156;
  assign n6158 = ~n5823 & ~n6157;
  assign n6159 = n5823 & n6157;
  assign n6160 = ~n6158 & ~n6159;
  assign n6161 = ~n6155 & ~n6160;
  assign n6162 = ~n6154 & ~n6161;
  assign n6163 = po47  & ~n6162;
  assign n6164 = ~po47  & n6162;
  assign n6165 = ~n5826 & ~n5827;
  assign n6166 = po28  & n6165;
  assign n6167 = ~n5832 & ~n6166;
  assign n6168 = n5832 & n6166;
  assign n6169 = ~n6167 & ~n6168;
  assign n6170 = ~n6164 & ~n6169;
  assign n6171 = ~n6163 & ~n6170;
  assign n6172 = po48  & ~n6171;
  assign n6173 = ~po48  & n6171;
  assign n6174 = ~n5835 & ~n5836;
  assign n6175 = po28  & n6174;
  assign n6176 = ~n5841 & ~n6175;
  assign n6177 = n5841 & n6175;
  assign n6178 = ~n6176 & ~n6177;
  assign n6179 = ~n6173 & ~n6178;
  assign n6180 = ~n6172 & ~n6179;
  assign n6181 = po49  & ~n6180;
  assign n6182 = ~po49  & n6180;
  assign n6183 = ~n5844 & ~n5845;
  assign n6184 = po28  & n6183;
  assign n6185 = ~n5850 & ~n6184;
  assign n6186 = n5850 & n6184;
  assign n6187 = ~n6185 & ~n6186;
  assign n6188 = ~n6182 & ~n6187;
  assign n6189 = ~n6181 & ~n6188;
  assign n6190 = po50  & ~n6189;
  assign n6191 = ~po50  & n6189;
  assign n6192 = ~n5853 & ~n5854;
  assign n6193 = po28  & n6192;
  assign n6194 = ~n5859 & ~n6193;
  assign n6195 = n5859 & n6193;
  assign n6196 = ~n6194 & ~n6195;
  assign n6197 = ~n6191 & ~n6196;
  assign n6198 = ~n6190 & ~n6197;
  assign n6199 = po51  & ~n6198;
  assign n6200 = ~po51  & n6198;
  assign n6201 = ~n5862 & ~n5863;
  assign n6202 = po28  & n6201;
  assign n6203 = ~n5868 & ~n6202;
  assign n6204 = n5868 & n6202;
  assign n6205 = ~n6203 & ~n6204;
  assign n6206 = ~n6200 & ~n6205;
  assign n6207 = ~n6199 & ~n6206;
  assign n6208 = po52  & ~n6207;
  assign n6209 = ~po52  & n6207;
  assign n6210 = ~n5871 & ~n5872;
  assign n6211 = po28  & n6210;
  assign n6212 = ~n5877 & ~n6211;
  assign n6213 = n5877 & n6211;
  assign n6214 = ~n6212 & ~n6213;
  assign n6215 = ~n6209 & ~n6214;
  assign n6216 = ~n6208 & ~n6215;
  assign n6217 = po53  & ~n6216;
  assign n6218 = ~po53  & n6216;
  assign n6219 = ~n5880 & ~n5881;
  assign n6220 = po28  & n6219;
  assign n6221 = ~n5886 & ~n6220;
  assign n6222 = n5886 & n6220;
  assign n6223 = ~n6221 & ~n6222;
  assign n6224 = ~n6218 & ~n6223;
  assign n6225 = ~n6217 & ~n6224;
  assign n6226 = po54  & ~n6225;
  assign n6227 = ~po54  & n6225;
  assign n6228 = ~n5889 & ~n5890;
  assign n6229 = po28  & n6228;
  assign n6230 = ~n5895 & ~n6229;
  assign n6231 = n5895 & n6229;
  assign n6232 = ~n6230 & ~n6231;
  assign n6233 = ~n6227 & ~n6232;
  assign n6234 = ~n6226 & ~n6233;
  assign n6235 = po55  & ~n6234;
  assign n6236 = ~po55  & n6234;
  assign n6237 = ~n5898 & ~n5899;
  assign n6238 = po28  & n6237;
  assign n6239 = ~n5904 & ~n6238;
  assign n6240 = n5904 & n6238;
  assign n6241 = ~n6239 & ~n6240;
  assign n6242 = ~n6236 & ~n6241;
  assign n6243 = ~n6235 & ~n6242;
  assign n6244 = po56  & ~n6243;
  assign n6245 = ~po56  & n6243;
  assign n6246 = ~n5907 & ~n5908;
  assign n6247 = po28  & n6246;
  assign n6248 = ~n5913 & ~n6247;
  assign n6249 = n5913 & n6247;
  assign n6250 = ~n6248 & ~n6249;
  assign n6251 = ~n6245 & ~n6250;
  assign n6252 = ~n6244 & ~n6251;
  assign n6253 = po57  & ~n6252;
  assign n6254 = ~po57  & n6252;
  assign n6255 = ~n5916 & ~n5917;
  assign n6256 = po28  & n6255;
  assign n6257 = ~n5922 & ~n6256;
  assign n6258 = n5922 & n6256;
  assign n6259 = ~n6257 & ~n6258;
  assign n6260 = ~n6254 & ~n6259;
  assign n6261 = ~n6253 & ~n6260;
  assign n6262 = po58  & ~n6261;
  assign n6263 = ~po58  & n6261;
  assign n6264 = ~n5925 & ~n5926;
  assign n6265 = po28  & n6264;
  assign n6266 = ~n5931 & ~n6265;
  assign n6267 = n5931 & n6265;
  assign n6268 = ~n6266 & ~n6267;
  assign n6269 = ~n6263 & ~n6268;
  assign n6270 = ~n6262 & ~n6269;
  assign n6271 = po59  & ~n6270;
  assign n6272 = ~po59  & n6270;
  assign n6273 = ~n5934 & ~n5935;
  assign n6274 = po28  & n6273;
  assign n6275 = ~n5940 & ~n6274;
  assign n6276 = n5940 & n6274;
  assign n6277 = ~n6275 & ~n6276;
  assign n6278 = ~n6272 & ~n6277;
  assign n6279 = ~n6271 & ~n6278;
  assign n6280 = po60  & ~n6279;
  assign n6281 = ~po60  & n6279;
  assign n6282 = ~n5943 & ~n5944;
  assign n6283 = po28  & n6282;
  assign n6284 = ~n5949 & ~n6283;
  assign n6285 = n5949 & n6283;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = ~n6281 & ~n6286;
  assign n6288 = ~n6280 & ~n6287;
  assign n6289 = po61  & ~n6288;
  assign n6290 = ~po61  & n6288;
  assign n6291 = ~n5952 & ~n5953;
  assign n6292 = po28  & n6291;
  assign n6293 = ~n5958 & ~n6292;
  assign n6294 = n5958 & n6292;
  assign n6295 = ~n6293 & ~n6294;
  assign n6296 = ~n6290 & ~n6295;
  assign n6297 = ~n6289 & ~n6296;
  assign n6298 = po62  & ~n6297;
  assign n6299 = ~po62  & n6297;
  assign n6300 = ~n5961 & ~n5962;
  assign n6301 = po28  & n6300;
  assign n6302 = ~n5967 & ~n6301;
  assign n6303 = n5967 & n6301;
  assign n6304 = ~n6302 & ~n6303;
  assign n6305 = ~n6299 & ~n6304;
  assign n6306 = ~n6298 & ~n6305;
  assign n6307 = n6002 & n6306;
  assign n6308 = ~n6002 & ~n6306;
  assign n6309 = n5980 & po28 ;
  assign n6310 = ~n5979 & ~n6309;
  assign n6311 = n6308 & n6310;
  assign n6312 = ~po63  & ~n6311;
  assign n6313 = ~n6307 & ~n6312;
  assign n6314 = ~n5997 & n6313;
  assign po27  = n5993 | ~n6314;
  assign n6316 = ~n6078 & ~n6079;
  assign n6317 = po27  & n6316;
  assign n6318 = ~n5992 & ~n6317;
  assign n6319 = n5992 & n6317;
  assign n6320 = ~n6318 & ~n6319;
  assign n6321 = n6002 & ~po27 ;
  assign n6322 = ~n6002 & po27 ;
  assign n6323 = n6306 & ~n6322;
  assign n6324 = po63  & ~n6323;
  assign n6325 = ~n6308 & n6324;
  assign n6326 = ~n6298 & ~n6299;
  assign n6327 = po27  & n6326;
  assign n6328 = ~n6304 & ~n6327;
  assign n6329 = n6304 & n6327;
  assign n6330 = ~n6328 & ~n6329;
  assign n6331 = pi54  & po27 ;
  assign n6332 = ~pi52  & ~pi53 ;
  assign n6333 = ~pi54  & n6332;
  assign n6334 = ~n6331 & ~n6333;
  assign n6335 = po28  & ~n6334;
  assign n6336 = ~po28  & n6334;
  assign n6337 = ~pi54  & po27 ;
  assign n6338 = pi55  & ~n6337;
  assign n6339 = n6004 & po27 ;
  assign n6340 = ~n6338 & ~n6339;
  assign n6341 = ~n6336 & n6340;
  assign n6342 = ~n6335 & ~n6341;
  assign n6343 = po29  & ~n6342;
  assign n6344 = ~po29  & n6342;
  assign n6345 = po28  & n6314;
  assign n6346 = ~n6339 & ~n6345;
  assign n6347 = pi56  & ~n6346;
  assign n6348 = ~pi56  & n6346;
  assign n6349 = ~n6347 & ~n6348;
  assign n6350 = ~n6344 & ~n6349;
  assign n6351 = ~n6343 & ~n6350;
  assign n6352 = po30  & ~n6351;
  assign n6353 = ~po30  & n6351;
  assign n6354 = ~n6007 & ~n6008;
  assign n6355 = po27  & n6354;
  assign n6356 = n6012 & ~n6355;
  assign n6357 = ~n6012 & n6355;
  assign n6358 = ~n6356 & ~n6357;
  assign n6359 = ~n6353 & ~n6358;
  assign n6360 = ~n6352 & ~n6359;
  assign n6361 = po31  & ~n6360;
  assign n6362 = ~po31  & n6360;
  assign n6363 = ~n6015 & ~n6016;
  assign n6364 = po27  & n6363;
  assign n6365 = ~n6021 & ~n6364;
  assign n6366 = n6021 & n6364;
  assign n6367 = ~n6365 & ~n6366;
  assign n6368 = ~n6362 & ~n6367;
  assign n6369 = ~n6361 & ~n6368;
  assign n6370 = po32  & ~n6369;
  assign n6371 = ~po32  & n6369;
  assign n6372 = ~n6024 & ~n6025;
  assign n6373 = po27  & n6372;
  assign n6374 = n6030 & n6373;
  assign n6375 = ~n6030 & ~n6373;
  assign n6376 = ~n6374 & ~n6375;
  assign n6377 = ~n6371 & ~n6376;
  assign n6378 = ~n6370 & ~n6377;
  assign n6379 = po33  & ~n6378;
  assign n6380 = ~po33  & n6378;
  assign n6381 = ~n6033 & ~n6034;
  assign n6382 = po27  & n6381;
  assign n6383 = ~n6039 & ~n6382;
  assign n6384 = n6039 & n6382;
  assign n6385 = ~n6383 & ~n6384;
  assign n6386 = ~n6380 & ~n6385;
  assign n6387 = ~n6379 & ~n6386;
  assign n6388 = po34  & ~n6387;
  assign n6389 = ~po34  & n6387;
  assign n6390 = ~n6042 & ~n6043;
  assign n6391 = po27  & n6390;
  assign n6392 = ~n6048 & ~n6391;
  assign n6393 = n6048 & n6391;
  assign n6394 = ~n6392 & ~n6393;
  assign n6395 = ~n6389 & ~n6394;
  assign n6396 = ~n6388 & ~n6395;
  assign n6397 = po35  & ~n6396;
  assign n6398 = ~po35  & n6396;
  assign n6399 = ~n6051 & ~n6052;
  assign n6400 = po27  & n6399;
  assign n6401 = ~n6057 & ~n6400;
  assign n6402 = n6057 & n6400;
  assign n6403 = ~n6401 & ~n6402;
  assign n6404 = ~n6398 & ~n6403;
  assign n6405 = ~n6397 & ~n6404;
  assign n6406 = po36  & ~n6405;
  assign n6407 = ~po36  & n6405;
  assign n6408 = ~n6060 & ~n6061;
  assign n6409 = po27  & n6408;
  assign n6410 = ~n6066 & ~n6409;
  assign n6411 = n6066 & n6409;
  assign n6412 = ~n6410 & ~n6411;
  assign n6413 = ~n6407 & ~n6412;
  assign n6414 = ~n6406 & ~n6413;
  assign n6415 = po37  & ~n6414;
  assign n6416 = ~n6069 & ~n6075;
  assign n6417 = po27  & n6416;
  assign n6418 = ~n6074 & ~n6417;
  assign n6419 = n6074 & n6417;
  assign n6420 = ~n6418 & ~n6419;
  assign n6421 = ~po37  & n6414;
  assign n6422 = ~n6420 & ~n6421;
  assign n6423 = ~n6415 & ~n6422;
  assign n6424 = po38  & ~n6423;
  assign n6425 = ~po38  & n6423;
  assign n6426 = ~n6320 & ~n6425;
  assign n6427 = ~n6424 & ~n6426;
  assign n6428 = po39  & ~n6427;
  assign n6429 = ~po39  & n6427;
  assign n6430 = ~n6082 & ~n6083;
  assign n6431 = po27  & n6430;
  assign n6432 = ~n6088 & ~n6431;
  assign n6433 = n6088 & n6431;
  assign n6434 = ~n6432 & ~n6433;
  assign n6435 = ~n6429 & ~n6434;
  assign n6436 = ~n6428 & ~n6435;
  assign n6437 = po40  & ~n6436;
  assign n6438 = ~po40  & n6436;
  assign n6439 = ~n6091 & ~n6092;
  assign n6440 = po27  & n6439;
  assign n6441 = ~n6097 & ~n6440;
  assign n6442 = n6097 & n6440;
  assign n6443 = ~n6441 & ~n6442;
  assign n6444 = ~n6438 & ~n6443;
  assign n6445 = ~n6437 & ~n6444;
  assign n6446 = po41  & ~n6445;
  assign n6447 = ~po41  & n6445;
  assign n6448 = ~n6100 & ~n6101;
  assign n6449 = po27  & n6448;
  assign n6450 = ~n6106 & ~n6449;
  assign n6451 = n6106 & n6449;
  assign n6452 = ~n6450 & ~n6451;
  assign n6453 = ~n6447 & ~n6452;
  assign n6454 = ~n6446 & ~n6453;
  assign n6455 = po42  & ~n6454;
  assign n6456 = ~po42  & n6454;
  assign n6457 = ~n6109 & ~n6110;
  assign n6458 = po27  & n6457;
  assign n6459 = ~n6115 & ~n6458;
  assign n6460 = n6115 & n6458;
  assign n6461 = ~n6459 & ~n6460;
  assign n6462 = ~n6456 & ~n6461;
  assign n6463 = ~n6455 & ~n6462;
  assign n6464 = po43  & ~n6463;
  assign n6465 = ~po43  & n6463;
  assign n6466 = ~n6118 & ~n6119;
  assign n6467 = po27  & n6466;
  assign n6468 = ~n6124 & ~n6467;
  assign n6469 = n6124 & n6467;
  assign n6470 = ~n6468 & ~n6469;
  assign n6471 = ~n6465 & ~n6470;
  assign n6472 = ~n6464 & ~n6471;
  assign n6473 = po44  & ~n6472;
  assign n6474 = ~po44  & n6472;
  assign n6475 = ~n6127 & ~n6128;
  assign n6476 = po27  & n6475;
  assign n6477 = ~n6133 & ~n6476;
  assign n6478 = n6133 & n6476;
  assign n6479 = ~n6477 & ~n6478;
  assign n6480 = ~n6474 & ~n6479;
  assign n6481 = ~n6473 & ~n6480;
  assign n6482 = po45  & ~n6481;
  assign n6483 = ~po45  & n6481;
  assign n6484 = ~n6136 & ~n6137;
  assign n6485 = po27  & n6484;
  assign n6486 = ~n6142 & ~n6485;
  assign n6487 = n6142 & n6485;
  assign n6488 = ~n6486 & ~n6487;
  assign n6489 = ~n6483 & ~n6488;
  assign n6490 = ~n6482 & ~n6489;
  assign n6491 = po46  & ~n6490;
  assign n6492 = ~po46  & n6490;
  assign n6493 = ~n6145 & ~n6146;
  assign n6494 = po27  & n6493;
  assign n6495 = ~n6151 & ~n6494;
  assign n6496 = n6151 & n6494;
  assign n6497 = ~n6495 & ~n6496;
  assign n6498 = ~n6492 & ~n6497;
  assign n6499 = ~n6491 & ~n6498;
  assign n6500 = po47  & ~n6499;
  assign n6501 = ~po47  & n6499;
  assign n6502 = ~n6154 & ~n6155;
  assign n6503 = po27  & n6502;
  assign n6504 = ~n6160 & ~n6503;
  assign n6505 = n6160 & n6503;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = ~n6501 & ~n6506;
  assign n6508 = ~n6500 & ~n6507;
  assign n6509 = po48  & ~n6508;
  assign n6510 = ~po48  & n6508;
  assign n6511 = ~n6163 & ~n6164;
  assign n6512 = po27  & n6511;
  assign n6513 = ~n6169 & ~n6512;
  assign n6514 = n6169 & n6512;
  assign n6515 = ~n6513 & ~n6514;
  assign n6516 = ~n6510 & ~n6515;
  assign n6517 = ~n6509 & ~n6516;
  assign n6518 = po49  & ~n6517;
  assign n6519 = ~po49  & n6517;
  assign n6520 = ~n6172 & ~n6173;
  assign n6521 = po27  & n6520;
  assign n6522 = ~n6178 & ~n6521;
  assign n6523 = n6178 & n6521;
  assign n6524 = ~n6522 & ~n6523;
  assign n6525 = ~n6519 & ~n6524;
  assign n6526 = ~n6518 & ~n6525;
  assign n6527 = po50  & ~n6526;
  assign n6528 = ~po50  & n6526;
  assign n6529 = ~n6181 & ~n6182;
  assign n6530 = po27  & n6529;
  assign n6531 = ~n6187 & ~n6530;
  assign n6532 = n6187 & n6530;
  assign n6533 = ~n6531 & ~n6532;
  assign n6534 = ~n6528 & ~n6533;
  assign n6535 = ~n6527 & ~n6534;
  assign n6536 = po51  & ~n6535;
  assign n6537 = ~po51  & n6535;
  assign n6538 = ~n6190 & ~n6191;
  assign n6539 = po27  & n6538;
  assign n6540 = ~n6196 & ~n6539;
  assign n6541 = n6196 & n6539;
  assign n6542 = ~n6540 & ~n6541;
  assign n6543 = ~n6537 & ~n6542;
  assign n6544 = ~n6536 & ~n6543;
  assign n6545 = po52  & ~n6544;
  assign n6546 = ~po52  & n6544;
  assign n6547 = ~n6199 & ~n6200;
  assign n6548 = po27  & n6547;
  assign n6549 = ~n6205 & ~n6548;
  assign n6550 = n6205 & n6548;
  assign n6551 = ~n6549 & ~n6550;
  assign n6552 = ~n6546 & ~n6551;
  assign n6553 = ~n6545 & ~n6552;
  assign n6554 = po53  & ~n6553;
  assign n6555 = ~po53  & n6553;
  assign n6556 = ~n6208 & ~n6209;
  assign n6557 = po27  & n6556;
  assign n6558 = ~n6214 & ~n6557;
  assign n6559 = n6214 & n6557;
  assign n6560 = ~n6558 & ~n6559;
  assign n6561 = ~n6555 & ~n6560;
  assign n6562 = ~n6554 & ~n6561;
  assign n6563 = po54  & ~n6562;
  assign n6564 = ~po54  & n6562;
  assign n6565 = ~n6217 & ~n6218;
  assign n6566 = po27  & n6565;
  assign n6567 = ~n6223 & ~n6566;
  assign n6568 = n6223 & n6566;
  assign n6569 = ~n6567 & ~n6568;
  assign n6570 = ~n6564 & ~n6569;
  assign n6571 = ~n6563 & ~n6570;
  assign n6572 = po55  & ~n6571;
  assign n6573 = ~po55  & n6571;
  assign n6574 = ~n6226 & ~n6227;
  assign n6575 = po27  & n6574;
  assign n6576 = ~n6232 & ~n6575;
  assign n6577 = n6232 & n6575;
  assign n6578 = ~n6576 & ~n6577;
  assign n6579 = ~n6573 & ~n6578;
  assign n6580 = ~n6572 & ~n6579;
  assign n6581 = po56  & ~n6580;
  assign n6582 = ~po56  & n6580;
  assign n6583 = ~n6235 & ~n6236;
  assign n6584 = po27  & n6583;
  assign n6585 = ~n6241 & ~n6584;
  assign n6586 = n6241 & n6584;
  assign n6587 = ~n6585 & ~n6586;
  assign n6588 = ~n6582 & ~n6587;
  assign n6589 = ~n6581 & ~n6588;
  assign n6590 = po57  & ~n6589;
  assign n6591 = ~po57  & n6589;
  assign n6592 = ~n6244 & ~n6245;
  assign n6593 = po27  & n6592;
  assign n6594 = ~n6250 & ~n6593;
  assign n6595 = n6250 & n6593;
  assign n6596 = ~n6594 & ~n6595;
  assign n6597 = ~n6591 & ~n6596;
  assign n6598 = ~n6590 & ~n6597;
  assign n6599 = po58  & ~n6598;
  assign n6600 = ~po58  & n6598;
  assign n6601 = ~n6253 & ~n6254;
  assign n6602 = po27  & n6601;
  assign n6603 = ~n6259 & ~n6602;
  assign n6604 = n6259 & n6602;
  assign n6605 = ~n6603 & ~n6604;
  assign n6606 = ~n6600 & ~n6605;
  assign n6607 = ~n6599 & ~n6606;
  assign n6608 = po59  & ~n6607;
  assign n6609 = ~po59  & n6607;
  assign n6610 = ~n6262 & ~n6263;
  assign n6611 = po27  & n6610;
  assign n6612 = ~n6268 & ~n6611;
  assign n6613 = n6268 & n6611;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = ~n6609 & ~n6614;
  assign n6616 = ~n6608 & ~n6615;
  assign n6617 = po60  & ~n6616;
  assign n6618 = ~po60  & n6616;
  assign n6619 = ~n6271 & ~n6272;
  assign n6620 = po27  & n6619;
  assign n6621 = ~n6277 & ~n6620;
  assign n6622 = n6277 & n6620;
  assign n6623 = ~n6621 & ~n6622;
  assign n6624 = ~n6618 & ~n6623;
  assign n6625 = ~n6617 & ~n6624;
  assign n6626 = po61  & ~n6625;
  assign n6627 = ~po61  & n6625;
  assign n6628 = ~n6280 & ~n6281;
  assign n6629 = po27  & n6628;
  assign n6630 = ~n6286 & ~n6629;
  assign n6631 = n6286 & n6629;
  assign n6632 = ~n6630 & ~n6631;
  assign n6633 = ~n6627 & ~n6632;
  assign n6634 = ~n6626 & ~n6633;
  assign n6635 = po62  & ~n6634;
  assign n6636 = ~po62  & n6634;
  assign n6637 = ~n6289 & ~n6290;
  assign n6638 = po27  & n6637;
  assign n6639 = ~n6295 & ~n6638;
  assign n6640 = n6295 & n6638;
  assign n6641 = ~n6639 & ~n6640;
  assign n6642 = ~n6636 & ~n6641;
  assign n6643 = ~n6635 & ~n6642;
  assign n6644 = n6330 & n6643;
  assign n6645 = ~n6330 & ~n6643;
  assign n6646 = n6308 & po27 ;
  assign n6647 = ~n6307 & ~n6646;
  assign n6648 = n6645 & n6647;
  assign n6649 = ~po63  & ~n6648;
  assign n6650 = ~n6644 & ~n6649;
  assign n6651 = ~n6325 & n6650;
  assign po26  = n6321 | ~n6651;
  assign n6653 = ~n6424 & ~n6425;
  assign n6654 = po26  & n6653;
  assign n6655 = ~n6320 & ~n6654;
  assign n6656 = n6320 & n6654;
  assign n6657 = ~n6655 & ~n6656;
  assign n6658 = n6330 & ~po26 ;
  assign n6659 = ~n6330 & po26 ;
  assign n6660 = n6643 & ~n6659;
  assign n6661 = po63  & ~n6660;
  assign n6662 = ~n6645 & n6661;
  assign n6663 = ~n6635 & ~n6636;
  assign n6664 = po26  & n6663;
  assign n6665 = ~n6641 & ~n6664;
  assign n6666 = n6641 & n6664;
  assign n6667 = ~n6665 & ~n6666;
  assign n6668 = pi52  & po26 ;
  assign n6669 = ~pi50  & ~pi51 ;
  assign n6670 = ~pi52  & n6669;
  assign n6671 = ~n6668 & ~n6670;
  assign n6672 = po27  & ~n6671;
  assign n6673 = ~po27  & n6671;
  assign n6674 = ~pi52  & po26 ;
  assign n6675 = pi53  & ~n6674;
  assign n6676 = n6332 & po26 ;
  assign n6677 = ~n6675 & ~n6676;
  assign n6678 = ~n6673 & n6677;
  assign n6679 = ~n6672 & ~n6678;
  assign n6680 = po28  & ~n6679;
  assign n6681 = ~po28  & n6679;
  assign n6682 = po27  & n6651;
  assign n6683 = ~n6676 & ~n6682;
  assign n6684 = pi54  & ~n6683;
  assign n6685 = ~pi54  & n6683;
  assign n6686 = ~n6684 & ~n6685;
  assign n6687 = ~n6681 & ~n6686;
  assign n6688 = ~n6680 & ~n6687;
  assign n6689 = po29  & ~n6688;
  assign n6690 = ~po29  & n6688;
  assign n6691 = ~n6335 & ~n6336;
  assign n6692 = po26  & n6691;
  assign n6693 = n6340 & ~n6692;
  assign n6694 = ~n6340 & n6692;
  assign n6695 = ~n6693 & ~n6694;
  assign n6696 = ~n6690 & ~n6695;
  assign n6697 = ~n6689 & ~n6696;
  assign n6698 = po30  & ~n6697;
  assign n6699 = ~po30  & n6697;
  assign n6700 = ~n6343 & ~n6344;
  assign n6701 = po26  & n6700;
  assign n6702 = ~n6349 & ~n6701;
  assign n6703 = n6349 & n6701;
  assign n6704 = ~n6702 & ~n6703;
  assign n6705 = ~n6699 & ~n6704;
  assign n6706 = ~n6698 & ~n6705;
  assign n6707 = po31  & ~n6706;
  assign n6708 = ~po31  & n6706;
  assign n6709 = ~n6352 & ~n6353;
  assign n6710 = po26  & n6709;
  assign n6711 = n6358 & n6710;
  assign n6712 = ~n6358 & ~n6710;
  assign n6713 = ~n6711 & ~n6712;
  assign n6714 = ~n6708 & ~n6713;
  assign n6715 = ~n6707 & ~n6714;
  assign n6716 = po32  & ~n6715;
  assign n6717 = ~po32  & n6715;
  assign n6718 = ~n6361 & ~n6362;
  assign n6719 = po26  & n6718;
  assign n6720 = ~n6367 & ~n6719;
  assign n6721 = n6367 & n6719;
  assign n6722 = ~n6720 & ~n6721;
  assign n6723 = ~n6717 & ~n6722;
  assign n6724 = ~n6716 & ~n6723;
  assign n6725 = po33  & ~n6724;
  assign n6726 = ~po33  & n6724;
  assign n6727 = ~n6370 & ~n6371;
  assign n6728 = po26  & n6727;
  assign n6729 = ~n6376 & ~n6728;
  assign n6730 = n6376 & n6728;
  assign n6731 = ~n6729 & ~n6730;
  assign n6732 = ~n6726 & ~n6731;
  assign n6733 = ~n6725 & ~n6732;
  assign n6734 = po34  & ~n6733;
  assign n6735 = ~po34  & n6733;
  assign n6736 = ~n6379 & ~n6380;
  assign n6737 = po26  & n6736;
  assign n6738 = ~n6385 & ~n6737;
  assign n6739 = n6385 & n6737;
  assign n6740 = ~n6738 & ~n6739;
  assign n6741 = ~n6735 & ~n6740;
  assign n6742 = ~n6734 & ~n6741;
  assign n6743 = po35  & ~n6742;
  assign n6744 = ~po35  & n6742;
  assign n6745 = ~n6388 & ~n6389;
  assign n6746 = po26  & n6745;
  assign n6747 = ~n6394 & ~n6746;
  assign n6748 = n6394 & n6746;
  assign n6749 = ~n6747 & ~n6748;
  assign n6750 = ~n6744 & ~n6749;
  assign n6751 = ~n6743 & ~n6750;
  assign n6752 = po36  & ~n6751;
  assign n6753 = ~po36  & n6751;
  assign n6754 = ~n6397 & ~n6398;
  assign n6755 = po26  & n6754;
  assign n6756 = ~n6403 & ~n6755;
  assign n6757 = n6403 & n6755;
  assign n6758 = ~n6756 & ~n6757;
  assign n6759 = ~n6753 & ~n6758;
  assign n6760 = ~n6752 & ~n6759;
  assign n6761 = po37  & ~n6760;
  assign n6762 = ~po37  & n6760;
  assign n6763 = ~n6406 & ~n6407;
  assign n6764 = po26  & n6763;
  assign n6765 = ~n6412 & ~n6764;
  assign n6766 = n6412 & n6764;
  assign n6767 = ~n6765 & ~n6766;
  assign n6768 = ~n6762 & ~n6767;
  assign n6769 = ~n6761 & ~n6768;
  assign n6770 = po38  & ~n6769;
  assign n6771 = ~n6415 & ~n6421;
  assign n6772 = po26  & n6771;
  assign n6773 = ~n6420 & ~n6772;
  assign n6774 = n6420 & n6772;
  assign n6775 = ~n6773 & ~n6774;
  assign n6776 = ~po38  & n6769;
  assign n6777 = ~n6775 & ~n6776;
  assign n6778 = ~n6770 & ~n6777;
  assign n6779 = po39  & ~n6778;
  assign n6780 = ~po39  & n6778;
  assign n6781 = ~n6657 & ~n6780;
  assign n6782 = ~n6779 & ~n6781;
  assign n6783 = po40  & ~n6782;
  assign n6784 = ~po40  & n6782;
  assign n6785 = ~n6428 & ~n6429;
  assign n6786 = po26  & n6785;
  assign n6787 = ~n6434 & ~n6786;
  assign n6788 = n6434 & n6786;
  assign n6789 = ~n6787 & ~n6788;
  assign n6790 = ~n6784 & ~n6789;
  assign n6791 = ~n6783 & ~n6790;
  assign n6792 = po41  & ~n6791;
  assign n6793 = ~po41  & n6791;
  assign n6794 = ~n6437 & ~n6438;
  assign n6795 = po26  & n6794;
  assign n6796 = ~n6443 & ~n6795;
  assign n6797 = n6443 & n6795;
  assign n6798 = ~n6796 & ~n6797;
  assign n6799 = ~n6793 & ~n6798;
  assign n6800 = ~n6792 & ~n6799;
  assign n6801 = po42  & ~n6800;
  assign n6802 = ~po42  & n6800;
  assign n6803 = ~n6446 & ~n6447;
  assign n6804 = po26  & n6803;
  assign n6805 = ~n6452 & ~n6804;
  assign n6806 = n6452 & n6804;
  assign n6807 = ~n6805 & ~n6806;
  assign n6808 = ~n6802 & ~n6807;
  assign n6809 = ~n6801 & ~n6808;
  assign n6810 = po43  & ~n6809;
  assign n6811 = ~po43  & n6809;
  assign n6812 = ~n6455 & ~n6456;
  assign n6813 = po26  & n6812;
  assign n6814 = ~n6461 & ~n6813;
  assign n6815 = n6461 & n6813;
  assign n6816 = ~n6814 & ~n6815;
  assign n6817 = ~n6811 & ~n6816;
  assign n6818 = ~n6810 & ~n6817;
  assign n6819 = po44  & ~n6818;
  assign n6820 = ~po44  & n6818;
  assign n6821 = ~n6464 & ~n6465;
  assign n6822 = po26  & n6821;
  assign n6823 = ~n6470 & ~n6822;
  assign n6824 = n6470 & n6822;
  assign n6825 = ~n6823 & ~n6824;
  assign n6826 = ~n6820 & ~n6825;
  assign n6827 = ~n6819 & ~n6826;
  assign n6828 = po45  & ~n6827;
  assign n6829 = ~po45  & n6827;
  assign n6830 = ~n6473 & ~n6474;
  assign n6831 = po26  & n6830;
  assign n6832 = ~n6479 & ~n6831;
  assign n6833 = n6479 & n6831;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = ~n6829 & ~n6834;
  assign n6836 = ~n6828 & ~n6835;
  assign n6837 = po46  & ~n6836;
  assign n6838 = ~po46  & n6836;
  assign n6839 = ~n6482 & ~n6483;
  assign n6840 = po26  & n6839;
  assign n6841 = ~n6488 & ~n6840;
  assign n6842 = n6488 & n6840;
  assign n6843 = ~n6841 & ~n6842;
  assign n6844 = ~n6838 & ~n6843;
  assign n6845 = ~n6837 & ~n6844;
  assign n6846 = po47  & ~n6845;
  assign n6847 = ~po47  & n6845;
  assign n6848 = ~n6491 & ~n6492;
  assign n6849 = po26  & n6848;
  assign n6850 = ~n6497 & ~n6849;
  assign n6851 = n6497 & n6849;
  assign n6852 = ~n6850 & ~n6851;
  assign n6853 = ~n6847 & ~n6852;
  assign n6854 = ~n6846 & ~n6853;
  assign n6855 = po48  & ~n6854;
  assign n6856 = ~po48  & n6854;
  assign n6857 = ~n6500 & ~n6501;
  assign n6858 = po26  & n6857;
  assign n6859 = ~n6506 & ~n6858;
  assign n6860 = n6506 & n6858;
  assign n6861 = ~n6859 & ~n6860;
  assign n6862 = ~n6856 & ~n6861;
  assign n6863 = ~n6855 & ~n6862;
  assign n6864 = po49  & ~n6863;
  assign n6865 = ~po49  & n6863;
  assign n6866 = ~n6509 & ~n6510;
  assign n6867 = po26  & n6866;
  assign n6868 = ~n6515 & ~n6867;
  assign n6869 = n6515 & n6867;
  assign n6870 = ~n6868 & ~n6869;
  assign n6871 = ~n6865 & ~n6870;
  assign n6872 = ~n6864 & ~n6871;
  assign n6873 = po50  & ~n6872;
  assign n6874 = ~po50  & n6872;
  assign n6875 = ~n6518 & ~n6519;
  assign n6876 = po26  & n6875;
  assign n6877 = ~n6524 & ~n6876;
  assign n6878 = n6524 & n6876;
  assign n6879 = ~n6877 & ~n6878;
  assign n6880 = ~n6874 & ~n6879;
  assign n6881 = ~n6873 & ~n6880;
  assign n6882 = po51  & ~n6881;
  assign n6883 = ~po51  & n6881;
  assign n6884 = ~n6527 & ~n6528;
  assign n6885 = po26  & n6884;
  assign n6886 = ~n6533 & ~n6885;
  assign n6887 = n6533 & n6885;
  assign n6888 = ~n6886 & ~n6887;
  assign n6889 = ~n6883 & ~n6888;
  assign n6890 = ~n6882 & ~n6889;
  assign n6891 = po52  & ~n6890;
  assign n6892 = ~po52  & n6890;
  assign n6893 = ~n6536 & ~n6537;
  assign n6894 = po26  & n6893;
  assign n6895 = ~n6542 & ~n6894;
  assign n6896 = n6542 & n6894;
  assign n6897 = ~n6895 & ~n6896;
  assign n6898 = ~n6892 & ~n6897;
  assign n6899 = ~n6891 & ~n6898;
  assign n6900 = po53  & ~n6899;
  assign n6901 = ~po53  & n6899;
  assign n6902 = ~n6545 & ~n6546;
  assign n6903 = po26  & n6902;
  assign n6904 = ~n6551 & ~n6903;
  assign n6905 = n6551 & n6903;
  assign n6906 = ~n6904 & ~n6905;
  assign n6907 = ~n6901 & ~n6906;
  assign n6908 = ~n6900 & ~n6907;
  assign n6909 = po54  & ~n6908;
  assign n6910 = ~po54  & n6908;
  assign n6911 = ~n6554 & ~n6555;
  assign n6912 = po26  & n6911;
  assign n6913 = ~n6560 & ~n6912;
  assign n6914 = n6560 & n6912;
  assign n6915 = ~n6913 & ~n6914;
  assign n6916 = ~n6910 & ~n6915;
  assign n6917 = ~n6909 & ~n6916;
  assign n6918 = po55  & ~n6917;
  assign n6919 = ~po55  & n6917;
  assign n6920 = ~n6563 & ~n6564;
  assign n6921 = po26  & n6920;
  assign n6922 = ~n6569 & ~n6921;
  assign n6923 = n6569 & n6921;
  assign n6924 = ~n6922 & ~n6923;
  assign n6925 = ~n6919 & ~n6924;
  assign n6926 = ~n6918 & ~n6925;
  assign n6927 = po56  & ~n6926;
  assign n6928 = ~po56  & n6926;
  assign n6929 = ~n6572 & ~n6573;
  assign n6930 = po26  & n6929;
  assign n6931 = ~n6578 & ~n6930;
  assign n6932 = n6578 & n6930;
  assign n6933 = ~n6931 & ~n6932;
  assign n6934 = ~n6928 & ~n6933;
  assign n6935 = ~n6927 & ~n6934;
  assign n6936 = po57  & ~n6935;
  assign n6937 = ~po57  & n6935;
  assign n6938 = ~n6581 & ~n6582;
  assign n6939 = po26  & n6938;
  assign n6940 = ~n6587 & ~n6939;
  assign n6941 = n6587 & n6939;
  assign n6942 = ~n6940 & ~n6941;
  assign n6943 = ~n6937 & ~n6942;
  assign n6944 = ~n6936 & ~n6943;
  assign n6945 = po58  & ~n6944;
  assign n6946 = ~po58  & n6944;
  assign n6947 = ~n6590 & ~n6591;
  assign n6948 = po26  & n6947;
  assign n6949 = ~n6596 & ~n6948;
  assign n6950 = n6596 & n6948;
  assign n6951 = ~n6949 & ~n6950;
  assign n6952 = ~n6946 & ~n6951;
  assign n6953 = ~n6945 & ~n6952;
  assign n6954 = po59  & ~n6953;
  assign n6955 = ~po59  & n6953;
  assign n6956 = ~n6599 & ~n6600;
  assign n6957 = po26  & n6956;
  assign n6958 = ~n6605 & ~n6957;
  assign n6959 = n6605 & n6957;
  assign n6960 = ~n6958 & ~n6959;
  assign n6961 = ~n6955 & ~n6960;
  assign n6962 = ~n6954 & ~n6961;
  assign n6963 = po60  & ~n6962;
  assign n6964 = ~po60  & n6962;
  assign n6965 = ~n6608 & ~n6609;
  assign n6966 = po26  & n6965;
  assign n6967 = ~n6614 & ~n6966;
  assign n6968 = n6614 & n6966;
  assign n6969 = ~n6967 & ~n6968;
  assign n6970 = ~n6964 & ~n6969;
  assign n6971 = ~n6963 & ~n6970;
  assign n6972 = po61  & ~n6971;
  assign n6973 = ~po61  & n6971;
  assign n6974 = ~n6617 & ~n6618;
  assign n6975 = po26  & n6974;
  assign n6976 = ~n6623 & ~n6975;
  assign n6977 = n6623 & n6975;
  assign n6978 = ~n6976 & ~n6977;
  assign n6979 = ~n6973 & ~n6978;
  assign n6980 = ~n6972 & ~n6979;
  assign n6981 = po62  & ~n6980;
  assign n6982 = ~po62  & n6980;
  assign n6983 = ~n6626 & ~n6627;
  assign n6984 = po26  & n6983;
  assign n6985 = ~n6632 & ~n6984;
  assign n6986 = n6632 & n6984;
  assign n6987 = ~n6985 & ~n6986;
  assign n6988 = ~n6982 & ~n6987;
  assign n6989 = ~n6981 & ~n6988;
  assign n6990 = n6667 & n6989;
  assign n6991 = ~n6667 & ~n6989;
  assign n6992 = n6645 & po26 ;
  assign n6993 = ~n6644 & ~n6992;
  assign n6994 = n6991 & n6993;
  assign n6995 = ~po63  & ~n6994;
  assign n6996 = ~n6990 & ~n6995;
  assign n6997 = ~n6662 & n6996;
  assign po25  = n6658 | ~n6997;
  assign n6999 = ~n6779 & ~n6780;
  assign n7000 = po25  & n6999;
  assign n7001 = ~n6657 & ~n7000;
  assign n7002 = n6657 & n7000;
  assign n7003 = ~n7001 & ~n7002;
  assign n7004 = n6667 & ~po25 ;
  assign n7005 = ~n6667 & po25 ;
  assign n7006 = n6989 & ~n7005;
  assign n7007 = po63  & ~n7006;
  assign n7008 = ~n6991 & n7007;
  assign n7009 = ~n6981 & ~n6982;
  assign n7010 = po25  & n7009;
  assign n7011 = ~n6987 & ~n7010;
  assign n7012 = n6987 & n7010;
  assign n7013 = ~n7011 & ~n7012;
  assign n7014 = pi50  & po25 ;
  assign n7015 = ~pi48  & ~pi49 ;
  assign n7016 = ~pi50  & n7015;
  assign n7017 = ~n7014 & ~n7016;
  assign n7018 = po26  & ~n7017;
  assign n7019 = ~po26  & n7017;
  assign n7020 = ~pi50  & po25 ;
  assign n7021 = pi51  & ~n7020;
  assign n7022 = n6669 & po25 ;
  assign n7023 = ~n7021 & ~n7022;
  assign n7024 = ~n7019 & n7023;
  assign n7025 = ~n7018 & ~n7024;
  assign n7026 = po27  & ~n7025;
  assign n7027 = ~po27  & n7025;
  assign n7028 = po26  & n6997;
  assign n7029 = ~n7022 & ~n7028;
  assign n7030 = pi52  & ~n7029;
  assign n7031 = ~pi52  & n7029;
  assign n7032 = ~n7030 & ~n7031;
  assign n7033 = ~n7027 & ~n7032;
  assign n7034 = ~n7026 & ~n7033;
  assign n7035 = po28  & ~n7034;
  assign n7036 = ~po28  & n7034;
  assign n7037 = ~n6672 & ~n6673;
  assign n7038 = po25  & n7037;
  assign n7039 = n6677 & ~n7038;
  assign n7040 = ~n6677 & n7038;
  assign n7041 = ~n7039 & ~n7040;
  assign n7042 = ~n7036 & ~n7041;
  assign n7043 = ~n7035 & ~n7042;
  assign n7044 = po29  & ~n7043;
  assign n7045 = ~po29  & n7043;
  assign n7046 = ~n6680 & ~n6681;
  assign n7047 = po25  & n7046;
  assign n7048 = ~n6686 & ~n7047;
  assign n7049 = n6686 & n7047;
  assign n7050 = ~n7048 & ~n7049;
  assign n7051 = ~n7045 & ~n7050;
  assign n7052 = ~n7044 & ~n7051;
  assign n7053 = po30  & ~n7052;
  assign n7054 = ~po30  & n7052;
  assign n7055 = ~n6689 & ~n6690;
  assign n7056 = po25  & n7055;
  assign n7057 = n6695 & n7056;
  assign n7058 = ~n6695 & ~n7056;
  assign n7059 = ~n7057 & ~n7058;
  assign n7060 = ~n7054 & ~n7059;
  assign n7061 = ~n7053 & ~n7060;
  assign n7062 = po31  & ~n7061;
  assign n7063 = ~po31  & n7061;
  assign n7064 = ~n6698 & ~n6699;
  assign n7065 = po25  & n7064;
  assign n7066 = ~n6704 & ~n7065;
  assign n7067 = n6704 & n7065;
  assign n7068 = ~n7066 & ~n7067;
  assign n7069 = ~n7063 & ~n7068;
  assign n7070 = ~n7062 & ~n7069;
  assign n7071 = po32  & ~n7070;
  assign n7072 = ~po32  & n7070;
  assign n7073 = ~n6707 & ~n6708;
  assign n7074 = po25  & n7073;
  assign n7075 = ~n6713 & ~n7074;
  assign n7076 = n6713 & n7074;
  assign n7077 = ~n7075 & ~n7076;
  assign n7078 = ~n7072 & ~n7077;
  assign n7079 = ~n7071 & ~n7078;
  assign n7080 = po33  & ~n7079;
  assign n7081 = ~po33  & n7079;
  assign n7082 = ~n6716 & ~n6717;
  assign n7083 = po25  & n7082;
  assign n7084 = ~n6722 & ~n7083;
  assign n7085 = n6722 & n7083;
  assign n7086 = ~n7084 & ~n7085;
  assign n7087 = ~n7081 & ~n7086;
  assign n7088 = ~n7080 & ~n7087;
  assign n7089 = po34  & ~n7088;
  assign n7090 = ~po34  & n7088;
  assign n7091 = ~n6725 & ~n6726;
  assign n7092 = po25  & n7091;
  assign n7093 = ~n6731 & ~n7092;
  assign n7094 = n6731 & n7092;
  assign n7095 = ~n7093 & ~n7094;
  assign n7096 = ~n7090 & ~n7095;
  assign n7097 = ~n7089 & ~n7096;
  assign n7098 = po35  & ~n7097;
  assign n7099 = ~po35  & n7097;
  assign n7100 = ~n6734 & ~n6735;
  assign n7101 = po25  & n7100;
  assign n7102 = ~n6740 & ~n7101;
  assign n7103 = n6740 & n7101;
  assign n7104 = ~n7102 & ~n7103;
  assign n7105 = ~n7099 & ~n7104;
  assign n7106 = ~n7098 & ~n7105;
  assign n7107 = po36  & ~n7106;
  assign n7108 = ~po36  & n7106;
  assign n7109 = ~n6743 & ~n6744;
  assign n7110 = po25  & n7109;
  assign n7111 = ~n6749 & ~n7110;
  assign n7112 = n6749 & n7110;
  assign n7113 = ~n7111 & ~n7112;
  assign n7114 = ~n7108 & ~n7113;
  assign n7115 = ~n7107 & ~n7114;
  assign n7116 = po37  & ~n7115;
  assign n7117 = ~po37  & n7115;
  assign n7118 = ~n6752 & ~n6753;
  assign n7119 = po25  & n7118;
  assign n7120 = ~n6758 & ~n7119;
  assign n7121 = n6758 & n7119;
  assign n7122 = ~n7120 & ~n7121;
  assign n7123 = ~n7117 & ~n7122;
  assign n7124 = ~n7116 & ~n7123;
  assign n7125 = po38  & ~n7124;
  assign n7126 = ~po38  & n7124;
  assign n7127 = ~n6761 & ~n6762;
  assign n7128 = po25  & n7127;
  assign n7129 = ~n6767 & ~n7128;
  assign n7130 = n6767 & n7128;
  assign n7131 = ~n7129 & ~n7130;
  assign n7132 = ~n7126 & ~n7131;
  assign n7133 = ~n7125 & ~n7132;
  assign n7134 = po39  & ~n7133;
  assign n7135 = ~n6770 & ~n6776;
  assign n7136 = po25  & n7135;
  assign n7137 = ~n6775 & ~n7136;
  assign n7138 = n6775 & n7136;
  assign n7139 = ~n7137 & ~n7138;
  assign n7140 = ~po39  & n7133;
  assign n7141 = ~n7139 & ~n7140;
  assign n7142 = ~n7134 & ~n7141;
  assign n7143 = po40  & ~n7142;
  assign n7144 = ~po40  & n7142;
  assign n7145 = ~n7003 & ~n7144;
  assign n7146 = ~n7143 & ~n7145;
  assign n7147 = po41  & ~n7146;
  assign n7148 = ~po41  & n7146;
  assign n7149 = ~n6783 & ~n6784;
  assign n7150 = po25  & n7149;
  assign n7151 = ~n6789 & ~n7150;
  assign n7152 = n6789 & n7150;
  assign n7153 = ~n7151 & ~n7152;
  assign n7154 = ~n7148 & ~n7153;
  assign n7155 = ~n7147 & ~n7154;
  assign n7156 = po42  & ~n7155;
  assign n7157 = ~po42  & n7155;
  assign n7158 = ~n6792 & ~n6793;
  assign n7159 = po25  & n7158;
  assign n7160 = ~n6798 & ~n7159;
  assign n7161 = n6798 & n7159;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = ~n7157 & ~n7162;
  assign n7164 = ~n7156 & ~n7163;
  assign n7165 = po43  & ~n7164;
  assign n7166 = ~po43  & n7164;
  assign n7167 = ~n6801 & ~n6802;
  assign n7168 = po25  & n7167;
  assign n7169 = ~n6807 & ~n7168;
  assign n7170 = n6807 & n7168;
  assign n7171 = ~n7169 & ~n7170;
  assign n7172 = ~n7166 & ~n7171;
  assign n7173 = ~n7165 & ~n7172;
  assign n7174 = po44  & ~n7173;
  assign n7175 = ~po44  & n7173;
  assign n7176 = ~n6810 & ~n6811;
  assign n7177 = po25  & n7176;
  assign n7178 = ~n6816 & ~n7177;
  assign n7179 = n6816 & n7177;
  assign n7180 = ~n7178 & ~n7179;
  assign n7181 = ~n7175 & ~n7180;
  assign n7182 = ~n7174 & ~n7181;
  assign n7183 = po45  & ~n7182;
  assign n7184 = ~po45  & n7182;
  assign n7185 = ~n6819 & ~n6820;
  assign n7186 = po25  & n7185;
  assign n7187 = ~n6825 & ~n7186;
  assign n7188 = n6825 & n7186;
  assign n7189 = ~n7187 & ~n7188;
  assign n7190 = ~n7184 & ~n7189;
  assign n7191 = ~n7183 & ~n7190;
  assign n7192 = po46  & ~n7191;
  assign n7193 = ~po46  & n7191;
  assign n7194 = ~n6828 & ~n6829;
  assign n7195 = po25  & n7194;
  assign n7196 = ~n6834 & ~n7195;
  assign n7197 = n6834 & n7195;
  assign n7198 = ~n7196 & ~n7197;
  assign n7199 = ~n7193 & ~n7198;
  assign n7200 = ~n7192 & ~n7199;
  assign n7201 = po47  & ~n7200;
  assign n7202 = ~po47  & n7200;
  assign n7203 = ~n6837 & ~n6838;
  assign n7204 = po25  & n7203;
  assign n7205 = ~n6843 & ~n7204;
  assign n7206 = n6843 & n7204;
  assign n7207 = ~n7205 & ~n7206;
  assign n7208 = ~n7202 & ~n7207;
  assign n7209 = ~n7201 & ~n7208;
  assign n7210 = po48  & ~n7209;
  assign n7211 = ~po48  & n7209;
  assign n7212 = ~n6846 & ~n6847;
  assign n7213 = po25  & n7212;
  assign n7214 = ~n6852 & ~n7213;
  assign n7215 = n6852 & n7213;
  assign n7216 = ~n7214 & ~n7215;
  assign n7217 = ~n7211 & ~n7216;
  assign n7218 = ~n7210 & ~n7217;
  assign n7219 = po49  & ~n7218;
  assign n7220 = ~po49  & n7218;
  assign n7221 = ~n6855 & ~n6856;
  assign n7222 = po25  & n7221;
  assign n7223 = ~n6861 & ~n7222;
  assign n7224 = n6861 & n7222;
  assign n7225 = ~n7223 & ~n7224;
  assign n7226 = ~n7220 & ~n7225;
  assign n7227 = ~n7219 & ~n7226;
  assign n7228 = po50  & ~n7227;
  assign n7229 = ~po50  & n7227;
  assign n7230 = ~n6864 & ~n6865;
  assign n7231 = po25  & n7230;
  assign n7232 = ~n6870 & ~n7231;
  assign n7233 = n6870 & n7231;
  assign n7234 = ~n7232 & ~n7233;
  assign n7235 = ~n7229 & ~n7234;
  assign n7236 = ~n7228 & ~n7235;
  assign n7237 = po51  & ~n7236;
  assign n7238 = ~po51  & n7236;
  assign n7239 = ~n6873 & ~n6874;
  assign n7240 = po25  & n7239;
  assign n7241 = ~n6879 & ~n7240;
  assign n7242 = n6879 & n7240;
  assign n7243 = ~n7241 & ~n7242;
  assign n7244 = ~n7238 & ~n7243;
  assign n7245 = ~n7237 & ~n7244;
  assign n7246 = po52  & ~n7245;
  assign n7247 = ~po52  & n7245;
  assign n7248 = ~n6882 & ~n6883;
  assign n7249 = po25  & n7248;
  assign n7250 = ~n6888 & ~n7249;
  assign n7251 = n6888 & n7249;
  assign n7252 = ~n7250 & ~n7251;
  assign n7253 = ~n7247 & ~n7252;
  assign n7254 = ~n7246 & ~n7253;
  assign n7255 = po53  & ~n7254;
  assign n7256 = ~po53  & n7254;
  assign n7257 = ~n6891 & ~n6892;
  assign n7258 = po25  & n7257;
  assign n7259 = ~n6897 & ~n7258;
  assign n7260 = n6897 & n7258;
  assign n7261 = ~n7259 & ~n7260;
  assign n7262 = ~n7256 & ~n7261;
  assign n7263 = ~n7255 & ~n7262;
  assign n7264 = po54  & ~n7263;
  assign n7265 = ~po54  & n7263;
  assign n7266 = ~n6900 & ~n6901;
  assign n7267 = po25  & n7266;
  assign n7268 = ~n6906 & ~n7267;
  assign n7269 = n6906 & n7267;
  assign n7270 = ~n7268 & ~n7269;
  assign n7271 = ~n7265 & ~n7270;
  assign n7272 = ~n7264 & ~n7271;
  assign n7273 = po55  & ~n7272;
  assign n7274 = ~po55  & n7272;
  assign n7275 = ~n6909 & ~n6910;
  assign n7276 = po25  & n7275;
  assign n7277 = ~n6915 & ~n7276;
  assign n7278 = n6915 & n7276;
  assign n7279 = ~n7277 & ~n7278;
  assign n7280 = ~n7274 & ~n7279;
  assign n7281 = ~n7273 & ~n7280;
  assign n7282 = po56  & ~n7281;
  assign n7283 = ~po56  & n7281;
  assign n7284 = ~n6918 & ~n6919;
  assign n7285 = po25  & n7284;
  assign n7286 = ~n6924 & ~n7285;
  assign n7287 = n6924 & n7285;
  assign n7288 = ~n7286 & ~n7287;
  assign n7289 = ~n7283 & ~n7288;
  assign n7290 = ~n7282 & ~n7289;
  assign n7291 = po57  & ~n7290;
  assign n7292 = ~po57  & n7290;
  assign n7293 = ~n6927 & ~n6928;
  assign n7294 = po25  & n7293;
  assign n7295 = ~n6933 & ~n7294;
  assign n7296 = n6933 & n7294;
  assign n7297 = ~n7295 & ~n7296;
  assign n7298 = ~n7292 & ~n7297;
  assign n7299 = ~n7291 & ~n7298;
  assign n7300 = po58  & ~n7299;
  assign n7301 = ~po58  & n7299;
  assign n7302 = ~n6936 & ~n6937;
  assign n7303 = po25  & n7302;
  assign n7304 = ~n6942 & ~n7303;
  assign n7305 = n6942 & n7303;
  assign n7306 = ~n7304 & ~n7305;
  assign n7307 = ~n7301 & ~n7306;
  assign n7308 = ~n7300 & ~n7307;
  assign n7309 = po59  & ~n7308;
  assign n7310 = ~po59  & n7308;
  assign n7311 = ~n6945 & ~n6946;
  assign n7312 = po25  & n7311;
  assign n7313 = ~n6951 & ~n7312;
  assign n7314 = n6951 & n7312;
  assign n7315 = ~n7313 & ~n7314;
  assign n7316 = ~n7310 & ~n7315;
  assign n7317 = ~n7309 & ~n7316;
  assign n7318 = po60  & ~n7317;
  assign n7319 = ~po60  & n7317;
  assign n7320 = ~n6954 & ~n6955;
  assign n7321 = po25  & n7320;
  assign n7322 = ~n6960 & ~n7321;
  assign n7323 = n6960 & n7321;
  assign n7324 = ~n7322 & ~n7323;
  assign n7325 = ~n7319 & ~n7324;
  assign n7326 = ~n7318 & ~n7325;
  assign n7327 = po61  & ~n7326;
  assign n7328 = ~po61  & n7326;
  assign n7329 = ~n6963 & ~n6964;
  assign n7330 = po25  & n7329;
  assign n7331 = ~n6969 & ~n7330;
  assign n7332 = n6969 & n7330;
  assign n7333 = ~n7331 & ~n7332;
  assign n7334 = ~n7328 & ~n7333;
  assign n7335 = ~n7327 & ~n7334;
  assign n7336 = po62  & ~n7335;
  assign n7337 = ~po62  & n7335;
  assign n7338 = ~n6972 & ~n6973;
  assign n7339 = po25  & n7338;
  assign n7340 = ~n6978 & ~n7339;
  assign n7341 = n6978 & n7339;
  assign n7342 = ~n7340 & ~n7341;
  assign n7343 = ~n7337 & ~n7342;
  assign n7344 = ~n7336 & ~n7343;
  assign n7345 = n7013 & n7344;
  assign n7346 = ~n7013 & ~n7344;
  assign n7347 = n6991 & po25 ;
  assign n7348 = ~n6990 & ~n7347;
  assign n7349 = n7346 & n7348;
  assign n7350 = ~po63  & ~n7349;
  assign n7351 = ~n7345 & ~n7350;
  assign n7352 = ~n7008 & n7351;
  assign po24  = n7004 | ~n7352;
  assign n7354 = ~n7143 & ~n7144;
  assign n7355 = po24  & n7354;
  assign n7356 = ~n7003 & ~n7355;
  assign n7357 = n7003 & n7355;
  assign n7358 = ~n7356 & ~n7357;
  assign n7359 = n7013 & ~po24 ;
  assign n7360 = ~n7013 & po24 ;
  assign n7361 = n7344 & ~n7360;
  assign n7362 = po63  & ~n7361;
  assign n7363 = ~n7346 & n7362;
  assign n7364 = ~n7336 & ~n7337;
  assign n7365 = po24  & n7364;
  assign n7366 = ~n7342 & ~n7365;
  assign n7367 = n7342 & n7365;
  assign n7368 = ~n7366 & ~n7367;
  assign n7369 = pi48  & po24 ;
  assign n7370 = ~pi46  & ~pi47 ;
  assign n7371 = ~pi48  & n7370;
  assign n7372 = ~n7369 & ~n7371;
  assign n7373 = po25  & ~n7372;
  assign n7374 = ~po25  & n7372;
  assign n7375 = ~pi48  & po24 ;
  assign n7376 = pi49  & ~n7375;
  assign n7377 = n7015 & po24 ;
  assign n7378 = ~n7376 & ~n7377;
  assign n7379 = ~n7374 & n7378;
  assign n7380 = ~n7373 & ~n7379;
  assign n7381 = po26  & ~n7380;
  assign n7382 = ~po26  & n7380;
  assign n7383 = po25  & n7352;
  assign n7384 = ~n7377 & ~n7383;
  assign n7385 = pi50  & ~n7384;
  assign n7386 = ~pi50  & n7384;
  assign n7387 = ~n7385 & ~n7386;
  assign n7388 = ~n7382 & ~n7387;
  assign n7389 = ~n7381 & ~n7388;
  assign n7390 = po27  & ~n7389;
  assign n7391 = ~po27  & n7389;
  assign n7392 = ~n7018 & ~n7019;
  assign n7393 = po24  & n7392;
  assign n7394 = n7023 & ~n7393;
  assign n7395 = ~n7023 & n7393;
  assign n7396 = ~n7394 & ~n7395;
  assign n7397 = ~n7391 & ~n7396;
  assign n7398 = ~n7390 & ~n7397;
  assign n7399 = po28  & ~n7398;
  assign n7400 = ~po28  & n7398;
  assign n7401 = ~n7026 & ~n7027;
  assign n7402 = po24  & n7401;
  assign n7403 = ~n7032 & ~n7402;
  assign n7404 = n7032 & n7402;
  assign n7405 = ~n7403 & ~n7404;
  assign n7406 = ~n7400 & ~n7405;
  assign n7407 = ~n7399 & ~n7406;
  assign n7408 = po29  & ~n7407;
  assign n7409 = ~po29  & n7407;
  assign n7410 = ~n7035 & ~n7036;
  assign n7411 = po24  & n7410;
  assign n7412 = n7041 & n7411;
  assign n7413 = ~n7041 & ~n7411;
  assign n7414 = ~n7412 & ~n7413;
  assign n7415 = ~n7409 & ~n7414;
  assign n7416 = ~n7408 & ~n7415;
  assign n7417 = po30  & ~n7416;
  assign n7418 = ~po30  & n7416;
  assign n7419 = ~n7044 & ~n7045;
  assign n7420 = po24  & n7419;
  assign n7421 = ~n7050 & ~n7420;
  assign n7422 = n7050 & n7420;
  assign n7423 = ~n7421 & ~n7422;
  assign n7424 = ~n7418 & ~n7423;
  assign n7425 = ~n7417 & ~n7424;
  assign n7426 = po31  & ~n7425;
  assign n7427 = ~po31  & n7425;
  assign n7428 = ~n7053 & ~n7054;
  assign n7429 = po24  & n7428;
  assign n7430 = ~n7059 & ~n7429;
  assign n7431 = n7059 & n7429;
  assign n7432 = ~n7430 & ~n7431;
  assign n7433 = ~n7427 & ~n7432;
  assign n7434 = ~n7426 & ~n7433;
  assign n7435 = po32  & ~n7434;
  assign n7436 = ~po32  & n7434;
  assign n7437 = ~n7062 & ~n7063;
  assign n7438 = po24  & n7437;
  assign n7439 = ~n7068 & ~n7438;
  assign n7440 = n7068 & n7438;
  assign n7441 = ~n7439 & ~n7440;
  assign n7442 = ~n7436 & ~n7441;
  assign n7443 = ~n7435 & ~n7442;
  assign n7444 = po33  & ~n7443;
  assign n7445 = ~po33  & n7443;
  assign n7446 = ~n7071 & ~n7072;
  assign n7447 = po24  & n7446;
  assign n7448 = ~n7077 & ~n7447;
  assign n7449 = n7077 & n7447;
  assign n7450 = ~n7448 & ~n7449;
  assign n7451 = ~n7445 & ~n7450;
  assign n7452 = ~n7444 & ~n7451;
  assign n7453 = po34  & ~n7452;
  assign n7454 = ~po34  & n7452;
  assign n7455 = ~n7080 & ~n7081;
  assign n7456 = po24  & n7455;
  assign n7457 = ~n7086 & ~n7456;
  assign n7458 = n7086 & n7456;
  assign n7459 = ~n7457 & ~n7458;
  assign n7460 = ~n7454 & ~n7459;
  assign n7461 = ~n7453 & ~n7460;
  assign n7462 = po35  & ~n7461;
  assign n7463 = ~po35  & n7461;
  assign n7464 = ~n7089 & ~n7090;
  assign n7465 = po24  & n7464;
  assign n7466 = ~n7095 & ~n7465;
  assign n7467 = n7095 & n7465;
  assign n7468 = ~n7466 & ~n7467;
  assign n7469 = ~n7463 & ~n7468;
  assign n7470 = ~n7462 & ~n7469;
  assign n7471 = po36  & ~n7470;
  assign n7472 = ~po36  & n7470;
  assign n7473 = ~n7098 & ~n7099;
  assign n7474 = po24  & n7473;
  assign n7475 = ~n7104 & ~n7474;
  assign n7476 = n7104 & n7474;
  assign n7477 = ~n7475 & ~n7476;
  assign n7478 = ~n7472 & ~n7477;
  assign n7479 = ~n7471 & ~n7478;
  assign n7480 = po37  & ~n7479;
  assign n7481 = ~po37  & n7479;
  assign n7482 = ~n7107 & ~n7108;
  assign n7483 = po24  & n7482;
  assign n7484 = ~n7113 & ~n7483;
  assign n7485 = n7113 & n7483;
  assign n7486 = ~n7484 & ~n7485;
  assign n7487 = ~n7481 & ~n7486;
  assign n7488 = ~n7480 & ~n7487;
  assign n7489 = po38  & ~n7488;
  assign n7490 = ~po38  & n7488;
  assign n7491 = ~n7116 & ~n7117;
  assign n7492 = po24  & n7491;
  assign n7493 = ~n7122 & ~n7492;
  assign n7494 = n7122 & n7492;
  assign n7495 = ~n7493 & ~n7494;
  assign n7496 = ~n7490 & ~n7495;
  assign n7497 = ~n7489 & ~n7496;
  assign n7498 = po39  & ~n7497;
  assign n7499 = ~po39  & n7497;
  assign n7500 = ~n7125 & ~n7126;
  assign n7501 = po24  & n7500;
  assign n7502 = ~n7131 & ~n7501;
  assign n7503 = n7131 & n7501;
  assign n7504 = ~n7502 & ~n7503;
  assign n7505 = ~n7499 & ~n7504;
  assign n7506 = ~n7498 & ~n7505;
  assign n7507 = po40  & ~n7506;
  assign n7508 = ~n7134 & ~n7140;
  assign n7509 = po24  & n7508;
  assign n7510 = ~n7139 & ~n7509;
  assign n7511 = n7139 & n7509;
  assign n7512 = ~n7510 & ~n7511;
  assign n7513 = ~po40  & n7506;
  assign n7514 = ~n7512 & ~n7513;
  assign n7515 = ~n7507 & ~n7514;
  assign n7516 = po41  & ~n7515;
  assign n7517 = ~po41  & n7515;
  assign n7518 = ~n7358 & ~n7517;
  assign n7519 = ~n7516 & ~n7518;
  assign n7520 = po42  & ~n7519;
  assign n7521 = ~po42  & n7519;
  assign n7522 = ~n7147 & ~n7148;
  assign n7523 = po24  & n7522;
  assign n7524 = ~n7153 & ~n7523;
  assign n7525 = n7153 & n7523;
  assign n7526 = ~n7524 & ~n7525;
  assign n7527 = ~n7521 & ~n7526;
  assign n7528 = ~n7520 & ~n7527;
  assign n7529 = po43  & ~n7528;
  assign n7530 = ~po43  & n7528;
  assign n7531 = ~n7156 & ~n7157;
  assign n7532 = po24  & n7531;
  assign n7533 = ~n7162 & ~n7532;
  assign n7534 = n7162 & n7532;
  assign n7535 = ~n7533 & ~n7534;
  assign n7536 = ~n7530 & ~n7535;
  assign n7537 = ~n7529 & ~n7536;
  assign n7538 = po44  & ~n7537;
  assign n7539 = ~po44  & n7537;
  assign n7540 = ~n7165 & ~n7166;
  assign n7541 = po24  & n7540;
  assign n7542 = ~n7171 & ~n7541;
  assign n7543 = n7171 & n7541;
  assign n7544 = ~n7542 & ~n7543;
  assign n7545 = ~n7539 & ~n7544;
  assign n7546 = ~n7538 & ~n7545;
  assign n7547 = po45  & ~n7546;
  assign n7548 = ~po45  & n7546;
  assign n7549 = ~n7174 & ~n7175;
  assign n7550 = po24  & n7549;
  assign n7551 = ~n7180 & ~n7550;
  assign n7552 = n7180 & n7550;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = ~n7548 & ~n7553;
  assign n7555 = ~n7547 & ~n7554;
  assign n7556 = po46  & ~n7555;
  assign n7557 = ~po46  & n7555;
  assign n7558 = ~n7183 & ~n7184;
  assign n7559 = po24  & n7558;
  assign n7560 = ~n7189 & ~n7559;
  assign n7561 = n7189 & n7559;
  assign n7562 = ~n7560 & ~n7561;
  assign n7563 = ~n7557 & ~n7562;
  assign n7564 = ~n7556 & ~n7563;
  assign n7565 = po47  & ~n7564;
  assign n7566 = ~po47  & n7564;
  assign n7567 = ~n7192 & ~n7193;
  assign n7568 = po24  & n7567;
  assign n7569 = ~n7198 & ~n7568;
  assign n7570 = n7198 & n7568;
  assign n7571 = ~n7569 & ~n7570;
  assign n7572 = ~n7566 & ~n7571;
  assign n7573 = ~n7565 & ~n7572;
  assign n7574 = po48  & ~n7573;
  assign n7575 = ~po48  & n7573;
  assign n7576 = ~n7201 & ~n7202;
  assign n7577 = po24  & n7576;
  assign n7578 = ~n7207 & ~n7577;
  assign n7579 = n7207 & n7577;
  assign n7580 = ~n7578 & ~n7579;
  assign n7581 = ~n7575 & ~n7580;
  assign n7582 = ~n7574 & ~n7581;
  assign n7583 = po49  & ~n7582;
  assign n7584 = ~po49  & n7582;
  assign n7585 = ~n7210 & ~n7211;
  assign n7586 = po24  & n7585;
  assign n7587 = ~n7216 & ~n7586;
  assign n7588 = n7216 & n7586;
  assign n7589 = ~n7587 & ~n7588;
  assign n7590 = ~n7584 & ~n7589;
  assign n7591 = ~n7583 & ~n7590;
  assign n7592 = po50  & ~n7591;
  assign n7593 = ~po50  & n7591;
  assign n7594 = ~n7219 & ~n7220;
  assign n7595 = po24  & n7594;
  assign n7596 = ~n7225 & ~n7595;
  assign n7597 = n7225 & n7595;
  assign n7598 = ~n7596 & ~n7597;
  assign n7599 = ~n7593 & ~n7598;
  assign n7600 = ~n7592 & ~n7599;
  assign n7601 = po51  & ~n7600;
  assign n7602 = ~po51  & n7600;
  assign n7603 = ~n7228 & ~n7229;
  assign n7604 = po24  & n7603;
  assign n7605 = ~n7234 & ~n7604;
  assign n7606 = n7234 & n7604;
  assign n7607 = ~n7605 & ~n7606;
  assign n7608 = ~n7602 & ~n7607;
  assign n7609 = ~n7601 & ~n7608;
  assign n7610 = po52  & ~n7609;
  assign n7611 = ~po52  & n7609;
  assign n7612 = ~n7237 & ~n7238;
  assign n7613 = po24  & n7612;
  assign n7614 = ~n7243 & ~n7613;
  assign n7615 = n7243 & n7613;
  assign n7616 = ~n7614 & ~n7615;
  assign n7617 = ~n7611 & ~n7616;
  assign n7618 = ~n7610 & ~n7617;
  assign n7619 = po53  & ~n7618;
  assign n7620 = ~po53  & n7618;
  assign n7621 = ~n7246 & ~n7247;
  assign n7622 = po24  & n7621;
  assign n7623 = ~n7252 & ~n7622;
  assign n7624 = n7252 & n7622;
  assign n7625 = ~n7623 & ~n7624;
  assign n7626 = ~n7620 & ~n7625;
  assign n7627 = ~n7619 & ~n7626;
  assign n7628 = po54  & ~n7627;
  assign n7629 = ~po54  & n7627;
  assign n7630 = ~n7255 & ~n7256;
  assign n7631 = po24  & n7630;
  assign n7632 = ~n7261 & ~n7631;
  assign n7633 = n7261 & n7631;
  assign n7634 = ~n7632 & ~n7633;
  assign n7635 = ~n7629 & ~n7634;
  assign n7636 = ~n7628 & ~n7635;
  assign n7637 = po55  & ~n7636;
  assign n7638 = ~po55  & n7636;
  assign n7639 = ~n7264 & ~n7265;
  assign n7640 = po24  & n7639;
  assign n7641 = ~n7270 & ~n7640;
  assign n7642 = n7270 & n7640;
  assign n7643 = ~n7641 & ~n7642;
  assign n7644 = ~n7638 & ~n7643;
  assign n7645 = ~n7637 & ~n7644;
  assign n7646 = po56  & ~n7645;
  assign n7647 = ~po56  & n7645;
  assign n7648 = ~n7273 & ~n7274;
  assign n7649 = po24  & n7648;
  assign n7650 = ~n7279 & ~n7649;
  assign n7651 = n7279 & n7649;
  assign n7652 = ~n7650 & ~n7651;
  assign n7653 = ~n7647 & ~n7652;
  assign n7654 = ~n7646 & ~n7653;
  assign n7655 = po57  & ~n7654;
  assign n7656 = ~po57  & n7654;
  assign n7657 = ~n7282 & ~n7283;
  assign n7658 = po24  & n7657;
  assign n7659 = ~n7288 & ~n7658;
  assign n7660 = n7288 & n7658;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = ~n7656 & ~n7661;
  assign n7663 = ~n7655 & ~n7662;
  assign n7664 = po58  & ~n7663;
  assign n7665 = ~po58  & n7663;
  assign n7666 = ~n7291 & ~n7292;
  assign n7667 = po24  & n7666;
  assign n7668 = ~n7297 & ~n7667;
  assign n7669 = n7297 & n7667;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~n7665 & ~n7670;
  assign n7672 = ~n7664 & ~n7671;
  assign n7673 = po59  & ~n7672;
  assign n7674 = ~po59  & n7672;
  assign n7675 = ~n7300 & ~n7301;
  assign n7676 = po24  & n7675;
  assign n7677 = ~n7306 & ~n7676;
  assign n7678 = n7306 & n7676;
  assign n7679 = ~n7677 & ~n7678;
  assign n7680 = ~n7674 & ~n7679;
  assign n7681 = ~n7673 & ~n7680;
  assign n7682 = po60  & ~n7681;
  assign n7683 = ~po60  & n7681;
  assign n7684 = ~n7309 & ~n7310;
  assign n7685 = po24  & n7684;
  assign n7686 = ~n7315 & ~n7685;
  assign n7687 = n7315 & n7685;
  assign n7688 = ~n7686 & ~n7687;
  assign n7689 = ~n7683 & ~n7688;
  assign n7690 = ~n7682 & ~n7689;
  assign n7691 = po61  & ~n7690;
  assign n7692 = ~po61  & n7690;
  assign n7693 = ~n7318 & ~n7319;
  assign n7694 = po24  & n7693;
  assign n7695 = ~n7324 & ~n7694;
  assign n7696 = n7324 & n7694;
  assign n7697 = ~n7695 & ~n7696;
  assign n7698 = ~n7692 & ~n7697;
  assign n7699 = ~n7691 & ~n7698;
  assign n7700 = po62  & ~n7699;
  assign n7701 = ~po62  & n7699;
  assign n7702 = ~n7327 & ~n7328;
  assign n7703 = po24  & n7702;
  assign n7704 = ~n7333 & ~n7703;
  assign n7705 = n7333 & n7703;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = ~n7701 & ~n7706;
  assign n7708 = ~n7700 & ~n7707;
  assign n7709 = n7368 & n7708;
  assign n7710 = ~n7368 & ~n7708;
  assign n7711 = n7346 & po24 ;
  assign n7712 = ~n7345 & ~n7711;
  assign n7713 = n7710 & n7712;
  assign n7714 = ~po63  & ~n7713;
  assign n7715 = ~n7709 & ~n7714;
  assign n7716 = ~n7363 & n7715;
  assign po23  = n7359 | ~n7716;
  assign n7718 = ~n7516 & ~n7517;
  assign n7719 = po23  & n7718;
  assign n7720 = ~n7358 & ~n7719;
  assign n7721 = n7358 & n7719;
  assign n7722 = ~n7720 & ~n7721;
  assign n7723 = n7368 & ~po23 ;
  assign n7724 = ~n7368 & po23 ;
  assign n7725 = n7708 & ~n7724;
  assign n7726 = po63  & ~n7725;
  assign n7727 = ~n7710 & n7726;
  assign n7728 = ~n7700 & ~n7701;
  assign n7729 = po23  & n7728;
  assign n7730 = ~n7706 & ~n7729;
  assign n7731 = n7706 & n7729;
  assign n7732 = ~n7730 & ~n7731;
  assign n7733 = pi46  & po23 ;
  assign n7734 = ~pi44  & ~pi45 ;
  assign n7735 = ~pi46  & n7734;
  assign n7736 = ~n7733 & ~n7735;
  assign n7737 = po24  & ~n7736;
  assign n7738 = ~po24  & n7736;
  assign n7739 = ~pi46  & po23 ;
  assign n7740 = pi47  & ~n7739;
  assign n7741 = n7370 & po23 ;
  assign n7742 = ~n7740 & ~n7741;
  assign n7743 = ~n7738 & n7742;
  assign n7744 = ~n7737 & ~n7743;
  assign n7745 = po25  & ~n7744;
  assign n7746 = ~po25  & n7744;
  assign n7747 = po24  & n7716;
  assign n7748 = ~n7741 & ~n7747;
  assign n7749 = pi48  & ~n7748;
  assign n7750 = ~pi48  & n7748;
  assign n7751 = ~n7749 & ~n7750;
  assign n7752 = ~n7746 & ~n7751;
  assign n7753 = ~n7745 & ~n7752;
  assign n7754 = po26  & ~n7753;
  assign n7755 = ~po26  & n7753;
  assign n7756 = ~n7373 & ~n7374;
  assign n7757 = po23  & n7756;
  assign n7758 = n7378 & ~n7757;
  assign n7759 = ~n7378 & n7757;
  assign n7760 = ~n7758 & ~n7759;
  assign n7761 = ~n7755 & ~n7760;
  assign n7762 = ~n7754 & ~n7761;
  assign n7763 = po27  & ~n7762;
  assign n7764 = ~po27  & n7762;
  assign n7765 = ~n7381 & ~n7382;
  assign n7766 = po23  & n7765;
  assign n7767 = ~n7387 & ~n7766;
  assign n7768 = n7387 & n7766;
  assign n7769 = ~n7767 & ~n7768;
  assign n7770 = ~n7764 & ~n7769;
  assign n7771 = ~n7763 & ~n7770;
  assign n7772 = po28  & ~n7771;
  assign n7773 = ~po28  & n7771;
  assign n7774 = ~n7390 & ~n7391;
  assign n7775 = po23  & n7774;
  assign n7776 = n7396 & n7775;
  assign n7777 = ~n7396 & ~n7775;
  assign n7778 = ~n7776 & ~n7777;
  assign n7779 = ~n7773 & ~n7778;
  assign n7780 = ~n7772 & ~n7779;
  assign n7781 = po29  & ~n7780;
  assign n7782 = ~po29  & n7780;
  assign n7783 = ~n7399 & ~n7400;
  assign n7784 = po23  & n7783;
  assign n7785 = ~n7405 & ~n7784;
  assign n7786 = n7405 & n7784;
  assign n7787 = ~n7785 & ~n7786;
  assign n7788 = ~n7782 & ~n7787;
  assign n7789 = ~n7781 & ~n7788;
  assign n7790 = po30  & ~n7789;
  assign n7791 = ~po30  & n7789;
  assign n7792 = ~n7408 & ~n7409;
  assign n7793 = po23  & n7792;
  assign n7794 = ~n7414 & ~n7793;
  assign n7795 = n7414 & n7793;
  assign n7796 = ~n7794 & ~n7795;
  assign n7797 = ~n7791 & ~n7796;
  assign n7798 = ~n7790 & ~n7797;
  assign n7799 = po31  & ~n7798;
  assign n7800 = ~po31  & n7798;
  assign n7801 = ~n7417 & ~n7418;
  assign n7802 = po23  & n7801;
  assign n7803 = ~n7423 & ~n7802;
  assign n7804 = n7423 & n7802;
  assign n7805 = ~n7803 & ~n7804;
  assign n7806 = ~n7800 & ~n7805;
  assign n7807 = ~n7799 & ~n7806;
  assign n7808 = po32  & ~n7807;
  assign n7809 = ~po32  & n7807;
  assign n7810 = ~n7426 & ~n7427;
  assign n7811 = po23  & n7810;
  assign n7812 = ~n7432 & ~n7811;
  assign n7813 = n7432 & n7811;
  assign n7814 = ~n7812 & ~n7813;
  assign n7815 = ~n7809 & ~n7814;
  assign n7816 = ~n7808 & ~n7815;
  assign n7817 = po33  & ~n7816;
  assign n7818 = ~po33  & n7816;
  assign n7819 = ~n7435 & ~n7436;
  assign n7820 = po23  & n7819;
  assign n7821 = ~n7441 & ~n7820;
  assign n7822 = n7441 & n7820;
  assign n7823 = ~n7821 & ~n7822;
  assign n7824 = ~n7818 & ~n7823;
  assign n7825 = ~n7817 & ~n7824;
  assign n7826 = po34  & ~n7825;
  assign n7827 = ~po34  & n7825;
  assign n7828 = ~n7444 & ~n7445;
  assign n7829 = po23  & n7828;
  assign n7830 = ~n7450 & ~n7829;
  assign n7831 = n7450 & n7829;
  assign n7832 = ~n7830 & ~n7831;
  assign n7833 = ~n7827 & ~n7832;
  assign n7834 = ~n7826 & ~n7833;
  assign n7835 = po35  & ~n7834;
  assign n7836 = ~po35  & n7834;
  assign n7837 = ~n7453 & ~n7454;
  assign n7838 = po23  & n7837;
  assign n7839 = ~n7459 & ~n7838;
  assign n7840 = n7459 & n7838;
  assign n7841 = ~n7839 & ~n7840;
  assign n7842 = ~n7836 & ~n7841;
  assign n7843 = ~n7835 & ~n7842;
  assign n7844 = po36  & ~n7843;
  assign n7845 = ~po36  & n7843;
  assign n7846 = ~n7462 & ~n7463;
  assign n7847 = po23  & n7846;
  assign n7848 = ~n7468 & ~n7847;
  assign n7849 = n7468 & n7847;
  assign n7850 = ~n7848 & ~n7849;
  assign n7851 = ~n7845 & ~n7850;
  assign n7852 = ~n7844 & ~n7851;
  assign n7853 = po37  & ~n7852;
  assign n7854 = ~po37  & n7852;
  assign n7855 = ~n7471 & ~n7472;
  assign n7856 = po23  & n7855;
  assign n7857 = ~n7477 & ~n7856;
  assign n7858 = n7477 & n7856;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = ~n7854 & ~n7859;
  assign n7861 = ~n7853 & ~n7860;
  assign n7862 = po38  & ~n7861;
  assign n7863 = ~po38  & n7861;
  assign n7864 = ~n7480 & ~n7481;
  assign n7865 = po23  & n7864;
  assign n7866 = ~n7486 & ~n7865;
  assign n7867 = n7486 & n7865;
  assign n7868 = ~n7866 & ~n7867;
  assign n7869 = ~n7863 & ~n7868;
  assign n7870 = ~n7862 & ~n7869;
  assign n7871 = po39  & ~n7870;
  assign n7872 = ~po39  & n7870;
  assign n7873 = ~n7489 & ~n7490;
  assign n7874 = po23  & n7873;
  assign n7875 = ~n7495 & ~n7874;
  assign n7876 = n7495 & n7874;
  assign n7877 = ~n7875 & ~n7876;
  assign n7878 = ~n7872 & ~n7877;
  assign n7879 = ~n7871 & ~n7878;
  assign n7880 = po40  & ~n7879;
  assign n7881 = ~po40  & n7879;
  assign n7882 = ~n7498 & ~n7499;
  assign n7883 = po23  & n7882;
  assign n7884 = ~n7504 & ~n7883;
  assign n7885 = n7504 & n7883;
  assign n7886 = ~n7884 & ~n7885;
  assign n7887 = ~n7881 & ~n7886;
  assign n7888 = ~n7880 & ~n7887;
  assign n7889 = po41  & ~n7888;
  assign n7890 = ~n7507 & ~n7513;
  assign n7891 = po23  & n7890;
  assign n7892 = ~n7512 & ~n7891;
  assign n7893 = n7512 & n7891;
  assign n7894 = ~n7892 & ~n7893;
  assign n7895 = ~po41  & n7888;
  assign n7896 = ~n7894 & ~n7895;
  assign n7897 = ~n7889 & ~n7896;
  assign n7898 = po42  & ~n7897;
  assign n7899 = ~po42  & n7897;
  assign n7900 = ~n7722 & ~n7899;
  assign n7901 = ~n7898 & ~n7900;
  assign n7902 = po43  & ~n7901;
  assign n7903 = ~po43  & n7901;
  assign n7904 = ~n7520 & ~n7521;
  assign n7905 = po23  & n7904;
  assign n7906 = ~n7526 & ~n7905;
  assign n7907 = n7526 & n7905;
  assign n7908 = ~n7906 & ~n7907;
  assign n7909 = ~n7903 & ~n7908;
  assign n7910 = ~n7902 & ~n7909;
  assign n7911 = po44  & ~n7910;
  assign n7912 = ~po44  & n7910;
  assign n7913 = ~n7529 & ~n7530;
  assign n7914 = po23  & n7913;
  assign n7915 = ~n7535 & ~n7914;
  assign n7916 = n7535 & n7914;
  assign n7917 = ~n7915 & ~n7916;
  assign n7918 = ~n7912 & ~n7917;
  assign n7919 = ~n7911 & ~n7918;
  assign n7920 = po45  & ~n7919;
  assign n7921 = ~po45  & n7919;
  assign n7922 = ~n7538 & ~n7539;
  assign n7923 = po23  & n7922;
  assign n7924 = ~n7544 & ~n7923;
  assign n7925 = n7544 & n7923;
  assign n7926 = ~n7924 & ~n7925;
  assign n7927 = ~n7921 & ~n7926;
  assign n7928 = ~n7920 & ~n7927;
  assign n7929 = po46  & ~n7928;
  assign n7930 = ~po46  & n7928;
  assign n7931 = ~n7547 & ~n7548;
  assign n7932 = po23  & n7931;
  assign n7933 = ~n7553 & ~n7932;
  assign n7934 = n7553 & n7932;
  assign n7935 = ~n7933 & ~n7934;
  assign n7936 = ~n7930 & ~n7935;
  assign n7937 = ~n7929 & ~n7936;
  assign n7938 = po47  & ~n7937;
  assign n7939 = ~po47  & n7937;
  assign n7940 = ~n7556 & ~n7557;
  assign n7941 = po23  & n7940;
  assign n7942 = ~n7562 & ~n7941;
  assign n7943 = n7562 & n7941;
  assign n7944 = ~n7942 & ~n7943;
  assign n7945 = ~n7939 & ~n7944;
  assign n7946 = ~n7938 & ~n7945;
  assign n7947 = po48  & ~n7946;
  assign n7948 = ~po48  & n7946;
  assign n7949 = ~n7565 & ~n7566;
  assign n7950 = po23  & n7949;
  assign n7951 = ~n7571 & ~n7950;
  assign n7952 = n7571 & n7950;
  assign n7953 = ~n7951 & ~n7952;
  assign n7954 = ~n7948 & ~n7953;
  assign n7955 = ~n7947 & ~n7954;
  assign n7956 = po49  & ~n7955;
  assign n7957 = ~po49  & n7955;
  assign n7958 = ~n7574 & ~n7575;
  assign n7959 = po23  & n7958;
  assign n7960 = ~n7580 & ~n7959;
  assign n7961 = n7580 & n7959;
  assign n7962 = ~n7960 & ~n7961;
  assign n7963 = ~n7957 & ~n7962;
  assign n7964 = ~n7956 & ~n7963;
  assign n7965 = po50  & ~n7964;
  assign n7966 = ~po50  & n7964;
  assign n7967 = ~n7583 & ~n7584;
  assign n7968 = po23  & n7967;
  assign n7969 = ~n7589 & ~n7968;
  assign n7970 = n7589 & n7968;
  assign n7971 = ~n7969 & ~n7970;
  assign n7972 = ~n7966 & ~n7971;
  assign n7973 = ~n7965 & ~n7972;
  assign n7974 = po51  & ~n7973;
  assign n7975 = ~po51  & n7973;
  assign n7976 = ~n7592 & ~n7593;
  assign n7977 = po23  & n7976;
  assign n7978 = ~n7598 & ~n7977;
  assign n7979 = n7598 & n7977;
  assign n7980 = ~n7978 & ~n7979;
  assign n7981 = ~n7975 & ~n7980;
  assign n7982 = ~n7974 & ~n7981;
  assign n7983 = po52  & ~n7982;
  assign n7984 = ~po52  & n7982;
  assign n7985 = ~n7601 & ~n7602;
  assign n7986 = po23  & n7985;
  assign n7987 = ~n7607 & ~n7986;
  assign n7988 = n7607 & n7986;
  assign n7989 = ~n7987 & ~n7988;
  assign n7990 = ~n7984 & ~n7989;
  assign n7991 = ~n7983 & ~n7990;
  assign n7992 = po53  & ~n7991;
  assign n7993 = ~po53  & n7991;
  assign n7994 = ~n7610 & ~n7611;
  assign n7995 = po23  & n7994;
  assign n7996 = ~n7616 & ~n7995;
  assign n7997 = n7616 & n7995;
  assign n7998 = ~n7996 & ~n7997;
  assign n7999 = ~n7993 & ~n7998;
  assign n8000 = ~n7992 & ~n7999;
  assign n8001 = po54  & ~n8000;
  assign n8002 = ~po54  & n8000;
  assign n8003 = ~n7619 & ~n7620;
  assign n8004 = po23  & n8003;
  assign n8005 = ~n7625 & ~n8004;
  assign n8006 = n7625 & n8004;
  assign n8007 = ~n8005 & ~n8006;
  assign n8008 = ~n8002 & ~n8007;
  assign n8009 = ~n8001 & ~n8008;
  assign n8010 = po55  & ~n8009;
  assign n8011 = ~po55  & n8009;
  assign n8012 = ~n7628 & ~n7629;
  assign n8013 = po23  & n8012;
  assign n8014 = ~n7634 & ~n8013;
  assign n8015 = n7634 & n8013;
  assign n8016 = ~n8014 & ~n8015;
  assign n8017 = ~n8011 & ~n8016;
  assign n8018 = ~n8010 & ~n8017;
  assign n8019 = po56  & ~n8018;
  assign n8020 = ~po56  & n8018;
  assign n8021 = ~n7637 & ~n7638;
  assign n8022 = po23  & n8021;
  assign n8023 = ~n7643 & ~n8022;
  assign n8024 = n7643 & n8022;
  assign n8025 = ~n8023 & ~n8024;
  assign n8026 = ~n8020 & ~n8025;
  assign n8027 = ~n8019 & ~n8026;
  assign n8028 = po57  & ~n8027;
  assign n8029 = ~po57  & n8027;
  assign n8030 = ~n7646 & ~n7647;
  assign n8031 = po23  & n8030;
  assign n8032 = ~n7652 & ~n8031;
  assign n8033 = n7652 & n8031;
  assign n8034 = ~n8032 & ~n8033;
  assign n8035 = ~n8029 & ~n8034;
  assign n8036 = ~n8028 & ~n8035;
  assign n8037 = po58  & ~n8036;
  assign n8038 = ~po58  & n8036;
  assign n8039 = ~n7655 & ~n7656;
  assign n8040 = po23  & n8039;
  assign n8041 = ~n7661 & ~n8040;
  assign n8042 = n7661 & n8040;
  assign n8043 = ~n8041 & ~n8042;
  assign n8044 = ~n8038 & ~n8043;
  assign n8045 = ~n8037 & ~n8044;
  assign n8046 = po59  & ~n8045;
  assign n8047 = ~po59  & n8045;
  assign n8048 = ~n7664 & ~n7665;
  assign n8049 = po23  & n8048;
  assign n8050 = ~n7670 & ~n8049;
  assign n8051 = n7670 & n8049;
  assign n8052 = ~n8050 & ~n8051;
  assign n8053 = ~n8047 & ~n8052;
  assign n8054 = ~n8046 & ~n8053;
  assign n8055 = po60  & ~n8054;
  assign n8056 = ~po60  & n8054;
  assign n8057 = ~n7673 & ~n7674;
  assign n8058 = po23  & n8057;
  assign n8059 = ~n7679 & ~n8058;
  assign n8060 = n7679 & n8058;
  assign n8061 = ~n8059 & ~n8060;
  assign n8062 = ~n8056 & ~n8061;
  assign n8063 = ~n8055 & ~n8062;
  assign n8064 = po61  & ~n8063;
  assign n8065 = ~po61  & n8063;
  assign n8066 = ~n7682 & ~n7683;
  assign n8067 = po23  & n8066;
  assign n8068 = ~n7688 & ~n8067;
  assign n8069 = n7688 & n8067;
  assign n8070 = ~n8068 & ~n8069;
  assign n8071 = ~n8065 & ~n8070;
  assign n8072 = ~n8064 & ~n8071;
  assign n8073 = po62  & ~n8072;
  assign n8074 = ~po62  & n8072;
  assign n8075 = ~n7691 & ~n7692;
  assign n8076 = po23  & n8075;
  assign n8077 = ~n7697 & ~n8076;
  assign n8078 = n7697 & n8076;
  assign n8079 = ~n8077 & ~n8078;
  assign n8080 = ~n8074 & ~n8079;
  assign n8081 = ~n8073 & ~n8080;
  assign n8082 = n7732 & n8081;
  assign n8083 = ~n7732 & ~n8081;
  assign n8084 = n7710 & po23 ;
  assign n8085 = ~n7709 & ~n8084;
  assign n8086 = n8083 & n8085;
  assign n8087 = ~po63  & ~n8086;
  assign n8088 = ~n8082 & ~n8087;
  assign n8089 = ~n7727 & n8088;
  assign po22  = n7723 | ~n8089;
  assign n8091 = ~n7898 & ~n7899;
  assign n8092 = po22  & n8091;
  assign n8093 = ~n7722 & ~n8092;
  assign n8094 = n7722 & n8092;
  assign n8095 = ~n8093 & ~n8094;
  assign n8096 = n7732 & ~po22 ;
  assign n8097 = ~n7732 & po22 ;
  assign n8098 = n8081 & ~n8097;
  assign n8099 = po63  & ~n8098;
  assign n8100 = ~n8083 & n8099;
  assign n8101 = ~n8073 & ~n8074;
  assign n8102 = po22  & n8101;
  assign n8103 = ~n8079 & ~n8102;
  assign n8104 = n8079 & n8102;
  assign n8105 = ~n8103 & ~n8104;
  assign n8106 = pi44  & po22 ;
  assign n8107 = ~pi42  & ~pi43 ;
  assign n8108 = ~pi44  & n8107;
  assign n8109 = ~n8106 & ~n8108;
  assign n8110 = po23  & ~n8109;
  assign n8111 = ~po23  & n8109;
  assign n8112 = ~pi44  & po22 ;
  assign n8113 = pi45  & ~n8112;
  assign n8114 = n7734 & po22 ;
  assign n8115 = ~n8113 & ~n8114;
  assign n8116 = ~n8111 & n8115;
  assign n8117 = ~n8110 & ~n8116;
  assign n8118 = po24  & ~n8117;
  assign n8119 = ~po24  & n8117;
  assign n8120 = po23  & n8089;
  assign n8121 = ~n8114 & ~n8120;
  assign n8122 = pi46  & ~n8121;
  assign n8123 = ~pi46  & n8121;
  assign n8124 = ~n8122 & ~n8123;
  assign n8125 = ~n8119 & ~n8124;
  assign n8126 = ~n8118 & ~n8125;
  assign n8127 = po25  & ~n8126;
  assign n8128 = ~po25  & n8126;
  assign n8129 = ~n7737 & ~n7738;
  assign n8130 = po22  & n8129;
  assign n8131 = n7742 & ~n8130;
  assign n8132 = ~n7742 & n8130;
  assign n8133 = ~n8131 & ~n8132;
  assign n8134 = ~n8128 & ~n8133;
  assign n8135 = ~n8127 & ~n8134;
  assign n8136 = po26  & ~n8135;
  assign n8137 = ~po26  & n8135;
  assign n8138 = ~n7745 & ~n7746;
  assign n8139 = po22  & n8138;
  assign n8140 = ~n7751 & ~n8139;
  assign n8141 = n7751 & n8139;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = ~n8137 & ~n8142;
  assign n8144 = ~n8136 & ~n8143;
  assign n8145 = po27  & ~n8144;
  assign n8146 = ~po27  & n8144;
  assign n8147 = ~n7754 & ~n7755;
  assign n8148 = po22  & n8147;
  assign n8149 = n7760 & n8148;
  assign n8150 = ~n7760 & ~n8148;
  assign n8151 = ~n8149 & ~n8150;
  assign n8152 = ~n8146 & ~n8151;
  assign n8153 = ~n8145 & ~n8152;
  assign n8154 = po28  & ~n8153;
  assign n8155 = ~po28  & n8153;
  assign n8156 = ~n7763 & ~n7764;
  assign n8157 = po22  & n8156;
  assign n8158 = ~n7769 & ~n8157;
  assign n8159 = n7769 & n8157;
  assign n8160 = ~n8158 & ~n8159;
  assign n8161 = ~n8155 & ~n8160;
  assign n8162 = ~n8154 & ~n8161;
  assign n8163 = po29  & ~n8162;
  assign n8164 = ~po29  & n8162;
  assign n8165 = ~n7772 & ~n7773;
  assign n8166 = po22  & n8165;
  assign n8167 = ~n7778 & ~n8166;
  assign n8168 = n7778 & n8166;
  assign n8169 = ~n8167 & ~n8168;
  assign n8170 = ~n8164 & ~n8169;
  assign n8171 = ~n8163 & ~n8170;
  assign n8172 = po30  & ~n8171;
  assign n8173 = ~po30  & n8171;
  assign n8174 = ~n7781 & ~n7782;
  assign n8175 = po22  & n8174;
  assign n8176 = ~n7787 & ~n8175;
  assign n8177 = n7787 & n8175;
  assign n8178 = ~n8176 & ~n8177;
  assign n8179 = ~n8173 & ~n8178;
  assign n8180 = ~n8172 & ~n8179;
  assign n8181 = po31  & ~n8180;
  assign n8182 = ~po31  & n8180;
  assign n8183 = ~n7790 & ~n7791;
  assign n8184 = po22  & n8183;
  assign n8185 = ~n7796 & ~n8184;
  assign n8186 = n7796 & n8184;
  assign n8187 = ~n8185 & ~n8186;
  assign n8188 = ~n8182 & ~n8187;
  assign n8189 = ~n8181 & ~n8188;
  assign n8190 = po32  & ~n8189;
  assign n8191 = ~po32  & n8189;
  assign n8192 = ~n7799 & ~n7800;
  assign n8193 = po22  & n8192;
  assign n8194 = ~n7805 & ~n8193;
  assign n8195 = n7805 & n8193;
  assign n8196 = ~n8194 & ~n8195;
  assign n8197 = ~n8191 & ~n8196;
  assign n8198 = ~n8190 & ~n8197;
  assign n8199 = po33  & ~n8198;
  assign n8200 = ~po33  & n8198;
  assign n8201 = ~n7808 & ~n7809;
  assign n8202 = po22  & n8201;
  assign n8203 = ~n7814 & ~n8202;
  assign n8204 = n7814 & n8202;
  assign n8205 = ~n8203 & ~n8204;
  assign n8206 = ~n8200 & ~n8205;
  assign n8207 = ~n8199 & ~n8206;
  assign n8208 = po34  & ~n8207;
  assign n8209 = ~po34  & n8207;
  assign n8210 = ~n7817 & ~n7818;
  assign n8211 = po22  & n8210;
  assign n8212 = ~n7823 & ~n8211;
  assign n8213 = n7823 & n8211;
  assign n8214 = ~n8212 & ~n8213;
  assign n8215 = ~n8209 & ~n8214;
  assign n8216 = ~n8208 & ~n8215;
  assign n8217 = po35  & ~n8216;
  assign n8218 = ~po35  & n8216;
  assign n8219 = ~n7826 & ~n7827;
  assign n8220 = po22  & n8219;
  assign n8221 = ~n7832 & ~n8220;
  assign n8222 = n7832 & n8220;
  assign n8223 = ~n8221 & ~n8222;
  assign n8224 = ~n8218 & ~n8223;
  assign n8225 = ~n8217 & ~n8224;
  assign n8226 = po36  & ~n8225;
  assign n8227 = ~po36  & n8225;
  assign n8228 = ~n7835 & ~n7836;
  assign n8229 = po22  & n8228;
  assign n8230 = ~n7841 & ~n8229;
  assign n8231 = n7841 & n8229;
  assign n8232 = ~n8230 & ~n8231;
  assign n8233 = ~n8227 & ~n8232;
  assign n8234 = ~n8226 & ~n8233;
  assign n8235 = po37  & ~n8234;
  assign n8236 = ~po37  & n8234;
  assign n8237 = ~n7844 & ~n7845;
  assign n8238 = po22  & n8237;
  assign n8239 = ~n7850 & ~n8238;
  assign n8240 = n7850 & n8238;
  assign n8241 = ~n8239 & ~n8240;
  assign n8242 = ~n8236 & ~n8241;
  assign n8243 = ~n8235 & ~n8242;
  assign n8244 = po38  & ~n8243;
  assign n8245 = ~po38  & n8243;
  assign n8246 = ~n7853 & ~n7854;
  assign n8247 = po22  & n8246;
  assign n8248 = ~n7859 & ~n8247;
  assign n8249 = n7859 & n8247;
  assign n8250 = ~n8248 & ~n8249;
  assign n8251 = ~n8245 & ~n8250;
  assign n8252 = ~n8244 & ~n8251;
  assign n8253 = po39  & ~n8252;
  assign n8254 = ~po39  & n8252;
  assign n8255 = ~n7862 & ~n7863;
  assign n8256 = po22  & n8255;
  assign n8257 = ~n7868 & ~n8256;
  assign n8258 = n7868 & n8256;
  assign n8259 = ~n8257 & ~n8258;
  assign n8260 = ~n8254 & ~n8259;
  assign n8261 = ~n8253 & ~n8260;
  assign n8262 = po40  & ~n8261;
  assign n8263 = ~po40  & n8261;
  assign n8264 = ~n7871 & ~n7872;
  assign n8265 = po22  & n8264;
  assign n8266 = ~n7877 & ~n8265;
  assign n8267 = n7877 & n8265;
  assign n8268 = ~n8266 & ~n8267;
  assign n8269 = ~n8263 & ~n8268;
  assign n8270 = ~n8262 & ~n8269;
  assign n8271 = po41  & ~n8270;
  assign n8272 = ~po41  & n8270;
  assign n8273 = ~n7880 & ~n7881;
  assign n8274 = po22  & n8273;
  assign n8275 = ~n7886 & ~n8274;
  assign n8276 = n7886 & n8274;
  assign n8277 = ~n8275 & ~n8276;
  assign n8278 = ~n8272 & ~n8277;
  assign n8279 = ~n8271 & ~n8278;
  assign n8280 = po42  & ~n8279;
  assign n8281 = ~n7889 & ~n7895;
  assign n8282 = po22  & n8281;
  assign n8283 = ~n7894 & ~n8282;
  assign n8284 = n7894 & n8282;
  assign n8285 = ~n8283 & ~n8284;
  assign n8286 = ~po42  & n8279;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = ~n8280 & ~n8287;
  assign n8289 = po43  & ~n8288;
  assign n8290 = ~po43  & n8288;
  assign n8291 = ~n8095 & ~n8290;
  assign n8292 = ~n8289 & ~n8291;
  assign n8293 = po44  & ~n8292;
  assign n8294 = ~po44  & n8292;
  assign n8295 = ~n7902 & ~n7903;
  assign n8296 = po22  & n8295;
  assign n8297 = ~n7908 & ~n8296;
  assign n8298 = n7908 & n8296;
  assign n8299 = ~n8297 & ~n8298;
  assign n8300 = ~n8294 & ~n8299;
  assign n8301 = ~n8293 & ~n8300;
  assign n8302 = po45  & ~n8301;
  assign n8303 = ~po45  & n8301;
  assign n8304 = ~n7911 & ~n7912;
  assign n8305 = po22  & n8304;
  assign n8306 = ~n7917 & ~n8305;
  assign n8307 = n7917 & n8305;
  assign n8308 = ~n8306 & ~n8307;
  assign n8309 = ~n8303 & ~n8308;
  assign n8310 = ~n8302 & ~n8309;
  assign n8311 = po46  & ~n8310;
  assign n8312 = ~po46  & n8310;
  assign n8313 = ~n7920 & ~n7921;
  assign n8314 = po22  & n8313;
  assign n8315 = ~n7926 & ~n8314;
  assign n8316 = n7926 & n8314;
  assign n8317 = ~n8315 & ~n8316;
  assign n8318 = ~n8312 & ~n8317;
  assign n8319 = ~n8311 & ~n8318;
  assign n8320 = po47  & ~n8319;
  assign n8321 = ~po47  & n8319;
  assign n8322 = ~n7929 & ~n7930;
  assign n8323 = po22  & n8322;
  assign n8324 = ~n7935 & ~n8323;
  assign n8325 = n7935 & n8323;
  assign n8326 = ~n8324 & ~n8325;
  assign n8327 = ~n8321 & ~n8326;
  assign n8328 = ~n8320 & ~n8327;
  assign n8329 = po48  & ~n8328;
  assign n8330 = ~po48  & n8328;
  assign n8331 = ~n7938 & ~n7939;
  assign n8332 = po22  & n8331;
  assign n8333 = ~n7944 & ~n8332;
  assign n8334 = n7944 & n8332;
  assign n8335 = ~n8333 & ~n8334;
  assign n8336 = ~n8330 & ~n8335;
  assign n8337 = ~n8329 & ~n8336;
  assign n8338 = po49  & ~n8337;
  assign n8339 = ~po49  & n8337;
  assign n8340 = ~n7947 & ~n7948;
  assign n8341 = po22  & n8340;
  assign n8342 = ~n7953 & ~n8341;
  assign n8343 = n7953 & n8341;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = ~n8339 & ~n8344;
  assign n8346 = ~n8338 & ~n8345;
  assign n8347 = po50  & ~n8346;
  assign n8348 = ~po50  & n8346;
  assign n8349 = ~n7956 & ~n7957;
  assign n8350 = po22  & n8349;
  assign n8351 = ~n7962 & ~n8350;
  assign n8352 = n7962 & n8350;
  assign n8353 = ~n8351 & ~n8352;
  assign n8354 = ~n8348 & ~n8353;
  assign n8355 = ~n8347 & ~n8354;
  assign n8356 = po51  & ~n8355;
  assign n8357 = ~po51  & n8355;
  assign n8358 = ~n7965 & ~n7966;
  assign n8359 = po22  & n8358;
  assign n8360 = ~n7971 & ~n8359;
  assign n8361 = n7971 & n8359;
  assign n8362 = ~n8360 & ~n8361;
  assign n8363 = ~n8357 & ~n8362;
  assign n8364 = ~n8356 & ~n8363;
  assign n8365 = po52  & ~n8364;
  assign n8366 = ~po52  & n8364;
  assign n8367 = ~n7974 & ~n7975;
  assign n8368 = po22  & n8367;
  assign n8369 = ~n7980 & ~n8368;
  assign n8370 = n7980 & n8368;
  assign n8371 = ~n8369 & ~n8370;
  assign n8372 = ~n8366 & ~n8371;
  assign n8373 = ~n8365 & ~n8372;
  assign n8374 = po53  & ~n8373;
  assign n8375 = ~po53  & n8373;
  assign n8376 = ~n7983 & ~n7984;
  assign n8377 = po22  & n8376;
  assign n8378 = ~n7989 & ~n8377;
  assign n8379 = n7989 & n8377;
  assign n8380 = ~n8378 & ~n8379;
  assign n8381 = ~n8375 & ~n8380;
  assign n8382 = ~n8374 & ~n8381;
  assign n8383 = po54  & ~n8382;
  assign n8384 = ~po54  & n8382;
  assign n8385 = ~n7992 & ~n7993;
  assign n8386 = po22  & n8385;
  assign n8387 = ~n7998 & ~n8386;
  assign n8388 = n7998 & n8386;
  assign n8389 = ~n8387 & ~n8388;
  assign n8390 = ~n8384 & ~n8389;
  assign n8391 = ~n8383 & ~n8390;
  assign n8392 = po55  & ~n8391;
  assign n8393 = ~po55  & n8391;
  assign n8394 = ~n8001 & ~n8002;
  assign n8395 = po22  & n8394;
  assign n8396 = ~n8007 & ~n8395;
  assign n8397 = n8007 & n8395;
  assign n8398 = ~n8396 & ~n8397;
  assign n8399 = ~n8393 & ~n8398;
  assign n8400 = ~n8392 & ~n8399;
  assign n8401 = po56  & ~n8400;
  assign n8402 = ~po56  & n8400;
  assign n8403 = ~n8010 & ~n8011;
  assign n8404 = po22  & n8403;
  assign n8405 = ~n8016 & ~n8404;
  assign n8406 = n8016 & n8404;
  assign n8407 = ~n8405 & ~n8406;
  assign n8408 = ~n8402 & ~n8407;
  assign n8409 = ~n8401 & ~n8408;
  assign n8410 = po57  & ~n8409;
  assign n8411 = ~po57  & n8409;
  assign n8412 = ~n8019 & ~n8020;
  assign n8413 = po22  & n8412;
  assign n8414 = ~n8025 & ~n8413;
  assign n8415 = n8025 & n8413;
  assign n8416 = ~n8414 & ~n8415;
  assign n8417 = ~n8411 & ~n8416;
  assign n8418 = ~n8410 & ~n8417;
  assign n8419 = po58  & ~n8418;
  assign n8420 = ~po58  & n8418;
  assign n8421 = ~n8028 & ~n8029;
  assign n8422 = po22  & n8421;
  assign n8423 = ~n8034 & ~n8422;
  assign n8424 = n8034 & n8422;
  assign n8425 = ~n8423 & ~n8424;
  assign n8426 = ~n8420 & ~n8425;
  assign n8427 = ~n8419 & ~n8426;
  assign n8428 = po59  & ~n8427;
  assign n8429 = ~po59  & n8427;
  assign n8430 = ~n8037 & ~n8038;
  assign n8431 = po22  & n8430;
  assign n8432 = ~n8043 & ~n8431;
  assign n8433 = n8043 & n8431;
  assign n8434 = ~n8432 & ~n8433;
  assign n8435 = ~n8429 & ~n8434;
  assign n8436 = ~n8428 & ~n8435;
  assign n8437 = po60  & ~n8436;
  assign n8438 = ~po60  & n8436;
  assign n8439 = ~n8046 & ~n8047;
  assign n8440 = po22  & n8439;
  assign n8441 = ~n8052 & ~n8440;
  assign n8442 = n8052 & n8440;
  assign n8443 = ~n8441 & ~n8442;
  assign n8444 = ~n8438 & ~n8443;
  assign n8445 = ~n8437 & ~n8444;
  assign n8446 = po61  & ~n8445;
  assign n8447 = ~po61  & n8445;
  assign n8448 = ~n8055 & ~n8056;
  assign n8449 = po22  & n8448;
  assign n8450 = ~n8061 & ~n8449;
  assign n8451 = n8061 & n8449;
  assign n8452 = ~n8450 & ~n8451;
  assign n8453 = ~n8447 & ~n8452;
  assign n8454 = ~n8446 & ~n8453;
  assign n8455 = po62  & ~n8454;
  assign n8456 = ~po62  & n8454;
  assign n8457 = ~n8064 & ~n8065;
  assign n8458 = po22  & n8457;
  assign n8459 = ~n8070 & ~n8458;
  assign n8460 = n8070 & n8458;
  assign n8461 = ~n8459 & ~n8460;
  assign n8462 = ~n8456 & ~n8461;
  assign n8463 = ~n8455 & ~n8462;
  assign n8464 = n8105 & n8463;
  assign n8465 = ~n8105 & ~n8463;
  assign n8466 = n8083 & po22 ;
  assign n8467 = ~n8082 & ~n8466;
  assign n8468 = n8465 & n8467;
  assign n8469 = ~po63  & ~n8468;
  assign n8470 = ~n8464 & ~n8469;
  assign n8471 = ~n8100 & n8470;
  assign po21  = n8096 | ~n8471;
  assign n8473 = ~n8289 & ~n8290;
  assign n8474 = po21  & n8473;
  assign n8475 = ~n8095 & ~n8474;
  assign n8476 = n8095 & n8474;
  assign n8477 = ~n8475 & ~n8476;
  assign n8478 = n8105 & ~po21 ;
  assign n8479 = ~n8105 & po21 ;
  assign n8480 = n8463 & ~n8479;
  assign n8481 = po63  & ~n8480;
  assign n8482 = ~n8465 & n8481;
  assign n8483 = ~n8455 & ~n8456;
  assign n8484 = po21  & n8483;
  assign n8485 = ~n8461 & ~n8484;
  assign n8486 = n8461 & n8484;
  assign n8487 = ~n8485 & ~n8486;
  assign n8488 = pi42  & po21 ;
  assign n8489 = ~pi40  & ~pi41 ;
  assign n8490 = ~pi42  & n8489;
  assign n8491 = ~n8488 & ~n8490;
  assign n8492 = po22  & ~n8491;
  assign n8493 = ~po22  & n8491;
  assign n8494 = ~pi42  & po21 ;
  assign n8495 = pi43  & ~n8494;
  assign n8496 = n8107 & po21 ;
  assign n8497 = ~n8495 & ~n8496;
  assign n8498 = ~n8493 & n8497;
  assign n8499 = ~n8492 & ~n8498;
  assign n8500 = po23  & ~n8499;
  assign n8501 = ~po23  & n8499;
  assign n8502 = po22  & n8471;
  assign n8503 = ~n8496 & ~n8502;
  assign n8504 = pi44  & ~n8503;
  assign n8505 = ~pi44  & n8503;
  assign n8506 = ~n8504 & ~n8505;
  assign n8507 = ~n8501 & ~n8506;
  assign n8508 = ~n8500 & ~n8507;
  assign n8509 = po24  & ~n8508;
  assign n8510 = ~po24  & n8508;
  assign n8511 = ~n8110 & ~n8111;
  assign n8512 = po21  & n8511;
  assign n8513 = n8115 & ~n8512;
  assign n8514 = ~n8115 & n8512;
  assign n8515 = ~n8513 & ~n8514;
  assign n8516 = ~n8510 & ~n8515;
  assign n8517 = ~n8509 & ~n8516;
  assign n8518 = po25  & ~n8517;
  assign n8519 = ~po25  & n8517;
  assign n8520 = ~n8118 & ~n8119;
  assign n8521 = po21  & n8520;
  assign n8522 = ~n8124 & ~n8521;
  assign n8523 = n8124 & n8521;
  assign n8524 = ~n8522 & ~n8523;
  assign n8525 = ~n8519 & ~n8524;
  assign n8526 = ~n8518 & ~n8525;
  assign n8527 = po26  & ~n8526;
  assign n8528 = ~po26  & n8526;
  assign n8529 = ~n8127 & ~n8128;
  assign n8530 = po21  & n8529;
  assign n8531 = n8133 & n8530;
  assign n8532 = ~n8133 & ~n8530;
  assign n8533 = ~n8531 & ~n8532;
  assign n8534 = ~n8528 & ~n8533;
  assign n8535 = ~n8527 & ~n8534;
  assign n8536 = po27  & ~n8535;
  assign n8537 = ~po27  & n8535;
  assign n8538 = ~n8136 & ~n8137;
  assign n8539 = po21  & n8538;
  assign n8540 = ~n8142 & ~n8539;
  assign n8541 = n8142 & n8539;
  assign n8542 = ~n8540 & ~n8541;
  assign n8543 = ~n8537 & ~n8542;
  assign n8544 = ~n8536 & ~n8543;
  assign n8545 = po28  & ~n8544;
  assign n8546 = ~po28  & n8544;
  assign n8547 = ~n8145 & ~n8146;
  assign n8548 = po21  & n8547;
  assign n8549 = ~n8151 & ~n8548;
  assign n8550 = n8151 & n8548;
  assign n8551 = ~n8549 & ~n8550;
  assign n8552 = ~n8546 & ~n8551;
  assign n8553 = ~n8545 & ~n8552;
  assign n8554 = po29  & ~n8553;
  assign n8555 = ~po29  & n8553;
  assign n8556 = ~n8154 & ~n8155;
  assign n8557 = po21  & n8556;
  assign n8558 = ~n8160 & ~n8557;
  assign n8559 = n8160 & n8557;
  assign n8560 = ~n8558 & ~n8559;
  assign n8561 = ~n8555 & ~n8560;
  assign n8562 = ~n8554 & ~n8561;
  assign n8563 = po30  & ~n8562;
  assign n8564 = ~po30  & n8562;
  assign n8565 = ~n8163 & ~n8164;
  assign n8566 = po21  & n8565;
  assign n8567 = ~n8169 & ~n8566;
  assign n8568 = n8169 & n8566;
  assign n8569 = ~n8567 & ~n8568;
  assign n8570 = ~n8564 & ~n8569;
  assign n8571 = ~n8563 & ~n8570;
  assign n8572 = po31  & ~n8571;
  assign n8573 = ~po31  & n8571;
  assign n8574 = ~n8172 & ~n8173;
  assign n8575 = po21  & n8574;
  assign n8576 = ~n8178 & ~n8575;
  assign n8577 = n8178 & n8575;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = ~n8573 & ~n8578;
  assign n8580 = ~n8572 & ~n8579;
  assign n8581 = po32  & ~n8580;
  assign n8582 = ~po32  & n8580;
  assign n8583 = ~n8181 & ~n8182;
  assign n8584 = po21  & n8583;
  assign n8585 = ~n8187 & ~n8584;
  assign n8586 = n8187 & n8584;
  assign n8587 = ~n8585 & ~n8586;
  assign n8588 = ~n8582 & ~n8587;
  assign n8589 = ~n8581 & ~n8588;
  assign n8590 = po33  & ~n8589;
  assign n8591 = ~po33  & n8589;
  assign n8592 = ~n8190 & ~n8191;
  assign n8593 = po21  & n8592;
  assign n8594 = ~n8196 & ~n8593;
  assign n8595 = n8196 & n8593;
  assign n8596 = ~n8594 & ~n8595;
  assign n8597 = ~n8591 & ~n8596;
  assign n8598 = ~n8590 & ~n8597;
  assign n8599 = po34  & ~n8598;
  assign n8600 = ~po34  & n8598;
  assign n8601 = ~n8199 & ~n8200;
  assign n8602 = po21  & n8601;
  assign n8603 = ~n8205 & ~n8602;
  assign n8604 = n8205 & n8602;
  assign n8605 = ~n8603 & ~n8604;
  assign n8606 = ~n8600 & ~n8605;
  assign n8607 = ~n8599 & ~n8606;
  assign n8608 = po35  & ~n8607;
  assign n8609 = ~po35  & n8607;
  assign n8610 = ~n8208 & ~n8209;
  assign n8611 = po21  & n8610;
  assign n8612 = ~n8214 & ~n8611;
  assign n8613 = n8214 & n8611;
  assign n8614 = ~n8612 & ~n8613;
  assign n8615 = ~n8609 & ~n8614;
  assign n8616 = ~n8608 & ~n8615;
  assign n8617 = po36  & ~n8616;
  assign n8618 = ~po36  & n8616;
  assign n8619 = ~n8217 & ~n8218;
  assign n8620 = po21  & n8619;
  assign n8621 = ~n8223 & ~n8620;
  assign n8622 = n8223 & n8620;
  assign n8623 = ~n8621 & ~n8622;
  assign n8624 = ~n8618 & ~n8623;
  assign n8625 = ~n8617 & ~n8624;
  assign n8626 = po37  & ~n8625;
  assign n8627 = ~po37  & n8625;
  assign n8628 = ~n8226 & ~n8227;
  assign n8629 = po21  & n8628;
  assign n8630 = ~n8232 & ~n8629;
  assign n8631 = n8232 & n8629;
  assign n8632 = ~n8630 & ~n8631;
  assign n8633 = ~n8627 & ~n8632;
  assign n8634 = ~n8626 & ~n8633;
  assign n8635 = po38  & ~n8634;
  assign n8636 = ~po38  & n8634;
  assign n8637 = ~n8235 & ~n8236;
  assign n8638 = po21  & n8637;
  assign n8639 = ~n8241 & ~n8638;
  assign n8640 = n8241 & n8638;
  assign n8641 = ~n8639 & ~n8640;
  assign n8642 = ~n8636 & ~n8641;
  assign n8643 = ~n8635 & ~n8642;
  assign n8644 = po39  & ~n8643;
  assign n8645 = ~po39  & n8643;
  assign n8646 = ~n8244 & ~n8245;
  assign n8647 = po21  & n8646;
  assign n8648 = ~n8250 & ~n8647;
  assign n8649 = n8250 & n8647;
  assign n8650 = ~n8648 & ~n8649;
  assign n8651 = ~n8645 & ~n8650;
  assign n8652 = ~n8644 & ~n8651;
  assign n8653 = po40  & ~n8652;
  assign n8654 = ~po40  & n8652;
  assign n8655 = ~n8253 & ~n8254;
  assign n8656 = po21  & n8655;
  assign n8657 = ~n8259 & ~n8656;
  assign n8658 = n8259 & n8656;
  assign n8659 = ~n8657 & ~n8658;
  assign n8660 = ~n8654 & ~n8659;
  assign n8661 = ~n8653 & ~n8660;
  assign n8662 = po41  & ~n8661;
  assign n8663 = ~po41  & n8661;
  assign n8664 = ~n8262 & ~n8263;
  assign n8665 = po21  & n8664;
  assign n8666 = ~n8268 & ~n8665;
  assign n8667 = n8268 & n8665;
  assign n8668 = ~n8666 & ~n8667;
  assign n8669 = ~n8663 & ~n8668;
  assign n8670 = ~n8662 & ~n8669;
  assign n8671 = po42  & ~n8670;
  assign n8672 = ~po42  & n8670;
  assign n8673 = ~n8271 & ~n8272;
  assign n8674 = po21  & n8673;
  assign n8675 = ~n8277 & ~n8674;
  assign n8676 = n8277 & n8674;
  assign n8677 = ~n8675 & ~n8676;
  assign n8678 = ~n8672 & ~n8677;
  assign n8679 = ~n8671 & ~n8678;
  assign n8680 = po43  & ~n8679;
  assign n8681 = ~n8280 & ~n8286;
  assign n8682 = po21  & n8681;
  assign n8683 = ~n8285 & ~n8682;
  assign n8684 = n8285 & n8682;
  assign n8685 = ~n8683 & ~n8684;
  assign n8686 = ~po43  & n8679;
  assign n8687 = ~n8685 & ~n8686;
  assign n8688 = ~n8680 & ~n8687;
  assign n8689 = po44  & ~n8688;
  assign n8690 = ~po44  & n8688;
  assign n8691 = ~n8477 & ~n8690;
  assign n8692 = ~n8689 & ~n8691;
  assign n8693 = po45  & ~n8692;
  assign n8694 = ~po45  & n8692;
  assign n8695 = ~n8293 & ~n8294;
  assign n8696 = po21  & n8695;
  assign n8697 = ~n8299 & ~n8696;
  assign n8698 = n8299 & n8696;
  assign n8699 = ~n8697 & ~n8698;
  assign n8700 = ~n8694 & ~n8699;
  assign n8701 = ~n8693 & ~n8700;
  assign n8702 = po46  & ~n8701;
  assign n8703 = ~po46  & n8701;
  assign n8704 = ~n8302 & ~n8303;
  assign n8705 = po21  & n8704;
  assign n8706 = ~n8308 & ~n8705;
  assign n8707 = n8308 & n8705;
  assign n8708 = ~n8706 & ~n8707;
  assign n8709 = ~n8703 & ~n8708;
  assign n8710 = ~n8702 & ~n8709;
  assign n8711 = po47  & ~n8710;
  assign n8712 = ~po47  & n8710;
  assign n8713 = ~n8311 & ~n8312;
  assign n8714 = po21  & n8713;
  assign n8715 = ~n8317 & ~n8714;
  assign n8716 = n8317 & n8714;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = ~n8712 & ~n8717;
  assign n8719 = ~n8711 & ~n8718;
  assign n8720 = po48  & ~n8719;
  assign n8721 = ~po48  & n8719;
  assign n8722 = ~n8320 & ~n8321;
  assign n8723 = po21  & n8722;
  assign n8724 = ~n8326 & ~n8723;
  assign n8725 = n8326 & n8723;
  assign n8726 = ~n8724 & ~n8725;
  assign n8727 = ~n8721 & ~n8726;
  assign n8728 = ~n8720 & ~n8727;
  assign n8729 = po49  & ~n8728;
  assign n8730 = ~po49  & n8728;
  assign n8731 = ~n8329 & ~n8330;
  assign n8732 = po21  & n8731;
  assign n8733 = ~n8335 & ~n8732;
  assign n8734 = n8335 & n8732;
  assign n8735 = ~n8733 & ~n8734;
  assign n8736 = ~n8730 & ~n8735;
  assign n8737 = ~n8729 & ~n8736;
  assign n8738 = po50  & ~n8737;
  assign n8739 = ~po50  & n8737;
  assign n8740 = ~n8338 & ~n8339;
  assign n8741 = po21  & n8740;
  assign n8742 = ~n8344 & ~n8741;
  assign n8743 = n8344 & n8741;
  assign n8744 = ~n8742 & ~n8743;
  assign n8745 = ~n8739 & ~n8744;
  assign n8746 = ~n8738 & ~n8745;
  assign n8747 = po51  & ~n8746;
  assign n8748 = ~po51  & n8746;
  assign n8749 = ~n8347 & ~n8348;
  assign n8750 = po21  & n8749;
  assign n8751 = ~n8353 & ~n8750;
  assign n8752 = n8353 & n8750;
  assign n8753 = ~n8751 & ~n8752;
  assign n8754 = ~n8748 & ~n8753;
  assign n8755 = ~n8747 & ~n8754;
  assign n8756 = po52  & ~n8755;
  assign n8757 = ~po52  & n8755;
  assign n8758 = ~n8356 & ~n8357;
  assign n8759 = po21  & n8758;
  assign n8760 = ~n8362 & ~n8759;
  assign n8761 = n8362 & n8759;
  assign n8762 = ~n8760 & ~n8761;
  assign n8763 = ~n8757 & ~n8762;
  assign n8764 = ~n8756 & ~n8763;
  assign n8765 = po53  & ~n8764;
  assign n8766 = ~po53  & n8764;
  assign n8767 = ~n8365 & ~n8366;
  assign n8768 = po21  & n8767;
  assign n8769 = ~n8371 & ~n8768;
  assign n8770 = n8371 & n8768;
  assign n8771 = ~n8769 & ~n8770;
  assign n8772 = ~n8766 & ~n8771;
  assign n8773 = ~n8765 & ~n8772;
  assign n8774 = po54  & ~n8773;
  assign n8775 = ~po54  & n8773;
  assign n8776 = ~n8374 & ~n8375;
  assign n8777 = po21  & n8776;
  assign n8778 = ~n8380 & ~n8777;
  assign n8779 = n8380 & n8777;
  assign n8780 = ~n8778 & ~n8779;
  assign n8781 = ~n8775 & ~n8780;
  assign n8782 = ~n8774 & ~n8781;
  assign n8783 = po55  & ~n8782;
  assign n8784 = ~po55  & n8782;
  assign n8785 = ~n8383 & ~n8384;
  assign n8786 = po21  & n8785;
  assign n8787 = ~n8389 & ~n8786;
  assign n8788 = n8389 & n8786;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = ~n8784 & ~n8789;
  assign n8791 = ~n8783 & ~n8790;
  assign n8792 = po56  & ~n8791;
  assign n8793 = ~po56  & n8791;
  assign n8794 = ~n8392 & ~n8393;
  assign n8795 = po21  & n8794;
  assign n8796 = ~n8398 & ~n8795;
  assign n8797 = n8398 & n8795;
  assign n8798 = ~n8796 & ~n8797;
  assign n8799 = ~n8793 & ~n8798;
  assign n8800 = ~n8792 & ~n8799;
  assign n8801 = po57  & ~n8800;
  assign n8802 = ~po57  & n8800;
  assign n8803 = ~n8401 & ~n8402;
  assign n8804 = po21  & n8803;
  assign n8805 = ~n8407 & ~n8804;
  assign n8806 = n8407 & n8804;
  assign n8807 = ~n8805 & ~n8806;
  assign n8808 = ~n8802 & ~n8807;
  assign n8809 = ~n8801 & ~n8808;
  assign n8810 = po58  & ~n8809;
  assign n8811 = ~po58  & n8809;
  assign n8812 = ~n8410 & ~n8411;
  assign n8813 = po21  & n8812;
  assign n8814 = ~n8416 & ~n8813;
  assign n8815 = n8416 & n8813;
  assign n8816 = ~n8814 & ~n8815;
  assign n8817 = ~n8811 & ~n8816;
  assign n8818 = ~n8810 & ~n8817;
  assign n8819 = po59  & ~n8818;
  assign n8820 = ~po59  & n8818;
  assign n8821 = ~n8419 & ~n8420;
  assign n8822 = po21  & n8821;
  assign n8823 = ~n8425 & ~n8822;
  assign n8824 = n8425 & n8822;
  assign n8825 = ~n8823 & ~n8824;
  assign n8826 = ~n8820 & ~n8825;
  assign n8827 = ~n8819 & ~n8826;
  assign n8828 = po60  & ~n8827;
  assign n8829 = ~po60  & n8827;
  assign n8830 = ~n8428 & ~n8429;
  assign n8831 = po21  & n8830;
  assign n8832 = ~n8434 & ~n8831;
  assign n8833 = n8434 & n8831;
  assign n8834 = ~n8832 & ~n8833;
  assign n8835 = ~n8829 & ~n8834;
  assign n8836 = ~n8828 & ~n8835;
  assign n8837 = po61  & ~n8836;
  assign n8838 = ~po61  & n8836;
  assign n8839 = ~n8437 & ~n8438;
  assign n8840 = po21  & n8839;
  assign n8841 = ~n8443 & ~n8840;
  assign n8842 = n8443 & n8840;
  assign n8843 = ~n8841 & ~n8842;
  assign n8844 = ~n8838 & ~n8843;
  assign n8845 = ~n8837 & ~n8844;
  assign n8846 = po62  & ~n8845;
  assign n8847 = ~po62  & n8845;
  assign n8848 = ~n8446 & ~n8447;
  assign n8849 = po21  & n8848;
  assign n8850 = ~n8452 & ~n8849;
  assign n8851 = n8452 & n8849;
  assign n8852 = ~n8850 & ~n8851;
  assign n8853 = ~n8847 & ~n8852;
  assign n8854 = ~n8846 & ~n8853;
  assign n8855 = n8487 & n8854;
  assign n8856 = ~n8487 & ~n8854;
  assign n8857 = n8465 & po21 ;
  assign n8858 = ~n8464 & ~n8857;
  assign n8859 = n8856 & n8858;
  assign n8860 = ~po63  & ~n8859;
  assign n8861 = ~n8855 & ~n8860;
  assign n8862 = ~n8482 & n8861;
  assign po20  = n8478 | ~n8862;
  assign n8864 = ~n8689 & ~n8690;
  assign n8865 = po20  & n8864;
  assign n8866 = ~n8477 & ~n8865;
  assign n8867 = n8477 & n8865;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = n8487 & ~po20 ;
  assign n8870 = ~n8487 & po20 ;
  assign n8871 = n8854 & ~n8870;
  assign n8872 = po63  & ~n8871;
  assign n8873 = ~n8856 & n8872;
  assign n8874 = ~n8846 & ~n8847;
  assign n8875 = po20  & n8874;
  assign n8876 = ~n8852 & ~n8875;
  assign n8877 = n8852 & n8875;
  assign n8878 = ~n8876 & ~n8877;
  assign n8879 = pi40  & po20 ;
  assign n8880 = ~pi38  & ~pi39 ;
  assign n8881 = ~pi40  & n8880;
  assign n8882 = ~n8879 & ~n8881;
  assign n8883 = po21  & ~n8882;
  assign n8884 = ~po21  & n8882;
  assign n8885 = ~pi40  & po20 ;
  assign n8886 = pi41  & ~n8885;
  assign n8887 = n8489 & po20 ;
  assign n8888 = ~n8886 & ~n8887;
  assign n8889 = ~n8884 & n8888;
  assign n8890 = ~n8883 & ~n8889;
  assign n8891 = po22  & ~n8890;
  assign n8892 = ~po22  & n8890;
  assign n8893 = po21  & n8862;
  assign n8894 = ~n8887 & ~n8893;
  assign n8895 = pi42  & ~n8894;
  assign n8896 = ~pi42  & n8894;
  assign n8897 = ~n8895 & ~n8896;
  assign n8898 = ~n8892 & ~n8897;
  assign n8899 = ~n8891 & ~n8898;
  assign n8900 = po23  & ~n8899;
  assign n8901 = ~po23  & n8899;
  assign n8902 = ~n8492 & ~n8493;
  assign n8903 = po20  & n8902;
  assign n8904 = n8497 & ~n8903;
  assign n8905 = ~n8497 & n8903;
  assign n8906 = ~n8904 & ~n8905;
  assign n8907 = ~n8901 & ~n8906;
  assign n8908 = ~n8900 & ~n8907;
  assign n8909 = po24  & ~n8908;
  assign n8910 = ~po24  & n8908;
  assign n8911 = ~n8500 & ~n8501;
  assign n8912 = po20  & n8911;
  assign n8913 = ~n8506 & ~n8912;
  assign n8914 = n8506 & n8912;
  assign n8915 = ~n8913 & ~n8914;
  assign n8916 = ~n8910 & ~n8915;
  assign n8917 = ~n8909 & ~n8916;
  assign n8918 = po25  & ~n8917;
  assign n8919 = ~po25  & n8917;
  assign n8920 = ~n8509 & ~n8510;
  assign n8921 = po20  & n8920;
  assign n8922 = n8515 & n8921;
  assign n8923 = ~n8515 & ~n8921;
  assign n8924 = ~n8922 & ~n8923;
  assign n8925 = ~n8919 & ~n8924;
  assign n8926 = ~n8918 & ~n8925;
  assign n8927 = po26  & ~n8926;
  assign n8928 = ~po26  & n8926;
  assign n8929 = ~n8518 & ~n8519;
  assign n8930 = po20  & n8929;
  assign n8931 = ~n8524 & ~n8930;
  assign n8932 = n8524 & n8930;
  assign n8933 = ~n8931 & ~n8932;
  assign n8934 = ~n8928 & ~n8933;
  assign n8935 = ~n8927 & ~n8934;
  assign n8936 = po27  & ~n8935;
  assign n8937 = ~po27  & n8935;
  assign n8938 = ~n8527 & ~n8528;
  assign n8939 = po20  & n8938;
  assign n8940 = ~n8533 & ~n8939;
  assign n8941 = n8533 & n8939;
  assign n8942 = ~n8940 & ~n8941;
  assign n8943 = ~n8937 & ~n8942;
  assign n8944 = ~n8936 & ~n8943;
  assign n8945 = po28  & ~n8944;
  assign n8946 = ~po28  & n8944;
  assign n8947 = ~n8536 & ~n8537;
  assign n8948 = po20  & n8947;
  assign n8949 = ~n8542 & ~n8948;
  assign n8950 = n8542 & n8948;
  assign n8951 = ~n8949 & ~n8950;
  assign n8952 = ~n8946 & ~n8951;
  assign n8953 = ~n8945 & ~n8952;
  assign n8954 = po29  & ~n8953;
  assign n8955 = ~po29  & n8953;
  assign n8956 = ~n8545 & ~n8546;
  assign n8957 = po20  & n8956;
  assign n8958 = ~n8551 & ~n8957;
  assign n8959 = n8551 & n8957;
  assign n8960 = ~n8958 & ~n8959;
  assign n8961 = ~n8955 & ~n8960;
  assign n8962 = ~n8954 & ~n8961;
  assign n8963 = po30  & ~n8962;
  assign n8964 = ~po30  & n8962;
  assign n8965 = ~n8554 & ~n8555;
  assign n8966 = po20  & n8965;
  assign n8967 = ~n8560 & ~n8966;
  assign n8968 = n8560 & n8966;
  assign n8969 = ~n8967 & ~n8968;
  assign n8970 = ~n8964 & ~n8969;
  assign n8971 = ~n8963 & ~n8970;
  assign n8972 = po31  & ~n8971;
  assign n8973 = ~po31  & n8971;
  assign n8974 = ~n8563 & ~n8564;
  assign n8975 = po20  & n8974;
  assign n8976 = ~n8569 & ~n8975;
  assign n8977 = n8569 & n8975;
  assign n8978 = ~n8976 & ~n8977;
  assign n8979 = ~n8973 & ~n8978;
  assign n8980 = ~n8972 & ~n8979;
  assign n8981 = po32  & ~n8980;
  assign n8982 = ~po32  & n8980;
  assign n8983 = ~n8572 & ~n8573;
  assign n8984 = po20  & n8983;
  assign n8985 = ~n8578 & ~n8984;
  assign n8986 = n8578 & n8984;
  assign n8987 = ~n8985 & ~n8986;
  assign n8988 = ~n8982 & ~n8987;
  assign n8989 = ~n8981 & ~n8988;
  assign n8990 = po33  & ~n8989;
  assign n8991 = ~po33  & n8989;
  assign n8992 = ~n8581 & ~n8582;
  assign n8993 = po20  & n8992;
  assign n8994 = ~n8587 & ~n8993;
  assign n8995 = n8587 & n8993;
  assign n8996 = ~n8994 & ~n8995;
  assign n8997 = ~n8991 & ~n8996;
  assign n8998 = ~n8990 & ~n8997;
  assign n8999 = po34  & ~n8998;
  assign n9000 = ~po34  & n8998;
  assign n9001 = ~n8590 & ~n8591;
  assign n9002 = po20  & n9001;
  assign n9003 = ~n8596 & ~n9002;
  assign n9004 = n8596 & n9002;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = ~n9000 & ~n9005;
  assign n9007 = ~n8999 & ~n9006;
  assign n9008 = po35  & ~n9007;
  assign n9009 = ~po35  & n9007;
  assign n9010 = ~n8599 & ~n8600;
  assign n9011 = po20  & n9010;
  assign n9012 = ~n8605 & ~n9011;
  assign n9013 = n8605 & n9011;
  assign n9014 = ~n9012 & ~n9013;
  assign n9015 = ~n9009 & ~n9014;
  assign n9016 = ~n9008 & ~n9015;
  assign n9017 = po36  & ~n9016;
  assign n9018 = ~po36  & n9016;
  assign n9019 = ~n8608 & ~n8609;
  assign n9020 = po20  & n9019;
  assign n9021 = ~n8614 & ~n9020;
  assign n9022 = n8614 & n9020;
  assign n9023 = ~n9021 & ~n9022;
  assign n9024 = ~n9018 & ~n9023;
  assign n9025 = ~n9017 & ~n9024;
  assign n9026 = po37  & ~n9025;
  assign n9027 = ~po37  & n9025;
  assign n9028 = ~n8617 & ~n8618;
  assign n9029 = po20  & n9028;
  assign n9030 = ~n8623 & ~n9029;
  assign n9031 = n8623 & n9029;
  assign n9032 = ~n9030 & ~n9031;
  assign n9033 = ~n9027 & ~n9032;
  assign n9034 = ~n9026 & ~n9033;
  assign n9035 = po38  & ~n9034;
  assign n9036 = ~po38  & n9034;
  assign n9037 = ~n8626 & ~n8627;
  assign n9038 = po20  & n9037;
  assign n9039 = ~n8632 & ~n9038;
  assign n9040 = n8632 & n9038;
  assign n9041 = ~n9039 & ~n9040;
  assign n9042 = ~n9036 & ~n9041;
  assign n9043 = ~n9035 & ~n9042;
  assign n9044 = po39  & ~n9043;
  assign n9045 = ~po39  & n9043;
  assign n9046 = ~n8635 & ~n8636;
  assign n9047 = po20  & n9046;
  assign n9048 = ~n8641 & ~n9047;
  assign n9049 = n8641 & n9047;
  assign n9050 = ~n9048 & ~n9049;
  assign n9051 = ~n9045 & ~n9050;
  assign n9052 = ~n9044 & ~n9051;
  assign n9053 = po40  & ~n9052;
  assign n9054 = ~po40  & n9052;
  assign n9055 = ~n8644 & ~n8645;
  assign n9056 = po20  & n9055;
  assign n9057 = ~n8650 & ~n9056;
  assign n9058 = n8650 & n9056;
  assign n9059 = ~n9057 & ~n9058;
  assign n9060 = ~n9054 & ~n9059;
  assign n9061 = ~n9053 & ~n9060;
  assign n9062 = po41  & ~n9061;
  assign n9063 = ~po41  & n9061;
  assign n9064 = ~n8653 & ~n8654;
  assign n9065 = po20  & n9064;
  assign n9066 = ~n8659 & ~n9065;
  assign n9067 = n8659 & n9065;
  assign n9068 = ~n9066 & ~n9067;
  assign n9069 = ~n9063 & ~n9068;
  assign n9070 = ~n9062 & ~n9069;
  assign n9071 = po42  & ~n9070;
  assign n9072 = ~po42  & n9070;
  assign n9073 = ~n8662 & ~n8663;
  assign n9074 = po20  & n9073;
  assign n9075 = ~n8668 & ~n9074;
  assign n9076 = n8668 & n9074;
  assign n9077 = ~n9075 & ~n9076;
  assign n9078 = ~n9072 & ~n9077;
  assign n9079 = ~n9071 & ~n9078;
  assign n9080 = po43  & ~n9079;
  assign n9081 = ~po43  & n9079;
  assign n9082 = ~n8671 & ~n8672;
  assign n9083 = po20  & n9082;
  assign n9084 = ~n8677 & ~n9083;
  assign n9085 = n8677 & n9083;
  assign n9086 = ~n9084 & ~n9085;
  assign n9087 = ~n9081 & ~n9086;
  assign n9088 = ~n9080 & ~n9087;
  assign n9089 = po44  & ~n9088;
  assign n9090 = ~n8680 & ~n8686;
  assign n9091 = po20  & n9090;
  assign n9092 = ~n8685 & ~n9091;
  assign n9093 = n8685 & n9091;
  assign n9094 = ~n9092 & ~n9093;
  assign n9095 = ~po44  & n9088;
  assign n9096 = ~n9094 & ~n9095;
  assign n9097 = ~n9089 & ~n9096;
  assign n9098 = po45  & ~n9097;
  assign n9099 = ~po45  & n9097;
  assign n9100 = ~n8868 & ~n9099;
  assign n9101 = ~n9098 & ~n9100;
  assign n9102 = po46  & ~n9101;
  assign n9103 = ~po46  & n9101;
  assign n9104 = ~n8693 & ~n8694;
  assign n9105 = po20  & n9104;
  assign n9106 = ~n8699 & ~n9105;
  assign n9107 = n8699 & n9105;
  assign n9108 = ~n9106 & ~n9107;
  assign n9109 = ~n9103 & ~n9108;
  assign n9110 = ~n9102 & ~n9109;
  assign n9111 = po47  & ~n9110;
  assign n9112 = ~po47  & n9110;
  assign n9113 = ~n8702 & ~n8703;
  assign n9114 = po20  & n9113;
  assign n9115 = ~n8708 & ~n9114;
  assign n9116 = n8708 & n9114;
  assign n9117 = ~n9115 & ~n9116;
  assign n9118 = ~n9112 & ~n9117;
  assign n9119 = ~n9111 & ~n9118;
  assign n9120 = po48  & ~n9119;
  assign n9121 = ~po48  & n9119;
  assign n9122 = ~n8711 & ~n8712;
  assign n9123 = po20  & n9122;
  assign n9124 = ~n8717 & ~n9123;
  assign n9125 = n8717 & n9123;
  assign n9126 = ~n9124 & ~n9125;
  assign n9127 = ~n9121 & ~n9126;
  assign n9128 = ~n9120 & ~n9127;
  assign n9129 = po49  & ~n9128;
  assign n9130 = ~po49  & n9128;
  assign n9131 = ~n8720 & ~n8721;
  assign n9132 = po20  & n9131;
  assign n9133 = ~n8726 & ~n9132;
  assign n9134 = n8726 & n9132;
  assign n9135 = ~n9133 & ~n9134;
  assign n9136 = ~n9130 & ~n9135;
  assign n9137 = ~n9129 & ~n9136;
  assign n9138 = po50  & ~n9137;
  assign n9139 = ~po50  & n9137;
  assign n9140 = ~n8729 & ~n8730;
  assign n9141 = po20  & n9140;
  assign n9142 = ~n8735 & ~n9141;
  assign n9143 = n8735 & n9141;
  assign n9144 = ~n9142 & ~n9143;
  assign n9145 = ~n9139 & ~n9144;
  assign n9146 = ~n9138 & ~n9145;
  assign n9147 = po51  & ~n9146;
  assign n9148 = ~po51  & n9146;
  assign n9149 = ~n8738 & ~n8739;
  assign n9150 = po20  & n9149;
  assign n9151 = ~n8744 & ~n9150;
  assign n9152 = n8744 & n9150;
  assign n9153 = ~n9151 & ~n9152;
  assign n9154 = ~n9148 & ~n9153;
  assign n9155 = ~n9147 & ~n9154;
  assign n9156 = po52  & ~n9155;
  assign n9157 = ~po52  & n9155;
  assign n9158 = ~n8747 & ~n8748;
  assign n9159 = po20  & n9158;
  assign n9160 = ~n8753 & ~n9159;
  assign n9161 = n8753 & n9159;
  assign n9162 = ~n9160 & ~n9161;
  assign n9163 = ~n9157 & ~n9162;
  assign n9164 = ~n9156 & ~n9163;
  assign n9165 = po53  & ~n9164;
  assign n9166 = ~po53  & n9164;
  assign n9167 = ~n8756 & ~n8757;
  assign n9168 = po20  & n9167;
  assign n9169 = ~n8762 & ~n9168;
  assign n9170 = n8762 & n9168;
  assign n9171 = ~n9169 & ~n9170;
  assign n9172 = ~n9166 & ~n9171;
  assign n9173 = ~n9165 & ~n9172;
  assign n9174 = po54  & ~n9173;
  assign n9175 = ~po54  & n9173;
  assign n9176 = ~n8765 & ~n8766;
  assign n9177 = po20  & n9176;
  assign n9178 = ~n8771 & ~n9177;
  assign n9179 = n8771 & n9177;
  assign n9180 = ~n9178 & ~n9179;
  assign n9181 = ~n9175 & ~n9180;
  assign n9182 = ~n9174 & ~n9181;
  assign n9183 = po55  & ~n9182;
  assign n9184 = ~po55  & n9182;
  assign n9185 = ~n8774 & ~n8775;
  assign n9186 = po20  & n9185;
  assign n9187 = ~n8780 & ~n9186;
  assign n9188 = n8780 & n9186;
  assign n9189 = ~n9187 & ~n9188;
  assign n9190 = ~n9184 & ~n9189;
  assign n9191 = ~n9183 & ~n9190;
  assign n9192 = po56  & ~n9191;
  assign n9193 = ~po56  & n9191;
  assign n9194 = ~n8783 & ~n8784;
  assign n9195 = po20  & n9194;
  assign n9196 = ~n8789 & ~n9195;
  assign n9197 = n8789 & n9195;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = ~n9193 & ~n9198;
  assign n9200 = ~n9192 & ~n9199;
  assign n9201 = po57  & ~n9200;
  assign n9202 = ~po57  & n9200;
  assign n9203 = ~n8792 & ~n8793;
  assign n9204 = po20  & n9203;
  assign n9205 = ~n8798 & ~n9204;
  assign n9206 = n8798 & n9204;
  assign n9207 = ~n9205 & ~n9206;
  assign n9208 = ~n9202 & ~n9207;
  assign n9209 = ~n9201 & ~n9208;
  assign n9210 = po58  & ~n9209;
  assign n9211 = ~po58  & n9209;
  assign n9212 = ~n8801 & ~n8802;
  assign n9213 = po20  & n9212;
  assign n9214 = ~n8807 & ~n9213;
  assign n9215 = n8807 & n9213;
  assign n9216 = ~n9214 & ~n9215;
  assign n9217 = ~n9211 & ~n9216;
  assign n9218 = ~n9210 & ~n9217;
  assign n9219 = po59  & ~n9218;
  assign n9220 = ~po59  & n9218;
  assign n9221 = ~n8810 & ~n8811;
  assign n9222 = po20  & n9221;
  assign n9223 = ~n8816 & ~n9222;
  assign n9224 = n8816 & n9222;
  assign n9225 = ~n9223 & ~n9224;
  assign n9226 = ~n9220 & ~n9225;
  assign n9227 = ~n9219 & ~n9226;
  assign n9228 = po60  & ~n9227;
  assign n9229 = ~po60  & n9227;
  assign n9230 = ~n8819 & ~n8820;
  assign n9231 = po20  & n9230;
  assign n9232 = ~n8825 & ~n9231;
  assign n9233 = n8825 & n9231;
  assign n9234 = ~n9232 & ~n9233;
  assign n9235 = ~n9229 & ~n9234;
  assign n9236 = ~n9228 & ~n9235;
  assign n9237 = po61  & ~n9236;
  assign n9238 = ~po61  & n9236;
  assign n9239 = ~n8828 & ~n8829;
  assign n9240 = po20  & n9239;
  assign n9241 = ~n8834 & ~n9240;
  assign n9242 = n8834 & n9240;
  assign n9243 = ~n9241 & ~n9242;
  assign n9244 = ~n9238 & ~n9243;
  assign n9245 = ~n9237 & ~n9244;
  assign n9246 = po62  & ~n9245;
  assign n9247 = ~po62  & n9245;
  assign n9248 = ~n8837 & ~n8838;
  assign n9249 = po20  & n9248;
  assign n9250 = ~n8843 & ~n9249;
  assign n9251 = n8843 & n9249;
  assign n9252 = ~n9250 & ~n9251;
  assign n9253 = ~n9247 & ~n9252;
  assign n9254 = ~n9246 & ~n9253;
  assign n9255 = n8878 & n9254;
  assign n9256 = ~n8878 & ~n9254;
  assign n9257 = n8856 & po20 ;
  assign n9258 = ~n8855 & ~n9257;
  assign n9259 = n9256 & n9258;
  assign n9260 = ~po63  & ~n9259;
  assign n9261 = ~n9255 & ~n9260;
  assign n9262 = ~n8873 & n9261;
  assign po19  = n8869 | ~n9262;
  assign n9264 = ~n9098 & ~n9099;
  assign n9265 = po19  & n9264;
  assign n9266 = ~n8868 & ~n9265;
  assign n9267 = n8868 & n9265;
  assign n9268 = ~n9266 & ~n9267;
  assign n9269 = n8878 & ~po19 ;
  assign n9270 = ~n8878 & po19 ;
  assign n9271 = n9254 & ~n9270;
  assign n9272 = po63  & ~n9271;
  assign n9273 = ~n9256 & n9272;
  assign n9274 = ~n9246 & ~n9247;
  assign n9275 = po19  & n9274;
  assign n9276 = ~n9252 & ~n9275;
  assign n9277 = n9252 & n9275;
  assign n9278 = ~n9276 & ~n9277;
  assign n9279 = pi38  & po19 ;
  assign n9280 = ~pi36  & ~pi37 ;
  assign n9281 = ~pi38  & n9280;
  assign n9282 = ~n9279 & ~n9281;
  assign n9283 = po20  & ~n9282;
  assign n9284 = ~po20  & n9282;
  assign n9285 = ~pi38  & po19 ;
  assign n9286 = pi39  & ~n9285;
  assign n9287 = n8880 & po19 ;
  assign n9288 = ~n9286 & ~n9287;
  assign n9289 = ~n9284 & n9288;
  assign n9290 = ~n9283 & ~n9289;
  assign n9291 = po21  & ~n9290;
  assign n9292 = ~po21  & n9290;
  assign n9293 = po20  & n9262;
  assign n9294 = ~n9287 & ~n9293;
  assign n9295 = pi40  & ~n9294;
  assign n9296 = ~pi40  & n9294;
  assign n9297 = ~n9295 & ~n9296;
  assign n9298 = ~n9292 & ~n9297;
  assign n9299 = ~n9291 & ~n9298;
  assign n9300 = po22  & ~n9299;
  assign n9301 = ~po22  & n9299;
  assign n9302 = ~n8883 & ~n8884;
  assign n9303 = po19  & n9302;
  assign n9304 = n8888 & ~n9303;
  assign n9305 = ~n8888 & n9303;
  assign n9306 = ~n9304 & ~n9305;
  assign n9307 = ~n9301 & ~n9306;
  assign n9308 = ~n9300 & ~n9307;
  assign n9309 = po23  & ~n9308;
  assign n9310 = ~po23  & n9308;
  assign n9311 = ~n8891 & ~n8892;
  assign n9312 = po19  & n9311;
  assign n9313 = ~n8897 & ~n9312;
  assign n9314 = n8897 & n9312;
  assign n9315 = ~n9313 & ~n9314;
  assign n9316 = ~n9310 & ~n9315;
  assign n9317 = ~n9309 & ~n9316;
  assign n9318 = po24  & ~n9317;
  assign n9319 = ~po24  & n9317;
  assign n9320 = ~n8900 & ~n8901;
  assign n9321 = po19  & n9320;
  assign n9322 = n8906 & n9321;
  assign n9323 = ~n8906 & ~n9321;
  assign n9324 = ~n9322 & ~n9323;
  assign n9325 = ~n9319 & ~n9324;
  assign n9326 = ~n9318 & ~n9325;
  assign n9327 = po25  & ~n9326;
  assign n9328 = ~po25  & n9326;
  assign n9329 = ~n8909 & ~n8910;
  assign n9330 = po19  & n9329;
  assign n9331 = ~n8915 & ~n9330;
  assign n9332 = n8915 & n9330;
  assign n9333 = ~n9331 & ~n9332;
  assign n9334 = ~n9328 & ~n9333;
  assign n9335 = ~n9327 & ~n9334;
  assign n9336 = po26  & ~n9335;
  assign n9337 = ~po26  & n9335;
  assign n9338 = ~n8918 & ~n8919;
  assign n9339 = po19  & n9338;
  assign n9340 = ~n8924 & ~n9339;
  assign n9341 = n8924 & n9339;
  assign n9342 = ~n9340 & ~n9341;
  assign n9343 = ~n9337 & ~n9342;
  assign n9344 = ~n9336 & ~n9343;
  assign n9345 = po27  & ~n9344;
  assign n9346 = ~po27  & n9344;
  assign n9347 = ~n8927 & ~n8928;
  assign n9348 = po19  & n9347;
  assign n9349 = ~n8933 & ~n9348;
  assign n9350 = n8933 & n9348;
  assign n9351 = ~n9349 & ~n9350;
  assign n9352 = ~n9346 & ~n9351;
  assign n9353 = ~n9345 & ~n9352;
  assign n9354 = po28  & ~n9353;
  assign n9355 = ~po28  & n9353;
  assign n9356 = ~n8936 & ~n8937;
  assign n9357 = po19  & n9356;
  assign n9358 = ~n8942 & ~n9357;
  assign n9359 = n8942 & n9357;
  assign n9360 = ~n9358 & ~n9359;
  assign n9361 = ~n9355 & ~n9360;
  assign n9362 = ~n9354 & ~n9361;
  assign n9363 = po29  & ~n9362;
  assign n9364 = ~po29  & n9362;
  assign n9365 = ~n8945 & ~n8946;
  assign n9366 = po19  & n9365;
  assign n9367 = ~n8951 & ~n9366;
  assign n9368 = n8951 & n9366;
  assign n9369 = ~n9367 & ~n9368;
  assign n9370 = ~n9364 & ~n9369;
  assign n9371 = ~n9363 & ~n9370;
  assign n9372 = po30  & ~n9371;
  assign n9373 = ~po30  & n9371;
  assign n9374 = ~n8954 & ~n8955;
  assign n9375 = po19  & n9374;
  assign n9376 = ~n8960 & ~n9375;
  assign n9377 = n8960 & n9375;
  assign n9378 = ~n9376 & ~n9377;
  assign n9379 = ~n9373 & ~n9378;
  assign n9380 = ~n9372 & ~n9379;
  assign n9381 = po31  & ~n9380;
  assign n9382 = ~po31  & n9380;
  assign n9383 = ~n8963 & ~n8964;
  assign n9384 = po19  & n9383;
  assign n9385 = ~n8969 & ~n9384;
  assign n9386 = n8969 & n9384;
  assign n9387 = ~n9385 & ~n9386;
  assign n9388 = ~n9382 & ~n9387;
  assign n9389 = ~n9381 & ~n9388;
  assign n9390 = po32  & ~n9389;
  assign n9391 = ~po32  & n9389;
  assign n9392 = ~n8972 & ~n8973;
  assign n9393 = po19  & n9392;
  assign n9394 = ~n8978 & ~n9393;
  assign n9395 = n8978 & n9393;
  assign n9396 = ~n9394 & ~n9395;
  assign n9397 = ~n9391 & ~n9396;
  assign n9398 = ~n9390 & ~n9397;
  assign n9399 = po33  & ~n9398;
  assign n9400 = ~po33  & n9398;
  assign n9401 = ~n8981 & ~n8982;
  assign n9402 = po19  & n9401;
  assign n9403 = ~n8987 & ~n9402;
  assign n9404 = n8987 & n9402;
  assign n9405 = ~n9403 & ~n9404;
  assign n9406 = ~n9400 & ~n9405;
  assign n9407 = ~n9399 & ~n9406;
  assign n9408 = po34  & ~n9407;
  assign n9409 = ~po34  & n9407;
  assign n9410 = ~n8990 & ~n8991;
  assign n9411 = po19  & n9410;
  assign n9412 = ~n8996 & ~n9411;
  assign n9413 = n8996 & n9411;
  assign n9414 = ~n9412 & ~n9413;
  assign n9415 = ~n9409 & ~n9414;
  assign n9416 = ~n9408 & ~n9415;
  assign n9417 = po35  & ~n9416;
  assign n9418 = ~po35  & n9416;
  assign n9419 = ~n8999 & ~n9000;
  assign n9420 = po19  & n9419;
  assign n9421 = ~n9005 & ~n9420;
  assign n9422 = n9005 & n9420;
  assign n9423 = ~n9421 & ~n9422;
  assign n9424 = ~n9418 & ~n9423;
  assign n9425 = ~n9417 & ~n9424;
  assign n9426 = po36  & ~n9425;
  assign n9427 = ~po36  & n9425;
  assign n9428 = ~n9008 & ~n9009;
  assign n9429 = po19  & n9428;
  assign n9430 = ~n9014 & ~n9429;
  assign n9431 = n9014 & n9429;
  assign n9432 = ~n9430 & ~n9431;
  assign n9433 = ~n9427 & ~n9432;
  assign n9434 = ~n9426 & ~n9433;
  assign n9435 = po37  & ~n9434;
  assign n9436 = ~po37  & n9434;
  assign n9437 = ~n9017 & ~n9018;
  assign n9438 = po19  & n9437;
  assign n9439 = ~n9023 & ~n9438;
  assign n9440 = n9023 & n9438;
  assign n9441 = ~n9439 & ~n9440;
  assign n9442 = ~n9436 & ~n9441;
  assign n9443 = ~n9435 & ~n9442;
  assign n9444 = po38  & ~n9443;
  assign n9445 = ~po38  & n9443;
  assign n9446 = ~n9026 & ~n9027;
  assign n9447 = po19  & n9446;
  assign n9448 = ~n9032 & ~n9447;
  assign n9449 = n9032 & n9447;
  assign n9450 = ~n9448 & ~n9449;
  assign n9451 = ~n9445 & ~n9450;
  assign n9452 = ~n9444 & ~n9451;
  assign n9453 = po39  & ~n9452;
  assign n9454 = ~po39  & n9452;
  assign n9455 = ~n9035 & ~n9036;
  assign n9456 = po19  & n9455;
  assign n9457 = ~n9041 & ~n9456;
  assign n9458 = n9041 & n9456;
  assign n9459 = ~n9457 & ~n9458;
  assign n9460 = ~n9454 & ~n9459;
  assign n9461 = ~n9453 & ~n9460;
  assign n9462 = po40  & ~n9461;
  assign n9463 = ~po40  & n9461;
  assign n9464 = ~n9044 & ~n9045;
  assign n9465 = po19  & n9464;
  assign n9466 = ~n9050 & ~n9465;
  assign n9467 = n9050 & n9465;
  assign n9468 = ~n9466 & ~n9467;
  assign n9469 = ~n9463 & ~n9468;
  assign n9470 = ~n9462 & ~n9469;
  assign n9471 = po41  & ~n9470;
  assign n9472 = ~po41  & n9470;
  assign n9473 = ~n9053 & ~n9054;
  assign n9474 = po19  & n9473;
  assign n9475 = ~n9059 & ~n9474;
  assign n9476 = n9059 & n9474;
  assign n9477 = ~n9475 & ~n9476;
  assign n9478 = ~n9472 & ~n9477;
  assign n9479 = ~n9471 & ~n9478;
  assign n9480 = po42  & ~n9479;
  assign n9481 = ~po42  & n9479;
  assign n9482 = ~n9062 & ~n9063;
  assign n9483 = po19  & n9482;
  assign n9484 = ~n9068 & ~n9483;
  assign n9485 = n9068 & n9483;
  assign n9486 = ~n9484 & ~n9485;
  assign n9487 = ~n9481 & ~n9486;
  assign n9488 = ~n9480 & ~n9487;
  assign n9489 = po43  & ~n9488;
  assign n9490 = ~po43  & n9488;
  assign n9491 = ~n9071 & ~n9072;
  assign n9492 = po19  & n9491;
  assign n9493 = ~n9077 & ~n9492;
  assign n9494 = n9077 & n9492;
  assign n9495 = ~n9493 & ~n9494;
  assign n9496 = ~n9490 & ~n9495;
  assign n9497 = ~n9489 & ~n9496;
  assign n9498 = po44  & ~n9497;
  assign n9499 = ~po44  & n9497;
  assign n9500 = ~n9080 & ~n9081;
  assign n9501 = po19  & n9500;
  assign n9502 = ~n9086 & ~n9501;
  assign n9503 = n9086 & n9501;
  assign n9504 = ~n9502 & ~n9503;
  assign n9505 = ~n9499 & ~n9504;
  assign n9506 = ~n9498 & ~n9505;
  assign n9507 = po45  & ~n9506;
  assign n9508 = ~n9089 & ~n9095;
  assign n9509 = po19  & n9508;
  assign n9510 = ~n9094 & ~n9509;
  assign n9511 = n9094 & n9509;
  assign n9512 = ~n9510 & ~n9511;
  assign n9513 = ~po45  & n9506;
  assign n9514 = ~n9512 & ~n9513;
  assign n9515 = ~n9507 & ~n9514;
  assign n9516 = po46  & ~n9515;
  assign n9517 = ~po46  & n9515;
  assign n9518 = ~n9268 & ~n9517;
  assign n9519 = ~n9516 & ~n9518;
  assign n9520 = po47  & ~n9519;
  assign n9521 = ~po47  & n9519;
  assign n9522 = ~n9102 & ~n9103;
  assign n9523 = po19  & n9522;
  assign n9524 = ~n9108 & ~n9523;
  assign n9525 = n9108 & n9523;
  assign n9526 = ~n9524 & ~n9525;
  assign n9527 = ~n9521 & ~n9526;
  assign n9528 = ~n9520 & ~n9527;
  assign n9529 = po48  & ~n9528;
  assign n9530 = ~po48  & n9528;
  assign n9531 = ~n9111 & ~n9112;
  assign n9532 = po19  & n9531;
  assign n9533 = ~n9117 & ~n9532;
  assign n9534 = n9117 & n9532;
  assign n9535 = ~n9533 & ~n9534;
  assign n9536 = ~n9530 & ~n9535;
  assign n9537 = ~n9529 & ~n9536;
  assign n9538 = po49  & ~n9537;
  assign n9539 = ~po49  & n9537;
  assign n9540 = ~n9120 & ~n9121;
  assign n9541 = po19  & n9540;
  assign n9542 = ~n9126 & ~n9541;
  assign n9543 = n9126 & n9541;
  assign n9544 = ~n9542 & ~n9543;
  assign n9545 = ~n9539 & ~n9544;
  assign n9546 = ~n9538 & ~n9545;
  assign n9547 = po50  & ~n9546;
  assign n9548 = ~po50  & n9546;
  assign n9549 = ~n9129 & ~n9130;
  assign n9550 = po19  & n9549;
  assign n9551 = ~n9135 & ~n9550;
  assign n9552 = n9135 & n9550;
  assign n9553 = ~n9551 & ~n9552;
  assign n9554 = ~n9548 & ~n9553;
  assign n9555 = ~n9547 & ~n9554;
  assign n9556 = po51  & ~n9555;
  assign n9557 = ~po51  & n9555;
  assign n9558 = ~n9138 & ~n9139;
  assign n9559 = po19  & n9558;
  assign n9560 = ~n9144 & ~n9559;
  assign n9561 = n9144 & n9559;
  assign n9562 = ~n9560 & ~n9561;
  assign n9563 = ~n9557 & ~n9562;
  assign n9564 = ~n9556 & ~n9563;
  assign n9565 = po52  & ~n9564;
  assign n9566 = ~po52  & n9564;
  assign n9567 = ~n9147 & ~n9148;
  assign n9568 = po19  & n9567;
  assign n9569 = ~n9153 & ~n9568;
  assign n9570 = n9153 & n9568;
  assign n9571 = ~n9569 & ~n9570;
  assign n9572 = ~n9566 & ~n9571;
  assign n9573 = ~n9565 & ~n9572;
  assign n9574 = po53  & ~n9573;
  assign n9575 = ~po53  & n9573;
  assign n9576 = ~n9156 & ~n9157;
  assign n9577 = po19  & n9576;
  assign n9578 = ~n9162 & ~n9577;
  assign n9579 = n9162 & n9577;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = ~n9575 & ~n9580;
  assign n9582 = ~n9574 & ~n9581;
  assign n9583 = po54  & ~n9582;
  assign n9584 = ~po54  & n9582;
  assign n9585 = ~n9165 & ~n9166;
  assign n9586 = po19  & n9585;
  assign n9587 = ~n9171 & ~n9586;
  assign n9588 = n9171 & n9586;
  assign n9589 = ~n9587 & ~n9588;
  assign n9590 = ~n9584 & ~n9589;
  assign n9591 = ~n9583 & ~n9590;
  assign n9592 = po55  & ~n9591;
  assign n9593 = ~po55  & n9591;
  assign n9594 = ~n9174 & ~n9175;
  assign n9595 = po19  & n9594;
  assign n9596 = ~n9180 & ~n9595;
  assign n9597 = n9180 & n9595;
  assign n9598 = ~n9596 & ~n9597;
  assign n9599 = ~n9593 & ~n9598;
  assign n9600 = ~n9592 & ~n9599;
  assign n9601 = po56  & ~n9600;
  assign n9602 = ~po56  & n9600;
  assign n9603 = ~n9183 & ~n9184;
  assign n9604 = po19  & n9603;
  assign n9605 = ~n9189 & ~n9604;
  assign n9606 = n9189 & n9604;
  assign n9607 = ~n9605 & ~n9606;
  assign n9608 = ~n9602 & ~n9607;
  assign n9609 = ~n9601 & ~n9608;
  assign n9610 = po57  & ~n9609;
  assign n9611 = ~po57  & n9609;
  assign n9612 = ~n9192 & ~n9193;
  assign n9613 = po19  & n9612;
  assign n9614 = ~n9198 & ~n9613;
  assign n9615 = n9198 & n9613;
  assign n9616 = ~n9614 & ~n9615;
  assign n9617 = ~n9611 & ~n9616;
  assign n9618 = ~n9610 & ~n9617;
  assign n9619 = po58  & ~n9618;
  assign n9620 = ~po58  & n9618;
  assign n9621 = ~n9201 & ~n9202;
  assign n9622 = po19  & n9621;
  assign n9623 = ~n9207 & ~n9622;
  assign n9624 = n9207 & n9622;
  assign n9625 = ~n9623 & ~n9624;
  assign n9626 = ~n9620 & ~n9625;
  assign n9627 = ~n9619 & ~n9626;
  assign n9628 = po59  & ~n9627;
  assign n9629 = ~po59  & n9627;
  assign n9630 = ~n9210 & ~n9211;
  assign n9631 = po19  & n9630;
  assign n9632 = ~n9216 & ~n9631;
  assign n9633 = n9216 & n9631;
  assign n9634 = ~n9632 & ~n9633;
  assign n9635 = ~n9629 & ~n9634;
  assign n9636 = ~n9628 & ~n9635;
  assign n9637 = po60  & ~n9636;
  assign n9638 = ~po60  & n9636;
  assign n9639 = ~n9219 & ~n9220;
  assign n9640 = po19  & n9639;
  assign n9641 = ~n9225 & ~n9640;
  assign n9642 = n9225 & n9640;
  assign n9643 = ~n9641 & ~n9642;
  assign n9644 = ~n9638 & ~n9643;
  assign n9645 = ~n9637 & ~n9644;
  assign n9646 = po61  & ~n9645;
  assign n9647 = ~po61  & n9645;
  assign n9648 = ~n9228 & ~n9229;
  assign n9649 = po19  & n9648;
  assign n9650 = ~n9234 & ~n9649;
  assign n9651 = n9234 & n9649;
  assign n9652 = ~n9650 & ~n9651;
  assign n9653 = ~n9647 & ~n9652;
  assign n9654 = ~n9646 & ~n9653;
  assign n9655 = po62  & ~n9654;
  assign n9656 = ~po62  & n9654;
  assign n9657 = ~n9237 & ~n9238;
  assign n9658 = po19  & n9657;
  assign n9659 = ~n9243 & ~n9658;
  assign n9660 = n9243 & n9658;
  assign n9661 = ~n9659 & ~n9660;
  assign n9662 = ~n9656 & ~n9661;
  assign n9663 = ~n9655 & ~n9662;
  assign n9664 = n9278 & n9663;
  assign n9665 = ~n9278 & ~n9663;
  assign n9666 = n9256 & po19 ;
  assign n9667 = ~n9255 & ~n9666;
  assign n9668 = n9665 & n9667;
  assign n9669 = ~po63  & ~n9668;
  assign n9670 = ~n9664 & ~n9669;
  assign n9671 = ~n9273 & n9670;
  assign po18  = n9269 | ~n9671;
  assign n9673 = ~n9516 & ~n9517;
  assign n9674 = po18  & n9673;
  assign n9675 = ~n9268 & ~n9674;
  assign n9676 = n9268 & n9674;
  assign n9677 = ~n9675 & ~n9676;
  assign n9678 = n9278 & ~po18 ;
  assign n9679 = ~n9278 & po18 ;
  assign n9680 = n9663 & ~n9679;
  assign n9681 = po63  & ~n9680;
  assign n9682 = ~n9665 & n9681;
  assign n9683 = ~n9655 & ~n9656;
  assign n9684 = po18  & n9683;
  assign n9685 = ~n9661 & ~n9684;
  assign n9686 = n9661 & n9684;
  assign n9687 = ~n9685 & ~n9686;
  assign n9688 = pi36  & po18 ;
  assign n9689 = ~pi34  & ~pi35 ;
  assign n9690 = ~pi36  & n9689;
  assign n9691 = ~n9688 & ~n9690;
  assign n9692 = po19  & ~n9691;
  assign n9693 = ~po19  & n9691;
  assign n9694 = ~pi36  & po18 ;
  assign n9695 = pi37  & ~n9694;
  assign n9696 = n9280 & po18 ;
  assign n9697 = ~n9695 & ~n9696;
  assign n9698 = ~n9693 & n9697;
  assign n9699 = ~n9692 & ~n9698;
  assign n9700 = po20  & ~n9699;
  assign n9701 = ~po20  & n9699;
  assign n9702 = po19  & n9671;
  assign n9703 = ~n9696 & ~n9702;
  assign n9704 = pi38  & ~n9703;
  assign n9705 = ~pi38  & n9703;
  assign n9706 = ~n9704 & ~n9705;
  assign n9707 = ~n9701 & ~n9706;
  assign n9708 = ~n9700 & ~n9707;
  assign n9709 = po21  & ~n9708;
  assign n9710 = ~po21  & n9708;
  assign n9711 = ~n9283 & ~n9284;
  assign n9712 = po18  & n9711;
  assign n9713 = n9288 & ~n9712;
  assign n9714 = ~n9288 & n9712;
  assign n9715 = ~n9713 & ~n9714;
  assign n9716 = ~n9710 & ~n9715;
  assign n9717 = ~n9709 & ~n9716;
  assign n9718 = po22  & ~n9717;
  assign n9719 = ~po22  & n9717;
  assign n9720 = ~n9291 & ~n9292;
  assign n9721 = po18  & n9720;
  assign n9722 = ~n9297 & ~n9721;
  assign n9723 = n9297 & n9721;
  assign n9724 = ~n9722 & ~n9723;
  assign n9725 = ~n9719 & ~n9724;
  assign n9726 = ~n9718 & ~n9725;
  assign n9727 = po23  & ~n9726;
  assign n9728 = ~po23  & n9726;
  assign n9729 = ~n9300 & ~n9301;
  assign n9730 = po18  & n9729;
  assign n9731 = n9306 & n9730;
  assign n9732 = ~n9306 & ~n9730;
  assign n9733 = ~n9731 & ~n9732;
  assign n9734 = ~n9728 & ~n9733;
  assign n9735 = ~n9727 & ~n9734;
  assign n9736 = po24  & ~n9735;
  assign n9737 = ~po24  & n9735;
  assign n9738 = ~n9309 & ~n9310;
  assign n9739 = po18  & n9738;
  assign n9740 = ~n9315 & ~n9739;
  assign n9741 = n9315 & n9739;
  assign n9742 = ~n9740 & ~n9741;
  assign n9743 = ~n9737 & ~n9742;
  assign n9744 = ~n9736 & ~n9743;
  assign n9745 = po25  & ~n9744;
  assign n9746 = ~po25  & n9744;
  assign n9747 = ~n9318 & ~n9319;
  assign n9748 = po18  & n9747;
  assign n9749 = ~n9324 & ~n9748;
  assign n9750 = n9324 & n9748;
  assign n9751 = ~n9749 & ~n9750;
  assign n9752 = ~n9746 & ~n9751;
  assign n9753 = ~n9745 & ~n9752;
  assign n9754 = po26  & ~n9753;
  assign n9755 = ~po26  & n9753;
  assign n9756 = ~n9327 & ~n9328;
  assign n9757 = po18  & n9756;
  assign n9758 = ~n9333 & ~n9757;
  assign n9759 = n9333 & n9757;
  assign n9760 = ~n9758 & ~n9759;
  assign n9761 = ~n9755 & ~n9760;
  assign n9762 = ~n9754 & ~n9761;
  assign n9763 = po27  & ~n9762;
  assign n9764 = ~po27  & n9762;
  assign n9765 = ~n9336 & ~n9337;
  assign n9766 = po18  & n9765;
  assign n9767 = ~n9342 & ~n9766;
  assign n9768 = n9342 & n9766;
  assign n9769 = ~n9767 & ~n9768;
  assign n9770 = ~n9764 & ~n9769;
  assign n9771 = ~n9763 & ~n9770;
  assign n9772 = po28  & ~n9771;
  assign n9773 = ~po28  & n9771;
  assign n9774 = ~n9345 & ~n9346;
  assign n9775 = po18  & n9774;
  assign n9776 = ~n9351 & ~n9775;
  assign n9777 = n9351 & n9775;
  assign n9778 = ~n9776 & ~n9777;
  assign n9779 = ~n9773 & ~n9778;
  assign n9780 = ~n9772 & ~n9779;
  assign n9781 = po29  & ~n9780;
  assign n9782 = ~po29  & n9780;
  assign n9783 = ~n9354 & ~n9355;
  assign n9784 = po18  & n9783;
  assign n9785 = ~n9360 & ~n9784;
  assign n9786 = n9360 & n9784;
  assign n9787 = ~n9785 & ~n9786;
  assign n9788 = ~n9782 & ~n9787;
  assign n9789 = ~n9781 & ~n9788;
  assign n9790 = po30  & ~n9789;
  assign n9791 = ~po30  & n9789;
  assign n9792 = ~n9363 & ~n9364;
  assign n9793 = po18  & n9792;
  assign n9794 = ~n9369 & ~n9793;
  assign n9795 = n9369 & n9793;
  assign n9796 = ~n9794 & ~n9795;
  assign n9797 = ~n9791 & ~n9796;
  assign n9798 = ~n9790 & ~n9797;
  assign n9799 = po31  & ~n9798;
  assign n9800 = ~po31  & n9798;
  assign n9801 = ~n9372 & ~n9373;
  assign n9802 = po18  & n9801;
  assign n9803 = ~n9378 & ~n9802;
  assign n9804 = n9378 & n9802;
  assign n9805 = ~n9803 & ~n9804;
  assign n9806 = ~n9800 & ~n9805;
  assign n9807 = ~n9799 & ~n9806;
  assign n9808 = po32  & ~n9807;
  assign n9809 = ~po32  & n9807;
  assign n9810 = ~n9381 & ~n9382;
  assign n9811 = po18  & n9810;
  assign n9812 = ~n9387 & ~n9811;
  assign n9813 = n9387 & n9811;
  assign n9814 = ~n9812 & ~n9813;
  assign n9815 = ~n9809 & ~n9814;
  assign n9816 = ~n9808 & ~n9815;
  assign n9817 = po33  & ~n9816;
  assign n9818 = ~po33  & n9816;
  assign n9819 = ~n9390 & ~n9391;
  assign n9820 = po18  & n9819;
  assign n9821 = ~n9396 & ~n9820;
  assign n9822 = n9396 & n9820;
  assign n9823 = ~n9821 & ~n9822;
  assign n9824 = ~n9818 & ~n9823;
  assign n9825 = ~n9817 & ~n9824;
  assign n9826 = po34  & ~n9825;
  assign n9827 = ~po34  & n9825;
  assign n9828 = ~n9399 & ~n9400;
  assign n9829 = po18  & n9828;
  assign n9830 = ~n9405 & ~n9829;
  assign n9831 = n9405 & n9829;
  assign n9832 = ~n9830 & ~n9831;
  assign n9833 = ~n9827 & ~n9832;
  assign n9834 = ~n9826 & ~n9833;
  assign n9835 = po35  & ~n9834;
  assign n9836 = ~po35  & n9834;
  assign n9837 = ~n9408 & ~n9409;
  assign n9838 = po18  & n9837;
  assign n9839 = ~n9414 & ~n9838;
  assign n9840 = n9414 & n9838;
  assign n9841 = ~n9839 & ~n9840;
  assign n9842 = ~n9836 & ~n9841;
  assign n9843 = ~n9835 & ~n9842;
  assign n9844 = po36  & ~n9843;
  assign n9845 = ~po36  & n9843;
  assign n9846 = ~n9417 & ~n9418;
  assign n9847 = po18  & n9846;
  assign n9848 = ~n9423 & ~n9847;
  assign n9849 = n9423 & n9847;
  assign n9850 = ~n9848 & ~n9849;
  assign n9851 = ~n9845 & ~n9850;
  assign n9852 = ~n9844 & ~n9851;
  assign n9853 = po37  & ~n9852;
  assign n9854 = ~po37  & n9852;
  assign n9855 = ~n9426 & ~n9427;
  assign n9856 = po18  & n9855;
  assign n9857 = ~n9432 & ~n9856;
  assign n9858 = n9432 & n9856;
  assign n9859 = ~n9857 & ~n9858;
  assign n9860 = ~n9854 & ~n9859;
  assign n9861 = ~n9853 & ~n9860;
  assign n9862 = po38  & ~n9861;
  assign n9863 = ~po38  & n9861;
  assign n9864 = ~n9435 & ~n9436;
  assign n9865 = po18  & n9864;
  assign n9866 = ~n9441 & ~n9865;
  assign n9867 = n9441 & n9865;
  assign n9868 = ~n9866 & ~n9867;
  assign n9869 = ~n9863 & ~n9868;
  assign n9870 = ~n9862 & ~n9869;
  assign n9871 = po39  & ~n9870;
  assign n9872 = ~po39  & n9870;
  assign n9873 = ~n9444 & ~n9445;
  assign n9874 = po18  & n9873;
  assign n9875 = ~n9450 & ~n9874;
  assign n9876 = n9450 & n9874;
  assign n9877 = ~n9875 & ~n9876;
  assign n9878 = ~n9872 & ~n9877;
  assign n9879 = ~n9871 & ~n9878;
  assign n9880 = po40  & ~n9879;
  assign n9881 = ~po40  & n9879;
  assign n9882 = ~n9453 & ~n9454;
  assign n9883 = po18  & n9882;
  assign n9884 = ~n9459 & ~n9883;
  assign n9885 = n9459 & n9883;
  assign n9886 = ~n9884 & ~n9885;
  assign n9887 = ~n9881 & ~n9886;
  assign n9888 = ~n9880 & ~n9887;
  assign n9889 = po41  & ~n9888;
  assign n9890 = ~po41  & n9888;
  assign n9891 = ~n9462 & ~n9463;
  assign n9892 = po18  & n9891;
  assign n9893 = ~n9468 & ~n9892;
  assign n9894 = n9468 & n9892;
  assign n9895 = ~n9893 & ~n9894;
  assign n9896 = ~n9890 & ~n9895;
  assign n9897 = ~n9889 & ~n9896;
  assign n9898 = po42  & ~n9897;
  assign n9899 = ~po42  & n9897;
  assign n9900 = ~n9471 & ~n9472;
  assign n9901 = po18  & n9900;
  assign n9902 = ~n9477 & ~n9901;
  assign n9903 = n9477 & n9901;
  assign n9904 = ~n9902 & ~n9903;
  assign n9905 = ~n9899 & ~n9904;
  assign n9906 = ~n9898 & ~n9905;
  assign n9907 = po43  & ~n9906;
  assign n9908 = ~po43  & n9906;
  assign n9909 = ~n9480 & ~n9481;
  assign n9910 = po18  & n9909;
  assign n9911 = ~n9486 & ~n9910;
  assign n9912 = n9486 & n9910;
  assign n9913 = ~n9911 & ~n9912;
  assign n9914 = ~n9908 & ~n9913;
  assign n9915 = ~n9907 & ~n9914;
  assign n9916 = po44  & ~n9915;
  assign n9917 = ~po44  & n9915;
  assign n9918 = ~n9489 & ~n9490;
  assign n9919 = po18  & n9918;
  assign n9920 = ~n9495 & ~n9919;
  assign n9921 = n9495 & n9919;
  assign n9922 = ~n9920 & ~n9921;
  assign n9923 = ~n9917 & ~n9922;
  assign n9924 = ~n9916 & ~n9923;
  assign n9925 = po45  & ~n9924;
  assign n9926 = ~po45  & n9924;
  assign n9927 = ~n9498 & ~n9499;
  assign n9928 = po18  & n9927;
  assign n9929 = ~n9504 & ~n9928;
  assign n9930 = n9504 & n9928;
  assign n9931 = ~n9929 & ~n9930;
  assign n9932 = ~n9926 & ~n9931;
  assign n9933 = ~n9925 & ~n9932;
  assign n9934 = po46  & ~n9933;
  assign n9935 = ~n9507 & ~n9513;
  assign n9936 = po18  & n9935;
  assign n9937 = ~n9512 & ~n9936;
  assign n9938 = n9512 & n9936;
  assign n9939 = ~n9937 & ~n9938;
  assign n9940 = ~po46  & n9933;
  assign n9941 = ~n9939 & ~n9940;
  assign n9942 = ~n9934 & ~n9941;
  assign n9943 = po47  & ~n9942;
  assign n9944 = ~po47  & n9942;
  assign n9945 = ~n9677 & ~n9944;
  assign n9946 = ~n9943 & ~n9945;
  assign n9947 = po48  & ~n9946;
  assign n9948 = ~po48  & n9946;
  assign n9949 = ~n9520 & ~n9521;
  assign n9950 = po18  & n9949;
  assign n9951 = ~n9526 & ~n9950;
  assign n9952 = n9526 & n9950;
  assign n9953 = ~n9951 & ~n9952;
  assign n9954 = ~n9948 & ~n9953;
  assign n9955 = ~n9947 & ~n9954;
  assign n9956 = po49  & ~n9955;
  assign n9957 = ~po49  & n9955;
  assign n9958 = ~n9529 & ~n9530;
  assign n9959 = po18  & n9958;
  assign n9960 = ~n9535 & ~n9959;
  assign n9961 = n9535 & n9959;
  assign n9962 = ~n9960 & ~n9961;
  assign n9963 = ~n9957 & ~n9962;
  assign n9964 = ~n9956 & ~n9963;
  assign n9965 = po50  & ~n9964;
  assign n9966 = ~po50  & n9964;
  assign n9967 = ~n9538 & ~n9539;
  assign n9968 = po18  & n9967;
  assign n9969 = ~n9544 & ~n9968;
  assign n9970 = n9544 & n9968;
  assign n9971 = ~n9969 & ~n9970;
  assign n9972 = ~n9966 & ~n9971;
  assign n9973 = ~n9965 & ~n9972;
  assign n9974 = po51  & ~n9973;
  assign n9975 = ~po51  & n9973;
  assign n9976 = ~n9547 & ~n9548;
  assign n9977 = po18  & n9976;
  assign n9978 = ~n9553 & ~n9977;
  assign n9979 = n9553 & n9977;
  assign n9980 = ~n9978 & ~n9979;
  assign n9981 = ~n9975 & ~n9980;
  assign n9982 = ~n9974 & ~n9981;
  assign n9983 = po52  & ~n9982;
  assign n9984 = ~po52  & n9982;
  assign n9985 = ~n9556 & ~n9557;
  assign n9986 = po18  & n9985;
  assign n9987 = ~n9562 & ~n9986;
  assign n9988 = n9562 & n9986;
  assign n9989 = ~n9987 & ~n9988;
  assign n9990 = ~n9984 & ~n9989;
  assign n9991 = ~n9983 & ~n9990;
  assign n9992 = po53  & ~n9991;
  assign n9993 = ~po53  & n9991;
  assign n9994 = ~n9565 & ~n9566;
  assign n9995 = po18  & n9994;
  assign n9996 = ~n9571 & ~n9995;
  assign n9997 = n9571 & n9995;
  assign n9998 = ~n9996 & ~n9997;
  assign n9999 = ~n9993 & ~n9998;
  assign n10000 = ~n9992 & ~n9999;
  assign n10001 = po54  & ~n10000;
  assign n10002 = ~po54  & n10000;
  assign n10003 = ~n9574 & ~n9575;
  assign n10004 = po18  & n10003;
  assign n10005 = ~n9580 & ~n10004;
  assign n10006 = n9580 & n10004;
  assign n10007 = ~n10005 & ~n10006;
  assign n10008 = ~n10002 & ~n10007;
  assign n10009 = ~n10001 & ~n10008;
  assign n10010 = po55  & ~n10009;
  assign n10011 = ~po55  & n10009;
  assign n10012 = ~n9583 & ~n9584;
  assign n10013 = po18  & n10012;
  assign n10014 = ~n9589 & ~n10013;
  assign n10015 = n9589 & n10013;
  assign n10016 = ~n10014 & ~n10015;
  assign n10017 = ~n10011 & ~n10016;
  assign n10018 = ~n10010 & ~n10017;
  assign n10019 = po56  & ~n10018;
  assign n10020 = ~po56  & n10018;
  assign n10021 = ~n9592 & ~n9593;
  assign n10022 = po18  & n10021;
  assign n10023 = ~n9598 & ~n10022;
  assign n10024 = n9598 & n10022;
  assign n10025 = ~n10023 & ~n10024;
  assign n10026 = ~n10020 & ~n10025;
  assign n10027 = ~n10019 & ~n10026;
  assign n10028 = po57  & ~n10027;
  assign n10029 = ~po57  & n10027;
  assign n10030 = ~n9601 & ~n9602;
  assign n10031 = po18  & n10030;
  assign n10032 = ~n9607 & ~n10031;
  assign n10033 = n9607 & n10031;
  assign n10034 = ~n10032 & ~n10033;
  assign n10035 = ~n10029 & ~n10034;
  assign n10036 = ~n10028 & ~n10035;
  assign n10037 = po58  & ~n10036;
  assign n10038 = ~po58  & n10036;
  assign n10039 = ~n9610 & ~n9611;
  assign n10040 = po18  & n10039;
  assign n10041 = ~n9616 & ~n10040;
  assign n10042 = n9616 & n10040;
  assign n10043 = ~n10041 & ~n10042;
  assign n10044 = ~n10038 & ~n10043;
  assign n10045 = ~n10037 & ~n10044;
  assign n10046 = po59  & ~n10045;
  assign n10047 = ~po59  & n10045;
  assign n10048 = ~n9619 & ~n9620;
  assign n10049 = po18  & n10048;
  assign n10050 = ~n9625 & ~n10049;
  assign n10051 = n9625 & n10049;
  assign n10052 = ~n10050 & ~n10051;
  assign n10053 = ~n10047 & ~n10052;
  assign n10054 = ~n10046 & ~n10053;
  assign n10055 = po60  & ~n10054;
  assign n10056 = ~po60  & n10054;
  assign n10057 = ~n9628 & ~n9629;
  assign n10058 = po18  & n10057;
  assign n10059 = ~n9634 & ~n10058;
  assign n10060 = n9634 & n10058;
  assign n10061 = ~n10059 & ~n10060;
  assign n10062 = ~n10056 & ~n10061;
  assign n10063 = ~n10055 & ~n10062;
  assign n10064 = po61  & ~n10063;
  assign n10065 = ~po61  & n10063;
  assign n10066 = ~n9637 & ~n9638;
  assign n10067 = po18  & n10066;
  assign n10068 = ~n9643 & ~n10067;
  assign n10069 = n9643 & n10067;
  assign n10070 = ~n10068 & ~n10069;
  assign n10071 = ~n10065 & ~n10070;
  assign n10072 = ~n10064 & ~n10071;
  assign n10073 = po62  & ~n10072;
  assign n10074 = ~po62  & n10072;
  assign n10075 = ~n9646 & ~n9647;
  assign n10076 = po18  & n10075;
  assign n10077 = ~n9652 & ~n10076;
  assign n10078 = n9652 & n10076;
  assign n10079 = ~n10077 & ~n10078;
  assign n10080 = ~n10074 & ~n10079;
  assign n10081 = ~n10073 & ~n10080;
  assign n10082 = n9687 & n10081;
  assign n10083 = ~n9687 & ~n10081;
  assign n10084 = n9665 & po18 ;
  assign n10085 = ~n9664 & ~n10084;
  assign n10086 = n10083 & n10085;
  assign n10087 = ~po63  & ~n10086;
  assign n10088 = ~n10082 & ~n10087;
  assign n10089 = ~n9682 & n10088;
  assign po17  = n9678 | ~n10089;
  assign n10091 = ~n9943 & ~n9944;
  assign n10092 = po17  & n10091;
  assign n10093 = ~n9677 & ~n10092;
  assign n10094 = n9677 & n10092;
  assign n10095 = ~n10093 & ~n10094;
  assign n10096 = n9687 & ~po17 ;
  assign n10097 = ~n9687 & po17 ;
  assign n10098 = n10081 & ~n10097;
  assign n10099 = po63  & ~n10098;
  assign n10100 = ~n10083 & n10099;
  assign n10101 = ~n10073 & ~n10074;
  assign n10102 = po17  & n10101;
  assign n10103 = ~n10079 & ~n10102;
  assign n10104 = n10079 & n10102;
  assign n10105 = ~n10103 & ~n10104;
  assign n10106 = pi34  & po17 ;
  assign n10107 = ~pi32  & ~pi33 ;
  assign n10108 = ~pi34  & n10107;
  assign n10109 = ~n10106 & ~n10108;
  assign n10110 = po18  & ~n10109;
  assign n10111 = ~po18  & n10109;
  assign n10112 = ~pi34  & po17 ;
  assign n10113 = pi35  & ~n10112;
  assign n10114 = n9689 & po17 ;
  assign n10115 = ~n10113 & ~n10114;
  assign n10116 = ~n10111 & n10115;
  assign n10117 = ~n10110 & ~n10116;
  assign n10118 = po19  & ~n10117;
  assign n10119 = ~po19  & n10117;
  assign n10120 = po18  & n10089;
  assign n10121 = ~n10114 & ~n10120;
  assign n10122 = pi36  & ~n10121;
  assign n10123 = ~pi36  & n10121;
  assign n10124 = ~n10122 & ~n10123;
  assign n10125 = ~n10119 & ~n10124;
  assign n10126 = ~n10118 & ~n10125;
  assign n10127 = po20  & ~n10126;
  assign n10128 = ~po20  & n10126;
  assign n10129 = ~n9692 & ~n9693;
  assign n10130 = po17  & n10129;
  assign n10131 = n9697 & ~n10130;
  assign n10132 = ~n9697 & n10130;
  assign n10133 = ~n10131 & ~n10132;
  assign n10134 = ~n10128 & ~n10133;
  assign n10135 = ~n10127 & ~n10134;
  assign n10136 = po21  & ~n10135;
  assign n10137 = ~po21  & n10135;
  assign n10138 = ~n9700 & ~n9701;
  assign n10139 = po17  & n10138;
  assign n10140 = ~n9706 & ~n10139;
  assign n10141 = n9706 & n10139;
  assign n10142 = ~n10140 & ~n10141;
  assign n10143 = ~n10137 & ~n10142;
  assign n10144 = ~n10136 & ~n10143;
  assign n10145 = po22  & ~n10144;
  assign n10146 = ~po22  & n10144;
  assign n10147 = ~n9709 & ~n9710;
  assign n10148 = po17  & n10147;
  assign n10149 = n9715 & n10148;
  assign n10150 = ~n9715 & ~n10148;
  assign n10151 = ~n10149 & ~n10150;
  assign n10152 = ~n10146 & ~n10151;
  assign n10153 = ~n10145 & ~n10152;
  assign n10154 = po23  & ~n10153;
  assign n10155 = ~po23  & n10153;
  assign n10156 = ~n9718 & ~n9719;
  assign n10157 = po17  & n10156;
  assign n10158 = ~n9724 & ~n10157;
  assign n10159 = n9724 & n10157;
  assign n10160 = ~n10158 & ~n10159;
  assign n10161 = ~n10155 & ~n10160;
  assign n10162 = ~n10154 & ~n10161;
  assign n10163 = po24  & ~n10162;
  assign n10164 = ~po24  & n10162;
  assign n10165 = ~n9727 & ~n9728;
  assign n10166 = po17  & n10165;
  assign n10167 = ~n9733 & ~n10166;
  assign n10168 = n9733 & n10166;
  assign n10169 = ~n10167 & ~n10168;
  assign n10170 = ~n10164 & ~n10169;
  assign n10171 = ~n10163 & ~n10170;
  assign n10172 = po25  & ~n10171;
  assign n10173 = ~po25  & n10171;
  assign n10174 = ~n9736 & ~n9737;
  assign n10175 = po17  & n10174;
  assign n10176 = ~n9742 & ~n10175;
  assign n10177 = n9742 & n10175;
  assign n10178 = ~n10176 & ~n10177;
  assign n10179 = ~n10173 & ~n10178;
  assign n10180 = ~n10172 & ~n10179;
  assign n10181 = po26  & ~n10180;
  assign n10182 = ~po26  & n10180;
  assign n10183 = ~n9745 & ~n9746;
  assign n10184 = po17  & n10183;
  assign n10185 = ~n9751 & ~n10184;
  assign n10186 = n9751 & n10184;
  assign n10187 = ~n10185 & ~n10186;
  assign n10188 = ~n10182 & ~n10187;
  assign n10189 = ~n10181 & ~n10188;
  assign n10190 = po27  & ~n10189;
  assign n10191 = ~po27  & n10189;
  assign n10192 = ~n9754 & ~n9755;
  assign n10193 = po17  & n10192;
  assign n10194 = ~n9760 & ~n10193;
  assign n10195 = n9760 & n10193;
  assign n10196 = ~n10194 & ~n10195;
  assign n10197 = ~n10191 & ~n10196;
  assign n10198 = ~n10190 & ~n10197;
  assign n10199 = po28  & ~n10198;
  assign n10200 = ~po28  & n10198;
  assign n10201 = ~n9763 & ~n9764;
  assign n10202 = po17  & n10201;
  assign n10203 = ~n9769 & ~n10202;
  assign n10204 = n9769 & n10202;
  assign n10205 = ~n10203 & ~n10204;
  assign n10206 = ~n10200 & ~n10205;
  assign n10207 = ~n10199 & ~n10206;
  assign n10208 = po29  & ~n10207;
  assign n10209 = ~po29  & n10207;
  assign n10210 = ~n9772 & ~n9773;
  assign n10211 = po17  & n10210;
  assign n10212 = ~n9778 & ~n10211;
  assign n10213 = n9778 & n10211;
  assign n10214 = ~n10212 & ~n10213;
  assign n10215 = ~n10209 & ~n10214;
  assign n10216 = ~n10208 & ~n10215;
  assign n10217 = po30  & ~n10216;
  assign n10218 = ~po30  & n10216;
  assign n10219 = ~n9781 & ~n9782;
  assign n10220 = po17  & n10219;
  assign n10221 = ~n9787 & ~n10220;
  assign n10222 = n9787 & n10220;
  assign n10223 = ~n10221 & ~n10222;
  assign n10224 = ~n10218 & ~n10223;
  assign n10225 = ~n10217 & ~n10224;
  assign n10226 = po31  & ~n10225;
  assign n10227 = ~po31  & n10225;
  assign n10228 = ~n9790 & ~n9791;
  assign n10229 = po17  & n10228;
  assign n10230 = ~n9796 & ~n10229;
  assign n10231 = n9796 & n10229;
  assign n10232 = ~n10230 & ~n10231;
  assign n10233 = ~n10227 & ~n10232;
  assign n10234 = ~n10226 & ~n10233;
  assign n10235 = po32  & ~n10234;
  assign n10236 = ~po32  & n10234;
  assign n10237 = ~n9799 & ~n9800;
  assign n10238 = po17  & n10237;
  assign n10239 = ~n9805 & ~n10238;
  assign n10240 = n9805 & n10238;
  assign n10241 = ~n10239 & ~n10240;
  assign n10242 = ~n10236 & ~n10241;
  assign n10243 = ~n10235 & ~n10242;
  assign n10244 = po33  & ~n10243;
  assign n10245 = ~po33  & n10243;
  assign n10246 = ~n9808 & ~n9809;
  assign n10247 = po17  & n10246;
  assign n10248 = ~n9814 & ~n10247;
  assign n10249 = n9814 & n10247;
  assign n10250 = ~n10248 & ~n10249;
  assign n10251 = ~n10245 & ~n10250;
  assign n10252 = ~n10244 & ~n10251;
  assign n10253 = po34  & ~n10252;
  assign n10254 = ~po34  & n10252;
  assign n10255 = ~n9817 & ~n9818;
  assign n10256 = po17  & n10255;
  assign n10257 = ~n9823 & ~n10256;
  assign n10258 = n9823 & n10256;
  assign n10259 = ~n10257 & ~n10258;
  assign n10260 = ~n10254 & ~n10259;
  assign n10261 = ~n10253 & ~n10260;
  assign n10262 = po35  & ~n10261;
  assign n10263 = ~po35  & n10261;
  assign n10264 = ~n9826 & ~n9827;
  assign n10265 = po17  & n10264;
  assign n10266 = ~n9832 & ~n10265;
  assign n10267 = n9832 & n10265;
  assign n10268 = ~n10266 & ~n10267;
  assign n10269 = ~n10263 & ~n10268;
  assign n10270 = ~n10262 & ~n10269;
  assign n10271 = po36  & ~n10270;
  assign n10272 = ~po36  & n10270;
  assign n10273 = ~n9835 & ~n9836;
  assign n10274 = po17  & n10273;
  assign n10275 = ~n9841 & ~n10274;
  assign n10276 = n9841 & n10274;
  assign n10277 = ~n10275 & ~n10276;
  assign n10278 = ~n10272 & ~n10277;
  assign n10279 = ~n10271 & ~n10278;
  assign n10280 = po37  & ~n10279;
  assign n10281 = ~po37  & n10279;
  assign n10282 = ~n9844 & ~n9845;
  assign n10283 = po17  & n10282;
  assign n10284 = ~n9850 & ~n10283;
  assign n10285 = n9850 & n10283;
  assign n10286 = ~n10284 & ~n10285;
  assign n10287 = ~n10281 & ~n10286;
  assign n10288 = ~n10280 & ~n10287;
  assign n10289 = po38  & ~n10288;
  assign n10290 = ~po38  & n10288;
  assign n10291 = ~n9853 & ~n9854;
  assign n10292 = po17  & n10291;
  assign n10293 = ~n9859 & ~n10292;
  assign n10294 = n9859 & n10292;
  assign n10295 = ~n10293 & ~n10294;
  assign n10296 = ~n10290 & ~n10295;
  assign n10297 = ~n10289 & ~n10296;
  assign n10298 = po39  & ~n10297;
  assign n10299 = ~po39  & n10297;
  assign n10300 = ~n9862 & ~n9863;
  assign n10301 = po17  & n10300;
  assign n10302 = ~n9868 & ~n10301;
  assign n10303 = n9868 & n10301;
  assign n10304 = ~n10302 & ~n10303;
  assign n10305 = ~n10299 & ~n10304;
  assign n10306 = ~n10298 & ~n10305;
  assign n10307 = po40  & ~n10306;
  assign n10308 = ~po40  & n10306;
  assign n10309 = ~n9871 & ~n9872;
  assign n10310 = po17  & n10309;
  assign n10311 = ~n9877 & ~n10310;
  assign n10312 = n9877 & n10310;
  assign n10313 = ~n10311 & ~n10312;
  assign n10314 = ~n10308 & ~n10313;
  assign n10315 = ~n10307 & ~n10314;
  assign n10316 = po41  & ~n10315;
  assign n10317 = ~po41  & n10315;
  assign n10318 = ~n9880 & ~n9881;
  assign n10319 = po17  & n10318;
  assign n10320 = ~n9886 & ~n10319;
  assign n10321 = n9886 & n10319;
  assign n10322 = ~n10320 & ~n10321;
  assign n10323 = ~n10317 & ~n10322;
  assign n10324 = ~n10316 & ~n10323;
  assign n10325 = po42  & ~n10324;
  assign n10326 = ~po42  & n10324;
  assign n10327 = ~n9889 & ~n9890;
  assign n10328 = po17  & n10327;
  assign n10329 = ~n9895 & ~n10328;
  assign n10330 = n9895 & n10328;
  assign n10331 = ~n10329 & ~n10330;
  assign n10332 = ~n10326 & ~n10331;
  assign n10333 = ~n10325 & ~n10332;
  assign n10334 = po43  & ~n10333;
  assign n10335 = ~po43  & n10333;
  assign n10336 = ~n9898 & ~n9899;
  assign n10337 = po17  & n10336;
  assign n10338 = ~n9904 & ~n10337;
  assign n10339 = n9904 & n10337;
  assign n10340 = ~n10338 & ~n10339;
  assign n10341 = ~n10335 & ~n10340;
  assign n10342 = ~n10334 & ~n10341;
  assign n10343 = po44  & ~n10342;
  assign n10344 = ~po44  & n10342;
  assign n10345 = ~n9907 & ~n9908;
  assign n10346 = po17  & n10345;
  assign n10347 = ~n9913 & ~n10346;
  assign n10348 = n9913 & n10346;
  assign n10349 = ~n10347 & ~n10348;
  assign n10350 = ~n10344 & ~n10349;
  assign n10351 = ~n10343 & ~n10350;
  assign n10352 = po45  & ~n10351;
  assign n10353 = ~po45  & n10351;
  assign n10354 = ~n9916 & ~n9917;
  assign n10355 = po17  & n10354;
  assign n10356 = ~n9922 & ~n10355;
  assign n10357 = n9922 & n10355;
  assign n10358 = ~n10356 & ~n10357;
  assign n10359 = ~n10353 & ~n10358;
  assign n10360 = ~n10352 & ~n10359;
  assign n10361 = po46  & ~n10360;
  assign n10362 = ~po46  & n10360;
  assign n10363 = ~n9925 & ~n9926;
  assign n10364 = po17  & n10363;
  assign n10365 = ~n9931 & ~n10364;
  assign n10366 = n9931 & n10364;
  assign n10367 = ~n10365 & ~n10366;
  assign n10368 = ~n10362 & ~n10367;
  assign n10369 = ~n10361 & ~n10368;
  assign n10370 = po47  & ~n10369;
  assign n10371 = ~n9934 & ~n9940;
  assign n10372 = po17  & n10371;
  assign n10373 = ~n9939 & ~n10372;
  assign n10374 = n9939 & n10372;
  assign n10375 = ~n10373 & ~n10374;
  assign n10376 = ~po47  & n10369;
  assign n10377 = ~n10375 & ~n10376;
  assign n10378 = ~n10370 & ~n10377;
  assign n10379 = po48  & ~n10378;
  assign n10380 = ~po48  & n10378;
  assign n10381 = ~n10095 & ~n10380;
  assign n10382 = ~n10379 & ~n10381;
  assign n10383 = po49  & ~n10382;
  assign n10384 = ~po49  & n10382;
  assign n10385 = ~n9947 & ~n9948;
  assign n10386 = po17  & n10385;
  assign n10387 = ~n9953 & ~n10386;
  assign n10388 = n9953 & n10386;
  assign n10389 = ~n10387 & ~n10388;
  assign n10390 = ~n10384 & ~n10389;
  assign n10391 = ~n10383 & ~n10390;
  assign n10392 = po50  & ~n10391;
  assign n10393 = ~po50  & n10391;
  assign n10394 = ~n9956 & ~n9957;
  assign n10395 = po17  & n10394;
  assign n10396 = ~n9962 & ~n10395;
  assign n10397 = n9962 & n10395;
  assign n10398 = ~n10396 & ~n10397;
  assign n10399 = ~n10393 & ~n10398;
  assign n10400 = ~n10392 & ~n10399;
  assign n10401 = po51  & ~n10400;
  assign n10402 = ~po51  & n10400;
  assign n10403 = ~n9965 & ~n9966;
  assign n10404 = po17  & n10403;
  assign n10405 = ~n9971 & ~n10404;
  assign n10406 = n9971 & n10404;
  assign n10407 = ~n10405 & ~n10406;
  assign n10408 = ~n10402 & ~n10407;
  assign n10409 = ~n10401 & ~n10408;
  assign n10410 = po52  & ~n10409;
  assign n10411 = ~po52  & n10409;
  assign n10412 = ~n9974 & ~n9975;
  assign n10413 = po17  & n10412;
  assign n10414 = ~n9980 & ~n10413;
  assign n10415 = n9980 & n10413;
  assign n10416 = ~n10414 & ~n10415;
  assign n10417 = ~n10411 & ~n10416;
  assign n10418 = ~n10410 & ~n10417;
  assign n10419 = po53  & ~n10418;
  assign n10420 = ~po53  & n10418;
  assign n10421 = ~n9983 & ~n9984;
  assign n10422 = po17  & n10421;
  assign n10423 = ~n9989 & ~n10422;
  assign n10424 = n9989 & n10422;
  assign n10425 = ~n10423 & ~n10424;
  assign n10426 = ~n10420 & ~n10425;
  assign n10427 = ~n10419 & ~n10426;
  assign n10428 = po54  & ~n10427;
  assign n10429 = ~po54  & n10427;
  assign n10430 = ~n9992 & ~n9993;
  assign n10431 = po17  & n10430;
  assign n10432 = ~n9998 & ~n10431;
  assign n10433 = n9998 & n10431;
  assign n10434 = ~n10432 & ~n10433;
  assign n10435 = ~n10429 & ~n10434;
  assign n10436 = ~n10428 & ~n10435;
  assign n10437 = po55  & ~n10436;
  assign n10438 = ~po55  & n10436;
  assign n10439 = ~n10001 & ~n10002;
  assign n10440 = po17  & n10439;
  assign n10441 = ~n10007 & ~n10440;
  assign n10442 = n10007 & n10440;
  assign n10443 = ~n10441 & ~n10442;
  assign n10444 = ~n10438 & ~n10443;
  assign n10445 = ~n10437 & ~n10444;
  assign n10446 = po56  & ~n10445;
  assign n10447 = ~po56  & n10445;
  assign n10448 = ~n10010 & ~n10011;
  assign n10449 = po17  & n10448;
  assign n10450 = ~n10016 & ~n10449;
  assign n10451 = n10016 & n10449;
  assign n10452 = ~n10450 & ~n10451;
  assign n10453 = ~n10447 & ~n10452;
  assign n10454 = ~n10446 & ~n10453;
  assign n10455 = po57  & ~n10454;
  assign n10456 = ~po57  & n10454;
  assign n10457 = ~n10019 & ~n10020;
  assign n10458 = po17  & n10457;
  assign n10459 = ~n10025 & ~n10458;
  assign n10460 = n10025 & n10458;
  assign n10461 = ~n10459 & ~n10460;
  assign n10462 = ~n10456 & ~n10461;
  assign n10463 = ~n10455 & ~n10462;
  assign n10464 = po58  & ~n10463;
  assign n10465 = ~po58  & n10463;
  assign n10466 = ~n10028 & ~n10029;
  assign n10467 = po17  & n10466;
  assign n10468 = ~n10034 & ~n10467;
  assign n10469 = n10034 & n10467;
  assign n10470 = ~n10468 & ~n10469;
  assign n10471 = ~n10465 & ~n10470;
  assign n10472 = ~n10464 & ~n10471;
  assign n10473 = po59  & ~n10472;
  assign n10474 = ~po59  & n10472;
  assign n10475 = ~n10037 & ~n10038;
  assign n10476 = po17  & n10475;
  assign n10477 = ~n10043 & ~n10476;
  assign n10478 = n10043 & n10476;
  assign n10479 = ~n10477 & ~n10478;
  assign n10480 = ~n10474 & ~n10479;
  assign n10481 = ~n10473 & ~n10480;
  assign n10482 = po60  & ~n10481;
  assign n10483 = ~po60  & n10481;
  assign n10484 = ~n10046 & ~n10047;
  assign n10485 = po17  & n10484;
  assign n10486 = ~n10052 & ~n10485;
  assign n10487 = n10052 & n10485;
  assign n10488 = ~n10486 & ~n10487;
  assign n10489 = ~n10483 & ~n10488;
  assign n10490 = ~n10482 & ~n10489;
  assign n10491 = po61  & ~n10490;
  assign n10492 = ~po61  & n10490;
  assign n10493 = ~n10055 & ~n10056;
  assign n10494 = po17  & n10493;
  assign n10495 = ~n10061 & ~n10494;
  assign n10496 = n10061 & n10494;
  assign n10497 = ~n10495 & ~n10496;
  assign n10498 = ~n10492 & ~n10497;
  assign n10499 = ~n10491 & ~n10498;
  assign n10500 = po62  & ~n10499;
  assign n10501 = ~po62  & n10499;
  assign n10502 = ~n10064 & ~n10065;
  assign n10503 = po17  & n10502;
  assign n10504 = ~n10070 & ~n10503;
  assign n10505 = n10070 & n10503;
  assign n10506 = ~n10504 & ~n10505;
  assign n10507 = ~n10501 & ~n10506;
  assign n10508 = ~n10500 & ~n10507;
  assign n10509 = n10105 & n10508;
  assign n10510 = ~n10105 & ~n10508;
  assign n10511 = n10083 & po17 ;
  assign n10512 = ~n10082 & ~n10511;
  assign n10513 = n10510 & n10512;
  assign n10514 = ~po63  & ~n10513;
  assign n10515 = ~n10509 & ~n10514;
  assign n10516 = ~n10100 & n10515;
  assign po16  = n10096 | ~n10516;
  assign n10518 = ~n10379 & ~n10380;
  assign n10519 = po16  & n10518;
  assign n10520 = ~n10095 & ~n10519;
  assign n10521 = n10095 & n10519;
  assign n10522 = ~n10520 & ~n10521;
  assign n10523 = n10105 & ~po16 ;
  assign n10524 = ~n10105 & po16 ;
  assign n10525 = n10508 & ~n10524;
  assign n10526 = po63  & ~n10525;
  assign n10527 = ~n10510 & n10526;
  assign n10528 = ~n10500 & ~n10501;
  assign n10529 = po16  & n10528;
  assign n10530 = ~n10506 & ~n10529;
  assign n10531 = n10506 & n10529;
  assign n10532 = ~n10530 & ~n10531;
  assign n10533 = pi32  & po16 ;
  assign n10534 = ~pi30  & ~pi31 ;
  assign n10535 = ~pi32  & n10534;
  assign n10536 = ~n10533 & ~n10535;
  assign n10537 = po17  & ~n10536;
  assign n10538 = ~po17  & n10536;
  assign n10539 = ~pi32  & po16 ;
  assign n10540 = pi33  & ~n10539;
  assign n10541 = n10107 & po16 ;
  assign n10542 = ~n10540 & ~n10541;
  assign n10543 = ~n10538 & n10542;
  assign n10544 = ~n10537 & ~n10543;
  assign n10545 = po18  & ~n10544;
  assign n10546 = ~po18  & n10544;
  assign n10547 = po17  & n10516;
  assign n10548 = ~n10541 & ~n10547;
  assign n10549 = pi34  & ~n10548;
  assign n10550 = ~pi34  & n10548;
  assign n10551 = ~n10549 & ~n10550;
  assign n10552 = ~n10546 & ~n10551;
  assign n10553 = ~n10545 & ~n10552;
  assign n10554 = po19  & ~n10553;
  assign n10555 = ~po19  & n10553;
  assign n10556 = ~n10110 & ~n10111;
  assign n10557 = po16  & n10556;
  assign n10558 = n10115 & ~n10557;
  assign n10559 = ~n10115 & n10557;
  assign n10560 = ~n10558 & ~n10559;
  assign n10561 = ~n10555 & ~n10560;
  assign n10562 = ~n10554 & ~n10561;
  assign n10563 = po20  & ~n10562;
  assign n10564 = ~po20  & n10562;
  assign n10565 = ~n10118 & ~n10119;
  assign n10566 = po16  & n10565;
  assign n10567 = ~n10124 & ~n10566;
  assign n10568 = n10124 & n10566;
  assign n10569 = ~n10567 & ~n10568;
  assign n10570 = ~n10564 & ~n10569;
  assign n10571 = ~n10563 & ~n10570;
  assign n10572 = po21  & ~n10571;
  assign n10573 = ~po21  & n10571;
  assign n10574 = ~n10127 & ~n10128;
  assign n10575 = po16  & n10574;
  assign n10576 = n10133 & n10575;
  assign n10577 = ~n10133 & ~n10575;
  assign n10578 = ~n10576 & ~n10577;
  assign n10579 = ~n10573 & ~n10578;
  assign n10580 = ~n10572 & ~n10579;
  assign n10581 = po22  & ~n10580;
  assign n10582 = ~po22  & n10580;
  assign n10583 = ~n10136 & ~n10137;
  assign n10584 = po16  & n10583;
  assign n10585 = ~n10142 & ~n10584;
  assign n10586 = n10142 & n10584;
  assign n10587 = ~n10585 & ~n10586;
  assign n10588 = ~n10582 & ~n10587;
  assign n10589 = ~n10581 & ~n10588;
  assign n10590 = po23  & ~n10589;
  assign n10591 = ~po23  & n10589;
  assign n10592 = ~n10145 & ~n10146;
  assign n10593 = po16  & n10592;
  assign n10594 = ~n10151 & ~n10593;
  assign n10595 = n10151 & n10593;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = ~n10591 & ~n10596;
  assign n10598 = ~n10590 & ~n10597;
  assign n10599 = po24  & ~n10598;
  assign n10600 = ~po24  & n10598;
  assign n10601 = ~n10154 & ~n10155;
  assign n10602 = po16  & n10601;
  assign n10603 = ~n10160 & ~n10602;
  assign n10604 = n10160 & n10602;
  assign n10605 = ~n10603 & ~n10604;
  assign n10606 = ~n10600 & ~n10605;
  assign n10607 = ~n10599 & ~n10606;
  assign n10608 = po25  & ~n10607;
  assign n10609 = ~po25  & n10607;
  assign n10610 = ~n10163 & ~n10164;
  assign n10611 = po16  & n10610;
  assign n10612 = ~n10169 & ~n10611;
  assign n10613 = n10169 & n10611;
  assign n10614 = ~n10612 & ~n10613;
  assign n10615 = ~n10609 & ~n10614;
  assign n10616 = ~n10608 & ~n10615;
  assign n10617 = po26  & ~n10616;
  assign n10618 = ~po26  & n10616;
  assign n10619 = ~n10172 & ~n10173;
  assign n10620 = po16  & n10619;
  assign n10621 = ~n10178 & ~n10620;
  assign n10622 = n10178 & n10620;
  assign n10623 = ~n10621 & ~n10622;
  assign n10624 = ~n10618 & ~n10623;
  assign n10625 = ~n10617 & ~n10624;
  assign n10626 = po27  & ~n10625;
  assign n10627 = ~po27  & n10625;
  assign n10628 = ~n10181 & ~n10182;
  assign n10629 = po16  & n10628;
  assign n10630 = ~n10187 & ~n10629;
  assign n10631 = n10187 & n10629;
  assign n10632 = ~n10630 & ~n10631;
  assign n10633 = ~n10627 & ~n10632;
  assign n10634 = ~n10626 & ~n10633;
  assign n10635 = po28  & ~n10634;
  assign n10636 = ~po28  & n10634;
  assign n10637 = ~n10190 & ~n10191;
  assign n10638 = po16  & n10637;
  assign n10639 = ~n10196 & ~n10638;
  assign n10640 = n10196 & n10638;
  assign n10641 = ~n10639 & ~n10640;
  assign n10642 = ~n10636 & ~n10641;
  assign n10643 = ~n10635 & ~n10642;
  assign n10644 = po29  & ~n10643;
  assign n10645 = ~po29  & n10643;
  assign n10646 = ~n10199 & ~n10200;
  assign n10647 = po16  & n10646;
  assign n10648 = ~n10205 & ~n10647;
  assign n10649 = n10205 & n10647;
  assign n10650 = ~n10648 & ~n10649;
  assign n10651 = ~n10645 & ~n10650;
  assign n10652 = ~n10644 & ~n10651;
  assign n10653 = po30  & ~n10652;
  assign n10654 = ~po30  & n10652;
  assign n10655 = ~n10208 & ~n10209;
  assign n10656 = po16  & n10655;
  assign n10657 = ~n10214 & ~n10656;
  assign n10658 = n10214 & n10656;
  assign n10659 = ~n10657 & ~n10658;
  assign n10660 = ~n10654 & ~n10659;
  assign n10661 = ~n10653 & ~n10660;
  assign n10662 = po31  & ~n10661;
  assign n10663 = ~po31  & n10661;
  assign n10664 = ~n10217 & ~n10218;
  assign n10665 = po16  & n10664;
  assign n10666 = ~n10223 & ~n10665;
  assign n10667 = n10223 & n10665;
  assign n10668 = ~n10666 & ~n10667;
  assign n10669 = ~n10663 & ~n10668;
  assign n10670 = ~n10662 & ~n10669;
  assign n10671 = po32  & ~n10670;
  assign n10672 = ~po32  & n10670;
  assign n10673 = ~n10226 & ~n10227;
  assign n10674 = po16  & n10673;
  assign n10675 = ~n10232 & ~n10674;
  assign n10676 = n10232 & n10674;
  assign n10677 = ~n10675 & ~n10676;
  assign n10678 = ~n10672 & ~n10677;
  assign n10679 = ~n10671 & ~n10678;
  assign n10680 = po33  & ~n10679;
  assign n10681 = ~po33  & n10679;
  assign n10682 = ~n10235 & ~n10236;
  assign n10683 = po16  & n10682;
  assign n10684 = ~n10241 & ~n10683;
  assign n10685 = n10241 & n10683;
  assign n10686 = ~n10684 & ~n10685;
  assign n10687 = ~n10681 & ~n10686;
  assign n10688 = ~n10680 & ~n10687;
  assign n10689 = po34  & ~n10688;
  assign n10690 = ~po34  & n10688;
  assign n10691 = ~n10244 & ~n10245;
  assign n10692 = po16  & n10691;
  assign n10693 = ~n10250 & ~n10692;
  assign n10694 = n10250 & n10692;
  assign n10695 = ~n10693 & ~n10694;
  assign n10696 = ~n10690 & ~n10695;
  assign n10697 = ~n10689 & ~n10696;
  assign n10698 = po35  & ~n10697;
  assign n10699 = ~po35  & n10697;
  assign n10700 = ~n10253 & ~n10254;
  assign n10701 = po16  & n10700;
  assign n10702 = ~n10259 & ~n10701;
  assign n10703 = n10259 & n10701;
  assign n10704 = ~n10702 & ~n10703;
  assign n10705 = ~n10699 & ~n10704;
  assign n10706 = ~n10698 & ~n10705;
  assign n10707 = po36  & ~n10706;
  assign n10708 = ~po36  & n10706;
  assign n10709 = ~n10262 & ~n10263;
  assign n10710 = po16  & n10709;
  assign n10711 = ~n10268 & ~n10710;
  assign n10712 = n10268 & n10710;
  assign n10713 = ~n10711 & ~n10712;
  assign n10714 = ~n10708 & ~n10713;
  assign n10715 = ~n10707 & ~n10714;
  assign n10716 = po37  & ~n10715;
  assign n10717 = ~po37  & n10715;
  assign n10718 = ~n10271 & ~n10272;
  assign n10719 = po16  & n10718;
  assign n10720 = ~n10277 & ~n10719;
  assign n10721 = n10277 & n10719;
  assign n10722 = ~n10720 & ~n10721;
  assign n10723 = ~n10717 & ~n10722;
  assign n10724 = ~n10716 & ~n10723;
  assign n10725 = po38  & ~n10724;
  assign n10726 = ~po38  & n10724;
  assign n10727 = ~n10280 & ~n10281;
  assign n10728 = po16  & n10727;
  assign n10729 = ~n10286 & ~n10728;
  assign n10730 = n10286 & n10728;
  assign n10731 = ~n10729 & ~n10730;
  assign n10732 = ~n10726 & ~n10731;
  assign n10733 = ~n10725 & ~n10732;
  assign n10734 = po39  & ~n10733;
  assign n10735 = ~po39  & n10733;
  assign n10736 = ~n10289 & ~n10290;
  assign n10737 = po16  & n10736;
  assign n10738 = ~n10295 & ~n10737;
  assign n10739 = n10295 & n10737;
  assign n10740 = ~n10738 & ~n10739;
  assign n10741 = ~n10735 & ~n10740;
  assign n10742 = ~n10734 & ~n10741;
  assign n10743 = po40  & ~n10742;
  assign n10744 = ~po40  & n10742;
  assign n10745 = ~n10298 & ~n10299;
  assign n10746 = po16  & n10745;
  assign n10747 = ~n10304 & ~n10746;
  assign n10748 = n10304 & n10746;
  assign n10749 = ~n10747 & ~n10748;
  assign n10750 = ~n10744 & ~n10749;
  assign n10751 = ~n10743 & ~n10750;
  assign n10752 = po41  & ~n10751;
  assign n10753 = ~po41  & n10751;
  assign n10754 = ~n10307 & ~n10308;
  assign n10755 = po16  & n10754;
  assign n10756 = ~n10313 & ~n10755;
  assign n10757 = n10313 & n10755;
  assign n10758 = ~n10756 & ~n10757;
  assign n10759 = ~n10753 & ~n10758;
  assign n10760 = ~n10752 & ~n10759;
  assign n10761 = po42  & ~n10760;
  assign n10762 = ~po42  & n10760;
  assign n10763 = ~n10316 & ~n10317;
  assign n10764 = po16  & n10763;
  assign n10765 = ~n10322 & ~n10764;
  assign n10766 = n10322 & n10764;
  assign n10767 = ~n10765 & ~n10766;
  assign n10768 = ~n10762 & ~n10767;
  assign n10769 = ~n10761 & ~n10768;
  assign n10770 = po43  & ~n10769;
  assign n10771 = ~po43  & n10769;
  assign n10772 = ~n10325 & ~n10326;
  assign n10773 = po16  & n10772;
  assign n10774 = ~n10331 & ~n10773;
  assign n10775 = n10331 & n10773;
  assign n10776 = ~n10774 & ~n10775;
  assign n10777 = ~n10771 & ~n10776;
  assign n10778 = ~n10770 & ~n10777;
  assign n10779 = po44  & ~n10778;
  assign n10780 = ~po44  & n10778;
  assign n10781 = ~n10334 & ~n10335;
  assign n10782 = po16  & n10781;
  assign n10783 = ~n10340 & ~n10782;
  assign n10784 = n10340 & n10782;
  assign n10785 = ~n10783 & ~n10784;
  assign n10786 = ~n10780 & ~n10785;
  assign n10787 = ~n10779 & ~n10786;
  assign n10788 = po45  & ~n10787;
  assign n10789 = ~po45  & n10787;
  assign n10790 = ~n10343 & ~n10344;
  assign n10791 = po16  & n10790;
  assign n10792 = ~n10349 & ~n10791;
  assign n10793 = n10349 & n10791;
  assign n10794 = ~n10792 & ~n10793;
  assign n10795 = ~n10789 & ~n10794;
  assign n10796 = ~n10788 & ~n10795;
  assign n10797 = po46  & ~n10796;
  assign n10798 = ~po46  & n10796;
  assign n10799 = ~n10352 & ~n10353;
  assign n10800 = po16  & n10799;
  assign n10801 = ~n10358 & ~n10800;
  assign n10802 = n10358 & n10800;
  assign n10803 = ~n10801 & ~n10802;
  assign n10804 = ~n10798 & ~n10803;
  assign n10805 = ~n10797 & ~n10804;
  assign n10806 = po47  & ~n10805;
  assign n10807 = ~po47  & n10805;
  assign n10808 = ~n10361 & ~n10362;
  assign n10809 = po16  & n10808;
  assign n10810 = ~n10367 & ~n10809;
  assign n10811 = n10367 & n10809;
  assign n10812 = ~n10810 & ~n10811;
  assign n10813 = ~n10807 & ~n10812;
  assign n10814 = ~n10806 & ~n10813;
  assign n10815 = po48  & ~n10814;
  assign n10816 = ~n10370 & ~n10376;
  assign n10817 = po16  & n10816;
  assign n10818 = ~n10375 & ~n10817;
  assign n10819 = n10375 & n10817;
  assign n10820 = ~n10818 & ~n10819;
  assign n10821 = ~po48  & n10814;
  assign n10822 = ~n10820 & ~n10821;
  assign n10823 = ~n10815 & ~n10822;
  assign n10824 = po49  & ~n10823;
  assign n10825 = ~po49  & n10823;
  assign n10826 = ~n10522 & ~n10825;
  assign n10827 = ~n10824 & ~n10826;
  assign n10828 = po50  & ~n10827;
  assign n10829 = ~po50  & n10827;
  assign n10830 = ~n10383 & ~n10384;
  assign n10831 = po16  & n10830;
  assign n10832 = ~n10389 & ~n10831;
  assign n10833 = n10389 & n10831;
  assign n10834 = ~n10832 & ~n10833;
  assign n10835 = ~n10829 & ~n10834;
  assign n10836 = ~n10828 & ~n10835;
  assign n10837 = po51  & ~n10836;
  assign n10838 = ~po51  & n10836;
  assign n10839 = ~n10392 & ~n10393;
  assign n10840 = po16  & n10839;
  assign n10841 = ~n10398 & ~n10840;
  assign n10842 = n10398 & n10840;
  assign n10843 = ~n10841 & ~n10842;
  assign n10844 = ~n10838 & ~n10843;
  assign n10845 = ~n10837 & ~n10844;
  assign n10846 = po52  & ~n10845;
  assign n10847 = ~po52  & n10845;
  assign n10848 = ~n10401 & ~n10402;
  assign n10849 = po16  & n10848;
  assign n10850 = ~n10407 & ~n10849;
  assign n10851 = n10407 & n10849;
  assign n10852 = ~n10850 & ~n10851;
  assign n10853 = ~n10847 & ~n10852;
  assign n10854 = ~n10846 & ~n10853;
  assign n10855 = po53  & ~n10854;
  assign n10856 = ~po53  & n10854;
  assign n10857 = ~n10410 & ~n10411;
  assign n10858 = po16  & n10857;
  assign n10859 = ~n10416 & ~n10858;
  assign n10860 = n10416 & n10858;
  assign n10861 = ~n10859 & ~n10860;
  assign n10862 = ~n10856 & ~n10861;
  assign n10863 = ~n10855 & ~n10862;
  assign n10864 = po54  & ~n10863;
  assign n10865 = ~po54  & n10863;
  assign n10866 = ~n10419 & ~n10420;
  assign n10867 = po16  & n10866;
  assign n10868 = ~n10425 & ~n10867;
  assign n10869 = n10425 & n10867;
  assign n10870 = ~n10868 & ~n10869;
  assign n10871 = ~n10865 & ~n10870;
  assign n10872 = ~n10864 & ~n10871;
  assign n10873 = po55  & ~n10872;
  assign n10874 = ~po55  & n10872;
  assign n10875 = ~n10428 & ~n10429;
  assign n10876 = po16  & n10875;
  assign n10877 = ~n10434 & ~n10876;
  assign n10878 = n10434 & n10876;
  assign n10879 = ~n10877 & ~n10878;
  assign n10880 = ~n10874 & ~n10879;
  assign n10881 = ~n10873 & ~n10880;
  assign n10882 = po56  & ~n10881;
  assign n10883 = ~po56  & n10881;
  assign n10884 = ~n10437 & ~n10438;
  assign n10885 = po16  & n10884;
  assign n10886 = ~n10443 & ~n10885;
  assign n10887 = n10443 & n10885;
  assign n10888 = ~n10886 & ~n10887;
  assign n10889 = ~n10883 & ~n10888;
  assign n10890 = ~n10882 & ~n10889;
  assign n10891 = po57  & ~n10890;
  assign n10892 = ~po57  & n10890;
  assign n10893 = ~n10446 & ~n10447;
  assign n10894 = po16  & n10893;
  assign n10895 = ~n10452 & ~n10894;
  assign n10896 = n10452 & n10894;
  assign n10897 = ~n10895 & ~n10896;
  assign n10898 = ~n10892 & ~n10897;
  assign n10899 = ~n10891 & ~n10898;
  assign n10900 = po58  & ~n10899;
  assign n10901 = ~po58  & n10899;
  assign n10902 = ~n10455 & ~n10456;
  assign n10903 = po16  & n10902;
  assign n10904 = ~n10461 & ~n10903;
  assign n10905 = n10461 & n10903;
  assign n10906 = ~n10904 & ~n10905;
  assign n10907 = ~n10901 & ~n10906;
  assign n10908 = ~n10900 & ~n10907;
  assign n10909 = po59  & ~n10908;
  assign n10910 = ~po59  & n10908;
  assign n10911 = ~n10464 & ~n10465;
  assign n10912 = po16  & n10911;
  assign n10913 = ~n10470 & ~n10912;
  assign n10914 = n10470 & n10912;
  assign n10915 = ~n10913 & ~n10914;
  assign n10916 = ~n10910 & ~n10915;
  assign n10917 = ~n10909 & ~n10916;
  assign n10918 = po60  & ~n10917;
  assign n10919 = ~po60  & n10917;
  assign n10920 = ~n10473 & ~n10474;
  assign n10921 = po16  & n10920;
  assign n10922 = ~n10479 & ~n10921;
  assign n10923 = n10479 & n10921;
  assign n10924 = ~n10922 & ~n10923;
  assign n10925 = ~n10919 & ~n10924;
  assign n10926 = ~n10918 & ~n10925;
  assign n10927 = po61  & ~n10926;
  assign n10928 = ~po61  & n10926;
  assign n10929 = ~n10482 & ~n10483;
  assign n10930 = po16  & n10929;
  assign n10931 = ~n10488 & ~n10930;
  assign n10932 = n10488 & n10930;
  assign n10933 = ~n10931 & ~n10932;
  assign n10934 = ~n10928 & ~n10933;
  assign n10935 = ~n10927 & ~n10934;
  assign n10936 = po62  & ~n10935;
  assign n10937 = ~po62  & n10935;
  assign n10938 = ~n10491 & ~n10492;
  assign n10939 = po16  & n10938;
  assign n10940 = ~n10497 & ~n10939;
  assign n10941 = n10497 & n10939;
  assign n10942 = ~n10940 & ~n10941;
  assign n10943 = ~n10937 & ~n10942;
  assign n10944 = ~n10936 & ~n10943;
  assign n10945 = n10532 & n10944;
  assign n10946 = ~n10532 & ~n10944;
  assign n10947 = n10510 & po16 ;
  assign n10948 = ~n10509 & ~n10947;
  assign n10949 = n10946 & n10948;
  assign n10950 = ~po63  & ~n10949;
  assign n10951 = ~n10945 & ~n10950;
  assign n10952 = ~n10527 & n10951;
  assign po15  = n10523 | ~n10952;
  assign n10954 = ~n10824 & ~n10825;
  assign n10955 = po15  & n10954;
  assign n10956 = ~n10522 & ~n10955;
  assign n10957 = n10522 & n10955;
  assign n10958 = ~n10956 & ~n10957;
  assign n10959 = n10532 & ~po15 ;
  assign n10960 = ~n10532 & po15 ;
  assign n10961 = n10944 & ~n10960;
  assign n10962 = po63  & ~n10961;
  assign n10963 = ~n10946 & n10962;
  assign n10964 = ~n10936 & ~n10937;
  assign n10965 = po15  & n10964;
  assign n10966 = ~n10942 & ~n10965;
  assign n10967 = n10942 & n10965;
  assign n10968 = ~n10966 & ~n10967;
  assign n10969 = pi30  & po15 ;
  assign n10970 = ~pi28  & ~pi29 ;
  assign n10971 = ~pi30  & n10970;
  assign n10972 = ~n10969 & ~n10971;
  assign n10973 = po16  & ~n10972;
  assign n10974 = ~po16  & n10972;
  assign n10975 = ~pi30  & po15 ;
  assign n10976 = pi31  & ~n10975;
  assign n10977 = n10534 & po15 ;
  assign n10978 = ~n10976 & ~n10977;
  assign n10979 = ~n10974 & n10978;
  assign n10980 = ~n10973 & ~n10979;
  assign n10981 = po17  & ~n10980;
  assign n10982 = ~po17  & n10980;
  assign n10983 = po16  & n10952;
  assign n10984 = ~n10977 & ~n10983;
  assign n10985 = pi32  & ~n10984;
  assign n10986 = ~pi32  & n10984;
  assign n10987 = ~n10985 & ~n10986;
  assign n10988 = ~n10982 & ~n10987;
  assign n10989 = ~n10981 & ~n10988;
  assign n10990 = po18  & ~n10989;
  assign n10991 = ~po18  & n10989;
  assign n10992 = ~n10537 & ~n10538;
  assign n10993 = po15  & n10992;
  assign n10994 = n10542 & ~n10993;
  assign n10995 = ~n10542 & n10993;
  assign n10996 = ~n10994 & ~n10995;
  assign n10997 = ~n10991 & ~n10996;
  assign n10998 = ~n10990 & ~n10997;
  assign n10999 = po19  & ~n10998;
  assign n11000 = ~po19  & n10998;
  assign n11001 = ~n10545 & ~n10546;
  assign n11002 = po15  & n11001;
  assign n11003 = ~n10551 & ~n11002;
  assign n11004 = n10551 & n11002;
  assign n11005 = ~n11003 & ~n11004;
  assign n11006 = ~n11000 & ~n11005;
  assign n11007 = ~n10999 & ~n11006;
  assign n11008 = po20  & ~n11007;
  assign n11009 = ~po20  & n11007;
  assign n11010 = ~n10554 & ~n10555;
  assign n11011 = po15  & n11010;
  assign n11012 = n10560 & n11011;
  assign n11013 = ~n10560 & ~n11011;
  assign n11014 = ~n11012 & ~n11013;
  assign n11015 = ~n11009 & ~n11014;
  assign n11016 = ~n11008 & ~n11015;
  assign n11017 = po21  & ~n11016;
  assign n11018 = ~po21  & n11016;
  assign n11019 = ~n10563 & ~n10564;
  assign n11020 = po15  & n11019;
  assign n11021 = ~n10569 & ~n11020;
  assign n11022 = n10569 & n11020;
  assign n11023 = ~n11021 & ~n11022;
  assign n11024 = ~n11018 & ~n11023;
  assign n11025 = ~n11017 & ~n11024;
  assign n11026 = po22  & ~n11025;
  assign n11027 = ~po22  & n11025;
  assign n11028 = ~n10572 & ~n10573;
  assign n11029 = po15  & n11028;
  assign n11030 = ~n10578 & ~n11029;
  assign n11031 = n10578 & n11029;
  assign n11032 = ~n11030 & ~n11031;
  assign n11033 = ~n11027 & ~n11032;
  assign n11034 = ~n11026 & ~n11033;
  assign n11035 = po23  & ~n11034;
  assign n11036 = ~po23  & n11034;
  assign n11037 = ~n10581 & ~n10582;
  assign n11038 = po15  & n11037;
  assign n11039 = ~n10587 & ~n11038;
  assign n11040 = n10587 & n11038;
  assign n11041 = ~n11039 & ~n11040;
  assign n11042 = ~n11036 & ~n11041;
  assign n11043 = ~n11035 & ~n11042;
  assign n11044 = po24  & ~n11043;
  assign n11045 = ~po24  & n11043;
  assign n11046 = ~n10590 & ~n10591;
  assign n11047 = po15  & n11046;
  assign n11048 = ~n10596 & ~n11047;
  assign n11049 = n10596 & n11047;
  assign n11050 = ~n11048 & ~n11049;
  assign n11051 = ~n11045 & ~n11050;
  assign n11052 = ~n11044 & ~n11051;
  assign n11053 = po25  & ~n11052;
  assign n11054 = ~po25  & n11052;
  assign n11055 = ~n10599 & ~n10600;
  assign n11056 = po15  & n11055;
  assign n11057 = ~n10605 & ~n11056;
  assign n11058 = n10605 & n11056;
  assign n11059 = ~n11057 & ~n11058;
  assign n11060 = ~n11054 & ~n11059;
  assign n11061 = ~n11053 & ~n11060;
  assign n11062 = po26  & ~n11061;
  assign n11063 = ~po26  & n11061;
  assign n11064 = ~n10608 & ~n10609;
  assign n11065 = po15  & n11064;
  assign n11066 = ~n10614 & ~n11065;
  assign n11067 = n10614 & n11065;
  assign n11068 = ~n11066 & ~n11067;
  assign n11069 = ~n11063 & ~n11068;
  assign n11070 = ~n11062 & ~n11069;
  assign n11071 = po27  & ~n11070;
  assign n11072 = ~po27  & n11070;
  assign n11073 = ~n10617 & ~n10618;
  assign n11074 = po15  & n11073;
  assign n11075 = ~n10623 & ~n11074;
  assign n11076 = n10623 & n11074;
  assign n11077 = ~n11075 & ~n11076;
  assign n11078 = ~n11072 & ~n11077;
  assign n11079 = ~n11071 & ~n11078;
  assign n11080 = po28  & ~n11079;
  assign n11081 = ~po28  & n11079;
  assign n11082 = ~n10626 & ~n10627;
  assign n11083 = po15  & n11082;
  assign n11084 = ~n10632 & ~n11083;
  assign n11085 = n10632 & n11083;
  assign n11086 = ~n11084 & ~n11085;
  assign n11087 = ~n11081 & ~n11086;
  assign n11088 = ~n11080 & ~n11087;
  assign n11089 = po29  & ~n11088;
  assign n11090 = ~po29  & n11088;
  assign n11091 = ~n10635 & ~n10636;
  assign n11092 = po15  & n11091;
  assign n11093 = ~n10641 & ~n11092;
  assign n11094 = n10641 & n11092;
  assign n11095 = ~n11093 & ~n11094;
  assign n11096 = ~n11090 & ~n11095;
  assign n11097 = ~n11089 & ~n11096;
  assign n11098 = po30  & ~n11097;
  assign n11099 = ~po30  & n11097;
  assign n11100 = ~n10644 & ~n10645;
  assign n11101 = po15  & n11100;
  assign n11102 = ~n10650 & ~n11101;
  assign n11103 = n10650 & n11101;
  assign n11104 = ~n11102 & ~n11103;
  assign n11105 = ~n11099 & ~n11104;
  assign n11106 = ~n11098 & ~n11105;
  assign n11107 = po31  & ~n11106;
  assign n11108 = ~po31  & n11106;
  assign n11109 = ~n10653 & ~n10654;
  assign n11110 = po15  & n11109;
  assign n11111 = ~n10659 & ~n11110;
  assign n11112 = n10659 & n11110;
  assign n11113 = ~n11111 & ~n11112;
  assign n11114 = ~n11108 & ~n11113;
  assign n11115 = ~n11107 & ~n11114;
  assign n11116 = po32  & ~n11115;
  assign n11117 = ~po32  & n11115;
  assign n11118 = ~n10662 & ~n10663;
  assign n11119 = po15  & n11118;
  assign n11120 = ~n10668 & ~n11119;
  assign n11121 = n10668 & n11119;
  assign n11122 = ~n11120 & ~n11121;
  assign n11123 = ~n11117 & ~n11122;
  assign n11124 = ~n11116 & ~n11123;
  assign n11125 = po33  & ~n11124;
  assign n11126 = ~po33  & n11124;
  assign n11127 = ~n10671 & ~n10672;
  assign n11128 = po15  & n11127;
  assign n11129 = ~n10677 & ~n11128;
  assign n11130 = n10677 & n11128;
  assign n11131 = ~n11129 & ~n11130;
  assign n11132 = ~n11126 & ~n11131;
  assign n11133 = ~n11125 & ~n11132;
  assign n11134 = po34  & ~n11133;
  assign n11135 = ~po34  & n11133;
  assign n11136 = ~n10680 & ~n10681;
  assign n11137 = po15  & n11136;
  assign n11138 = ~n10686 & ~n11137;
  assign n11139 = n10686 & n11137;
  assign n11140 = ~n11138 & ~n11139;
  assign n11141 = ~n11135 & ~n11140;
  assign n11142 = ~n11134 & ~n11141;
  assign n11143 = po35  & ~n11142;
  assign n11144 = ~po35  & n11142;
  assign n11145 = ~n10689 & ~n10690;
  assign n11146 = po15  & n11145;
  assign n11147 = ~n10695 & ~n11146;
  assign n11148 = n10695 & n11146;
  assign n11149 = ~n11147 & ~n11148;
  assign n11150 = ~n11144 & ~n11149;
  assign n11151 = ~n11143 & ~n11150;
  assign n11152 = po36  & ~n11151;
  assign n11153 = ~po36  & n11151;
  assign n11154 = ~n10698 & ~n10699;
  assign n11155 = po15  & n11154;
  assign n11156 = ~n10704 & ~n11155;
  assign n11157 = n10704 & n11155;
  assign n11158 = ~n11156 & ~n11157;
  assign n11159 = ~n11153 & ~n11158;
  assign n11160 = ~n11152 & ~n11159;
  assign n11161 = po37  & ~n11160;
  assign n11162 = ~po37  & n11160;
  assign n11163 = ~n10707 & ~n10708;
  assign n11164 = po15  & n11163;
  assign n11165 = ~n10713 & ~n11164;
  assign n11166 = n10713 & n11164;
  assign n11167 = ~n11165 & ~n11166;
  assign n11168 = ~n11162 & ~n11167;
  assign n11169 = ~n11161 & ~n11168;
  assign n11170 = po38  & ~n11169;
  assign n11171 = ~po38  & n11169;
  assign n11172 = ~n10716 & ~n10717;
  assign n11173 = po15  & n11172;
  assign n11174 = ~n10722 & ~n11173;
  assign n11175 = n10722 & n11173;
  assign n11176 = ~n11174 & ~n11175;
  assign n11177 = ~n11171 & ~n11176;
  assign n11178 = ~n11170 & ~n11177;
  assign n11179 = po39  & ~n11178;
  assign n11180 = ~po39  & n11178;
  assign n11181 = ~n10725 & ~n10726;
  assign n11182 = po15  & n11181;
  assign n11183 = ~n10731 & ~n11182;
  assign n11184 = n10731 & n11182;
  assign n11185 = ~n11183 & ~n11184;
  assign n11186 = ~n11180 & ~n11185;
  assign n11187 = ~n11179 & ~n11186;
  assign n11188 = po40  & ~n11187;
  assign n11189 = ~po40  & n11187;
  assign n11190 = ~n10734 & ~n10735;
  assign n11191 = po15  & n11190;
  assign n11192 = ~n10740 & ~n11191;
  assign n11193 = n10740 & n11191;
  assign n11194 = ~n11192 & ~n11193;
  assign n11195 = ~n11189 & ~n11194;
  assign n11196 = ~n11188 & ~n11195;
  assign n11197 = po41  & ~n11196;
  assign n11198 = ~po41  & n11196;
  assign n11199 = ~n10743 & ~n10744;
  assign n11200 = po15  & n11199;
  assign n11201 = ~n10749 & ~n11200;
  assign n11202 = n10749 & n11200;
  assign n11203 = ~n11201 & ~n11202;
  assign n11204 = ~n11198 & ~n11203;
  assign n11205 = ~n11197 & ~n11204;
  assign n11206 = po42  & ~n11205;
  assign n11207 = ~po42  & n11205;
  assign n11208 = ~n10752 & ~n10753;
  assign n11209 = po15  & n11208;
  assign n11210 = ~n10758 & ~n11209;
  assign n11211 = n10758 & n11209;
  assign n11212 = ~n11210 & ~n11211;
  assign n11213 = ~n11207 & ~n11212;
  assign n11214 = ~n11206 & ~n11213;
  assign n11215 = po43  & ~n11214;
  assign n11216 = ~po43  & n11214;
  assign n11217 = ~n10761 & ~n10762;
  assign n11218 = po15  & n11217;
  assign n11219 = ~n10767 & ~n11218;
  assign n11220 = n10767 & n11218;
  assign n11221 = ~n11219 & ~n11220;
  assign n11222 = ~n11216 & ~n11221;
  assign n11223 = ~n11215 & ~n11222;
  assign n11224 = po44  & ~n11223;
  assign n11225 = ~po44  & n11223;
  assign n11226 = ~n10770 & ~n10771;
  assign n11227 = po15  & n11226;
  assign n11228 = ~n10776 & ~n11227;
  assign n11229 = n10776 & n11227;
  assign n11230 = ~n11228 & ~n11229;
  assign n11231 = ~n11225 & ~n11230;
  assign n11232 = ~n11224 & ~n11231;
  assign n11233 = po45  & ~n11232;
  assign n11234 = ~po45  & n11232;
  assign n11235 = ~n10779 & ~n10780;
  assign n11236 = po15  & n11235;
  assign n11237 = ~n10785 & ~n11236;
  assign n11238 = n10785 & n11236;
  assign n11239 = ~n11237 & ~n11238;
  assign n11240 = ~n11234 & ~n11239;
  assign n11241 = ~n11233 & ~n11240;
  assign n11242 = po46  & ~n11241;
  assign n11243 = ~po46  & n11241;
  assign n11244 = ~n10788 & ~n10789;
  assign n11245 = po15  & n11244;
  assign n11246 = ~n10794 & ~n11245;
  assign n11247 = n10794 & n11245;
  assign n11248 = ~n11246 & ~n11247;
  assign n11249 = ~n11243 & ~n11248;
  assign n11250 = ~n11242 & ~n11249;
  assign n11251 = po47  & ~n11250;
  assign n11252 = ~po47  & n11250;
  assign n11253 = ~n10797 & ~n10798;
  assign n11254 = po15  & n11253;
  assign n11255 = ~n10803 & ~n11254;
  assign n11256 = n10803 & n11254;
  assign n11257 = ~n11255 & ~n11256;
  assign n11258 = ~n11252 & ~n11257;
  assign n11259 = ~n11251 & ~n11258;
  assign n11260 = po48  & ~n11259;
  assign n11261 = ~po48  & n11259;
  assign n11262 = ~n10806 & ~n10807;
  assign n11263 = po15  & n11262;
  assign n11264 = ~n10812 & ~n11263;
  assign n11265 = n10812 & n11263;
  assign n11266 = ~n11264 & ~n11265;
  assign n11267 = ~n11261 & ~n11266;
  assign n11268 = ~n11260 & ~n11267;
  assign n11269 = po49  & ~n11268;
  assign n11270 = ~n10815 & ~n10821;
  assign n11271 = po15  & n11270;
  assign n11272 = ~n10820 & ~n11271;
  assign n11273 = n10820 & n11271;
  assign n11274 = ~n11272 & ~n11273;
  assign n11275 = ~po49  & n11268;
  assign n11276 = ~n11274 & ~n11275;
  assign n11277 = ~n11269 & ~n11276;
  assign n11278 = po50  & ~n11277;
  assign n11279 = ~po50  & n11277;
  assign n11280 = ~n10958 & ~n11279;
  assign n11281 = ~n11278 & ~n11280;
  assign n11282 = po51  & ~n11281;
  assign n11283 = ~po51  & n11281;
  assign n11284 = ~n10828 & ~n10829;
  assign n11285 = po15  & n11284;
  assign n11286 = ~n10834 & ~n11285;
  assign n11287 = n10834 & n11285;
  assign n11288 = ~n11286 & ~n11287;
  assign n11289 = ~n11283 & ~n11288;
  assign n11290 = ~n11282 & ~n11289;
  assign n11291 = po52  & ~n11290;
  assign n11292 = ~po52  & n11290;
  assign n11293 = ~n10837 & ~n10838;
  assign n11294 = po15  & n11293;
  assign n11295 = ~n10843 & ~n11294;
  assign n11296 = n10843 & n11294;
  assign n11297 = ~n11295 & ~n11296;
  assign n11298 = ~n11292 & ~n11297;
  assign n11299 = ~n11291 & ~n11298;
  assign n11300 = po53  & ~n11299;
  assign n11301 = ~po53  & n11299;
  assign n11302 = ~n10846 & ~n10847;
  assign n11303 = po15  & n11302;
  assign n11304 = ~n10852 & ~n11303;
  assign n11305 = n10852 & n11303;
  assign n11306 = ~n11304 & ~n11305;
  assign n11307 = ~n11301 & ~n11306;
  assign n11308 = ~n11300 & ~n11307;
  assign n11309 = po54  & ~n11308;
  assign n11310 = ~po54  & n11308;
  assign n11311 = ~n10855 & ~n10856;
  assign n11312 = po15  & n11311;
  assign n11313 = ~n10861 & ~n11312;
  assign n11314 = n10861 & n11312;
  assign n11315 = ~n11313 & ~n11314;
  assign n11316 = ~n11310 & ~n11315;
  assign n11317 = ~n11309 & ~n11316;
  assign n11318 = po55  & ~n11317;
  assign n11319 = ~po55  & n11317;
  assign n11320 = ~n10864 & ~n10865;
  assign n11321 = po15  & n11320;
  assign n11322 = ~n10870 & ~n11321;
  assign n11323 = n10870 & n11321;
  assign n11324 = ~n11322 & ~n11323;
  assign n11325 = ~n11319 & ~n11324;
  assign n11326 = ~n11318 & ~n11325;
  assign n11327 = po56  & ~n11326;
  assign n11328 = ~po56  & n11326;
  assign n11329 = ~n10873 & ~n10874;
  assign n11330 = po15  & n11329;
  assign n11331 = ~n10879 & ~n11330;
  assign n11332 = n10879 & n11330;
  assign n11333 = ~n11331 & ~n11332;
  assign n11334 = ~n11328 & ~n11333;
  assign n11335 = ~n11327 & ~n11334;
  assign n11336 = po57  & ~n11335;
  assign n11337 = ~po57  & n11335;
  assign n11338 = ~n10882 & ~n10883;
  assign n11339 = po15  & n11338;
  assign n11340 = ~n10888 & ~n11339;
  assign n11341 = n10888 & n11339;
  assign n11342 = ~n11340 & ~n11341;
  assign n11343 = ~n11337 & ~n11342;
  assign n11344 = ~n11336 & ~n11343;
  assign n11345 = po58  & ~n11344;
  assign n11346 = ~po58  & n11344;
  assign n11347 = ~n10891 & ~n10892;
  assign n11348 = po15  & n11347;
  assign n11349 = ~n10897 & ~n11348;
  assign n11350 = n10897 & n11348;
  assign n11351 = ~n11349 & ~n11350;
  assign n11352 = ~n11346 & ~n11351;
  assign n11353 = ~n11345 & ~n11352;
  assign n11354 = po59  & ~n11353;
  assign n11355 = ~po59  & n11353;
  assign n11356 = ~n10900 & ~n10901;
  assign n11357 = po15  & n11356;
  assign n11358 = ~n10906 & ~n11357;
  assign n11359 = n10906 & n11357;
  assign n11360 = ~n11358 & ~n11359;
  assign n11361 = ~n11355 & ~n11360;
  assign n11362 = ~n11354 & ~n11361;
  assign n11363 = po60  & ~n11362;
  assign n11364 = ~po60  & n11362;
  assign n11365 = ~n10909 & ~n10910;
  assign n11366 = po15  & n11365;
  assign n11367 = ~n10915 & ~n11366;
  assign n11368 = n10915 & n11366;
  assign n11369 = ~n11367 & ~n11368;
  assign n11370 = ~n11364 & ~n11369;
  assign n11371 = ~n11363 & ~n11370;
  assign n11372 = po61  & ~n11371;
  assign n11373 = ~po61  & n11371;
  assign n11374 = ~n10918 & ~n10919;
  assign n11375 = po15  & n11374;
  assign n11376 = ~n10924 & ~n11375;
  assign n11377 = n10924 & n11375;
  assign n11378 = ~n11376 & ~n11377;
  assign n11379 = ~n11373 & ~n11378;
  assign n11380 = ~n11372 & ~n11379;
  assign n11381 = po62  & ~n11380;
  assign n11382 = ~po62  & n11380;
  assign n11383 = ~n10927 & ~n10928;
  assign n11384 = po15  & n11383;
  assign n11385 = ~n10933 & ~n11384;
  assign n11386 = n10933 & n11384;
  assign n11387 = ~n11385 & ~n11386;
  assign n11388 = ~n11382 & ~n11387;
  assign n11389 = ~n11381 & ~n11388;
  assign n11390 = n10968 & n11389;
  assign n11391 = ~n10968 & ~n11389;
  assign n11392 = n10946 & po15 ;
  assign n11393 = ~n10945 & ~n11392;
  assign n11394 = n11391 & n11393;
  assign n11395 = ~po63  & ~n11394;
  assign n11396 = ~n11390 & ~n11395;
  assign n11397 = ~n10963 & n11396;
  assign po14  = n10959 | ~n11397;
  assign n11399 = ~n11278 & ~n11279;
  assign n11400 = po14  & n11399;
  assign n11401 = ~n10958 & ~n11400;
  assign n11402 = n10958 & n11400;
  assign n11403 = ~n11401 & ~n11402;
  assign n11404 = n10968 & ~po14 ;
  assign n11405 = ~n10968 & po14 ;
  assign n11406 = n11389 & ~n11405;
  assign n11407 = po63  & ~n11406;
  assign n11408 = ~n11391 & n11407;
  assign n11409 = ~n11381 & ~n11382;
  assign n11410 = po14  & n11409;
  assign n11411 = ~n11387 & ~n11410;
  assign n11412 = n11387 & n11410;
  assign n11413 = ~n11411 & ~n11412;
  assign n11414 = pi28  & po14 ;
  assign n11415 = ~pi26  & ~pi27 ;
  assign n11416 = ~pi28  & n11415;
  assign n11417 = ~n11414 & ~n11416;
  assign n11418 = po15  & ~n11417;
  assign n11419 = ~po15  & n11417;
  assign n11420 = ~pi28  & po14 ;
  assign n11421 = pi29  & ~n11420;
  assign n11422 = n10970 & po14 ;
  assign n11423 = ~n11421 & ~n11422;
  assign n11424 = ~n11419 & n11423;
  assign n11425 = ~n11418 & ~n11424;
  assign n11426 = po16  & ~n11425;
  assign n11427 = ~po16  & n11425;
  assign n11428 = po15  & n11397;
  assign n11429 = ~n11422 & ~n11428;
  assign n11430 = pi30  & ~n11429;
  assign n11431 = ~pi30  & n11429;
  assign n11432 = ~n11430 & ~n11431;
  assign n11433 = ~n11427 & ~n11432;
  assign n11434 = ~n11426 & ~n11433;
  assign n11435 = po17  & ~n11434;
  assign n11436 = ~po17  & n11434;
  assign n11437 = ~n10973 & ~n10974;
  assign n11438 = po14  & n11437;
  assign n11439 = n10978 & ~n11438;
  assign n11440 = ~n10978 & n11438;
  assign n11441 = ~n11439 & ~n11440;
  assign n11442 = ~n11436 & ~n11441;
  assign n11443 = ~n11435 & ~n11442;
  assign n11444 = po18  & ~n11443;
  assign n11445 = ~po18  & n11443;
  assign n11446 = ~n10981 & ~n10982;
  assign n11447 = po14  & n11446;
  assign n11448 = ~n10987 & ~n11447;
  assign n11449 = n10987 & n11447;
  assign n11450 = ~n11448 & ~n11449;
  assign n11451 = ~n11445 & ~n11450;
  assign n11452 = ~n11444 & ~n11451;
  assign n11453 = po19  & ~n11452;
  assign n11454 = ~po19  & n11452;
  assign n11455 = ~n10990 & ~n10991;
  assign n11456 = po14  & n11455;
  assign n11457 = n10996 & n11456;
  assign n11458 = ~n10996 & ~n11456;
  assign n11459 = ~n11457 & ~n11458;
  assign n11460 = ~n11454 & ~n11459;
  assign n11461 = ~n11453 & ~n11460;
  assign n11462 = po20  & ~n11461;
  assign n11463 = ~po20  & n11461;
  assign n11464 = ~n10999 & ~n11000;
  assign n11465 = po14  & n11464;
  assign n11466 = ~n11005 & ~n11465;
  assign n11467 = n11005 & n11465;
  assign n11468 = ~n11466 & ~n11467;
  assign n11469 = ~n11463 & ~n11468;
  assign n11470 = ~n11462 & ~n11469;
  assign n11471 = po21  & ~n11470;
  assign n11472 = ~po21  & n11470;
  assign n11473 = ~n11008 & ~n11009;
  assign n11474 = po14  & n11473;
  assign n11475 = ~n11014 & ~n11474;
  assign n11476 = n11014 & n11474;
  assign n11477 = ~n11475 & ~n11476;
  assign n11478 = ~n11472 & ~n11477;
  assign n11479 = ~n11471 & ~n11478;
  assign n11480 = po22  & ~n11479;
  assign n11481 = ~po22  & n11479;
  assign n11482 = ~n11017 & ~n11018;
  assign n11483 = po14  & n11482;
  assign n11484 = ~n11023 & ~n11483;
  assign n11485 = n11023 & n11483;
  assign n11486 = ~n11484 & ~n11485;
  assign n11487 = ~n11481 & ~n11486;
  assign n11488 = ~n11480 & ~n11487;
  assign n11489 = po23  & ~n11488;
  assign n11490 = ~po23  & n11488;
  assign n11491 = ~n11026 & ~n11027;
  assign n11492 = po14  & n11491;
  assign n11493 = ~n11032 & ~n11492;
  assign n11494 = n11032 & n11492;
  assign n11495 = ~n11493 & ~n11494;
  assign n11496 = ~n11490 & ~n11495;
  assign n11497 = ~n11489 & ~n11496;
  assign n11498 = po24  & ~n11497;
  assign n11499 = ~po24  & n11497;
  assign n11500 = ~n11035 & ~n11036;
  assign n11501 = po14  & n11500;
  assign n11502 = ~n11041 & ~n11501;
  assign n11503 = n11041 & n11501;
  assign n11504 = ~n11502 & ~n11503;
  assign n11505 = ~n11499 & ~n11504;
  assign n11506 = ~n11498 & ~n11505;
  assign n11507 = po25  & ~n11506;
  assign n11508 = ~po25  & n11506;
  assign n11509 = ~n11044 & ~n11045;
  assign n11510 = po14  & n11509;
  assign n11511 = ~n11050 & ~n11510;
  assign n11512 = n11050 & n11510;
  assign n11513 = ~n11511 & ~n11512;
  assign n11514 = ~n11508 & ~n11513;
  assign n11515 = ~n11507 & ~n11514;
  assign n11516 = po26  & ~n11515;
  assign n11517 = ~po26  & n11515;
  assign n11518 = ~n11053 & ~n11054;
  assign n11519 = po14  & n11518;
  assign n11520 = ~n11059 & ~n11519;
  assign n11521 = n11059 & n11519;
  assign n11522 = ~n11520 & ~n11521;
  assign n11523 = ~n11517 & ~n11522;
  assign n11524 = ~n11516 & ~n11523;
  assign n11525 = po27  & ~n11524;
  assign n11526 = ~po27  & n11524;
  assign n11527 = ~n11062 & ~n11063;
  assign n11528 = po14  & n11527;
  assign n11529 = ~n11068 & ~n11528;
  assign n11530 = n11068 & n11528;
  assign n11531 = ~n11529 & ~n11530;
  assign n11532 = ~n11526 & ~n11531;
  assign n11533 = ~n11525 & ~n11532;
  assign n11534 = po28  & ~n11533;
  assign n11535 = ~po28  & n11533;
  assign n11536 = ~n11071 & ~n11072;
  assign n11537 = po14  & n11536;
  assign n11538 = ~n11077 & ~n11537;
  assign n11539 = n11077 & n11537;
  assign n11540 = ~n11538 & ~n11539;
  assign n11541 = ~n11535 & ~n11540;
  assign n11542 = ~n11534 & ~n11541;
  assign n11543 = po29  & ~n11542;
  assign n11544 = ~po29  & n11542;
  assign n11545 = ~n11080 & ~n11081;
  assign n11546 = po14  & n11545;
  assign n11547 = ~n11086 & ~n11546;
  assign n11548 = n11086 & n11546;
  assign n11549 = ~n11547 & ~n11548;
  assign n11550 = ~n11544 & ~n11549;
  assign n11551 = ~n11543 & ~n11550;
  assign n11552 = po30  & ~n11551;
  assign n11553 = ~po30  & n11551;
  assign n11554 = ~n11089 & ~n11090;
  assign n11555 = po14  & n11554;
  assign n11556 = ~n11095 & ~n11555;
  assign n11557 = n11095 & n11555;
  assign n11558 = ~n11556 & ~n11557;
  assign n11559 = ~n11553 & ~n11558;
  assign n11560 = ~n11552 & ~n11559;
  assign n11561 = po31  & ~n11560;
  assign n11562 = ~po31  & n11560;
  assign n11563 = ~n11098 & ~n11099;
  assign n11564 = po14  & n11563;
  assign n11565 = ~n11104 & ~n11564;
  assign n11566 = n11104 & n11564;
  assign n11567 = ~n11565 & ~n11566;
  assign n11568 = ~n11562 & ~n11567;
  assign n11569 = ~n11561 & ~n11568;
  assign n11570 = po32  & ~n11569;
  assign n11571 = ~po32  & n11569;
  assign n11572 = ~n11107 & ~n11108;
  assign n11573 = po14  & n11572;
  assign n11574 = ~n11113 & ~n11573;
  assign n11575 = n11113 & n11573;
  assign n11576 = ~n11574 & ~n11575;
  assign n11577 = ~n11571 & ~n11576;
  assign n11578 = ~n11570 & ~n11577;
  assign n11579 = po33  & ~n11578;
  assign n11580 = ~po33  & n11578;
  assign n11581 = ~n11116 & ~n11117;
  assign n11582 = po14  & n11581;
  assign n11583 = ~n11122 & ~n11582;
  assign n11584 = n11122 & n11582;
  assign n11585 = ~n11583 & ~n11584;
  assign n11586 = ~n11580 & ~n11585;
  assign n11587 = ~n11579 & ~n11586;
  assign n11588 = po34  & ~n11587;
  assign n11589 = ~po34  & n11587;
  assign n11590 = ~n11125 & ~n11126;
  assign n11591 = po14  & n11590;
  assign n11592 = ~n11131 & ~n11591;
  assign n11593 = n11131 & n11591;
  assign n11594 = ~n11592 & ~n11593;
  assign n11595 = ~n11589 & ~n11594;
  assign n11596 = ~n11588 & ~n11595;
  assign n11597 = po35  & ~n11596;
  assign n11598 = ~po35  & n11596;
  assign n11599 = ~n11134 & ~n11135;
  assign n11600 = po14  & n11599;
  assign n11601 = ~n11140 & ~n11600;
  assign n11602 = n11140 & n11600;
  assign n11603 = ~n11601 & ~n11602;
  assign n11604 = ~n11598 & ~n11603;
  assign n11605 = ~n11597 & ~n11604;
  assign n11606 = po36  & ~n11605;
  assign n11607 = ~po36  & n11605;
  assign n11608 = ~n11143 & ~n11144;
  assign n11609 = po14  & n11608;
  assign n11610 = ~n11149 & ~n11609;
  assign n11611 = n11149 & n11609;
  assign n11612 = ~n11610 & ~n11611;
  assign n11613 = ~n11607 & ~n11612;
  assign n11614 = ~n11606 & ~n11613;
  assign n11615 = po37  & ~n11614;
  assign n11616 = ~po37  & n11614;
  assign n11617 = ~n11152 & ~n11153;
  assign n11618 = po14  & n11617;
  assign n11619 = ~n11158 & ~n11618;
  assign n11620 = n11158 & n11618;
  assign n11621 = ~n11619 & ~n11620;
  assign n11622 = ~n11616 & ~n11621;
  assign n11623 = ~n11615 & ~n11622;
  assign n11624 = po38  & ~n11623;
  assign n11625 = ~po38  & n11623;
  assign n11626 = ~n11161 & ~n11162;
  assign n11627 = po14  & n11626;
  assign n11628 = ~n11167 & ~n11627;
  assign n11629 = n11167 & n11627;
  assign n11630 = ~n11628 & ~n11629;
  assign n11631 = ~n11625 & ~n11630;
  assign n11632 = ~n11624 & ~n11631;
  assign n11633 = po39  & ~n11632;
  assign n11634 = ~po39  & n11632;
  assign n11635 = ~n11170 & ~n11171;
  assign n11636 = po14  & n11635;
  assign n11637 = ~n11176 & ~n11636;
  assign n11638 = n11176 & n11636;
  assign n11639 = ~n11637 & ~n11638;
  assign n11640 = ~n11634 & ~n11639;
  assign n11641 = ~n11633 & ~n11640;
  assign n11642 = po40  & ~n11641;
  assign n11643 = ~po40  & n11641;
  assign n11644 = ~n11179 & ~n11180;
  assign n11645 = po14  & n11644;
  assign n11646 = ~n11185 & ~n11645;
  assign n11647 = n11185 & n11645;
  assign n11648 = ~n11646 & ~n11647;
  assign n11649 = ~n11643 & ~n11648;
  assign n11650 = ~n11642 & ~n11649;
  assign n11651 = po41  & ~n11650;
  assign n11652 = ~po41  & n11650;
  assign n11653 = ~n11188 & ~n11189;
  assign n11654 = po14  & n11653;
  assign n11655 = ~n11194 & ~n11654;
  assign n11656 = n11194 & n11654;
  assign n11657 = ~n11655 & ~n11656;
  assign n11658 = ~n11652 & ~n11657;
  assign n11659 = ~n11651 & ~n11658;
  assign n11660 = po42  & ~n11659;
  assign n11661 = ~po42  & n11659;
  assign n11662 = ~n11197 & ~n11198;
  assign n11663 = po14  & n11662;
  assign n11664 = ~n11203 & ~n11663;
  assign n11665 = n11203 & n11663;
  assign n11666 = ~n11664 & ~n11665;
  assign n11667 = ~n11661 & ~n11666;
  assign n11668 = ~n11660 & ~n11667;
  assign n11669 = po43  & ~n11668;
  assign n11670 = ~po43  & n11668;
  assign n11671 = ~n11206 & ~n11207;
  assign n11672 = po14  & n11671;
  assign n11673 = ~n11212 & ~n11672;
  assign n11674 = n11212 & n11672;
  assign n11675 = ~n11673 & ~n11674;
  assign n11676 = ~n11670 & ~n11675;
  assign n11677 = ~n11669 & ~n11676;
  assign n11678 = po44  & ~n11677;
  assign n11679 = ~po44  & n11677;
  assign n11680 = ~n11215 & ~n11216;
  assign n11681 = po14  & n11680;
  assign n11682 = ~n11221 & ~n11681;
  assign n11683 = n11221 & n11681;
  assign n11684 = ~n11682 & ~n11683;
  assign n11685 = ~n11679 & ~n11684;
  assign n11686 = ~n11678 & ~n11685;
  assign n11687 = po45  & ~n11686;
  assign n11688 = ~po45  & n11686;
  assign n11689 = ~n11224 & ~n11225;
  assign n11690 = po14  & n11689;
  assign n11691 = ~n11230 & ~n11690;
  assign n11692 = n11230 & n11690;
  assign n11693 = ~n11691 & ~n11692;
  assign n11694 = ~n11688 & ~n11693;
  assign n11695 = ~n11687 & ~n11694;
  assign n11696 = po46  & ~n11695;
  assign n11697 = ~po46  & n11695;
  assign n11698 = ~n11233 & ~n11234;
  assign n11699 = po14  & n11698;
  assign n11700 = ~n11239 & ~n11699;
  assign n11701 = n11239 & n11699;
  assign n11702 = ~n11700 & ~n11701;
  assign n11703 = ~n11697 & ~n11702;
  assign n11704 = ~n11696 & ~n11703;
  assign n11705 = po47  & ~n11704;
  assign n11706 = ~po47  & n11704;
  assign n11707 = ~n11242 & ~n11243;
  assign n11708 = po14  & n11707;
  assign n11709 = ~n11248 & ~n11708;
  assign n11710 = n11248 & n11708;
  assign n11711 = ~n11709 & ~n11710;
  assign n11712 = ~n11706 & ~n11711;
  assign n11713 = ~n11705 & ~n11712;
  assign n11714 = po48  & ~n11713;
  assign n11715 = ~po48  & n11713;
  assign n11716 = ~n11251 & ~n11252;
  assign n11717 = po14  & n11716;
  assign n11718 = ~n11257 & ~n11717;
  assign n11719 = n11257 & n11717;
  assign n11720 = ~n11718 & ~n11719;
  assign n11721 = ~n11715 & ~n11720;
  assign n11722 = ~n11714 & ~n11721;
  assign n11723 = po49  & ~n11722;
  assign n11724 = ~po49  & n11722;
  assign n11725 = ~n11260 & ~n11261;
  assign n11726 = po14  & n11725;
  assign n11727 = ~n11266 & ~n11726;
  assign n11728 = n11266 & n11726;
  assign n11729 = ~n11727 & ~n11728;
  assign n11730 = ~n11724 & ~n11729;
  assign n11731 = ~n11723 & ~n11730;
  assign n11732 = po50  & ~n11731;
  assign n11733 = ~n11269 & ~n11275;
  assign n11734 = po14  & n11733;
  assign n11735 = ~n11274 & ~n11734;
  assign n11736 = n11274 & n11734;
  assign n11737 = ~n11735 & ~n11736;
  assign n11738 = ~po50  & n11731;
  assign n11739 = ~n11737 & ~n11738;
  assign n11740 = ~n11732 & ~n11739;
  assign n11741 = po51  & ~n11740;
  assign n11742 = ~po51  & n11740;
  assign n11743 = ~n11403 & ~n11742;
  assign n11744 = ~n11741 & ~n11743;
  assign n11745 = po52  & ~n11744;
  assign n11746 = ~po52  & n11744;
  assign n11747 = ~n11282 & ~n11283;
  assign n11748 = po14  & n11747;
  assign n11749 = ~n11288 & ~n11748;
  assign n11750 = n11288 & n11748;
  assign n11751 = ~n11749 & ~n11750;
  assign n11752 = ~n11746 & ~n11751;
  assign n11753 = ~n11745 & ~n11752;
  assign n11754 = po53  & ~n11753;
  assign n11755 = ~po53  & n11753;
  assign n11756 = ~n11291 & ~n11292;
  assign n11757 = po14  & n11756;
  assign n11758 = ~n11297 & ~n11757;
  assign n11759 = n11297 & n11757;
  assign n11760 = ~n11758 & ~n11759;
  assign n11761 = ~n11755 & ~n11760;
  assign n11762 = ~n11754 & ~n11761;
  assign n11763 = po54  & ~n11762;
  assign n11764 = ~po54  & n11762;
  assign n11765 = ~n11300 & ~n11301;
  assign n11766 = po14  & n11765;
  assign n11767 = ~n11306 & ~n11766;
  assign n11768 = n11306 & n11766;
  assign n11769 = ~n11767 & ~n11768;
  assign n11770 = ~n11764 & ~n11769;
  assign n11771 = ~n11763 & ~n11770;
  assign n11772 = po55  & ~n11771;
  assign n11773 = ~po55  & n11771;
  assign n11774 = ~n11309 & ~n11310;
  assign n11775 = po14  & n11774;
  assign n11776 = ~n11315 & ~n11775;
  assign n11777 = n11315 & n11775;
  assign n11778 = ~n11776 & ~n11777;
  assign n11779 = ~n11773 & ~n11778;
  assign n11780 = ~n11772 & ~n11779;
  assign n11781 = po56  & ~n11780;
  assign n11782 = ~po56  & n11780;
  assign n11783 = ~n11318 & ~n11319;
  assign n11784 = po14  & n11783;
  assign n11785 = ~n11324 & ~n11784;
  assign n11786 = n11324 & n11784;
  assign n11787 = ~n11785 & ~n11786;
  assign n11788 = ~n11782 & ~n11787;
  assign n11789 = ~n11781 & ~n11788;
  assign n11790 = po57  & ~n11789;
  assign n11791 = ~po57  & n11789;
  assign n11792 = ~n11327 & ~n11328;
  assign n11793 = po14  & n11792;
  assign n11794 = ~n11333 & ~n11793;
  assign n11795 = n11333 & n11793;
  assign n11796 = ~n11794 & ~n11795;
  assign n11797 = ~n11791 & ~n11796;
  assign n11798 = ~n11790 & ~n11797;
  assign n11799 = po58  & ~n11798;
  assign n11800 = ~po58  & n11798;
  assign n11801 = ~n11336 & ~n11337;
  assign n11802 = po14  & n11801;
  assign n11803 = ~n11342 & ~n11802;
  assign n11804 = n11342 & n11802;
  assign n11805 = ~n11803 & ~n11804;
  assign n11806 = ~n11800 & ~n11805;
  assign n11807 = ~n11799 & ~n11806;
  assign n11808 = po59  & ~n11807;
  assign n11809 = ~po59  & n11807;
  assign n11810 = ~n11345 & ~n11346;
  assign n11811 = po14  & n11810;
  assign n11812 = ~n11351 & ~n11811;
  assign n11813 = n11351 & n11811;
  assign n11814 = ~n11812 & ~n11813;
  assign n11815 = ~n11809 & ~n11814;
  assign n11816 = ~n11808 & ~n11815;
  assign n11817 = po60  & ~n11816;
  assign n11818 = ~po60  & n11816;
  assign n11819 = ~n11354 & ~n11355;
  assign n11820 = po14  & n11819;
  assign n11821 = ~n11360 & ~n11820;
  assign n11822 = n11360 & n11820;
  assign n11823 = ~n11821 & ~n11822;
  assign n11824 = ~n11818 & ~n11823;
  assign n11825 = ~n11817 & ~n11824;
  assign n11826 = po61  & ~n11825;
  assign n11827 = ~po61  & n11825;
  assign n11828 = ~n11363 & ~n11364;
  assign n11829 = po14  & n11828;
  assign n11830 = ~n11369 & ~n11829;
  assign n11831 = n11369 & n11829;
  assign n11832 = ~n11830 & ~n11831;
  assign n11833 = ~n11827 & ~n11832;
  assign n11834 = ~n11826 & ~n11833;
  assign n11835 = po62  & ~n11834;
  assign n11836 = ~po62  & n11834;
  assign n11837 = ~n11372 & ~n11373;
  assign n11838 = po14  & n11837;
  assign n11839 = ~n11378 & ~n11838;
  assign n11840 = n11378 & n11838;
  assign n11841 = ~n11839 & ~n11840;
  assign n11842 = ~n11836 & ~n11841;
  assign n11843 = ~n11835 & ~n11842;
  assign n11844 = n11413 & n11843;
  assign n11845 = ~n11413 & ~n11843;
  assign n11846 = n11391 & po14 ;
  assign n11847 = ~n11390 & ~n11846;
  assign n11848 = n11845 & n11847;
  assign n11849 = ~po63  & ~n11848;
  assign n11850 = ~n11844 & ~n11849;
  assign n11851 = ~n11408 & n11850;
  assign po13  = n11404 | ~n11851;
  assign n11853 = ~n11741 & ~n11742;
  assign n11854 = po13  & n11853;
  assign n11855 = ~n11403 & ~n11854;
  assign n11856 = n11403 & n11854;
  assign n11857 = ~n11855 & ~n11856;
  assign n11858 = n11413 & ~po13 ;
  assign n11859 = ~n11413 & po13 ;
  assign n11860 = n11843 & ~n11859;
  assign n11861 = po63  & ~n11860;
  assign n11862 = ~n11845 & n11861;
  assign n11863 = ~n11835 & ~n11836;
  assign n11864 = po13  & n11863;
  assign n11865 = ~n11841 & ~n11864;
  assign n11866 = n11841 & n11864;
  assign n11867 = ~n11865 & ~n11866;
  assign n11868 = pi26  & po13 ;
  assign n11869 = ~pi24  & ~pi25 ;
  assign n11870 = ~pi26  & n11869;
  assign n11871 = ~n11868 & ~n11870;
  assign n11872 = po14  & ~n11871;
  assign n11873 = ~po14  & n11871;
  assign n11874 = ~pi26  & po13 ;
  assign n11875 = pi27  & ~n11874;
  assign n11876 = n11415 & po13 ;
  assign n11877 = ~n11875 & ~n11876;
  assign n11878 = ~n11873 & n11877;
  assign n11879 = ~n11872 & ~n11878;
  assign n11880 = po15  & ~n11879;
  assign n11881 = ~po15  & n11879;
  assign n11882 = po14  & n11851;
  assign n11883 = ~n11876 & ~n11882;
  assign n11884 = pi28  & ~n11883;
  assign n11885 = ~pi28  & n11883;
  assign n11886 = ~n11884 & ~n11885;
  assign n11887 = ~n11881 & ~n11886;
  assign n11888 = ~n11880 & ~n11887;
  assign n11889 = po16  & ~n11888;
  assign n11890 = ~po16  & n11888;
  assign n11891 = ~n11418 & ~n11419;
  assign n11892 = po13  & n11891;
  assign n11893 = n11423 & ~n11892;
  assign n11894 = ~n11423 & n11892;
  assign n11895 = ~n11893 & ~n11894;
  assign n11896 = ~n11890 & ~n11895;
  assign n11897 = ~n11889 & ~n11896;
  assign n11898 = po17  & ~n11897;
  assign n11899 = ~po17  & n11897;
  assign n11900 = ~n11426 & ~n11427;
  assign n11901 = po13  & n11900;
  assign n11902 = ~n11432 & ~n11901;
  assign n11903 = n11432 & n11901;
  assign n11904 = ~n11902 & ~n11903;
  assign n11905 = ~n11899 & ~n11904;
  assign n11906 = ~n11898 & ~n11905;
  assign n11907 = po18  & ~n11906;
  assign n11908 = ~po18  & n11906;
  assign n11909 = ~n11435 & ~n11436;
  assign n11910 = po13  & n11909;
  assign n11911 = n11441 & n11910;
  assign n11912 = ~n11441 & ~n11910;
  assign n11913 = ~n11911 & ~n11912;
  assign n11914 = ~n11908 & ~n11913;
  assign n11915 = ~n11907 & ~n11914;
  assign n11916 = po19  & ~n11915;
  assign n11917 = ~po19  & n11915;
  assign n11918 = ~n11444 & ~n11445;
  assign n11919 = po13  & n11918;
  assign n11920 = ~n11450 & ~n11919;
  assign n11921 = n11450 & n11919;
  assign n11922 = ~n11920 & ~n11921;
  assign n11923 = ~n11917 & ~n11922;
  assign n11924 = ~n11916 & ~n11923;
  assign n11925 = po20  & ~n11924;
  assign n11926 = ~po20  & n11924;
  assign n11927 = ~n11453 & ~n11454;
  assign n11928 = po13  & n11927;
  assign n11929 = ~n11459 & ~n11928;
  assign n11930 = n11459 & n11928;
  assign n11931 = ~n11929 & ~n11930;
  assign n11932 = ~n11926 & ~n11931;
  assign n11933 = ~n11925 & ~n11932;
  assign n11934 = po21  & ~n11933;
  assign n11935 = ~po21  & n11933;
  assign n11936 = ~n11462 & ~n11463;
  assign n11937 = po13  & n11936;
  assign n11938 = ~n11468 & ~n11937;
  assign n11939 = n11468 & n11937;
  assign n11940 = ~n11938 & ~n11939;
  assign n11941 = ~n11935 & ~n11940;
  assign n11942 = ~n11934 & ~n11941;
  assign n11943 = po22  & ~n11942;
  assign n11944 = ~po22  & n11942;
  assign n11945 = ~n11471 & ~n11472;
  assign n11946 = po13  & n11945;
  assign n11947 = ~n11477 & ~n11946;
  assign n11948 = n11477 & n11946;
  assign n11949 = ~n11947 & ~n11948;
  assign n11950 = ~n11944 & ~n11949;
  assign n11951 = ~n11943 & ~n11950;
  assign n11952 = po23  & ~n11951;
  assign n11953 = ~po23  & n11951;
  assign n11954 = ~n11480 & ~n11481;
  assign n11955 = po13  & n11954;
  assign n11956 = ~n11486 & ~n11955;
  assign n11957 = n11486 & n11955;
  assign n11958 = ~n11956 & ~n11957;
  assign n11959 = ~n11953 & ~n11958;
  assign n11960 = ~n11952 & ~n11959;
  assign n11961 = po24  & ~n11960;
  assign n11962 = ~po24  & n11960;
  assign n11963 = ~n11489 & ~n11490;
  assign n11964 = po13  & n11963;
  assign n11965 = ~n11495 & ~n11964;
  assign n11966 = n11495 & n11964;
  assign n11967 = ~n11965 & ~n11966;
  assign n11968 = ~n11962 & ~n11967;
  assign n11969 = ~n11961 & ~n11968;
  assign n11970 = po25  & ~n11969;
  assign n11971 = ~po25  & n11969;
  assign n11972 = ~n11498 & ~n11499;
  assign n11973 = po13  & n11972;
  assign n11974 = ~n11504 & ~n11973;
  assign n11975 = n11504 & n11973;
  assign n11976 = ~n11974 & ~n11975;
  assign n11977 = ~n11971 & ~n11976;
  assign n11978 = ~n11970 & ~n11977;
  assign n11979 = po26  & ~n11978;
  assign n11980 = ~po26  & n11978;
  assign n11981 = ~n11507 & ~n11508;
  assign n11982 = po13  & n11981;
  assign n11983 = ~n11513 & ~n11982;
  assign n11984 = n11513 & n11982;
  assign n11985 = ~n11983 & ~n11984;
  assign n11986 = ~n11980 & ~n11985;
  assign n11987 = ~n11979 & ~n11986;
  assign n11988 = po27  & ~n11987;
  assign n11989 = ~po27  & n11987;
  assign n11990 = ~n11516 & ~n11517;
  assign n11991 = po13  & n11990;
  assign n11992 = ~n11522 & ~n11991;
  assign n11993 = n11522 & n11991;
  assign n11994 = ~n11992 & ~n11993;
  assign n11995 = ~n11989 & ~n11994;
  assign n11996 = ~n11988 & ~n11995;
  assign n11997 = po28  & ~n11996;
  assign n11998 = ~po28  & n11996;
  assign n11999 = ~n11525 & ~n11526;
  assign n12000 = po13  & n11999;
  assign n12001 = ~n11531 & ~n12000;
  assign n12002 = n11531 & n12000;
  assign n12003 = ~n12001 & ~n12002;
  assign n12004 = ~n11998 & ~n12003;
  assign n12005 = ~n11997 & ~n12004;
  assign n12006 = po29  & ~n12005;
  assign n12007 = ~po29  & n12005;
  assign n12008 = ~n11534 & ~n11535;
  assign n12009 = po13  & n12008;
  assign n12010 = ~n11540 & ~n12009;
  assign n12011 = n11540 & n12009;
  assign n12012 = ~n12010 & ~n12011;
  assign n12013 = ~n12007 & ~n12012;
  assign n12014 = ~n12006 & ~n12013;
  assign n12015 = po30  & ~n12014;
  assign n12016 = ~po30  & n12014;
  assign n12017 = ~n11543 & ~n11544;
  assign n12018 = po13  & n12017;
  assign n12019 = ~n11549 & ~n12018;
  assign n12020 = n11549 & n12018;
  assign n12021 = ~n12019 & ~n12020;
  assign n12022 = ~n12016 & ~n12021;
  assign n12023 = ~n12015 & ~n12022;
  assign n12024 = po31  & ~n12023;
  assign n12025 = ~po31  & n12023;
  assign n12026 = ~n11552 & ~n11553;
  assign n12027 = po13  & n12026;
  assign n12028 = ~n11558 & ~n12027;
  assign n12029 = n11558 & n12027;
  assign n12030 = ~n12028 & ~n12029;
  assign n12031 = ~n12025 & ~n12030;
  assign n12032 = ~n12024 & ~n12031;
  assign n12033 = po32  & ~n12032;
  assign n12034 = ~po32  & n12032;
  assign n12035 = ~n11561 & ~n11562;
  assign n12036 = po13  & n12035;
  assign n12037 = ~n11567 & ~n12036;
  assign n12038 = n11567 & n12036;
  assign n12039 = ~n12037 & ~n12038;
  assign n12040 = ~n12034 & ~n12039;
  assign n12041 = ~n12033 & ~n12040;
  assign n12042 = po33  & ~n12041;
  assign n12043 = ~po33  & n12041;
  assign n12044 = ~n11570 & ~n11571;
  assign n12045 = po13  & n12044;
  assign n12046 = ~n11576 & ~n12045;
  assign n12047 = n11576 & n12045;
  assign n12048 = ~n12046 & ~n12047;
  assign n12049 = ~n12043 & ~n12048;
  assign n12050 = ~n12042 & ~n12049;
  assign n12051 = po34  & ~n12050;
  assign n12052 = ~po34  & n12050;
  assign n12053 = ~n11579 & ~n11580;
  assign n12054 = po13  & n12053;
  assign n12055 = ~n11585 & ~n12054;
  assign n12056 = n11585 & n12054;
  assign n12057 = ~n12055 & ~n12056;
  assign n12058 = ~n12052 & ~n12057;
  assign n12059 = ~n12051 & ~n12058;
  assign n12060 = po35  & ~n12059;
  assign n12061 = ~po35  & n12059;
  assign n12062 = ~n11588 & ~n11589;
  assign n12063 = po13  & n12062;
  assign n12064 = ~n11594 & ~n12063;
  assign n12065 = n11594 & n12063;
  assign n12066 = ~n12064 & ~n12065;
  assign n12067 = ~n12061 & ~n12066;
  assign n12068 = ~n12060 & ~n12067;
  assign n12069 = po36  & ~n12068;
  assign n12070 = ~po36  & n12068;
  assign n12071 = ~n11597 & ~n11598;
  assign n12072 = po13  & n12071;
  assign n12073 = ~n11603 & ~n12072;
  assign n12074 = n11603 & n12072;
  assign n12075 = ~n12073 & ~n12074;
  assign n12076 = ~n12070 & ~n12075;
  assign n12077 = ~n12069 & ~n12076;
  assign n12078 = po37  & ~n12077;
  assign n12079 = ~po37  & n12077;
  assign n12080 = ~n11606 & ~n11607;
  assign n12081 = po13  & n12080;
  assign n12082 = ~n11612 & ~n12081;
  assign n12083 = n11612 & n12081;
  assign n12084 = ~n12082 & ~n12083;
  assign n12085 = ~n12079 & ~n12084;
  assign n12086 = ~n12078 & ~n12085;
  assign n12087 = po38  & ~n12086;
  assign n12088 = ~po38  & n12086;
  assign n12089 = ~n11615 & ~n11616;
  assign n12090 = po13  & n12089;
  assign n12091 = ~n11621 & ~n12090;
  assign n12092 = n11621 & n12090;
  assign n12093 = ~n12091 & ~n12092;
  assign n12094 = ~n12088 & ~n12093;
  assign n12095 = ~n12087 & ~n12094;
  assign n12096 = po39  & ~n12095;
  assign n12097 = ~po39  & n12095;
  assign n12098 = ~n11624 & ~n11625;
  assign n12099 = po13  & n12098;
  assign n12100 = ~n11630 & ~n12099;
  assign n12101 = n11630 & n12099;
  assign n12102 = ~n12100 & ~n12101;
  assign n12103 = ~n12097 & ~n12102;
  assign n12104 = ~n12096 & ~n12103;
  assign n12105 = po40  & ~n12104;
  assign n12106 = ~po40  & n12104;
  assign n12107 = ~n11633 & ~n11634;
  assign n12108 = po13  & n12107;
  assign n12109 = ~n11639 & ~n12108;
  assign n12110 = n11639 & n12108;
  assign n12111 = ~n12109 & ~n12110;
  assign n12112 = ~n12106 & ~n12111;
  assign n12113 = ~n12105 & ~n12112;
  assign n12114 = po41  & ~n12113;
  assign n12115 = ~po41  & n12113;
  assign n12116 = ~n11642 & ~n11643;
  assign n12117 = po13  & n12116;
  assign n12118 = ~n11648 & ~n12117;
  assign n12119 = n11648 & n12117;
  assign n12120 = ~n12118 & ~n12119;
  assign n12121 = ~n12115 & ~n12120;
  assign n12122 = ~n12114 & ~n12121;
  assign n12123 = po42  & ~n12122;
  assign n12124 = ~po42  & n12122;
  assign n12125 = ~n11651 & ~n11652;
  assign n12126 = po13  & n12125;
  assign n12127 = ~n11657 & ~n12126;
  assign n12128 = n11657 & n12126;
  assign n12129 = ~n12127 & ~n12128;
  assign n12130 = ~n12124 & ~n12129;
  assign n12131 = ~n12123 & ~n12130;
  assign n12132 = po43  & ~n12131;
  assign n12133 = ~po43  & n12131;
  assign n12134 = ~n11660 & ~n11661;
  assign n12135 = po13  & n12134;
  assign n12136 = ~n11666 & ~n12135;
  assign n12137 = n11666 & n12135;
  assign n12138 = ~n12136 & ~n12137;
  assign n12139 = ~n12133 & ~n12138;
  assign n12140 = ~n12132 & ~n12139;
  assign n12141 = po44  & ~n12140;
  assign n12142 = ~po44  & n12140;
  assign n12143 = ~n11669 & ~n11670;
  assign n12144 = po13  & n12143;
  assign n12145 = ~n11675 & ~n12144;
  assign n12146 = n11675 & n12144;
  assign n12147 = ~n12145 & ~n12146;
  assign n12148 = ~n12142 & ~n12147;
  assign n12149 = ~n12141 & ~n12148;
  assign n12150 = po45  & ~n12149;
  assign n12151 = ~po45  & n12149;
  assign n12152 = ~n11678 & ~n11679;
  assign n12153 = po13  & n12152;
  assign n12154 = ~n11684 & ~n12153;
  assign n12155 = n11684 & n12153;
  assign n12156 = ~n12154 & ~n12155;
  assign n12157 = ~n12151 & ~n12156;
  assign n12158 = ~n12150 & ~n12157;
  assign n12159 = po46  & ~n12158;
  assign n12160 = ~po46  & n12158;
  assign n12161 = ~n11687 & ~n11688;
  assign n12162 = po13  & n12161;
  assign n12163 = ~n11693 & ~n12162;
  assign n12164 = n11693 & n12162;
  assign n12165 = ~n12163 & ~n12164;
  assign n12166 = ~n12160 & ~n12165;
  assign n12167 = ~n12159 & ~n12166;
  assign n12168 = po47  & ~n12167;
  assign n12169 = ~po47  & n12167;
  assign n12170 = ~n11696 & ~n11697;
  assign n12171 = po13  & n12170;
  assign n12172 = ~n11702 & ~n12171;
  assign n12173 = n11702 & n12171;
  assign n12174 = ~n12172 & ~n12173;
  assign n12175 = ~n12169 & ~n12174;
  assign n12176 = ~n12168 & ~n12175;
  assign n12177 = po48  & ~n12176;
  assign n12178 = ~po48  & n12176;
  assign n12179 = ~n11705 & ~n11706;
  assign n12180 = po13  & n12179;
  assign n12181 = ~n11711 & ~n12180;
  assign n12182 = n11711 & n12180;
  assign n12183 = ~n12181 & ~n12182;
  assign n12184 = ~n12178 & ~n12183;
  assign n12185 = ~n12177 & ~n12184;
  assign n12186 = po49  & ~n12185;
  assign n12187 = ~po49  & n12185;
  assign n12188 = ~n11714 & ~n11715;
  assign n12189 = po13  & n12188;
  assign n12190 = ~n11720 & ~n12189;
  assign n12191 = n11720 & n12189;
  assign n12192 = ~n12190 & ~n12191;
  assign n12193 = ~n12187 & ~n12192;
  assign n12194 = ~n12186 & ~n12193;
  assign n12195 = po50  & ~n12194;
  assign n12196 = ~po50  & n12194;
  assign n12197 = ~n11723 & ~n11724;
  assign n12198 = po13  & n12197;
  assign n12199 = ~n11729 & ~n12198;
  assign n12200 = n11729 & n12198;
  assign n12201 = ~n12199 & ~n12200;
  assign n12202 = ~n12196 & ~n12201;
  assign n12203 = ~n12195 & ~n12202;
  assign n12204 = po51  & ~n12203;
  assign n12205 = ~n11732 & ~n11738;
  assign n12206 = po13  & n12205;
  assign n12207 = ~n11737 & ~n12206;
  assign n12208 = n11737 & n12206;
  assign n12209 = ~n12207 & ~n12208;
  assign n12210 = ~po51  & n12203;
  assign n12211 = ~n12209 & ~n12210;
  assign n12212 = ~n12204 & ~n12211;
  assign n12213 = po52  & ~n12212;
  assign n12214 = ~po52  & n12212;
  assign n12215 = ~n11857 & ~n12214;
  assign n12216 = ~n12213 & ~n12215;
  assign n12217 = po53  & ~n12216;
  assign n12218 = ~po53  & n12216;
  assign n12219 = ~n11745 & ~n11746;
  assign n12220 = po13  & n12219;
  assign n12221 = ~n11751 & ~n12220;
  assign n12222 = n11751 & n12220;
  assign n12223 = ~n12221 & ~n12222;
  assign n12224 = ~n12218 & ~n12223;
  assign n12225 = ~n12217 & ~n12224;
  assign n12226 = po54  & ~n12225;
  assign n12227 = ~po54  & n12225;
  assign n12228 = ~n11754 & ~n11755;
  assign n12229 = po13  & n12228;
  assign n12230 = ~n11760 & ~n12229;
  assign n12231 = n11760 & n12229;
  assign n12232 = ~n12230 & ~n12231;
  assign n12233 = ~n12227 & ~n12232;
  assign n12234 = ~n12226 & ~n12233;
  assign n12235 = po55  & ~n12234;
  assign n12236 = ~po55  & n12234;
  assign n12237 = ~n11763 & ~n11764;
  assign n12238 = po13  & n12237;
  assign n12239 = ~n11769 & ~n12238;
  assign n12240 = n11769 & n12238;
  assign n12241 = ~n12239 & ~n12240;
  assign n12242 = ~n12236 & ~n12241;
  assign n12243 = ~n12235 & ~n12242;
  assign n12244 = po56  & ~n12243;
  assign n12245 = ~po56  & n12243;
  assign n12246 = ~n11772 & ~n11773;
  assign n12247 = po13  & n12246;
  assign n12248 = ~n11778 & ~n12247;
  assign n12249 = n11778 & n12247;
  assign n12250 = ~n12248 & ~n12249;
  assign n12251 = ~n12245 & ~n12250;
  assign n12252 = ~n12244 & ~n12251;
  assign n12253 = po57  & ~n12252;
  assign n12254 = ~po57  & n12252;
  assign n12255 = ~n11781 & ~n11782;
  assign n12256 = po13  & n12255;
  assign n12257 = ~n11787 & ~n12256;
  assign n12258 = n11787 & n12256;
  assign n12259 = ~n12257 & ~n12258;
  assign n12260 = ~n12254 & ~n12259;
  assign n12261 = ~n12253 & ~n12260;
  assign n12262 = po58  & ~n12261;
  assign n12263 = ~po58  & n12261;
  assign n12264 = ~n11790 & ~n11791;
  assign n12265 = po13  & n12264;
  assign n12266 = ~n11796 & ~n12265;
  assign n12267 = n11796 & n12265;
  assign n12268 = ~n12266 & ~n12267;
  assign n12269 = ~n12263 & ~n12268;
  assign n12270 = ~n12262 & ~n12269;
  assign n12271 = po59  & ~n12270;
  assign n12272 = ~po59  & n12270;
  assign n12273 = ~n11799 & ~n11800;
  assign n12274 = po13  & n12273;
  assign n12275 = ~n11805 & ~n12274;
  assign n12276 = n11805 & n12274;
  assign n12277 = ~n12275 & ~n12276;
  assign n12278 = ~n12272 & ~n12277;
  assign n12279 = ~n12271 & ~n12278;
  assign n12280 = po60  & ~n12279;
  assign n12281 = ~po60  & n12279;
  assign n12282 = ~n11808 & ~n11809;
  assign n12283 = po13  & n12282;
  assign n12284 = ~n11814 & ~n12283;
  assign n12285 = n11814 & n12283;
  assign n12286 = ~n12284 & ~n12285;
  assign n12287 = ~n12281 & ~n12286;
  assign n12288 = ~n12280 & ~n12287;
  assign n12289 = po61  & ~n12288;
  assign n12290 = ~po61  & n12288;
  assign n12291 = ~n11817 & ~n11818;
  assign n12292 = po13  & n12291;
  assign n12293 = ~n11823 & ~n12292;
  assign n12294 = n11823 & n12292;
  assign n12295 = ~n12293 & ~n12294;
  assign n12296 = ~n12290 & ~n12295;
  assign n12297 = ~n12289 & ~n12296;
  assign n12298 = po62  & ~n12297;
  assign n12299 = ~po62  & n12297;
  assign n12300 = ~n11826 & ~n11827;
  assign n12301 = po13  & n12300;
  assign n12302 = ~n11832 & ~n12301;
  assign n12303 = n11832 & n12301;
  assign n12304 = ~n12302 & ~n12303;
  assign n12305 = ~n12299 & ~n12304;
  assign n12306 = ~n12298 & ~n12305;
  assign n12307 = n11867 & n12306;
  assign n12308 = ~n11867 & ~n12306;
  assign n12309 = n11845 & po13 ;
  assign n12310 = ~n11844 & ~n12309;
  assign n12311 = n12308 & n12310;
  assign n12312 = ~po63  & ~n12311;
  assign n12313 = ~n12307 & ~n12312;
  assign n12314 = ~n11862 & n12313;
  assign po12  = n11858 | ~n12314;
  assign n12316 = ~n12213 & ~n12214;
  assign n12317 = po12  & n12316;
  assign n12318 = ~n11857 & ~n12317;
  assign n12319 = n11857 & n12317;
  assign n12320 = ~n12318 & ~n12319;
  assign n12321 = n11867 & ~po12 ;
  assign n12322 = ~n11867 & po12 ;
  assign n12323 = n12306 & ~n12322;
  assign n12324 = po63  & ~n12323;
  assign n12325 = ~n12308 & n12324;
  assign n12326 = ~n12298 & ~n12299;
  assign n12327 = po12  & n12326;
  assign n12328 = ~n12304 & ~n12327;
  assign n12329 = n12304 & n12327;
  assign n12330 = ~n12328 & ~n12329;
  assign n12331 = pi24  & po12 ;
  assign n12332 = ~pi22  & ~pi23 ;
  assign n12333 = ~pi24  & n12332;
  assign n12334 = ~n12331 & ~n12333;
  assign n12335 = po13  & ~n12334;
  assign n12336 = ~po13  & n12334;
  assign n12337 = ~pi24  & po12 ;
  assign n12338 = pi25  & ~n12337;
  assign n12339 = n11869 & po12 ;
  assign n12340 = ~n12338 & ~n12339;
  assign n12341 = ~n12336 & n12340;
  assign n12342 = ~n12335 & ~n12341;
  assign n12343 = po14  & ~n12342;
  assign n12344 = ~po14  & n12342;
  assign n12345 = po13  & n12314;
  assign n12346 = ~n12339 & ~n12345;
  assign n12347 = pi26  & ~n12346;
  assign n12348 = ~pi26  & n12346;
  assign n12349 = ~n12347 & ~n12348;
  assign n12350 = ~n12344 & ~n12349;
  assign n12351 = ~n12343 & ~n12350;
  assign n12352 = po15  & ~n12351;
  assign n12353 = ~po15  & n12351;
  assign n12354 = ~n11872 & ~n11873;
  assign n12355 = po12  & n12354;
  assign n12356 = n11877 & ~n12355;
  assign n12357 = ~n11877 & n12355;
  assign n12358 = ~n12356 & ~n12357;
  assign n12359 = ~n12353 & ~n12358;
  assign n12360 = ~n12352 & ~n12359;
  assign n12361 = po16  & ~n12360;
  assign n12362 = ~po16  & n12360;
  assign n12363 = ~n11880 & ~n11881;
  assign n12364 = po12  & n12363;
  assign n12365 = ~n11886 & ~n12364;
  assign n12366 = n11886 & n12364;
  assign n12367 = ~n12365 & ~n12366;
  assign n12368 = ~n12362 & ~n12367;
  assign n12369 = ~n12361 & ~n12368;
  assign n12370 = po17  & ~n12369;
  assign n12371 = ~po17  & n12369;
  assign n12372 = ~n11889 & ~n11890;
  assign n12373 = po12  & n12372;
  assign n12374 = n11895 & n12373;
  assign n12375 = ~n11895 & ~n12373;
  assign n12376 = ~n12374 & ~n12375;
  assign n12377 = ~n12371 & ~n12376;
  assign n12378 = ~n12370 & ~n12377;
  assign n12379 = po18  & ~n12378;
  assign n12380 = ~po18  & n12378;
  assign n12381 = ~n11898 & ~n11899;
  assign n12382 = po12  & n12381;
  assign n12383 = ~n11904 & ~n12382;
  assign n12384 = n11904 & n12382;
  assign n12385 = ~n12383 & ~n12384;
  assign n12386 = ~n12380 & ~n12385;
  assign n12387 = ~n12379 & ~n12386;
  assign n12388 = po19  & ~n12387;
  assign n12389 = ~po19  & n12387;
  assign n12390 = ~n11907 & ~n11908;
  assign n12391 = po12  & n12390;
  assign n12392 = ~n11913 & ~n12391;
  assign n12393 = n11913 & n12391;
  assign n12394 = ~n12392 & ~n12393;
  assign n12395 = ~n12389 & ~n12394;
  assign n12396 = ~n12388 & ~n12395;
  assign n12397 = po20  & ~n12396;
  assign n12398 = ~po20  & n12396;
  assign n12399 = ~n11916 & ~n11917;
  assign n12400 = po12  & n12399;
  assign n12401 = ~n11922 & ~n12400;
  assign n12402 = n11922 & n12400;
  assign n12403 = ~n12401 & ~n12402;
  assign n12404 = ~n12398 & ~n12403;
  assign n12405 = ~n12397 & ~n12404;
  assign n12406 = po21  & ~n12405;
  assign n12407 = ~po21  & n12405;
  assign n12408 = ~n11925 & ~n11926;
  assign n12409 = po12  & n12408;
  assign n12410 = ~n11931 & ~n12409;
  assign n12411 = n11931 & n12409;
  assign n12412 = ~n12410 & ~n12411;
  assign n12413 = ~n12407 & ~n12412;
  assign n12414 = ~n12406 & ~n12413;
  assign n12415 = po22  & ~n12414;
  assign n12416 = ~po22  & n12414;
  assign n12417 = ~n11934 & ~n11935;
  assign n12418 = po12  & n12417;
  assign n12419 = ~n11940 & ~n12418;
  assign n12420 = n11940 & n12418;
  assign n12421 = ~n12419 & ~n12420;
  assign n12422 = ~n12416 & ~n12421;
  assign n12423 = ~n12415 & ~n12422;
  assign n12424 = po23  & ~n12423;
  assign n12425 = ~po23  & n12423;
  assign n12426 = ~n11943 & ~n11944;
  assign n12427 = po12  & n12426;
  assign n12428 = ~n11949 & ~n12427;
  assign n12429 = n11949 & n12427;
  assign n12430 = ~n12428 & ~n12429;
  assign n12431 = ~n12425 & ~n12430;
  assign n12432 = ~n12424 & ~n12431;
  assign n12433 = po24  & ~n12432;
  assign n12434 = ~po24  & n12432;
  assign n12435 = ~n11952 & ~n11953;
  assign n12436 = po12  & n12435;
  assign n12437 = ~n11958 & ~n12436;
  assign n12438 = n11958 & n12436;
  assign n12439 = ~n12437 & ~n12438;
  assign n12440 = ~n12434 & ~n12439;
  assign n12441 = ~n12433 & ~n12440;
  assign n12442 = po25  & ~n12441;
  assign n12443 = ~po25  & n12441;
  assign n12444 = ~n11961 & ~n11962;
  assign n12445 = po12  & n12444;
  assign n12446 = ~n11967 & ~n12445;
  assign n12447 = n11967 & n12445;
  assign n12448 = ~n12446 & ~n12447;
  assign n12449 = ~n12443 & ~n12448;
  assign n12450 = ~n12442 & ~n12449;
  assign n12451 = po26  & ~n12450;
  assign n12452 = ~po26  & n12450;
  assign n12453 = ~n11970 & ~n11971;
  assign n12454 = po12  & n12453;
  assign n12455 = ~n11976 & ~n12454;
  assign n12456 = n11976 & n12454;
  assign n12457 = ~n12455 & ~n12456;
  assign n12458 = ~n12452 & ~n12457;
  assign n12459 = ~n12451 & ~n12458;
  assign n12460 = po27  & ~n12459;
  assign n12461 = ~po27  & n12459;
  assign n12462 = ~n11979 & ~n11980;
  assign n12463 = po12  & n12462;
  assign n12464 = ~n11985 & ~n12463;
  assign n12465 = n11985 & n12463;
  assign n12466 = ~n12464 & ~n12465;
  assign n12467 = ~n12461 & ~n12466;
  assign n12468 = ~n12460 & ~n12467;
  assign n12469 = po28  & ~n12468;
  assign n12470 = ~po28  & n12468;
  assign n12471 = ~n11988 & ~n11989;
  assign n12472 = po12  & n12471;
  assign n12473 = ~n11994 & ~n12472;
  assign n12474 = n11994 & n12472;
  assign n12475 = ~n12473 & ~n12474;
  assign n12476 = ~n12470 & ~n12475;
  assign n12477 = ~n12469 & ~n12476;
  assign n12478 = po29  & ~n12477;
  assign n12479 = ~po29  & n12477;
  assign n12480 = ~n11997 & ~n11998;
  assign n12481 = po12  & n12480;
  assign n12482 = ~n12003 & ~n12481;
  assign n12483 = n12003 & n12481;
  assign n12484 = ~n12482 & ~n12483;
  assign n12485 = ~n12479 & ~n12484;
  assign n12486 = ~n12478 & ~n12485;
  assign n12487 = po30  & ~n12486;
  assign n12488 = ~po30  & n12486;
  assign n12489 = ~n12006 & ~n12007;
  assign n12490 = po12  & n12489;
  assign n12491 = ~n12012 & ~n12490;
  assign n12492 = n12012 & n12490;
  assign n12493 = ~n12491 & ~n12492;
  assign n12494 = ~n12488 & ~n12493;
  assign n12495 = ~n12487 & ~n12494;
  assign n12496 = po31  & ~n12495;
  assign n12497 = ~po31  & n12495;
  assign n12498 = ~n12015 & ~n12016;
  assign n12499 = po12  & n12498;
  assign n12500 = ~n12021 & ~n12499;
  assign n12501 = n12021 & n12499;
  assign n12502 = ~n12500 & ~n12501;
  assign n12503 = ~n12497 & ~n12502;
  assign n12504 = ~n12496 & ~n12503;
  assign n12505 = po32  & ~n12504;
  assign n12506 = ~po32  & n12504;
  assign n12507 = ~n12024 & ~n12025;
  assign n12508 = po12  & n12507;
  assign n12509 = ~n12030 & ~n12508;
  assign n12510 = n12030 & n12508;
  assign n12511 = ~n12509 & ~n12510;
  assign n12512 = ~n12506 & ~n12511;
  assign n12513 = ~n12505 & ~n12512;
  assign n12514 = po33  & ~n12513;
  assign n12515 = ~po33  & n12513;
  assign n12516 = ~n12033 & ~n12034;
  assign n12517 = po12  & n12516;
  assign n12518 = ~n12039 & ~n12517;
  assign n12519 = n12039 & n12517;
  assign n12520 = ~n12518 & ~n12519;
  assign n12521 = ~n12515 & ~n12520;
  assign n12522 = ~n12514 & ~n12521;
  assign n12523 = po34  & ~n12522;
  assign n12524 = ~po34  & n12522;
  assign n12525 = ~n12042 & ~n12043;
  assign n12526 = po12  & n12525;
  assign n12527 = ~n12048 & ~n12526;
  assign n12528 = n12048 & n12526;
  assign n12529 = ~n12527 & ~n12528;
  assign n12530 = ~n12524 & ~n12529;
  assign n12531 = ~n12523 & ~n12530;
  assign n12532 = po35  & ~n12531;
  assign n12533 = ~po35  & n12531;
  assign n12534 = ~n12051 & ~n12052;
  assign n12535 = po12  & n12534;
  assign n12536 = ~n12057 & ~n12535;
  assign n12537 = n12057 & n12535;
  assign n12538 = ~n12536 & ~n12537;
  assign n12539 = ~n12533 & ~n12538;
  assign n12540 = ~n12532 & ~n12539;
  assign n12541 = po36  & ~n12540;
  assign n12542 = ~po36  & n12540;
  assign n12543 = ~n12060 & ~n12061;
  assign n12544 = po12  & n12543;
  assign n12545 = ~n12066 & ~n12544;
  assign n12546 = n12066 & n12544;
  assign n12547 = ~n12545 & ~n12546;
  assign n12548 = ~n12542 & ~n12547;
  assign n12549 = ~n12541 & ~n12548;
  assign n12550 = po37  & ~n12549;
  assign n12551 = ~po37  & n12549;
  assign n12552 = ~n12069 & ~n12070;
  assign n12553 = po12  & n12552;
  assign n12554 = ~n12075 & ~n12553;
  assign n12555 = n12075 & n12553;
  assign n12556 = ~n12554 & ~n12555;
  assign n12557 = ~n12551 & ~n12556;
  assign n12558 = ~n12550 & ~n12557;
  assign n12559 = po38  & ~n12558;
  assign n12560 = ~po38  & n12558;
  assign n12561 = ~n12078 & ~n12079;
  assign n12562 = po12  & n12561;
  assign n12563 = ~n12084 & ~n12562;
  assign n12564 = n12084 & n12562;
  assign n12565 = ~n12563 & ~n12564;
  assign n12566 = ~n12560 & ~n12565;
  assign n12567 = ~n12559 & ~n12566;
  assign n12568 = po39  & ~n12567;
  assign n12569 = ~po39  & n12567;
  assign n12570 = ~n12087 & ~n12088;
  assign n12571 = po12  & n12570;
  assign n12572 = ~n12093 & ~n12571;
  assign n12573 = n12093 & n12571;
  assign n12574 = ~n12572 & ~n12573;
  assign n12575 = ~n12569 & ~n12574;
  assign n12576 = ~n12568 & ~n12575;
  assign n12577 = po40  & ~n12576;
  assign n12578 = ~po40  & n12576;
  assign n12579 = ~n12096 & ~n12097;
  assign n12580 = po12  & n12579;
  assign n12581 = ~n12102 & ~n12580;
  assign n12582 = n12102 & n12580;
  assign n12583 = ~n12581 & ~n12582;
  assign n12584 = ~n12578 & ~n12583;
  assign n12585 = ~n12577 & ~n12584;
  assign n12586 = po41  & ~n12585;
  assign n12587 = ~po41  & n12585;
  assign n12588 = ~n12105 & ~n12106;
  assign n12589 = po12  & n12588;
  assign n12590 = ~n12111 & ~n12589;
  assign n12591 = n12111 & n12589;
  assign n12592 = ~n12590 & ~n12591;
  assign n12593 = ~n12587 & ~n12592;
  assign n12594 = ~n12586 & ~n12593;
  assign n12595 = po42  & ~n12594;
  assign n12596 = ~po42  & n12594;
  assign n12597 = ~n12114 & ~n12115;
  assign n12598 = po12  & n12597;
  assign n12599 = ~n12120 & ~n12598;
  assign n12600 = n12120 & n12598;
  assign n12601 = ~n12599 & ~n12600;
  assign n12602 = ~n12596 & ~n12601;
  assign n12603 = ~n12595 & ~n12602;
  assign n12604 = po43  & ~n12603;
  assign n12605 = ~po43  & n12603;
  assign n12606 = ~n12123 & ~n12124;
  assign n12607 = po12  & n12606;
  assign n12608 = ~n12129 & ~n12607;
  assign n12609 = n12129 & n12607;
  assign n12610 = ~n12608 & ~n12609;
  assign n12611 = ~n12605 & ~n12610;
  assign n12612 = ~n12604 & ~n12611;
  assign n12613 = po44  & ~n12612;
  assign n12614 = ~po44  & n12612;
  assign n12615 = ~n12132 & ~n12133;
  assign n12616 = po12  & n12615;
  assign n12617 = ~n12138 & ~n12616;
  assign n12618 = n12138 & n12616;
  assign n12619 = ~n12617 & ~n12618;
  assign n12620 = ~n12614 & ~n12619;
  assign n12621 = ~n12613 & ~n12620;
  assign n12622 = po45  & ~n12621;
  assign n12623 = ~po45  & n12621;
  assign n12624 = ~n12141 & ~n12142;
  assign n12625 = po12  & n12624;
  assign n12626 = ~n12147 & ~n12625;
  assign n12627 = n12147 & n12625;
  assign n12628 = ~n12626 & ~n12627;
  assign n12629 = ~n12623 & ~n12628;
  assign n12630 = ~n12622 & ~n12629;
  assign n12631 = po46  & ~n12630;
  assign n12632 = ~po46  & n12630;
  assign n12633 = ~n12150 & ~n12151;
  assign n12634 = po12  & n12633;
  assign n12635 = ~n12156 & ~n12634;
  assign n12636 = n12156 & n12634;
  assign n12637 = ~n12635 & ~n12636;
  assign n12638 = ~n12632 & ~n12637;
  assign n12639 = ~n12631 & ~n12638;
  assign n12640 = po47  & ~n12639;
  assign n12641 = ~po47  & n12639;
  assign n12642 = ~n12159 & ~n12160;
  assign n12643 = po12  & n12642;
  assign n12644 = ~n12165 & ~n12643;
  assign n12645 = n12165 & n12643;
  assign n12646 = ~n12644 & ~n12645;
  assign n12647 = ~n12641 & ~n12646;
  assign n12648 = ~n12640 & ~n12647;
  assign n12649 = po48  & ~n12648;
  assign n12650 = ~po48  & n12648;
  assign n12651 = ~n12168 & ~n12169;
  assign n12652 = po12  & n12651;
  assign n12653 = ~n12174 & ~n12652;
  assign n12654 = n12174 & n12652;
  assign n12655 = ~n12653 & ~n12654;
  assign n12656 = ~n12650 & ~n12655;
  assign n12657 = ~n12649 & ~n12656;
  assign n12658 = po49  & ~n12657;
  assign n12659 = ~po49  & n12657;
  assign n12660 = ~n12177 & ~n12178;
  assign n12661 = po12  & n12660;
  assign n12662 = ~n12183 & ~n12661;
  assign n12663 = n12183 & n12661;
  assign n12664 = ~n12662 & ~n12663;
  assign n12665 = ~n12659 & ~n12664;
  assign n12666 = ~n12658 & ~n12665;
  assign n12667 = po50  & ~n12666;
  assign n12668 = ~po50  & n12666;
  assign n12669 = ~n12186 & ~n12187;
  assign n12670 = po12  & n12669;
  assign n12671 = ~n12192 & ~n12670;
  assign n12672 = n12192 & n12670;
  assign n12673 = ~n12671 & ~n12672;
  assign n12674 = ~n12668 & ~n12673;
  assign n12675 = ~n12667 & ~n12674;
  assign n12676 = po51  & ~n12675;
  assign n12677 = ~po51  & n12675;
  assign n12678 = ~n12195 & ~n12196;
  assign n12679 = po12  & n12678;
  assign n12680 = ~n12201 & ~n12679;
  assign n12681 = n12201 & n12679;
  assign n12682 = ~n12680 & ~n12681;
  assign n12683 = ~n12677 & ~n12682;
  assign n12684 = ~n12676 & ~n12683;
  assign n12685 = po52  & ~n12684;
  assign n12686 = ~n12204 & ~n12210;
  assign n12687 = po12  & n12686;
  assign n12688 = ~n12209 & ~n12687;
  assign n12689 = n12209 & n12687;
  assign n12690 = ~n12688 & ~n12689;
  assign n12691 = ~po52  & n12684;
  assign n12692 = ~n12690 & ~n12691;
  assign n12693 = ~n12685 & ~n12692;
  assign n12694 = po53  & ~n12693;
  assign n12695 = ~po53  & n12693;
  assign n12696 = ~n12320 & ~n12695;
  assign n12697 = ~n12694 & ~n12696;
  assign n12698 = po54  & ~n12697;
  assign n12699 = ~po54  & n12697;
  assign n12700 = ~n12217 & ~n12218;
  assign n12701 = po12  & n12700;
  assign n12702 = ~n12223 & ~n12701;
  assign n12703 = n12223 & n12701;
  assign n12704 = ~n12702 & ~n12703;
  assign n12705 = ~n12699 & ~n12704;
  assign n12706 = ~n12698 & ~n12705;
  assign n12707 = po55  & ~n12706;
  assign n12708 = ~po55  & n12706;
  assign n12709 = ~n12226 & ~n12227;
  assign n12710 = po12  & n12709;
  assign n12711 = ~n12232 & ~n12710;
  assign n12712 = n12232 & n12710;
  assign n12713 = ~n12711 & ~n12712;
  assign n12714 = ~n12708 & ~n12713;
  assign n12715 = ~n12707 & ~n12714;
  assign n12716 = po56  & ~n12715;
  assign n12717 = ~po56  & n12715;
  assign n12718 = ~n12235 & ~n12236;
  assign n12719 = po12  & n12718;
  assign n12720 = ~n12241 & ~n12719;
  assign n12721 = n12241 & n12719;
  assign n12722 = ~n12720 & ~n12721;
  assign n12723 = ~n12717 & ~n12722;
  assign n12724 = ~n12716 & ~n12723;
  assign n12725 = po57  & ~n12724;
  assign n12726 = ~po57  & n12724;
  assign n12727 = ~n12244 & ~n12245;
  assign n12728 = po12  & n12727;
  assign n12729 = ~n12250 & ~n12728;
  assign n12730 = n12250 & n12728;
  assign n12731 = ~n12729 & ~n12730;
  assign n12732 = ~n12726 & ~n12731;
  assign n12733 = ~n12725 & ~n12732;
  assign n12734 = po58  & ~n12733;
  assign n12735 = ~po58  & n12733;
  assign n12736 = ~n12253 & ~n12254;
  assign n12737 = po12  & n12736;
  assign n12738 = ~n12259 & ~n12737;
  assign n12739 = n12259 & n12737;
  assign n12740 = ~n12738 & ~n12739;
  assign n12741 = ~n12735 & ~n12740;
  assign n12742 = ~n12734 & ~n12741;
  assign n12743 = po59  & ~n12742;
  assign n12744 = ~po59  & n12742;
  assign n12745 = ~n12262 & ~n12263;
  assign n12746 = po12  & n12745;
  assign n12747 = ~n12268 & ~n12746;
  assign n12748 = n12268 & n12746;
  assign n12749 = ~n12747 & ~n12748;
  assign n12750 = ~n12744 & ~n12749;
  assign n12751 = ~n12743 & ~n12750;
  assign n12752 = po60  & ~n12751;
  assign n12753 = ~po60  & n12751;
  assign n12754 = ~n12271 & ~n12272;
  assign n12755 = po12  & n12754;
  assign n12756 = ~n12277 & ~n12755;
  assign n12757 = n12277 & n12755;
  assign n12758 = ~n12756 & ~n12757;
  assign n12759 = ~n12753 & ~n12758;
  assign n12760 = ~n12752 & ~n12759;
  assign n12761 = po61  & ~n12760;
  assign n12762 = ~po61  & n12760;
  assign n12763 = ~n12280 & ~n12281;
  assign n12764 = po12  & n12763;
  assign n12765 = ~n12286 & ~n12764;
  assign n12766 = n12286 & n12764;
  assign n12767 = ~n12765 & ~n12766;
  assign n12768 = ~n12762 & ~n12767;
  assign n12769 = ~n12761 & ~n12768;
  assign n12770 = po62  & ~n12769;
  assign n12771 = ~po62  & n12769;
  assign n12772 = ~n12289 & ~n12290;
  assign n12773 = po12  & n12772;
  assign n12774 = ~n12295 & ~n12773;
  assign n12775 = n12295 & n12773;
  assign n12776 = ~n12774 & ~n12775;
  assign n12777 = ~n12771 & ~n12776;
  assign n12778 = ~n12770 & ~n12777;
  assign n12779 = n12330 & n12778;
  assign n12780 = ~n12330 & ~n12778;
  assign n12781 = n12308 & po12 ;
  assign n12782 = ~n12307 & ~n12781;
  assign n12783 = n12780 & n12782;
  assign n12784 = ~po63  & ~n12783;
  assign n12785 = ~n12779 & ~n12784;
  assign n12786 = ~n12325 & n12785;
  assign po11  = n12321 | ~n12786;
  assign n12788 = ~n12694 & ~n12695;
  assign n12789 = po11  & n12788;
  assign n12790 = ~n12320 & ~n12789;
  assign n12791 = n12320 & n12789;
  assign n12792 = ~n12790 & ~n12791;
  assign n12793 = n12330 & ~po11 ;
  assign n12794 = ~n12330 & po11 ;
  assign n12795 = n12778 & ~n12794;
  assign n12796 = po63  & ~n12795;
  assign n12797 = ~n12780 & n12796;
  assign n12798 = ~n12770 & ~n12771;
  assign n12799 = po11  & n12798;
  assign n12800 = ~n12776 & ~n12799;
  assign n12801 = n12776 & n12799;
  assign n12802 = ~n12800 & ~n12801;
  assign n12803 = pi22  & po11 ;
  assign n12804 = ~pi20  & ~pi21 ;
  assign n12805 = ~pi22  & n12804;
  assign n12806 = ~n12803 & ~n12805;
  assign n12807 = po12  & ~n12806;
  assign n12808 = ~po12  & n12806;
  assign n12809 = ~pi22  & po11 ;
  assign n12810 = pi23  & ~n12809;
  assign n12811 = n12332 & po11 ;
  assign n12812 = ~n12810 & ~n12811;
  assign n12813 = ~n12808 & n12812;
  assign n12814 = ~n12807 & ~n12813;
  assign n12815 = po13  & ~n12814;
  assign n12816 = ~po13  & n12814;
  assign n12817 = po12  & n12786;
  assign n12818 = ~n12811 & ~n12817;
  assign n12819 = pi24  & ~n12818;
  assign n12820 = ~pi24  & n12818;
  assign n12821 = ~n12819 & ~n12820;
  assign n12822 = ~n12816 & ~n12821;
  assign n12823 = ~n12815 & ~n12822;
  assign n12824 = po14  & ~n12823;
  assign n12825 = ~po14  & n12823;
  assign n12826 = ~n12335 & ~n12336;
  assign n12827 = po11  & n12826;
  assign n12828 = n12340 & ~n12827;
  assign n12829 = ~n12340 & n12827;
  assign n12830 = ~n12828 & ~n12829;
  assign n12831 = ~n12825 & ~n12830;
  assign n12832 = ~n12824 & ~n12831;
  assign n12833 = po15  & ~n12832;
  assign n12834 = ~po15  & n12832;
  assign n12835 = ~n12343 & ~n12344;
  assign n12836 = po11  & n12835;
  assign n12837 = ~n12349 & ~n12836;
  assign n12838 = n12349 & n12836;
  assign n12839 = ~n12837 & ~n12838;
  assign n12840 = ~n12834 & ~n12839;
  assign n12841 = ~n12833 & ~n12840;
  assign n12842 = po16  & ~n12841;
  assign n12843 = ~po16  & n12841;
  assign n12844 = ~n12352 & ~n12353;
  assign n12845 = po11  & n12844;
  assign n12846 = n12358 & n12845;
  assign n12847 = ~n12358 & ~n12845;
  assign n12848 = ~n12846 & ~n12847;
  assign n12849 = ~n12843 & ~n12848;
  assign n12850 = ~n12842 & ~n12849;
  assign n12851 = po17  & ~n12850;
  assign n12852 = ~po17  & n12850;
  assign n12853 = ~n12361 & ~n12362;
  assign n12854 = po11  & n12853;
  assign n12855 = ~n12367 & ~n12854;
  assign n12856 = n12367 & n12854;
  assign n12857 = ~n12855 & ~n12856;
  assign n12858 = ~n12852 & ~n12857;
  assign n12859 = ~n12851 & ~n12858;
  assign n12860 = po18  & ~n12859;
  assign n12861 = ~po18  & n12859;
  assign n12862 = ~n12370 & ~n12371;
  assign n12863 = po11  & n12862;
  assign n12864 = ~n12376 & ~n12863;
  assign n12865 = n12376 & n12863;
  assign n12866 = ~n12864 & ~n12865;
  assign n12867 = ~n12861 & ~n12866;
  assign n12868 = ~n12860 & ~n12867;
  assign n12869 = po19  & ~n12868;
  assign n12870 = ~po19  & n12868;
  assign n12871 = ~n12379 & ~n12380;
  assign n12872 = po11  & n12871;
  assign n12873 = ~n12385 & ~n12872;
  assign n12874 = n12385 & n12872;
  assign n12875 = ~n12873 & ~n12874;
  assign n12876 = ~n12870 & ~n12875;
  assign n12877 = ~n12869 & ~n12876;
  assign n12878 = po20  & ~n12877;
  assign n12879 = ~po20  & n12877;
  assign n12880 = ~n12388 & ~n12389;
  assign n12881 = po11  & n12880;
  assign n12882 = ~n12394 & ~n12881;
  assign n12883 = n12394 & n12881;
  assign n12884 = ~n12882 & ~n12883;
  assign n12885 = ~n12879 & ~n12884;
  assign n12886 = ~n12878 & ~n12885;
  assign n12887 = po21  & ~n12886;
  assign n12888 = ~po21  & n12886;
  assign n12889 = ~n12397 & ~n12398;
  assign n12890 = po11  & n12889;
  assign n12891 = ~n12403 & ~n12890;
  assign n12892 = n12403 & n12890;
  assign n12893 = ~n12891 & ~n12892;
  assign n12894 = ~n12888 & ~n12893;
  assign n12895 = ~n12887 & ~n12894;
  assign n12896 = po22  & ~n12895;
  assign n12897 = ~po22  & n12895;
  assign n12898 = ~n12406 & ~n12407;
  assign n12899 = po11  & n12898;
  assign n12900 = ~n12412 & ~n12899;
  assign n12901 = n12412 & n12899;
  assign n12902 = ~n12900 & ~n12901;
  assign n12903 = ~n12897 & ~n12902;
  assign n12904 = ~n12896 & ~n12903;
  assign n12905 = po23  & ~n12904;
  assign n12906 = ~po23  & n12904;
  assign n12907 = ~n12415 & ~n12416;
  assign n12908 = po11  & n12907;
  assign n12909 = ~n12421 & ~n12908;
  assign n12910 = n12421 & n12908;
  assign n12911 = ~n12909 & ~n12910;
  assign n12912 = ~n12906 & ~n12911;
  assign n12913 = ~n12905 & ~n12912;
  assign n12914 = po24  & ~n12913;
  assign n12915 = ~po24  & n12913;
  assign n12916 = ~n12424 & ~n12425;
  assign n12917 = po11  & n12916;
  assign n12918 = ~n12430 & ~n12917;
  assign n12919 = n12430 & n12917;
  assign n12920 = ~n12918 & ~n12919;
  assign n12921 = ~n12915 & ~n12920;
  assign n12922 = ~n12914 & ~n12921;
  assign n12923 = po25  & ~n12922;
  assign n12924 = ~po25  & n12922;
  assign n12925 = ~n12433 & ~n12434;
  assign n12926 = po11  & n12925;
  assign n12927 = ~n12439 & ~n12926;
  assign n12928 = n12439 & n12926;
  assign n12929 = ~n12927 & ~n12928;
  assign n12930 = ~n12924 & ~n12929;
  assign n12931 = ~n12923 & ~n12930;
  assign n12932 = po26  & ~n12931;
  assign n12933 = ~po26  & n12931;
  assign n12934 = ~n12442 & ~n12443;
  assign n12935 = po11  & n12934;
  assign n12936 = ~n12448 & ~n12935;
  assign n12937 = n12448 & n12935;
  assign n12938 = ~n12936 & ~n12937;
  assign n12939 = ~n12933 & ~n12938;
  assign n12940 = ~n12932 & ~n12939;
  assign n12941 = po27  & ~n12940;
  assign n12942 = ~po27  & n12940;
  assign n12943 = ~n12451 & ~n12452;
  assign n12944 = po11  & n12943;
  assign n12945 = ~n12457 & ~n12944;
  assign n12946 = n12457 & n12944;
  assign n12947 = ~n12945 & ~n12946;
  assign n12948 = ~n12942 & ~n12947;
  assign n12949 = ~n12941 & ~n12948;
  assign n12950 = po28  & ~n12949;
  assign n12951 = ~po28  & n12949;
  assign n12952 = ~n12460 & ~n12461;
  assign n12953 = po11  & n12952;
  assign n12954 = ~n12466 & ~n12953;
  assign n12955 = n12466 & n12953;
  assign n12956 = ~n12954 & ~n12955;
  assign n12957 = ~n12951 & ~n12956;
  assign n12958 = ~n12950 & ~n12957;
  assign n12959 = po29  & ~n12958;
  assign n12960 = ~po29  & n12958;
  assign n12961 = ~n12469 & ~n12470;
  assign n12962 = po11  & n12961;
  assign n12963 = ~n12475 & ~n12962;
  assign n12964 = n12475 & n12962;
  assign n12965 = ~n12963 & ~n12964;
  assign n12966 = ~n12960 & ~n12965;
  assign n12967 = ~n12959 & ~n12966;
  assign n12968 = po30  & ~n12967;
  assign n12969 = ~po30  & n12967;
  assign n12970 = ~n12478 & ~n12479;
  assign n12971 = po11  & n12970;
  assign n12972 = ~n12484 & ~n12971;
  assign n12973 = n12484 & n12971;
  assign n12974 = ~n12972 & ~n12973;
  assign n12975 = ~n12969 & ~n12974;
  assign n12976 = ~n12968 & ~n12975;
  assign n12977 = po31  & ~n12976;
  assign n12978 = ~po31  & n12976;
  assign n12979 = ~n12487 & ~n12488;
  assign n12980 = po11  & n12979;
  assign n12981 = ~n12493 & ~n12980;
  assign n12982 = n12493 & n12980;
  assign n12983 = ~n12981 & ~n12982;
  assign n12984 = ~n12978 & ~n12983;
  assign n12985 = ~n12977 & ~n12984;
  assign n12986 = po32  & ~n12985;
  assign n12987 = ~po32  & n12985;
  assign n12988 = ~n12496 & ~n12497;
  assign n12989 = po11  & n12988;
  assign n12990 = ~n12502 & ~n12989;
  assign n12991 = n12502 & n12989;
  assign n12992 = ~n12990 & ~n12991;
  assign n12993 = ~n12987 & ~n12992;
  assign n12994 = ~n12986 & ~n12993;
  assign n12995 = po33  & ~n12994;
  assign n12996 = ~po33  & n12994;
  assign n12997 = ~n12505 & ~n12506;
  assign n12998 = po11  & n12997;
  assign n12999 = ~n12511 & ~n12998;
  assign n13000 = n12511 & n12998;
  assign n13001 = ~n12999 & ~n13000;
  assign n13002 = ~n12996 & ~n13001;
  assign n13003 = ~n12995 & ~n13002;
  assign n13004 = po34  & ~n13003;
  assign n13005 = ~po34  & n13003;
  assign n13006 = ~n12514 & ~n12515;
  assign n13007 = po11  & n13006;
  assign n13008 = ~n12520 & ~n13007;
  assign n13009 = n12520 & n13007;
  assign n13010 = ~n13008 & ~n13009;
  assign n13011 = ~n13005 & ~n13010;
  assign n13012 = ~n13004 & ~n13011;
  assign n13013 = po35  & ~n13012;
  assign n13014 = ~po35  & n13012;
  assign n13015 = ~n12523 & ~n12524;
  assign n13016 = po11  & n13015;
  assign n13017 = ~n12529 & ~n13016;
  assign n13018 = n12529 & n13016;
  assign n13019 = ~n13017 & ~n13018;
  assign n13020 = ~n13014 & ~n13019;
  assign n13021 = ~n13013 & ~n13020;
  assign n13022 = po36  & ~n13021;
  assign n13023 = ~po36  & n13021;
  assign n13024 = ~n12532 & ~n12533;
  assign n13025 = po11  & n13024;
  assign n13026 = ~n12538 & ~n13025;
  assign n13027 = n12538 & n13025;
  assign n13028 = ~n13026 & ~n13027;
  assign n13029 = ~n13023 & ~n13028;
  assign n13030 = ~n13022 & ~n13029;
  assign n13031 = po37  & ~n13030;
  assign n13032 = ~po37  & n13030;
  assign n13033 = ~n12541 & ~n12542;
  assign n13034 = po11  & n13033;
  assign n13035 = ~n12547 & ~n13034;
  assign n13036 = n12547 & n13034;
  assign n13037 = ~n13035 & ~n13036;
  assign n13038 = ~n13032 & ~n13037;
  assign n13039 = ~n13031 & ~n13038;
  assign n13040 = po38  & ~n13039;
  assign n13041 = ~po38  & n13039;
  assign n13042 = ~n12550 & ~n12551;
  assign n13043 = po11  & n13042;
  assign n13044 = ~n12556 & ~n13043;
  assign n13045 = n12556 & n13043;
  assign n13046 = ~n13044 & ~n13045;
  assign n13047 = ~n13041 & ~n13046;
  assign n13048 = ~n13040 & ~n13047;
  assign n13049 = po39  & ~n13048;
  assign n13050 = ~po39  & n13048;
  assign n13051 = ~n12559 & ~n12560;
  assign n13052 = po11  & n13051;
  assign n13053 = ~n12565 & ~n13052;
  assign n13054 = n12565 & n13052;
  assign n13055 = ~n13053 & ~n13054;
  assign n13056 = ~n13050 & ~n13055;
  assign n13057 = ~n13049 & ~n13056;
  assign n13058 = po40  & ~n13057;
  assign n13059 = ~po40  & n13057;
  assign n13060 = ~n12568 & ~n12569;
  assign n13061 = po11  & n13060;
  assign n13062 = ~n12574 & ~n13061;
  assign n13063 = n12574 & n13061;
  assign n13064 = ~n13062 & ~n13063;
  assign n13065 = ~n13059 & ~n13064;
  assign n13066 = ~n13058 & ~n13065;
  assign n13067 = po41  & ~n13066;
  assign n13068 = ~po41  & n13066;
  assign n13069 = ~n12577 & ~n12578;
  assign n13070 = po11  & n13069;
  assign n13071 = ~n12583 & ~n13070;
  assign n13072 = n12583 & n13070;
  assign n13073 = ~n13071 & ~n13072;
  assign n13074 = ~n13068 & ~n13073;
  assign n13075 = ~n13067 & ~n13074;
  assign n13076 = po42  & ~n13075;
  assign n13077 = ~po42  & n13075;
  assign n13078 = ~n12586 & ~n12587;
  assign n13079 = po11  & n13078;
  assign n13080 = ~n12592 & ~n13079;
  assign n13081 = n12592 & n13079;
  assign n13082 = ~n13080 & ~n13081;
  assign n13083 = ~n13077 & ~n13082;
  assign n13084 = ~n13076 & ~n13083;
  assign n13085 = po43  & ~n13084;
  assign n13086 = ~po43  & n13084;
  assign n13087 = ~n12595 & ~n12596;
  assign n13088 = po11  & n13087;
  assign n13089 = ~n12601 & ~n13088;
  assign n13090 = n12601 & n13088;
  assign n13091 = ~n13089 & ~n13090;
  assign n13092 = ~n13086 & ~n13091;
  assign n13093 = ~n13085 & ~n13092;
  assign n13094 = po44  & ~n13093;
  assign n13095 = ~po44  & n13093;
  assign n13096 = ~n12604 & ~n12605;
  assign n13097 = po11  & n13096;
  assign n13098 = ~n12610 & ~n13097;
  assign n13099 = n12610 & n13097;
  assign n13100 = ~n13098 & ~n13099;
  assign n13101 = ~n13095 & ~n13100;
  assign n13102 = ~n13094 & ~n13101;
  assign n13103 = po45  & ~n13102;
  assign n13104 = ~po45  & n13102;
  assign n13105 = ~n12613 & ~n12614;
  assign n13106 = po11  & n13105;
  assign n13107 = ~n12619 & ~n13106;
  assign n13108 = n12619 & n13106;
  assign n13109 = ~n13107 & ~n13108;
  assign n13110 = ~n13104 & ~n13109;
  assign n13111 = ~n13103 & ~n13110;
  assign n13112 = po46  & ~n13111;
  assign n13113 = ~po46  & n13111;
  assign n13114 = ~n12622 & ~n12623;
  assign n13115 = po11  & n13114;
  assign n13116 = ~n12628 & ~n13115;
  assign n13117 = n12628 & n13115;
  assign n13118 = ~n13116 & ~n13117;
  assign n13119 = ~n13113 & ~n13118;
  assign n13120 = ~n13112 & ~n13119;
  assign n13121 = po47  & ~n13120;
  assign n13122 = ~po47  & n13120;
  assign n13123 = ~n12631 & ~n12632;
  assign n13124 = po11  & n13123;
  assign n13125 = ~n12637 & ~n13124;
  assign n13126 = n12637 & n13124;
  assign n13127 = ~n13125 & ~n13126;
  assign n13128 = ~n13122 & ~n13127;
  assign n13129 = ~n13121 & ~n13128;
  assign n13130 = po48  & ~n13129;
  assign n13131 = ~po48  & n13129;
  assign n13132 = ~n12640 & ~n12641;
  assign n13133 = po11  & n13132;
  assign n13134 = ~n12646 & ~n13133;
  assign n13135 = n12646 & n13133;
  assign n13136 = ~n13134 & ~n13135;
  assign n13137 = ~n13131 & ~n13136;
  assign n13138 = ~n13130 & ~n13137;
  assign n13139 = po49  & ~n13138;
  assign n13140 = ~po49  & n13138;
  assign n13141 = ~n12649 & ~n12650;
  assign n13142 = po11  & n13141;
  assign n13143 = ~n12655 & ~n13142;
  assign n13144 = n12655 & n13142;
  assign n13145 = ~n13143 & ~n13144;
  assign n13146 = ~n13140 & ~n13145;
  assign n13147 = ~n13139 & ~n13146;
  assign n13148 = po50  & ~n13147;
  assign n13149 = ~po50  & n13147;
  assign n13150 = ~n12658 & ~n12659;
  assign n13151 = po11  & n13150;
  assign n13152 = ~n12664 & ~n13151;
  assign n13153 = n12664 & n13151;
  assign n13154 = ~n13152 & ~n13153;
  assign n13155 = ~n13149 & ~n13154;
  assign n13156 = ~n13148 & ~n13155;
  assign n13157 = po51  & ~n13156;
  assign n13158 = ~po51  & n13156;
  assign n13159 = ~n12667 & ~n12668;
  assign n13160 = po11  & n13159;
  assign n13161 = ~n12673 & ~n13160;
  assign n13162 = n12673 & n13160;
  assign n13163 = ~n13161 & ~n13162;
  assign n13164 = ~n13158 & ~n13163;
  assign n13165 = ~n13157 & ~n13164;
  assign n13166 = po52  & ~n13165;
  assign n13167 = ~po52  & n13165;
  assign n13168 = ~n12676 & ~n12677;
  assign n13169 = po11  & n13168;
  assign n13170 = ~n12682 & ~n13169;
  assign n13171 = n12682 & n13169;
  assign n13172 = ~n13170 & ~n13171;
  assign n13173 = ~n13167 & ~n13172;
  assign n13174 = ~n13166 & ~n13173;
  assign n13175 = po53  & ~n13174;
  assign n13176 = ~n12685 & ~n12691;
  assign n13177 = po11  & n13176;
  assign n13178 = ~n12690 & ~n13177;
  assign n13179 = n12690 & n13177;
  assign n13180 = ~n13178 & ~n13179;
  assign n13181 = ~po53  & n13174;
  assign n13182 = ~n13180 & ~n13181;
  assign n13183 = ~n13175 & ~n13182;
  assign n13184 = po54  & ~n13183;
  assign n13185 = ~po54  & n13183;
  assign n13186 = ~n12792 & ~n13185;
  assign n13187 = ~n13184 & ~n13186;
  assign n13188 = po55  & ~n13187;
  assign n13189 = ~po55  & n13187;
  assign n13190 = ~n12698 & ~n12699;
  assign n13191 = po11  & n13190;
  assign n13192 = ~n12704 & ~n13191;
  assign n13193 = n12704 & n13191;
  assign n13194 = ~n13192 & ~n13193;
  assign n13195 = ~n13189 & ~n13194;
  assign n13196 = ~n13188 & ~n13195;
  assign n13197 = po56  & ~n13196;
  assign n13198 = ~po56  & n13196;
  assign n13199 = ~n12707 & ~n12708;
  assign n13200 = po11  & n13199;
  assign n13201 = ~n12713 & ~n13200;
  assign n13202 = n12713 & n13200;
  assign n13203 = ~n13201 & ~n13202;
  assign n13204 = ~n13198 & ~n13203;
  assign n13205 = ~n13197 & ~n13204;
  assign n13206 = po57  & ~n13205;
  assign n13207 = ~po57  & n13205;
  assign n13208 = ~n12716 & ~n12717;
  assign n13209 = po11  & n13208;
  assign n13210 = ~n12722 & ~n13209;
  assign n13211 = n12722 & n13209;
  assign n13212 = ~n13210 & ~n13211;
  assign n13213 = ~n13207 & ~n13212;
  assign n13214 = ~n13206 & ~n13213;
  assign n13215 = po58  & ~n13214;
  assign n13216 = ~po58  & n13214;
  assign n13217 = ~n12725 & ~n12726;
  assign n13218 = po11  & n13217;
  assign n13219 = ~n12731 & ~n13218;
  assign n13220 = n12731 & n13218;
  assign n13221 = ~n13219 & ~n13220;
  assign n13222 = ~n13216 & ~n13221;
  assign n13223 = ~n13215 & ~n13222;
  assign n13224 = po59  & ~n13223;
  assign n13225 = ~po59  & n13223;
  assign n13226 = ~n12734 & ~n12735;
  assign n13227 = po11  & n13226;
  assign n13228 = ~n12740 & ~n13227;
  assign n13229 = n12740 & n13227;
  assign n13230 = ~n13228 & ~n13229;
  assign n13231 = ~n13225 & ~n13230;
  assign n13232 = ~n13224 & ~n13231;
  assign n13233 = po60  & ~n13232;
  assign n13234 = ~po60  & n13232;
  assign n13235 = ~n12743 & ~n12744;
  assign n13236 = po11  & n13235;
  assign n13237 = ~n12749 & ~n13236;
  assign n13238 = n12749 & n13236;
  assign n13239 = ~n13237 & ~n13238;
  assign n13240 = ~n13234 & ~n13239;
  assign n13241 = ~n13233 & ~n13240;
  assign n13242 = po61  & ~n13241;
  assign n13243 = ~po61  & n13241;
  assign n13244 = ~n12752 & ~n12753;
  assign n13245 = po11  & n13244;
  assign n13246 = ~n12758 & ~n13245;
  assign n13247 = n12758 & n13245;
  assign n13248 = ~n13246 & ~n13247;
  assign n13249 = ~n13243 & ~n13248;
  assign n13250 = ~n13242 & ~n13249;
  assign n13251 = po62  & ~n13250;
  assign n13252 = ~po62  & n13250;
  assign n13253 = ~n12761 & ~n12762;
  assign n13254 = po11  & n13253;
  assign n13255 = ~n12767 & ~n13254;
  assign n13256 = n12767 & n13254;
  assign n13257 = ~n13255 & ~n13256;
  assign n13258 = ~n13252 & ~n13257;
  assign n13259 = ~n13251 & ~n13258;
  assign n13260 = n12802 & n13259;
  assign n13261 = ~n12802 & ~n13259;
  assign n13262 = n12780 & po11 ;
  assign n13263 = ~n12779 & ~n13262;
  assign n13264 = n13261 & n13263;
  assign n13265 = ~po63  & ~n13264;
  assign n13266 = ~n13260 & ~n13265;
  assign n13267 = ~n12797 & n13266;
  assign po10  = n12793 | ~n13267;
  assign n13269 = ~n13184 & ~n13185;
  assign n13270 = po10  & n13269;
  assign n13271 = ~n12792 & ~n13270;
  assign n13272 = n12792 & n13270;
  assign n13273 = ~n13271 & ~n13272;
  assign n13274 = n12802 & ~po10 ;
  assign n13275 = ~n12802 & po10 ;
  assign n13276 = n13259 & ~n13275;
  assign n13277 = po63  & ~n13276;
  assign n13278 = ~n13261 & n13277;
  assign n13279 = ~n13251 & ~n13252;
  assign n13280 = po10  & n13279;
  assign n13281 = ~n13257 & ~n13280;
  assign n13282 = n13257 & n13280;
  assign n13283 = ~n13281 & ~n13282;
  assign n13284 = pi20  & po10 ;
  assign n13285 = ~pi18  & ~pi19 ;
  assign n13286 = ~pi20  & n13285;
  assign n13287 = ~n13284 & ~n13286;
  assign n13288 = po11  & ~n13287;
  assign n13289 = ~po11  & n13287;
  assign n13290 = ~pi20  & po10 ;
  assign n13291 = pi21  & ~n13290;
  assign n13292 = n12804 & po10 ;
  assign n13293 = ~n13291 & ~n13292;
  assign n13294 = ~n13289 & n13293;
  assign n13295 = ~n13288 & ~n13294;
  assign n13296 = po12  & ~n13295;
  assign n13297 = ~po12  & n13295;
  assign n13298 = po11  & n13267;
  assign n13299 = ~n13292 & ~n13298;
  assign n13300 = pi22  & ~n13299;
  assign n13301 = ~pi22  & n13299;
  assign n13302 = ~n13300 & ~n13301;
  assign n13303 = ~n13297 & ~n13302;
  assign n13304 = ~n13296 & ~n13303;
  assign n13305 = po13  & ~n13304;
  assign n13306 = ~po13  & n13304;
  assign n13307 = ~n12807 & ~n12808;
  assign n13308 = po10  & n13307;
  assign n13309 = n12812 & ~n13308;
  assign n13310 = ~n12812 & n13308;
  assign n13311 = ~n13309 & ~n13310;
  assign n13312 = ~n13306 & ~n13311;
  assign n13313 = ~n13305 & ~n13312;
  assign n13314 = po14  & ~n13313;
  assign n13315 = ~po14  & n13313;
  assign n13316 = ~n12815 & ~n12816;
  assign n13317 = po10  & n13316;
  assign n13318 = ~n12821 & ~n13317;
  assign n13319 = n12821 & n13317;
  assign n13320 = ~n13318 & ~n13319;
  assign n13321 = ~n13315 & ~n13320;
  assign n13322 = ~n13314 & ~n13321;
  assign n13323 = po15  & ~n13322;
  assign n13324 = ~po15  & n13322;
  assign n13325 = ~n12824 & ~n12825;
  assign n13326 = po10  & n13325;
  assign n13327 = n12830 & n13326;
  assign n13328 = ~n12830 & ~n13326;
  assign n13329 = ~n13327 & ~n13328;
  assign n13330 = ~n13324 & ~n13329;
  assign n13331 = ~n13323 & ~n13330;
  assign n13332 = po16  & ~n13331;
  assign n13333 = ~po16  & n13331;
  assign n13334 = ~n12833 & ~n12834;
  assign n13335 = po10  & n13334;
  assign n13336 = ~n12839 & ~n13335;
  assign n13337 = n12839 & n13335;
  assign n13338 = ~n13336 & ~n13337;
  assign n13339 = ~n13333 & ~n13338;
  assign n13340 = ~n13332 & ~n13339;
  assign n13341 = po17  & ~n13340;
  assign n13342 = ~po17  & n13340;
  assign n13343 = ~n12842 & ~n12843;
  assign n13344 = po10  & n13343;
  assign n13345 = ~n12848 & ~n13344;
  assign n13346 = n12848 & n13344;
  assign n13347 = ~n13345 & ~n13346;
  assign n13348 = ~n13342 & ~n13347;
  assign n13349 = ~n13341 & ~n13348;
  assign n13350 = po18  & ~n13349;
  assign n13351 = ~po18  & n13349;
  assign n13352 = ~n12851 & ~n12852;
  assign n13353 = po10  & n13352;
  assign n13354 = ~n12857 & ~n13353;
  assign n13355 = n12857 & n13353;
  assign n13356 = ~n13354 & ~n13355;
  assign n13357 = ~n13351 & ~n13356;
  assign n13358 = ~n13350 & ~n13357;
  assign n13359 = po19  & ~n13358;
  assign n13360 = ~po19  & n13358;
  assign n13361 = ~n12860 & ~n12861;
  assign n13362 = po10  & n13361;
  assign n13363 = ~n12866 & ~n13362;
  assign n13364 = n12866 & n13362;
  assign n13365 = ~n13363 & ~n13364;
  assign n13366 = ~n13360 & ~n13365;
  assign n13367 = ~n13359 & ~n13366;
  assign n13368 = po20  & ~n13367;
  assign n13369 = ~po20  & n13367;
  assign n13370 = ~n12869 & ~n12870;
  assign n13371 = po10  & n13370;
  assign n13372 = ~n12875 & ~n13371;
  assign n13373 = n12875 & n13371;
  assign n13374 = ~n13372 & ~n13373;
  assign n13375 = ~n13369 & ~n13374;
  assign n13376 = ~n13368 & ~n13375;
  assign n13377 = po21  & ~n13376;
  assign n13378 = ~po21  & n13376;
  assign n13379 = ~n12878 & ~n12879;
  assign n13380 = po10  & n13379;
  assign n13381 = ~n12884 & ~n13380;
  assign n13382 = n12884 & n13380;
  assign n13383 = ~n13381 & ~n13382;
  assign n13384 = ~n13378 & ~n13383;
  assign n13385 = ~n13377 & ~n13384;
  assign n13386 = po22  & ~n13385;
  assign n13387 = ~po22  & n13385;
  assign n13388 = ~n12887 & ~n12888;
  assign n13389 = po10  & n13388;
  assign n13390 = ~n12893 & ~n13389;
  assign n13391 = n12893 & n13389;
  assign n13392 = ~n13390 & ~n13391;
  assign n13393 = ~n13387 & ~n13392;
  assign n13394 = ~n13386 & ~n13393;
  assign n13395 = po23  & ~n13394;
  assign n13396 = ~po23  & n13394;
  assign n13397 = ~n12896 & ~n12897;
  assign n13398 = po10  & n13397;
  assign n13399 = ~n12902 & ~n13398;
  assign n13400 = n12902 & n13398;
  assign n13401 = ~n13399 & ~n13400;
  assign n13402 = ~n13396 & ~n13401;
  assign n13403 = ~n13395 & ~n13402;
  assign n13404 = po24  & ~n13403;
  assign n13405 = ~po24  & n13403;
  assign n13406 = ~n12905 & ~n12906;
  assign n13407 = po10  & n13406;
  assign n13408 = ~n12911 & ~n13407;
  assign n13409 = n12911 & n13407;
  assign n13410 = ~n13408 & ~n13409;
  assign n13411 = ~n13405 & ~n13410;
  assign n13412 = ~n13404 & ~n13411;
  assign n13413 = po25  & ~n13412;
  assign n13414 = ~po25  & n13412;
  assign n13415 = ~n12914 & ~n12915;
  assign n13416 = po10  & n13415;
  assign n13417 = ~n12920 & ~n13416;
  assign n13418 = n12920 & n13416;
  assign n13419 = ~n13417 & ~n13418;
  assign n13420 = ~n13414 & ~n13419;
  assign n13421 = ~n13413 & ~n13420;
  assign n13422 = po26  & ~n13421;
  assign n13423 = ~po26  & n13421;
  assign n13424 = ~n12923 & ~n12924;
  assign n13425 = po10  & n13424;
  assign n13426 = ~n12929 & ~n13425;
  assign n13427 = n12929 & n13425;
  assign n13428 = ~n13426 & ~n13427;
  assign n13429 = ~n13423 & ~n13428;
  assign n13430 = ~n13422 & ~n13429;
  assign n13431 = po27  & ~n13430;
  assign n13432 = ~po27  & n13430;
  assign n13433 = ~n12932 & ~n12933;
  assign n13434 = po10  & n13433;
  assign n13435 = ~n12938 & ~n13434;
  assign n13436 = n12938 & n13434;
  assign n13437 = ~n13435 & ~n13436;
  assign n13438 = ~n13432 & ~n13437;
  assign n13439 = ~n13431 & ~n13438;
  assign n13440 = po28  & ~n13439;
  assign n13441 = ~po28  & n13439;
  assign n13442 = ~n12941 & ~n12942;
  assign n13443 = po10  & n13442;
  assign n13444 = ~n12947 & ~n13443;
  assign n13445 = n12947 & n13443;
  assign n13446 = ~n13444 & ~n13445;
  assign n13447 = ~n13441 & ~n13446;
  assign n13448 = ~n13440 & ~n13447;
  assign n13449 = po29  & ~n13448;
  assign n13450 = ~po29  & n13448;
  assign n13451 = ~n12950 & ~n12951;
  assign n13452 = po10  & n13451;
  assign n13453 = ~n12956 & ~n13452;
  assign n13454 = n12956 & n13452;
  assign n13455 = ~n13453 & ~n13454;
  assign n13456 = ~n13450 & ~n13455;
  assign n13457 = ~n13449 & ~n13456;
  assign n13458 = po30  & ~n13457;
  assign n13459 = ~po30  & n13457;
  assign n13460 = ~n12959 & ~n12960;
  assign n13461 = po10  & n13460;
  assign n13462 = ~n12965 & ~n13461;
  assign n13463 = n12965 & n13461;
  assign n13464 = ~n13462 & ~n13463;
  assign n13465 = ~n13459 & ~n13464;
  assign n13466 = ~n13458 & ~n13465;
  assign n13467 = po31  & ~n13466;
  assign n13468 = ~po31  & n13466;
  assign n13469 = ~n12968 & ~n12969;
  assign n13470 = po10  & n13469;
  assign n13471 = ~n12974 & ~n13470;
  assign n13472 = n12974 & n13470;
  assign n13473 = ~n13471 & ~n13472;
  assign n13474 = ~n13468 & ~n13473;
  assign n13475 = ~n13467 & ~n13474;
  assign n13476 = po32  & ~n13475;
  assign n13477 = ~po32  & n13475;
  assign n13478 = ~n12977 & ~n12978;
  assign n13479 = po10  & n13478;
  assign n13480 = ~n12983 & ~n13479;
  assign n13481 = n12983 & n13479;
  assign n13482 = ~n13480 & ~n13481;
  assign n13483 = ~n13477 & ~n13482;
  assign n13484 = ~n13476 & ~n13483;
  assign n13485 = po33  & ~n13484;
  assign n13486 = ~po33  & n13484;
  assign n13487 = ~n12986 & ~n12987;
  assign n13488 = po10  & n13487;
  assign n13489 = ~n12992 & ~n13488;
  assign n13490 = n12992 & n13488;
  assign n13491 = ~n13489 & ~n13490;
  assign n13492 = ~n13486 & ~n13491;
  assign n13493 = ~n13485 & ~n13492;
  assign n13494 = po34  & ~n13493;
  assign n13495 = ~po34  & n13493;
  assign n13496 = ~n12995 & ~n12996;
  assign n13497 = po10  & n13496;
  assign n13498 = ~n13001 & ~n13497;
  assign n13499 = n13001 & n13497;
  assign n13500 = ~n13498 & ~n13499;
  assign n13501 = ~n13495 & ~n13500;
  assign n13502 = ~n13494 & ~n13501;
  assign n13503 = po35  & ~n13502;
  assign n13504 = ~po35  & n13502;
  assign n13505 = ~n13004 & ~n13005;
  assign n13506 = po10  & n13505;
  assign n13507 = ~n13010 & ~n13506;
  assign n13508 = n13010 & n13506;
  assign n13509 = ~n13507 & ~n13508;
  assign n13510 = ~n13504 & ~n13509;
  assign n13511 = ~n13503 & ~n13510;
  assign n13512 = po36  & ~n13511;
  assign n13513 = ~po36  & n13511;
  assign n13514 = ~n13013 & ~n13014;
  assign n13515 = po10  & n13514;
  assign n13516 = ~n13019 & ~n13515;
  assign n13517 = n13019 & n13515;
  assign n13518 = ~n13516 & ~n13517;
  assign n13519 = ~n13513 & ~n13518;
  assign n13520 = ~n13512 & ~n13519;
  assign n13521 = po37  & ~n13520;
  assign n13522 = ~po37  & n13520;
  assign n13523 = ~n13022 & ~n13023;
  assign n13524 = po10  & n13523;
  assign n13525 = ~n13028 & ~n13524;
  assign n13526 = n13028 & n13524;
  assign n13527 = ~n13525 & ~n13526;
  assign n13528 = ~n13522 & ~n13527;
  assign n13529 = ~n13521 & ~n13528;
  assign n13530 = po38  & ~n13529;
  assign n13531 = ~po38  & n13529;
  assign n13532 = ~n13031 & ~n13032;
  assign n13533 = po10  & n13532;
  assign n13534 = ~n13037 & ~n13533;
  assign n13535 = n13037 & n13533;
  assign n13536 = ~n13534 & ~n13535;
  assign n13537 = ~n13531 & ~n13536;
  assign n13538 = ~n13530 & ~n13537;
  assign n13539 = po39  & ~n13538;
  assign n13540 = ~po39  & n13538;
  assign n13541 = ~n13040 & ~n13041;
  assign n13542 = po10  & n13541;
  assign n13543 = ~n13046 & ~n13542;
  assign n13544 = n13046 & n13542;
  assign n13545 = ~n13543 & ~n13544;
  assign n13546 = ~n13540 & ~n13545;
  assign n13547 = ~n13539 & ~n13546;
  assign n13548 = po40  & ~n13547;
  assign n13549 = ~po40  & n13547;
  assign n13550 = ~n13049 & ~n13050;
  assign n13551 = po10  & n13550;
  assign n13552 = ~n13055 & ~n13551;
  assign n13553 = n13055 & n13551;
  assign n13554 = ~n13552 & ~n13553;
  assign n13555 = ~n13549 & ~n13554;
  assign n13556 = ~n13548 & ~n13555;
  assign n13557 = po41  & ~n13556;
  assign n13558 = ~po41  & n13556;
  assign n13559 = ~n13058 & ~n13059;
  assign n13560 = po10  & n13559;
  assign n13561 = ~n13064 & ~n13560;
  assign n13562 = n13064 & n13560;
  assign n13563 = ~n13561 & ~n13562;
  assign n13564 = ~n13558 & ~n13563;
  assign n13565 = ~n13557 & ~n13564;
  assign n13566 = po42  & ~n13565;
  assign n13567 = ~po42  & n13565;
  assign n13568 = ~n13067 & ~n13068;
  assign n13569 = po10  & n13568;
  assign n13570 = ~n13073 & ~n13569;
  assign n13571 = n13073 & n13569;
  assign n13572 = ~n13570 & ~n13571;
  assign n13573 = ~n13567 & ~n13572;
  assign n13574 = ~n13566 & ~n13573;
  assign n13575 = po43  & ~n13574;
  assign n13576 = ~po43  & n13574;
  assign n13577 = ~n13076 & ~n13077;
  assign n13578 = po10  & n13577;
  assign n13579 = ~n13082 & ~n13578;
  assign n13580 = n13082 & n13578;
  assign n13581 = ~n13579 & ~n13580;
  assign n13582 = ~n13576 & ~n13581;
  assign n13583 = ~n13575 & ~n13582;
  assign n13584 = po44  & ~n13583;
  assign n13585 = ~po44  & n13583;
  assign n13586 = ~n13085 & ~n13086;
  assign n13587 = po10  & n13586;
  assign n13588 = ~n13091 & ~n13587;
  assign n13589 = n13091 & n13587;
  assign n13590 = ~n13588 & ~n13589;
  assign n13591 = ~n13585 & ~n13590;
  assign n13592 = ~n13584 & ~n13591;
  assign n13593 = po45  & ~n13592;
  assign n13594 = ~po45  & n13592;
  assign n13595 = ~n13094 & ~n13095;
  assign n13596 = po10  & n13595;
  assign n13597 = ~n13100 & ~n13596;
  assign n13598 = n13100 & n13596;
  assign n13599 = ~n13597 & ~n13598;
  assign n13600 = ~n13594 & ~n13599;
  assign n13601 = ~n13593 & ~n13600;
  assign n13602 = po46  & ~n13601;
  assign n13603 = ~po46  & n13601;
  assign n13604 = ~n13103 & ~n13104;
  assign n13605 = po10  & n13604;
  assign n13606 = ~n13109 & ~n13605;
  assign n13607 = n13109 & n13605;
  assign n13608 = ~n13606 & ~n13607;
  assign n13609 = ~n13603 & ~n13608;
  assign n13610 = ~n13602 & ~n13609;
  assign n13611 = po47  & ~n13610;
  assign n13612 = ~po47  & n13610;
  assign n13613 = ~n13112 & ~n13113;
  assign n13614 = po10  & n13613;
  assign n13615 = ~n13118 & ~n13614;
  assign n13616 = n13118 & n13614;
  assign n13617 = ~n13615 & ~n13616;
  assign n13618 = ~n13612 & ~n13617;
  assign n13619 = ~n13611 & ~n13618;
  assign n13620 = po48  & ~n13619;
  assign n13621 = ~po48  & n13619;
  assign n13622 = ~n13121 & ~n13122;
  assign n13623 = po10  & n13622;
  assign n13624 = ~n13127 & ~n13623;
  assign n13625 = n13127 & n13623;
  assign n13626 = ~n13624 & ~n13625;
  assign n13627 = ~n13621 & ~n13626;
  assign n13628 = ~n13620 & ~n13627;
  assign n13629 = po49  & ~n13628;
  assign n13630 = ~po49  & n13628;
  assign n13631 = ~n13130 & ~n13131;
  assign n13632 = po10  & n13631;
  assign n13633 = ~n13136 & ~n13632;
  assign n13634 = n13136 & n13632;
  assign n13635 = ~n13633 & ~n13634;
  assign n13636 = ~n13630 & ~n13635;
  assign n13637 = ~n13629 & ~n13636;
  assign n13638 = po50  & ~n13637;
  assign n13639 = ~po50  & n13637;
  assign n13640 = ~n13139 & ~n13140;
  assign n13641 = po10  & n13640;
  assign n13642 = ~n13145 & ~n13641;
  assign n13643 = n13145 & n13641;
  assign n13644 = ~n13642 & ~n13643;
  assign n13645 = ~n13639 & ~n13644;
  assign n13646 = ~n13638 & ~n13645;
  assign n13647 = po51  & ~n13646;
  assign n13648 = ~po51  & n13646;
  assign n13649 = ~n13148 & ~n13149;
  assign n13650 = po10  & n13649;
  assign n13651 = ~n13154 & ~n13650;
  assign n13652 = n13154 & n13650;
  assign n13653 = ~n13651 & ~n13652;
  assign n13654 = ~n13648 & ~n13653;
  assign n13655 = ~n13647 & ~n13654;
  assign n13656 = po52  & ~n13655;
  assign n13657 = ~po52  & n13655;
  assign n13658 = ~n13157 & ~n13158;
  assign n13659 = po10  & n13658;
  assign n13660 = ~n13163 & ~n13659;
  assign n13661 = n13163 & n13659;
  assign n13662 = ~n13660 & ~n13661;
  assign n13663 = ~n13657 & ~n13662;
  assign n13664 = ~n13656 & ~n13663;
  assign n13665 = po53  & ~n13664;
  assign n13666 = ~po53  & n13664;
  assign n13667 = ~n13166 & ~n13167;
  assign n13668 = po10  & n13667;
  assign n13669 = ~n13172 & ~n13668;
  assign n13670 = n13172 & n13668;
  assign n13671 = ~n13669 & ~n13670;
  assign n13672 = ~n13666 & ~n13671;
  assign n13673 = ~n13665 & ~n13672;
  assign n13674 = po54  & ~n13673;
  assign n13675 = ~n13175 & ~n13181;
  assign n13676 = po10  & n13675;
  assign n13677 = ~n13180 & ~n13676;
  assign n13678 = n13180 & n13676;
  assign n13679 = ~n13677 & ~n13678;
  assign n13680 = ~po54  & n13673;
  assign n13681 = ~n13679 & ~n13680;
  assign n13682 = ~n13674 & ~n13681;
  assign n13683 = po55  & ~n13682;
  assign n13684 = ~po55  & n13682;
  assign n13685 = ~n13273 & ~n13684;
  assign n13686 = ~n13683 & ~n13685;
  assign n13687 = po56  & ~n13686;
  assign n13688 = ~po56  & n13686;
  assign n13689 = ~n13188 & ~n13189;
  assign n13690 = po10  & n13689;
  assign n13691 = ~n13194 & ~n13690;
  assign n13692 = n13194 & n13690;
  assign n13693 = ~n13691 & ~n13692;
  assign n13694 = ~n13688 & ~n13693;
  assign n13695 = ~n13687 & ~n13694;
  assign n13696 = po57  & ~n13695;
  assign n13697 = ~po57  & n13695;
  assign n13698 = ~n13197 & ~n13198;
  assign n13699 = po10  & n13698;
  assign n13700 = ~n13203 & ~n13699;
  assign n13701 = n13203 & n13699;
  assign n13702 = ~n13700 & ~n13701;
  assign n13703 = ~n13697 & ~n13702;
  assign n13704 = ~n13696 & ~n13703;
  assign n13705 = po58  & ~n13704;
  assign n13706 = ~po58  & n13704;
  assign n13707 = ~n13206 & ~n13207;
  assign n13708 = po10  & n13707;
  assign n13709 = ~n13212 & ~n13708;
  assign n13710 = n13212 & n13708;
  assign n13711 = ~n13709 & ~n13710;
  assign n13712 = ~n13706 & ~n13711;
  assign n13713 = ~n13705 & ~n13712;
  assign n13714 = po59  & ~n13713;
  assign n13715 = ~po59  & n13713;
  assign n13716 = ~n13215 & ~n13216;
  assign n13717 = po10  & n13716;
  assign n13718 = ~n13221 & ~n13717;
  assign n13719 = n13221 & n13717;
  assign n13720 = ~n13718 & ~n13719;
  assign n13721 = ~n13715 & ~n13720;
  assign n13722 = ~n13714 & ~n13721;
  assign n13723 = po60  & ~n13722;
  assign n13724 = ~po60  & n13722;
  assign n13725 = ~n13224 & ~n13225;
  assign n13726 = po10  & n13725;
  assign n13727 = ~n13230 & ~n13726;
  assign n13728 = n13230 & n13726;
  assign n13729 = ~n13727 & ~n13728;
  assign n13730 = ~n13724 & ~n13729;
  assign n13731 = ~n13723 & ~n13730;
  assign n13732 = po61  & ~n13731;
  assign n13733 = ~po61  & n13731;
  assign n13734 = ~n13233 & ~n13234;
  assign n13735 = po10  & n13734;
  assign n13736 = ~n13239 & ~n13735;
  assign n13737 = n13239 & n13735;
  assign n13738 = ~n13736 & ~n13737;
  assign n13739 = ~n13733 & ~n13738;
  assign n13740 = ~n13732 & ~n13739;
  assign n13741 = po62  & ~n13740;
  assign n13742 = ~po62  & n13740;
  assign n13743 = ~n13242 & ~n13243;
  assign n13744 = po10  & n13743;
  assign n13745 = ~n13248 & ~n13744;
  assign n13746 = n13248 & n13744;
  assign n13747 = ~n13745 & ~n13746;
  assign n13748 = ~n13742 & ~n13747;
  assign n13749 = ~n13741 & ~n13748;
  assign n13750 = n13283 & n13749;
  assign n13751 = ~n13283 & ~n13749;
  assign n13752 = n13261 & po10 ;
  assign n13753 = ~n13260 & ~n13752;
  assign n13754 = n13751 & n13753;
  assign n13755 = ~po63  & ~n13754;
  assign n13756 = ~n13750 & ~n13755;
  assign n13757 = ~n13278 & n13756;
  assign po9  = n13274 | ~n13757;
  assign n13759 = ~n13683 & ~n13684;
  assign n13760 = po9  & n13759;
  assign n13761 = ~n13273 & ~n13760;
  assign n13762 = n13273 & n13760;
  assign n13763 = ~n13761 & ~n13762;
  assign n13764 = n13283 & ~po9 ;
  assign n13765 = ~n13283 & po9 ;
  assign n13766 = n13749 & ~n13765;
  assign n13767 = po63  & ~n13766;
  assign n13768 = ~n13751 & n13767;
  assign n13769 = ~n13741 & ~n13742;
  assign n13770 = po9  & n13769;
  assign n13771 = ~n13747 & ~n13770;
  assign n13772 = n13747 & n13770;
  assign n13773 = ~n13771 & ~n13772;
  assign n13774 = pi18  & po9 ;
  assign n13775 = ~pi16  & ~pi17 ;
  assign n13776 = ~pi18  & n13775;
  assign n13777 = ~n13774 & ~n13776;
  assign n13778 = po10  & ~n13777;
  assign n13779 = ~po10  & n13777;
  assign n13780 = ~pi18  & po9 ;
  assign n13781 = pi19  & ~n13780;
  assign n13782 = n13285 & po9 ;
  assign n13783 = ~n13781 & ~n13782;
  assign n13784 = ~n13779 & n13783;
  assign n13785 = ~n13778 & ~n13784;
  assign n13786 = po11  & ~n13785;
  assign n13787 = ~po11  & n13785;
  assign n13788 = po10  & n13757;
  assign n13789 = ~n13782 & ~n13788;
  assign n13790 = pi20  & ~n13789;
  assign n13791 = ~pi20  & n13789;
  assign n13792 = ~n13790 & ~n13791;
  assign n13793 = ~n13787 & ~n13792;
  assign n13794 = ~n13786 & ~n13793;
  assign n13795 = po12  & ~n13794;
  assign n13796 = ~po12  & n13794;
  assign n13797 = ~n13288 & ~n13289;
  assign n13798 = po9  & n13797;
  assign n13799 = n13293 & ~n13798;
  assign n13800 = ~n13293 & n13798;
  assign n13801 = ~n13799 & ~n13800;
  assign n13802 = ~n13796 & ~n13801;
  assign n13803 = ~n13795 & ~n13802;
  assign n13804 = po13  & ~n13803;
  assign n13805 = ~po13  & n13803;
  assign n13806 = ~n13296 & ~n13297;
  assign n13807 = po9  & n13806;
  assign n13808 = ~n13302 & ~n13807;
  assign n13809 = n13302 & n13807;
  assign n13810 = ~n13808 & ~n13809;
  assign n13811 = ~n13805 & ~n13810;
  assign n13812 = ~n13804 & ~n13811;
  assign n13813 = po14  & ~n13812;
  assign n13814 = ~po14  & n13812;
  assign n13815 = ~n13305 & ~n13306;
  assign n13816 = po9  & n13815;
  assign n13817 = n13311 & n13816;
  assign n13818 = ~n13311 & ~n13816;
  assign n13819 = ~n13817 & ~n13818;
  assign n13820 = ~n13814 & ~n13819;
  assign n13821 = ~n13813 & ~n13820;
  assign n13822 = po15  & ~n13821;
  assign n13823 = ~po15  & n13821;
  assign n13824 = ~n13314 & ~n13315;
  assign n13825 = po9  & n13824;
  assign n13826 = ~n13320 & ~n13825;
  assign n13827 = n13320 & n13825;
  assign n13828 = ~n13826 & ~n13827;
  assign n13829 = ~n13823 & ~n13828;
  assign n13830 = ~n13822 & ~n13829;
  assign n13831 = po16  & ~n13830;
  assign n13832 = ~po16  & n13830;
  assign n13833 = ~n13323 & ~n13324;
  assign n13834 = po9  & n13833;
  assign n13835 = ~n13329 & ~n13834;
  assign n13836 = n13329 & n13834;
  assign n13837 = ~n13835 & ~n13836;
  assign n13838 = ~n13832 & ~n13837;
  assign n13839 = ~n13831 & ~n13838;
  assign n13840 = po17  & ~n13839;
  assign n13841 = ~po17  & n13839;
  assign n13842 = ~n13332 & ~n13333;
  assign n13843 = po9  & n13842;
  assign n13844 = ~n13338 & ~n13843;
  assign n13845 = n13338 & n13843;
  assign n13846 = ~n13844 & ~n13845;
  assign n13847 = ~n13841 & ~n13846;
  assign n13848 = ~n13840 & ~n13847;
  assign n13849 = po18  & ~n13848;
  assign n13850 = ~po18  & n13848;
  assign n13851 = ~n13341 & ~n13342;
  assign n13852 = po9  & n13851;
  assign n13853 = ~n13347 & ~n13852;
  assign n13854 = n13347 & n13852;
  assign n13855 = ~n13853 & ~n13854;
  assign n13856 = ~n13850 & ~n13855;
  assign n13857 = ~n13849 & ~n13856;
  assign n13858 = po19  & ~n13857;
  assign n13859 = ~po19  & n13857;
  assign n13860 = ~n13350 & ~n13351;
  assign n13861 = po9  & n13860;
  assign n13862 = ~n13356 & ~n13861;
  assign n13863 = n13356 & n13861;
  assign n13864 = ~n13862 & ~n13863;
  assign n13865 = ~n13859 & ~n13864;
  assign n13866 = ~n13858 & ~n13865;
  assign n13867 = po20  & ~n13866;
  assign n13868 = ~po20  & n13866;
  assign n13869 = ~n13359 & ~n13360;
  assign n13870 = po9  & n13869;
  assign n13871 = ~n13365 & ~n13870;
  assign n13872 = n13365 & n13870;
  assign n13873 = ~n13871 & ~n13872;
  assign n13874 = ~n13868 & ~n13873;
  assign n13875 = ~n13867 & ~n13874;
  assign n13876 = po21  & ~n13875;
  assign n13877 = ~po21  & n13875;
  assign n13878 = ~n13368 & ~n13369;
  assign n13879 = po9  & n13878;
  assign n13880 = ~n13374 & ~n13879;
  assign n13881 = n13374 & n13879;
  assign n13882 = ~n13880 & ~n13881;
  assign n13883 = ~n13877 & ~n13882;
  assign n13884 = ~n13876 & ~n13883;
  assign n13885 = po22  & ~n13884;
  assign n13886 = ~po22  & n13884;
  assign n13887 = ~n13377 & ~n13378;
  assign n13888 = po9  & n13887;
  assign n13889 = ~n13383 & ~n13888;
  assign n13890 = n13383 & n13888;
  assign n13891 = ~n13889 & ~n13890;
  assign n13892 = ~n13886 & ~n13891;
  assign n13893 = ~n13885 & ~n13892;
  assign n13894 = po23  & ~n13893;
  assign n13895 = ~po23  & n13893;
  assign n13896 = ~n13386 & ~n13387;
  assign n13897 = po9  & n13896;
  assign n13898 = ~n13392 & ~n13897;
  assign n13899 = n13392 & n13897;
  assign n13900 = ~n13898 & ~n13899;
  assign n13901 = ~n13895 & ~n13900;
  assign n13902 = ~n13894 & ~n13901;
  assign n13903 = po24  & ~n13902;
  assign n13904 = ~po24  & n13902;
  assign n13905 = ~n13395 & ~n13396;
  assign n13906 = po9  & n13905;
  assign n13907 = ~n13401 & ~n13906;
  assign n13908 = n13401 & n13906;
  assign n13909 = ~n13907 & ~n13908;
  assign n13910 = ~n13904 & ~n13909;
  assign n13911 = ~n13903 & ~n13910;
  assign n13912 = po25  & ~n13911;
  assign n13913 = ~po25  & n13911;
  assign n13914 = ~n13404 & ~n13405;
  assign n13915 = po9  & n13914;
  assign n13916 = ~n13410 & ~n13915;
  assign n13917 = n13410 & n13915;
  assign n13918 = ~n13916 & ~n13917;
  assign n13919 = ~n13913 & ~n13918;
  assign n13920 = ~n13912 & ~n13919;
  assign n13921 = po26  & ~n13920;
  assign n13922 = ~po26  & n13920;
  assign n13923 = ~n13413 & ~n13414;
  assign n13924 = po9  & n13923;
  assign n13925 = ~n13419 & ~n13924;
  assign n13926 = n13419 & n13924;
  assign n13927 = ~n13925 & ~n13926;
  assign n13928 = ~n13922 & ~n13927;
  assign n13929 = ~n13921 & ~n13928;
  assign n13930 = po27  & ~n13929;
  assign n13931 = ~po27  & n13929;
  assign n13932 = ~n13422 & ~n13423;
  assign n13933 = po9  & n13932;
  assign n13934 = ~n13428 & ~n13933;
  assign n13935 = n13428 & n13933;
  assign n13936 = ~n13934 & ~n13935;
  assign n13937 = ~n13931 & ~n13936;
  assign n13938 = ~n13930 & ~n13937;
  assign n13939 = po28  & ~n13938;
  assign n13940 = ~po28  & n13938;
  assign n13941 = ~n13431 & ~n13432;
  assign n13942 = po9  & n13941;
  assign n13943 = ~n13437 & ~n13942;
  assign n13944 = n13437 & n13942;
  assign n13945 = ~n13943 & ~n13944;
  assign n13946 = ~n13940 & ~n13945;
  assign n13947 = ~n13939 & ~n13946;
  assign n13948 = po29  & ~n13947;
  assign n13949 = ~po29  & n13947;
  assign n13950 = ~n13440 & ~n13441;
  assign n13951 = po9  & n13950;
  assign n13952 = ~n13446 & ~n13951;
  assign n13953 = n13446 & n13951;
  assign n13954 = ~n13952 & ~n13953;
  assign n13955 = ~n13949 & ~n13954;
  assign n13956 = ~n13948 & ~n13955;
  assign n13957 = po30  & ~n13956;
  assign n13958 = ~po30  & n13956;
  assign n13959 = ~n13449 & ~n13450;
  assign n13960 = po9  & n13959;
  assign n13961 = ~n13455 & ~n13960;
  assign n13962 = n13455 & n13960;
  assign n13963 = ~n13961 & ~n13962;
  assign n13964 = ~n13958 & ~n13963;
  assign n13965 = ~n13957 & ~n13964;
  assign n13966 = po31  & ~n13965;
  assign n13967 = ~po31  & n13965;
  assign n13968 = ~n13458 & ~n13459;
  assign n13969 = po9  & n13968;
  assign n13970 = ~n13464 & ~n13969;
  assign n13971 = n13464 & n13969;
  assign n13972 = ~n13970 & ~n13971;
  assign n13973 = ~n13967 & ~n13972;
  assign n13974 = ~n13966 & ~n13973;
  assign n13975 = po32  & ~n13974;
  assign n13976 = ~po32  & n13974;
  assign n13977 = ~n13467 & ~n13468;
  assign n13978 = po9  & n13977;
  assign n13979 = ~n13473 & ~n13978;
  assign n13980 = n13473 & n13978;
  assign n13981 = ~n13979 & ~n13980;
  assign n13982 = ~n13976 & ~n13981;
  assign n13983 = ~n13975 & ~n13982;
  assign n13984 = po33  & ~n13983;
  assign n13985 = ~po33  & n13983;
  assign n13986 = ~n13476 & ~n13477;
  assign n13987 = po9  & n13986;
  assign n13988 = ~n13482 & ~n13987;
  assign n13989 = n13482 & n13987;
  assign n13990 = ~n13988 & ~n13989;
  assign n13991 = ~n13985 & ~n13990;
  assign n13992 = ~n13984 & ~n13991;
  assign n13993 = po34  & ~n13992;
  assign n13994 = ~po34  & n13992;
  assign n13995 = ~n13485 & ~n13486;
  assign n13996 = po9  & n13995;
  assign n13997 = ~n13491 & ~n13996;
  assign n13998 = n13491 & n13996;
  assign n13999 = ~n13997 & ~n13998;
  assign n14000 = ~n13994 & ~n13999;
  assign n14001 = ~n13993 & ~n14000;
  assign n14002 = po35  & ~n14001;
  assign n14003 = ~po35  & n14001;
  assign n14004 = ~n13494 & ~n13495;
  assign n14005 = po9  & n14004;
  assign n14006 = ~n13500 & ~n14005;
  assign n14007 = n13500 & n14005;
  assign n14008 = ~n14006 & ~n14007;
  assign n14009 = ~n14003 & ~n14008;
  assign n14010 = ~n14002 & ~n14009;
  assign n14011 = po36  & ~n14010;
  assign n14012 = ~po36  & n14010;
  assign n14013 = ~n13503 & ~n13504;
  assign n14014 = po9  & n14013;
  assign n14015 = ~n13509 & ~n14014;
  assign n14016 = n13509 & n14014;
  assign n14017 = ~n14015 & ~n14016;
  assign n14018 = ~n14012 & ~n14017;
  assign n14019 = ~n14011 & ~n14018;
  assign n14020 = po37  & ~n14019;
  assign n14021 = ~po37  & n14019;
  assign n14022 = ~n13512 & ~n13513;
  assign n14023 = po9  & n14022;
  assign n14024 = ~n13518 & ~n14023;
  assign n14025 = n13518 & n14023;
  assign n14026 = ~n14024 & ~n14025;
  assign n14027 = ~n14021 & ~n14026;
  assign n14028 = ~n14020 & ~n14027;
  assign n14029 = po38  & ~n14028;
  assign n14030 = ~po38  & n14028;
  assign n14031 = ~n13521 & ~n13522;
  assign n14032 = po9  & n14031;
  assign n14033 = ~n13527 & ~n14032;
  assign n14034 = n13527 & n14032;
  assign n14035 = ~n14033 & ~n14034;
  assign n14036 = ~n14030 & ~n14035;
  assign n14037 = ~n14029 & ~n14036;
  assign n14038 = po39  & ~n14037;
  assign n14039 = ~po39  & n14037;
  assign n14040 = ~n13530 & ~n13531;
  assign n14041 = po9  & n14040;
  assign n14042 = ~n13536 & ~n14041;
  assign n14043 = n13536 & n14041;
  assign n14044 = ~n14042 & ~n14043;
  assign n14045 = ~n14039 & ~n14044;
  assign n14046 = ~n14038 & ~n14045;
  assign n14047 = po40  & ~n14046;
  assign n14048 = ~po40  & n14046;
  assign n14049 = ~n13539 & ~n13540;
  assign n14050 = po9  & n14049;
  assign n14051 = ~n13545 & ~n14050;
  assign n14052 = n13545 & n14050;
  assign n14053 = ~n14051 & ~n14052;
  assign n14054 = ~n14048 & ~n14053;
  assign n14055 = ~n14047 & ~n14054;
  assign n14056 = po41  & ~n14055;
  assign n14057 = ~po41  & n14055;
  assign n14058 = ~n13548 & ~n13549;
  assign n14059 = po9  & n14058;
  assign n14060 = ~n13554 & ~n14059;
  assign n14061 = n13554 & n14059;
  assign n14062 = ~n14060 & ~n14061;
  assign n14063 = ~n14057 & ~n14062;
  assign n14064 = ~n14056 & ~n14063;
  assign n14065 = po42  & ~n14064;
  assign n14066 = ~po42  & n14064;
  assign n14067 = ~n13557 & ~n13558;
  assign n14068 = po9  & n14067;
  assign n14069 = ~n13563 & ~n14068;
  assign n14070 = n13563 & n14068;
  assign n14071 = ~n14069 & ~n14070;
  assign n14072 = ~n14066 & ~n14071;
  assign n14073 = ~n14065 & ~n14072;
  assign n14074 = po43  & ~n14073;
  assign n14075 = ~po43  & n14073;
  assign n14076 = ~n13566 & ~n13567;
  assign n14077 = po9  & n14076;
  assign n14078 = ~n13572 & ~n14077;
  assign n14079 = n13572 & n14077;
  assign n14080 = ~n14078 & ~n14079;
  assign n14081 = ~n14075 & ~n14080;
  assign n14082 = ~n14074 & ~n14081;
  assign n14083 = po44  & ~n14082;
  assign n14084 = ~po44  & n14082;
  assign n14085 = ~n13575 & ~n13576;
  assign n14086 = po9  & n14085;
  assign n14087 = ~n13581 & ~n14086;
  assign n14088 = n13581 & n14086;
  assign n14089 = ~n14087 & ~n14088;
  assign n14090 = ~n14084 & ~n14089;
  assign n14091 = ~n14083 & ~n14090;
  assign n14092 = po45  & ~n14091;
  assign n14093 = ~po45  & n14091;
  assign n14094 = ~n13584 & ~n13585;
  assign n14095 = po9  & n14094;
  assign n14096 = ~n13590 & ~n14095;
  assign n14097 = n13590 & n14095;
  assign n14098 = ~n14096 & ~n14097;
  assign n14099 = ~n14093 & ~n14098;
  assign n14100 = ~n14092 & ~n14099;
  assign n14101 = po46  & ~n14100;
  assign n14102 = ~po46  & n14100;
  assign n14103 = ~n13593 & ~n13594;
  assign n14104 = po9  & n14103;
  assign n14105 = ~n13599 & ~n14104;
  assign n14106 = n13599 & n14104;
  assign n14107 = ~n14105 & ~n14106;
  assign n14108 = ~n14102 & ~n14107;
  assign n14109 = ~n14101 & ~n14108;
  assign n14110 = po47  & ~n14109;
  assign n14111 = ~po47  & n14109;
  assign n14112 = ~n13602 & ~n13603;
  assign n14113 = po9  & n14112;
  assign n14114 = ~n13608 & ~n14113;
  assign n14115 = n13608 & n14113;
  assign n14116 = ~n14114 & ~n14115;
  assign n14117 = ~n14111 & ~n14116;
  assign n14118 = ~n14110 & ~n14117;
  assign n14119 = po48  & ~n14118;
  assign n14120 = ~po48  & n14118;
  assign n14121 = ~n13611 & ~n13612;
  assign n14122 = po9  & n14121;
  assign n14123 = ~n13617 & ~n14122;
  assign n14124 = n13617 & n14122;
  assign n14125 = ~n14123 & ~n14124;
  assign n14126 = ~n14120 & ~n14125;
  assign n14127 = ~n14119 & ~n14126;
  assign n14128 = po49  & ~n14127;
  assign n14129 = ~po49  & n14127;
  assign n14130 = ~n13620 & ~n13621;
  assign n14131 = po9  & n14130;
  assign n14132 = ~n13626 & ~n14131;
  assign n14133 = n13626 & n14131;
  assign n14134 = ~n14132 & ~n14133;
  assign n14135 = ~n14129 & ~n14134;
  assign n14136 = ~n14128 & ~n14135;
  assign n14137 = po50  & ~n14136;
  assign n14138 = ~po50  & n14136;
  assign n14139 = ~n13629 & ~n13630;
  assign n14140 = po9  & n14139;
  assign n14141 = ~n13635 & ~n14140;
  assign n14142 = n13635 & n14140;
  assign n14143 = ~n14141 & ~n14142;
  assign n14144 = ~n14138 & ~n14143;
  assign n14145 = ~n14137 & ~n14144;
  assign n14146 = po51  & ~n14145;
  assign n14147 = ~po51  & n14145;
  assign n14148 = ~n13638 & ~n13639;
  assign n14149 = po9  & n14148;
  assign n14150 = ~n13644 & ~n14149;
  assign n14151 = n13644 & n14149;
  assign n14152 = ~n14150 & ~n14151;
  assign n14153 = ~n14147 & ~n14152;
  assign n14154 = ~n14146 & ~n14153;
  assign n14155 = po52  & ~n14154;
  assign n14156 = ~po52  & n14154;
  assign n14157 = ~n13647 & ~n13648;
  assign n14158 = po9  & n14157;
  assign n14159 = ~n13653 & ~n14158;
  assign n14160 = n13653 & n14158;
  assign n14161 = ~n14159 & ~n14160;
  assign n14162 = ~n14156 & ~n14161;
  assign n14163 = ~n14155 & ~n14162;
  assign n14164 = po53  & ~n14163;
  assign n14165 = ~po53  & n14163;
  assign n14166 = ~n13656 & ~n13657;
  assign n14167 = po9  & n14166;
  assign n14168 = ~n13662 & ~n14167;
  assign n14169 = n13662 & n14167;
  assign n14170 = ~n14168 & ~n14169;
  assign n14171 = ~n14165 & ~n14170;
  assign n14172 = ~n14164 & ~n14171;
  assign n14173 = po54  & ~n14172;
  assign n14174 = ~po54  & n14172;
  assign n14175 = ~n13665 & ~n13666;
  assign n14176 = po9  & n14175;
  assign n14177 = ~n13671 & ~n14176;
  assign n14178 = n13671 & n14176;
  assign n14179 = ~n14177 & ~n14178;
  assign n14180 = ~n14174 & ~n14179;
  assign n14181 = ~n14173 & ~n14180;
  assign n14182 = po55  & ~n14181;
  assign n14183 = ~n13674 & ~n13680;
  assign n14184 = po9  & n14183;
  assign n14185 = ~n13679 & ~n14184;
  assign n14186 = n13679 & n14184;
  assign n14187 = ~n14185 & ~n14186;
  assign n14188 = ~po55  & n14181;
  assign n14189 = ~n14187 & ~n14188;
  assign n14190 = ~n14182 & ~n14189;
  assign n14191 = po56  & ~n14190;
  assign n14192 = ~po56  & n14190;
  assign n14193 = ~n13763 & ~n14192;
  assign n14194 = ~n14191 & ~n14193;
  assign n14195 = po57  & ~n14194;
  assign n14196 = ~po57  & n14194;
  assign n14197 = ~n13687 & ~n13688;
  assign n14198 = po9  & n14197;
  assign n14199 = ~n13693 & ~n14198;
  assign n14200 = n13693 & n14198;
  assign n14201 = ~n14199 & ~n14200;
  assign n14202 = ~n14196 & ~n14201;
  assign n14203 = ~n14195 & ~n14202;
  assign n14204 = po58  & ~n14203;
  assign n14205 = ~po58  & n14203;
  assign n14206 = ~n13696 & ~n13697;
  assign n14207 = po9  & n14206;
  assign n14208 = ~n13702 & ~n14207;
  assign n14209 = n13702 & n14207;
  assign n14210 = ~n14208 & ~n14209;
  assign n14211 = ~n14205 & ~n14210;
  assign n14212 = ~n14204 & ~n14211;
  assign n14213 = po59  & ~n14212;
  assign n14214 = ~po59  & n14212;
  assign n14215 = ~n13705 & ~n13706;
  assign n14216 = po9  & n14215;
  assign n14217 = ~n13711 & ~n14216;
  assign n14218 = n13711 & n14216;
  assign n14219 = ~n14217 & ~n14218;
  assign n14220 = ~n14214 & ~n14219;
  assign n14221 = ~n14213 & ~n14220;
  assign n14222 = po60  & ~n14221;
  assign n14223 = ~po60  & n14221;
  assign n14224 = ~n13714 & ~n13715;
  assign n14225 = po9  & n14224;
  assign n14226 = ~n13720 & ~n14225;
  assign n14227 = n13720 & n14225;
  assign n14228 = ~n14226 & ~n14227;
  assign n14229 = ~n14223 & ~n14228;
  assign n14230 = ~n14222 & ~n14229;
  assign n14231 = po61  & ~n14230;
  assign n14232 = ~po61  & n14230;
  assign n14233 = ~n13723 & ~n13724;
  assign n14234 = po9  & n14233;
  assign n14235 = ~n13729 & ~n14234;
  assign n14236 = n13729 & n14234;
  assign n14237 = ~n14235 & ~n14236;
  assign n14238 = ~n14232 & ~n14237;
  assign n14239 = ~n14231 & ~n14238;
  assign n14240 = po62  & ~n14239;
  assign n14241 = ~po62  & n14239;
  assign n14242 = ~n13732 & ~n13733;
  assign n14243 = po9  & n14242;
  assign n14244 = ~n13738 & ~n14243;
  assign n14245 = n13738 & n14243;
  assign n14246 = ~n14244 & ~n14245;
  assign n14247 = ~n14241 & ~n14246;
  assign n14248 = ~n14240 & ~n14247;
  assign n14249 = n13773 & n14248;
  assign n14250 = ~n13773 & ~n14248;
  assign n14251 = n13751 & po9 ;
  assign n14252 = ~n13750 & ~n14251;
  assign n14253 = n14250 & n14252;
  assign n14254 = ~po63  & ~n14253;
  assign n14255 = ~n14249 & ~n14254;
  assign n14256 = ~n13768 & n14255;
  assign po8  = n13764 | ~n14256;
  assign n14258 = ~n14191 & ~n14192;
  assign n14259 = po8  & n14258;
  assign n14260 = ~n13763 & ~n14259;
  assign n14261 = n13763 & n14259;
  assign n14262 = ~n14260 & ~n14261;
  assign n14263 = n13773 & ~po8 ;
  assign n14264 = ~n13773 & po8 ;
  assign n14265 = n14248 & ~n14264;
  assign n14266 = po63  & ~n14265;
  assign n14267 = ~n14250 & n14266;
  assign n14268 = ~n14240 & ~n14241;
  assign n14269 = po8  & n14268;
  assign n14270 = ~n14246 & ~n14269;
  assign n14271 = n14246 & n14269;
  assign n14272 = ~n14270 & ~n14271;
  assign n14273 = pi16  & po8 ;
  assign n14274 = ~pi14  & ~pi15 ;
  assign n14275 = ~pi16  & n14274;
  assign n14276 = ~n14273 & ~n14275;
  assign n14277 = po9  & ~n14276;
  assign n14278 = ~po9  & n14276;
  assign n14279 = ~pi16  & po8 ;
  assign n14280 = pi17  & ~n14279;
  assign n14281 = n13775 & po8 ;
  assign n14282 = ~n14280 & ~n14281;
  assign n14283 = ~n14278 & n14282;
  assign n14284 = ~n14277 & ~n14283;
  assign n14285 = po10  & ~n14284;
  assign n14286 = ~po10  & n14284;
  assign n14287 = po9  & n14256;
  assign n14288 = ~n14281 & ~n14287;
  assign n14289 = pi18  & ~n14288;
  assign n14290 = ~pi18  & n14288;
  assign n14291 = ~n14289 & ~n14290;
  assign n14292 = ~n14286 & ~n14291;
  assign n14293 = ~n14285 & ~n14292;
  assign n14294 = po11  & ~n14293;
  assign n14295 = ~po11  & n14293;
  assign n14296 = ~n13778 & ~n13779;
  assign n14297 = po8  & n14296;
  assign n14298 = n13783 & ~n14297;
  assign n14299 = ~n13783 & n14297;
  assign n14300 = ~n14298 & ~n14299;
  assign n14301 = ~n14295 & ~n14300;
  assign n14302 = ~n14294 & ~n14301;
  assign n14303 = po12  & ~n14302;
  assign n14304 = ~po12  & n14302;
  assign n14305 = ~n13786 & ~n13787;
  assign n14306 = po8  & n14305;
  assign n14307 = ~n13792 & ~n14306;
  assign n14308 = n13792 & n14306;
  assign n14309 = ~n14307 & ~n14308;
  assign n14310 = ~n14304 & ~n14309;
  assign n14311 = ~n14303 & ~n14310;
  assign n14312 = po13  & ~n14311;
  assign n14313 = ~po13  & n14311;
  assign n14314 = ~n13795 & ~n13796;
  assign n14315 = po8  & n14314;
  assign n14316 = n13801 & n14315;
  assign n14317 = ~n13801 & ~n14315;
  assign n14318 = ~n14316 & ~n14317;
  assign n14319 = ~n14313 & ~n14318;
  assign n14320 = ~n14312 & ~n14319;
  assign n14321 = po14  & ~n14320;
  assign n14322 = ~po14  & n14320;
  assign n14323 = ~n13804 & ~n13805;
  assign n14324 = po8  & n14323;
  assign n14325 = ~n13810 & ~n14324;
  assign n14326 = n13810 & n14324;
  assign n14327 = ~n14325 & ~n14326;
  assign n14328 = ~n14322 & ~n14327;
  assign n14329 = ~n14321 & ~n14328;
  assign n14330 = po15  & ~n14329;
  assign n14331 = ~po15  & n14329;
  assign n14332 = ~n13813 & ~n13814;
  assign n14333 = po8  & n14332;
  assign n14334 = ~n13819 & ~n14333;
  assign n14335 = n13819 & n14333;
  assign n14336 = ~n14334 & ~n14335;
  assign n14337 = ~n14331 & ~n14336;
  assign n14338 = ~n14330 & ~n14337;
  assign n14339 = po16  & ~n14338;
  assign n14340 = ~po16  & n14338;
  assign n14341 = ~n13822 & ~n13823;
  assign n14342 = po8  & n14341;
  assign n14343 = ~n13828 & ~n14342;
  assign n14344 = n13828 & n14342;
  assign n14345 = ~n14343 & ~n14344;
  assign n14346 = ~n14340 & ~n14345;
  assign n14347 = ~n14339 & ~n14346;
  assign n14348 = po17  & ~n14347;
  assign n14349 = ~po17  & n14347;
  assign n14350 = ~n13831 & ~n13832;
  assign n14351 = po8  & n14350;
  assign n14352 = ~n13837 & ~n14351;
  assign n14353 = n13837 & n14351;
  assign n14354 = ~n14352 & ~n14353;
  assign n14355 = ~n14349 & ~n14354;
  assign n14356 = ~n14348 & ~n14355;
  assign n14357 = po18  & ~n14356;
  assign n14358 = ~po18  & n14356;
  assign n14359 = ~n13840 & ~n13841;
  assign n14360 = po8  & n14359;
  assign n14361 = ~n13846 & ~n14360;
  assign n14362 = n13846 & n14360;
  assign n14363 = ~n14361 & ~n14362;
  assign n14364 = ~n14358 & ~n14363;
  assign n14365 = ~n14357 & ~n14364;
  assign n14366 = po19  & ~n14365;
  assign n14367 = ~po19  & n14365;
  assign n14368 = ~n13849 & ~n13850;
  assign n14369 = po8  & n14368;
  assign n14370 = ~n13855 & ~n14369;
  assign n14371 = n13855 & n14369;
  assign n14372 = ~n14370 & ~n14371;
  assign n14373 = ~n14367 & ~n14372;
  assign n14374 = ~n14366 & ~n14373;
  assign n14375 = po20  & ~n14374;
  assign n14376 = ~po20  & n14374;
  assign n14377 = ~n13858 & ~n13859;
  assign n14378 = po8  & n14377;
  assign n14379 = ~n13864 & ~n14378;
  assign n14380 = n13864 & n14378;
  assign n14381 = ~n14379 & ~n14380;
  assign n14382 = ~n14376 & ~n14381;
  assign n14383 = ~n14375 & ~n14382;
  assign n14384 = po21  & ~n14383;
  assign n14385 = ~po21  & n14383;
  assign n14386 = ~n13867 & ~n13868;
  assign n14387 = po8  & n14386;
  assign n14388 = ~n13873 & ~n14387;
  assign n14389 = n13873 & n14387;
  assign n14390 = ~n14388 & ~n14389;
  assign n14391 = ~n14385 & ~n14390;
  assign n14392 = ~n14384 & ~n14391;
  assign n14393 = po22  & ~n14392;
  assign n14394 = ~po22  & n14392;
  assign n14395 = ~n13876 & ~n13877;
  assign n14396 = po8  & n14395;
  assign n14397 = ~n13882 & ~n14396;
  assign n14398 = n13882 & n14396;
  assign n14399 = ~n14397 & ~n14398;
  assign n14400 = ~n14394 & ~n14399;
  assign n14401 = ~n14393 & ~n14400;
  assign n14402 = po23  & ~n14401;
  assign n14403 = ~po23  & n14401;
  assign n14404 = ~n13885 & ~n13886;
  assign n14405 = po8  & n14404;
  assign n14406 = ~n13891 & ~n14405;
  assign n14407 = n13891 & n14405;
  assign n14408 = ~n14406 & ~n14407;
  assign n14409 = ~n14403 & ~n14408;
  assign n14410 = ~n14402 & ~n14409;
  assign n14411 = po24  & ~n14410;
  assign n14412 = ~po24  & n14410;
  assign n14413 = ~n13894 & ~n13895;
  assign n14414 = po8  & n14413;
  assign n14415 = ~n13900 & ~n14414;
  assign n14416 = n13900 & n14414;
  assign n14417 = ~n14415 & ~n14416;
  assign n14418 = ~n14412 & ~n14417;
  assign n14419 = ~n14411 & ~n14418;
  assign n14420 = po25  & ~n14419;
  assign n14421 = ~po25  & n14419;
  assign n14422 = ~n13903 & ~n13904;
  assign n14423 = po8  & n14422;
  assign n14424 = ~n13909 & ~n14423;
  assign n14425 = n13909 & n14423;
  assign n14426 = ~n14424 & ~n14425;
  assign n14427 = ~n14421 & ~n14426;
  assign n14428 = ~n14420 & ~n14427;
  assign n14429 = po26  & ~n14428;
  assign n14430 = ~po26  & n14428;
  assign n14431 = ~n13912 & ~n13913;
  assign n14432 = po8  & n14431;
  assign n14433 = ~n13918 & ~n14432;
  assign n14434 = n13918 & n14432;
  assign n14435 = ~n14433 & ~n14434;
  assign n14436 = ~n14430 & ~n14435;
  assign n14437 = ~n14429 & ~n14436;
  assign n14438 = po27  & ~n14437;
  assign n14439 = ~po27  & n14437;
  assign n14440 = ~n13921 & ~n13922;
  assign n14441 = po8  & n14440;
  assign n14442 = ~n13927 & ~n14441;
  assign n14443 = n13927 & n14441;
  assign n14444 = ~n14442 & ~n14443;
  assign n14445 = ~n14439 & ~n14444;
  assign n14446 = ~n14438 & ~n14445;
  assign n14447 = po28  & ~n14446;
  assign n14448 = ~po28  & n14446;
  assign n14449 = ~n13930 & ~n13931;
  assign n14450 = po8  & n14449;
  assign n14451 = ~n13936 & ~n14450;
  assign n14452 = n13936 & n14450;
  assign n14453 = ~n14451 & ~n14452;
  assign n14454 = ~n14448 & ~n14453;
  assign n14455 = ~n14447 & ~n14454;
  assign n14456 = po29  & ~n14455;
  assign n14457 = ~po29  & n14455;
  assign n14458 = ~n13939 & ~n13940;
  assign n14459 = po8  & n14458;
  assign n14460 = ~n13945 & ~n14459;
  assign n14461 = n13945 & n14459;
  assign n14462 = ~n14460 & ~n14461;
  assign n14463 = ~n14457 & ~n14462;
  assign n14464 = ~n14456 & ~n14463;
  assign n14465 = po30  & ~n14464;
  assign n14466 = ~po30  & n14464;
  assign n14467 = ~n13948 & ~n13949;
  assign n14468 = po8  & n14467;
  assign n14469 = ~n13954 & ~n14468;
  assign n14470 = n13954 & n14468;
  assign n14471 = ~n14469 & ~n14470;
  assign n14472 = ~n14466 & ~n14471;
  assign n14473 = ~n14465 & ~n14472;
  assign n14474 = po31  & ~n14473;
  assign n14475 = ~po31  & n14473;
  assign n14476 = ~n13957 & ~n13958;
  assign n14477 = po8  & n14476;
  assign n14478 = ~n13963 & ~n14477;
  assign n14479 = n13963 & n14477;
  assign n14480 = ~n14478 & ~n14479;
  assign n14481 = ~n14475 & ~n14480;
  assign n14482 = ~n14474 & ~n14481;
  assign n14483 = po32  & ~n14482;
  assign n14484 = ~po32  & n14482;
  assign n14485 = ~n13966 & ~n13967;
  assign n14486 = po8  & n14485;
  assign n14487 = ~n13972 & ~n14486;
  assign n14488 = n13972 & n14486;
  assign n14489 = ~n14487 & ~n14488;
  assign n14490 = ~n14484 & ~n14489;
  assign n14491 = ~n14483 & ~n14490;
  assign n14492 = po33  & ~n14491;
  assign n14493 = ~po33  & n14491;
  assign n14494 = ~n13975 & ~n13976;
  assign n14495 = po8  & n14494;
  assign n14496 = ~n13981 & ~n14495;
  assign n14497 = n13981 & n14495;
  assign n14498 = ~n14496 & ~n14497;
  assign n14499 = ~n14493 & ~n14498;
  assign n14500 = ~n14492 & ~n14499;
  assign n14501 = po34  & ~n14500;
  assign n14502 = ~po34  & n14500;
  assign n14503 = ~n13984 & ~n13985;
  assign n14504 = po8  & n14503;
  assign n14505 = ~n13990 & ~n14504;
  assign n14506 = n13990 & n14504;
  assign n14507 = ~n14505 & ~n14506;
  assign n14508 = ~n14502 & ~n14507;
  assign n14509 = ~n14501 & ~n14508;
  assign n14510 = po35  & ~n14509;
  assign n14511 = ~po35  & n14509;
  assign n14512 = ~n13993 & ~n13994;
  assign n14513 = po8  & n14512;
  assign n14514 = ~n13999 & ~n14513;
  assign n14515 = n13999 & n14513;
  assign n14516 = ~n14514 & ~n14515;
  assign n14517 = ~n14511 & ~n14516;
  assign n14518 = ~n14510 & ~n14517;
  assign n14519 = po36  & ~n14518;
  assign n14520 = ~po36  & n14518;
  assign n14521 = ~n14002 & ~n14003;
  assign n14522 = po8  & n14521;
  assign n14523 = ~n14008 & ~n14522;
  assign n14524 = n14008 & n14522;
  assign n14525 = ~n14523 & ~n14524;
  assign n14526 = ~n14520 & ~n14525;
  assign n14527 = ~n14519 & ~n14526;
  assign n14528 = po37  & ~n14527;
  assign n14529 = ~po37  & n14527;
  assign n14530 = ~n14011 & ~n14012;
  assign n14531 = po8  & n14530;
  assign n14532 = ~n14017 & ~n14531;
  assign n14533 = n14017 & n14531;
  assign n14534 = ~n14532 & ~n14533;
  assign n14535 = ~n14529 & ~n14534;
  assign n14536 = ~n14528 & ~n14535;
  assign n14537 = po38  & ~n14536;
  assign n14538 = ~po38  & n14536;
  assign n14539 = ~n14020 & ~n14021;
  assign n14540 = po8  & n14539;
  assign n14541 = ~n14026 & ~n14540;
  assign n14542 = n14026 & n14540;
  assign n14543 = ~n14541 & ~n14542;
  assign n14544 = ~n14538 & ~n14543;
  assign n14545 = ~n14537 & ~n14544;
  assign n14546 = po39  & ~n14545;
  assign n14547 = ~po39  & n14545;
  assign n14548 = ~n14029 & ~n14030;
  assign n14549 = po8  & n14548;
  assign n14550 = ~n14035 & ~n14549;
  assign n14551 = n14035 & n14549;
  assign n14552 = ~n14550 & ~n14551;
  assign n14553 = ~n14547 & ~n14552;
  assign n14554 = ~n14546 & ~n14553;
  assign n14555 = po40  & ~n14554;
  assign n14556 = ~po40  & n14554;
  assign n14557 = ~n14038 & ~n14039;
  assign n14558 = po8  & n14557;
  assign n14559 = ~n14044 & ~n14558;
  assign n14560 = n14044 & n14558;
  assign n14561 = ~n14559 & ~n14560;
  assign n14562 = ~n14556 & ~n14561;
  assign n14563 = ~n14555 & ~n14562;
  assign n14564 = po41  & ~n14563;
  assign n14565 = ~po41  & n14563;
  assign n14566 = ~n14047 & ~n14048;
  assign n14567 = po8  & n14566;
  assign n14568 = ~n14053 & ~n14567;
  assign n14569 = n14053 & n14567;
  assign n14570 = ~n14568 & ~n14569;
  assign n14571 = ~n14565 & ~n14570;
  assign n14572 = ~n14564 & ~n14571;
  assign n14573 = po42  & ~n14572;
  assign n14574 = ~po42  & n14572;
  assign n14575 = ~n14056 & ~n14057;
  assign n14576 = po8  & n14575;
  assign n14577 = ~n14062 & ~n14576;
  assign n14578 = n14062 & n14576;
  assign n14579 = ~n14577 & ~n14578;
  assign n14580 = ~n14574 & ~n14579;
  assign n14581 = ~n14573 & ~n14580;
  assign n14582 = po43  & ~n14581;
  assign n14583 = ~po43  & n14581;
  assign n14584 = ~n14065 & ~n14066;
  assign n14585 = po8  & n14584;
  assign n14586 = ~n14071 & ~n14585;
  assign n14587 = n14071 & n14585;
  assign n14588 = ~n14586 & ~n14587;
  assign n14589 = ~n14583 & ~n14588;
  assign n14590 = ~n14582 & ~n14589;
  assign n14591 = po44  & ~n14590;
  assign n14592 = ~po44  & n14590;
  assign n14593 = ~n14074 & ~n14075;
  assign n14594 = po8  & n14593;
  assign n14595 = ~n14080 & ~n14594;
  assign n14596 = n14080 & n14594;
  assign n14597 = ~n14595 & ~n14596;
  assign n14598 = ~n14592 & ~n14597;
  assign n14599 = ~n14591 & ~n14598;
  assign n14600 = po45  & ~n14599;
  assign n14601 = ~po45  & n14599;
  assign n14602 = ~n14083 & ~n14084;
  assign n14603 = po8  & n14602;
  assign n14604 = ~n14089 & ~n14603;
  assign n14605 = n14089 & n14603;
  assign n14606 = ~n14604 & ~n14605;
  assign n14607 = ~n14601 & ~n14606;
  assign n14608 = ~n14600 & ~n14607;
  assign n14609 = po46  & ~n14608;
  assign n14610 = ~po46  & n14608;
  assign n14611 = ~n14092 & ~n14093;
  assign n14612 = po8  & n14611;
  assign n14613 = ~n14098 & ~n14612;
  assign n14614 = n14098 & n14612;
  assign n14615 = ~n14613 & ~n14614;
  assign n14616 = ~n14610 & ~n14615;
  assign n14617 = ~n14609 & ~n14616;
  assign n14618 = po47  & ~n14617;
  assign n14619 = ~po47  & n14617;
  assign n14620 = ~n14101 & ~n14102;
  assign n14621 = po8  & n14620;
  assign n14622 = ~n14107 & ~n14621;
  assign n14623 = n14107 & n14621;
  assign n14624 = ~n14622 & ~n14623;
  assign n14625 = ~n14619 & ~n14624;
  assign n14626 = ~n14618 & ~n14625;
  assign n14627 = po48  & ~n14626;
  assign n14628 = ~po48  & n14626;
  assign n14629 = ~n14110 & ~n14111;
  assign n14630 = po8  & n14629;
  assign n14631 = ~n14116 & ~n14630;
  assign n14632 = n14116 & n14630;
  assign n14633 = ~n14631 & ~n14632;
  assign n14634 = ~n14628 & ~n14633;
  assign n14635 = ~n14627 & ~n14634;
  assign n14636 = po49  & ~n14635;
  assign n14637 = ~po49  & n14635;
  assign n14638 = ~n14119 & ~n14120;
  assign n14639 = po8  & n14638;
  assign n14640 = ~n14125 & ~n14639;
  assign n14641 = n14125 & n14639;
  assign n14642 = ~n14640 & ~n14641;
  assign n14643 = ~n14637 & ~n14642;
  assign n14644 = ~n14636 & ~n14643;
  assign n14645 = po50  & ~n14644;
  assign n14646 = ~po50  & n14644;
  assign n14647 = ~n14128 & ~n14129;
  assign n14648 = po8  & n14647;
  assign n14649 = ~n14134 & ~n14648;
  assign n14650 = n14134 & n14648;
  assign n14651 = ~n14649 & ~n14650;
  assign n14652 = ~n14646 & ~n14651;
  assign n14653 = ~n14645 & ~n14652;
  assign n14654 = po51  & ~n14653;
  assign n14655 = ~po51  & n14653;
  assign n14656 = ~n14137 & ~n14138;
  assign n14657 = po8  & n14656;
  assign n14658 = ~n14143 & ~n14657;
  assign n14659 = n14143 & n14657;
  assign n14660 = ~n14658 & ~n14659;
  assign n14661 = ~n14655 & ~n14660;
  assign n14662 = ~n14654 & ~n14661;
  assign n14663 = po52  & ~n14662;
  assign n14664 = ~po52  & n14662;
  assign n14665 = ~n14146 & ~n14147;
  assign n14666 = po8  & n14665;
  assign n14667 = ~n14152 & ~n14666;
  assign n14668 = n14152 & n14666;
  assign n14669 = ~n14667 & ~n14668;
  assign n14670 = ~n14664 & ~n14669;
  assign n14671 = ~n14663 & ~n14670;
  assign n14672 = po53  & ~n14671;
  assign n14673 = ~po53  & n14671;
  assign n14674 = ~n14155 & ~n14156;
  assign n14675 = po8  & n14674;
  assign n14676 = ~n14161 & ~n14675;
  assign n14677 = n14161 & n14675;
  assign n14678 = ~n14676 & ~n14677;
  assign n14679 = ~n14673 & ~n14678;
  assign n14680 = ~n14672 & ~n14679;
  assign n14681 = po54  & ~n14680;
  assign n14682 = ~po54  & n14680;
  assign n14683 = ~n14164 & ~n14165;
  assign n14684 = po8  & n14683;
  assign n14685 = ~n14170 & ~n14684;
  assign n14686 = n14170 & n14684;
  assign n14687 = ~n14685 & ~n14686;
  assign n14688 = ~n14682 & ~n14687;
  assign n14689 = ~n14681 & ~n14688;
  assign n14690 = po55  & ~n14689;
  assign n14691 = ~po55  & n14689;
  assign n14692 = ~n14173 & ~n14174;
  assign n14693 = po8  & n14692;
  assign n14694 = ~n14179 & ~n14693;
  assign n14695 = n14179 & n14693;
  assign n14696 = ~n14694 & ~n14695;
  assign n14697 = ~n14691 & ~n14696;
  assign n14698 = ~n14690 & ~n14697;
  assign n14699 = po56  & ~n14698;
  assign n14700 = ~n14182 & ~n14188;
  assign n14701 = po8  & n14700;
  assign n14702 = ~n14187 & ~n14701;
  assign n14703 = n14187 & n14701;
  assign n14704 = ~n14702 & ~n14703;
  assign n14705 = ~po56  & n14698;
  assign n14706 = ~n14704 & ~n14705;
  assign n14707 = ~n14699 & ~n14706;
  assign n14708 = po57  & ~n14707;
  assign n14709 = ~po57  & n14707;
  assign n14710 = ~n14262 & ~n14709;
  assign n14711 = ~n14708 & ~n14710;
  assign n14712 = po58  & ~n14711;
  assign n14713 = ~po58  & n14711;
  assign n14714 = ~n14195 & ~n14196;
  assign n14715 = po8  & n14714;
  assign n14716 = ~n14201 & ~n14715;
  assign n14717 = n14201 & n14715;
  assign n14718 = ~n14716 & ~n14717;
  assign n14719 = ~n14713 & ~n14718;
  assign n14720 = ~n14712 & ~n14719;
  assign n14721 = po59  & ~n14720;
  assign n14722 = ~po59  & n14720;
  assign n14723 = ~n14204 & ~n14205;
  assign n14724 = po8  & n14723;
  assign n14725 = ~n14210 & ~n14724;
  assign n14726 = n14210 & n14724;
  assign n14727 = ~n14725 & ~n14726;
  assign n14728 = ~n14722 & ~n14727;
  assign n14729 = ~n14721 & ~n14728;
  assign n14730 = po60  & ~n14729;
  assign n14731 = ~po60  & n14729;
  assign n14732 = ~n14213 & ~n14214;
  assign n14733 = po8  & n14732;
  assign n14734 = ~n14219 & ~n14733;
  assign n14735 = n14219 & n14733;
  assign n14736 = ~n14734 & ~n14735;
  assign n14737 = ~n14731 & ~n14736;
  assign n14738 = ~n14730 & ~n14737;
  assign n14739 = po61  & ~n14738;
  assign n14740 = ~po61  & n14738;
  assign n14741 = ~n14222 & ~n14223;
  assign n14742 = po8  & n14741;
  assign n14743 = ~n14228 & ~n14742;
  assign n14744 = n14228 & n14742;
  assign n14745 = ~n14743 & ~n14744;
  assign n14746 = ~n14740 & ~n14745;
  assign n14747 = ~n14739 & ~n14746;
  assign n14748 = po62  & ~n14747;
  assign n14749 = ~po62  & n14747;
  assign n14750 = ~n14231 & ~n14232;
  assign n14751 = po8  & n14750;
  assign n14752 = ~n14237 & ~n14751;
  assign n14753 = n14237 & n14751;
  assign n14754 = ~n14752 & ~n14753;
  assign n14755 = ~n14749 & ~n14754;
  assign n14756 = ~n14748 & ~n14755;
  assign n14757 = n14272 & n14756;
  assign n14758 = ~n14272 & ~n14756;
  assign n14759 = n14250 & po8 ;
  assign n14760 = ~n14249 & ~n14759;
  assign n14761 = n14758 & n14760;
  assign n14762 = ~po63  & ~n14761;
  assign n14763 = ~n14757 & ~n14762;
  assign n14764 = ~n14267 & n14763;
  assign po7  = n14263 | ~n14764;
  assign n14766 = ~n14708 & ~n14709;
  assign n14767 = po7  & n14766;
  assign n14768 = ~n14262 & ~n14767;
  assign n14769 = n14262 & n14767;
  assign n14770 = ~n14768 & ~n14769;
  assign n14771 = n14272 & ~po7 ;
  assign n14772 = ~n14272 & po7 ;
  assign n14773 = n14756 & ~n14772;
  assign n14774 = po63  & ~n14773;
  assign n14775 = ~n14758 & n14774;
  assign n14776 = ~n14748 & ~n14749;
  assign n14777 = po7  & n14776;
  assign n14778 = ~n14754 & ~n14777;
  assign n14779 = n14754 & n14777;
  assign n14780 = ~n14778 & ~n14779;
  assign n14781 = pi14  & po7 ;
  assign n14782 = ~pi12  & ~pi13 ;
  assign n14783 = ~pi14  & n14782;
  assign n14784 = ~n14781 & ~n14783;
  assign n14785 = po8  & ~n14784;
  assign n14786 = ~po8  & n14784;
  assign n14787 = ~pi14  & po7 ;
  assign n14788 = pi15  & ~n14787;
  assign n14789 = n14274 & po7 ;
  assign n14790 = ~n14788 & ~n14789;
  assign n14791 = ~n14786 & n14790;
  assign n14792 = ~n14785 & ~n14791;
  assign n14793 = po9  & ~n14792;
  assign n14794 = ~po9  & n14792;
  assign n14795 = po8  & n14764;
  assign n14796 = ~n14789 & ~n14795;
  assign n14797 = pi16  & ~n14796;
  assign n14798 = ~pi16  & n14796;
  assign n14799 = ~n14797 & ~n14798;
  assign n14800 = ~n14794 & ~n14799;
  assign n14801 = ~n14793 & ~n14800;
  assign n14802 = po10  & ~n14801;
  assign n14803 = ~po10  & n14801;
  assign n14804 = ~n14277 & ~n14278;
  assign n14805 = po7  & n14804;
  assign n14806 = n14282 & ~n14805;
  assign n14807 = ~n14282 & n14805;
  assign n14808 = ~n14806 & ~n14807;
  assign n14809 = ~n14803 & ~n14808;
  assign n14810 = ~n14802 & ~n14809;
  assign n14811 = po11  & ~n14810;
  assign n14812 = ~po11  & n14810;
  assign n14813 = ~n14285 & ~n14286;
  assign n14814 = po7  & n14813;
  assign n14815 = ~n14291 & ~n14814;
  assign n14816 = n14291 & n14814;
  assign n14817 = ~n14815 & ~n14816;
  assign n14818 = ~n14812 & ~n14817;
  assign n14819 = ~n14811 & ~n14818;
  assign n14820 = po12  & ~n14819;
  assign n14821 = ~po12  & n14819;
  assign n14822 = ~n14294 & ~n14295;
  assign n14823 = po7  & n14822;
  assign n14824 = n14300 & n14823;
  assign n14825 = ~n14300 & ~n14823;
  assign n14826 = ~n14824 & ~n14825;
  assign n14827 = ~n14821 & ~n14826;
  assign n14828 = ~n14820 & ~n14827;
  assign n14829 = po13  & ~n14828;
  assign n14830 = ~po13  & n14828;
  assign n14831 = ~n14303 & ~n14304;
  assign n14832 = po7  & n14831;
  assign n14833 = ~n14309 & ~n14832;
  assign n14834 = n14309 & n14832;
  assign n14835 = ~n14833 & ~n14834;
  assign n14836 = ~n14830 & ~n14835;
  assign n14837 = ~n14829 & ~n14836;
  assign n14838 = po14  & ~n14837;
  assign n14839 = ~po14  & n14837;
  assign n14840 = ~n14312 & ~n14313;
  assign n14841 = po7  & n14840;
  assign n14842 = ~n14318 & ~n14841;
  assign n14843 = n14318 & n14841;
  assign n14844 = ~n14842 & ~n14843;
  assign n14845 = ~n14839 & ~n14844;
  assign n14846 = ~n14838 & ~n14845;
  assign n14847 = po15  & ~n14846;
  assign n14848 = ~po15  & n14846;
  assign n14849 = ~n14321 & ~n14322;
  assign n14850 = po7  & n14849;
  assign n14851 = ~n14327 & ~n14850;
  assign n14852 = n14327 & n14850;
  assign n14853 = ~n14851 & ~n14852;
  assign n14854 = ~n14848 & ~n14853;
  assign n14855 = ~n14847 & ~n14854;
  assign n14856 = po16  & ~n14855;
  assign n14857 = ~po16  & n14855;
  assign n14858 = ~n14330 & ~n14331;
  assign n14859 = po7  & n14858;
  assign n14860 = ~n14336 & ~n14859;
  assign n14861 = n14336 & n14859;
  assign n14862 = ~n14860 & ~n14861;
  assign n14863 = ~n14857 & ~n14862;
  assign n14864 = ~n14856 & ~n14863;
  assign n14865 = po17  & ~n14864;
  assign n14866 = ~po17  & n14864;
  assign n14867 = ~n14339 & ~n14340;
  assign n14868 = po7  & n14867;
  assign n14869 = ~n14345 & ~n14868;
  assign n14870 = n14345 & n14868;
  assign n14871 = ~n14869 & ~n14870;
  assign n14872 = ~n14866 & ~n14871;
  assign n14873 = ~n14865 & ~n14872;
  assign n14874 = po18  & ~n14873;
  assign n14875 = ~po18  & n14873;
  assign n14876 = ~n14348 & ~n14349;
  assign n14877 = po7  & n14876;
  assign n14878 = ~n14354 & ~n14877;
  assign n14879 = n14354 & n14877;
  assign n14880 = ~n14878 & ~n14879;
  assign n14881 = ~n14875 & ~n14880;
  assign n14882 = ~n14874 & ~n14881;
  assign n14883 = po19  & ~n14882;
  assign n14884 = ~po19  & n14882;
  assign n14885 = ~n14357 & ~n14358;
  assign n14886 = po7  & n14885;
  assign n14887 = ~n14363 & ~n14886;
  assign n14888 = n14363 & n14886;
  assign n14889 = ~n14887 & ~n14888;
  assign n14890 = ~n14884 & ~n14889;
  assign n14891 = ~n14883 & ~n14890;
  assign n14892 = po20  & ~n14891;
  assign n14893 = ~po20  & n14891;
  assign n14894 = ~n14366 & ~n14367;
  assign n14895 = po7  & n14894;
  assign n14896 = ~n14372 & ~n14895;
  assign n14897 = n14372 & n14895;
  assign n14898 = ~n14896 & ~n14897;
  assign n14899 = ~n14893 & ~n14898;
  assign n14900 = ~n14892 & ~n14899;
  assign n14901 = po21  & ~n14900;
  assign n14902 = ~po21  & n14900;
  assign n14903 = ~n14375 & ~n14376;
  assign n14904 = po7  & n14903;
  assign n14905 = ~n14381 & ~n14904;
  assign n14906 = n14381 & n14904;
  assign n14907 = ~n14905 & ~n14906;
  assign n14908 = ~n14902 & ~n14907;
  assign n14909 = ~n14901 & ~n14908;
  assign n14910 = po22  & ~n14909;
  assign n14911 = ~po22  & n14909;
  assign n14912 = ~n14384 & ~n14385;
  assign n14913 = po7  & n14912;
  assign n14914 = ~n14390 & ~n14913;
  assign n14915 = n14390 & n14913;
  assign n14916 = ~n14914 & ~n14915;
  assign n14917 = ~n14911 & ~n14916;
  assign n14918 = ~n14910 & ~n14917;
  assign n14919 = po23  & ~n14918;
  assign n14920 = ~po23  & n14918;
  assign n14921 = ~n14393 & ~n14394;
  assign n14922 = po7  & n14921;
  assign n14923 = ~n14399 & ~n14922;
  assign n14924 = n14399 & n14922;
  assign n14925 = ~n14923 & ~n14924;
  assign n14926 = ~n14920 & ~n14925;
  assign n14927 = ~n14919 & ~n14926;
  assign n14928 = po24  & ~n14927;
  assign n14929 = ~po24  & n14927;
  assign n14930 = ~n14402 & ~n14403;
  assign n14931 = po7  & n14930;
  assign n14932 = ~n14408 & ~n14931;
  assign n14933 = n14408 & n14931;
  assign n14934 = ~n14932 & ~n14933;
  assign n14935 = ~n14929 & ~n14934;
  assign n14936 = ~n14928 & ~n14935;
  assign n14937 = po25  & ~n14936;
  assign n14938 = ~po25  & n14936;
  assign n14939 = ~n14411 & ~n14412;
  assign n14940 = po7  & n14939;
  assign n14941 = ~n14417 & ~n14940;
  assign n14942 = n14417 & n14940;
  assign n14943 = ~n14941 & ~n14942;
  assign n14944 = ~n14938 & ~n14943;
  assign n14945 = ~n14937 & ~n14944;
  assign n14946 = po26  & ~n14945;
  assign n14947 = ~po26  & n14945;
  assign n14948 = ~n14420 & ~n14421;
  assign n14949 = po7  & n14948;
  assign n14950 = ~n14426 & ~n14949;
  assign n14951 = n14426 & n14949;
  assign n14952 = ~n14950 & ~n14951;
  assign n14953 = ~n14947 & ~n14952;
  assign n14954 = ~n14946 & ~n14953;
  assign n14955 = po27  & ~n14954;
  assign n14956 = ~po27  & n14954;
  assign n14957 = ~n14429 & ~n14430;
  assign n14958 = po7  & n14957;
  assign n14959 = ~n14435 & ~n14958;
  assign n14960 = n14435 & n14958;
  assign n14961 = ~n14959 & ~n14960;
  assign n14962 = ~n14956 & ~n14961;
  assign n14963 = ~n14955 & ~n14962;
  assign n14964 = po28  & ~n14963;
  assign n14965 = ~po28  & n14963;
  assign n14966 = ~n14438 & ~n14439;
  assign n14967 = po7  & n14966;
  assign n14968 = ~n14444 & ~n14967;
  assign n14969 = n14444 & n14967;
  assign n14970 = ~n14968 & ~n14969;
  assign n14971 = ~n14965 & ~n14970;
  assign n14972 = ~n14964 & ~n14971;
  assign n14973 = po29  & ~n14972;
  assign n14974 = ~po29  & n14972;
  assign n14975 = ~n14447 & ~n14448;
  assign n14976 = po7  & n14975;
  assign n14977 = ~n14453 & ~n14976;
  assign n14978 = n14453 & n14976;
  assign n14979 = ~n14977 & ~n14978;
  assign n14980 = ~n14974 & ~n14979;
  assign n14981 = ~n14973 & ~n14980;
  assign n14982 = po30  & ~n14981;
  assign n14983 = ~po30  & n14981;
  assign n14984 = ~n14456 & ~n14457;
  assign n14985 = po7  & n14984;
  assign n14986 = ~n14462 & ~n14985;
  assign n14987 = n14462 & n14985;
  assign n14988 = ~n14986 & ~n14987;
  assign n14989 = ~n14983 & ~n14988;
  assign n14990 = ~n14982 & ~n14989;
  assign n14991 = po31  & ~n14990;
  assign n14992 = ~po31  & n14990;
  assign n14993 = ~n14465 & ~n14466;
  assign n14994 = po7  & n14993;
  assign n14995 = ~n14471 & ~n14994;
  assign n14996 = n14471 & n14994;
  assign n14997 = ~n14995 & ~n14996;
  assign n14998 = ~n14992 & ~n14997;
  assign n14999 = ~n14991 & ~n14998;
  assign n15000 = po32  & ~n14999;
  assign n15001 = ~po32  & n14999;
  assign n15002 = ~n14474 & ~n14475;
  assign n15003 = po7  & n15002;
  assign n15004 = ~n14480 & ~n15003;
  assign n15005 = n14480 & n15003;
  assign n15006 = ~n15004 & ~n15005;
  assign n15007 = ~n15001 & ~n15006;
  assign n15008 = ~n15000 & ~n15007;
  assign n15009 = po33  & ~n15008;
  assign n15010 = ~po33  & n15008;
  assign n15011 = ~n14483 & ~n14484;
  assign n15012 = po7  & n15011;
  assign n15013 = ~n14489 & ~n15012;
  assign n15014 = n14489 & n15012;
  assign n15015 = ~n15013 & ~n15014;
  assign n15016 = ~n15010 & ~n15015;
  assign n15017 = ~n15009 & ~n15016;
  assign n15018 = po34  & ~n15017;
  assign n15019 = ~po34  & n15017;
  assign n15020 = ~n14492 & ~n14493;
  assign n15021 = po7  & n15020;
  assign n15022 = ~n14498 & ~n15021;
  assign n15023 = n14498 & n15021;
  assign n15024 = ~n15022 & ~n15023;
  assign n15025 = ~n15019 & ~n15024;
  assign n15026 = ~n15018 & ~n15025;
  assign n15027 = po35  & ~n15026;
  assign n15028 = ~po35  & n15026;
  assign n15029 = ~n14501 & ~n14502;
  assign n15030 = po7  & n15029;
  assign n15031 = ~n14507 & ~n15030;
  assign n15032 = n14507 & n15030;
  assign n15033 = ~n15031 & ~n15032;
  assign n15034 = ~n15028 & ~n15033;
  assign n15035 = ~n15027 & ~n15034;
  assign n15036 = po36  & ~n15035;
  assign n15037 = ~po36  & n15035;
  assign n15038 = ~n14510 & ~n14511;
  assign n15039 = po7  & n15038;
  assign n15040 = ~n14516 & ~n15039;
  assign n15041 = n14516 & n15039;
  assign n15042 = ~n15040 & ~n15041;
  assign n15043 = ~n15037 & ~n15042;
  assign n15044 = ~n15036 & ~n15043;
  assign n15045 = po37  & ~n15044;
  assign n15046 = ~po37  & n15044;
  assign n15047 = ~n14519 & ~n14520;
  assign n15048 = po7  & n15047;
  assign n15049 = ~n14525 & ~n15048;
  assign n15050 = n14525 & n15048;
  assign n15051 = ~n15049 & ~n15050;
  assign n15052 = ~n15046 & ~n15051;
  assign n15053 = ~n15045 & ~n15052;
  assign n15054 = po38  & ~n15053;
  assign n15055 = ~po38  & n15053;
  assign n15056 = ~n14528 & ~n14529;
  assign n15057 = po7  & n15056;
  assign n15058 = ~n14534 & ~n15057;
  assign n15059 = n14534 & n15057;
  assign n15060 = ~n15058 & ~n15059;
  assign n15061 = ~n15055 & ~n15060;
  assign n15062 = ~n15054 & ~n15061;
  assign n15063 = po39  & ~n15062;
  assign n15064 = ~po39  & n15062;
  assign n15065 = ~n14537 & ~n14538;
  assign n15066 = po7  & n15065;
  assign n15067 = ~n14543 & ~n15066;
  assign n15068 = n14543 & n15066;
  assign n15069 = ~n15067 & ~n15068;
  assign n15070 = ~n15064 & ~n15069;
  assign n15071 = ~n15063 & ~n15070;
  assign n15072 = po40  & ~n15071;
  assign n15073 = ~po40  & n15071;
  assign n15074 = ~n14546 & ~n14547;
  assign n15075 = po7  & n15074;
  assign n15076 = ~n14552 & ~n15075;
  assign n15077 = n14552 & n15075;
  assign n15078 = ~n15076 & ~n15077;
  assign n15079 = ~n15073 & ~n15078;
  assign n15080 = ~n15072 & ~n15079;
  assign n15081 = po41  & ~n15080;
  assign n15082 = ~po41  & n15080;
  assign n15083 = ~n14555 & ~n14556;
  assign n15084 = po7  & n15083;
  assign n15085 = ~n14561 & ~n15084;
  assign n15086 = n14561 & n15084;
  assign n15087 = ~n15085 & ~n15086;
  assign n15088 = ~n15082 & ~n15087;
  assign n15089 = ~n15081 & ~n15088;
  assign n15090 = po42  & ~n15089;
  assign n15091 = ~po42  & n15089;
  assign n15092 = ~n14564 & ~n14565;
  assign n15093 = po7  & n15092;
  assign n15094 = ~n14570 & ~n15093;
  assign n15095 = n14570 & n15093;
  assign n15096 = ~n15094 & ~n15095;
  assign n15097 = ~n15091 & ~n15096;
  assign n15098 = ~n15090 & ~n15097;
  assign n15099 = po43  & ~n15098;
  assign n15100 = ~po43  & n15098;
  assign n15101 = ~n14573 & ~n14574;
  assign n15102 = po7  & n15101;
  assign n15103 = ~n14579 & ~n15102;
  assign n15104 = n14579 & n15102;
  assign n15105 = ~n15103 & ~n15104;
  assign n15106 = ~n15100 & ~n15105;
  assign n15107 = ~n15099 & ~n15106;
  assign n15108 = po44  & ~n15107;
  assign n15109 = ~po44  & n15107;
  assign n15110 = ~n14582 & ~n14583;
  assign n15111 = po7  & n15110;
  assign n15112 = ~n14588 & ~n15111;
  assign n15113 = n14588 & n15111;
  assign n15114 = ~n15112 & ~n15113;
  assign n15115 = ~n15109 & ~n15114;
  assign n15116 = ~n15108 & ~n15115;
  assign n15117 = po45  & ~n15116;
  assign n15118 = ~po45  & n15116;
  assign n15119 = ~n14591 & ~n14592;
  assign n15120 = po7  & n15119;
  assign n15121 = ~n14597 & ~n15120;
  assign n15122 = n14597 & n15120;
  assign n15123 = ~n15121 & ~n15122;
  assign n15124 = ~n15118 & ~n15123;
  assign n15125 = ~n15117 & ~n15124;
  assign n15126 = po46  & ~n15125;
  assign n15127 = ~po46  & n15125;
  assign n15128 = ~n14600 & ~n14601;
  assign n15129 = po7  & n15128;
  assign n15130 = ~n14606 & ~n15129;
  assign n15131 = n14606 & n15129;
  assign n15132 = ~n15130 & ~n15131;
  assign n15133 = ~n15127 & ~n15132;
  assign n15134 = ~n15126 & ~n15133;
  assign n15135 = po47  & ~n15134;
  assign n15136 = ~po47  & n15134;
  assign n15137 = ~n14609 & ~n14610;
  assign n15138 = po7  & n15137;
  assign n15139 = ~n14615 & ~n15138;
  assign n15140 = n14615 & n15138;
  assign n15141 = ~n15139 & ~n15140;
  assign n15142 = ~n15136 & ~n15141;
  assign n15143 = ~n15135 & ~n15142;
  assign n15144 = po48  & ~n15143;
  assign n15145 = ~po48  & n15143;
  assign n15146 = ~n14618 & ~n14619;
  assign n15147 = po7  & n15146;
  assign n15148 = ~n14624 & ~n15147;
  assign n15149 = n14624 & n15147;
  assign n15150 = ~n15148 & ~n15149;
  assign n15151 = ~n15145 & ~n15150;
  assign n15152 = ~n15144 & ~n15151;
  assign n15153 = po49  & ~n15152;
  assign n15154 = ~po49  & n15152;
  assign n15155 = ~n14627 & ~n14628;
  assign n15156 = po7  & n15155;
  assign n15157 = ~n14633 & ~n15156;
  assign n15158 = n14633 & n15156;
  assign n15159 = ~n15157 & ~n15158;
  assign n15160 = ~n15154 & ~n15159;
  assign n15161 = ~n15153 & ~n15160;
  assign n15162 = po50  & ~n15161;
  assign n15163 = ~po50  & n15161;
  assign n15164 = ~n14636 & ~n14637;
  assign n15165 = po7  & n15164;
  assign n15166 = ~n14642 & ~n15165;
  assign n15167 = n14642 & n15165;
  assign n15168 = ~n15166 & ~n15167;
  assign n15169 = ~n15163 & ~n15168;
  assign n15170 = ~n15162 & ~n15169;
  assign n15171 = po51  & ~n15170;
  assign n15172 = ~po51  & n15170;
  assign n15173 = ~n14645 & ~n14646;
  assign n15174 = po7  & n15173;
  assign n15175 = ~n14651 & ~n15174;
  assign n15176 = n14651 & n15174;
  assign n15177 = ~n15175 & ~n15176;
  assign n15178 = ~n15172 & ~n15177;
  assign n15179 = ~n15171 & ~n15178;
  assign n15180 = po52  & ~n15179;
  assign n15181 = ~po52  & n15179;
  assign n15182 = ~n14654 & ~n14655;
  assign n15183 = po7  & n15182;
  assign n15184 = ~n14660 & ~n15183;
  assign n15185 = n14660 & n15183;
  assign n15186 = ~n15184 & ~n15185;
  assign n15187 = ~n15181 & ~n15186;
  assign n15188 = ~n15180 & ~n15187;
  assign n15189 = po53  & ~n15188;
  assign n15190 = ~po53  & n15188;
  assign n15191 = ~n14663 & ~n14664;
  assign n15192 = po7  & n15191;
  assign n15193 = ~n14669 & ~n15192;
  assign n15194 = n14669 & n15192;
  assign n15195 = ~n15193 & ~n15194;
  assign n15196 = ~n15190 & ~n15195;
  assign n15197 = ~n15189 & ~n15196;
  assign n15198 = po54  & ~n15197;
  assign n15199 = ~po54  & n15197;
  assign n15200 = ~n14672 & ~n14673;
  assign n15201 = po7  & n15200;
  assign n15202 = ~n14678 & ~n15201;
  assign n15203 = n14678 & n15201;
  assign n15204 = ~n15202 & ~n15203;
  assign n15205 = ~n15199 & ~n15204;
  assign n15206 = ~n15198 & ~n15205;
  assign n15207 = po55  & ~n15206;
  assign n15208 = ~po55  & n15206;
  assign n15209 = ~n14681 & ~n14682;
  assign n15210 = po7  & n15209;
  assign n15211 = ~n14687 & ~n15210;
  assign n15212 = n14687 & n15210;
  assign n15213 = ~n15211 & ~n15212;
  assign n15214 = ~n15208 & ~n15213;
  assign n15215 = ~n15207 & ~n15214;
  assign n15216 = po56  & ~n15215;
  assign n15217 = ~po56  & n15215;
  assign n15218 = ~n14690 & ~n14691;
  assign n15219 = po7  & n15218;
  assign n15220 = ~n14696 & ~n15219;
  assign n15221 = n14696 & n15219;
  assign n15222 = ~n15220 & ~n15221;
  assign n15223 = ~n15217 & ~n15222;
  assign n15224 = ~n15216 & ~n15223;
  assign n15225 = po57  & ~n15224;
  assign n15226 = ~n14699 & ~n14705;
  assign n15227 = po7  & n15226;
  assign n15228 = ~n14704 & ~n15227;
  assign n15229 = n14704 & n15227;
  assign n15230 = ~n15228 & ~n15229;
  assign n15231 = ~po57  & n15224;
  assign n15232 = ~n15230 & ~n15231;
  assign n15233 = ~n15225 & ~n15232;
  assign n15234 = po58  & ~n15233;
  assign n15235 = ~po58  & n15233;
  assign n15236 = ~n14770 & ~n15235;
  assign n15237 = ~n15234 & ~n15236;
  assign n15238 = po59  & ~n15237;
  assign n15239 = ~po59  & n15237;
  assign n15240 = ~n14712 & ~n14713;
  assign n15241 = po7  & n15240;
  assign n15242 = ~n14718 & ~n15241;
  assign n15243 = n14718 & n15241;
  assign n15244 = ~n15242 & ~n15243;
  assign n15245 = ~n15239 & ~n15244;
  assign n15246 = ~n15238 & ~n15245;
  assign n15247 = po60  & ~n15246;
  assign n15248 = ~po60  & n15246;
  assign n15249 = ~n14721 & ~n14722;
  assign n15250 = po7  & n15249;
  assign n15251 = ~n14727 & ~n15250;
  assign n15252 = n14727 & n15250;
  assign n15253 = ~n15251 & ~n15252;
  assign n15254 = ~n15248 & ~n15253;
  assign n15255 = ~n15247 & ~n15254;
  assign n15256 = po61  & ~n15255;
  assign n15257 = ~po61  & n15255;
  assign n15258 = ~n14730 & ~n14731;
  assign n15259 = po7  & n15258;
  assign n15260 = ~n14736 & ~n15259;
  assign n15261 = n14736 & n15259;
  assign n15262 = ~n15260 & ~n15261;
  assign n15263 = ~n15257 & ~n15262;
  assign n15264 = ~n15256 & ~n15263;
  assign n15265 = po62  & ~n15264;
  assign n15266 = ~po62  & n15264;
  assign n15267 = ~n14739 & ~n14740;
  assign n15268 = po7  & n15267;
  assign n15269 = ~n14745 & ~n15268;
  assign n15270 = n14745 & n15268;
  assign n15271 = ~n15269 & ~n15270;
  assign n15272 = ~n15266 & ~n15271;
  assign n15273 = ~n15265 & ~n15272;
  assign n15274 = n14780 & n15273;
  assign n15275 = ~n14780 & ~n15273;
  assign n15276 = n14758 & po7 ;
  assign n15277 = ~n14757 & ~n15276;
  assign n15278 = n15275 & n15277;
  assign n15279 = ~po63  & ~n15278;
  assign n15280 = ~n15274 & ~n15279;
  assign n15281 = ~n14775 & n15280;
  assign po6  = n14771 | ~n15281;
  assign n15283 = ~n15234 & ~n15235;
  assign n15284 = po6  & n15283;
  assign n15285 = ~n14770 & ~n15284;
  assign n15286 = n14770 & n15284;
  assign n15287 = ~n15285 & ~n15286;
  assign n15288 = ~n15265 & ~n15266;
  assign n15289 = po6  & n15288;
  assign n15290 = ~n15271 & ~n15289;
  assign n15291 = n15271 & n15289;
  assign n15292 = ~n15290 & ~n15291;
  assign n15293 = pi12  & po6 ;
  assign n15294 = ~pi10  & ~pi11 ;
  assign n15295 = ~pi12  & n15294;
  assign n15296 = ~n15293 & ~n15295;
  assign n15297 = po7  & ~n15296;
  assign n15298 = ~po7  & n15296;
  assign n15299 = ~pi12  & po6 ;
  assign n15300 = pi13  & ~n15299;
  assign n15301 = n14782 & po6 ;
  assign n15302 = ~n15300 & ~n15301;
  assign n15303 = ~n15298 & n15302;
  assign n15304 = ~n15297 & ~n15303;
  assign n15305 = po8  & ~n15304;
  assign n15306 = ~po8  & n15304;
  assign n15307 = po7  & n15281;
  assign n15308 = ~n15301 & ~n15307;
  assign n15309 = pi14  & ~n15308;
  assign n15310 = ~pi14  & n15308;
  assign n15311 = ~n15309 & ~n15310;
  assign n15312 = ~n15306 & ~n15311;
  assign n15313 = ~n15305 & ~n15312;
  assign n15314 = po9  & ~n15313;
  assign n15315 = ~po9  & n15313;
  assign n15316 = ~n14785 & ~n14786;
  assign n15317 = po6  & n15316;
  assign n15318 = n14790 & ~n15317;
  assign n15319 = ~n14790 & n15317;
  assign n15320 = ~n15318 & ~n15319;
  assign n15321 = ~n15315 & ~n15320;
  assign n15322 = ~n15314 & ~n15321;
  assign n15323 = po10  & ~n15322;
  assign n15324 = ~po10  & n15322;
  assign n15325 = ~n14793 & ~n14794;
  assign n15326 = po6  & n15325;
  assign n15327 = ~n14799 & ~n15326;
  assign n15328 = n14799 & n15326;
  assign n15329 = ~n15327 & ~n15328;
  assign n15330 = ~n15324 & ~n15329;
  assign n15331 = ~n15323 & ~n15330;
  assign n15332 = po11  & ~n15331;
  assign n15333 = ~po11  & n15331;
  assign n15334 = ~n14802 & ~n14803;
  assign n15335 = po6  & n15334;
  assign n15336 = n14808 & n15335;
  assign n15337 = ~n14808 & ~n15335;
  assign n15338 = ~n15336 & ~n15337;
  assign n15339 = ~n15333 & ~n15338;
  assign n15340 = ~n15332 & ~n15339;
  assign n15341 = po12  & ~n15340;
  assign n15342 = ~po12  & n15340;
  assign n15343 = ~n14811 & ~n14812;
  assign n15344 = po6  & n15343;
  assign n15345 = ~n14817 & ~n15344;
  assign n15346 = n14817 & n15344;
  assign n15347 = ~n15345 & ~n15346;
  assign n15348 = ~n15342 & ~n15347;
  assign n15349 = ~n15341 & ~n15348;
  assign n15350 = po13  & ~n15349;
  assign n15351 = ~po13  & n15349;
  assign n15352 = ~n14820 & ~n14821;
  assign n15353 = po6  & n15352;
  assign n15354 = ~n14826 & ~n15353;
  assign n15355 = n14826 & n15353;
  assign n15356 = ~n15354 & ~n15355;
  assign n15357 = ~n15351 & ~n15356;
  assign n15358 = ~n15350 & ~n15357;
  assign n15359 = po14  & ~n15358;
  assign n15360 = ~po14  & n15358;
  assign n15361 = ~n14829 & ~n14830;
  assign n15362 = po6  & n15361;
  assign n15363 = ~n14835 & ~n15362;
  assign n15364 = n14835 & n15362;
  assign n15365 = ~n15363 & ~n15364;
  assign n15366 = ~n15360 & ~n15365;
  assign n15367 = ~n15359 & ~n15366;
  assign n15368 = po15  & ~n15367;
  assign n15369 = ~po15  & n15367;
  assign n15370 = ~n14838 & ~n14839;
  assign n15371 = po6  & n15370;
  assign n15372 = ~n14844 & ~n15371;
  assign n15373 = n14844 & n15371;
  assign n15374 = ~n15372 & ~n15373;
  assign n15375 = ~n15369 & ~n15374;
  assign n15376 = ~n15368 & ~n15375;
  assign n15377 = po16  & ~n15376;
  assign n15378 = ~po16  & n15376;
  assign n15379 = ~n14847 & ~n14848;
  assign n15380 = po6  & n15379;
  assign n15381 = ~n14853 & ~n15380;
  assign n15382 = n14853 & n15380;
  assign n15383 = ~n15381 & ~n15382;
  assign n15384 = ~n15378 & ~n15383;
  assign n15385 = ~n15377 & ~n15384;
  assign n15386 = po17  & ~n15385;
  assign n15387 = ~po17  & n15385;
  assign n15388 = ~n14856 & ~n14857;
  assign n15389 = po6  & n15388;
  assign n15390 = ~n14862 & ~n15389;
  assign n15391 = n14862 & n15389;
  assign n15392 = ~n15390 & ~n15391;
  assign n15393 = ~n15387 & ~n15392;
  assign n15394 = ~n15386 & ~n15393;
  assign n15395 = po18  & ~n15394;
  assign n15396 = ~po18  & n15394;
  assign n15397 = ~n14865 & ~n14866;
  assign n15398 = po6  & n15397;
  assign n15399 = ~n14871 & ~n15398;
  assign n15400 = n14871 & n15398;
  assign n15401 = ~n15399 & ~n15400;
  assign n15402 = ~n15396 & ~n15401;
  assign n15403 = ~n15395 & ~n15402;
  assign n15404 = po19  & ~n15403;
  assign n15405 = ~po19  & n15403;
  assign n15406 = ~n14874 & ~n14875;
  assign n15407 = po6  & n15406;
  assign n15408 = ~n14880 & ~n15407;
  assign n15409 = n14880 & n15407;
  assign n15410 = ~n15408 & ~n15409;
  assign n15411 = ~n15405 & ~n15410;
  assign n15412 = ~n15404 & ~n15411;
  assign n15413 = po20  & ~n15412;
  assign n15414 = ~po20  & n15412;
  assign n15415 = ~n14883 & ~n14884;
  assign n15416 = po6  & n15415;
  assign n15417 = ~n14889 & ~n15416;
  assign n15418 = n14889 & n15416;
  assign n15419 = ~n15417 & ~n15418;
  assign n15420 = ~n15414 & ~n15419;
  assign n15421 = ~n15413 & ~n15420;
  assign n15422 = po21  & ~n15421;
  assign n15423 = ~po21  & n15421;
  assign n15424 = ~n14892 & ~n14893;
  assign n15425 = po6  & n15424;
  assign n15426 = ~n14898 & ~n15425;
  assign n15427 = n14898 & n15425;
  assign n15428 = ~n15426 & ~n15427;
  assign n15429 = ~n15423 & ~n15428;
  assign n15430 = ~n15422 & ~n15429;
  assign n15431 = po22  & ~n15430;
  assign n15432 = ~po22  & n15430;
  assign n15433 = ~n14901 & ~n14902;
  assign n15434 = po6  & n15433;
  assign n15435 = ~n14907 & ~n15434;
  assign n15436 = n14907 & n15434;
  assign n15437 = ~n15435 & ~n15436;
  assign n15438 = ~n15432 & ~n15437;
  assign n15439 = ~n15431 & ~n15438;
  assign n15440 = po23  & ~n15439;
  assign n15441 = ~po23  & n15439;
  assign n15442 = ~n14910 & ~n14911;
  assign n15443 = po6  & n15442;
  assign n15444 = ~n14916 & ~n15443;
  assign n15445 = n14916 & n15443;
  assign n15446 = ~n15444 & ~n15445;
  assign n15447 = ~n15441 & ~n15446;
  assign n15448 = ~n15440 & ~n15447;
  assign n15449 = po24  & ~n15448;
  assign n15450 = ~po24  & n15448;
  assign n15451 = ~n14919 & ~n14920;
  assign n15452 = po6  & n15451;
  assign n15453 = ~n14925 & ~n15452;
  assign n15454 = n14925 & n15452;
  assign n15455 = ~n15453 & ~n15454;
  assign n15456 = ~n15450 & ~n15455;
  assign n15457 = ~n15449 & ~n15456;
  assign n15458 = po25  & ~n15457;
  assign n15459 = ~po25  & n15457;
  assign n15460 = ~n14928 & ~n14929;
  assign n15461 = po6  & n15460;
  assign n15462 = ~n14934 & ~n15461;
  assign n15463 = n14934 & n15461;
  assign n15464 = ~n15462 & ~n15463;
  assign n15465 = ~n15459 & ~n15464;
  assign n15466 = ~n15458 & ~n15465;
  assign n15467 = po26  & ~n15466;
  assign n15468 = ~po26  & n15466;
  assign n15469 = ~n14937 & ~n14938;
  assign n15470 = po6  & n15469;
  assign n15471 = ~n14943 & ~n15470;
  assign n15472 = n14943 & n15470;
  assign n15473 = ~n15471 & ~n15472;
  assign n15474 = ~n15468 & ~n15473;
  assign n15475 = ~n15467 & ~n15474;
  assign n15476 = po27  & ~n15475;
  assign n15477 = ~po27  & n15475;
  assign n15478 = ~n14946 & ~n14947;
  assign n15479 = po6  & n15478;
  assign n15480 = ~n14952 & ~n15479;
  assign n15481 = n14952 & n15479;
  assign n15482 = ~n15480 & ~n15481;
  assign n15483 = ~n15477 & ~n15482;
  assign n15484 = ~n15476 & ~n15483;
  assign n15485 = po28  & ~n15484;
  assign n15486 = ~po28  & n15484;
  assign n15487 = ~n14955 & ~n14956;
  assign n15488 = po6  & n15487;
  assign n15489 = ~n14961 & ~n15488;
  assign n15490 = n14961 & n15488;
  assign n15491 = ~n15489 & ~n15490;
  assign n15492 = ~n15486 & ~n15491;
  assign n15493 = ~n15485 & ~n15492;
  assign n15494 = po29  & ~n15493;
  assign n15495 = ~po29  & n15493;
  assign n15496 = ~n14964 & ~n14965;
  assign n15497 = po6  & n15496;
  assign n15498 = ~n14970 & ~n15497;
  assign n15499 = n14970 & n15497;
  assign n15500 = ~n15498 & ~n15499;
  assign n15501 = ~n15495 & ~n15500;
  assign n15502 = ~n15494 & ~n15501;
  assign n15503 = po30  & ~n15502;
  assign n15504 = ~po30  & n15502;
  assign n15505 = ~n14973 & ~n14974;
  assign n15506 = po6  & n15505;
  assign n15507 = ~n14979 & ~n15506;
  assign n15508 = n14979 & n15506;
  assign n15509 = ~n15507 & ~n15508;
  assign n15510 = ~n15504 & ~n15509;
  assign n15511 = ~n15503 & ~n15510;
  assign n15512 = po31  & ~n15511;
  assign n15513 = ~po31  & n15511;
  assign n15514 = ~n14982 & ~n14983;
  assign n15515 = po6  & n15514;
  assign n15516 = ~n14988 & ~n15515;
  assign n15517 = n14988 & n15515;
  assign n15518 = ~n15516 & ~n15517;
  assign n15519 = ~n15513 & ~n15518;
  assign n15520 = ~n15512 & ~n15519;
  assign n15521 = po32  & ~n15520;
  assign n15522 = ~po32  & n15520;
  assign n15523 = ~n14991 & ~n14992;
  assign n15524 = po6  & n15523;
  assign n15525 = ~n14997 & ~n15524;
  assign n15526 = n14997 & n15524;
  assign n15527 = ~n15525 & ~n15526;
  assign n15528 = ~n15522 & ~n15527;
  assign n15529 = ~n15521 & ~n15528;
  assign n15530 = po33  & ~n15529;
  assign n15531 = ~po33  & n15529;
  assign n15532 = ~n15000 & ~n15001;
  assign n15533 = po6  & n15532;
  assign n15534 = ~n15006 & ~n15533;
  assign n15535 = n15006 & n15533;
  assign n15536 = ~n15534 & ~n15535;
  assign n15537 = ~n15531 & ~n15536;
  assign n15538 = ~n15530 & ~n15537;
  assign n15539 = po34  & ~n15538;
  assign n15540 = ~po34  & n15538;
  assign n15541 = ~n15009 & ~n15010;
  assign n15542 = po6  & n15541;
  assign n15543 = ~n15015 & ~n15542;
  assign n15544 = n15015 & n15542;
  assign n15545 = ~n15543 & ~n15544;
  assign n15546 = ~n15540 & ~n15545;
  assign n15547 = ~n15539 & ~n15546;
  assign n15548 = po35  & ~n15547;
  assign n15549 = ~po35  & n15547;
  assign n15550 = ~n15018 & ~n15019;
  assign n15551 = po6  & n15550;
  assign n15552 = ~n15024 & ~n15551;
  assign n15553 = n15024 & n15551;
  assign n15554 = ~n15552 & ~n15553;
  assign n15555 = ~n15549 & ~n15554;
  assign n15556 = ~n15548 & ~n15555;
  assign n15557 = po36  & ~n15556;
  assign n15558 = ~po36  & n15556;
  assign n15559 = ~n15027 & ~n15028;
  assign n15560 = po6  & n15559;
  assign n15561 = ~n15033 & ~n15560;
  assign n15562 = n15033 & n15560;
  assign n15563 = ~n15561 & ~n15562;
  assign n15564 = ~n15558 & ~n15563;
  assign n15565 = ~n15557 & ~n15564;
  assign n15566 = po37  & ~n15565;
  assign n15567 = ~po37  & n15565;
  assign n15568 = ~n15036 & ~n15037;
  assign n15569 = po6  & n15568;
  assign n15570 = ~n15042 & ~n15569;
  assign n15571 = n15042 & n15569;
  assign n15572 = ~n15570 & ~n15571;
  assign n15573 = ~n15567 & ~n15572;
  assign n15574 = ~n15566 & ~n15573;
  assign n15575 = po38  & ~n15574;
  assign n15576 = ~po38  & n15574;
  assign n15577 = ~n15045 & ~n15046;
  assign n15578 = po6  & n15577;
  assign n15579 = ~n15051 & ~n15578;
  assign n15580 = n15051 & n15578;
  assign n15581 = ~n15579 & ~n15580;
  assign n15582 = ~n15576 & ~n15581;
  assign n15583 = ~n15575 & ~n15582;
  assign n15584 = po39  & ~n15583;
  assign n15585 = ~po39  & n15583;
  assign n15586 = ~n15054 & ~n15055;
  assign n15587 = po6  & n15586;
  assign n15588 = ~n15060 & ~n15587;
  assign n15589 = n15060 & n15587;
  assign n15590 = ~n15588 & ~n15589;
  assign n15591 = ~n15585 & ~n15590;
  assign n15592 = ~n15584 & ~n15591;
  assign n15593 = po40  & ~n15592;
  assign n15594 = ~po40  & n15592;
  assign n15595 = ~n15063 & ~n15064;
  assign n15596 = po6  & n15595;
  assign n15597 = ~n15069 & ~n15596;
  assign n15598 = n15069 & n15596;
  assign n15599 = ~n15597 & ~n15598;
  assign n15600 = ~n15594 & ~n15599;
  assign n15601 = ~n15593 & ~n15600;
  assign n15602 = po41  & ~n15601;
  assign n15603 = ~po41  & n15601;
  assign n15604 = ~n15072 & ~n15073;
  assign n15605 = po6  & n15604;
  assign n15606 = ~n15078 & ~n15605;
  assign n15607 = n15078 & n15605;
  assign n15608 = ~n15606 & ~n15607;
  assign n15609 = ~n15603 & ~n15608;
  assign n15610 = ~n15602 & ~n15609;
  assign n15611 = po42  & ~n15610;
  assign n15612 = ~po42  & n15610;
  assign n15613 = ~n15081 & ~n15082;
  assign n15614 = po6  & n15613;
  assign n15615 = ~n15087 & ~n15614;
  assign n15616 = n15087 & n15614;
  assign n15617 = ~n15615 & ~n15616;
  assign n15618 = ~n15612 & ~n15617;
  assign n15619 = ~n15611 & ~n15618;
  assign n15620 = po43  & ~n15619;
  assign n15621 = ~po43  & n15619;
  assign n15622 = ~n15090 & ~n15091;
  assign n15623 = po6  & n15622;
  assign n15624 = ~n15096 & ~n15623;
  assign n15625 = n15096 & n15623;
  assign n15626 = ~n15624 & ~n15625;
  assign n15627 = ~n15621 & ~n15626;
  assign n15628 = ~n15620 & ~n15627;
  assign n15629 = po44  & ~n15628;
  assign n15630 = ~po44  & n15628;
  assign n15631 = ~n15099 & ~n15100;
  assign n15632 = po6  & n15631;
  assign n15633 = ~n15105 & ~n15632;
  assign n15634 = n15105 & n15632;
  assign n15635 = ~n15633 & ~n15634;
  assign n15636 = ~n15630 & ~n15635;
  assign n15637 = ~n15629 & ~n15636;
  assign n15638 = po45  & ~n15637;
  assign n15639 = ~po45  & n15637;
  assign n15640 = ~n15108 & ~n15109;
  assign n15641 = po6  & n15640;
  assign n15642 = ~n15114 & ~n15641;
  assign n15643 = n15114 & n15641;
  assign n15644 = ~n15642 & ~n15643;
  assign n15645 = ~n15639 & ~n15644;
  assign n15646 = ~n15638 & ~n15645;
  assign n15647 = po46  & ~n15646;
  assign n15648 = ~po46  & n15646;
  assign n15649 = ~n15117 & ~n15118;
  assign n15650 = po6  & n15649;
  assign n15651 = ~n15123 & ~n15650;
  assign n15652 = n15123 & n15650;
  assign n15653 = ~n15651 & ~n15652;
  assign n15654 = ~n15648 & ~n15653;
  assign n15655 = ~n15647 & ~n15654;
  assign n15656 = po47  & ~n15655;
  assign n15657 = ~po47  & n15655;
  assign n15658 = ~n15126 & ~n15127;
  assign n15659 = po6  & n15658;
  assign n15660 = ~n15132 & ~n15659;
  assign n15661 = n15132 & n15659;
  assign n15662 = ~n15660 & ~n15661;
  assign n15663 = ~n15657 & ~n15662;
  assign n15664 = ~n15656 & ~n15663;
  assign n15665 = po48  & ~n15664;
  assign n15666 = ~po48  & n15664;
  assign n15667 = ~n15135 & ~n15136;
  assign n15668 = po6  & n15667;
  assign n15669 = ~n15141 & ~n15668;
  assign n15670 = n15141 & n15668;
  assign n15671 = ~n15669 & ~n15670;
  assign n15672 = ~n15666 & ~n15671;
  assign n15673 = ~n15665 & ~n15672;
  assign n15674 = po49  & ~n15673;
  assign n15675 = ~po49  & n15673;
  assign n15676 = ~n15144 & ~n15145;
  assign n15677 = po6  & n15676;
  assign n15678 = ~n15150 & ~n15677;
  assign n15679 = n15150 & n15677;
  assign n15680 = ~n15678 & ~n15679;
  assign n15681 = ~n15675 & ~n15680;
  assign n15682 = ~n15674 & ~n15681;
  assign n15683 = po50  & ~n15682;
  assign n15684 = ~po50  & n15682;
  assign n15685 = ~n15153 & ~n15154;
  assign n15686 = po6  & n15685;
  assign n15687 = ~n15159 & ~n15686;
  assign n15688 = n15159 & n15686;
  assign n15689 = ~n15687 & ~n15688;
  assign n15690 = ~n15684 & ~n15689;
  assign n15691 = ~n15683 & ~n15690;
  assign n15692 = po51  & ~n15691;
  assign n15693 = ~po51  & n15691;
  assign n15694 = ~n15162 & ~n15163;
  assign n15695 = po6  & n15694;
  assign n15696 = ~n15168 & ~n15695;
  assign n15697 = n15168 & n15695;
  assign n15698 = ~n15696 & ~n15697;
  assign n15699 = ~n15693 & ~n15698;
  assign n15700 = ~n15692 & ~n15699;
  assign n15701 = po52  & ~n15700;
  assign n15702 = ~po52  & n15700;
  assign n15703 = ~n15171 & ~n15172;
  assign n15704 = po6  & n15703;
  assign n15705 = ~n15177 & ~n15704;
  assign n15706 = n15177 & n15704;
  assign n15707 = ~n15705 & ~n15706;
  assign n15708 = ~n15702 & ~n15707;
  assign n15709 = ~n15701 & ~n15708;
  assign n15710 = po53  & ~n15709;
  assign n15711 = ~po53  & n15709;
  assign n15712 = ~n15180 & ~n15181;
  assign n15713 = po6  & n15712;
  assign n15714 = ~n15186 & ~n15713;
  assign n15715 = n15186 & n15713;
  assign n15716 = ~n15714 & ~n15715;
  assign n15717 = ~n15711 & ~n15716;
  assign n15718 = ~n15710 & ~n15717;
  assign n15719 = po54  & ~n15718;
  assign n15720 = ~po54  & n15718;
  assign n15721 = ~n15189 & ~n15190;
  assign n15722 = po6  & n15721;
  assign n15723 = ~n15195 & ~n15722;
  assign n15724 = n15195 & n15722;
  assign n15725 = ~n15723 & ~n15724;
  assign n15726 = ~n15720 & ~n15725;
  assign n15727 = ~n15719 & ~n15726;
  assign n15728 = po55  & ~n15727;
  assign n15729 = ~po55  & n15727;
  assign n15730 = ~n15198 & ~n15199;
  assign n15731 = po6  & n15730;
  assign n15732 = ~n15204 & ~n15731;
  assign n15733 = n15204 & n15731;
  assign n15734 = ~n15732 & ~n15733;
  assign n15735 = ~n15729 & ~n15734;
  assign n15736 = ~n15728 & ~n15735;
  assign n15737 = po56  & ~n15736;
  assign n15738 = ~po56  & n15736;
  assign n15739 = ~n15207 & ~n15208;
  assign n15740 = po6  & n15739;
  assign n15741 = ~n15213 & ~n15740;
  assign n15742 = n15213 & n15740;
  assign n15743 = ~n15741 & ~n15742;
  assign n15744 = ~n15738 & ~n15743;
  assign n15745 = ~n15737 & ~n15744;
  assign n15746 = po57  & ~n15745;
  assign n15747 = ~po57  & n15745;
  assign n15748 = ~n15216 & ~n15217;
  assign n15749 = po6  & n15748;
  assign n15750 = ~n15222 & ~n15749;
  assign n15751 = n15222 & n15749;
  assign n15752 = ~n15750 & ~n15751;
  assign n15753 = ~n15747 & ~n15752;
  assign n15754 = ~n15746 & ~n15753;
  assign n15755 = po58  & ~n15754;
  assign n15756 = ~n15225 & ~n15231;
  assign n15757 = po6  & n15756;
  assign n15758 = ~n15230 & ~n15757;
  assign n15759 = n15230 & n15757;
  assign n15760 = ~n15758 & ~n15759;
  assign n15761 = ~po58  & n15754;
  assign n15762 = ~n15760 & ~n15761;
  assign n15763 = ~n15755 & ~n15762;
  assign n15764 = po59  & ~n15763;
  assign n15765 = ~po59  & n15763;
  assign n15766 = ~n15287 & ~n15765;
  assign n15767 = ~n15764 & ~n15766;
  assign n15768 = po60  & ~n15767;
  assign n15769 = ~po60  & n15767;
  assign n15770 = ~n15238 & ~n15239;
  assign n15771 = po6  & n15770;
  assign n15772 = ~n15244 & ~n15771;
  assign n15773 = n15244 & n15771;
  assign n15774 = ~n15772 & ~n15773;
  assign n15775 = ~n15769 & ~n15774;
  assign n15776 = ~n15768 & ~n15775;
  assign n15777 = po61  & ~n15776;
  assign n15778 = ~po61  & n15776;
  assign n15779 = ~n15247 & ~n15248;
  assign n15780 = po6  & n15779;
  assign n15781 = ~n15253 & ~n15780;
  assign n15782 = n15253 & n15780;
  assign n15783 = ~n15781 & ~n15782;
  assign n15784 = ~n15778 & ~n15783;
  assign n15785 = ~n15777 & ~n15784;
  assign n15786 = po62  & ~n15785;
  assign n15787 = ~po62  & n15785;
  assign n15788 = ~n15256 & ~n15257;
  assign n15789 = po6  & n15788;
  assign n15790 = ~n15262 & ~n15789;
  assign n15791 = n15262 & n15789;
  assign n15792 = ~n15790 & ~n15791;
  assign n15793 = ~n15787 & ~n15792;
  assign n15794 = ~n15786 & ~n15793;
  assign n15795 = n15292 & n15794;
  assign n15796 = ~n15292 & ~n15794;
  assign n15797 = n15275 & po6 ;
  assign n15798 = ~n15274 & ~n15797;
  assign n15799 = n15796 & n15798;
  assign n15800 = ~po63  & ~n15799;
  assign n15801 = ~n14780 & po6 ;
  assign n15802 = n15273 & ~n15801;
  assign n15803 = po63  & ~n15275;
  assign n15804 = ~n15802 & n15803;
  assign n15805 = ~n15800 & ~n15804;
  assign po5  = n15795 | ~n15805;
  assign n15807 = ~n15764 & ~n15765;
  assign n15808 = po5  & n15807;
  assign n15809 = ~n15287 & ~n15808;
  assign n15810 = n15287 & n15808;
  assign n15811 = ~n15809 & ~n15810;
  assign n15812 = ~n15786 & ~n15787;
  assign n15813 = po5  & n15812;
  assign n15814 = ~n15792 & ~n15813;
  assign n15815 = n15792 & n15813;
  assign n15816 = ~n15814 & ~n15815;
  assign n15817 = pi10  & po5 ;
  assign n15818 = ~pi8  & ~pi9 ;
  assign n15819 = ~pi10  & n15818;
  assign n15820 = ~n15817 & ~n15819;
  assign n15821 = po6  & ~n15820;
  assign n15822 = ~po6  & n15820;
  assign n15823 = ~pi10  & po5 ;
  assign n15824 = pi11  & ~n15823;
  assign n15825 = n15294 & po5 ;
  assign n15826 = ~n15824 & ~n15825;
  assign n15827 = ~n15822 & n15826;
  assign n15828 = ~n15821 & ~n15827;
  assign n15829 = po7  & ~n15828;
  assign n15830 = ~po7  & n15828;
  assign n15831 = po6  & ~po5 ;
  assign n15832 = ~n15825 & ~n15831;
  assign n15833 = pi12  & ~n15832;
  assign n15834 = ~pi12  & n15832;
  assign n15835 = ~n15833 & ~n15834;
  assign n15836 = ~n15830 & ~n15835;
  assign n15837 = ~n15829 & ~n15836;
  assign n15838 = po8  & ~n15837;
  assign n15839 = ~po8  & n15837;
  assign n15840 = ~n15297 & ~n15298;
  assign n15841 = po5  & n15840;
  assign n15842 = n15302 & ~n15841;
  assign n15843 = ~n15302 & n15841;
  assign n15844 = ~n15842 & ~n15843;
  assign n15845 = ~n15839 & ~n15844;
  assign n15846 = ~n15838 & ~n15845;
  assign n15847 = po9  & ~n15846;
  assign n15848 = ~po9  & n15846;
  assign n15849 = ~n15305 & ~n15306;
  assign n15850 = po5  & n15849;
  assign n15851 = ~n15311 & ~n15850;
  assign n15852 = n15311 & n15850;
  assign n15853 = ~n15851 & ~n15852;
  assign n15854 = ~n15848 & ~n15853;
  assign n15855 = ~n15847 & ~n15854;
  assign n15856 = po10  & ~n15855;
  assign n15857 = ~po10  & n15855;
  assign n15858 = ~n15314 & ~n15315;
  assign n15859 = po5  & n15858;
  assign n15860 = n15320 & n15859;
  assign n15861 = ~n15320 & ~n15859;
  assign n15862 = ~n15860 & ~n15861;
  assign n15863 = ~n15857 & ~n15862;
  assign n15864 = ~n15856 & ~n15863;
  assign n15865 = po11  & ~n15864;
  assign n15866 = ~po11  & n15864;
  assign n15867 = ~n15323 & ~n15324;
  assign n15868 = po5  & n15867;
  assign n15869 = ~n15329 & ~n15868;
  assign n15870 = n15329 & n15868;
  assign n15871 = ~n15869 & ~n15870;
  assign n15872 = ~n15866 & ~n15871;
  assign n15873 = ~n15865 & ~n15872;
  assign n15874 = po12  & ~n15873;
  assign n15875 = ~po12  & n15873;
  assign n15876 = ~n15332 & ~n15333;
  assign n15877 = po5  & n15876;
  assign n15878 = ~n15338 & ~n15877;
  assign n15879 = n15338 & n15877;
  assign n15880 = ~n15878 & ~n15879;
  assign n15881 = ~n15875 & ~n15880;
  assign n15882 = ~n15874 & ~n15881;
  assign n15883 = po13  & ~n15882;
  assign n15884 = ~po13  & n15882;
  assign n15885 = ~n15341 & ~n15342;
  assign n15886 = po5  & n15885;
  assign n15887 = ~n15347 & ~n15886;
  assign n15888 = n15347 & n15886;
  assign n15889 = ~n15887 & ~n15888;
  assign n15890 = ~n15884 & ~n15889;
  assign n15891 = ~n15883 & ~n15890;
  assign n15892 = po14  & ~n15891;
  assign n15893 = ~po14  & n15891;
  assign n15894 = ~n15350 & ~n15351;
  assign n15895 = po5  & n15894;
  assign n15896 = ~n15356 & ~n15895;
  assign n15897 = n15356 & n15895;
  assign n15898 = ~n15896 & ~n15897;
  assign n15899 = ~n15893 & ~n15898;
  assign n15900 = ~n15892 & ~n15899;
  assign n15901 = po15  & ~n15900;
  assign n15902 = ~po15  & n15900;
  assign n15903 = ~n15359 & ~n15360;
  assign n15904 = po5  & n15903;
  assign n15905 = ~n15365 & ~n15904;
  assign n15906 = n15365 & n15904;
  assign n15907 = ~n15905 & ~n15906;
  assign n15908 = ~n15902 & ~n15907;
  assign n15909 = ~n15901 & ~n15908;
  assign n15910 = po16  & ~n15909;
  assign n15911 = ~po16  & n15909;
  assign n15912 = ~n15368 & ~n15369;
  assign n15913 = po5  & n15912;
  assign n15914 = ~n15374 & ~n15913;
  assign n15915 = n15374 & n15913;
  assign n15916 = ~n15914 & ~n15915;
  assign n15917 = ~n15911 & ~n15916;
  assign n15918 = ~n15910 & ~n15917;
  assign n15919 = po17  & ~n15918;
  assign n15920 = ~po17  & n15918;
  assign n15921 = ~n15377 & ~n15378;
  assign n15922 = po5  & n15921;
  assign n15923 = ~n15383 & ~n15922;
  assign n15924 = n15383 & n15922;
  assign n15925 = ~n15923 & ~n15924;
  assign n15926 = ~n15920 & ~n15925;
  assign n15927 = ~n15919 & ~n15926;
  assign n15928 = po18  & ~n15927;
  assign n15929 = ~po18  & n15927;
  assign n15930 = ~n15386 & ~n15387;
  assign n15931 = po5  & n15930;
  assign n15932 = ~n15392 & ~n15931;
  assign n15933 = n15392 & n15931;
  assign n15934 = ~n15932 & ~n15933;
  assign n15935 = ~n15929 & ~n15934;
  assign n15936 = ~n15928 & ~n15935;
  assign n15937 = po19  & ~n15936;
  assign n15938 = ~po19  & n15936;
  assign n15939 = ~n15395 & ~n15396;
  assign n15940 = po5  & n15939;
  assign n15941 = ~n15401 & ~n15940;
  assign n15942 = n15401 & n15940;
  assign n15943 = ~n15941 & ~n15942;
  assign n15944 = ~n15938 & ~n15943;
  assign n15945 = ~n15937 & ~n15944;
  assign n15946 = po20  & ~n15945;
  assign n15947 = ~po20  & n15945;
  assign n15948 = ~n15404 & ~n15405;
  assign n15949 = po5  & n15948;
  assign n15950 = ~n15410 & ~n15949;
  assign n15951 = n15410 & n15949;
  assign n15952 = ~n15950 & ~n15951;
  assign n15953 = ~n15947 & ~n15952;
  assign n15954 = ~n15946 & ~n15953;
  assign n15955 = po21  & ~n15954;
  assign n15956 = ~po21  & n15954;
  assign n15957 = ~n15413 & ~n15414;
  assign n15958 = po5  & n15957;
  assign n15959 = ~n15419 & ~n15958;
  assign n15960 = n15419 & n15958;
  assign n15961 = ~n15959 & ~n15960;
  assign n15962 = ~n15956 & ~n15961;
  assign n15963 = ~n15955 & ~n15962;
  assign n15964 = po22  & ~n15963;
  assign n15965 = ~po22  & n15963;
  assign n15966 = ~n15422 & ~n15423;
  assign n15967 = po5  & n15966;
  assign n15968 = ~n15428 & ~n15967;
  assign n15969 = n15428 & n15967;
  assign n15970 = ~n15968 & ~n15969;
  assign n15971 = ~n15965 & ~n15970;
  assign n15972 = ~n15964 & ~n15971;
  assign n15973 = po23  & ~n15972;
  assign n15974 = ~po23  & n15972;
  assign n15975 = ~n15431 & ~n15432;
  assign n15976 = po5  & n15975;
  assign n15977 = ~n15437 & ~n15976;
  assign n15978 = n15437 & n15976;
  assign n15979 = ~n15977 & ~n15978;
  assign n15980 = ~n15974 & ~n15979;
  assign n15981 = ~n15973 & ~n15980;
  assign n15982 = po24  & ~n15981;
  assign n15983 = ~po24  & n15981;
  assign n15984 = ~n15440 & ~n15441;
  assign n15985 = po5  & n15984;
  assign n15986 = ~n15446 & ~n15985;
  assign n15987 = n15446 & n15985;
  assign n15988 = ~n15986 & ~n15987;
  assign n15989 = ~n15983 & ~n15988;
  assign n15990 = ~n15982 & ~n15989;
  assign n15991 = po25  & ~n15990;
  assign n15992 = ~po25  & n15990;
  assign n15993 = ~n15449 & ~n15450;
  assign n15994 = po5  & n15993;
  assign n15995 = ~n15455 & ~n15994;
  assign n15996 = n15455 & n15994;
  assign n15997 = ~n15995 & ~n15996;
  assign n15998 = ~n15992 & ~n15997;
  assign n15999 = ~n15991 & ~n15998;
  assign n16000 = po26  & ~n15999;
  assign n16001 = ~po26  & n15999;
  assign n16002 = ~n15458 & ~n15459;
  assign n16003 = po5  & n16002;
  assign n16004 = ~n15464 & ~n16003;
  assign n16005 = n15464 & n16003;
  assign n16006 = ~n16004 & ~n16005;
  assign n16007 = ~n16001 & ~n16006;
  assign n16008 = ~n16000 & ~n16007;
  assign n16009 = po27  & ~n16008;
  assign n16010 = ~po27  & n16008;
  assign n16011 = ~n15467 & ~n15468;
  assign n16012 = po5  & n16011;
  assign n16013 = ~n15473 & ~n16012;
  assign n16014 = n15473 & n16012;
  assign n16015 = ~n16013 & ~n16014;
  assign n16016 = ~n16010 & ~n16015;
  assign n16017 = ~n16009 & ~n16016;
  assign n16018 = po28  & ~n16017;
  assign n16019 = ~po28  & n16017;
  assign n16020 = ~n15476 & ~n15477;
  assign n16021 = po5  & n16020;
  assign n16022 = ~n15482 & ~n16021;
  assign n16023 = n15482 & n16021;
  assign n16024 = ~n16022 & ~n16023;
  assign n16025 = ~n16019 & ~n16024;
  assign n16026 = ~n16018 & ~n16025;
  assign n16027 = po29  & ~n16026;
  assign n16028 = ~po29  & n16026;
  assign n16029 = ~n15485 & ~n15486;
  assign n16030 = po5  & n16029;
  assign n16031 = ~n15491 & ~n16030;
  assign n16032 = n15491 & n16030;
  assign n16033 = ~n16031 & ~n16032;
  assign n16034 = ~n16028 & ~n16033;
  assign n16035 = ~n16027 & ~n16034;
  assign n16036 = po30  & ~n16035;
  assign n16037 = ~po30  & n16035;
  assign n16038 = ~n15494 & ~n15495;
  assign n16039 = po5  & n16038;
  assign n16040 = ~n15500 & ~n16039;
  assign n16041 = n15500 & n16039;
  assign n16042 = ~n16040 & ~n16041;
  assign n16043 = ~n16037 & ~n16042;
  assign n16044 = ~n16036 & ~n16043;
  assign n16045 = po31  & ~n16044;
  assign n16046 = ~po31  & n16044;
  assign n16047 = ~n15503 & ~n15504;
  assign n16048 = po5  & n16047;
  assign n16049 = ~n15509 & ~n16048;
  assign n16050 = n15509 & n16048;
  assign n16051 = ~n16049 & ~n16050;
  assign n16052 = ~n16046 & ~n16051;
  assign n16053 = ~n16045 & ~n16052;
  assign n16054 = po32  & ~n16053;
  assign n16055 = ~po32  & n16053;
  assign n16056 = ~n15512 & ~n15513;
  assign n16057 = po5  & n16056;
  assign n16058 = ~n15518 & ~n16057;
  assign n16059 = n15518 & n16057;
  assign n16060 = ~n16058 & ~n16059;
  assign n16061 = ~n16055 & ~n16060;
  assign n16062 = ~n16054 & ~n16061;
  assign n16063 = po33  & ~n16062;
  assign n16064 = ~po33  & n16062;
  assign n16065 = ~n15521 & ~n15522;
  assign n16066 = po5  & n16065;
  assign n16067 = ~n15527 & ~n16066;
  assign n16068 = n15527 & n16066;
  assign n16069 = ~n16067 & ~n16068;
  assign n16070 = ~n16064 & ~n16069;
  assign n16071 = ~n16063 & ~n16070;
  assign n16072 = po34  & ~n16071;
  assign n16073 = ~po34  & n16071;
  assign n16074 = ~n15530 & ~n15531;
  assign n16075 = po5  & n16074;
  assign n16076 = ~n15536 & ~n16075;
  assign n16077 = n15536 & n16075;
  assign n16078 = ~n16076 & ~n16077;
  assign n16079 = ~n16073 & ~n16078;
  assign n16080 = ~n16072 & ~n16079;
  assign n16081 = po35  & ~n16080;
  assign n16082 = ~po35  & n16080;
  assign n16083 = ~n15539 & ~n15540;
  assign n16084 = po5  & n16083;
  assign n16085 = ~n15545 & ~n16084;
  assign n16086 = n15545 & n16084;
  assign n16087 = ~n16085 & ~n16086;
  assign n16088 = ~n16082 & ~n16087;
  assign n16089 = ~n16081 & ~n16088;
  assign n16090 = po36  & ~n16089;
  assign n16091 = ~po36  & n16089;
  assign n16092 = ~n15548 & ~n15549;
  assign n16093 = po5  & n16092;
  assign n16094 = ~n15554 & ~n16093;
  assign n16095 = n15554 & n16093;
  assign n16096 = ~n16094 & ~n16095;
  assign n16097 = ~n16091 & ~n16096;
  assign n16098 = ~n16090 & ~n16097;
  assign n16099 = po37  & ~n16098;
  assign n16100 = ~po37  & n16098;
  assign n16101 = ~n15557 & ~n15558;
  assign n16102 = po5  & n16101;
  assign n16103 = ~n15563 & ~n16102;
  assign n16104 = n15563 & n16102;
  assign n16105 = ~n16103 & ~n16104;
  assign n16106 = ~n16100 & ~n16105;
  assign n16107 = ~n16099 & ~n16106;
  assign n16108 = po38  & ~n16107;
  assign n16109 = ~po38  & n16107;
  assign n16110 = ~n15566 & ~n15567;
  assign n16111 = po5  & n16110;
  assign n16112 = ~n15572 & ~n16111;
  assign n16113 = n15572 & n16111;
  assign n16114 = ~n16112 & ~n16113;
  assign n16115 = ~n16109 & ~n16114;
  assign n16116 = ~n16108 & ~n16115;
  assign n16117 = po39  & ~n16116;
  assign n16118 = ~po39  & n16116;
  assign n16119 = ~n15575 & ~n15576;
  assign n16120 = po5  & n16119;
  assign n16121 = ~n15581 & ~n16120;
  assign n16122 = n15581 & n16120;
  assign n16123 = ~n16121 & ~n16122;
  assign n16124 = ~n16118 & ~n16123;
  assign n16125 = ~n16117 & ~n16124;
  assign n16126 = po40  & ~n16125;
  assign n16127 = ~po40  & n16125;
  assign n16128 = ~n15584 & ~n15585;
  assign n16129 = po5  & n16128;
  assign n16130 = ~n15590 & ~n16129;
  assign n16131 = n15590 & n16129;
  assign n16132 = ~n16130 & ~n16131;
  assign n16133 = ~n16127 & ~n16132;
  assign n16134 = ~n16126 & ~n16133;
  assign n16135 = po41  & ~n16134;
  assign n16136 = ~po41  & n16134;
  assign n16137 = ~n15593 & ~n15594;
  assign n16138 = po5  & n16137;
  assign n16139 = ~n15599 & ~n16138;
  assign n16140 = n15599 & n16138;
  assign n16141 = ~n16139 & ~n16140;
  assign n16142 = ~n16136 & ~n16141;
  assign n16143 = ~n16135 & ~n16142;
  assign n16144 = po42  & ~n16143;
  assign n16145 = ~po42  & n16143;
  assign n16146 = ~n15602 & ~n15603;
  assign n16147 = po5  & n16146;
  assign n16148 = ~n15608 & ~n16147;
  assign n16149 = n15608 & n16147;
  assign n16150 = ~n16148 & ~n16149;
  assign n16151 = ~n16145 & ~n16150;
  assign n16152 = ~n16144 & ~n16151;
  assign n16153 = po43  & ~n16152;
  assign n16154 = ~po43  & n16152;
  assign n16155 = ~n15611 & ~n15612;
  assign n16156 = po5  & n16155;
  assign n16157 = ~n15617 & ~n16156;
  assign n16158 = n15617 & n16156;
  assign n16159 = ~n16157 & ~n16158;
  assign n16160 = ~n16154 & ~n16159;
  assign n16161 = ~n16153 & ~n16160;
  assign n16162 = po44  & ~n16161;
  assign n16163 = ~po44  & n16161;
  assign n16164 = ~n15620 & ~n15621;
  assign n16165 = po5  & n16164;
  assign n16166 = ~n15626 & ~n16165;
  assign n16167 = n15626 & n16165;
  assign n16168 = ~n16166 & ~n16167;
  assign n16169 = ~n16163 & ~n16168;
  assign n16170 = ~n16162 & ~n16169;
  assign n16171 = po45  & ~n16170;
  assign n16172 = ~po45  & n16170;
  assign n16173 = ~n15629 & ~n15630;
  assign n16174 = po5  & n16173;
  assign n16175 = ~n15635 & ~n16174;
  assign n16176 = n15635 & n16174;
  assign n16177 = ~n16175 & ~n16176;
  assign n16178 = ~n16172 & ~n16177;
  assign n16179 = ~n16171 & ~n16178;
  assign n16180 = po46  & ~n16179;
  assign n16181 = ~po46  & n16179;
  assign n16182 = ~n15638 & ~n15639;
  assign n16183 = po5  & n16182;
  assign n16184 = ~n15644 & ~n16183;
  assign n16185 = n15644 & n16183;
  assign n16186 = ~n16184 & ~n16185;
  assign n16187 = ~n16181 & ~n16186;
  assign n16188 = ~n16180 & ~n16187;
  assign n16189 = po47  & ~n16188;
  assign n16190 = ~po47  & n16188;
  assign n16191 = ~n15647 & ~n15648;
  assign n16192 = po5  & n16191;
  assign n16193 = ~n15653 & ~n16192;
  assign n16194 = n15653 & n16192;
  assign n16195 = ~n16193 & ~n16194;
  assign n16196 = ~n16190 & ~n16195;
  assign n16197 = ~n16189 & ~n16196;
  assign n16198 = po48  & ~n16197;
  assign n16199 = ~po48  & n16197;
  assign n16200 = ~n15656 & ~n15657;
  assign n16201 = po5  & n16200;
  assign n16202 = ~n15662 & ~n16201;
  assign n16203 = n15662 & n16201;
  assign n16204 = ~n16202 & ~n16203;
  assign n16205 = ~n16199 & ~n16204;
  assign n16206 = ~n16198 & ~n16205;
  assign n16207 = po49  & ~n16206;
  assign n16208 = ~po49  & n16206;
  assign n16209 = ~n15665 & ~n15666;
  assign n16210 = po5  & n16209;
  assign n16211 = ~n15671 & ~n16210;
  assign n16212 = n15671 & n16210;
  assign n16213 = ~n16211 & ~n16212;
  assign n16214 = ~n16208 & ~n16213;
  assign n16215 = ~n16207 & ~n16214;
  assign n16216 = po50  & ~n16215;
  assign n16217 = ~po50  & n16215;
  assign n16218 = ~n15674 & ~n15675;
  assign n16219 = po5  & n16218;
  assign n16220 = ~n15680 & ~n16219;
  assign n16221 = n15680 & n16219;
  assign n16222 = ~n16220 & ~n16221;
  assign n16223 = ~n16217 & ~n16222;
  assign n16224 = ~n16216 & ~n16223;
  assign n16225 = po51  & ~n16224;
  assign n16226 = ~po51  & n16224;
  assign n16227 = ~n15683 & ~n15684;
  assign n16228 = po5  & n16227;
  assign n16229 = ~n15689 & ~n16228;
  assign n16230 = n15689 & n16228;
  assign n16231 = ~n16229 & ~n16230;
  assign n16232 = ~n16226 & ~n16231;
  assign n16233 = ~n16225 & ~n16232;
  assign n16234 = po52  & ~n16233;
  assign n16235 = ~po52  & n16233;
  assign n16236 = ~n15692 & ~n15693;
  assign n16237 = po5  & n16236;
  assign n16238 = ~n15698 & ~n16237;
  assign n16239 = n15698 & n16237;
  assign n16240 = ~n16238 & ~n16239;
  assign n16241 = ~n16235 & ~n16240;
  assign n16242 = ~n16234 & ~n16241;
  assign n16243 = po53  & ~n16242;
  assign n16244 = ~po53  & n16242;
  assign n16245 = ~n15701 & ~n15702;
  assign n16246 = po5  & n16245;
  assign n16247 = ~n15707 & ~n16246;
  assign n16248 = n15707 & n16246;
  assign n16249 = ~n16247 & ~n16248;
  assign n16250 = ~n16244 & ~n16249;
  assign n16251 = ~n16243 & ~n16250;
  assign n16252 = po54  & ~n16251;
  assign n16253 = ~po54  & n16251;
  assign n16254 = ~n15710 & ~n15711;
  assign n16255 = po5  & n16254;
  assign n16256 = ~n15716 & ~n16255;
  assign n16257 = n15716 & n16255;
  assign n16258 = ~n16256 & ~n16257;
  assign n16259 = ~n16253 & ~n16258;
  assign n16260 = ~n16252 & ~n16259;
  assign n16261 = po55  & ~n16260;
  assign n16262 = ~po55  & n16260;
  assign n16263 = ~n15719 & ~n15720;
  assign n16264 = po5  & n16263;
  assign n16265 = ~n15725 & ~n16264;
  assign n16266 = n15725 & n16264;
  assign n16267 = ~n16265 & ~n16266;
  assign n16268 = ~n16262 & ~n16267;
  assign n16269 = ~n16261 & ~n16268;
  assign n16270 = po56  & ~n16269;
  assign n16271 = ~po56  & n16269;
  assign n16272 = ~n15728 & ~n15729;
  assign n16273 = po5  & n16272;
  assign n16274 = ~n15734 & ~n16273;
  assign n16275 = n15734 & n16273;
  assign n16276 = ~n16274 & ~n16275;
  assign n16277 = ~n16271 & ~n16276;
  assign n16278 = ~n16270 & ~n16277;
  assign n16279 = po57  & ~n16278;
  assign n16280 = ~po57  & n16278;
  assign n16281 = ~n15737 & ~n15738;
  assign n16282 = po5  & n16281;
  assign n16283 = ~n15743 & ~n16282;
  assign n16284 = n15743 & n16282;
  assign n16285 = ~n16283 & ~n16284;
  assign n16286 = ~n16280 & ~n16285;
  assign n16287 = ~n16279 & ~n16286;
  assign n16288 = po58  & ~n16287;
  assign n16289 = ~po58  & n16287;
  assign n16290 = ~n15746 & ~n15747;
  assign n16291 = po5  & n16290;
  assign n16292 = ~n15752 & ~n16291;
  assign n16293 = n15752 & n16291;
  assign n16294 = ~n16292 & ~n16293;
  assign n16295 = ~n16289 & ~n16294;
  assign n16296 = ~n16288 & ~n16295;
  assign n16297 = po59  & ~n16296;
  assign n16298 = ~n15755 & ~n15761;
  assign n16299 = po5  & n16298;
  assign n16300 = ~n15760 & ~n16299;
  assign n16301 = n15760 & n16299;
  assign n16302 = ~n16300 & ~n16301;
  assign n16303 = ~po59  & n16296;
  assign n16304 = ~n16302 & ~n16303;
  assign n16305 = ~n16297 & ~n16304;
  assign n16306 = po60  & ~n16305;
  assign n16307 = ~po60  & n16305;
  assign n16308 = ~n15811 & ~n16307;
  assign n16309 = ~n16306 & ~n16308;
  assign n16310 = po61  & ~n16309;
  assign n16311 = ~po61  & n16309;
  assign n16312 = ~n15768 & ~n15769;
  assign n16313 = po5  & n16312;
  assign n16314 = ~n15774 & ~n16313;
  assign n16315 = n15774 & n16313;
  assign n16316 = ~n16314 & ~n16315;
  assign n16317 = ~n16311 & ~n16316;
  assign n16318 = ~n16310 & ~n16317;
  assign n16319 = po62  & ~n16318;
  assign n16320 = ~po62  & n16318;
  assign n16321 = ~n15777 & ~n15778;
  assign n16322 = po5  & n16321;
  assign n16323 = ~n15783 & ~n16322;
  assign n16324 = n15783 & n16322;
  assign n16325 = ~n16323 & ~n16324;
  assign n16326 = ~n16320 & ~n16325;
  assign n16327 = ~n16319 & ~n16326;
  assign n16328 = n15816 & n16327;
  assign n16329 = ~n15816 & ~n16327;
  assign n16330 = n15796 & ~n15805;
  assign n16331 = ~n15795 & ~n16330;
  assign n16332 = n16329 & n16331;
  assign n16333 = ~po63  & ~n16332;
  assign n16334 = ~n15292 & ~n15805;
  assign n16335 = n15794 & ~n16334;
  assign n16336 = po63  & ~n15796;
  assign n16337 = ~n16335 & n16336;
  assign n16338 = ~n16333 & ~n16337;
  assign po4  = n16328 | ~n16338;
  assign n16340 = ~n16306 & ~n16307;
  assign n16341 = po4  & n16340;
  assign n16342 = ~n15811 & ~n16341;
  assign n16343 = n15811 & n16341;
  assign n16344 = ~n16342 & ~n16343;
  assign n16345 = ~n16319 & ~n16320;
  assign n16346 = po4  & n16345;
  assign n16347 = ~n16325 & ~n16346;
  assign n16348 = n16325 & n16346;
  assign n16349 = ~n16347 & ~n16348;
  assign n16350 = pi8  & po4 ;
  assign n16351 = ~pi6  & ~pi7 ;
  assign n16352 = ~pi8  & n16351;
  assign n16353 = ~n16350 & ~n16352;
  assign n16354 = po5  & ~n16353;
  assign n16355 = ~po5  & n16353;
  assign n16356 = ~pi8  & po4 ;
  assign n16357 = pi9  & ~n16356;
  assign n16358 = n15818 & po4 ;
  assign n16359 = ~n16357 & ~n16358;
  assign n16360 = ~n16355 & n16359;
  assign n16361 = ~n16354 & ~n16360;
  assign n16362 = po6  & ~n16361;
  assign n16363 = ~po6  & n16361;
  assign n16364 = po5  & ~po4 ;
  assign n16365 = ~n16358 & ~n16364;
  assign n16366 = pi10  & ~n16365;
  assign n16367 = ~pi10  & n16365;
  assign n16368 = ~n16366 & ~n16367;
  assign n16369 = ~n16363 & ~n16368;
  assign n16370 = ~n16362 & ~n16369;
  assign n16371 = po7  & ~n16370;
  assign n16372 = ~po7  & n16370;
  assign n16373 = ~n15821 & ~n15822;
  assign n16374 = po4  & n16373;
  assign n16375 = n15826 & ~n16374;
  assign n16376 = ~n15826 & n16374;
  assign n16377 = ~n16375 & ~n16376;
  assign n16378 = ~n16372 & ~n16377;
  assign n16379 = ~n16371 & ~n16378;
  assign n16380 = po8  & ~n16379;
  assign n16381 = ~po8  & n16379;
  assign n16382 = ~n15829 & ~n15830;
  assign n16383 = po4  & n16382;
  assign n16384 = ~n15835 & ~n16383;
  assign n16385 = n15835 & n16383;
  assign n16386 = ~n16384 & ~n16385;
  assign n16387 = ~n16381 & ~n16386;
  assign n16388 = ~n16380 & ~n16387;
  assign n16389 = po9  & ~n16388;
  assign n16390 = ~po9  & n16388;
  assign n16391 = ~n15838 & ~n15839;
  assign n16392 = po4  & n16391;
  assign n16393 = n15844 & n16392;
  assign n16394 = ~n15844 & ~n16392;
  assign n16395 = ~n16393 & ~n16394;
  assign n16396 = ~n16390 & ~n16395;
  assign n16397 = ~n16389 & ~n16396;
  assign n16398 = po10  & ~n16397;
  assign n16399 = ~po10  & n16397;
  assign n16400 = ~n15847 & ~n15848;
  assign n16401 = po4  & n16400;
  assign n16402 = ~n15853 & ~n16401;
  assign n16403 = n15853 & n16401;
  assign n16404 = ~n16402 & ~n16403;
  assign n16405 = ~n16399 & ~n16404;
  assign n16406 = ~n16398 & ~n16405;
  assign n16407 = po11  & ~n16406;
  assign n16408 = ~po11  & n16406;
  assign n16409 = ~n15856 & ~n15857;
  assign n16410 = po4  & n16409;
  assign n16411 = ~n15862 & ~n16410;
  assign n16412 = n15862 & n16410;
  assign n16413 = ~n16411 & ~n16412;
  assign n16414 = ~n16408 & ~n16413;
  assign n16415 = ~n16407 & ~n16414;
  assign n16416 = po12  & ~n16415;
  assign n16417 = ~po12  & n16415;
  assign n16418 = ~n15865 & ~n15866;
  assign n16419 = po4  & n16418;
  assign n16420 = ~n15871 & ~n16419;
  assign n16421 = n15871 & n16419;
  assign n16422 = ~n16420 & ~n16421;
  assign n16423 = ~n16417 & ~n16422;
  assign n16424 = ~n16416 & ~n16423;
  assign n16425 = po13  & ~n16424;
  assign n16426 = ~po13  & n16424;
  assign n16427 = ~n15874 & ~n15875;
  assign n16428 = po4  & n16427;
  assign n16429 = ~n15880 & ~n16428;
  assign n16430 = n15880 & n16428;
  assign n16431 = ~n16429 & ~n16430;
  assign n16432 = ~n16426 & ~n16431;
  assign n16433 = ~n16425 & ~n16432;
  assign n16434 = po14  & ~n16433;
  assign n16435 = ~po14  & n16433;
  assign n16436 = ~n15883 & ~n15884;
  assign n16437 = po4  & n16436;
  assign n16438 = ~n15889 & ~n16437;
  assign n16439 = n15889 & n16437;
  assign n16440 = ~n16438 & ~n16439;
  assign n16441 = ~n16435 & ~n16440;
  assign n16442 = ~n16434 & ~n16441;
  assign n16443 = po15  & ~n16442;
  assign n16444 = ~po15  & n16442;
  assign n16445 = ~n15892 & ~n15893;
  assign n16446 = po4  & n16445;
  assign n16447 = ~n15898 & ~n16446;
  assign n16448 = n15898 & n16446;
  assign n16449 = ~n16447 & ~n16448;
  assign n16450 = ~n16444 & ~n16449;
  assign n16451 = ~n16443 & ~n16450;
  assign n16452 = po16  & ~n16451;
  assign n16453 = ~po16  & n16451;
  assign n16454 = ~n15901 & ~n15902;
  assign n16455 = po4  & n16454;
  assign n16456 = ~n15907 & ~n16455;
  assign n16457 = n15907 & n16455;
  assign n16458 = ~n16456 & ~n16457;
  assign n16459 = ~n16453 & ~n16458;
  assign n16460 = ~n16452 & ~n16459;
  assign n16461 = po17  & ~n16460;
  assign n16462 = ~po17  & n16460;
  assign n16463 = ~n15910 & ~n15911;
  assign n16464 = po4  & n16463;
  assign n16465 = ~n15916 & ~n16464;
  assign n16466 = n15916 & n16464;
  assign n16467 = ~n16465 & ~n16466;
  assign n16468 = ~n16462 & ~n16467;
  assign n16469 = ~n16461 & ~n16468;
  assign n16470 = po18  & ~n16469;
  assign n16471 = ~po18  & n16469;
  assign n16472 = ~n15919 & ~n15920;
  assign n16473 = po4  & n16472;
  assign n16474 = ~n15925 & ~n16473;
  assign n16475 = n15925 & n16473;
  assign n16476 = ~n16474 & ~n16475;
  assign n16477 = ~n16471 & ~n16476;
  assign n16478 = ~n16470 & ~n16477;
  assign n16479 = po19  & ~n16478;
  assign n16480 = ~po19  & n16478;
  assign n16481 = ~n15928 & ~n15929;
  assign n16482 = po4  & n16481;
  assign n16483 = ~n15934 & ~n16482;
  assign n16484 = n15934 & n16482;
  assign n16485 = ~n16483 & ~n16484;
  assign n16486 = ~n16480 & ~n16485;
  assign n16487 = ~n16479 & ~n16486;
  assign n16488 = po20  & ~n16487;
  assign n16489 = ~po20  & n16487;
  assign n16490 = ~n15937 & ~n15938;
  assign n16491 = po4  & n16490;
  assign n16492 = ~n15943 & ~n16491;
  assign n16493 = n15943 & n16491;
  assign n16494 = ~n16492 & ~n16493;
  assign n16495 = ~n16489 & ~n16494;
  assign n16496 = ~n16488 & ~n16495;
  assign n16497 = po21  & ~n16496;
  assign n16498 = ~po21  & n16496;
  assign n16499 = ~n15946 & ~n15947;
  assign n16500 = po4  & n16499;
  assign n16501 = ~n15952 & ~n16500;
  assign n16502 = n15952 & n16500;
  assign n16503 = ~n16501 & ~n16502;
  assign n16504 = ~n16498 & ~n16503;
  assign n16505 = ~n16497 & ~n16504;
  assign n16506 = po22  & ~n16505;
  assign n16507 = ~po22  & n16505;
  assign n16508 = ~n15955 & ~n15956;
  assign n16509 = po4  & n16508;
  assign n16510 = ~n15961 & ~n16509;
  assign n16511 = n15961 & n16509;
  assign n16512 = ~n16510 & ~n16511;
  assign n16513 = ~n16507 & ~n16512;
  assign n16514 = ~n16506 & ~n16513;
  assign n16515 = po23  & ~n16514;
  assign n16516 = ~po23  & n16514;
  assign n16517 = ~n15964 & ~n15965;
  assign n16518 = po4  & n16517;
  assign n16519 = ~n15970 & ~n16518;
  assign n16520 = n15970 & n16518;
  assign n16521 = ~n16519 & ~n16520;
  assign n16522 = ~n16516 & ~n16521;
  assign n16523 = ~n16515 & ~n16522;
  assign n16524 = po24  & ~n16523;
  assign n16525 = ~po24  & n16523;
  assign n16526 = ~n15973 & ~n15974;
  assign n16527 = po4  & n16526;
  assign n16528 = ~n15979 & ~n16527;
  assign n16529 = n15979 & n16527;
  assign n16530 = ~n16528 & ~n16529;
  assign n16531 = ~n16525 & ~n16530;
  assign n16532 = ~n16524 & ~n16531;
  assign n16533 = po25  & ~n16532;
  assign n16534 = ~po25  & n16532;
  assign n16535 = ~n15982 & ~n15983;
  assign n16536 = po4  & n16535;
  assign n16537 = ~n15988 & ~n16536;
  assign n16538 = n15988 & n16536;
  assign n16539 = ~n16537 & ~n16538;
  assign n16540 = ~n16534 & ~n16539;
  assign n16541 = ~n16533 & ~n16540;
  assign n16542 = po26  & ~n16541;
  assign n16543 = ~po26  & n16541;
  assign n16544 = ~n15991 & ~n15992;
  assign n16545 = po4  & n16544;
  assign n16546 = ~n15997 & ~n16545;
  assign n16547 = n15997 & n16545;
  assign n16548 = ~n16546 & ~n16547;
  assign n16549 = ~n16543 & ~n16548;
  assign n16550 = ~n16542 & ~n16549;
  assign n16551 = po27  & ~n16550;
  assign n16552 = ~po27  & n16550;
  assign n16553 = ~n16000 & ~n16001;
  assign n16554 = po4  & n16553;
  assign n16555 = ~n16006 & ~n16554;
  assign n16556 = n16006 & n16554;
  assign n16557 = ~n16555 & ~n16556;
  assign n16558 = ~n16552 & ~n16557;
  assign n16559 = ~n16551 & ~n16558;
  assign n16560 = po28  & ~n16559;
  assign n16561 = ~po28  & n16559;
  assign n16562 = ~n16009 & ~n16010;
  assign n16563 = po4  & n16562;
  assign n16564 = ~n16015 & ~n16563;
  assign n16565 = n16015 & n16563;
  assign n16566 = ~n16564 & ~n16565;
  assign n16567 = ~n16561 & ~n16566;
  assign n16568 = ~n16560 & ~n16567;
  assign n16569 = po29  & ~n16568;
  assign n16570 = ~po29  & n16568;
  assign n16571 = ~n16018 & ~n16019;
  assign n16572 = po4  & n16571;
  assign n16573 = ~n16024 & ~n16572;
  assign n16574 = n16024 & n16572;
  assign n16575 = ~n16573 & ~n16574;
  assign n16576 = ~n16570 & ~n16575;
  assign n16577 = ~n16569 & ~n16576;
  assign n16578 = po30  & ~n16577;
  assign n16579 = ~po30  & n16577;
  assign n16580 = ~n16027 & ~n16028;
  assign n16581 = po4  & n16580;
  assign n16582 = ~n16033 & ~n16581;
  assign n16583 = n16033 & n16581;
  assign n16584 = ~n16582 & ~n16583;
  assign n16585 = ~n16579 & ~n16584;
  assign n16586 = ~n16578 & ~n16585;
  assign n16587 = po31  & ~n16586;
  assign n16588 = ~po31  & n16586;
  assign n16589 = ~n16036 & ~n16037;
  assign n16590 = po4  & n16589;
  assign n16591 = ~n16042 & ~n16590;
  assign n16592 = n16042 & n16590;
  assign n16593 = ~n16591 & ~n16592;
  assign n16594 = ~n16588 & ~n16593;
  assign n16595 = ~n16587 & ~n16594;
  assign n16596 = po32  & ~n16595;
  assign n16597 = ~po32  & n16595;
  assign n16598 = ~n16045 & ~n16046;
  assign n16599 = po4  & n16598;
  assign n16600 = ~n16051 & ~n16599;
  assign n16601 = n16051 & n16599;
  assign n16602 = ~n16600 & ~n16601;
  assign n16603 = ~n16597 & ~n16602;
  assign n16604 = ~n16596 & ~n16603;
  assign n16605 = po33  & ~n16604;
  assign n16606 = ~po33  & n16604;
  assign n16607 = ~n16054 & ~n16055;
  assign n16608 = po4  & n16607;
  assign n16609 = ~n16060 & ~n16608;
  assign n16610 = n16060 & n16608;
  assign n16611 = ~n16609 & ~n16610;
  assign n16612 = ~n16606 & ~n16611;
  assign n16613 = ~n16605 & ~n16612;
  assign n16614 = po34  & ~n16613;
  assign n16615 = ~po34  & n16613;
  assign n16616 = ~n16063 & ~n16064;
  assign n16617 = po4  & n16616;
  assign n16618 = ~n16069 & ~n16617;
  assign n16619 = n16069 & n16617;
  assign n16620 = ~n16618 & ~n16619;
  assign n16621 = ~n16615 & ~n16620;
  assign n16622 = ~n16614 & ~n16621;
  assign n16623 = po35  & ~n16622;
  assign n16624 = ~po35  & n16622;
  assign n16625 = ~n16072 & ~n16073;
  assign n16626 = po4  & n16625;
  assign n16627 = ~n16078 & ~n16626;
  assign n16628 = n16078 & n16626;
  assign n16629 = ~n16627 & ~n16628;
  assign n16630 = ~n16624 & ~n16629;
  assign n16631 = ~n16623 & ~n16630;
  assign n16632 = po36  & ~n16631;
  assign n16633 = ~po36  & n16631;
  assign n16634 = ~n16081 & ~n16082;
  assign n16635 = po4  & n16634;
  assign n16636 = ~n16087 & ~n16635;
  assign n16637 = n16087 & n16635;
  assign n16638 = ~n16636 & ~n16637;
  assign n16639 = ~n16633 & ~n16638;
  assign n16640 = ~n16632 & ~n16639;
  assign n16641 = po37  & ~n16640;
  assign n16642 = ~po37  & n16640;
  assign n16643 = ~n16090 & ~n16091;
  assign n16644 = po4  & n16643;
  assign n16645 = ~n16096 & ~n16644;
  assign n16646 = n16096 & n16644;
  assign n16647 = ~n16645 & ~n16646;
  assign n16648 = ~n16642 & ~n16647;
  assign n16649 = ~n16641 & ~n16648;
  assign n16650 = po38  & ~n16649;
  assign n16651 = ~po38  & n16649;
  assign n16652 = ~n16099 & ~n16100;
  assign n16653 = po4  & n16652;
  assign n16654 = ~n16105 & ~n16653;
  assign n16655 = n16105 & n16653;
  assign n16656 = ~n16654 & ~n16655;
  assign n16657 = ~n16651 & ~n16656;
  assign n16658 = ~n16650 & ~n16657;
  assign n16659 = po39  & ~n16658;
  assign n16660 = ~po39  & n16658;
  assign n16661 = ~n16108 & ~n16109;
  assign n16662 = po4  & n16661;
  assign n16663 = ~n16114 & ~n16662;
  assign n16664 = n16114 & n16662;
  assign n16665 = ~n16663 & ~n16664;
  assign n16666 = ~n16660 & ~n16665;
  assign n16667 = ~n16659 & ~n16666;
  assign n16668 = po40  & ~n16667;
  assign n16669 = ~po40  & n16667;
  assign n16670 = ~n16117 & ~n16118;
  assign n16671 = po4  & n16670;
  assign n16672 = ~n16123 & ~n16671;
  assign n16673 = n16123 & n16671;
  assign n16674 = ~n16672 & ~n16673;
  assign n16675 = ~n16669 & ~n16674;
  assign n16676 = ~n16668 & ~n16675;
  assign n16677 = po41  & ~n16676;
  assign n16678 = ~po41  & n16676;
  assign n16679 = ~n16126 & ~n16127;
  assign n16680 = po4  & n16679;
  assign n16681 = ~n16132 & ~n16680;
  assign n16682 = n16132 & n16680;
  assign n16683 = ~n16681 & ~n16682;
  assign n16684 = ~n16678 & ~n16683;
  assign n16685 = ~n16677 & ~n16684;
  assign n16686 = po42  & ~n16685;
  assign n16687 = ~po42  & n16685;
  assign n16688 = ~n16135 & ~n16136;
  assign n16689 = po4  & n16688;
  assign n16690 = ~n16141 & ~n16689;
  assign n16691 = n16141 & n16689;
  assign n16692 = ~n16690 & ~n16691;
  assign n16693 = ~n16687 & ~n16692;
  assign n16694 = ~n16686 & ~n16693;
  assign n16695 = po43  & ~n16694;
  assign n16696 = ~po43  & n16694;
  assign n16697 = ~n16144 & ~n16145;
  assign n16698 = po4  & n16697;
  assign n16699 = ~n16150 & ~n16698;
  assign n16700 = n16150 & n16698;
  assign n16701 = ~n16699 & ~n16700;
  assign n16702 = ~n16696 & ~n16701;
  assign n16703 = ~n16695 & ~n16702;
  assign n16704 = po44  & ~n16703;
  assign n16705 = ~po44  & n16703;
  assign n16706 = ~n16153 & ~n16154;
  assign n16707 = po4  & n16706;
  assign n16708 = ~n16159 & ~n16707;
  assign n16709 = n16159 & n16707;
  assign n16710 = ~n16708 & ~n16709;
  assign n16711 = ~n16705 & ~n16710;
  assign n16712 = ~n16704 & ~n16711;
  assign n16713 = po45  & ~n16712;
  assign n16714 = ~po45  & n16712;
  assign n16715 = ~n16162 & ~n16163;
  assign n16716 = po4  & n16715;
  assign n16717 = ~n16168 & ~n16716;
  assign n16718 = n16168 & n16716;
  assign n16719 = ~n16717 & ~n16718;
  assign n16720 = ~n16714 & ~n16719;
  assign n16721 = ~n16713 & ~n16720;
  assign n16722 = po46  & ~n16721;
  assign n16723 = ~po46  & n16721;
  assign n16724 = ~n16171 & ~n16172;
  assign n16725 = po4  & n16724;
  assign n16726 = ~n16177 & ~n16725;
  assign n16727 = n16177 & n16725;
  assign n16728 = ~n16726 & ~n16727;
  assign n16729 = ~n16723 & ~n16728;
  assign n16730 = ~n16722 & ~n16729;
  assign n16731 = po47  & ~n16730;
  assign n16732 = ~po47  & n16730;
  assign n16733 = ~n16180 & ~n16181;
  assign n16734 = po4  & n16733;
  assign n16735 = ~n16186 & ~n16734;
  assign n16736 = n16186 & n16734;
  assign n16737 = ~n16735 & ~n16736;
  assign n16738 = ~n16732 & ~n16737;
  assign n16739 = ~n16731 & ~n16738;
  assign n16740 = po48  & ~n16739;
  assign n16741 = ~po48  & n16739;
  assign n16742 = ~n16189 & ~n16190;
  assign n16743 = po4  & n16742;
  assign n16744 = ~n16195 & ~n16743;
  assign n16745 = n16195 & n16743;
  assign n16746 = ~n16744 & ~n16745;
  assign n16747 = ~n16741 & ~n16746;
  assign n16748 = ~n16740 & ~n16747;
  assign n16749 = po49  & ~n16748;
  assign n16750 = ~po49  & n16748;
  assign n16751 = ~n16198 & ~n16199;
  assign n16752 = po4  & n16751;
  assign n16753 = ~n16204 & ~n16752;
  assign n16754 = n16204 & n16752;
  assign n16755 = ~n16753 & ~n16754;
  assign n16756 = ~n16750 & ~n16755;
  assign n16757 = ~n16749 & ~n16756;
  assign n16758 = po50  & ~n16757;
  assign n16759 = ~po50  & n16757;
  assign n16760 = ~n16207 & ~n16208;
  assign n16761 = po4  & n16760;
  assign n16762 = ~n16213 & ~n16761;
  assign n16763 = n16213 & n16761;
  assign n16764 = ~n16762 & ~n16763;
  assign n16765 = ~n16759 & ~n16764;
  assign n16766 = ~n16758 & ~n16765;
  assign n16767 = po51  & ~n16766;
  assign n16768 = ~po51  & n16766;
  assign n16769 = ~n16216 & ~n16217;
  assign n16770 = po4  & n16769;
  assign n16771 = ~n16222 & ~n16770;
  assign n16772 = n16222 & n16770;
  assign n16773 = ~n16771 & ~n16772;
  assign n16774 = ~n16768 & ~n16773;
  assign n16775 = ~n16767 & ~n16774;
  assign n16776 = po52  & ~n16775;
  assign n16777 = ~po52  & n16775;
  assign n16778 = ~n16225 & ~n16226;
  assign n16779 = po4  & n16778;
  assign n16780 = ~n16231 & ~n16779;
  assign n16781 = n16231 & n16779;
  assign n16782 = ~n16780 & ~n16781;
  assign n16783 = ~n16777 & ~n16782;
  assign n16784 = ~n16776 & ~n16783;
  assign n16785 = po53  & ~n16784;
  assign n16786 = ~po53  & n16784;
  assign n16787 = ~n16234 & ~n16235;
  assign n16788 = po4  & n16787;
  assign n16789 = ~n16240 & ~n16788;
  assign n16790 = n16240 & n16788;
  assign n16791 = ~n16789 & ~n16790;
  assign n16792 = ~n16786 & ~n16791;
  assign n16793 = ~n16785 & ~n16792;
  assign n16794 = po54  & ~n16793;
  assign n16795 = ~po54  & n16793;
  assign n16796 = ~n16243 & ~n16244;
  assign n16797 = po4  & n16796;
  assign n16798 = ~n16249 & ~n16797;
  assign n16799 = n16249 & n16797;
  assign n16800 = ~n16798 & ~n16799;
  assign n16801 = ~n16795 & ~n16800;
  assign n16802 = ~n16794 & ~n16801;
  assign n16803 = po55  & ~n16802;
  assign n16804 = ~po55  & n16802;
  assign n16805 = ~n16252 & ~n16253;
  assign n16806 = po4  & n16805;
  assign n16807 = ~n16258 & ~n16806;
  assign n16808 = n16258 & n16806;
  assign n16809 = ~n16807 & ~n16808;
  assign n16810 = ~n16804 & ~n16809;
  assign n16811 = ~n16803 & ~n16810;
  assign n16812 = po56  & ~n16811;
  assign n16813 = ~po56  & n16811;
  assign n16814 = ~n16261 & ~n16262;
  assign n16815 = po4  & n16814;
  assign n16816 = ~n16267 & ~n16815;
  assign n16817 = n16267 & n16815;
  assign n16818 = ~n16816 & ~n16817;
  assign n16819 = ~n16813 & ~n16818;
  assign n16820 = ~n16812 & ~n16819;
  assign n16821 = po57  & ~n16820;
  assign n16822 = ~po57  & n16820;
  assign n16823 = ~n16270 & ~n16271;
  assign n16824 = po4  & n16823;
  assign n16825 = ~n16276 & ~n16824;
  assign n16826 = n16276 & n16824;
  assign n16827 = ~n16825 & ~n16826;
  assign n16828 = ~n16822 & ~n16827;
  assign n16829 = ~n16821 & ~n16828;
  assign n16830 = po58  & ~n16829;
  assign n16831 = ~po58  & n16829;
  assign n16832 = ~n16279 & ~n16280;
  assign n16833 = po4  & n16832;
  assign n16834 = ~n16285 & ~n16833;
  assign n16835 = n16285 & n16833;
  assign n16836 = ~n16834 & ~n16835;
  assign n16837 = ~n16831 & ~n16836;
  assign n16838 = ~n16830 & ~n16837;
  assign n16839 = po59  & ~n16838;
  assign n16840 = ~po59  & n16838;
  assign n16841 = ~n16288 & ~n16289;
  assign n16842 = po4  & n16841;
  assign n16843 = ~n16294 & ~n16842;
  assign n16844 = n16294 & n16842;
  assign n16845 = ~n16843 & ~n16844;
  assign n16846 = ~n16840 & ~n16845;
  assign n16847 = ~n16839 & ~n16846;
  assign n16848 = po60  & ~n16847;
  assign n16849 = ~n16297 & ~n16303;
  assign n16850 = po4  & n16849;
  assign n16851 = ~n16302 & ~n16850;
  assign n16852 = n16302 & n16850;
  assign n16853 = ~n16851 & ~n16852;
  assign n16854 = ~po60  & n16847;
  assign n16855 = ~n16853 & ~n16854;
  assign n16856 = ~n16848 & ~n16855;
  assign n16857 = po61  & ~n16856;
  assign n16858 = ~po61  & n16856;
  assign n16859 = ~n16344 & ~n16858;
  assign n16860 = ~n16857 & ~n16859;
  assign n16861 = po62  & ~n16860;
  assign n16862 = ~po62  & n16860;
  assign n16863 = ~n16310 & ~n16311;
  assign n16864 = po4  & n16863;
  assign n16865 = ~n16316 & ~n16864;
  assign n16866 = n16316 & n16864;
  assign n16867 = ~n16865 & ~n16866;
  assign n16868 = ~n16862 & ~n16867;
  assign n16869 = ~n16861 & ~n16868;
  assign n16870 = n16349 & n16869;
  assign n16871 = ~n16349 & ~n16869;
  assign n16872 = n16329 & ~n16338;
  assign n16873 = ~n16328 & ~n16872;
  assign n16874 = n16871 & n16873;
  assign n16875 = ~po63  & ~n16874;
  assign n16876 = ~n15816 & ~n16338;
  assign n16877 = n16327 & ~n16876;
  assign n16878 = po63  & ~n16329;
  assign n16879 = ~n16877 & n16878;
  assign n16880 = ~n16875 & ~n16879;
  assign po3  = n16870 | ~n16880;
  assign n16882 = ~n16857 & ~n16858;
  assign n16883 = po3  & n16882;
  assign n16884 = ~n16344 & ~n16883;
  assign n16885 = n16344 & n16883;
  assign n16886 = ~n16884 & ~n16885;
  assign n16887 = ~n16861 & ~n16862;
  assign n16888 = po3  & n16887;
  assign n16889 = ~n16867 & ~n16888;
  assign n16890 = n16867 & n16888;
  assign n16891 = ~n16889 & ~n16890;
  assign n16892 = pi6  & po3 ;
  assign n16893 = ~pi4  & ~pi5 ;
  assign n16894 = ~pi6  & n16893;
  assign n16895 = ~n16892 & ~n16894;
  assign n16896 = po4  & ~n16895;
  assign n16897 = ~po4  & n16895;
  assign n16898 = ~pi6  & po3 ;
  assign n16899 = pi7  & ~n16898;
  assign n16900 = n16351 & po3 ;
  assign n16901 = ~n16899 & ~n16900;
  assign n16902 = ~n16897 & n16901;
  assign n16903 = ~n16896 & ~n16902;
  assign n16904 = po5  & ~n16903;
  assign n16905 = ~po5  & n16903;
  assign n16906 = po4  & ~po3 ;
  assign n16907 = ~n16900 & ~n16906;
  assign n16908 = pi8  & ~n16907;
  assign n16909 = ~pi8  & n16907;
  assign n16910 = ~n16908 & ~n16909;
  assign n16911 = ~n16905 & ~n16910;
  assign n16912 = ~n16904 & ~n16911;
  assign n16913 = po6  & ~n16912;
  assign n16914 = ~po6  & n16912;
  assign n16915 = ~n16354 & ~n16355;
  assign n16916 = po3  & n16915;
  assign n16917 = n16359 & ~n16916;
  assign n16918 = ~n16359 & n16916;
  assign n16919 = ~n16917 & ~n16918;
  assign n16920 = ~n16914 & ~n16919;
  assign n16921 = ~n16913 & ~n16920;
  assign n16922 = po7  & ~n16921;
  assign n16923 = ~po7  & n16921;
  assign n16924 = ~n16362 & ~n16363;
  assign n16925 = po3  & n16924;
  assign n16926 = ~n16368 & ~n16925;
  assign n16927 = n16368 & n16925;
  assign n16928 = ~n16926 & ~n16927;
  assign n16929 = ~n16923 & ~n16928;
  assign n16930 = ~n16922 & ~n16929;
  assign n16931 = po8  & ~n16930;
  assign n16932 = ~po8  & n16930;
  assign n16933 = ~n16371 & ~n16372;
  assign n16934 = po3  & n16933;
  assign n16935 = n16377 & n16934;
  assign n16936 = ~n16377 & ~n16934;
  assign n16937 = ~n16935 & ~n16936;
  assign n16938 = ~n16932 & ~n16937;
  assign n16939 = ~n16931 & ~n16938;
  assign n16940 = po9  & ~n16939;
  assign n16941 = ~po9  & n16939;
  assign n16942 = ~n16380 & ~n16381;
  assign n16943 = po3  & n16942;
  assign n16944 = ~n16386 & ~n16943;
  assign n16945 = n16386 & n16943;
  assign n16946 = ~n16944 & ~n16945;
  assign n16947 = ~n16941 & ~n16946;
  assign n16948 = ~n16940 & ~n16947;
  assign n16949 = po10  & ~n16948;
  assign n16950 = ~po10  & n16948;
  assign n16951 = ~n16389 & ~n16390;
  assign n16952 = po3  & n16951;
  assign n16953 = ~n16395 & ~n16952;
  assign n16954 = n16395 & n16952;
  assign n16955 = ~n16953 & ~n16954;
  assign n16956 = ~n16950 & ~n16955;
  assign n16957 = ~n16949 & ~n16956;
  assign n16958 = po11  & ~n16957;
  assign n16959 = ~po11  & n16957;
  assign n16960 = ~n16398 & ~n16399;
  assign n16961 = po3  & n16960;
  assign n16962 = ~n16404 & ~n16961;
  assign n16963 = n16404 & n16961;
  assign n16964 = ~n16962 & ~n16963;
  assign n16965 = ~n16959 & ~n16964;
  assign n16966 = ~n16958 & ~n16965;
  assign n16967 = po12  & ~n16966;
  assign n16968 = ~po12  & n16966;
  assign n16969 = ~n16407 & ~n16408;
  assign n16970 = po3  & n16969;
  assign n16971 = ~n16413 & ~n16970;
  assign n16972 = n16413 & n16970;
  assign n16973 = ~n16971 & ~n16972;
  assign n16974 = ~n16968 & ~n16973;
  assign n16975 = ~n16967 & ~n16974;
  assign n16976 = po13  & ~n16975;
  assign n16977 = ~po13  & n16975;
  assign n16978 = ~n16416 & ~n16417;
  assign n16979 = po3  & n16978;
  assign n16980 = ~n16422 & ~n16979;
  assign n16981 = n16422 & n16979;
  assign n16982 = ~n16980 & ~n16981;
  assign n16983 = ~n16977 & ~n16982;
  assign n16984 = ~n16976 & ~n16983;
  assign n16985 = po14  & ~n16984;
  assign n16986 = ~po14  & n16984;
  assign n16987 = ~n16425 & ~n16426;
  assign n16988 = po3  & n16987;
  assign n16989 = ~n16431 & ~n16988;
  assign n16990 = n16431 & n16988;
  assign n16991 = ~n16989 & ~n16990;
  assign n16992 = ~n16986 & ~n16991;
  assign n16993 = ~n16985 & ~n16992;
  assign n16994 = po15  & ~n16993;
  assign n16995 = ~po15  & n16993;
  assign n16996 = ~n16434 & ~n16435;
  assign n16997 = po3  & n16996;
  assign n16998 = ~n16440 & ~n16997;
  assign n16999 = n16440 & n16997;
  assign n17000 = ~n16998 & ~n16999;
  assign n17001 = ~n16995 & ~n17000;
  assign n17002 = ~n16994 & ~n17001;
  assign n17003 = po16  & ~n17002;
  assign n17004 = ~po16  & n17002;
  assign n17005 = ~n16443 & ~n16444;
  assign n17006 = po3  & n17005;
  assign n17007 = ~n16449 & ~n17006;
  assign n17008 = n16449 & n17006;
  assign n17009 = ~n17007 & ~n17008;
  assign n17010 = ~n17004 & ~n17009;
  assign n17011 = ~n17003 & ~n17010;
  assign n17012 = po17  & ~n17011;
  assign n17013 = ~po17  & n17011;
  assign n17014 = ~n16452 & ~n16453;
  assign n17015 = po3  & n17014;
  assign n17016 = ~n16458 & ~n17015;
  assign n17017 = n16458 & n17015;
  assign n17018 = ~n17016 & ~n17017;
  assign n17019 = ~n17013 & ~n17018;
  assign n17020 = ~n17012 & ~n17019;
  assign n17021 = po18  & ~n17020;
  assign n17022 = ~po18  & n17020;
  assign n17023 = ~n16461 & ~n16462;
  assign n17024 = po3  & n17023;
  assign n17025 = ~n16467 & ~n17024;
  assign n17026 = n16467 & n17024;
  assign n17027 = ~n17025 & ~n17026;
  assign n17028 = ~n17022 & ~n17027;
  assign n17029 = ~n17021 & ~n17028;
  assign n17030 = po19  & ~n17029;
  assign n17031 = ~po19  & n17029;
  assign n17032 = ~n16470 & ~n16471;
  assign n17033 = po3  & n17032;
  assign n17034 = ~n16476 & ~n17033;
  assign n17035 = n16476 & n17033;
  assign n17036 = ~n17034 & ~n17035;
  assign n17037 = ~n17031 & ~n17036;
  assign n17038 = ~n17030 & ~n17037;
  assign n17039 = po20  & ~n17038;
  assign n17040 = ~po20  & n17038;
  assign n17041 = ~n16479 & ~n16480;
  assign n17042 = po3  & n17041;
  assign n17043 = ~n16485 & ~n17042;
  assign n17044 = n16485 & n17042;
  assign n17045 = ~n17043 & ~n17044;
  assign n17046 = ~n17040 & ~n17045;
  assign n17047 = ~n17039 & ~n17046;
  assign n17048 = po21  & ~n17047;
  assign n17049 = ~po21  & n17047;
  assign n17050 = ~n16488 & ~n16489;
  assign n17051 = po3  & n17050;
  assign n17052 = ~n16494 & ~n17051;
  assign n17053 = n16494 & n17051;
  assign n17054 = ~n17052 & ~n17053;
  assign n17055 = ~n17049 & ~n17054;
  assign n17056 = ~n17048 & ~n17055;
  assign n17057 = po22  & ~n17056;
  assign n17058 = ~po22  & n17056;
  assign n17059 = ~n16497 & ~n16498;
  assign n17060 = po3  & n17059;
  assign n17061 = ~n16503 & ~n17060;
  assign n17062 = n16503 & n17060;
  assign n17063 = ~n17061 & ~n17062;
  assign n17064 = ~n17058 & ~n17063;
  assign n17065 = ~n17057 & ~n17064;
  assign n17066 = po23  & ~n17065;
  assign n17067 = ~po23  & n17065;
  assign n17068 = ~n16506 & ~n16507;
  assign n17069 = po3  & n17068;
  assign n17070 = ~n16512 & ~n17069;
  assign n17071 = n16512 & n17069;
  assign n17072 = ~n17070 & ~n17071;
  assign n17073 = ~n17067 & ~n17072;
  assign n17074 = ~n17066 & ~n17073;
  assign n17075 = po24  & ~n17074;
  assign n17076 = ~po24  & n17074;
  assign n17077 = ~n16515 & ~n16516;
  assign n17078 = po3  & n17077;
  assign n17079 = ~n16521 & ~n17078;
  assign n17080 = n16521 & n17078;
  assign n17081 = ~n17079 & ~n17080;
  assign n17082 = ~n17076 & ~n17081;
  assign n17083 = ~n17075 & ~n17082;
  assign n17084 = po25  & ~n17083;
  assign n17085 = ~po25  & n17083;
  assign n17086 = ~n16524 & ~n16525;
  assign n17087 = po3  & n17086;
  assign n17088 = ~n16530 & ~n17087;
  assign n17089 = n16530 & n17087;
  assign n17090 = ~n17088 & ~n17089;
  assign n17091 = ~n17085 & ~n17090;
  assign n17092 = ~n17084 & ~n17091;
  assign n17093 = po26  & ~n17092;
  assign n17094 = ~po26  & n17092;
  assign n17095 = ~n16533 & ~n16534;
  assign n17096 = po3  & n17095;
  assign n17097 = ~n16539 & ~n17096;
  assign n17098 = n16539 & n17096;
  assign n17099 = ~n17097 & ~n17098;
  assign n17100 = ~n17094 & ~n17099;
  assign n17101 = ~n17093 & ~n17100;
  assign n17102 = po27  & ~n17101;
  assign n17103 = ~po27  & n17101;
  assign n17104 = ~n16542 & ~n16543;
  assign n17105 = po3  & n17104;
  assign n17106 = ~n16548 & ~n17105;
  assign n17107 = n16548 & n17105;
  assign n17108 = ~n17106 & ~n17107;
  assign n17109 = ~n17103 & ~n17108;
  assign n17110 = ~n17102 & ~n17109;
  assign n17111 = po28  & ~n17110;
  assign n17112 = ~po28  & n17110;
  assign n17113 = ~n16551 & ~n16552;
  assign n17114 = po3  & n17113;
  assign n17115 = ~n16557 & ~n17114;
  assign n17116 = n16557 & n17114;
  assign n17117 = ~n17115 & ~n17116;
  assign n17118 = ~n17112 & ~n17117;
  assign n17119 = ~n17111 & ~n17118;
  assign n17120 = po29  & ~n17119;
  assign n17121 = ~po29  & n17119;
  assign n17122 = ~n16560 & ~n16561;
  assign n17123 = po3  & n17122;
  assign n17124 = ~n16566 & ~n17123;
  assign n17125 = n16566 & n17123;
  assign n17126 = ~n17124 & ~n17125;
  assign n17127 = ~n17121 & ~n17126;
  assign n17128 = ~n17120 & ~n17127;
  assign n17129 = po30  & ~n17128;
  assign n17130 = ~po30  & n17128;
  assign n17131 = ~n16569 & ~n16570;
  assign n17132 = po3  & n17131;
  assign n17133 = ~n16575 & ~n17132;
  assign n17134 = n16575 & n17132;
  assign n17135 = ~n17133 & ~n17134;
  assign n17136 = ~n17130 & ~n17135;
  assign n17137 = ~n17129 & ~n17136;
  assign n17138 = po31  & ~n17137;
  assign n17139 = ~po31  & n17137;
  assign n17140 = ~n16578 & ~n16579;
  assign n17141 = po3  & n17140;
  assign n17142 = ~n16584 & ~n17141;
  assign n17143 = n16584 & n17141;
  assign n17144 = ~n17142 & ~n17143;
  assign n17145 = ~n17139 & ~n17144;
  assign n17146 = ~n17138 & ~n17145;
  assign n17147 = po32  & ~n17146;
  assign n17148 = ~po32  & n17146;
  assign n17149 = ~n16587 & ~n16588;
  assign n17150 = po3  & n17149;
  assign n17151 = ~n16593 & ~n17150;
  assign n17152 = n16593 & n17150;
  assign n17153 = ~n17151 & ~n17152;
  assign n17154 = ~n17148 & ~n17153;
  assign n17155 = ~n17147 & ~n17154;
  assign n17156 = po33  & ~n17155;
  assign n17157 = ~po33  & n17155;
  assign n17158 = ~n16596 & ~n16597;
  assign n17159 = po3  & n17158;
  assign n17160 = ~n16602 & ~n17159;
  assign n17161 = n16602 & n17159;
  assign n17162 = ~n17160 & ~n17161;
  assign n17163 = ~n17157 & ~n17162;
  assign n17164 = ~n17156 & ~n17163;
  assign n17165 = po34  & ~n17164;
  assign n17166 = ~po34  & n17164;
  assign n17167 = ~n16605 & ~n16606;
  assign n17168 = po3  & n17167;
  assign n17169 = ~n16611 & ~n17168;
  assign n17170 = n16611 & n17168;
  assign n17171 = ~n17169 & ~n17170;
  assign n17172 = ~n17166 & ~n17171;
  assign n17173 = ~n17165 & ~n17172;
  assign n17174 = po35  & ~n17173;
  assign n17175 = ~po35  & n17173;
  assign n17176 = ~n16614 & ~n16615;
  assign n17177 = po3  & n17176;
  assign n17178 = ~n16620 & ~n17177;
  assign n17179 = n16620 & n17177;
  assign n17180 = ~n17178 & ~n17179;
  assign n17181 = ~n17175 & ~n17180;
  assign n17182 = ~n17174 & ~n17181;
  assign n17183 = po36  & ~n17182;
  assign n17184 = ~po36  & n17182;
  assign n17185 = ~n16623 & ~n16624;
  assign n17186 = po3  & n17185;
  assign n17187 = ~n16629 & ~n17186;
  assign n17188 = n16629 & n17186;
  assign n17189 = ~n17187 & ~n17188;
  assign n17190 = ~n17184 & ~n17189;
  assign n17191 = ~n17183 & ~n17190;
  assign n17192 = po37  & ~n17191;
  assign n17193 = ~po37  & n17191;
  assign n17194 = ~n16632 & ~n16633;
  assign n17195 = po3  & n17194;
  assign n17196 = ~n16638 & ~n17195;
  assign n17197 = n16638 & n17195;
  assign n17198 = ~n17196 & ~n17197;
  assign n17199 = ~n17193 & ~n17198;
  assign n17200 = ~n17192 & ~n17199;
  assign n17201 = po38  & ~n17200;
  assign n17202 = ~po38  & n17200;
  assign n17203 = ~n16641 & ~n16642;
  assign n17204 = po3  & n17203;
  assign n17205 = ~n16647 & ~n17204;
  assign n17206 = n16647 & n17204;
  assign n17207 = ~n17205 & ~n17206;
  assign n17208 = ~n17202 & ~n17207;
  assign n17209 = ~n17201 & ~n17208;
  assign n17210 = po39  & ~n17209;
  assign n17211 = ~po39  & n17209;
  assign n17212 = ~n16650 & ~n16651;
  assign n17213 = po3  & n17212;
  assign n17214 = ~n16656 & ~n17213;
  assign n17215 = n16656 & n17213;
  assign n17216 = ~n17214 & ~n17215;
  assign n17217 = ~n17211 & ~n17216;
  assign n17218 = ~n17210 & ~n17217;
  assign n17219 = po40  & ~n17218;
  assign n17220 = ~po40  & n17218;
  assign n17221 = ~n16659 & ~n16660;
  assign n17222 = po3  & n17221;
  assign n17223 = ~n16665 & ~n17222;
  assign n17224 = n16665 & n17222;
  assign n17225 = ~n17223 & ~n17224;
  assign n17226 = ~n17220 & ~n17225;
  assign n17227 = ~n17219 & ~n17226;
  assign n17228 = po41  & ~n17227;
  assign n17229 = ~po41  & n17227;
  assign n17230 = ~n16668 & ~n16669;
  assign n17231 = po3  & n17230;
  assign n17232 = ~n16674 & ~n17231;
  assign n17233 = n16674 & n17231;
  assign n17234 = ~n17232 & ~n17233;
  assign n17235 = ~n17229 & ~n17234;
  assign n17236 = ~n17228 & ~n17235;
  assign n17237 = po42  & ~n17236;
  assign n17238 = ~po42  & n17236;
  assign n17239 = ~n16677 & ~n16678;
  assign n17240 = po3  & n17239;
  assign n17241 = ~n16683 & ~n17240;
  assign n17242 = n16683 & n17240;
  assign n17243 = ~n17241 & ~n17242;
  assign n17244 = ~n17238 & ~n17243;
  assign n17245 = ~n17237 & ~n17244;
  assign n17246 = po43  & ~n17245;
  assign n17247 = ~po43  & n17245;
  assign n17248 = ~n16686 & ~n16687;
  assign n17249 = po3  & n17248;
  assign n17250 = ~n16692 & ~n17249;
  assign n17251 = n16692 & n17249;
  assign n17252 = ~n17250 & ~n17251;
  assign n17253 = ~n17247 & ~n17252;
  assign n17254 = ~n17246 & ~n17253;
  assign n17255 = po44  & ~n17254;
  assign n17256 = ~po44  & n17254;
  assign n17257 = ~n16695 & ~n16696;
  assign n17258 = po3  & n17257;
  assign n17259 = ~n16701 & ~n17258;
  assign n17260 = n16701 & n17258;
  assign n17261 = ~n17259 & ~n17260;
  assign n17262 = ~n17256 & ~n17261;
  assign n17263 = ~n17255 & ~n17262;
  assign n17264 = po45  & ~n17263;
  assign n17265 = ~po45  & n17263;
  assign n17266 = ~n16704 & ~n16705;
  assign n17267 = po3  & n17266;
  assign n17268 = ~n16710 & ~n17267;
  assign n17269 = n16710 & n17267;
  assign n17270 = ~n17268 & ~n17269;
  assign n17271 = ~n17265 & ~n17270;
  assign n17272 = ~n17264 & ~n17271;
  assign n17273 = po46  & ~n17272;
  assign n17274 = ~po46  & n17272;
  assign n17275 = ~n16713 & ~n16714;
  assign n17276 = po3  & n17275;
  assign n17277 = ~n16719 & ~n17276;
  assign n17278 = n16719 & n17276;
  assign n17279 = ~n17277 & ~n17278;
  assign n17280 = ~n17274 & ~n17279;
  assign n17281 = ~n17273 & ~n17280;
  assign n17282 = po47  & ~n17281;
  assign n17283 = ~po47  & n17281;
  assign n17284 = ~n16722 & ~n16723;
  assign n17285 = po3  & n17284;
  assign n17286 = ~n16728 & ~n17285;
  assign n17287 = n16728 & n17285;
  assign n17288 = ~n17286 & ~n17287;
  assign n17289 = ~n17283 & ~n17288;
  assign n17290 = ~n17282 & ~n17289;
  assign n17291 = po48  & ~n17290;
  assign n17292 = ~po48  & n17290;
  assign n17293 = ~n16731 & ~n16732;
  assign n17294 = po3  & n17293;
  assign n17295 = ~n16737 & ~n17294;
  assign n17296 = n16737 & n17294;
  assign n17297 = ~n17295 & ~n17296;
  assign n17298 = ~n17292 & ~n17297;
  assign n17299 = ~n17291 & ~n17298;
  assign n17300 = po49  & ~n17299;
  assign n17301 = ~po49  & n17299;
  assign n17302 = ~n16740 & ~n16741;
  assign n17303 = po3  & n17302;
  assign n17304 = ~n16746 & ~n17303;
  assign n17305 = n16746 & n17303;
  assign n17306 = ~n17304 & ~n17305;
  assign n17307 = ~n17301 & ~n17306;
  assign n17308 = ~n17300 & ~n17307;
  assign n17309 = po50  & ~n17308;
  assign n17310 = ~po50  & n17308;
  assign n17311 = ~n16749 & ~n16750;
  assign n17312 = po3  & n17311;
  assign n17313 = ~n16755 & ~n17312;
  assign n17314 = n16755 & n17312;
  assign n17315 = ~n17313 & ~n17314;
  assign n17316 = ~n17310 & ~n17315;
  assign n17317 = ~n17309 & ~n17316;
  assign n17318 = po51  & ~n17317;
  assign n17319 = ~po51  & n17317;
  assign n17320 = ~n16758 & ~n16759;
  assign n17321 = po3  & n17320;
  assign n17322 = ~n16764 & ~n17321;
  assign n17323 = n16764 & n17321;
  assign n17324 = ~n17322 & ~n17323;
  assign n17325 = ~n17319 & ~n17324;
  assign n17326 = ~n17318 & ~n17325;
  assign n17327 = po52  & ~n17326;
  assign n17328 = ~po52  & n17326;
  assign n17329 = ~n16767 & ~n16768;
  assign n17330 = po3  & n17329;
  assign n17331 = ~n16773 & ~n17330;
  assign n17332 = n16773 & n17330;
  assign n17333 = ~n17331 & ~n17332;
  assign n17334 = ~n17328 & ~n17333;
  assign n17335 = ~n17327 & ~n17334;
  assign n17336 = po53  & ~n17335;
  assign n17337 = ~po53  & n17335;
  assign n17338 = ~n16776 & ~n16777;
  assign n17339 = po3  & n17338;
  assign n17340 = ~n16782 & ~n17339;
  assign n17341 = n16782 & n17339;
  assign n17342 = ~n17340 & ~n17341;
  assign n17343 = ~n17337 & ~n17342;
  assign n17344 = ~n17336 & ~n17343;
  assign n17345 = po54  & ~n17344;
  assign n17346 = ~po54  & n17344;
  assign n17347 = ~n16785 & ~n16786;
  assign n17348 = po3  & n17347;
  assign n17349 = ~n16791 & ~n17348;
  assign n17350 = n16791 & n17348;
  assign n17351 = ~n17349 & ~n17350;
  assign n17352 = ~n17346 & ~n17351;
  assign n17353 = ~n17345 & ~n17352;
  assign n17354 = po55  & ~n17353;
  assign n17355 = ~po55  & n17353;
  assign n17356 = ~n16794 & ~n16795;
  assign n17357 = po3  & n17356;
  assign n17358 = ~n16800 & ~n17357;
  assign n17359 = n16800 & n17357;
  assign n17360 = ~n17358 & ~n17359;
  assign n17361 = ~n17355 & ~n17360;
  assign n17362 = ~n17354 & ~n17361;
  assign n17363 = po56  & ~n17362;
  assign n17364 = ~po56  & n17362;
  assign n17365 = ~n16803 & ~n16804;
  assign n17366 = po3  & n17365;
  assign n17367 = ~n16809 & ~n17366;
  assign n17368 = n16809 & n17366;
  assign n17369 = ~n17367 & ~n17368;
  assign n17370 = ~n17364 & ~n17369;
  assign n17371 = ~n17363 & ~n17370;
  assign n17372 = po57  & ~n17371;
  assign n17373 = ~po57  & n17371;
  assign n17374 = ~n16812 & ~n16813;
  assign n17375 = po3  & n17374;
  assign n17376 = ~n16818 & ~n17375;
  assign n17377 = n16818 & n17375;
  assign n17378 = ~n17376 & ~n17377;
  assign n17379 = ~n17373 & ~n17378;
  assign n17380 = ~n17372 & ~n17379;
  assign n17381 = po58  & ~n17380;
  assign n17382 = ~po58  & n17380;
  assign n17383 = ~n16821 & ~n16822;
  assign n17384 = po3  & n17383;
  assign n17385 = ~n16827 & ~n17384;
  assign n17386 = n16827 & n17384;
  assign n17387 = ~n17385 & ~n17386;
  assign n17388 = ~n17382 & ~n17387;
  assign n17389 = ~n17381 & ~n17388;
  assign n17390 = po59  & ~n17389;
  assign n17391 = ~po59  & n17389;
  assign n17392 = ~n16830 & ~n16831;
  assign n17393 = po3  & n17392;
  assign n17394 = ~n16836 & ~n17393;
  assign n17395 = n16836 & n17393;
  assign n17396 = ~n17394 & ~n17395;
  assign n17397 = ~n17391 & ~n17396;
  assign n17398 = ~n17390 & ~n17397;
  assign n17399 = po60  & ~n17398;
  assign n17400 = ~po60  & n17398;
  assign n17401 = ~n16839 & ~n16840;
  assign n17402 = po3  & n17401;
  assign n17403 = ~n16845 & ~n17402;
  assign n17404 = n16845 & n17402;
  assign n17405 = ~n17403 & ~n17404;
  assign n17406 = ~n17400 & ~n17405;
  assign n17407 = ~n17399 & ~n17406;
  assign n17408 = po61  & ~n17407;
  assign n17409 = ~n16848 & ~n16854;
  assign n17410 = po3  & n17409;
  assign n17411 = ~n16853 & ~n17410;
  assign n17412 = n16853 & n17410;
  assign n17413 = ~n17411 & ~n17412;
  assign n17414 = ~po61  & n17407;
  assign n17415 = ~n17413 & ~n17414;
  assign n17416 = ~n17408 & ~n17415;
  assign n17417 = po62  & ~n17416;
  assign n17418 = ~po62  & n17416;
  assign n17419 = ~n16886 & ~n17418;
  assign n17420 = ~n17417 & ~n17419;
  assign n17421 = n16891 & n17420;
  assign n17422 = ~n16891 & ~n17420;
  assign n17423 = n16871 & ~n16880;
  assign n17424 = ~n16870 & ~n17423;
  assign n17425 = n17422 & n17424;
  assign n17426 = ~po63  & ~n17425;
  assign n17427 = ~n16349 & ~n16880;
  assign n17428 = n16869 & ~n17427;
  assign n17429 = po63  & ~n16871;
  assign n17430 = ~n17428 & n17429;
  assign n17431 = ~n17426 & ~n17430;
  assign po2  = n17421 | ~n17431;
  assign n17433 = ~n17417 & ~n17418;
  assign n17434 = po2  & n17433;
  assign n17435 = ~n16886 & ~n17434;
  assign n17436 = n16886 & n17434;
  assign n17437 = ~n17435 & ~n17436;
  assign n17438 = pi4  & po2 ;
  assign n17439 = ~pi2  & ~pi3 ;
  assign n17440 = ~pi4  & n17439;
  assign n17441 = ~n17438 & ~n17440;
  assign n17442 = po3  & ~n17441;
  assign n17443 = ~po3  & n17441;
  assign n17444 = ~pi4  & po2 ;
  assign n17445 = pi5  & ~n17444;
  assign n17446 = n16893 & po2 ;
  assign n17447 = ~n17445 & ~n17446;
  assign n17448 = ~n17443 & n17447;
  assign n17449 = ~n17442 & ~n17448;
  assign n17450 = po4  & ~n17449;
  assign n17451 = ~po4  & n17449;
  assign n17452 = po3  & ~po2 ;
  assign n17453 = ~n17446 & ~n17452;
  assign n17454 = pi6  & ~n17453;
  assign n17455 = ~pi6  & n17453;
  assign n17456 = ~n17454 & ~n17455;
  assign n17457 = ~n17451 & ~n17456;
  assign n17458 = ~n17450 & ~n17457;
  assign n17459 = po5  & ~n17458;
  assign n17460 = ~po5  & n17458;
  assign n17461 = ~n16896 & ~n16897;
  assign n17462 = po2  & n17461;
  assign n17463 = n16901 & ~n17462;
  assign n17464 = ~n16901 & n17462;
  assign n17465 = ~n17463 & ~n17464;
  assign n17466 = ~n17460 & ~n17465;
  assign n17467 = ~n17459 & ~n17466;
  assign n17468 = po6  & ~n17467;
  assign n17469 = ~po6  & n17467;
  assign n17470 = ~n16904 & ~n16905;
  assign n17471 = po2  & n17470;
  assign n17472 = ~n16910 & ~n17471;
  assign n17473 = n16910 & n17471;
  assign n17474 = ~n17472 & ~n17473;
  assign n17475 = ~n17469 & ~n17474;
  assign n17476 = ~n17468 & ~n17475;
  assign n17477 = po7  & ~n17476;
  assign n17478 = ~po7  & n17476;
  assign n17479 = ~n16913 & ~n16914;
  assign n17480 = po2  & n17479;
  assign n17481 = n16919 & n17480;
  assign n17482 = ~n16919 & ~n17480;
  assign n17483 = ~n17481 & ~n17482;
  assign n17484 = ~n17478 & ~n17483;
  assign n17485 = ~n17477 & ~n17484;
  assign n17486 = po8  & ~n17485;
  assign n17487 = ~po8  & n17485;
  assign n17488 = ~n16922 & ~n16923;
  assign n17489 = po2  & n17488;
  assign n17490 = ~n16928 & ~n17489;
  assign n17491 = n16928 & n17489;
  assign n17492 = ~n17490 & ~n17491;
  assign n17493 = ~n17487 & ~n17492;
  assign n17494 = ~n17486 & ~n17493;
  assign n17495 = po9  & ~n17494;
  assign n17496 = ~po9  & n17494;
  assign n17497 = ~n16931 & ~n16932;
  assign n17498 = po2  & n17497;
  assign n17499 = ~n16937 & ~n17498;
  assign n17500 = n16937 & n17498;
  assign n17501 = ~n17499 & ~n17500;
  assign n17502 = ~n17496 & ~n17501;
  assign n17503 = ~n17495 & ~n17502;
  assign n17504 = po10  & ~n17503;
  assign n17505 = ~po10  & n17503;
  assign n17506 = ~n16940 & ~n16941;
  assign n17507 = po2  & n17506;
  assign n17508 = ~n16946 & ~n17507;
  assign n17509 = n16946 & n17507;
  assign n17510 = ~n17508 & ~n17509;
  assign n17511 = ~n17505 & ~n17510;
  assign n17512 = ~n17504 & ~n17511;
  assign n17513 = po11  & ~n17512;
  assign n17514 = ~po11  & n17512;
  assign n17515 = ~n16949 & ~n16950;
  assign n17516 = po2  & n17515;
  assign n17517 = ~n16955 & ~n17516;
  assign n17518 = n16955 & n17516;
  assign n17519 = ~n17517 & ~n17518;
  assign n17520 = ~n17514 & ~n17519;
  assign n17521 = ~n17513 & ~n17520;
  assign n17522 = po12  & ~n17521;
  assign n17523 = ~po12  & n17521;
  assign n17524 = ~n16958 & ~n16959;
  assign n17525 = po2  & n17524;
  assign n17526 = ~n16964 & ~n17525;
  assign n17527 = n16964 & n17525;
  assign n17528 = ~n17526 & ~n17527;
  assign n17529 = ~n17523 & ~n17528;
  assign n17530 = ~n17522 & ~n17529;
  assign n17531 = po13  & ~n17530;
  assign n17532 = ~po13  & n17530;
  assign n17533 = ~n16967 & ~n16968;
  assign n17534 = po2  & n17533;
  assign n17535 = ~n16973 & ~n17534;
  assign n17536 = n16973 & n17534;
  assign n17537 = ~n17535 & ~n17536;
  assign n17538 = ~n17532 & ~n17537;
  assign n17539 = ~n17531 & ~n17538;
  assign n17540 = po14  & ~n17539;
  assign n17541 = ~po14  & n17539;
  assign n17542 = ~n16976 & ~n16977;
  assign n17543 = po2  & n17542;
  assign n17544 = ~n16982 & ~n17543;
  assign n17545 = n16982 & n17543;
  assign n17546 = ~n17544 & ~n17545;
  assign n17547 = ~n17541 & ~n17546;
  assign n17548 = ~n17540 & ~n17547;
  assign n17549 = po15  & ~n17548;
  assign n17550 = ~po15  & n17548;
  assign n17551 = ~n16985 & ~n16986;
  assign n17552 = po2  & n17551;
  assign n17553 = ~n16991 & ~n17552;
  assign n17554 = n16991 & n17552;
  assign n17555 = ~n17553 & ~n17554;
  assign n17556 = ~n17550 & ~n17555;
  assign n17557 = ~n17549 & ~n17556;
  assign n17558 = po16  & ~n17557;
  assign n17559 = ~po16  & n17557;
  assign n17560 = ~n16994 & ~n16995;
  assign n17561 = po2  & n17560;
  assign n17562 = ~n17000 & ~n17561;
  assign n17563 = n17000 & n17561;
  assign n17564 = ~n17562 & ~n17563;
  assign n17565 = ~n17559 & ~n17564;
  assign n17566 = ~n17558 & ~n17565;
  assign n17567 = po17  & ~n17566;
  assign n17568 = ~po17  & n17566;
  assign n17569 = ~n17003 & ~n17004;
  assign n17570 = po2  & n17569;
  assign n17571 = ~n17009 & ~n17570;
  assign n17572 = n17009 & n17570;
  assign n17573 = ~n17571 & ~n17572;
  assign n17574 = ~n17568 & ~n17573;
  assign n17575 = ~n17567 & ~n17574;
  assign n17576 = po18  & ~n17575;
  assign n17577 = ~po18  & n17575;
  assign n17578 = ~n17012 & ~n17013;
  assign n17579 = po2  & n17578;
  assign n17580 = ~n17018 & ~n17579;
  assign n17581 = n17018 & n17579;
  assign n17582 = ~n17580 & ~n17581;
  assign n17583 = ~n17577 & ~n17582;
  assign n17584 = ~n17576 & ~n17583;
  assign n17585 = po19  & ~n17584;
  assign n17586 = ~po19  & n17584;
  assign n17587 = ~n17021 & ~n17022;
  assign n17588 = po2  & n17587;
  assign n17589 = ~n17027 & ~n17588;
  assign n17590 = n17027 & n17588;
  assign n17591 = ~n17589 & ~n17590;
  assign n17592 = ~n17586 & ~n17591;
  assign n17593 = ~n17585 & ~n17592;
  assign n17594 = po20  & ~n17593;
  assign n17595 = ~po20  & n17593;
  assign n17596 = ~n17030 & ~n17031;
  assign n17597 = po2  & n17596;
  assign n17598 = ~n17036 & ~n17597;
  assign n17599 = n17036 & n17597;
  assign n17600 = ~n17598 & ~n17599;
  assign n17601 = ~n17595 & ~n17600;
  assign n17602 = ~n17594 & ~n17601;
  assign n17603 = po21  & ~n17602;
  assign n17604 = ~po21  & n17602;
  assign n17605 = ~n17039 & ~n17040;
  assign n17606 = po2  & n17605;
  assign n17607 = ~n17045 & ~n17606;
  assign n17608 = n17045 & n17606;
  assign n17609 = ~n17607 & ~n17608;
  assign n17610 = ~n17604 & ~n17609;
  assign n17611 = ~n17603 & ~n17610;
  assign n17612 = po22  & ~n17611;
  assign n17613 = ~po22  & n17611;
  assign n17614 = ~n17048 & ~n17049;
  assign n17615 = po2  & n17614;
  assign n17616 = ~n17054 & ~n17615;
  assign n17617 = n17054 & n17615;
  assign n17618 = ~n17616 & ~n17617;
  assign n17619 = ~n17613 & ~n17618;
  assign n17620 = ~n17612 & ~n17619;
  assign n17621 = po23  & ~n17620;
  assign n17622 = ~po23  & n17620;
  assign n17623 = ~n17057 & ~n17058;
  assign n17624 = po2  & n17623;
  assign n17625 = ~n17063 & ~n17624;
  assign n17626 = n17063 & n17624;
  assign n17627 = ~n17625 & ~n17626;
  assign n17628 = ~n17622 & ~n17627;
  assign n17629 = ~n17621 & ~n17628;
  assign n17630 = po24  & ~n17629;
  assign n17631 = ~po24  & n17629;
  assign n17632 = ~n17066 & ~n17067;
  assign n17633 = po2  & n17632;
  assign n17634 = ~n17072 & ~n17633;
  assign n17635 = n17072 & n17633;
  assign n17636 = ~n17634 & ~n17635;
  assign n17637 = ~n17631 & ~n17636;
  assign n17638 = ~n17630 & ~n17637;
  assign n17639 = po25  & ~n17638;
  assign n17640 = ~po25  & n17638;
  assign n17641 = ~n17075 & ~n17076;
  assign n17642 = po2  & n17641;
  assign n17643 = ~n17081 & ~n17642;
  assign n17644 = n17081 & n17642;
  assign n17645 = ~n17643 & ~n17644;
  assign n17646 = ~n17640 & ~n17645;
  assign n17647 = ~n17639 & ~n17646;
  assign n17648 = po26  & ~n17647;
  assign n17649 = ~po26  & n17647;
  assign n17650 = ~n17084 & ~n17085;
  assign n17651 = po2  & n17650;
  assign n17652 = ~n17090 & ~n17651;
  assign n17653 = n17090 & n17651;
  assign n17654 = ~n17652 & ~n17653;
  assign n17655 = ~n17649 & ~n17654;
  assign n17656 = ~n17648 & ~n17655;
  assign n17657 = po27  & ~n17656;
  assign n17658 = ~po27  & n17656;
  assign n17659 = ~n17093 & ~n17094;
  assign n17660 = po2  & n17659;
  assign n17661 = ~n17099 & ~n17660;
  assign n17662 = n17099 & n17660;
  assign n17663 = ~n17661 & ~n17662;
  assign n17664 = ~n17658 & ~n17663;
  assign n17665 = ~n17657 & ~n17664;
  assign n17666 = po28  & ~n17665;
  assign n17667 = ~po28  & n17665;
  assign n17668 = ~n17102 & ~n17103;
  assign n17669 = po2  & n17668;
  assign n17670 = ~n17108 & ~n17669;
  assign n17671 = n17108 & n17669;
  assign n17672 = ~n17670 & ~n17671;
  assign n17673 = ~n17667 & ~n17672;
  assign n17674 = ~n17666 & ~n17673;
  assign n17675 = po29  & ~n17674;
  assign n17676 = ~po29  & n17674;
  assign n17677 = ~n17111 & ~n17112;
  assign n17678 = po2  & n17677;
  assign n17679 = ~n17117 & ~n17678;
  assign n17680 = n17117 & n17678;
  assign n17681 = ~n17679 & ~n17680;
  assign n17682 = ~n17676 & ~n17681;
  assign n17683 = ~n17675 & ~n17682;
  assign n17684 = po30  & ~n17683;
  assign n17685 = ~po30  & n17683;
  assign n17686 = ~n17120 & ~n17121;
  assign n17687 = po2  & n17686;
  assign n17688 = ~n17126 & ~n17687;
  assign n17689 = n17126 & n17687;
  assign n17690 = ~n17688 & ~n17689;
  assign n17691 = ~n17685 & ~n17690;
  assign n17692 = ~n17684 & ~n17691;
  assign n17693 = po31  & ~n17692;
  assign n17694 = ~po31  & n17692;
  assign n17695 = ~n17129 & ~n17130;
  assign n17696 = po2  & n17695;
  assign n17697 = ~n17135 & ~n17696;
  assign n17698 = n17135 & n17696;
  assign n17699 = ~n17697 & ~n17698;
  assign n17700 = ~n17694 & ~n17699;
  assign n17701 = ~n17693 & ~n17700;
  assign n17702 = po32  & ~n17701;
  assign n17703 = ~po32  & n17701;
  assign n17704 = ~n17138 & ~n17139;
  assign n17705 = po2  & n17704;
  assign n17706 = ~n17144 & ~n17705;
  assign n17707 = n17144 & n17705;
  assign n17708 = ~n17706 & ~n17707;
  assign n17709 = ~n17703 & ~n17708;
  assign n17710 = ~n17702 & ~n17709;
  assign n17711 = po33  & ~n17710;
  assign n17712 = ~po33  & n17710;
  assign n17713 = ~n17147 & ~n17148;
  assign n17714 = po2  & n17713;
  assign n17715 = ~n17153 & ~n17714;
  assign n17716 = n17153 & n17714;
  assign n17717 = ~n17715 & ~n17716;
  assign n17718 = ~n17712 & ~n17717;
  assign n17719 = ~n17711 & ~n17718;
  assign n17720 = po34  & ~n17719;
  assign n17721 = ~po34  & n17719;
  assign n17722 = ~n17156 & ~n17157;
  assign n17723 = po2  & n17722;
  assign n17724 = ~n17162 & ~n17723;
  assign n17725 = n17162 & n17723;
  assign n17726 = ~n17724 & ~n17725;
  assign n17727 = ~n17721 & ~n17726;
  assign n17728 = ~n17720 & ~n17727;
  assign n17729 = po35  & ~n17728;
  assign n17730 = ~po35  & n17728;
  assign n17731 = ~n17165 & ~n17166;
  assign n17732 = po2  & n17731;
  assign n17733 = ~n17171 & ~n17732;
  assign n17734 = n17171 & n17732;
  assign n17735 = ~n17733 & ~n17734;
  assign n17736 = ~n17730 & ~n17735;
  assign n17737 = ~n17729 & ~n17736;
  assign n17738 = po36  & ~n17737;
  assign n17739 = ~po36  & n17737;
  assign n17740 = ~n17174 & ~n17175;
  assign n17741 = po2  & n17740;
  assign n17742 = ~n17180 & ~n17741;
  assign n17743 = n17180 & n17741;
  assign n17744 = ~n17742 & ~n17743;
  assign n17745 = ~n17739 & ~n17744;
  assign n17746 = ~n17738 & ~n17745;
  assign n17747 = po37  & ~n17746;
  assign n17748 = ~po37  & n17746;
  assign n17749 = ~n17183 & ~n17184;
  assign n17750 = po2  & n17749;
  assign n17751 = ~n17189 & ~n17750;
  assign n17752 = n17189 & n17750;
  assign n17753 = ~n17751 & ~n17752;
  assign n17754 = ~n17748 & ~n17753;
  assign n17755 = ~n17747 & ~n17754;
  assign n17756 = po38  & ~n17755;
  assign n17757 = ~po38  & n17755;
  assign n17758 = ~n17192 & ~n17193;
  assign n17759 = po2  & n17758;
  assign n17760 = ~n17198 & ~n17759;
  assign n17761 = n17198 & n17759;
  assign n17762 = ~n17760 & ~n17761;
  assign n17763 = ~n17757 & ~n17762;
  assign n17764 = ~n17756 & ~n17763;
  assign n17765 = po39  & ~n17764;
  assign n17766 = ~po39  & n17764;
  assign n17767 = ~n17201 & ~n17202;
  assign n17768 = po2  & n17767;
  assign n17769 = ~n17207 & ~n17768;
  assign n17770 = n17207 & n17768;
  assign n17771 = ~n17769 & ~n17770;
  assign n17772 = ~n17766 & ~n17771;
  assign n17773 = ~n17765 & ~n17772;
  assign n17774 = po40  & ~n17773;
  assign n17775 = ~po40  & n17773;
  assign n17776 = ~n17210 & ~n17211;
  assign n17777 = po2  & n17776;
  assign n17778 = ~n17216 & ~n17777;
  assign n17779 = n17216 & n17777;
  assign n17780 = ~n17778 & ~n17779;
  assign n17781 = ~n17775 & ~n17780;
  assign n17782 = ~n17774 & ~n17781;
  assign n17783 = po41  & ~n17782;
  assign n17784 = ~po41  & n17782;
  assign n17785 = ~n17219 & ~n17220;
  assign n17786 = po2  & n17785;
  assign n17787 = ~n17225 & ~n17786;
  assign n17788 = n17225 & n17786;
  assign n17789 = ~n17787 & ~n17788;
  assign n17790 = ~n17784 & ~n17789;
  assign n17791 = ~n17783 & ~n17790;
  assign n17792 = po42  & ~n17791;
  assign n17793 = ~po42  & n17791;
  assign n17794 = ~n17228 & ~n17229;
  assign n17795 = po2  & n17794;
  assign n17796 = ~n17234 & ~n17795;
  assign n17797 = n17234 & n17795;
  assign n17798 = ~n17796 & ~n17797;
  assign n17799 = ~n17793 & ~n17798;
  assign n17800 = ~n17792 & ~n17799;
  assign n17801 = po43  & ~n17800;
  assign n17802 = ~po43  & n17800;
  assign n17803 = ~n17237 & ~n17238;
  assign n17804 = po2  & n17803;
  assign n17805 = ~n17243 & ~n17804;
  assign n17806 = n17243 & n17804;
  assign n17807 = ~n17805 & ~n17806;
  assign n17808 = ~n17802 & ~n17807;
  assign n17809 = ~n17801 & ~n17808;
  assign n17810 = po44  & ~n17809;
  assign n17811 = ~po44  & n17809;
  assign n17812 = ~n17246 & ~n17247;
  assign n17813 = po2  & n17812;
  assign n17814 = ~n17252 & ~n17813;
  assign n17815 = n17252 & n17813;
  assign n17816 = ~n17814 & ~n17815;
  assign n17817 = ~n17811 & ~n17816;
  assign n17818 = ~n17810 & ~n17817;
  assign n17819 = po45  & ~n17818;
  assign n17820 = ~po45  & n17818;
  assign n17821 = ~n17255 & ~n17256;
  assign n17822 = po2  & n17821;
  assign n17823 = ~n17261 & ~n17822;
  assign n17824 = n17261 & n17822;
  assign n17825 = ~n17823 & ~n17824;
  assign n17826 = ~n17820 & ~n17825;
  assign n17827 = ~n17819 & ~n17826;
  assign n17828 = po46  & ~n17827;
  assign n17829 = ~po46  & n17827;
  assign n17830 = ~n17264 & ~n17265;
  assign n17831 = po2  & n17830;
  assign n17832 = ~n17270 & ~n17831;
  assign n17833 = n17270 & n17831;
  assign n17834 = ~n17832 & ~n17833;
  assign n17835 = ~n17829 & ~n17834;
  assign n17836 = ~n17828 & ~n17835;
  assign n17837 = po47  & ~n17836;
  assign n17838 = ~po47  & n17836;
  assign n17839 = ~n17273 & ~n17274;
  assign n17840 = po2  & n17839;
  assign n17841 = ~n17279 & ~n17840;
  assign n17842 = n17279 & n17840;
  assign n17843 = ~n17841 & ~n17842;
  assign n17844 = ~n17838 & ~n17843;
  assign n17845 = ~n17837 & ~n17844;
  assign n17846 = po48  & ~n17845;
  assign n17847 = ~po48  & n17845;
  assign n17848 = ~n17282 & ~n17283;
  assign n17849 = po2  & n17848;
  assign n17850 = ~n17288 & ~n17849;
  assign n17851 = n17288 & n17849;
  assign n17852 = ~n17850 & ~n17851;
  assign n17853 = ~n17847 & ~n17852;
  assign n17854 = ~n17846 & ~n17853;
  assign n17855 = po49  & ~n17854;
  assign n17856 = ~po49  & n17854;
  assign n17857 = ~n17291 & ~n17292;
  assign n17858 = po2  & n17857;
  assign n17859 = ~n17297 & ~n17858;
  assign n17860 = n17297 & n17858;
  assign n17861 = ~n17859 & ~n17860;
  assign n17862 = ~n17856 & ~n17861;
  assign n17863 = ~n17855 & ~n17862;
  assign n17864 = po50  & ~n17863;
  assign n17865 = ~po50  & n17863;
  assign n17866 = ~n17300 & ~n17301;
  assign n17867 = po2  & n17866;
  assign n17868 = ~n17306 & ~n17867;
  assign n17869 = n17306 & n17867;
  assign n17870 = ~n17868 & ~n17869;
  assign n17871 = ~n17865 & ~n17870;
  assign n17872 = ~n17864 & ~n17871;
  assign n17873 = po51  & ~n17872;
  assign n17874 = ~po51  & n17872;
  assign n17875 = ~n17309 & ~n17310;
  assign n17876 = po2  & n17875;
  assign n17877 = ~n17315 & ~n17876;
  assign n17878 = n17315 & n17876;
  assign n17879 = ~n17877 & ~n17878;
  assign n17880 = ~n17874 & ~n17879;
  assign n17881 = ~n17873 & ~n17880;
  assign n17882 = po52  & ~n17881;
  assign n17883 = ~po52  & n17881;
  assign n17884 = ~n17318 & ~n17319;
  assign n17885 = po2  & n17884;
  assign n17886 = ~n17324 & ~n17885;
  assign n17887 = n17324 & n17885;
  assign n17888 = ~n17886 & ~n17887;
  assign n17889 = ~n17883 & ~n17888;
  assign n17890 = ~n17882 & ~n17889;
  assign n17891 = po53  & ~n17890;
  assign n17892 = ~po53  & n17890;
  assign n17893 = ~n17327 & ~n17328;
  assign n17894 = po2  & n17893;
  assign n17895 = ~n17333 & ~n17894;
  assign n17896 = n17333 & n17894;
  assign n17897 = ~n17895 & ~n17896;
  assign n17898 = ~n17892 & ~n17897;
  assign n17899 = ~n17891 & ~n17898;
  assign n17900 = po54  & ~n17899;
  assign n17901 = ~po54  & n17899;
  assign n17902 = ~n17336 & ~n17337;
  assign n17903 = po2  & n17902;
  assign n17904 = ~n17342 & ~n17903;
  assign n17905 = n17342 & n17903;
  assign n17906 = ~n17904 & ~n17905;
  assign n17907 = ~n17901 & ~n17906;
  assign n17908 = ~n17900 & ~n17907;
  assign n17909 = po55  & ~n17908;
  assign n17910 = ~po55  & n17908;
  assign n17911 = ~n17345 & ~n17346;
  assign n17912 = po2  & n17911;
  assign n17913 = ~n17351 & ~n17912;
  assign n17914 = n17351 & n17912;
  assign n17915 = ~n17913 & ~n17914;
  assign n17916 = ~n17910 & ~n17915;
  assign n17917 = ~n17909 & ~n17916;
  assign n17918 = po56  & ~n17917;
  assign n17919 = ~po56  & n17917;
  assign n17920 = ~n17354 & ~n17355;
  assign n17921 = po2  & n17920;
  assign n17922 = ~n17360 & ~n17921;
  assign n17923 = n17360 & n17921;
  assign n17924 = ~n17922 & ~n17923;
  assign n17925 = ~n17919 & ~n17924;
  assign n17926 = ~n17918 & ~n17925;
  assign n17927 = po57  & ~n17926;
  assign n17928 = ~po57  & n17926;
  assign n17929 = ~n17363 & ~n17364;
  assign n17930 = po2  & n17929;
  assign n17931 = ~n17369 & ~n17930;
  assign n17932 = n17369 & n17930;
  assign n17933 = ~n17931 & ~n17932;
  assign n17934 = ~n17928 & ~n17933;
  assign n17935 = ~n17927 & ~n17934;
  assign n17936 = po58  & ~n17935;
  assign n17937 = ~po58  & n17935;
  assign n17938 = ~n17372 & ~n17373;
  assign n17939 = po2  & n17938;
  assign n17940 = ~n17378 & ~n17939;
  assign n17941 = n17378 & n17939;
  assign n17942 = ~n17940 & ~n17941;
  assign n17943 = ~n17937 & ~n17942;
  assign n17944 = ~n17936 & ~n17943;
  assign n17945 = po59  & ~n17944;
  assign n17946 = ~po59  & n17944;
  assign n17947 = ~n17381 & ~n17382;
  assign n17948 = po2  & n17947;
  assign n17949 = ~n17387 & ~n17948;
  assign n17950 = n17387 & n17948;
  assign n17951 = ~n17949 & ~n17950;
  assign n17952 = ~n17946 & ~n17951;
  assign n17953 = ~n17945 & ~n17952;
  assign n17954 = po60  & ~n17953;
  assign n17955 = ~po60  & n17953;
  assign n17956 = ~n17390 & ~n17391;
  assign n17957 = po2  & n17956;
  assign n17958 = ~n17396 & ~n17957;
  assign n17959 = n17396 & n17957;
  assign n17960 = ~n17958 & ~n17959;
  assign n17961 = ~n17955 & ~n17960;
  assign n17962 = ~n17954 & ~n17961;
  assign n17963 = po61  & ~n17962;
  assign n17964 = ~po61  & n17962;
  assign n17965 = ~n17399 & ~n17400;
  assign n17966 = po2  & n17965;
  assign n17967 = ~n17405 & ~n17966;
  assign n17968 = n17405 & n17966;
  assign n17969 = ~n17967 & ~n17968;
  assign n17970 = ~n17964 & ~n17969;
  assign n17971 = ~n17963 & ~n17970;
  assign n17972 = po62  & ~n17971;
  assign n17973 = ~n17408 & ~n17414;
  assign n17974 = po2  & n17973;
  assign n17975 = ~n17413 & ~n17974;
  assign n17976 = n17413 & n17974;
  assign n17977 = ~n17975 & ~n17976;
  assign n17978 = ~po62  & n17971;
  assign n17979 = ~n17977 & ~n17978;
  assign n17980 = ~n17972 & ~n17979;
  assign n17981 = ~n17437 & ~n17980;
  assign n17982 = n17422 & ~n17431;
  assign n17983 = ~n17421 & ~n17982;
  assign n17984 = n17981 & n17983;
  assign n17985 = ~po63  & ~n17984;
  assign n17986 = ~n16891 & ~n17431;
  assign n17987 = n17420 & ~n17986;
  assign n17988 = po63  & ~n17422;
  assign n17989 = ~n17987 & n17988;
  assign n17990 = ~n17985 & ~n17989;
  assign n17991 = ~n17437 & ~n17990;
  assign n17992 = n17980 & ~n17991;
  assign n17993 = po63  & ~n17981;
  assign n17994 = ~n17992 & n17993;
  assign n17995 = n17437 & n17980;
  assign po1  = ~n17990 | n17995;
  assign n17997 = ~n17972 & ~n17978;
  assign n17998 = po1  & n17997;
  assign n17999 = ~n17977 & ~n17998;
  assign n18000 = n17977 & n17998;
  assign n18001 = ~n17999 & ~n18000;
  assign n18002 = ~pi0  & ~pi1 ;
  assign n18003 = ~pi2  & ~n18002;
  assign n18004 = pi2  & ~po1 ;
  assign n18005 = ~n18003 & ~n18004;
  assign n18006 = ~pi2  & po1 ;
  assign n18007 = pi3  & ~n18006;
  assign n18008 = n17439 & po1 ;
  assign n18009 = ~n18007 & ~n18008;
  assign n18010 = ~po2  & ~n18009;
  assign n18011 = n18005 & ~n18010;
  assign n18012 = po2  & n18009;
  assign n18013 = ~n18011 & ~n18012;
  assign n18014 = po2  & ~po1 ;
  assign n18015 = ~n18008 & ~n18014;
  assign n18016 = pi4  & ~n18015;
  assign n18017 = ~pi4  & n18015;
  assign n18018 = ~n18016 & ~n18017;
  assign n18019 = ~po3  & n18018;
  assign n18020 = ~n18013 & ~n18019;
  assign n18021 = po3  & ~n18018;
  assign n18022 = ~n18020 & ~n18021;
  assign n18023 = ~n17442 & ~n17443;
  assign n18024 = po1  & n18023;
  assign n18025 = n17447 & ~n18024;
  assign n18026 = ~n17447 & n18024;
  assign n18027 = ~n18025 & ~n18026;
  assign n18028 = ~po4  & n18027;
  assign n18029 = ~n18022 & ~n18028;
  assign n18030 = po4  & ~n18027;
  assign n18031 = ~n18029 & ~n18030;
  assign n18032 = ~n17450 & ~n17451;
  assign n18033 = po1  & n18032;
  assign n18034 = ~n17456 & ~n18033;
  assign n18035 = n17456 & n18033;
  assign n18036 = ~n18034 & ~n18035;
  assign n18037 = ~po5  & n18036;
  assign n18038 = ~n18031 & ~n18037;
  assign n18039 = po5  & ~n18036;
  assign n18040 = ~n18038 & ~n18039;
  assign n18041 = ~n17459 & ~n17460;
  assign n18042 = po1  & n18041;
  assign n18043 = n17465 & n18042;
  assign n18044 = ~n17465 & ~n18042;
  assign n18045 = ~n18043 & ~n18044;
  assign n18046 = ~po6  & n18045;
  assign n18047 = ~n18040 & ~n18046;
  assign n18048 = po6  & ~n18045;
  assign n18049 = ~n18047 & ~n18048;
  assign n18050 = ~n17468 & ~n17469;
  assign n18051 = po1  & n18050;
  assign n18052 = ~n17474 & ~n18051;
  assign n18053 = n17474 & n18051;
  assign n18054 = ~n18052 & ~n18053;
  assign n18055 = ~po7  & n18054;
  assign n18056 = ~n18049 & ~n18055;
  assign n18057 = po7  & ~n18054;
  assign n18058 = ~n18056 & ~n18057;
  assign n18059 = ~n17477 & ~n17478;
  assign n18060 = po1  & n18059;
  assign n18061 = ~n17483 & ~n18060;
  assign n18062 = n17483 & n18060;
  assign n18063 = ~n18061 & ~n18062;
  assign n18064 = ~po8  & n18063;
  assign n18065 = ~n18058 & ~n18064;
  assign n18066 = po8  & ~n18063;
  assign n18067 = ~n18065 & ~n18066;
  assign n18068 = ~n17486 & ~n17487;
  assign n18069 = po1  & n18068;
  assign n18070 = ~n17492 & ~n18069;
  assign n18071 = n17492 & n18069;
  assign n18072 = ~n18070 & ~n18071;
  assign n18073 = ~po9  & n18072;
  assign n18074 = ~n18067 & ~n18073;
  assign n18075 = po9  & ~n18072;
  assign n18076 = ~n18074 & ~n18075;
  assign n18077 = ~n17495 & ~n17496;
  assign n18078 = po1  & n18077;
  assign n18079 = ~n17501 & ~n18078;
  assign n18080 = n17501 & n18078;
  assign n18081 = ~n18079 & ~n18080;
  assign n18082 = ~po10  & n18081;
  assign n18083 = ~n18076 & ~n18082;
  assign n18084 = po10  & ~n18081;
  assign n18085 = ~n18083 & ~n18084;
  assign n18086 = ~n17504 & ~n17505;
  assign n18087 = po1  & n18086;
  assign n18088 = ~n17510 & ~n18087;
  assign n18089 = n17510 & n18087;
  assign n18090 = ~n18088 & ~n18089;
  assign n18091 = ~po11  & n18090;
  assign n18092 = ~n18085 & ~n18091;
  assign n18093 = po11  & ~n18090;
  assign n18094 = ~n18092 & ~n18093;
  assign n18095 = ~n17513 & ~n17514;
  assign n18096 = po1  & n18095;
  assign n18097 = ~n17519 & ~n18096;
  assign n18098 = n17519 & n18096;
  assign n18099 = ~n18097 & ~n18098;
  assign n18100 = ~po12  & n18099;
  assign n18101 = ~n18094 & ~n18100;
  assign n18102 = po12  & ~n18099;
  assign n18103 = ~n18101 & ~n18102;
  assign n18104 = ~n17522 & ~n17523;
  assign n18105 = po1  & n18104;
  assign n18106 = ~n17528 & ~n18105;
  assign n18107 = n17528 & n18105;
  assign n18108 = ~n18106 & ~n18107;
  assign n18109 = ~po13  & n18108;
  assign n18110 = ~n18103 & ~n18109;
  assign n18111 = po13  & ~n18108;
  assign n18112 = ~n18110 & ~n18111;
  assign n18113 = ~n17531 & ~n17532;
  assign n18114 = po1  & n18113;
  assign n18115 = ~n17537 & ~n18114;
  assign n18116 = n17537 & n18114;
  assign n18117 = ~n18115 & ~n18116;
  assign n18118 = ~po14  & n18117;
  assign n18119 = ~n18112 & ~n18118;
  assign n18120 = po14  & ~n18117;
  assign n18121 = ~n18119 & ~n18120;
  assign n18122 = ~n17540 & ~n17541;
  assign n18123 = po1  & n18122;
  assign n18124 = ~n17546 & ~n18123;
  assign n18125 = n17546 & n18123;
  assign n18126 = ~n18124 & ~n18125;
  assign n18127 = ~po15  & n18126;
  assign n18128 = ~n18121 & ~n18127;
  assign n18129 = po15  & ~n18126;
  assign n18130 = ~n18128 & ~n18129;
  assign n18131 = ~n17549 & ~n17550;
  assign n18132 = po1  & n18131;
  assign n18133 = ~n17555 & ~n18132;
  assign n18134 = n17555 & n18132;
  assign n18135 = ~n18133 & ~n18134;
  assign n18136 = ~po16  & n18135;
  assign n18137 = ~n18130 & ~n18136;
  assign n18138 = po16  & ~n18135;
  assign n18139 = ~n18137 & ~n18138;
  assign n18140 = ~n17558 & ~n17559;
  assign n18141 = po1  & n18140;
  assign n18142 = ~n17564 & ~n18141;
  assign n18143 = n17564 & n18141;
  assign n18144 = ~n18142 & ~n18143;
  assign n18145 = ~po17  & n18144;
  assign n18146 = ~n18139 & ~n18145;
  assign n18147 = po17  & ~n18144;
  assign n18148 = ~n18146 & ~n18147;
  assign n18149 = ~n17567 & ~n17568;
  assign n18150 = po1  & n18149;
  assign n18151 = ~n17573 & ~n18150;
  assign n18152 = n17573 & n18150;
  assign n18153 = ~n18151 & ~n18152;
  assign n18154 = ~po18  & n18153;
  assign n18155 = ~n18148 & ~n18154;
  assign n18156 = po18  & ~n18153;
  assign n18157 = ~n18155 & ~n18156;
  assign n18158 = ~n17576 & ~n17577;
  assign n18159 = po1  & n18158;
  assign n18160 = ~n17582 & ~n18159;
  assign n18161 = n17582 & n18159;
  assign n18162 = ~n18160 & ~n18161;
  assign n18163 = ~po19  & n18162;
  assign n18164 = ~n18157 & ~n18163;
  assign n18165 = po19  & ~n18162;
  assign n18166 = ~n18164 & ~n18165;
  assign n18167 = ~n17585 & ~n17586;
  assign n18168 = po1  & n18167;
  assign n18169 = ~n17591 & ~n18168;
  assign n18170 = n17591 & n18168;
  assign n18171 = ~n18169 & ~n18170;
  assign n18172 = ~po20  & n18171;
  assign n18173 = ~n18166 & ~n18172;
  assign n18174 = po20  & ~n18171;
  assign n18175 = ~n18173 & ~n18174;
  assign n18176 = ~n17594 & ~n17595;
  assign n18177 = po1  & n18176;
  assign n18178 = ~n17600 & ~n18177;
  assign n18179 = n17600 & n18177;
  assign n18180 = ~n18178 & ~n18179;
  assign n18181 = ~po21  & n18180;
  assign n18182 = ~n18175 & ~n18181;
  assign n18183 = po21  & ~n18180;
  assign n18184 = ~n18182 & ~n18183;
  assign n18185 = ~n17603 & ~n17604;
  assign n18186 = po1  & n18185;
  assign n18187 = ~n17609 & ~n18186;
  assign n18188 = n17609 & n18186;
  assign n18189 = ~n18187 & ~n18188;
  assign n18190 = ~po22  & n18189;
  assign n18191 = ~n18184 & ~n18190;
  assign n18192 = po22  & ~n18189;
  assign n18193 = ~n18191 & ~n18192;
  assign n18194 = ~n17612 & ~n17613;
  assign n18195 = po1  & n18194;
  assign n18196 = ~n17618 & ~n18195;
  assign n18197 = n17618 & n18195;
  assign n18198 = ~n18196 & ~n18197;
  assign n18199 = ~po23  & n18198;
  assign n18200 = ~n18193 & ~n18199;
  assign n18201 = po23  & ~n18198;
  assign n18202 = ~n18200 & ~n18201;
  assign n18203 = ~n17621 & ~n17622;
  assign n18204 = po1  & n18203;
  assign n18205 = ~n17627 & ~n18204;
  assign n18206 = n17627 & n18204;
  assign n18207 = ~n18205 & ~n18206;
  assign n18208 = ~po24  & n18207;
  assign n18209 = ~n18202 & ~n18208;
  assign n18210 = po24  & ~n18207;
  assign n18211 = ~n18209 & ~n18210;
  assign n18212 = ~n17630 & ~n17631;
  assign n18213 = po1  & n18212;
  assign n18214 = ~n17636 & ~n18213;
  assign n18215 = n17636 & n18213;
  assign n18216 = ~n18214 & ~n18215;
  assign n18217 = ~po25  & n18216;
  assign n18218 = ~n18211 & ~n18217;
  assign n18219 = po25  & ~n18216;
  assign n18220 = ~n18218 & ~n18219;
  assign n18221 = ~n17639 & ~n17640;
  assign n18222 = po1  & n18221;
  assign n18223 = ~n17645 & ~n18222;
  assign n18224 = n17645 & n18222;
  assign n18225 = ~n18223 & ~n18224;
  assign n18226 = ~po26  & n18225;
  assign n18227 = ~n18220 & ~n18226;
  assign n18228 = po26  & ~n18225;
  assign n18229 = ~n18227 & ~n18228;
  assign n18230 = ~n17648 & ~n17649;
  assign n18231 = po1  & n18230;
  assign n18232 = ~n17654 & ~n18231;
  assign n18233 = n17654 & n18231;
  assign n18234 = ~n18232 & ~n18233;
  assign n18235 = ~po27  & n18234;
  assign n18236 = ~n18229 & ~n18235;
  assign n18237 = po27  & ~n18234;
  assign n18238 = ~n18236 & ~n18237;
  assign n18239 = ~n17657 & ~n17658;
  assign n18240 = po1  & n18239;
  assign n18241 = ~n17663 & ~n18240;
  assign n18242 = n17663 & n18240;
  assign n18243 = ~n18241 & ~n18242;
  assign n18244 = ~po28  & n18243;
  assign n18245 = ~n18238 & ~n18244;
  assign n18246 = po28  & ~n18243;
  assign n18247 = ~n18245 & ~n18246;
  assign n18248 = ~n17666 & ~n17667;
  assign n18249 = po1  & n18248;
  assign n18250 = ~n17672 & ~n18249;
  assign n18251 = n17672 & n18249;
  assign n18252 = ~n18250 & ~n18251;
  assign n18253 = ~po29  & n18252;
  assign n18254 = ~n18247 & ~n18253;
  assign n18255 = po29  & ~n18252;
  assign n18256 = ~n18254 & ~n18255;
  assign n18257 = ~n17675 & ~n17676;
  assign n18258 = po1  & n18257;
  assign n18259 = ~n17681 & ~n18258;
  assign n18260 = n17681 & n18258;
  assign n18261 = ~n18259 & ~n18260;
  assign n18262 = ~po30  & n18261;
  assign n18263 = ~n18256 & ~n18262;
  assign n18264 = po30  & ~n18261;
  assign n18265 = ~n18263 & ~n18264;
  assign n18266 = ~n17684 & ~n17685;
  assign n18267 = po1  & n18266;
  assign n18268 = ~n17690 & ~n18267;
  assign n18269 = n17690 & n18267;
  assign n18270 = ~n18268 & ~n18269;
  assign n18271 = ~po31  & n18270;
  assign n18272 = ~n18265 & ~n18271;
  assign n18273 = po31  & ~n18270;
  assign n18274 = ~n18272 & ~n18273;
  assign n18275 = ~n17693 & ~n17694;
  assign n18276 = po1  & n18275;
  assign n18277 = ~n17699 & ~n18276;
  assign n18278 = n17699 & n18276;
  assign n18279 = ~n18277 & ~n18278;
  assign n18280 = ~po32  & n18279;
  assign n18281 = ~n18274 & ~n18280;
  assign n18282 = po32  & ~n18279;
  assign n18283 = ~n18281 & ~n18282;
  assign n18284 = ~n17702 & ~n17703;
  assign n18285 = po1  & n18284;
  assign n18286 = ~n17708 & ~n18285;
  assign n18287 = n17708 & n18285;
  assign n18288 = ~n18286 & ~n18287;
  assign n18289 = ~po33  & n18288;
  assign n18290 = ~n18283 & ~n18289;
  assign n18291 = po33  & ~n18288;
  assign n18292 = ~n18290 & ~n18291;
  assign n18293 = ~n17711 & ~n17712;
  assign n18294 = po1  & n18293;
  assign n18295 = ~n17717 & ~n18294;
  assign n18296 = n17717 & n18294;
  assign n18297 = ~n18295 & ~n18296;
  assign n18298 = ~po34  & n18297;
  assign n18299 = ~n18292 & ~n18298;
  assign n18300 = po34  & ~n18297;
  assign n18301 = ~n18299 & ~n18300;
  assign n18302 = ~n17720 & ~n17721;
  assign n18303 = po1  & n18302;
  assign n18304 = ~n17726 & ~n18303;
  assign n18305 = n17726 & n18303;
  assign n18306 = ~n18304 & ~n18305;
  assign n18307 = ~po35  & n18306;
  assign n18308 = ~n18301 & ~n18307;
  assign n18309 = po35  & ~n18306;
  assign n18310 = ~n18308 & ~n18309;
  assign n18311 = ~n17729 & ~n17730;
  assign n18312 = po1  & n18311;
  assign n18313 = ~n17735 & ~n18312;
  assign n18314 = n17735 & n18312;
  assign n18315 = ~n18313 & ~n18314;
  assign n18316 = ~po36  & n18315;
  assign n18317 = ~n18310 & ~n18316;
  assign n18318 = po36  & ~n18315;
  assign n18319 = ~n18317 & ~n18318;
  assign n18320 = ~n17738 & ~n17739;
  assign n18321 = po1  & n18320;
  assign n18322 = ~n17744 & ~n18321;
  assign n18323 = n17744 & n18321;
  assign n18324 = ~n18322 & ~n18323;
  assign n18325 = ~po37  & n18324;
  assign n18326 = ~n18319 & ~n18325;
  assign n18327 = po37  & ~n18324;
  assign n18328 = ~n18326 & ~n18327;
  assign n18329 = ~n17747 & ~n17748;
  assign n18330 = po1  & n18329;
  assign n18331 = ~n17753 & ~n18330;
  assign n18332 = n17753 & n18330;
  assign n18333 = ~n18331 & ~n18332;
  assign n18334 = ~po38  & n18333;
  assign n18335 = ~n18328 & ~n18334;
  assign n18336 = po38  & ~n18333;
  assign n18337 = ~n18335 & ~n18336;
  assign n18338 = ~n17756 & ~n17757;
  assign n18339 = po1  & n18338;
  assign n18340 = ~n17762 & ~n18339;
  assign n18341 = n17762 & n18339;
  assign n18342 = ~n18340 & ~n18341;
  assign n18343 = ~po39  & n18342;
  assign n18344 = ~n18337 & ~n18343;
  assign n18345 = po39  & ~n18342;
  assign n18346 = ~n18344 & ~n18345;
  assign n18347 = ~n17765 & ~n17766;
  assign n18348 = po1  & n18347;
  assign n18349 = ~n17771 & ~n18348;
  assign n18350 = n17771 & n18348;
  assign n18351 = ~n18349 & ~n18350;
  assign n18352 = ~po40  & n18351;
  assign n18353 = ~n18346 & ~n18352;
  assign n18354 = po40  & ~n18351;
  assign n18355 = ~n18353 & ~n18354;
  assign n18356 = ~n17774 & ~n17775;
  assign n18357 = po1  & n18356;
  assign n18358 = ~n17780 & ~n18357;
  assign n18359 = n17780 & n18357;
  assign n18360 = ~n18358 & ~n18359;
  assign n18361 = ~po41  & n18360;
  assign n18362 = ~n18355 & ~n18361;
  assign n18363 = po41  & ~n18360;
  assign n18364 = ~n18362 & ~n18363;
  assign n18365 = ~n17783 & ~n17784;
  assign n18366 = po1  & n18365;
  assign n18367 = ~n17789 & ~n18366;
  assign n18368 = n17789 & n18366;
  assign n18369 = ~n18367 & ~n18368;
  assign n18370 = ~po42  & n18369;
  assign n18371 = ~n18364 & ~n18370;
  assign n18372 = po42  & ~n18369;
  assign n18373 = ~n18371 & ~n18372;
  assign n18374 = ~n17792 & ~n17793;
  assign n18375 = po1  & n18374;
  assign n18376 = ~n17798 & ~n18375;
  assign n18377 = n17798 & n18375;
  assign n18378 = ~n18376 & ~n18377;
  assign n18379 = ~po43  & n18378;
  assign n18380 = ~n18373 & ~n18379;
  assign n18381 = po43  & ~n18378;
  assign n18382 = ~n18380 & ~n18381;
  assign n18383 = ~n17801 & ~n17802;
  assign n18384 = po1  & n18383;
  assign n18385 = ~n17807 & ~n18384;
  assign n18386 = n17807 & n18384;
  assign n18387 = ~n18385 & ~n18386;
  assign n18388 = ~po44  & n18387;
  assign n18389 = ~n18382 & ~n18388;
  assign n18390 = po44  & ~n18387;
  assign n18391 = ~n18389 & ~n18390;
  assign n18392 = ~n17810 & ~n17811;
  assign n18393 = po1  & n18392;
  assign n18394 = ~n17816 & ~n18393;
  assign n18395 = n17816 & n18393;
  assign n18396 = ~n18394 & ~n18395;
  assign n18397 = ~po45  & n18396;
  assign n18398 = ~n18391 & ~n18397;
  assign n18399 = po45  & ~n18396;
  assign n18400 = ~n18398 & ~n18399;
  assign n18401 = ~n17819 & ~n17820;
  assign n18402 = po1  & n18401;
  assign n18403 = ~n17825 & ~n18402;
  assign n18404 = n17825 & n18402;
  assign n18405 = ~n18403 & ~n18404;
  assign n18406 = ~po46  & n18405;
  assign n18407 = ~n18400 & ~n18406;
  assign n18408 = po46  & ~n18405;
  assign n18409 = ~n18407 & ~n18408;
  assign n18410 = ~n17828 & ~n17829;
  assign n18411 = po1  & n18410;
  assign n18412 = ~n17834 & ~n18411;
  assign n18413 = n17834 & n18411;
  assign n18414 = ~n18412 & ~n18413;
  assign n18415 = ~po47  & n18414;
  assign n18416 = ~n18409 & ~n18415;
  assign n18417 = po47  & ~n18414;
  assign n18418 = ~n18416 & ~n18417;
  assign n18419 = ~n17837 & ~n17838;
  assign n18420 = po1  & n18419;
  assign n18421 = ~n17843 & ~n18420;
  assign n18422 = n17843 & n18420;
  assign n18423 = ~n18421 & ~n18422;
  assign n18424 = ~po48  & n18423;
  assign n18425 = ~n18418 & ~n18424;
  assign n18426 = po48  & ~n18423;
  assign n18427 = ~n18425 & ~n18426;
  assign n18428 = ~n17846 & ~n17847;
  assign n18429 = po1  & n18428;
  assign n18430 = ~n17852 & ~n18429;
  assign n18431 = n17852 & n18429;
  assign n18432 = ~n18430 & ~n18431;
  assign n18433 = ~po49  & n18432;
  assign n18434 = ~n18427 & ~n18433;
  assign n18435 = po49  & ~n18432;
  assign n18436 = ~n18434 & ~n18435;
  assign n18437 = ~n17855 & ~n17856;
  assign n18438 = po1  & n18437;
  assign n18439 = ~n17861 & ~n18438;
  assign n18440 = n17861 & n18438;
  assign n18441 = ~n18439 & ~n18440;
  assign n18442 = ~po50  & n18441;
  assign n18443 = ~n18436 & ~n18442;
  assign n18444 = po50  & ~n18441;
  assign n18445 = ~n18443 & ~n18444;
  assign n18446 = ~n17864 & ~n17865;
  assign n18447 = po1  & n18446;
  assign n18448 = ~n17870 & ~n18447;
  assign n18449 = n17870 & n18447;
  assign n18450 = ~n18448 & ~n18449;
  assign n18451 = ~po51  & n18450;
  assign n18452 = ~n18445 & ~n18451;
  assign n18453 = po51  & ~n18450;
  assign n18454 = ~n18452 & ~n18453;
  assign n18455 = ~n17873 & ~n17874;
  assign n18456 = po1  & n18455;
  assign n18457 = ~n17879 & ~n18456;
  assign n18458 = n17879 & n18456;
  assign n18459 = ~n18457 & ~n18458;
  assign n18460 = ~po52  & n18459;
  assign n18461 = ~n18454 & ~n18460;
  assign n18462 = po52  & ~n18459;
  assign n18463 = ~n18461 & ~n18462;
  assign n18464 = ~n17882 & ~n17883;
  assign n18465 = po1  & n18464;
  assign n18466 = ~n17888 & ~n18465;
  assign n18467 = n17888 & n18465;
  assign n18468 = ~n18466 & ~n18467;
  assign n18469 = ~po53  & n18468;
  assign n18470 = ~n18463 & ~n18469;
  assign n18471 = po53  & ~n18468;
  assign n18472 = ~n18470 & ~n18471;
  assign n18473 = ~n17891 & ~n17892;
  assign n18474 = po1  & n18473;
  assign n18475 = ~n17897 & ~n18474;
  assign n18476 = n17897 & n18474;
  assign n18477 = ~n18475 & ~n18476;
  assign n18478 = ~po54  & n18477;
  assign n18479 = ~n18472 & ~n18478;
  assign n18480 = po54  & ~n18477;
  assign n18481 = ~n18479 & ~n18480;
  assign n18482 = ~n17900 & ~n17901;
  assign n18483 = po1  & n18482;
  assign n18484 = ~n17906 & ~n18483;
  assign n18485 = n17906 & n18483;
  assign n18486 = ~n18484 & ~n18485;
  assign n18487 = ~po55  & n18486;
  assign n18488 = ~n18481 & ~n18487;
  assign n18489 = po55  & ~n18486;
  assign n18490 = ~n18488 & ~n18489;
  assign n18491 = ~n17909 & ~n17910;
  assign n18492 = po1  & n18491;
  assign n18493 = ~n17915 & ~n18492;
  assign n18494 = n17915 & n18492;
  assign n18495 = ~n18493 & ~n18494;
  assign n18496 = ~po56  & n18495;
  assign n18497 = ~n18490 & ~n18496;
  assign n18498 = po56  & ~n18495;
  assign n18499 = ~n18497 & ~n18498;
  assign n18500 = ~n17918 & ~n17919;
  assign n18501 = po1  & n18500;
  assign n18502 = ~n17924 & ~n18501;
  assign n18503 = n17924 & n18501;
  assign n18504 = ~n18502 & ~n18503;
  assign n18505 = ~po57  & n18504;
  assign n18506 = ~n18499 & ~n18505;
  assign n18507 = po57  & ~n18504;
  assign n18508 = ~n18506 & ~n18507;
  assign n18509 = ~n17927 & ~n17928;
  assign n18510 = po1  & n18509;
  assign n18511 = ~n17933 & ~n18510;
  assign n18512 = n17933 & n18510;
  assign n18513 = ~n18511 & ~n18512;
  assign n18514 = ~po58  & n18513;
  assign n18515 = ~n18508 & ~n18514;
  assign n18516 = po58  & ~n18513;
  assign n18517 = ~n18515 & ~n18516;
  assign n18518 = ~n17936 & ~n17937;
  assign n18519 = po1  & n18518;
  assign n18520 = ~n17942 & ~n18519;
  assign n18521 = n17942 & n18519;
  assign n18522 = ~n18520 & ~n18521;
  assign n18523 = ~po59  & n18522;
  assign n18524 = ~n18517 & ~n18523;
  assign n18525 = po59  & ~n18522;
  assign n18526 = ~n18524 & ~n18525;
  assign n18527 = ~n17945 & ~n17946;
  assign n18528 = po1  & n18527;
  assign n18529 = ~n17951 & ~n18528;
  assign n18530 = n17951 & n18528;
  assign n18531 = ~n18529 & ~n18530;
  assign n18532 = ~po60  & n18531;
  assign n18533 = ~n18526 & ~n18532;
  assign n18534 = po60  & ~n18531;
  assign n18535 = ~n18533 & ~n18534;
  assign n18536 = ~n17954 & ~n17955;
  assign n18537 = po1  & n18536;
  assign n18538 = ~n17960 & ~n18537;
  assign n18539 = n17960 & n18537;
  assign n18540 = ~n18538 & ~n18539;
  assign n18541 = ~po61  & n18540;
  assign n18542 = ~n18535 & ~n18541;
  assign n18543 = po61  & ~n18540;
  assign n18544 = ~n18542 & ~n18543;
  assign n18545 = ~n17963 & ~n17964;
  assign n18546 = po1  & n18545;
  assign n18547 = ~n17969 & ~n18546;
  assign n18548 = n17969 & n18546;
  assign n18549 = ~n18547 & ~n18548;
  assign n18550 = ~po62  & n18549;
  assign n18551 = ~n18544 & ~n18550;
  assign n18552 = po62  & ~n18549;
  assign n18553 = ~n18551 & ~n18552;
  assign n18554 = n18001 & n18553;
  assign n18555 = ~n17995 & ~n18553;
  assign n18556 = ~n17980 & n17991;
  assign n18557 = ~n18001 & ~n18556;
  assign n18558 = n18555 & n18557;
  assign n18559 = ~po63  & ~n18558;
  assign n18560 = ~n18554 & ~n18559;
  assign po0  = n17994 | ~n18560;
endmodule
