module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7;
  wire n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n707,
    n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n735, n736,
    n737, n738, n739, n740, n741, n742, n745,
    n746, n747, n748, n749, n750, n751;
  assign n137 = pi1  & ~pi2 ;
  assign n138 = pi125  & ~pi126 ;
  assign n139 = ~pi127  & ~n138;
  assign n140 = ~pi124  & ~pi125 ;
  assign n141 = ~pi126  & ~pi127 ;
  assign n142 = n140 & n141;
  assign n143 = pi123  & n142;
  assign n144 = n139 & ~n143;
  assign n145 = ~pi121  & ~n144;
  assign n146 = ~pi122  & n142;
  assign n147 = n144 & ~n146;
  assign n148 = pi121  & ~n147;
  assign n149 = ~n145 & ~n148;
  assign n150 = ~pi122  & ~pi123 ;
  assign n151 = ~pi120  & ~pi121 ;
  assign n152 = n150 & n151;
  assign n153 = n142 & n152;
  assign n154 = n149 & ~n153;
  assign n155 = ~pi118  & ~n154;
  assign n156 = pi117  & n155;
  assign n157 = pi119  & n153;
  assign n158 = n149 & ~n157;
  assign n159 = ~n156 & n158;
  assign n160 = ~pi116  & n155;
  assign n161 = pi115  & n160;
  assign n162 = n159 & ~n161;
  assign n163 = ~pi114  & n160;
  assign n164 = n162 & ~n163;
  assign n165 = ~pi112  & ~n164;
  assign n166 = ~pi110  & n165;
  assign n167 = ~pi113  & ~n162;
  assign n168 = pi113  & ~n164;
  assign n169 = ~n167 & ~n168;
  assign n170 = pi111  & n165;
  assign n171 = n169 & ~n170;
  assign n172 = ~n166 & n171;
  assign n173 = ~pi110  & ~pi111 ;
  assign n174 = ~pi109  & n173;
  assign n175 = n169 & n174;
  assign n176 = pi108  & n175;
  assign n177 = ~n172 & ~n176;
  assign n178 = ~pi106  & n177;
  assign n179 = ~pi107  & n175;
  assign n180 = n177 & ~n179;
  assign n181 = pi106  & n180;
  assign n182 = ~n178 & ~n181;
  assign n183 = ~pi106  & ~pi107 ;
  assign n184 = ~pi105  & n183;
  assign n185 = n175 & n184;
  assign n186 = ~n182 & ~n185;
  assign n187 = ~pi104  & ~n182;
  assign n188 = pi103  & n187;
  assign n189 = ~n186 & ~n188;
  assign n190 = ~pi102  & n187;
  assign n191 = n189 & ~n190;
  assign n192 = ~pi102  & ~pi103 ;
  assign n193 = ~pi101  & n192;
  assign n194 = n185 & n193;
  assign n195 = ~n191 & ~n194;
  assign n196 = ~pi100  & ~n191;
  assign n197 = pi99  & n196;
  assign n198 = ~n195 & ~n197;
  assign n199 = ~pi98  & n196;
  assign n200 = n198 & ~n199;
  assign n201 = ~pi98  & ~pi99 ;
  assign n202 = ~pi97  & n201;
  assign n203 = n194 & n202;
  assign n204 = ~n200 & ~n203;
  assign n205 = ~pi96  & ~n200;
  assign n206 = pi95  & n205;
  assign n207 = ~n204 & ~n206;
  assign n208 = ~pi94  & n205;
  assign n209 = n207 & ~n208;
  assign n210 = ~pi94  & ~pi95 ;
  assign n211 = ~pi93  & n210;
  assign n212 = n203 & n211;
  assign n213 = ~n209 & ~n212;
  assign n214 = ~pi92  & ~n209;
  assign n215 = pi91  & n214;
  assign n216 = ~n213 & ~n215;
  assign n217 = ~pi90  & n214;
  assign n218 = n216 & ~n217;
  assign n219 = ~pi90  & ~pi91 ;
  assign n220 = ~pi89  & n219;
  assign n221 = n212 & n220;
  assign n222 = ~n218 & ~n221;
  assign n223 = ~pi88  & ~n218;
  assign n224 = pi87  & n223;
  assign n225 = ~n222 & ~n224;
  assign n226 = ~pi86  & n223;
  assign n227 = n225 & ~n226;
  assign n228 = ~pi86  & ~pi87 ;
  assign n229 = ~pi85  & n228;
  assign n230 = n221 & n229;
  assign n231 = ~n227 & ~n230;
  assign n232 = ~pi84  & ~n227;
  assign n233 = pi83  & n232;
  assign n234 = ~n231 & ~n233;
  assign n235 = ~pi82  & n232;
  assign n236 = n234 & ~n235;
  assign n237 = ~pi82  & ~pi83 ;
  assign n238 = ~pi81  & n237;
  assign n239 = n230 & n238;
  assign n240 = ~n236 & ~n239;
  assign n241 = ~pi80  & ~n236;
  assign n242 = pi79  & n241;
  assign n243 = ~n240 & ~n242;
  assign n244 = ~pi78  & n241;
  assign n245 = n243 & ~n244;
  assign n246 = ~pi78  & ~pi79 ;
  assign n247 = ~pi77  & n246;
  assign n248 = n239 & n247;
  assign n249 = ~n245 & ~n248;
  assign n250 = ~pi76  & ~n245;
  assign n251 = pi75  & n250;
  assign n252 = ~n249 & ~n251;
  assign n253 = ~pi74  & n250;
  assign n254 = n252 & ~n253;
  assign n255 = ~pi74  & ~pi75 ;
  assign n256 = ~pi73  & n255;
  assign n257 = n248 & n256;
  assign n258 = ~n254 & ~n257;
  assign n259 = ~pi72  & ~n254;
  assign n260 = pi71  & n259;
  assign n261 = ~n258 & ~n260;
  assign n262 = ~pi70  & n259;
  assign n263 = n261 & ~n262;
  assign n264 = ~pi70  & ~pi71 ;
  assign n265 = ~pi69  & n264;
  assign n266 = n257 & n265;
  assign n267 = ~n263 & ~n266;
  assign n268 = ~pi68  & ~n263;
  assign n269 = pi67  & n268;
  assign n270 = ~n267 & ~n269;
  assign n271 = ~pi66  & n268;
  assign n272 = n270 & ~n271;
  assign n273 = ~pi66  & ~pi67 ;
  assign n274 = ~pi65  & n273;
  assign n275 = n266 & n274;
  assign n276 = ~n272 & ~n275;
  assign n277 = ~pi64  & ~n272;
  assign n278 = pi63  & n277;
  assign n279 = ~n276 & ~n278;
  assign n280 = ~pi62  & n277;
  assign n281 = n279 & ~n280;
  assign n282 = ~pi62  & ~pi63 ;
  assign n283 = ~pi61  & n282;
  assign n284 = n275 & n283;
  assign n285 = ~n281 & ~n284;
  assign n286 = ~pi60  & ~n281;
  assign n287 = pi59  & n286;
  assign n288 = ~n285 & ~n287;
  assign n289 = ~pi58  & n286;
  assign n290 = n288 & ~n289;
  assign n291 = ~pi58  & ~pi59 ;
  assign n292 = ~pi57  & n291;
  assign n293 = n284 & n292;
  assign n294 = ~n290 & ~n293;
  assign n295 = ~pi56  & ~n290;
  assign n296 = pi55  & n295;
  assign n297 = ~n294 & ~n296;
  assign n298 = ~pi54  & n295;
  assign n299 = n297 & ~n298;
  assign n300 = ~pi54  & ~pi55 ;
  assign n301 = ~pi53  & n300;
  assign n302 = n293 & n301;
  assign n303 = ~n299 & ~n302;
  assign n304 = ~pi52  & ~n299;
  assign n305 = pi51  & n304;
  assign n306 = ~n303 & ~n305;
  assign n307 = ~pi50  & n304;
  assign n308 = n306 & ~n307;
  assign n309 = ~pi50  & ~pi51 ;
  assign n310 = ~pi49  & n309;
  assign n311 = n302 & n310;
  assign n312 = ~n308 & ~n311;
  assign n313 = ~pi48  & ~n308;
  assign n314 = pi47  & n313;
  assign n315 = ~n312 & ~n314;
  assign n316 = ~pi46  & n313;
  assign n317 = n315 & ~n316;
  assign n318 = ~pi46  & ~pi47 ;
  assign n319 = ~pi45  & n318;
  assign n320 = n311 & n319;
  assign n321 = ~n317 & ~n320;
  assign n322 = ~pi44  & ~n317;
  assign n323 = pi43  & n322;
  assign n324 = ~n321 & ~n323;
  assign n325 = ~pi42  & n322;
  assign n326 = n324 & ~n325;
  assign n327 = ~pi42  & ~pi43 ;
  assign n328 = ~pi41  & n327;
  assign n329 = n320 & n328;
  assign n330 = ~n326 & ~n329;
  assign n331 = ~pi40  & ~n326;
  assign n332 = pi39  & n331;
  assign n333 = ~n330 & ~n332;
  assign n334 = ~pi38  & n331;
  assign n335 = n333 & ~n334;
  assign n336 = ~pi38  & ~pi39 ;
  assign n337 = ~pi37  & n336;
  assign n338 = n329 & n337;
  assign n339 = ~n335 & ~n338;
  assign n340 = ~pi36  & ~n335;
  assign n341 = pi35  & n340;
  assign n342 = ~n339 & ~n341;
  assign n343 = ~pi34  & n340;
  assign n344 = n342 & ~n343;
  assign n345 = ~pi34  & ~pi35 ;
  assign n346 = ~pi33  & n345;
  assign n347 = n338 & n346;
  assign n348 = ~n344 & ~n347;
  assign n349 = ~pi32  & ~n344;
  assign n350 = pi31  & n349;
  assign n351 = ~n348 & ~n350;
  assign n352 = ~pi30  & n349;
  assign n353 = n351 & ~n352;
  assign n354 = ~pi30  & ~pi31 ;
  assign n355 = ~pi29  & n354;
  assign n356 = n347 & n355;
  assign n357 = ~n353 & ~n356;
  assign n358 = ~pi28  & ~n353;
  assign n359 = pi27  & n358;
  assign n360 = ~n357 & ~n359;
  assign n361 = ~pi26  & n358;
  assign n362 = n360 & ~n361;
  assign n363 = ~pi26  & ~pi27 ;
  assign n364 = ~pi25  & n363;
  assign n365 = n356 & n364;
  assign n366 = ~n362 & ~n365;
  assign n367 = ~pi24  & ~n362;
  assign n368 = pi23  & n367;
  assign n369 = ~n366 & ~n368;
  assign n370 = ~pi22  & n367;
  assign n371 = n369 & ~n370;
  assign n372 = ~pi22  & ~pi23 ;
  assign n373 = ~pi21  & n372;
  assign n374 = n365 & n373;
  assign n375 = ~n371 & ~n374;
  assign n376 = ~pi20  & ~n371;
  assign n377 = pi19  & n376;
  assign n378 = ~n375 & ~n377;
  assign n379 = ~pi18  & n376;
  assign n380 = n378 & ~n379;
  assign n381 = ~pi18  & ~pi19 ;
  assign n382 = ~pi17  & n381;
  assign n383 = n374 & n382;
  assign n384 = ~n380 & ~n383;
  assign n385 = ~pi16  & ~n380;
  assign n386 = pi15  & n385;
  assign n387 = ~n384 & ~n386;
  assign n388 = ~pi14  & n385;
  assign n389 = n387 & ~n388;
  assign n390 = ~pi14  & ~pi15 ;
  assign n391 = ~pi13  & n390;
  assign n392 = n383 & n391;
  assign n393 = ~n389 & ~n392;
  assign n394 = ~pi12  & ~n389;
  assign n395 = pi11  & n394;
  assign n396 = ~n393 & ~n395;
  assign n397 = ~pi10  & n394;
  assign n398 = n396 & ~n397;
  assign n399 = ~pi10  & ~pi11 ;
  assign n400 = ~pi9  & n399;
  assign n401 = n392 & n400;
  assign n402 = ~n398 & ~n401;
  assign n403 = ~pi8  & ~n398;
  assign n404 = pi7  & n403;
  assign n405 = ~n402 & ~n404;
  assign n406 = ~pi6  & n403;
  assign n407 = n405 & ~n406;
  assign n408 = ~pi6  & ~pi7 ;
  assign n409 = ~pi5  & n408;
  assign n410 = n401 & n409;
  assign n411 = ~n407 & ~n410;
  assign n412 = ~pi4  & ~n407;
  assign n413 = pi3  & n412;
  assign n414 = ~n411 & ~n413;
  assign n415 = ~n137 & n414;
  assign n416 = ~n411 & ~n412;
  assign n417 = n137 & n416;
  assign po0  = ~n415 & ~n417;
  assign n419 = ~pi2  & ~pi3 ;
  assign n420 = n140 & ~n150;
  assign n421 = n141 & ~n420;
  assign n422 = ~n153 & n421;
  assign n423 = ~pi116  & ~pi117 ;
  assign n424 = ~pi118  & ~pi119 ;
  assign n425 = n153 & n424;
  assign n426 = ~n423 & n425;
  assign n427 = ~n422 & ~n426;
  assign n428 = ~pi112  & ~pi113 ;
  assign n429 = ~pi114  & ~pi115 ;
  assign n430 = n425 & n429;
  assign n431 = ~n428 & n430;
  assign n432 = n427 & ~n431;
  assign n433 = n173 & n430;
  assign n434 = ~pi108  & n174;
  assign n435 = n433 & ~n434;
  assign n436 = n432 & ~n435;
  assign n437 = ~pi104  & ~pi105 ;
  assign n438 = n436 & n437;
  assign n439 = ~n192 & n438;
  assign n440 = n183 & n433;
  assign n441 = n436 & ~n440;
  assign n442 = ~n439 & ~n441;
  assign n443 = ~pi100  & ~pi101 ;
  assign n444 = n438 & n443;
  assign n445 = n442 & ~n444;
  assign n446 = n201 & n442;
  assign n447 = ~pi96  & ~pi97 ;
  assign n448 = n446 & ~n447;
  assign n449 = ~n445 & ~n448;
  assign n450 = ~pi92  & ~pi93 ;
  assign n451 = ~n445 & ~n446;
  assign n452 = n210 & ~n451;
  assign n453 = ~n450 & n452;
  assign n454 = n449 & ~n453;
  assign n455 = ~pi88  & ~pi89 ;
  assign n456 = n219 & n452;
  assign n457 = ~n455 & n456;
  assign n458 = n454 & ~n457;
  assign n459 = ~pi84  & ~pi85 ;
  assign n460 = n458 & n459;
  assign n461 = ~n237 & n460;
  assign n462 = n228 & n456;
  assign n463 = n458 & ~n462;
  assign n464 = ~n461 & ~n463;
  assign n465 = ~pi80  & ~pi81 ;
  assign n466 = n460 & n465;
  assign n467 = n464 & ~n466;
  assign n468 = n246 & n464;
  assign n469 = ~pi76  & ~pi77 ;
  assign n470 = n468 & ~n469;
  assign n471 = ~n467 & ~n470;
  assign n472 = ~pi72  & ~pi73 ;
  assign n473 = ~n467 & ~n468;
  assign n474 = n255 & ~n473;
  assign n475 = ~n472 & n474;
  assign n476 = n471 & ~n475;
  assign n477 = ~pi68  & ~pi69 ;
  assign n478 = n264 & n474;
  assign n479 = ~n477 & n478;
  assign n480 = n476 & ~n479;
  assign n481 = ~pi64  & ~pi65 ;
  assign n482 = n480 & n481;
  assign n483 = ~n282 & n482;
  assign n484 = n273 & n478;
  assign n485 = n480 & ~n484;
  assign n486 = ~n483 & ~n485;
  assign n487 = ~pi60  & ~pi61 ;
  assign n488 = n482 & n487;
  assign n489 = n486 & ~n488;
  assign n490 = n291 & n486;
  assign n491 = ~pi56  & ~pi57 ;
  assign n492 = n490 & ~n491;
  assign n493 = ~n489 & ~n492;
  assign n494 = ~pi52  & ~pi53 ;
  assign n495 = ~n489 & ~n490;
  assign n496 = n300 & ~n495;
  assign n497 = ~n494 & n496;
  assign n498 = n493 & ~n497;
  assign n499 = ~pi48  & ~pi49 ;
  assign n500 = n309 & n496;
  assign n501 = ~n499 & n500;
  assign n502 = n498 & ~n501;
  assign n503 = ~pi44  & ~pi45 ;
  assign n504 = n502 & n503;
  assign n505 = ~n327 & n504;
  assign n506 = n318 & n500;
  assign n507 = n502 & ~n506;
  assign n508 = ~n505 & ~n507;
  assign n509 = ~pi40  & ~pi41 ;
  assign n510 = n504 & n509;
  assign n511 = n508 & ~n510;
  assign n512 = n336 & n508;
  assign n513 = ~pi36  & ~pi37 ;
  assign n514 = n512 & ~n513;
  assign n515 = ~n511 & ~n514;
  assign n516 = ~pi32  & ~pi33 ;
  assign n517 = ~n511 & ~n512;
  assign n518 = n345 & ~n517;
  assign n519 = ~n516 & n518;
  assign n520 = n515 & ~n519;
  assign n521 = ~pi28  & ~pi29 ;
  assign n522 = n354 & n518;
  assign n523 = ~n521 & n522;
  assign n524 = n520 & ~n523;
  assign n525 = ~pi24  & ~pi25 ;
  assign n526 = n524 & n525;
  assign n527 = ~n372 & n526;
  assign n528 = n363 & n522;
  assign n529 = n524 & ~n528;
  assign n530 = ~n527 & ~n529;
  assign n531 = ~pi20  & ~pi21 ;
  assign n532 = n526 & n531;
  assign n533 = n530 & ~n532;
  assign n534 = n381 & n530;
  assign n535 = ~pi16  & ~pi17 ;
  assign n536 = n534 & ~n535;
  assign n537 = ~n533 & ~n536;
  assign n538 = ~pi12  & ~pi13 ;
  assign n539 = ~n533 & ~n534;
  assign n540 = n390 & ~n539;
  assign n541 = ~n538 & n540;
  assign n542 = n537 & ~n541;
  assign n543 = ~pi8  & ~pi9 ;
  assign n544 = n399 & n540;
  assign n545 = ~n543 & n544;
  assign n546 = n542 & ~n545;
  assign n547 = ~pi4  & ~pi5 ;
  assign n548 = n408 & n544;
  assign n549 = ~n547 & n548;
  assign n550 = n546 & ~n549;
  assign n551 = ~n419 & ~n550;
  assign n552 = n546 & ~n548;
  assign n553 = n419 & ~n552;
  assign po1  = ~n551 & ~n553;
  assign n555 = ~pi60  & n283;
  assign n556 = n423 & n424;
  assign n557 = n152 & ~n556;
  assign n558 = n142 & ~n557;
  assign n559 = n428 & n429;
  assign n560 = n556 & n559;
  assign n561 = n153 & n560;
  assign n562 = n558 & ~n561;
  assign n563 = ~pi104  & n184;
  assign n564 = n434 & n561;
  assign n565 = ~n563 & n564;
  assign n566 = ~n562 & ~n565;
  assign n567 = ~pi96  & n202;
  assign n568 = ~pi100  & n193;
  assign n569 = n564 & n568;
  assign n570 = ~n567 & n569;
  assign n571 = n566 & ~n570;
  assign n572 = ~pi88  & n220;
  assign n573 = ~pi92  & n211;
  assign n574 = n569 & n573;
  assign n575 = ~n572 & n574;
  assign n576 = n571 & ~n575;
  assign n577 = ~pi80  & n238;
  assign n578 = ~pi84  & n229;
  assign n579 = n574 & n578;
  assign n580 = ~n577 & n579;
  assign n581 = n576 & ~n580;
  assign n582 = ~pi72  & n256;
  assign n583 = ~pi76  & n247;
  assign n584 = n579 & n583;
  assign n585 = ~n582 & n584;
  assign n586 = n581 & ~n585;
  assign n587 = ~pi64  & n274;
  assign n588 = ~pi68  & n265;
  assign n589 = n584 & n588;
  assign n590 = ~n587 & n589;
  assign n591 = n586 & ~n590;
  assign n592 = ~n555 & n591;
  assign n593 = n586 & ~n589;
  assign n594 = n555 & n593;
  assign n595 = ~n592 & ~n594;
  assign n596 = ~pi56  & n292;
  assign n597 = n595 & ~n596;
  assign n598 = ~n591 & n596;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~pi52  & n301;
  assign n601 = n599 & ~n600;
  assign n602 = ~n595 & n600;
  assign n603 = ~n601 & ~n602;
  assign n604 = ~pi48  & n310;
  assign n605 = n603 & ~n604;
  assign n606 = ~n599 & n604;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~pi44  & n319;
  assign n609 = n607 & ~n608;
  assign n610 = ~n603 & n608;
  assign n611 = ~n609 & ~n610;
  assign n612 = ~pi40  & n328;
  assign n613 = n611 & ~n612;
  assign n614 = ~n607 & n612;
  assign n615 = ~n613 & ~n614;
  assign n616 = ~pi36  & n337;
  assign n617 = n615 & ~n616;
  assign n618 = ~n611 & n616;
  assign n619 = ~n617 & ~n618;
  assign n620 = ~pi32  & n346;
  assign n621 = n619 & ~n620;
  assign n622 = ~n615 & n620;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~pi28  & n355;
  assign n625 = n623 & ~n624;
  assign n626 = ~n619 & n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = ~pi24  & n364;
  assign n629 = n627 & ~n628;
  assign n630 = ~n623 & n628;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~pi20  & n373;
  assign n633 = n631 & ~n632;
  assign n634 = ~n627 & n632;
  assign n635 = ~n633 & ~n634;
  assign n636 = ~pi16  & n382;
  assign n637 = n635 & ~n636;
  assign n638 = ~n631 & n636;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~pi12  & n391;
  assign n641 = n639 & ~n640;
  assign n642 = ~n635 & n640;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~pi8  & n400;
  assign n645 = n643 & ~n644;
  assign n646 = ~n639 & n644;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~pi4  & n409;
  assign n649 = n647 & ~n648;
  assign n650 = ~n643 & n648;
  assign po2  = n649 | n650;
  assign n652 = n434 & n563;
  assign n653 = n560 & ~n652;
  assign n654 = n153 & ~n653;
  assign n655 = ~pi102  & n443;
  assign n656 = n567 & n655;
  assign n657 = n654 & ~n656;
  assign n658 = pi103  & n652;
  assign n659 = n560 & ~n658;
  assign n660 = n153 & ~n659;
  assign n661 = n656 & n660;
  assign n662 = ~n657 & ~n661;
  assign n663 = n572 & n573;
  assign n664 = n662 & ~n663;
  assign n665 = ~n654 & n663;
  assign n666 = ~n664 & ~n665;
  assign n667 = n577 & n578;
  assign n668 = n666 & ~n667;
  assign n669 = ~n662 & n667;
  assign n670 = ~n668 & ~n669;
  assign n671 = n582 & n583;
  assign n672 = n670 & ~n671;
  assign n673 = ~n666 & n671;
  assign n674 = ~n672 & ~n673;
  assign n675 = n587 & n588;
  assign n676 = n674 & ~n675;
  assign n677 = ~n670 & n675;
  assign n678 = ~n676 & ~n677;
  assign n679 = n555 & n596;
  assign n680 = n678 & ~n679;
  assign n681 = ~n674 & n679;
  assign n682 = ~n680 & ~n681;
  assign n683 = n600 & n604;
  assign n684 = n682 & ~n683;
  assign n685 = ~n678 & n683;
  assign n686 = ~n684 & ~n685;
  assign n687 = n608 & n612;
  assign n688 = n686 & ~n687;
  assign n689 = ~n682 & n687;
  assign n690 = ~n688 & ~n689;
  assign n691 = n616 & n620;
  assign n692 = n690 & ~n691;
  assign n693 = ~n686 & n691;
  assign n694 = ~n692 & ~n693;
  assign n695 = n624 & n628;
  assign n696 = n694 & ~n695;
  assign n697 = ~n690 & n695;
  assign n698 = ~n696 & ~n697;
  assign n699 = n632 & n636;
  assign n700 = n698 & ~n699;
  assign n701 = ~n694 & n699;
  assign n702 = ~n700 & ~n701;
  assign n703 = n640 & n644;
  assign n704 = n702 & ~n703;
  assign n705 = ~n698 & n703;
  assign po3  = n704 | n705;
  assign n707 = ~pi99  & n568;
  assign n708 = ~pi98  & n447;
  assign n709 = n652 & n708;
  assign n710 = n707 & n709;
  assign n711 = n663 & n667;
  assign n712 = n710 & ~n711;
  assign n713 = n561 & ~n712;
  assign n714 = ~pi78  & n469;
  assign n715 = n582 & n714;
  assign n716 = n675 & n715;
  assign n717 = n713 & ~n716;
  assign n718 = pi79  & n711;
  assign n719 = n710 & ~n718;
  assign n720 = n561 & ~n719;
  assign n721 = n716 & n720;
  assign n722 = ~n717 & ~n721;
  assign n723 = n679 & n683;
  assign n724 = n722 & ~n723;
  assign n725 = ~n713 & n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = n687 & n691;
  assign n728 = n726 & ~n727;
  assign n729 = ~n722 & n727;
  assign n730 = ~n728 & ~n729;
  assign n731 = n695 & n699;
  assign n732 = n730 & ~n731;
  assign n733 = ~n726 & n731;
  assign po4  = n732 | n733;
  assign n735 = n561 & n710;
  assign n736 = ~pi71  & n671;
  assign n737 = ~pi70  & n477;
  assign n738 = n587 & n737;
  assign n739 = n711 & n738;
  assign n740 = n736 & n739;
  assign n741 = n723 & n727;
  assign n742 = n740 & ~n741;
  assign po5  = ~n735 | n742;
  assign po6  = ~n735 | ~n740;
  assign n745 = ~pi0  & ~po6 ;
  assign n746 = n703 & n745;
  assign n747 = ~pi3  & n746;
  assign n748 = ~pi2  & n747;
  assign n749 = n731 & n741;
  assign n750 = n648 & n749;
  assign n751 = ~pi1  & n750;
  assign po7 = ~n748 | ~n751;
endmodule
