module alu4_cl ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    po0, po1, po2, po3, po4, po5  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9;
  output po0, po1, po2, po3, po4, po5;
  wire n17, n18, n19, n20, n21, n22, n23,
    n24, n25, n26, n27, n28, n29, n30, n31,
    n32, n33, n34, n35, n36, n37, n38, n39,
    n40, n41, n42, n43, n44, n45, n46, n47,
    n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63,
    n64, n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102,
    n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172,
    n174, n175, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216,
    n217, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287,
    n288, n289, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n344,
    n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372,
    n373, n374;
  assign n17 = ~pi2 & pi6;
  assign n18 = pi0 & pi2;
  assign n19 = ~pi5 & pi6;
  assign n20 = ~pi7 & n19;
  assign n21 = ~pi4 & n20;
  assign n22 = ~pi6 & pi7;
  assign n23 = ~pi4 & pi5;
  assign n24 = pi5 & pi9;
  assign n25 = ~pi4 & pi9;
  assign n26 = ~n24 & ~n25;
  assign n27 = ~n23 & ~n26;
  assign n28 = n22 & n27;
  assign n29 = ~n21 & ~n28;
  assign n30 = n18 & ~n29;
  assign n31 = pi0 & ~pi2;
  assign n32 = pi6 & ~pi7;
  assign n33 = ~pi0 & pi2;
  assign n34 = n32 & n33;
  assign n35 = ~n31 & ~n34;
  assign n36 = n24 & ~n35;
  assign n37 = pi6 & pi9;
  assign n38 = ~pi7 & ~pi9;
  assign n39 = ~pi6 & n38;
  assign n40 = ~n37 & ~n39;
  assign n41 = ~pi5 & ~pi6;
  assign n42 = n40 & ~n41;
  assign n43 = ~pi9 & ~n42;
  assign n44 = ~pi0 & n43;
  assign n45 = ~n36 & ~n44;
  assign n46 = ~pi4 & ~n45;
  assign n47 = ~pi0 & ~pi2;
  assign n48 = pi4 & ~pi5;
  assign n49 = ~n40 & n48;
  assign n50 = ~n47 & n49;
  assign n51 = pi4 & pi5;
  assign n52 = n32 & n51;
  assign n53 = n24 & ~n32;
  assign n54 = ~pi4 & n53;
  assign n55 = pi4 & ~pi9;
  assign n56 = pi7 & n19;
  assign n57 = n55 & n56;
  assign n58 = ~n54 & ~n57;
  assign n59 = ~n52 & n58;
  assign n60 = ~pi2 & ~n59;
  assign n61 = ~n50 & ~n60;
  assign n62 = ~n46 & n61;
  assign n63 = ~n30 & n62;
  assign n64 = ~pi6 & n63;
  assign n65 = ~n17 & ~n64;
  assign n66 = pi4 & ~n65;
  assign n67 = ~pi7 & n66;
  assign n68 = pi6 & ~n63;
  assign n69 = pi4 & ~pi6;
  assign n70 = n33 & n69;
  assign n71 = ~n68 & ~n70;
  assign n72 = pi0 & ~pi4;
  assign n73 = ~pi4 & pi6;
  assign n74 = ~n72 & ~n73;
  assign n75 = ~n31 & n74;
  assign n76 = n71 & n75;
  assign n77 = pi7 & ~n76;
  assign n78 = ~n64 & ~n68;
  assign n79 = ~pi4 & n78;
  assign n80 = ~n77 & ~n79;
  assign n81 = ~n67 & n80;
  assign n82 = ~pi5 & ~n81;
  assign n83 = pi0 & pi6;
  assign n84 = pi5 & n18;
  assign n85 = ~n83 & ~n84;
  assign n86 = pi7 & ~n85;
  assign n87 = ~pi6 & ~n63;
  assign n88 = ~pi4 & n87;
  assign n89 = ~pi4 & pi7;
  assign n90 = pi5 & n89;
  assign n91 = ~n88 & ~n90;
  assign n92 = pi2 & ~n91;
  assign n93 = n32 & n47;
  assign n94 = ~pi4 & n93;
  assign n95 = n18 & n73;
  assign n96 = pi0 & ~n63;
  assign n97 = pi6 & n96;
  assign n98 = pi4 & n97;
  assign n99 = ~n95 & ~n98;
  assign n100 = ~n94 & n99;
  assign n101 = pi5 & ~n100;
  assign n102 = ~n92 & ~n101;
  assign n103 = ~n86 & n102;
  assign n104 = ~n82 & n103;
  assign n105 = ~pi9 & ~n104;
  assign n106 = n63 & n83;
  assign n107 = pi7 & n106;
  assign n108 = pi0 & ~pi7;
  assign n109 = ~pi6 & n108;
  assign n110 = ~n107 & ~n109;
  assign n111 = ~n51 & ~n110;
  assign n112 = pi6 & n51;
  assign n113 = ~pi0 & pi7;
  assign n114 = n24 & n89;
  assign n115 = ~pi0 & n63;
  assign n116 = n114 & ~n115;
  assign n117 = pi9 & n32;
  assign n118 = n51 & n96;
  assign n119 = n18 & n48;
  assign n120 = ~pi4 & ~pi5;
  assign n121 = n63 & n120;
  assign n122 = ~n119 & ~n121;
  assign n123 = ~n118 & n122;
  assign n124 = n117 & ~n123;
  assign n125 = ~n116 & ~n124;
  assign n126 = ~pi7 & n125;
  assign n127 = ~n113 & ~n126;
  assign n128 = n112 & ~n127;
  assign n129 = n48 & n117;
  assign n130 = n125 & n129;
  assign n131 = n64 & n116;
  assign n132 = ~n130 & ~n131;
  assign n133 = n23 & n132;
  assign n134 = n22 & n133;
  assign n135 = ~pi6 & ~n120;
  assign n136 = ~pi0 & ~n135;
  assign n137 = n21 & n136;
  assign n138 = ~n134 & ~n137;
  assign n139 = ~n125 & ~n138;
  assign n140 = ~n63 & n136;
  assign n141 = n51 & n64;
  assign n142 = ~n140 & ~n141;
  assign n143 = pi7 & ~n142;
  assign n144 = pi4 & ~n132;
  assign n145 = n20 & n144;
  assign n146 = n41 & n72;
  assign n147 = ~n145 & ~n146;
  assign n148 = n63 & ~n147;
  assign n149 = ~n18 & ~n47;
  assign n150 = n69 & n149;
  assign n151 = n72 & n126;
  assign n152 = ~n150 & ~n151;
  assign n153 = ~pi5 & ~n152;
  assign n154 = n23 & n78;
  assign n155 = n48 & n68;
  assign n156 = ~n130 & n155;
  assign n157 = ~n154 & ~n156;
  assign n158 = ~pi7 & ~n157;
  assign n159 = ~n153 & ~n158;
  assign n160 = ~n148 & n159;
  assign n161 = ~n143 & n160;
  assign n162 = ~n139 & n161;
  assign n163 = ~n128 & n162;
  assign n164 = ~n111 & n163;
  assign n165 = pi9 & ~n164;
  assign n166 = pi8 & n165;
  assign n167 = ~pi8 & ~n165;
  assign n168 = ~pi6 & n51;
  assign n169 = ~pi7 & n168;
  assign n170 = ~n167 & ~n169;
  assign n171 = ~n166 & n170;
  assign n172 = pi9 & ~n171;
  assign po0 = n105 | n172;
  assign n174 = ~pi5 & n69;
  assign n175 = n18 & n174;
  assign po3 = pi1 & pi3;
  assign n177 = ~pi1 & ~pi3;
  assign n178 = pi7 & n177;
  assign n179 = ~po3 & ~n178;
  assign n180 = n175 & ~n179;
  assign n181 = n20 & po3;
  assign n182 = ~n55 & n181;
  assign n183 = ~pi6 & po3;
  assign n184 = n27 & n183;
  assign n185 = ~pi5 & n83;
  assign n186 = n25 & n185;
  assign n187 = ~n184 & ~n186;
  assign n188 = pi7 & ~n187;
  assign n189 = n33 & po3;
  assign n190 = ~pi1 & pi3;
  assign n191 = pi5 & n190;
  assign n192 = ~n33 & n191;
  assign n193 = ~n189 & ~n192;
  assign n194 = n32 & ~n193;
  assign n195 = n33 & n177;
  assign n196 = pi1 & ~pi3;
  assign n197 = ~n33 & n196;
  assign n198 = ~n195 & ~n197;
  assign n199 = pi5 & ~n198;
  assign n200 = ~n194 & ~n199;
  assign n201 = pi9 & ~n200;
  assign n202 = ~pi1 & n43;
  assign n203 = ~n201 & ~n202;
  assign n204 = ~pi4 & ~n203;
  assign n205 = ~pi3 & ~n59;
  assign n206 = n49 & ~n177;
  assign n207 = ~n205 & ~n206;
  assign n208 = ~n204 & n207;
  assign n209 = ~n188 & n208;
  assign n210 = ~n182 & n209;
  assign n211 = n96 & ~n210;
  assign n212 = ~n96 & n210;
  assign n213 = ~n211 & ~n212;
  assign n214 = ~n51 & ~n135;
  assign n215 = pi1 & ~n32;
  assign n216 = n214 & n215;
  assign n217 = ~n213 & n216;
  assign po2 = po3 | n177;
  assign n219 = ~n18 & ~po2;
  assign n220 = pi3 & ~pi7;
  assign n221 = ~n219 & ~n220;
  assign n222 = n174 & ~n221;
  assign n223 = n23 & ~n210;
  assign n224 = pi1 & ~n51;
  assign n225 = ~n223 & ~n224;
  assign n226 = ~pi6 & ~n225;
  assign n227 = n63 & n210;
  assign n228 = pi6 & n227;
  assign n229 = ~n63 & ~n210;
  assign n230 = ~n228 & ~n229;
  assign n231 = n23 & ~n230;
  assign n232 = n114 & n183;
  assign n233 = ~pi1 & n210;
  assign n234 = n114 & ~n233;
  assign n235 = pi1 & ~n210;
  assign n236 = n51 & n235;
  assign n237 = n120 & n210;
  assign n238 = n48 & po3;
  assign n239 = ~n237 & ~n238;
  assign n240 = ~n236 & n239;
  assign n241 = n117 & ~n240;
  assign n242 = ~n234 & ~n241;
  assign n243 = n129 & n242;
  assign n244 = ~n232 & ~n243;
  assign n245 = ~n63 & ~n132;
  assign n246 = n244 & ~n245;
  assign n247 = n125 & n242;
  assign n248 = ~n63 & n247;
  assign n249 = ~n246 & ~n248;
  assign n250 = ~n210 & ~n249;
  assign n251 = n210 & n249;
  assign n252 = ~n250 & ~n251;
  assign n253 = n48 & ~n252;
  assign n254 = pi0 & ~n125;
  assign n255 = ~n242 & ~n254;
  assign n256 = n242 & n254;
  assign n257 = ~n255 & ~n256;
  assign n258 = ~pi1 & n120;
  assign n259 = ~n257 & n258;
  assign n260 = n51 & n247;
  assign n261 = ~n125 & ~n242;
  assign n262 = n51 & n261;
  assign n263 = ~n260 & ~n262;
  assign n264 = ~n259 & n263;
  assign n265 = ~n253 & n264;
  assign n266 = pi6 & ~n265;
  assign n267 = pi1 & ~pi4;
  assign n268 = ~pi5 & n257;
  assign n269 = n267 & n268;
  assign n270 = ~n266 & ~n269;
  assign n271 = ~n231 & n270;
  assign n272 = ~n226 & n271;
  assign n273 = ~pi7 & ~n272;
  assign n274 = n213 & n214;
  assign n275 = n51 & n136;
  assign n276 = ~n274 & ~n275;
  assign n277 = ~pi1 & ~n276;
  assign n278 = n131 & ~n244;
  assign n279 = ~n131 & n244;
  assign n280 = ~n278 & ~n279;
  assign n281 = ~n242 & ~n280;
  assign n282 = n242 & n280;
  assign n283 = ~n281 & ~n282;
  assign n284 = n23 & ~n283;
  assign n285 = n51 & n227;
  assign n286 = ~n284 & ~n285;
  assign n287 = ~pi6 & ~n286;
  assign n288 = n87 & ~n210;
  assign n289 = pi1 & n83;
  assign n290 = ~n288 & ~n289;
  assign n291 = n51 & ~n290;
  assign n292 = ~n287 & ~n291;
  assign n293 = ~n277 & n292;
  assign n294 = pi7 & ~n293;
  assign n295 = ~n273 & ~n294;
  assign n296 = ~n222 & n295;
  assign n297 = ~n217 & n296;
  assign n298 = ~n180 & n297;
  assign n299 = pi9 & ~n298;
  assign n300 = ~pi8 & n165;
  assign n301 = n299 & ~n300;
  assign n302 = ~n299 & n300;
  assign n303 = ~n169 & ~n302;
  assign n304 = ~n301 & n303;
  assign n305 = pi9 & ~n304;
  assign n306 = ~pi3 & pi6;
  assign n307 = ~pi6 & n210;
  assign n308 = ~n306 & ~n307;
  assign n309 = pi4 & ~n308;
  assign n310 = ~pi7 & n309;
  assign n311 = ~pi7 & ~n210;
  assign n312 = n73 & ~n311;
  assign n313 = ~pi4 & ~pi6;
  assign n314 = ~n210 & n313;
  assign n315 = pi6 & ~n210;
  assign n316 = ~n196 & ~n315;
  assign n317 = n69 & n190;
  assign n318 = ~n267 & ~n317;
  assign n319 = n316 & n318;
  assign n320 = pi7 & ~n319;
  assign n321 = ~n314 & ~n320;
  assign n322 = ~n312 & n321;
  assign n323 = ~n310 & n322;
  assign n324 = ~pi5 & ~n323;
  assign n325 = pi1 & pi6;
  assign n326 = pi5 & po3;
  assign n327 = ~n325 & ~n326;
  assign n328 = pi7 & ~n327;
  assign n329 = ~n90 & ~n314;
  assign n330 = pi3 & ~n329;
  assign n331 = pi4 & n235;
  assign n332 = pi6 & n331;
  assign n333 = n32 & n177;
  assign n334 = ~pi4 & n333;
  assign n335 = n73 & po3;
  assign n336 = ~n334 & ~n335;
  assign n337 = ~n332 & n336;
  assign n338 = pi5 & ~n337;
  assign n339 = ~n330 & ~n338;
  assign n340 = ~n328 & n339;
  assign n341 = ~n324 & n340;
  assign n342 = ~pi9 & ~n341;
  assign po1 = n305 | n342;
  assign n344 = n23 & n32;
  assign n345 = ~n168 & ~n344;
  assign n346 = n227 & ~n345;
  assign n347 = ~pi1 & ~n254;
  assign n348 = ~pi4 & ~n347;
  assign n349 = ~n242 & n348;
  assign n350 = ~n246 & ~n251;
  assign n351 = pi4 & n350;
  assign n352 = n254 & n267;
  assign n353 = ~n351 & ~n352;
  assign n354 = ~n349 & n353;
  assign n355 = n19 & ~n354;
  assign n356 = ~n168 & ~n260;
  assign n357 = ~n355 & n356;
  assign n358 = ~pi7 & ~n357;
  assign n359 = ~n279 & ~n282;
  assign n360 = n23 & n359;
  assign n361 = n96 & ~n233;
  assign n362 = ~n235 & ~n361;
  assign n363 = n214 & ~n362;
  assign n364 = n175 & ~n177;
  assign n365 = ~n238 & ~n275;
  assign n366 = ~n325 & ~n365;
  assign n367 = ~n364 & ~n366;
  assign n368 = ~n363 & n367;
  assign n369 = ~n360 & n368;
  assign n370 = pi7 & ~n369;
  assign n371 = n299 & n300;
  assign n372 = ~n370 & ~n371;
  assign n373 = ~n358 & n372;
  assign n374 = ~n346 & n373;
  assign po4 = pi9 & ~n374;
  assign po5 = ~n149 & po2;
endmodule
