module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n415, n416, n417, n418,
    n419, n420, n422, n423, n424, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504,
    n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639,
    n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n677, n678, n679, n680, n681, n682;
  assign n22 = ~pi5  & pi7 ;
  assign n23 = pi8  & n22;
  assign n24 = ~pi7  & pi9 ;
  assign n25 = ~n23 & ~n24;
  assign n26 = pi1  & ~n25;
  assign n27 = pi1  & ~pi7 ;
  assign n28 = ~pi5  & ~pi9 ;
  assign n29 = ~n27 & n28;
  assign n30 = ~n26 & ~n29;
  assign n31 = pi0  & ~pi2 ;
  assign n32 = ~n30 & n31;
  assign n33 = ~pi0  & ~pi1 ;
  assign n34 = pi2  & ~pi9 ;
  assign n35 = n33 & n34;
  assign n36 = n23 & n35;
  assign n37 = ~n32 & ~n36;
  assign n38 = ~pi3  & ~n37;
  assign n39 = ~pi3  & ~pi5 ;
  assign n40 = ~pi0  & pi9 ;
  assign n41 = pi1  & ~n40;
  assign n42 = ~pi1  & pi9 ;
  assign n43 = n39 & ~n42;
  assign n44 = ~n41 & n43;
  assign n45 = pi0  & ~pi9 ;
  assign n46 = ~pi1  & ~n45;
  assign n47 = pi1  & ~pi9 ;
  assign n48 = ~pi7  & ~n47;
  assign n49 = ~n46 & n48;
  assign n50 = ~n44 & ~n49;
  assign n51 = ~pi2  & ~n50;
  assign n52 = ~pi2  & ~pi3 ;
  assign n53 = pi9  & ~n52;
  assign n54 = pi0  & pi3 ;
  assign n55 = ~n53 & ~n54;
  assign n56 = ~pi1  & ~n55;
  assign n57 = pi1  & ~pi3 ;
  assign n58 = pi1  & pi2 ;
  assign n59 = ~pi2  & ~pi5 ;
  assign n60 = ~pi0  & ~n59;
  assign n61 = ~n58 & ~n60;
  assign n62 = ~pi9  & ~n61;
  assign n63 = ~n56 & ~n57;
  assign n64 = ~n62 & n63;
  assign n65 = ~pi7  & ~n64;
  assign n66 = ~n51 & ~n65;
  assign n67 = ~pi8  & ~n66;
  assign n68 = ~n38 & ~n67;
  assign n69 = ~pi6  & ~n68;
  assign n70 = ~pi1  & ~pi9 ;
  assign n71 = ~pi8  & n70;
  assign n72 = ~pi0  & n52;
  assign n73 = n71 & n72;
  assign n74 = ~pi0  & ~pi2 ;
  assign n75 = n42 & n74;
  assign n76 = ~pi5  & ~n75;
  assign n77 = pi6  & ~n76;
  assign n78 = ~n40 & ~n45;
  assign n79 = pi1  & pi5 ;
  assign n80 = pi2  & n79;
  assign n81 = n78 & n80;
  assign n82 = ~n77 & ~n81;
  assign n83 = pi8  & ~n82;
  assign n84 = ~pi1  & ~n40;
  assign n85 = ~pi8  & ~n84;
  assign n86 = ~pi1  & pi2 ;
  assign n87 = n45 & n86;
  assign n88 = ~n85 & ~n87;
  assign n89 = ~pi5  & ~n88;
  assign n90 = ~n83 & ~n89;
  assign n91 = pi3  & ~n90;
  assign n92 = pi1  & ~pi8 ;
  assign n93 = pi2  & ~pi3 ;
  assign n94 = n42 & n93;
  assign n95 = ~n92 & ~n94;
  assign n96 = ~pi0  & ~n95;
  assign n97 = pi2  & pi9 ;
  assign n98 = ~pi2  & pi6 ;
  assign n99 = pi3  & ~n98;
  assign n100 = n70 & ~n99;
  assign n101 = ~n97 & ~n100;
  assign n102 = ~pi8  & ~n101;
  assign n103 = ~n96 & ~n102;
  assign n104 = ~pi5  & ~n103;
  assign n105 = ~pi2  & ~n45;
  assign n106 = ~pi6  & ~n105;
  assign n107 = ~pi3  & n41;
  assign n108 = n105 & ~n107;
  assign n109 = pi5  & ~n106;
  assign n110 = ~n108 & n109;
  assign n111 = ~pi2  & n47;
  assign n112 = ~n97 & ~n111;
  assign n113 = ~pi0  & ~pi3 ;
  assign n114 = pi6  & n113;
  assign n115 = ~n112 & n114;
  assign n116 = ~n110 & ~n115;
  assign n117 = pi8  & ~n116;
  assign n118 = ~n73 & ~n104;
  assign n119 = ~n117 & n118;
  assign n120 = ~n91 & n119;
  assign n121 = ~pi7  & ~n120;
  assign n122 = ~n69 & ~n121;
  assign n123 = ~pi4  & ~n122;
  assign n124 = ~pi1  & ~pi3 ;
  assign n125 = ~pi6  & pi8 ;
  assign n126 = pi5  & ~n125;
  assign n127 = pi4  & pi8 ;
  assign n128 = ~pi6  & ~pi9 ;
  assign n129 = ~n127 & ~n128;
  assign n130 = n126 & ~n129;
  assign n131 = pi6  & ~pi9 ;
  assign n132 = pi4  & pi9 ;
  assign n133 = ~n131 & ~n132;
  assign n134 = pi5  & pi6 ;
  assign n135 = ~pi8  & ~n134;
  assign n136 = ~n133 & n135;
  assign n137 = ~n130 & ~n136;
  assign n138 = ~pi7  & n74;
  assign n139 = n124 & n138;
  assign n140 = ~n137 & n139;
  assign po0  = n123 | n140;
  assign n142 = n34 & n125;
  assign n143 = ~pi2  & ~pi8 ;
  assign n144 = ~pi0  & ~pi9 ;
  assign n145 = n143 & n144;
  assign n146 = pi0  & pi8 ;
  assign n147 = pi9  & n146;
  assign n148 = pi2  & n147;
  assign n149 = ~n145 & ~n148;
  assign n150 = pi5  & ~n149;
  assign n151 = ~pi8  & n28;
  assign n152 = ~pi5  & pi8 ;
  assign n153 = pi6  & pi9 ;
  assign n154 = ~n152 & ~n153;
  assign n155 = ~pi0  & ~n154;
  assign n156 = pi6  & pi8 ;
  assign n157 = pi9  & n156;
  assign n158 = ~n151 & ~n157;
  assign n159 = ~n155 & n158;
  assign n160 = pi2  & ~n159;
  assign n161 = ~n150 & ~n160;
  assign n162 = ~pi1  & ~n161;
  assign n163 = ~pi0  & pi5 ;
  assign n164 = ~pi8  & pi9 ;
  assign n165 = n163 & n164;
  assign n166 = pi0  & ~n156;
  assign n167 = ~n154 & n166;
  assign n168 = ~n165 & ~n167;
  assign n169 = ~pi2  & ~n168;
  assign n170 = ~pi6  & ~pi8 ;
  assign n171 = ~pi0  & pi6 ;
  assign n172 = ~pi2  & ~n171;
  assign n173 = n152 & ~n172;
  assign n174 = ~n170 & ~n173;
  assign n175 = ~pi9  & ~n174;
  assign n176 = ~n169 & ~n175;
  assign n177 = pi1  & ~n176;
  assign n178 = ~n142 & ~n162;
  assign n179 = ~n177 & n178;
  assign n180 = ~pi4  & ~n179;
  assign n181 = ~pi2  & n33;
  assign n182 = pi5  & ~pi8 ;
  assign n183 = ~n127 & ~n182;
  assign n184 = n128 & ~n183;
  assign n185 = pi4  & n153;
  assign n186 = ~n184 & ~n185;
  assign n187 = n181 & ~n186;
  assign n188 = ~n180 & ~n187;
  assign n189 = ~pi3  & ~n188;
  assign n190 = pi3  & pi8 ;
  assign n191 = ~pi2  & ~n190;
  assign n192 = ~pi0  & ~n191;
  assign n193 = pi5  & n143;
  assign n194 = ~pi3  & ~pi8 ;
  assign n195 = ~n152 & ~n194;
  assign n196 = pi0  & n195;
  assign n197 = ~n193 & ~n196;
  assign n198 = ~pi1  & ~n197;
  assign n199 = ~pi2  & pi8 ;
  assign n200 = pi0  & n199;
  assign n201 = pi0  & ~pi5 ;
  assign n202 = ~n163 & ~n201;
  assign n203 = ~n200 & n202;
  assign n204 = pi1  & ~n203;
  assign n205 = ~n192 & ~n204;
  assign n206 = ~n198 & n205;
  assign n207 = ~pi6  & ~n206;
  assign n208 = ~pi1  & ~pi8 ;
  assign n209 = ~pi2  & ~n208;
  assign n210 = ~pi1  & pi8 ;
  assign n211 = pi6  & n210;
  assign n212 = ~n209 & ~n211;
  assign n213 = pi3  & ~n212;
  assign n214 = ~pi0  & pi8 ;
  assign n215 = pi0  & pi1 ;
  assign n216 = ~pi1  & ~pi6 ;
  assign n217 = ~pi2  & ~n214;
  assign n218 = ~n215 & ~n216;
  assign n219 = n217 & n218;
  assign n220 = ~n213 & ~n219;
  assign n221 = ~pi5  & ~n220;
  assign n222 = ~pi9  & ~n221;
  assign n223 = ~n207 & n222;
  assign n224 = ~pi1  & ~pi2 ;
  assign n225 = pi3  & ~pi8 ;
  assign n226 = n224 & n225;
  assign n227 = ~n79 & ~n226;
  assign n228 = pi0  & ~n227;
  assign n229 = pi3  & n58;
  assign n230 = ~pi5  & ~n229;
  assign n231 = ~n52 & ~n230;
  assign n232 = ~n228 & ~n231;
  assign n233 = pi6  & ~n232;
  assign n234 = n182 & n229;
  assign n235 = pi9  & ~n234;
  assign n236 = ~n233 & n235;
  assign n237 = ~pi4  & ~n236;
  assign n238 = ~n223 & n237;
  assign n239 = ~n189 & ~n238;
  assign n240 = ~pi7  & ~n239;
  assign n241 = ~pi6  & n39;
  assign n242 = n47 & n199;
  assign n243 = n105 & ~n215;
  assign n244 = pi2  & ~n33;
  assign n245 = ~pi8  & ~n244;
  assign n246 = ~n243 & n245;
  assign n247 = ~n242 & ~n246;
  assign n248 = pi7  & ~n247;
  assign n249 = ~n35 & ~n248;
  assign n250 = ~pi4  & n241;
  assign n251 = ~n249 & n250;
  assign po1  = n240 | n251;
  assign n253 = ~pi8  & ~pi9 ;
  assign n254 = pi8  & pi9 ;
  assign n255 = ~n253 & ~n254;
  assign n256 = ~n70 & ~n255;
  assign n257 = pi2  & ~n256;
  assign n258 = ~pi5  & ~n97;
  assign n259 = pi5  & ~n253;
  assign n260 = ~n147 & n259;
  assign n261 = pi1  & ~n258;
  assign n262 = ~n260 & n261;
  assign n263 = ~n257 & ~n262;
  assign n264 = ~pi3  & ~n263;
  assign n265 = n53 & n210;
  assign n266 = ~pi1  & pi3 ;
  assign n267 = pi5  & ~n266;
  assign n268 = ~pi2  & n253;
  assign n269 = ~n267 & n268;
  assign n270 = ~n265 & ~n269;
  assign n271 = pi0  & ~n270;
  assign n272 = ~n264 & ~n271;
  assign n273 = ~pi6  & ~n272;
  assign n274 = pi6  & ~n42;
  assign n275 = ~n47 & ~n274;
  assign n276 = pi8  & ~n275;
  assign n277 = pi1  & pi9 ;
  assign n278 = ~n70 & ~n277;
  assign n279 = n194 & ~n278;
  assign n280 = ~n276 & ~n279;
  assign n281 = ~pi2  & ~n280;
  assign n282 = pi8  & ~n34;
  assign n283 = pi2  & n277;
  assign n284 = ~n210 & ~n283;
  assign n285 = pi6  & ~n284;
  assign n286 = pi2  & n253;
  assign n287 = ~n282 & ~n286;
  assign n288 = ~n285 & n287;
  assign n289 = pi3  & ~n288;
  assign n290 = ~n281 & ~n289;
  assign n291 = n201 & ~n290;
  assign n292 = ~n273 & ~n291;
  assign n293 = ~pi4  & ~n292;
  assign n294 = pi3  & ~n199;
  assign n295 = pi5  & ~n294;
  assign n296 = pi2  & ~pi5 ;
  assign n297 = pi3  & ~n296;
  assign n298 = pi8  & ~n297;
  assign n299 = ~n295 & ~n298;
  assign n300 = pi1  & ~n299;
  assign n301 = ~pi5  & pi6 ;
  assign n302 = ~pi3  & n301;
  assign n303 = n208 & n302;
  assign n304 = ~n300 & ~n303;
  assign n305 = ~pi9  & ~n304;
  assign n306 = pi1  & pi8 ;
  assign n307 = pi6  & ~n306;
  assign n308 = ~pi9  & ~n307;
  assign n309 = ~pi2  & ~n308;
  assign n310 = ~pi8  & n42;
  assign n311 = ~n309 & ~n310;
  assign n312 = pi3  & ~n311;
  assign n313 = pi6  & ~pi8 ;
  assign n314 = ~pi3  & pi9 ;
  assign n315 = pi1  & n314;
  assign n316 = n313 & n315;
  assign n317 = pi3  & ~pi9 ;
  assign n318 = ~n47 & ~n225;
  assign n319 = ~pi6  & ~n317;
  assign n320 = ~n318 & n319;
  assign n321 = pi2  & ~n125;
  assign n322 = pi1  & ~n321;
  assign n323 = pi5  & ~n191;
  assign n324 = ~n322 & n323;
  assign n325 = ~n316 & ~n320;
  assign n326 = ~n324 & n325;
  assign n327 = ~n312 & n326;
  assign n328 = ~n305 & n327;
  assign n329 = ~pi4  & ~n328;
  assign n330 = ~pi3  & pi4 ;
  assign n331 = ~n254 & ~n313;
  assign n332 = ~pi5  & ~n331;
  assign n333 = n224 & n330;
  assign n334 = ~n332 & n333;
  assign n335 = ~n329 & ~n334;
  assign n336 = ~pi0  & ~n335;
  assign n337 = ~n293 & ~n336;
  assign n338 = ~pi7  & ~n337;
  assign n339 = pi7  & n254;
  assign n340 = pi0  & ~n339;
  assign n341 = n41 & ~n340;
  assign n342 = n45 & n208;
  assign n343 = ~n341 & ~n342;
  assign n344 = ~pi5  & ~pi6 ;
  assign n345 = ~pi4  & n52;
  assign n346 = n344 & n345;
  assign n347 = ~n343 & n346;
  assign po2  = n338 | n347;
  assign n349 = pi2  & n301;
  assign n350 = pi5  & pi9 ;
  assign n351 = pi8  & n350;
  assign n352 = ~pi6  & n351;
  assign n353 = ~n151 & ~n352;
  assign n354 = pi2  & ~n353;
  assign n355 = ~pi3  & ~n313;
  assign n356 = ~n126 & ~n355;
  assign n357 = ~n354 & ~n356;
  assign n358 = pi1  & ~n357;
  assign n359 = pi6  & ~n52;
  assign n360 = ~n317 & ~n359;
  assign n361 = ~pi1  & ~n360;
  assign n362 = ~n349 & ~n361;
  assign n363 = ~n358 & n362;
  assign n364 = ~pi4  & ~n363;
  assign n365 = ~pi5  & ~n254;
  assign n366 = ~n134 & ~n344;
  assign n367 = n333 & ~n365;
  assign n368 = ~n366 & n367;
  assign n369 = ~n364 & ~n368;
  assign n370 = ~pi0  & ~n369;
  assign n371 = ~pi9  & n301;
  assign n372 = n306 & n371;
  assign n373 = pi2  & ~n195;
  assign n374 = ~pi2  & pi5 ;
  assign n375 = pi8  & n374;
  assign n376 = ~n373 & ~n375;
  assign n377 = ~pi9  & ~n376;
  assign n378 = pi5  & n164;
  assign n379 = ~pi3  & ~n378;
  assign n380 = ~pi2  & ~n379;
  assign n381 = ~pi6  & ~n225;
  assign n382 = pi3  & ~pi5 ;
  assign n383 = ~n381 & ~n382;
  assign n384 = ~n380 & ~n383;
  assign n385 = ~n377 & n384;
  assign n386 = pi1  & ~n385;
  assign n387 = n193 & n216;
  assign n388 = ~n302 & ~n387;
  assign n389 = ~pi9  & ~n388;
  assign n390 = ~n386 & ~n389;
  assign n391 = pi0  & ~n390;
  assign n392 = ~n28 & ~n170;
  assign n393 = ~pi2  & ~n392;
  assign n394 = ~pi6  & ~n350;
  assign n395 = pi5  & pi8 ;
  assign n396 = ~n277 & ~n395;
  assign n397 = n394 & ~n396;
  assign n398 = ~n393 & ~n397;
  assign n399 = pi3  & ~n398;
  assign n400 = pi3  & ~pi6 ;
  assign n401 = pi2  & n400;
  assign n402 = ~n52 & n301;
  assign n403 = ~n401 & ~n402;
  assign n404 = pi9  & ~n403;
  assign n405 = ~n371 & ~n400;
  assign n406 = ~pi8  & ~n405;
  assign n407 = ~n404 & ~n406;
  assign n408 = ~pi1  & ~n407;
  assign n409 = ~n372 & ~n399;
  assign n410 = ~n408 & n409;
  assign n411 = ~n391 & n410;
  assign n412 = ~pi4  & ~n411;
  assign n413 = ~n370 & ~n412;
  assign po3  = ~pi7  & ~n413;
  assign n415 = ~pi4  & n244;
  assign n416 = pi3  & ~pi4 ;
  assign n417 = ~n330 & ~n416;
  assign n418 = n181 & ~n417;
  assign n419 = ~n415 & ~n418;
  assign n420 = ~pi7  & n134;
  assign po4  = ~n419 & n420;
  assign n422 = ~n181 & n416;
  assign n423 = n181 & n330;
  assign n424 = ~n422 & ~n423;
  assign po5  = n420 & ~n424;
  assign n426 = pi4  & n33;
  assign n427 = n52 & n426;
  assign n428 = ~n134 & ~n427;
  assign n429 = ~pi7  & ~n428;
  assign n430 = pi7  & ~pi9 ;
  assign n431 = pi8  & ~n430;
  assign n432 = n86 & ~n431;
  assign n433 = ~n111 & ~n432;
  assign n434 = ~pi0  & ~n433;
  assign n435 = pi1  & n147;
  assign n436 = ~n253 & ~n435;
  assign n437 = ~pi2  & pi7 ;
  assign n438 = ~n436 & n437;
  assign n439 = ~n434 & ~n438;
  assign n440 = n344 & ~n439;
  assign n441 = pi2  & pi8 ;
  assign n442 = ~n143 & ~n441;
  assign n443 = pi6  & ~n255;
  assign n444 = ~n442 & n443;
  assign n445 = ~pi1  & ~pi5 ;
  assign n446 = pi2  & ~n445;
  assign n447 = n128 & ~n446;
  assign n448 = pi5  & n277;
  assign n449 = ~n447 & ~n448;
  assign n450 = pi0  & ~n449;
  assign n451 = ~pi0  & pi2 ;
  assign n452 = ~n28 & n451;
  assign n453 = ~n450 & ~n452;
  assign n454 = pi8  & ~n453;
  assign n455 = pi9  & n451;
  assign n456 = ~n71 & ~n455;
  assign n457 = pi5  & ~n456;
  assign n458 = ~n444 & ~n457;
  assign n459 = ~n454 & n458;
  assign n460 = ~pi7  & ~n459;
  assign n461 = ~n440 & ~n460;
  assign n462 = ~pi3  & ~n461;
  assign n463 = n40 & n441;
  assign n464 = ~pi2  & ~pi9 ;
  assign n465 = ~pi0  & ~n313;
  assign n466 = ~n395 & n464;
  assign n467 = ~n465 & n466;
  assign n468 = ~n463 & ~n467;
  assign n469 = ~pi1  & ~n468;
  assign n470 = n78 & n374;
  assign n471 = ~pi6  & ~n296;
  assign n472 = n40 & ~n471;
  assign n473 = ~n470 & ~n472;
  assign n474 = ~pi8  & ~n473;
  assign n475 = pi2  & ~n253;
  assign n476 = ~n147 & ~n475;
  assign n477 = pi6  & ~n476;
  assign n478 = ~n474 & ~n477;
  assign n479 = pi1  & ~n478;
  assign n480 = n92 & ~n451;
  assign n481 = pi0  & n156;
  assign n482 = ~pi2  & n481;
  assign n483 = ~n480 & ~n482;
  assign n484 = pi9  & ~n483;
  assign n485 = ~pi0  & ~pi6 ;
  assign n486 = ~n208 & n485;
  assign n487 = ~n58 & ~n486;
  assign n488 = n278 & ~n487;
  assign n489 = ~pi1  & ~n253;
  assign n490 = pi0  & ~n489;
  assign n491 = ~n47 & n490;
  assign n492 = ~n488 & ~n491;
  assign n493 = ~pi5  & ~n492;
  assign n494 = ~pi0  & ~pi8 ;
  assign n495 = n47 & ~n201;
  assign n496 = ~n494 & n495;
  assign n497 = ~n484 & ~n496;
  assign n498 = ~n493 & n497;
  assign n499 = pi3  & ~n498;
  assign n500 = ~n469 & ~n479;
  assign n501 = ~n499 & n500;
  assign n502 = ~pi7  & ~n501;
  assign n503 = ~n462 & ~n502;
  assign n504 = ~pi4  & ~n503;
  assign po6  = ~n429 & ~n504;
  assign n506 = n128 & n194;
  assign n507 = n214 & n400;
  assign n508 = ~n313 & ~n507;
  assign n509 = pi9  & ~n508;
  assign n510 = ~pi8  & ~n153;
  assign n511 = pi0  & ~n400;
  assign n512 = ~n131 & ~n511;
  assign n513 = ~n510 & ~n512;
  assign n514 = ~pi2  & ~n509;
  assign n515 = ~n513 & n514;
  assign n516 = ~pi3  & n254;
  assign n517 = pi3  & ~n254;
  assign n518 = ~n146 & ~n517;
  assign n519 = ~pi6  & ~n518;
  assign n520 = pi2  & ~n516;
  assign n521 = ~n519 & n520;
  assign n522 = ~n515 & ~n521;
  assign n523 = pi1  & ~n506;
  assign n524 = ~n522 & n523;
  assign n525 = n171 & ~n255;
  assign n526 = ~pi6  & ~n254;
  assign n527 = n105 & n526;
  assign n528 = ~n525 & ~n527;
  assign n529 = pi3  & ~n528;
  assign n530 = ~pi0  & n143;
  assign n531 = ~n481 & ~n530;
  assign n532 = ~pi9  & ~n531;
  assign n533 = ~pi6  & ~n194;
  assign n534 = n475 & ~n533;
  assign n535 = ~pi1  & ~n534;
  assign n536 = ~n532 & n535;
  assign n537 = ~n529 & n536;
  assign n538 = ~n524 & ~n537;
  assign n539 = pi3  & n143;
  assign n540 = n131 & n539;
  assign n541 = ~n538 & ~n540;
  assign n542 = ~pi5  & ~n541;
  assign n543 = pi2  & pi3 ;
  assign n544 = n351 & n543;
  assign n545 = pi3  & pi5 ;
  assign n546 = ~n34 & ~n545;
  assign n547 = ~pi0  & ~n546;
  assign n548 = pi3  & n374;
  assign n549 = ~n547 & ~n548;
  assign n550 = ~pi8  & ~n549;
  assign n551 = pi0  & ~n97;
  assign n552 = ~n464 & n551;
  assign n553 = ~pi9  & n163;
  assign n554 = ~n552 & ~n553;
  assign n555 = pi8  & ~n554;
  assign n556 = n97 & n182;
  assign n557 = ~n555 & ~n556;
  assign n558 = ~pi3  & ~n557;
  assign n559 = n464 & n545;
  assign n560 = pi1  & ~n559;
  assign n561 = ~n550 & n560;
  assign n562 = ~n558 & n561;
  assign n563 = n54 & n286;
  assign n564 = n255 & ~n543;
  assign n565 = ~pi2  & ~n54;
  assign n566 = pi5  & ~n565;
  assign n567 = ~n564 & n566;
  assign n568 = ~pi1  & ~n563;
  assign n569 = ~n567 & n568;
  assign n570 = ~n562 & ~n569;
  assign n571 = ~n544 & ~n570;
  assign n572 = ~pi6  & ~n571;
  assign n573 = ~n542 & ~n572;
  assign n574 = ~pi7  & ~n573;
  assign n575 = n255 & n451;
  assign n576 = pi8  & n31;
  assign n577 = n430 & n576;
  assign n578 = ~n575 & ~n577;
  assign n579 = n124 & n344;
  assign n580 = ~n578 & n579;
  assign n581 = ~n574 & ~n580;
  assign n582 = ~pi4  & ~n581;
  assign n583 = ~pi5  & ~pi7 ;
  assign n584 = n485 & n583;
  assign n585 = n333 & n584;
  assign po7  = ~n582 & ~n585;
  assign n587 = n124 & n201;
  assign n588 = ~n79 & ~n382;
  assign n589 = ~pi2  & ~n113;
  assign n590 = n588 & n589;
  assign n591 = ~n587 & ~n590;
  assign n592 = pi8  & ~n591;
  assign n593 = ~pi5  & ~n214;
  assign n594 = n58 & ~n545;
  assign n595 = ~n593 & n594;
  assign n596 = ~n592 & ~n595;
  assign n597 = ~pi9  & ~n596;
  assign n598 = ~n296 & ~n545;
  assign n599 = pi1  & ~n294;
  assign n600 = ~n598 & n599;
  assign n601 = ~n163 & n199;
  assign n602 = n266 & n601;
  assign n603 = ~n600 & ~n602;
  assign n604 = pi9  & ~n603;
  assign n605 = n70 & n374;
  assign n606 = ~n315 & ~n605;
  assign n607 = ~pi0  & ~n606;
  assign n608 = n278 & ~n445;
  assign n609 = n93 & ~n608;
  assign n610 = ~pi2  & ~n70;
  assign n611 = ~n314 & n610;
  assign n612 = n588 & n611;
  assign n613 = ~n607 & ~n609;
  assign n614 = ~n612 & n613;
  assign n615 = ~pi8  & ~n614;
  assign n616 = ~n597 & ~n604;
  assign n617 = ~n615 & n616;
  assign n618 = ~pi6  & ~n617;
  assign n619 = ~n47 & n214;
  assign n620 = n274 & ~n619;
  assign n621 = ~pi2  & ~n620;
  assign n622 = ~pi6  & ~n92;
  assign n623 = ~n490 & n622;
  assign n624 = n382 & ~n621;
  assign n625 = ~n623 & n624;
  assign n626 = ~n618 & ~n625;
  assign n627 = ~pi7  & ~n626;
  assign n628 = ~pi0  & ~n442;
  assign n629 = ~n200 & ~n628;
  assign n630 = ~pi9  & ~n629;
  assign n631 = ~pi8  & n455;
  assign n632 = ~n630 & ~n631;
  assign n633 = ~pi1  & ~n632;
  assign n634 = n277 & n530;
  assign n635 = ~n633 & ~n634;
  assign n636 = n241 & ~n635;
  assign n637 = ~n627 & ~n636;
  assign n638 = ~pi4  & ~n637;
  assign n639 = n423 & n583;
  assign po8  = ~n638 & ~n639;
  assign n641 = ~pi2  & n124;
  assign n642 = pi4  & ~n641;
  assign n643 = n365 & n401;
  assign n644 = ~pi6  & ~n351;
  assign n645 = ~pi3  & ~n644;
  assign n646 = ~pi3  & ~n28;
  assign n647 = pi3  & ~n153;
  assign n648 = n214 & ~n647;
  assign n649 = ~n646 & ~n648;
  assign n650 = ~pi2  & ~n649;
  assign n651 = ~n643 & ~n645;
  assign n652 = ~n650 & n651;
  assign n653 = pi1  & ~n652;
  assign n654 = n330 & ~n344;
  assign n655 = n214 & ~n394;
  assign n656 = n647 & ~n655;
  assign n657 = ~pi2  & ~n654;
  assign n658 = ~n656 & n657;
  assign n659 = n93 & ~n253;
  assign n660 = ~n365 & n659;
  assign n661 = ~n658 & ~n660;
  assign n662 = ~pi1  & ~n661;
  assign n663 = n201 & n401;
  assign n664 = ~pi7  & ~n663;
  assign n665 = ~n489 & ~n664;
  assign n666 = pi7  & ~n93;
  assign n667 = ~pi7  & ~n641;
  assign n668 = pi0  & ~n667;
  assign n669 = ~pi5  & ~n93;
  assign n670 = pi6  & ~n669;
  assign n671 = ~n642 & ~n666;
  assign n672 = ~n670 & n671;
  assign n673 = ~n668 & n672;
  assign n674 = ~n665 & n673;
  assign n675 = ~n653 & n674;
  assign po9  = ~n662 & n675;
  assign n677 = pi8  & ~n41;
  assign n678 = pi2  & n416;
  assign n679 = ~n46 & n678;
  assign n680 = ~n677 & n679;
  assign n681 = ~n423 & ~n680;
  assign n682 = ~pi7  & n344;
  assign po10  = ~n681 & n682;
endmodule
