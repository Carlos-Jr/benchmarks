module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 ;
  wire n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102,
    n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396,
    n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426,
    n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894,
    n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924,
    n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170,
    n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182,
    n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200,
    n3201, n3202, n3203, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212,
    n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242,
    n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272,
    n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302,
    n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332,
    n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362,
    n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3390, n3391, n3392,
    n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416,
    n3417, n3418, n3419, n3420, n3421, n3422,
    n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3439, n3440,
    n3441, n3442, n3443, n3444, n3445, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476,
    n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722,
    n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782,
    n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052,
    n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292,
    n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334,
    n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346,
    n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382,
    n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412,
    n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430,
    n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442,
    n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466,
    n4467, n4468, n4469, n4470, n4471, n4472,
    n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496,
    n4497, n4498, n4499, n4500, n4501, n4502,
    n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526,
    n4527, n4528, n4529, n4530, n4531, n4532,
    n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562,
    n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586,
    n4587, n4588, n4589, n4590, n4591, n4592,
    n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622,
    n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700,
    n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708, n4709, n4710, n4711, n4712,
    n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5040, n5041, n5042,
    n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072,
    n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372,
    n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390,
    n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402,
    n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414,
    n5415, n5416, n5417, n5418, n5419, n5420,
    n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5436, n5437, n5438,
    n5439, n5440, n5441, n5442, n5443, n5444,
    n5445, n5446, n5447, n5448, n5449, n5450,
    n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5460, n5461, n5462,
    n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5470, n5471, n5472, n5473, n5474,
    n5475, n5476, n5477, n5478, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528,
    n5529, n5530, n5531, n5532, n5533, n5534,
    n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5542, n5543, n5544, n5545, n5546,
    n5547, n5548, n5549, n5550, n5551, n5552,
    n5553, n5554, n5555, n5556, n5557, n5558,
    n5559, n5560, n5561, n5562, n5563, n5564,
    n5565, n5566, n5567, n5568, n5569, n5570,
    n5571, n5572, n5573, n5574, n5575, n5576,
    n5577, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588,
    n5589, n5590, n5591, n5592, n5593, n5594,
    n5595, n5596, n5597, n5598, n5599, n5600,
    n5601, n5602, n5603, n5604, n5605, n5606,
    n5607, n5608, n5609, n5610, n5611, n5612,
    n5613, n5614, n5615, n5616, n5617, n5618,
    n5619, n5620, n5621, n5622, n5623, n5624,
    n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636,
    n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648,
    n5649, n5650, n5651, n5652, n5653, n5654,
    n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678,
    n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708,
    n5709, n5710, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5718, n5719, n5720,
    n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732,
    n5733, n5734, n5735, n5736, n5737, n5738,
    n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750,
    n5751, n5752, n5753, n5754, n5755, n5756,
    n5757, n5758, n5759, n5760, n5761, n5762,
    n5763, n5764, n5765, n5766, n5767, n5768,
    n5769, n5770, n5771, n5772, n5773, n5774,
    n5775, n5776, n5777, n5778, n5779, n5780,
    n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792,
    n5793, n5794, n5795, n5796, n5797, n5798,
    n5799, n5800, n5801, n5802, n5803, n5804,
    n5805, n5806, n5807, n5808, n5809, n5810,
    n5811, n5812, n5813, n5814, n5815, n5816,
    n5817, n5818, n5819, n5820, n5821, n5822,
    n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5834,
    n5835, n5836, n5837, n5838, n5839, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846,
    n5847, n5848, n5849, n5850, n5851, n5852,
    n5853, n5854, n5855, n5856, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864,
    n5865, n5866, n5867, n5868, n5869, n5870,
    n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882,
    n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894,
    n5895, n5896, n5897, n5898, n5899, n5900,
    n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912,
    n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924,
    n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954,
    n5955, n5956, n5957, n5958, n5959, n5960,
    n5961, n5962, n5963, n5964, n5965, n5966,
    n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5986, n5987, n5988, n5989, n5990,
    n5991, n5992, n5993, n5994, n5995, n5996,
    n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020,
    n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050,
    n6051, n6052, n6053, n6054, n6055, n6056,
    n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074,
    n6075, n6076, n6077, n6078, n6079, n6080,
    n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110,
    n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122,
    n6123, n6124, n6125, n6126, n6127, n6128,
    n6129, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140,
    n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236,
    n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266,
    n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278,
    n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296,
    n6297, n6298, n6299, n6300, n6301, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326,
    n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362,
    n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386,
    n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398,
    n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416,
    n6417, n6418, n6419, n6420, n6421, n6422,
    n6423, n6424, n6425, n6426, n6427, n6428,
    n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446,
    n6447, n6448, n6449, n6450, n6451, n6452,
    n6453, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470,
    n6471, n6472, n6473, n6474, n6475, n6476,
    n6477, n6478, n6479, n6480, n6481, n6482,
    n6483, n6484, n6485, n6486, n6487, n6488,
    n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500,
    n6501, n6502, n6503, n6504, n6505, n6506,
    n6507, n6508, n6509, n6510, n6511, n6512,
    n6513, n6514, n6515, n6516, n6517, n6518,
    n6519, n6520, n6521, n6522, n6523, n6524,
    n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6533, n6534, n6535, n6536,
    n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548,
    n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566,
    n6567, n6568, n6569, n6570, n6571, n6572,
    n6573, n6574, n6575, n6576, n6577, n6578,
    n6579, n6580, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6588, n6589, n6590,
    n6591, n6592, n6593, n6594, n6595, n6596,
    n6597, n6598, n6599, n6600, n6601, n6602,
    n6603, n6604, n6605, n6606, n6607, n6608,
    n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620,
    n6621, n6622, n6623, n6624, n6625, n6626,
    n6627, n6628, n6629, n6630, n6631, n6632,
    n6633, n6634, n6635, n6636, n6637, n6638,
    n6639, n6640, n6641, n6642, n6643, n6644,
    n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902,
    n6903, n6904, n6905, n6906, n6907, n6908,
    n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6937, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962,
    n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992,
    n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112,
    n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136,
    n7137, n7138, n7139, n7140, n7141, n7142,
    n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154,
    n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172,
    n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214,
    n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370,
    n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400,
    n7401, n7402, n7403, n7404, n7405, n7406,
    n7407, n7408, n7409, n7410, n7411, n7412,
    n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430,
    n7431, n7432, n7433, n7434, n7435, n7436,
    n7437, n7438, n7439, n7440, n7441, n7442,
    n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472,
    n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496,
    n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562,
    n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580,
    n7581, n7582, n7583, n7584, n7585, n7586,
    n7587, n7588, n7589, n7590, n7591, n7592,
    n7593, n7594, n7595, n7596, n7597, n7598,
    n7599, n7600, n7601, n7602, n7603, n7604,
    n7605, n7606, n7607, n7608, n7609, n7610,
    n7611, n7612, n7613, n7614, n7615, n7616,
    n7617, n7618, n7619, n7620, n7621, n7622,
    n7623, n7624, n7625, n7626, n7627, n7628,
    n7629, n7630, n7631, n7632, n7633, n7634,
    n7635, n7636, n7637, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7645, n7646,
    n7647, n7648, n7649, n7650, n7651, n7652,
    n7653, n7654, n7655, n7656, n7657, n7658,
    n7659, n7660, n7661, n7662, n7663, n7664,
    n7665, n7666, n7667, n7668, n7669, n7670,
    n7671, n7672, n7673, n7674, n7675, n7676,
    n7677, n7678, n7679, n7680, n7681, n7682,
    n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694,
    n7695, n7696, n7697, n7698, n7699, n7700,
    n7701, n7702, n7703, n7704, n7705, n7706,
    n7707, n7708, n7709, n7710, n7711, n7712,
    n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724,
    n7725, n7726, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7735, n7736,
    n7737, n7738, n7739, n7740, n7741, n7742,
    n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7760,
    n7761, n7762, n7763, n7764, n7765, n7766,
    n7767, n7768, n7769, n7770, n7771, n7772,
    n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790,
    n7791, n7792, n7793, n7794, n7795, n7796,
    n7797, n7798, n7799, n7800, n7801, n7802,
    n7803, n7804, n7805, n7806, n7807, n7808,
    n7809, n7810, n7811, n7812, n7813, n7814,
    n7815, n7816, n7817, n7818, n7819, n7820,
    n7821, n7822, n7823, n7824, n7825, n7826,
    n7827, n7828, n7829, n7830, n7831, n7832,
    n7833, n7834, n7835, n7836, n7837, n7838,
    n7839, n7840, n7841, n7842, n7843, n7844,
    n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7854, n7855, n7856,
    n7857, n7858, n7859, n7860, n7861, n7862,
    n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886,
    n7887, n7888, n7889, n7890, n7891, n7892,
    n7893, n7894, n7895, n7896, n7897, n7898,
    n7899, n7900, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922,
    n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7948, n7949, n7950, n7951, n7952,
    n7953, n7954, n7955, n7956, n7957, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976,
    n7977, n7978, n7979, n7980, n7981, n7982,
    n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012,
    n8013, n8014, n8015, n8016, n8017, n8018,
    n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042,
    n8043, n8044, n8045, n8046, n8047, n8048,
    n8049, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066,
    n8067, n8068, n8069, n8070, n8071, n8072,
    n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084,
    n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102,
    n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114,
    n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126,
    n8127, n8128, n8129, n8130, n8131, n8132,
    n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144,
    n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156,
    n8157, n8158, n8159, n8160, n8161, n8162,
    n8163, n8164, n8165, n8166, n8167, n8168,
    n8169, n8170, n8171, n8172, n8173, n8174,
    n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186,
    n8187, n8188, n8189, n8190, n8191, n8192,
    n8193, n8194, n8195, n8196, n8197, n8198,
    n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8219, n8220, n8221, n8222,
    n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246,
    n8247, n8248, n8249, n8250, n8251, n8252,
    n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8278, n8279, n8280, n8281, n8282,
    n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8290, n8291, n8292, n8293, n8294,
    n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306,
    n8307, n8308, n8309, n8310, n8311, n8312,
    n8313, n8314, n8315, n8316, n8317, n8318,
    n8319, n8320, n8321, n8322, n8323, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336,
    n8337, n8338, n8339, n8340, n8341, n8342,
    n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366,
    n8367, n8368, n8369, n8370, n8371, n8372,
    n8373, n8374, n8375, n8376, n8377, n8378,
    n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396,
    n8397, n8398, n8399, n8400, n8401, n8402,
    n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456,
    n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486,
    n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564,
    n8565, n8566, n8567, n8568, n8569, n8570,
    n8571, n8572, n8573, n8574, n8575, n8576,
    n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8593, n8594,
    n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606,
    n8607, n8608, n8609, n8610, n8611, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618,
    n8619, n8620, n8621, n8622, n8623, n8624,
    n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648,
    n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678,
    n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708,
    n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726,
    n8727, n8728, n8729, n8730, n8731, n8732,
    n8733, n8734, n8735, n8736, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756,
    n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768,
    n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786,
    n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816,
    n8817, n8818, n8819, n8820, n8821, n8822,
    n8823, n8824, n8825, n8826, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8834,
    n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846,
    n8847, n8848, n8849, n8850, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864,
    n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876,
    n8877, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888,
    n8889, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8902, n8903, n8904, n8905, n8906,
    n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936,
    n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966,
    n8967, n8968, n8969, n8970, n8971, n8972,
    n8973, n8974, n8975, n8976, n8977, n8978,
    n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n8993, n8994, n8995, n8996,
    n8997, n8998, n8999, n9000, n9001, n9002,
    n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9026,
    n9027, n9028, n9029, n9030, n9031, n9032,
    n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050,
    n9051, n9052, n9053, n9054, n9055, n9056,
    n9057, n9058, n9059, n9060, n9061, n9062,
    n9063, n9064, n9065, n9066, n9067, n9068,
    n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9080,
    n9081, n9082, n9083, n9084, n9085, n9086,
    n9087, n9088, n9089, n9090, n9091, n9092,
    n9093, n9094, n9095, n9096, n9097, n9098,
    n9099, n9100, n9101, n9102, n9103, n9104,
    n9105, n9106, n9107, n9108, n9109, n9110,
    n9111, n9112, n9113, n9114, n9115, n9116,
    n9117, n9118, n9119, n9120, n9121, n9122,
    n9123, n9124, n9125, n9126, n9127, n9128,
    n9129, n9130, n9131, n9132, n9133, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140,
    n9141, n9142, n9143, n9144, n9145, n9146,
    n9147, n9148, n9149, n9150, n9151, n9152,
    n9153, n9154, n9155, n9156, n9157, n9158,
    n9159, n9160, n9161, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170,
    n9171, n9172, n9173, n9174, n9175, n9176,
    n9177, n9178, n9179, n9180, n9181, n9182,
    n9183, n9184, n9185, n9186, n9187, n9188,
    n9189, n9190, n9191, n9192, n9193, n9194,
    n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206,
    n9207, n9208, n9209, n9210, n9211, n9212,
    n9213, n9214, n9215, n9216, n9217, n9218,
    n9219, n9220, n9221, n9222, n9223, n9224,
    n9225, n9226, n9227, n9228, n9229, n9230,
    n9231, n9232, n9233, n9234, n9235, n9236,
    n9237, n9238, n9239, n9240, n9241, n9242,
    n9243, n9244, n9245, n9246, n9247, n9248,
    n9249, n9250, n9251, n9252, n9253, n9254,
    n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266,
    n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296,
    n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326,
    n9327, n9328, n9329, n9330, n9331, n9332,
    n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386,
    n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416,
    n9417, n9418, n9419, n9420, n9421, n9422,
    n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446,
    n9447, n9448, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052,
    n10053, n10054, n10055, n10056, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064,
    n10065, n10066, n10067, n10068, n10069, n10070,
    n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10082,
    n10083, n10084, n10085, n10086, n10087, n10088,
    n10089, n10090, n10091, n10092, n10093, n10094,
    n10095, n10096, n10097, n10098, n10099, n10100,
    n10101, n10102, n10103, n10104, n10105, n10106,
    n10107, n10108, n10109, n10110, n10111, n10112,
    n10113, n10114, n10115, n10116, n10117, n10118,
    n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10128, n10129, n10130,
    n10131, n10132, n10133, n10134, n10135, n10136,
    n10137, n10138, n10139, n10140, n10141, n10142,
    n10143, n10144, n10145, n10146, n10147, n10148,
    n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10158, n10159, n10160,
    n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10169, n10170, n10171, n10172,
    n10173, n10174, n10175, n10176, n10177, n10178,
    n10179, n10180, n10181, n10182, n10183, n10184,
    n10185, n10186, n10187, n10188, n10189, n10190,
    n10191, n10192, n10193, n10194, n10195, n10196,
    n10197, n10198, n10199, n10200, n10201, n10202,
    n10203, n10204, n10205, n10206, n10207, n10208,
    n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10222, n10223, n10224, n10225, n10226,
    n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238,
    n10239, n10240, n10241, n10242, n10243, n10244,
    n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256,
    n10257, n10258, n10259, n10260, n10261, n10262,
    n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292,
    n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328,
    n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10370,
    n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382,
    n10383, n10384, n10385, n10386, n10387, n10388,
    n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406,
    n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424,
    n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442,
    n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460,
    n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472,
    n10473, n10474, n10475, n10476, n10477, n10478,
    n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490,
    n10491, n10492, n10493, n10494, n10495, n10496,
    n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514,
    n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532,
    n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10546, n10547, n10548, n10549, n10550,
    n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562,
    n10563, n10564, n10565, n10566, n10567, n10568,
    n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580,
    n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598,
    n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10651, n10652,
    n10653, n10654, n10655, n10656, n10657, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664,
    n10665, n10666, n10667, n10668, n10669, n10670,
    n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706,
    n10707, n10708, n10709, n10710, n10711, n10712,
    n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724,
    n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742,
    n10743, n10744, n10745, n10746, n10747, n10748,
    n10749, n10750, n10751, n10752, n10753, n10754,
    n10755, n10756, n10757, n10758, n10759, n10760,
    n10761, n10762, n10763, n10764, n10765, n10766,
    n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778,
    n10779, n10780, n10781, n10782, n10783, n10784,
    n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868,
    n10869, n10870, n10871, n10872, n10873, n10874,
    n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892,
    n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904,
    n10905, n10906, n10907, n10908, n10909, n10910,
    n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922,
    n10923, n10924, n10925, n10926, n10927, n10928,
    n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940,
    n10941, n10942, n10943, n10944, n10945, n10946,
    n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054,
    n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066,
    n11067, n11068, n11069, n11070, n11071, n11072,
    n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084,
    n11085, n11086, n11087, n11088, n11089, n11090,
    n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108,
    n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126,
    n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144,
    n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156,
    n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174,
    n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11189, n11190, n11191, n11192,
    n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204,
    n11205, n11206, n11207, n11208, n11209, n11210,
    n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222,
    n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11242, n11243, n11244, n11245, n11246,
    n11247, n11248, n11249, n11250, n11251, n11252,
    n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264,
    n11265, n11266, n11267, n11268, n11269, n11270,
    n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282,
    n11283, n11284, n11285, n11286, n11287, n11288,
    n11289, n11290, n11291, n11292, n11293, n11294,
    n11295, n11296, n11297, n11298, n11299, n11300,
    n11301, n11302, n11303, n11304, n11305, n11306,
    n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318,
    n11319, n11320, n11321, n11322, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336,
    n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354,
    n11355, n11356, n11357, n11358, n11359, n11360,
    n11361, n11362, n11363, n11364, n11365, n11366,
    n11367, n11368, n11369, n11370, n11371, n11372,
    n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11394, n11395, n11396,
    n11397, n11398, n11399, n11400, n11401, n11402,
    n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414,
    n11415, n11416, n11417, n11418, n11419, n11420,
    n11421, n11422, n11423, n11424, n11425, n11426,
    n11427, n11428, n11429, n11430, n11431, n11432,
    n11433, n11434, n11435, n11436, n11437, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444,
    n11445, n11446, n11447, n11448, n11449, n11450,
    n11451, n11452, n11453, n11454, n11455, n11456,
    n11457, n11458, n11459, n11460, n11461, n11462,
    n11463, n11464, n11465, n11466, n11467, n11468,
    n11469, n11470, n11471, n11472, n11473, n11474,
    n11475, n11476, n11477, n11478, n11479, n11480,
    n11481, n11482, n11483, n11484, n11485, n11486,
    n11487, n11488, n11489, n11490, n11491, n11492,
    n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504,
    n11505, n11506, n11507, n11508, n11509, n11510,
    n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11520, n11521, n11522,
    n11523, n11524, n11525, n11526, n11527, n11528,
    n11529, n11530, n11531, n11532, n11533, n11534,
    n11535, n11536, n11537, n11538, n11539, n11540,
    n11541, n11542, n11543, n11544, n11545, n11546,
    n11547, n11548, n11549, n11550, n11551, n11552,
    n11553, n11554, n11555, n11556, n11557, n11558,
    n11559, n11560, n11561, n11562, n11563, n11564,
    n11565, n11566, n11567, n11568, n11569, n11570,
    n11571, n11572, n11573, n11574, n11575, n11576,
    n11577, n11578, n11579, n11580, n11581, n11582,
    n11583, n11584, n11585, n11586, n11587, n11588,
    n11589, n11590, n11591, n11592, n11593, n11594,
    n11595, n11596, n11597, n11598, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618,
    n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630,
    n11631, n11632, n11633, n11634, n11635, n11636,
    n11637, n11638, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11648,
    n11649, n11650, n11651, n11652, n11653, n11654,
    n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666,
    n11667, n11668, n11669, n11670, n11671, n11672,
    n11673, n11674, n11675, n11676, n11677, n11678,
    n11679, n11680, n11681, n11682, n11683, n11684,
    n11685, n11686, n11687, n11688, n11689, n11690,
    n11691, n11692, n11693, n11694, n11695, n11696,
    n11697, n11698, n11699, n11700, n11701, n11702,
    n11703, n11704, n11705, n11706, n11707, n11708,
    n11709, n11710, n11711, n11712, n11713, n11714,
    n11715, n11716, n11717, n11718, n11719, n11720,
    n11721, n11722, n11723, n11724, n11725, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756,
    n11757, n11758, n11759, n11760, n11761, n11762,
    n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774,
    n11775, n11776, n11777, n11778, n11779, n11780,
    n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792,
    n11793, n11794, n11795, n11796, n11797, n11798,
    n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810,
    n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218,
    n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236,
    n12237, n12238, n12239, n12240, n12241, n12242,
    n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254,
    n12255, n12256, n12257, n12258, n12259, n12260,
    n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272,
    n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290,
    n12291, n12292, n12293, n12294, n12295, n12296,
    n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314,
    n12315, n12316, n12317, n12318, n12319, n12320,
    n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12340, n12341, n12342, n12343, n12344,
    n12345, n12346, n12347, n12348, n12349, n12350,
    n12351, n12352, n12353, n12354, n12355, n12356,
    n12357, n12358, n12359, n12360, n12361, n12362,
    n12363, n12364, n12365, n12366, n12367, n12368,
    n12369, n12370, n12371, n12372, n12373, n12374,
    n12375, n12376, n12377, n12378, n12379, n12380,
    n12381, n12382, n12383, n12384, n12385, n12386,
    n12387, n12388, n12389, n12390, n12391, n12392,
    n12393, n12394, n12395, n12396, n12397, n12398,
    n12399, n12400, n12401, n12402, n12403, n12404,
    n12405, n12406, n12407, n12408, n12409, n12410,
    n12411, n12412, n12413, n12414, n12415, n12416,
    n12417, n12418, n12419, n12420, n12421, n12422,
    n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434,
    n12435, n12436, n12437, n12438, n12439, n12440,
    n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452,
    n12453, n12454, n12455, n12456, n12457, n12458,
    n12459, n12460, n12461, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470,
    n12471, n12472, n12473, n12474, n12475, n12476,
    n12477, n12478, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488,
    n12489, n12490, n12491, n12492, n12493, n12494,
    n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506,
    n12507, n12508, n12509, n12510, n12511, n12512,
    n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524,
    n12525, n12526, n12527, n12528, n12529, n12530,
    n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542,
    n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560,
    n12561, n12562, n12563, n12564, n12565, n12566,
    n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578,
    n12579, n12580, n12581, n12582, n12583, n12584,
    n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596,
    n12597, n12598, n12599, n12600, n12601, n12602,
    n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614,
    n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632,
    n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650,
    n12651, n12652, n12653, n12654, n12655, n12656,
    n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668,
    n12669, n12670, n12671, n12672, n12673, n12674,
    n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12691, n12692,
    n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704,
    n12705, n12706, n12707, n12708, n12709, n12710,
    n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722,
    n12723, n12724, n12725, n12726, n12727, n12728,
    n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740,
    n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758,
    n12759, n12760, n12761, n12762, n12763, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776,
    n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794,
    n12795, n12796, n12797, n12798, n12799, n12800,
    n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812,
    n12813, n12814, n12815, n12816, n12817, n12818,
    n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12830,
    n12831, n12832, n12833, n12834, n12835, n12836,
    n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848,
    n12849, n12850, n12851, n12852, n12853, n12854,
    n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866,
    n12867, n12868, n12869, n12870, n12871, n12872,
    n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884,
    n12885, n12886, n12887, n12888, n12889, n12890,
    n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902,
    n12903, n12904, n12905, n12906, n12907, n12908,
    n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920,
    n12921, n12922, n12923, n12924, n12925, n12926,
    n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938,
    n12939, n12940, n12941, n12942, n12943, n12944,
    n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956,
    n12957, n12958, n12959, n12960, n12961, n12962,
    n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974,
    n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010,
    n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028,
    n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046,
    n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058,
    n13059, n13060, n13061, n13062, n13063, n13064,
    n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13073, n13074, n13075, n13076,
    n13077, n13078, n13079, n13080, n13081, n13082,
    n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100,
    n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112,
    n13113, n13114, n13115, n13116, n13117, n13118,
    n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130,
    n13131, n13132, n13133, n13134, n13135, n13136,
    n13137, n13138, n13139, n13140, n13141, n13142,
    n13143, n13144, n13145, n13146, n13147, n13148,
    n13149, n13150, n13151, n13152, n13153, n13154,
    n13155, n13156, n13157, n13158, n13159, n13160,
    n13161, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232,
    n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322,
    n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13354, n13355, n13356, n13357, n13358,
    n13359, n13360, n13361, n13362, n13363, n13364,
    n13365, n13366, n13367, n13368, n13369, n13370,
    n13371, n13372, n13373, n13374, n13375, n13376,
    n13377, n13378, n13379, n13380, n13381, n13382,
    n13383, n13384, n13385, n13386, n13387, n13388,
    n13389, n13390, n13391, n13392, n13393, n13394,
    n13395, n13396, n13397, n13398, n13399, n13400,
    n13401, n13402, n13403, n13404, n13405, n13406,
    n13407, n13408, n13409, n13410, n13411, n13412,
    n13413, n13414, n13415, n13416, n13417, n13418,
    n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430,
    n13431, n13432, n13433, n13434, n13435, n13436,
    n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448,
    n13449, n13450, n13451, n13452, n13453, n13454,
    n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13464, n13465, n13466,
    n13467, n13468, n13469, n13470, n13471, n13472,
    n13473, n13474, n13475, n13476, n13477, n13478,
    n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13486, n13487, n13488, n13489, n13490,
    n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502,
    n13503, n13504, n13505, n13506, n13507, n13508,
    n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13516, n13517, n13518, n13519, n13520,
    n13521, n13522, n13523, n13524, n13525, n13526,
    n13527, n13528, n13529, n13530, n13531, n13532,
    n13533, n13534, n13535, n13536, n13537, n13538,
    n13539, n13540, n13541, n13542, n13543, n13544,
    n13545, n13546, n13547, n13548, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562,
    n13563, n13564, n13565, n13566, n13567, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580,
    n13581, n13582, n13583, n13584, n13585, n13586,
    n13587, n13588, n13589, n13590, n13591, n13592,
    n13593, n13594, n13595, n13596, n13597, n13598,
    n13599, n13600, n13601, n13602, n13603, n13604,
    n13605, n13606, n13607, n13608, n13609, n13610,
    n13611, n13612, n13613, n13614, n13615, n13616,
    n13617, n13618, n13619, n13620, n13621, n13622,
    n13623, n13624, n13625, n13626, n13627, n13628,
    n13629, n13630, n13631, n13632, n13633, n13634,
    n13635, n13636, n13637, n13638, n13639, n13640,
    n13641, n13642, n13643, n13644, n13645, n13646,
    n13647, n13648, n13649, n13650, n13651, n13652,
    n13653, n13654, n13655, n13656, n13657, n13658,
    n13659, n13660, n13661, n13662, n13663, n13664,
    n13665, n13666, n13667, n13668, n13669, n13670,
    n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682,
    n13683, n13684, n13685, n13686, n13687, n13688,
    n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700,
    n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718,
    n13719, n13720, n13721, n13722, n13723, n13724,
    n13725, n13726, n13727, n13728, n13729, n13730,
    n13731, n13732, n13733, n13734, n13735, n13736,
    n13737, n13738, n13739, n13740, n13741, n13742,
    n13743, n13744, n13745, n13746, n13747, n13748,
    n13749, n13750, n13751, n13752, n13753, n13754,
    n13755, n13756, n13757, n13758, n13759, n13760,
    n13761, n13762, n13763, n13764, n13765, n13766,
    n13767, n13768, n13769, n13770, n13771, n13772,
    n13773, n13774, n13775, n13776, n13777, n13778,
    n13779, n13780, n13781, n13782, n13783, n13784,
    n13785, n13786, n13787, n13788, n13789, n13790,
    n13791, n13792, n13793, n13794, n13795, n13796,
    n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808,
    n13809, n13810, n13811, n13812, n13813, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826,
    n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844,
    n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862,
    n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880,
    n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898,
    n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916,
    n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934,
    n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952,
    n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970,
    n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988,
    n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006,
    n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060,
    n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078,
    n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144,
    n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330,
    n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348,
    n14349, n14350, n14351, n14352, n14353, n14354,
    n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372,
    n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14381, n14382, n14383, n14384,
    n14385, n14386, n14387, n14388, n14389, n14390,
    n14391, n14392, n14393, n14394, n14395, n14396,
    n14397, n14398, n14399, n14400, n14401, n14402,
    n14403, n14404, n14405, n14406, n14407, n14408,
    n14409, n14410, n14411, n14412, n14413, n14414,
    n14415, n14416, n14417, n14418, n14419, n14420,
    n14421, n14422, n14423, n14424, n14425, n14426,
    n14427, n14428, n14429, n14430, n14431, n14432,
    n14433, n14434, n14435, n14436, n14437, n14438,
    n14439, n14440, n14441, n14442, n14443, n14444,
    n14445, n14446, n14447, n14448, n14449, n14450,
    n14451, n14452, n14453, n14454, n14455, n14456,
    n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468,
    n14469, n14470, n14471, n14472, n14473, n14474,
    n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486,
    n14487, n14488, n14489, n14490, n14491, n14492,
    n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504,
    n14505, n14506, n14507, n14508, n14509, n14510,
    n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522,
    n14523, n14524, n14525, n14526, n14527, n14528,
    n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540,
    n14541, n14542, n14543, n14544, n14545, n14546,
    n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558,
    n14559, n14560, n14561, n14562, n14563, n14564,
    n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576,
    n14577, n14578, n14579, n14580, n14581, n14582,
    n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594,
    n14595, n14596, n14597, n14598, n14599, n14600,
    n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612,
    n14613, n14614, n14615, n14616, n14617, n14618,
    n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630,
    n14631, n14632, n14633, n14634, n14635, n14636,
    n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648,
    n14649, n14650, n14651, n14652, n14653, n14654,
    n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666,
    n14667, n14668, n14669, n14670, n14671, n14672,
    n14673, n14674, n14675, n14676, n14677, n14678,
    n14679, n14680, n14681, n14682, n14683, n14684,
    n14685, n14686, n14687, n14688, n14689, n14690,
    n14691, n14692, n14693, n14694, n14695, n14696,
    n14697, n14698, n14699, n14700, n14701, n14702,
    n14703, n14704, n14705, n14706, n14707, n14708,
    n14709, n14710, n14711, n14712, n14713, n14714,
    n14715, n14716, n14717, n14718, n14719, n14720,
    n14721, n14722, n14723, n14724, n14725, n14726,
    n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738,
    n14739, n14740, n14741, n14742, n14743, n14744,
    n14745, n14746, n14747, n14748, n14749, n14750,
    n14751, n14752, n14753, n14754, n14755, n14756,
    n14757, n14758, n14759, n14760, n14761, n14762,
    n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816,
    n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834,
    n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846,
    n14847, n14848, n14849, n14850, n14851, n14852,
    n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864,
    n14865, n14866, n14867, n14868, n14869, n14870,
    n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882,
    n14883, n14884, n14885, n14886, n14887, n14888,
    n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906,
    n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924,
    n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942,
    n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978,
    n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996,
    n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014,
    n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032,
    n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050,
    n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068,
    n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086,
    n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122,
    n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194,
    n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230,
    n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248,
    n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15281, n15282, n15283, n15284,
    n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302,
    n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314,
    n15315, n15316, n15317, n15318, n15319, n15320,
    n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338,
    n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15355, n15356,
    n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368,
    n15369, n15370, n15371, n15372, n15373, n15374,
    n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392,
    n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404,
    n15405, n15406, n15407, n15408, n15409, n15410,
    n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422,
    n15423, n15424, n15425, n15426, n15427, n15428,
    n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440,
    n15441, n15442, n15443, n15444, n15445, n15446,
    n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458,
    n15459, n15460, n15461, n15462, n15463, n15464,
    n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476,
    n15477, n15478, n15479, n15480, n15481, n15482,
    n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494,
    n15495, n15496, n15497, n15498, n15499, n15500,
    n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512,
    n15513, n15514, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530,
    n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15768, n15769, n15770,
    n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782,
    n15783, n15784, n15785, n15786, n15787, n15788,
    n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800,
    n15801, n15802, n15803, n15804, n15805, n15806,
    n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824,
    n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854,
    n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872,
    n15873, n15874, n15875, n15876, n15877, n15878,
    n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890,
    n15891, n15892, n15893, n15894, n15895, n15896,
    n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908,
    n15909, n15910, n15911, n15912, n15913, n15914,
    n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926,
    n15927, n15928, n15929, n15930, n15931, n15932,
    n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944,
    n15945, n15946, n15947, n15948, n15949, n15950,
    n15951, n15952, n15953, n15954, n15955, n15956,
    n15957, n15958, n15959, n15960, n15961, n15962,
    n15963, n15964, n15965, n15966, n15967, n15968,
    n15969, n15970, n15971, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980,
    n15981, n15982, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998,
    n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016,
    n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034,
    n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106,
    n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178,
    n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196,
    n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214,
    n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232,
    n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250,
    n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262,
    n16263, n16264, n16265, n16266, n16267, n16268,
    n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280,
    n16281, n16282, n16283, n16284, n16285, n16286,
    n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16302, n16303, n16304,
    n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316,
    n16317, n16318, n16319, n16320, n16321, n16322,
    n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334,
    n16335, n16336, n16337, n16338, n16339, n16340,
    n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352,
    n16353, n16354, n16355, n16356, n16357, n16358,
    n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370,
    n16371, n16372, n16373, n16374, n16375, n16376,
    n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388,
    n16389, n16390, n16391, n16392, n16393, n16394,
    n16395, n16396, n16397, n16398, n16399, n16400,
    n16401, n16402, n16403, n16404, n16405, n16406,
    n16407, n16408, n16409, n16410, n16411, n16412,
    n16413, n16414, n16415, n16416, n16417, n16418,
    n16419, n16420, n16421, n16422, n16423, n16424,
    n16425, n16426, n16427, n16428, n16429, n16430,
    n16431, n16432, n16433, n16434, n16435, n16436,
    n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448,
    n16449, n16450, n16451, n16452, n16453, n16454,
    n16455, n16456, n16457, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466,
    n16467, n16468, n16469, n16470, n16471, n16472,
    n16473, n16474, n16475, n16476, n16477, n16478,
    n16479, n16480, n16481, n16482, n16483, n16484,
    n16485, n16486, n16487, n16488, n16489, n16490,
    n16491, n16492, n16493, n16494, n16495, n16496,
    n16497, n16498, n16499, n16500, n16501, n16502,
    n16503, n16504, n16505, n16506, n16507, n16508,
    n16509, n16510, n16511, n16512, n16513, n16514,
    n16515, n16516, n16517, n16518, n16519, n16520,
    n16521, n16522, n16523, n16524, n16525, n16526,
    n16527, n16528, n16529, n16530, n16531, n16532,
    n16533, n16534, n16535, n16536, n16537, n16538,
    n16539, n16540, n16541, n16542, n16543, n16544,
    n16545, n16546, n16547, n16548, n16549, n16550,
    n16551, n16552, n16553, n16554, n16555, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562,
    n16563, n16564, n16565, n16566, n16567, n16568,
    n16569, n16570, n16571, n16572, n16573, n16574,
    n16575, n16576, n16577, n16578, n16579, n16580,
    n16581, n16582, n16583, n16584, n16585, n16586,
    n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598,
    n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652,
    n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670,
    n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16687, n16688,
    n16689, n16690, n16691, n16692, n16693, n16694,
    n16695, n16696, n16697, n16698, n16699, n16700,
    n16701, n16702, n16703, n16704, n16705, n16706,
    n16707, n16708, n16709, n16710, n16711, n16712,
    n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724,
    n16725, n16726, n16727, n16728, n16729, n16730,
    n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742,
    n16743, n16744, n16745, n16746, n16747, n16748,
    n16749, n16750, n16751, n16752, n16753, n16754,
    n16755, n16756, n16757, n16758, n16759, n16760,
    n16761, n16762, n16763, n16764, n16765, n16766,
    n16767, n16768, n16769, n16770, n16771, n16772,
    n16773, n16774, n16775, n16776, n16777, n16778,
    n16779, n16780, n16781, n16782, n16783, n16784,
    n16785, n16786, n16787, n16788, n16789, n16790,
    n16791, n16792, n16793, n16794, n16795, n16796,
    n16797, n16798, n16799, n16800, n16801, n16802,
    n16803, n16804, n16805, n16806, n16807, n16808,
    n16809, n16810, n16811, n16812, n16813, n16814,
    n16815, n16816, n16817, n16818, n16819, n16820,
    n16821, n16822, n16823, n16824, n16825, n16826,
    n16827, n16828, n16829, n16830, n16831, n16832,
    n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844,
    n16845, n16846, n16847, n16848, n16849, n16850,
    n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16868,
    n16869, n16870, n16871, n16872, n16873, n16874,
    n16875, n16876, n16877, n16878, n16879, n16880,
    n16881, n16882, n16883, n16884, n16885, n16886,
    n16887, n16888, n16889, n16890, n16891, n16892,
    n16893, n16894, n16895, n16896, n16897, n16898,
    n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16906, n16907, n16908, n16909, n16910,
    n16911, n16912, n16913, n16914, n16915, n16916,
    n16917, n16918, n16919, n16920, n16921, n16922,
    n16923, n16924, n16925, n16926, n16927, n16928,
    n16929, n16930, n16931, n16932, n16933, n16934,
    n16935, n16936, n16937, n16938, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16952,
    n16953, n16954, n16955, n16956, n16957, n16958,
    n16959, n16960, n16961, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976,
    n16977, n16978, n16979, n16980, n16981, n16982,
    n16983, n16984, n16985, n16986, n16987, n16988,
    n16989, n16990, n16991, n16992, n16993, n16994,
    n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17004, n17005, n17006,
    n17007, n17008, n17009, n17010, n17011, n17012,
    n17013, n17014, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024,
    n17025, n17026, n17027, n17028, n17029, n17030,
    n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042,
    n17043, n17044, n17045, n17046, n17047, n17048,
    n17049, n17050, n17051, n17052, n17053, n17054,
    n17055, n17056, n17057, n17058, n17059, n17060,
    n17061, n17062, n17063, n17064, n17065, n17066,
    n17067, n17068, n17069, n17070, n17071, n17072,
    n17073, n17074, n17075, n17076, n17077, n17078,
    n17079, n17080, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090,
    n17091, n17092, n17093, n17094, n17095, n17096,
    n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17114,
    n17115, n17116, n17117, n17118, n17119, n17120,
    n17121, n17122, n17123, n17124, n17125, n17126,
    n17127, n17128, n17129, n17130, n17131, n17132,
    n17133, n17134, n17135, n17136, n17137, n17138,
    n17139, n17140, n17141, n17142, n17143, n17144,
    n17145, n17146, n17147, n17148, n17149, n17150,
    n17151, n17152, n17153, n17154, n17155, n17156,
    n17157, n17158, n17159, n17160, n17161, n17162,
    n17163, n17164, n17165, n17166, n17167, n17168,
    n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180,
    n17181, n17182, n17183, n17184, n17185, n17186,
    n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204,
    n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222,
    n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240,
    n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258,
    n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276,
    n17277, n17278, n17279, n17280, n17281, n17282,
    n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294,
    n17295, n17296, n17297, n17298, n17299, n17300,
    n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312,
    n17313, n17314, n17315, n17316, n17317, n17318,
    n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330,
    n17331, n17332, n17333, n17334, n17335, n17336,
    n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348,
    n17349, n17350, n17351, n17352, n17353, n17354,
    n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366,
    n17367, n17368, n17369, n17370, n17371, n17372,
    n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384,
    n17385, n17386, n17387, n17388, n17389, n17390,
    n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402,
    n17403, n17404, n17405, n17406, n17407, n17408,
    n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420,
    n17421, n17422, n17423, n17424, n17425, n17426,
    n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438,
    n17439, n17440, n17441, n17442, n17443, n17444,
    n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456,
    n17457, n17458, n17459, n17460, n17461, n17462,
    n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474,
    n17475, n17476, n17477, n17478, n17479, n17480,
    n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492,
    n17493, n17494, n17495, n17496, n17497, n17498,
    n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510,
    n17511, n17512, n17513, n17514, n17515, n17516,
    n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528,
    n17529, n17530, n17531, n17532, n17533, n17534,
    n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546,
    n17547, n17548, n17549, n17550, n17551, n17552,
    n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564,
    n17565, n17566, n17567, n17568, n17569, n17570,
    n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582,
    n17583, n17584, n17585, n17586, n17587, n17588,
    n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624,
    n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672,
    n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696,
    n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708,
    n17709, n17710, n17711, n17712, n17713, n17714,
    n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726,
    n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744,
    n17745, n17746, n17747, n17748, n17749, n17750,
    n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762,
    n17763, n17764, n17765, n17766, n17767, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780,
    n17781, n17782, n17783, n17784, n17785, n17786,
    n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798,
    n17799, n17800, n17801, n17802, n17803, n17804,
    n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816,
    n17817, n17818, n17819, n17820, n17821, n17822,
    n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834,
    n17835, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852,
    n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888,
    n17889, n17890, n17891, n17892, n17893, n17894,
    n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906,
    n17907, n17908, n17909, n17910, n17911, n17912,
    n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17923, n17924,
    n17925, n17926, n17927, n17928, n17929, n17930,
    n17931, n17932, n17933, n17934, n17935, n17936,
    n17937, n17938, n17939, n17940, n17941, n17942,
    n17943, n17944, n17945, n17946, n17947, n17948,
    n17949, n17950, n17951, n17952, n17953, n17954,
    n17955, n17956, n17957, n17958, n17959, n17960,
    n17961, n17962, n17963, n17964, n17965, n17966,
    n17967, n17968, n17969, n17970, n17971, n17972,
    n17973, n17974, n17975, n17976, n17977, n17978,
    n17979, n17980, n17981, n17982, n17983, n17984,
    n17985, n17986, n17987, n17988, n17989, n17990,
    n17991, n17992, n17993, n17994, n17995, n17996,
    n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014,
    n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032,
    n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050,
    n18051, n18052, n18053, n18054, n18055, n18056,
    n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068,
    n18069, n18070, n18071, n18072, n18073, n18074,
    n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086,
    n18087, n18088, n18089, n18090, n18091, n18092,
    n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104,
    n18105, n18106, n18107, n18108, n18109, n18110,
    n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122,
    n18123, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140,
    n18141, n18142, n18143, n18144, n18145, n18146,
    n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158,
    n18159, n18160, n18161, n18162, n18163, n18164,
    n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176,
    n18177, n18178, n18179, n18180, n18181, n18182,
    n18183, n18184, n18185, n18186, n18187, n18188,
    n18189, n18190, n18191, n18192, n18193, n18194,
    n18195, n18196, n18197, n18198, n18199, n18200,
    n18201, n18202, n18203, n18204, n18205, n18206,
    n18207, n18208, n18209, n18210, n18211, n18212,
    n18213, n18214, n18215, n18216, n18217, n18218,
    n18219, n18220, n18221, n18222, n18223, n18224,
    n18225, n18226, n18227, n18228, n18229, n18230,
    n18231, n18232, n18233, n18234, n18235, n18236,
    n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18248,
    n18249, n18250, n18251, n18252, n18253, n18254,
    n18255, n18256, n18257, n18258, n18259, n18260,
    n18261, n18262, n18263, n18264, n18265, n18266,
    n18267, n18268, n18269, n18270, n18271, n18272,
    n18273, n18274, n18275, n18276, n18277, n18278,
    n18279, n18280, n18281, n18282, n18283, n18284,
    n18285, n18286, n18287, n18288, n18289, n18290,
    n18291, n18292, n18293, n18294, n18295, n18296,
    n18297, n18298, n18299, n18300, n18301, n18302,
    n18303, n18304, n18305, n18306, n18307, n18308,
    n18309, n18310, n18311, n18312, n18313, n18314,
    n18315, n18316, n18317, n18318, n18319, n18320,
    n18321, n18322, n18323, n18324, n18325, n18326,
    n18327, n18328, n18329, n18330, n18331, n18332,
    n18333, n18334, n18335, n18336, n18337, n18338,
    n18339, n18340, n18341, n18342, n18343, n18344,
    n18345, n18346, n18347, n18348, n18349, n18350,
    n18351, n18352, n18353, n18354, n18355, n18356,
    n18357, n18358, n18359, n18360, n18361, n18362,
    n18363, n18364, n18365, n18366, n18367, n18368,
    n18369, n18370, n18371, n18372, n18373, n18374,
    n18375, n18376, n18377, n18378, n18379, n18380,
    n18381, n18382, n18383, n18384, n18385, n18386,
    n18387, n18388, n18389, n18390, n18391, n18392,
    n18393, n18394, n18395, n18396, n18397, n18398,
    n18399, n18400, n18401, n18402, n18403, n18404,
    n18405, n18406, n18407, n18408, n18409, n18410,
    n18411, n18412, n18413, n18414, n18415, n18416,
    n18417, n18418, n18419, n18420, n18421, n18422,
    n18423, n18424, n18425, n18426, n18427, n18428,
    n18429, n18430, n18431, n18432, n18433, n18434,
    n18435, n18436, n18437, n18438, n18439, n18440,
    n18441, n18442, n18443, n18444, n18445, n18446,
    n18447, n18448, n18449, n18450, n18451, n18452,
    n18453, n18454, n18455, n18456, n18457, n18458,
    n18459, n18460, n18461, n18462, n18463, n18464,
    n18465, n18466, n18467, n18468, n18469, n18470,
    n18471, n18472, n18473, n18474, n18475, n18476,
    n18477, n18478, n18479, n18480, n18481, n18482,
    n18483, n18484, n18485, n18486, n18487, n18488,
    n18489, n18490, n18491, n18492, n18493, n18494,
    n18495, n18496, n18497, n18498, n18499, n18500,
    n18501, n18502, n18503, n18504, n18505, n18506,
    n18507, n18508, n18509, n18510, n18511, n18512,
    n18513, n18514, n18515, n18516, n18517, n18518,
    n18519, n18520, n18521, n18522, n18523, n18524,
    n18525, n18526, n18527, n18528, n18529, n18530,
    n18531, n18532, n18533, n18534, n18535, n18536,
    n18537, n18538, n18539, n18540, n18541, n18542,
    n18543, n18544, n18545, n18546, n18547, n18548,
    n18549, n18550, n18551, n18552, n18553, n18554,
    n18555, n18556, n18557, n18558, n18559, n18560,
    n18561, n18562, n18563, n18564, n18565, n18566,
    n18567, n18568, n18569, n18570, n18571, n18572,
    n18573, n18574, n18575, n18576, n18577, n18578,
    n18579, n18580, n18581, n18582, n18583, n18584,
    n18585, n18586, n18587, n18588, n18589, n18590,
    n18591, n18592, n18593, n18594, n18595, n18596,
    n18597, n18598, n18599, n18600, n18601, n18602,
    n18603, n18604, n18605, n18606, n18607, n18608,
    n18609, n18610, n18611, n18612, n18613, n18614,
    n18615, n18616, n18617, n18618, n18619, n18620,
    n18621, n18622, n18623, n18624, n18625, n18626,
    n18627, n18628, n18629, n18630, n18631, n18632,
    n18633, n18634, n18635, n18636, n18637, n18638,
    n18639, n18640, n18641, n18642, n18643, n18644,
    n18645, n18646, n18647, n18648, n18649, n18650,
    n18651, n18652, n18653, n18654, n18655, n18656,
    n18657, n18658, n18659, n18660, n18661, n18662,
    n18663, n18664, n18665, n18666, n18667, n18668,
    n18669, n18670, n18671, n18672, n18673, n18674,
    n18675, n18676, n18677, n18678, n18679, n18680,
    n18681, n18682, n18683, n18684, n18685, n18686,
    n18687, n18688, n18689, n18690, n18691, n18692,
    n18693, n18694, n18695, n18696, n18697, n18698,
    n18699, n18700, n18701, n18702, n18703, n18704,
    n18705, n18706, n18707, n18708, n18709, n18710,
    n18711, n18712, n18713, n18714, n18715, n18716,
    n18717, n18718, n18719, n18720, n18721, n18722,
    n18723, n18724, n18725, n18726, n18727, n18728,
    n18729, n18730, n18731, n18732, n18733, n18734,
    n18735, n18736, n18737, n18738, n18739, n18740,
    n18741, n18742, n18743, n18744, n18745, n18746,
    n18747, n18748, n18749, n18750, n18751, n18752,
    n18753, n18754, n18755, n18756, n18757, n18758,
    n18759, n18760, n18761, n18762, n18763, n18764,
    n18765, n18766, n18767, n18768, n18769, n18770,
    n18771, n18772, n18773, n18774, n18775, n18776,
    n18777, n18778, n18779, n18780, n18781, n18782,
    n18783, n18784, n18785, n18786, n18787, n18788,
    n18789, n18790, n18791, n18792, n18793, n18794,
    n18795, n18796, n18797, n18798, n18799, n18800,
    n18801, n18802, n18803, n18804, n18805, n18806,
    n18807, n18808, n18809, n18810, n18811, n18812,
    n18813, n18814, n18815, n18816, n18817, n18818,
    n18819, n18820, n18821, n18822, n18823, n18824,
    n18825, n18826, n18827, n18828, n18829, n18830,
    n18831, n18832, n18833, n18834, n18835, n18836,
    n18837, n18838, n18839, n18840, n18841, n18842,
    n18843, n18844, n18845, n18846, n18847, n18848,
    n18849, n18850, n18851, n18852, n18853, n18854,
    n18855, n18856, n18857, n18858, n18859, n18860,
    n18861, n18862, n18863, n18864, n18865, n18866,
    n18867, n18868, n18869, n18870, n18871, n18872,
    n18873, n18874, n18875, n18876, n18877, n18878,
    n18879, n18880, n18881, n18882, n18883, n18884,
    n18885, n18886, n18887, n18888, n18889, n18890,
    n18891, n18892, n18893, n18894, n18895, n18896,
    n18897, n18898, n18899, n18900, n18901, n18902,
    n18903, n18904, n18905, n18906, n18907, n18908,
    n18909, n18910, n18911, n18912, n18913, n18914,
    n18915, n18916, n18917, n18918, n18919, n18920,
    n18921, n18922, n18923, n18924, n18925, n18926,
    n18927, n18928, n18929, n18930, n18931, n18932,
    n18933, n18934, n18935, n18936, n18937, n18938,
    n18939, n18940, n18941, n18942, n18943, n18944,
    n18945, n18946, n18947, n18948, n18949, n18950,
    n18951, n18952, n18953, n18954, n18955, n18956,
    n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968,
    n18969, n18970, n18971, n18972, n18973, n18974,
    n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986,
    n18987, n18988, n18989, n18990, n18991, n18992,
    n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004,
    n19005, n19006, n19007, n19008, n19009, n19010,
    n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022,
    n19023, n19024, n19025, n19026, n19027, n19028,
    n19029, n19030, n19031, n19032, n19033, n19034,
    n19035, n19036, n19037, n19038, n19039, n19040,
    n19041, n19042, n19043, n19044, n19045, n19046,
    n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058,
    n19059, n19060, n19061, n19062, n19063, n19064,
    n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076,
    n19077, n19078, n19079, n19080, n19081, n19082,
    n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094,
    n19095, n19096, n19097, n19098, n19099, n19100,
    n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112,
    n19113, n19114, n19115, n19116, n19117, n19118,
    n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130,
    n19131, n19132, n19133, n19134, n19135, n19136,
    n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148,
    n19149, n19150, n19151, n19152, n19153, n19154,
    n19155, n19156, n19157, n19158, n19159, n19160,
    n19161, n19162, n19163, n19164, n19165, n19166,
    n19167, n19168, n19169, n19170, n19171, n19172,
    n19173, n19174, n19175, n19176, n19177, n19178,
    n19179, n19180, n19181, n19182, n19183, n19184,
    n19185, n19186, n19187, n19188, n19189, n19190,
    n19191, n19192, n19193, n19194, n19195, n19196,
    n19197, n19198, n19199, n19200, n19201, n19202,
    n19203, n19204, n19205, n19206, n19207, n19208,
    n19209, n19210, n19211, n19212, n19213, n19214,
    n19215, n19216, n19217, n19218, n19219, n19220,
    n19221, n19222, n19223, n19224, n19225, n19226,
    n19227, n19228, n19229, n19230, n19231, n19232,
    n19233, n19234, n19235, n19236, n19237, n19238,
    n19239, n19240, n19241, n19242, n19243, n19244,
    n19245, n19246, n19247, n19248, n19249, n19250,
    n19251, n19252, n19253, n19254, n19255, n19256,
    n19257, n19258, n19259, n19260, n19261, n19262,
    n19263, n19264, n19265, n19266, n19267, n19268,
    n19269, n19270, n19271, n19272, n19273, n19274,
    n19275, n19276, n19277, n19278, n19279, n19280,
    n19281, n19282, n19283, n19284, n19285, n19286,
    n19287, n19288, n19289, n19290, n19291, n19292,
    n19293, n19294, n19295, n19296, n19297, n19298,
    n19299, n19300, n19301, n19302, n19303, n19304,
    n19305, n19306, n19307, n19308, n19309, n19310,
    n19311, n19312, n19313, n19314, n19315, n19316,
    n19317, n19318, n19319, n19320, n19321, n19322,
    n19323, n19324, n19325, n19326, n19327, n19328,
    n19329, n19330, n19331, n19332, n19333, n19334,
    n19335, n19336, n19337, n19338, n19339, n19340,
    n19341, n19342, n19343, n19344, n19345, n19346,
    n19347, n19348, n19349, n19350, n19351, n19352,
    n19353, n19354, n19355, n19356, n19357, n19358,
    n19359, n19360, n19361, n19362, n19363, n19364,
    n19365, n19366, n19367, n19368, n19369, n19370,
    n19371, n19372, n19373, n19374, n19375, n19376,
    n19377, n19378, n19379, n19380, n19381, n19382,
    n19383, n19384, n19385, n19386, n19387, n19388,
    n19389, n19390, n19391, n19392, n19393, n19394,
    n19395, n19396, n19397, n19398, n19399, n19400,
    n19401, n19402, n19403, n19404, n19405, n19406,
    n19407, n19408, n19409, n19410, n19411, n19412,
    n19413, n19414, n19415, n19416, n19417, n19418,
    n19419, n19420, n19421, n19422, n19423, n19424,
    n19425, n19426, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19435, n19436,
    n19437, n19438, n19439, n19440, n19441, n19442,
    n19443, n19444, n19445, n19446, n19447, n19448,
    n19449, n19450, n19451, n19452, n19453, n19454,
    n19455, n19456, n19457, n19458, n19459, n19460,
    n19461, n19462, n19463, n19464, n19465, n19466,
    n19467, n19468, n19469, n19470, n19471, n19472,
    n19473, n19474, n19475, n19476, n19477, n19478,
    n19479, n19480, n19481, n19482, n19483, n19484,
    n19485, n19486, n19487, n19488, n19489, n19490,
    n19491, n19492, n19493, n19494, n19495, n19496,
    n19497, n19498, n19499, n19500, n19501, n19502,
    n19503, n19504, n19505, n19506, n19507, n19508,
    n19509, n19510, n19511, n19512, n19513, n19514,
    n19515, n19516, n19517, n19518, n19519, n19520,
    n19521, n19522, n19523, n19524, n19525, n19526,
    n19527, n19528, n19529, n19530, n19531, n19532,
    n19533, n19534, n19535, n19536, n19537, n19538,
    n19539, n19540, n19541, n19542, n19543, n19544,
    n19545, n19546, n19547, n19548, n19549, n19550,
    n19551, n19552, n19553, n19554, n19555, n19556,
    n19557, n19558, n19559, n19560, n19561, n19562,
    n19563, n19564, n19565, n19566, n19567, n19568,
    n19569, n19570, n19571, n19572, n19573, n19574,
    n19575, n19576, n19577, n19578, n19579, n19580,
    n19581, n19582, n19583, n19584, n19585, n19586,
    n19587, n19588, n19589, n19590, n19591, n19592,
    n19593, n19594, n19595, n19596, n19597, n19598,
    n19599, n19600, n19601, n19602, n19603, n19604,
    n19605, n19606, n19607, n19608, n19609, n19610,
    n19611, n19612, n19613, n19614, n19615, n19616,
    n19617, n19618, n19619, n19620, n19621, n19622,
    n19623, n19624, n19625, n19626, n19627, n19628,
    n19629, n19630, n19631, n19632, n19633, n19634,
    n19635, n19636, n19637, n19638, n19639, n19640,
    n19641, n19642, n19643, n19644, n19645, n19646,
    n19647, n19648, n19649, n19650, n19651, n19652,
    n19653, n19654, n19655, n19656, n19657, n19658,
    n19659, n19660, n19661, n19662, n19663, n19664,
    n19665, n19666, n19667, n19668, n19669, n19670,
    n19671, n19672, n19673, n19674, n19675, n19676,
    n19677, n19678, n19679, n19680, n19681, n19682,
    n19683, n19684, n19685, n19686, n19687, n19688,
    n19689, n19690, n19691, n19692, n19693, n19694,
    n19695, n19696, n19697, n19698, n19699, n19700,
    n19701, n19702, n19703, n19704, n19705, n19706,
    n19707, n19708, n19709, n19710, n19711, n19712,
    n19713, n19714, n19715, n19716, n19717, n19718,
    n19719, n19720, n19721, n19722, n19723, n19724,
    n19725, n19726, n19727, n19728, n19729, n19730,
    n19731, n19732, n19733, n19734, n19735, n19736,
    n19737, n19738, n19739, n19740, n19741, n19742,
    n19743, n19744, n19745, n19746, n19747, n19748,
    n19749, n19750, n19751, n19752, n19753, n19754,
    n19755, n19756, n19757, n19758, n19759, n19760,
    n19761, n19762, n19763, n19764, n19765, n19766,
    n19767, n19768, n19769, n19770, n19771, n19772,
    n19773, n19774, n19775, n19776, n19777, n19778,
    n19779, n19780, n19781, n19782, n19783, n19784,
    n19785, n19786, n19787, n19788, n19789, n19790,
    n19791, n19792, n19793, n19794, n19795, n19796,
    n19797, n19798, n19799, n19800, n19801, n19802,
    n19803, n19804, n19805, n19806, n19807, n19808,
    n19809, n19810, n19811, n19812, n19813, n19814,
    n19815, n19816, n19817, n19818, n19819, n19820,
    n19821, n19822, n19823, n19824, n19825, n19826,
    n19827, n19828, n19829, n19830, n19831, n19832,
    n19833, n19834, n19835, n19836, n19837, n19838,
    n19839, n19840, n19841, n19842, n19843, n19844,
    n19845, n19846, n19847, n19848, n19849, n19850,
    n19851, n19852, n19853, n19854, n19855, n19856,
    n19857, n19858, n19859, n19860, n19861, n19862,
    n19863, n19864, n19865, n19866, n19867, n19868,
    n19869, n19870, n19871, n19872, n19873, n19874,
    n19875, n19876, n19877, n19878, n19879, n19880,
    n19881, n19882, n19883, n19884, n19885, n19886,
    n19887, n19888, n19889, n19890, n19891, n19892,
    n19893, n19894, n19895, n19896, n19897, n19898,
    n19899, n19900, n19901, n19902, n19903, n19904,
    n19905, n19906, n19907, n19908, n19909, n19910,
    n19911, n19912, n19913, n19914, n19915, n19916,
    n19917, n19918, n19919, n19920, n19921, n19922,
    n19923, n19924, n19925, n19926, n19927, n19928,
    n19929, n19930, n19931, n19932, n19933, n19934,
    n19935, n19936, n19937, n19938, n19939, n19940,
    n19941, n19942, n19943, n19944, n19945, n19946,
    n19947, n19948, n19949, n19950, n19951, n19952,
    n19953, n19954, n19955, n19956, n19957, n19958,
    n19959, n19960, n19961, n19962, n19963, n19964,
    n19965, n19966, n19967, n19968, n19969, n19970,
    n19971, n19972, n19973, n19974, n19975, n19976,
    n19977, n19978, n19979, n19980, n19981, n19982,
    n19983, n19984, n19985, n19986, n19987, n19988,
    n19989, n19990, n19991, n19992, n19993, n19994,
    n19995, n19996, n19997, n19998, n19999, n20000,
    n20001, n20002, n20003, n20004, n20005, n20006,
    n20007, n20008, n20009, n20010, n20011, n20012,
    n20013, n20014, n20015, n20016, n20017, n20018,
    n20019, n20020, n20021, n20022, n20023, n20024,
    n20025, n20026, n20027, n20028, n20029, n20030,
    n20031, n20032, n20033, n20034, n20035, n20036,
    n20037, n20038, n20039, n20040, n20041, n20042,
    n20043, n20044, n20045, n20046, n20047, n20048,
    n20049, n20050, n20051, n20052, n20053, n20054,
    n20055, n20056, n20057, n20058, n20059, n20060,
    n20061, n20062, n20063, n20064, n20065, n20066,
    n20067, n20068, n20069, n20070, n20071, n20072,
    n20073, n20074, n20075, n20076, n20077, n20078,
    n20079, n20080, n20081, n20082, n20083, n20084,
    n20085, n20086, n20087, n20088, n20089, n20090,
    n20091, n20092, n20093, n20094, n20095, n20096,
    n20097, n20098, n20099, n20100, n20101, n20102,
    n20103, n20104, n20105, n20106, n20107, n20108,
    n20109, n20110, n20111, n20112, n20113, n20114,
    n20115, n20116, n20117, n20118, n20119, n20120,
    n20121, n20122, n20123, n20124, n20125, n20126,
    n20127, n20128, n20129, n20130, n20131, n20132,
    n20133, n20134, n20135, n20136, n20137, n20138,
    n20139, n20140, n20141, n20142, n20143, n20144,
    n20145, n20146, n20147, n20148, n20149, n20150,
    n20151, n20152, n20153, n20154, n20155, n20156,
    n20157, n20158, n20159, n20160, n20161, n20162,
    n20163, n20164, n20165, n20166, n20167, n20168,
    n20169, n20170, n20171, n20172, n20173, n20174,
    n20175, n20176, n20177, n20178, n20179, n20180,
    n20181, n20182, n20183, n20184, n20185, n20186,
    n20187, n20188, n20189, n20190, n20191, n20192,
    n20193, n20194, n20195, n20196, n20197, n20198,
    n20199, n20200, n20201, n20202, n20203, n20204,
    n20205, n20206, n20207, n20208, n20209, n20210,
    n20211, n20212, n20213, n20214, n20215, n20216,
    n20217, n20218, n20219, n20220, n20221, n20222,
    n20223, n20224, n20225, n20226, n20227, n20228,
    n20229, n20230, n20231, n20232, n20233, n20234,
    n20235, n20236, n20237, n20238, n20239, n20240,
    n20241, n20242, n20243, n20244, n20245, n20246,
    n20247, n20248, n20249, n20250, n20251, n20252,
    n20253, n20254, n20255, n20256, n20257, n20258,
    n20259, n20260, n20261, n20262, n20263, n20264,
    n20265, n20266, n20267, n20268, n20269, n20270,
    n20271, n20272, n20273, n20274, n20275, n20276,
    n20277, n20278, n20279, n20280, n20281, n20282,
    n20283, n20284, n20285, n20286, n20287, n20288,
    n20289, n20290, n20291, n20292, n20293, n20294,
    n20295, n20296, n20297, n20298, n20299, n20300,
    n20301, n20302, n20303, n20304, n20305, n20306,
    n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318,
    n20319, n20320, n20321, n20322, n20323, n20324,
    n20325, n20326, n20327, n20328, n20329, n20330,
    n20331, n20332, n20333, n20334, n20335, n20336,
    n20337, n20338, n20339, n20340, n20341, n20342,
    n20343, n20344, n20345, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354,
    n20355, n20356, n20357, n20358, n20359, n20360,
    n20361, n20362, n20363, n20364, n20365, n20366,
    n20367, n20368, n20369, n20370, n20371, n20372,
    n20373, n20374, n20375, n20376, n20377, n20378,
    n20379, n20380, n20381, n20382, n20383, n20384,
    n20385, n20386, n20387, n20388, n20389, n20390,
    n20391, n20392, n20393, n20394, n20395, n20396,
    n20397, n20398, n20399, n20400, n20401, n20402,
    n20403, n20404, n20405, n20406, n20407, n20408,
    n20409, n20410, n20411, n20412, n20413, n20414,
    n20415, n20416, n20417, n20418, n20419, n20420,
    n20421, n20422, n20423, n20424, n20425, n20426,
    n20427, n20428, n20429, n20430, n20431, n20432,
    n20433, n20434, n20435, n20436, n20437, n20438,
    n20439, n20440, n20441, n20442, n20443, n20444,
    n20445, n20446, n20447, n20448, n20449, n20450,
    n20451, n20452, n20453, n20454, n20455, n20456,
    n20457, n20458, n20459, n20460, n20461, n20462,
    n20463, n20464, n20465, n20466, n20467, n20468,
    n20469, n20470, n20471, n20472, n20473, n20474,
    n20475, n20476, n20477, n20478, n20479, n20480,
    n20481, n20482, n20483, n20484, n20485, n20486,
    n20487, n20488, n20489, n20490, n20491, n20492,
    n20493, n20494, n20495, n20496, n20497, n20498,
    n20499, n20500, n20501, n20502, n20503, n20504,
    n20505, n20506, n20507, n20508, n20509, n20510,
    n20511, n20512, n20513, n20514, n20515, n20516,
    n20517, n20518, n20519, n20520, n20521, n20522,
    n20523, n20524, n20525, n20526, n20527, n20528,
    n20529, n20530, n20531, n20532, n20533, n20534,
    n20535, n20536, n20537, n20538, n20539, n20540,
    n20541, n20542, n20543, n20544, n20545, n20546,
    n20547, n20548, n20549, n20550, n20551, n20552,
    n20553, n20554, n20555, n20556, n20557, n20558,
    n20559, n20560, n20561, n20562, n20563, n20564,
    n20565, n20566, n20567, n20568, n20569, n20570,
    n20571, n20572, n20573, n20574, n20575, n20576,
    n20577, n20578, n20579, n20580, n20581, n20582,
    n20583, n20584, n20585, n20586, n20587, n20588,
    n20589, n20590, n20591, n20592, n20593, n20594,
    n20595, n20596, n20597, n20598, n20599, n20600,
    n20601, n20602, n20603, n20604, n20605, n20606,
    n20607, n20608, n20609, n20610, n20611, n20612,
    n20613, n20614, n20615, n20616, n20617, n20618,
    n20619, n20620, n20621, n20622, n20623, n20624,
    n20625, n20626, n20627, n20628, n20629, n20630,
    n20631, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20645, n20646, n20647, n20648,
    n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660,
    n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20675, n20676, n20677, n20678,
    n20679, n20680, n20681, n20682, n20683, n20684,
    n20685, n20686, n20687, n20688, n20689, n20690,
    n20691, n20692, n20693, n20694, n20695, n20696,
    n20697, n20698, n20699, n20700, n20701, n20702,
    n20703, n20704, n20705, n20706, n20707, n20708,
    n20709, n20710, n20711, n20712, n20713, n20714,
    n20715, n20716, n20717, n20718, n20719, n20720,
    n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732,
    n20733, n20734, n20735, n20736, n20737, n20738,
    n20739, n20740, n20741, n20742, n20743, n20744,
    n20745, n20746, n20747, n20748, n20749, n20750,
    n20751, n20752, n20753, n20754, n20755, n20756,
    n20757, n20758, n20759, n20760, n20761, n20762,
    n20763, n20764, n20765, n20766, n20767, n20768,
    n20769, n20770, n20771, n20772, n20773, n20774,
    n20775, n20776, n20777, n20778, n20779, n20780,
    n20781, n20782, n20783, n20784, n20785, n20786,
    n20787, n20788, n20789, n20790, n20791, n20792,
    n20793, n20794, n20795, n20796, n20797, n20798,
    n20799, n20800, n20801, n20802, n20803, n20804,
    n20805, n20806, n20807, n20808, n20809, n20810,
    n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822,
    n20823, n20824, n20825, n20826, n20827, n20828,
    n20829, n20830, n20831, n20832, n20833, n20834,
    n20835, n20836, n20837, n20838, n20839, n20840,
    n20841, n20842, n20843, n20844, n20845, n20846,
    n20847, n20848, n20849, n20850, n20851, n20852,
    n20853, n20854, n20855, n20856, n20857, n20858,
    n20859, n20860, n20861, n20862, n20863, n20864,
    n20865, n20866, n20867, n20868, n20869, n20870,
    n20871, n20872, n20873, n20874, n20875, n20876,
    n20877, n20878, n20879, n20880, n20881, n20882,
    n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20892, n20893, n20894,
    n20895, n20896, n20897, n20898, n20899, n20900,
    n20901, n20902, n20903, n20904, n20905, n20906,
    n20907, n20908, n20909, n20910, n20911, n20912,
    n20913, n20914, n20915, n20916, n20917, n20918,
    n20919, n20920, n20921, n20922, n20923, n20924,
    n20925, n20926, n20927, n20928, n20929, n20930,
    n20931, n20932, n20933, n20934, n20935, n20936,
    n20937, n20938, n20939, n20940, n20941, n20942,
    n20943, n20944, n20945, n20946, n20947, n20948,
    n20949, n20950, n20951, n20952, n20953, n20954,
    n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972,
    n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984,
    n20985, n20986, n20987, n20988, n20989, n20990,
    n20991, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008,
    n21009, n21010, n21011, n21012, n21013, n21014,
    n21015, n21016, n21017, n21018, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026,
    n21027, n21028, n21029, n21030, n21031, n21032,
    n21033, n21034, n21035, n21036, n21037, n21038,
    n21039, n21040, n21041, n21042, n21043, n21044,
    n21045, n21046, n21047, n21048, n21049, n21050,
    n21051, n21052, n21053, n21054, n21055, n21056,
    n21057, n21058, n21059, n21060, n21061, n21062,
    n21063, n21064, n21065, n21066, n21067, n21068,
    n21069, n21070, n21071, n21072, n21073, n21074,
    n21075, n21076, n21077, n21078, n21079, n21080,
    n21081, n21082, n21083, n21084, n21085, n21086,
    n21087, n21088, n21089, n21090, n21091, n21092,
    n21093, n21094, n21095, n21096, n21097, n21098,
    n21099, n21100, n21101, n21102, n21103, n21104,
    n21105, n21106, n21107, n21108, n21109, n21110,
    n21111, n21112, n21113, n21114, n21115, n21116,
    n21117, n21118, n21119, n21120, n21121, n21122,
    n21123, n21124, n21125, n21126, n21127, n21128,
    n21129, n21130, n21131, n21132, n21133, n21134,
    n21135, n21136, n21137, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21145, n21146,
    n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158,
    n21159, n21160, n21161, n21162, n21163, n21164,
    n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176,
    n21177, n21178, n21179, n21180, n21181, n21182,
    n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200,
    n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218,
    n21219, n21220, n21221, n21222, n21223, n21224,
    n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236,
    n21237, n21238, n21239, n21240, n21241, n21242,
    n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260,
    n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21278,
    n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290,
    n21291, n21292, n21293, n21294, n21295, n21296,
    n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314,
    n21315, n21316, n21317, n21318, n21319, n21320,
    n21321, n21322, n21323, n21324, n21325, n21326,
    n21327, n21328, n21329, n21330, n21331, n21332,
    n21333, n21334, n21335, n21336, n21337, n21338,
    n21339, n21340, n21341, n21342, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350,
    n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368,
    n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428,
    n21429, n21430, n21431, n21432, n21433, n21434,
    n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21446,
    n21447, n21448, n21449, n21450, n21451, n21452,
    n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464,
    n21465, n21466, n21467, n21468, n21469, n21470,
    n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482,
    n21483, n21484, n21485, n21486, n21487, n21488,
    n21489, n21490, n21491, n21492, n21493, n21494,
    n21495, n21496, n21497, n21498, n21499, n21500,
    n21501, n21502, n21503, n21504, n21505, n21506,
    n21507, n21508, n21509, n21510, n21511, n21512,
    n21513, n21514, n21515, n21516, n21517, n21518,
    n21519, n21520, n21521, n21522, n21523, n21524,
    n21525, n21526, n21527, n21528, n21529, n21530,
    n21531, n21532, n21533, n21534, n21535, n21536,
    n21537, n21538, n21539, n21540, n21541, n21542,
    n21543, n21544, n21545, n21546, n21547, n21548,
    n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560,
    n21561, n21562, n21563, n21564, n21565, n21566,
    n21567, n21568, n21569, n21570, n21571, n21572,
    n21573, n21574, n21575, n21576, n21577, n21578,
    n21579, n21580, n21581, n21582, n21583, n21584,
    n21585, n21586, n21587, n21588, n21589, n21590,
    n21591, n21592, n21593, n21594, n21595, n21596,
    n21597, n21598, n21599, n21600, n21601, n21602,
    n21603, n21604, n21605, n21606, n21607, n21608,
    n21609, n21610, n21611, n21612, n21613, n21614,
    n21615, n21616, n21617, n21618, n21619, n21620,
    n21621, n21622, n21623, n21624, n21625, n21626,
    n21627, n21628, n21629, n21630, n21631, n21632,
    n21633, n21634, n21635, n21636, n21637, n21638,
    n21639, n21640, n21641, n21642, n21643, n21644,
    n21645, n21646, n21647, n21648, n21649, n21650,
    n21651, n21652, n21653, n21654, n21655, n21656,
    n21657, n21658, n21659, n21660, n21661, n21662,
    n21663, n21664, n21665, n21666, n21667, n21668,
    n21669, n21670, n21671, n21672, n21673, n21674,
    n21675, n21676, n21677, n21678, n21679, n21680,
    n21681, n21682, n21683, n21684, n21685, n21686,
    n21687, n21688, n21689, n21690, n21691, n21692,
    n21693, n21694, n21695, n21696, n21697, n21698,
    n21699, n21700, n21701, n21702, n21703, n21704,
    n21705, n21706, n21707, n21708, n21709, n21710,
    n21711, n21712, n21713, n21714, n21715, n21716,
    n21717, n21718, n21719, n21720, n21721, n21722,
    n21723, n21724, n21725, n21726, n21727, n21728,
    n21729, n21730, n21731, n21732, n21733, n21734,
    n21735, n21736, n21737, n21738, n21739, n21740,
    n21741, n21742, n21743, n21744, n21745, n21746,
    n21747, n21748, n21749, n21750, n21751, n21752,
    n21753, n21754, n21755, n21756, n21757, n21758,
    n21759, n21760, n21761, n21762, n21763, n21764,
    n21765, n21766, n21767, n21768, n21769, n21770,
    n21771, n21772, n21773, n21774, n21775, n21776,
    n21777, n21778, n21779, n21780, n21781, n21782,
    n21783, n21784, n21785, n21786, n21787, n21788,
    n21789, n21790, n21791, n21792, n21793, n21794,
    n21795, n21796, n21797, n21798, n21799, n21800,
    n21801, n21802, n21803, n21804, n21805, n21806,
    n21807, n21808, n21809, n21810, n21811, n21812,
    n21813, n21814, n21815, n21816, n21817, n21818,
    n21819, n21820, n21821, n21822, n21823, n21824,
    n21825, n21826, n21827, n21828, n21829, n21830,
    n21831, n21832, n21833, n21834, n21835, n21836,
    n21837, n21838, n21839, n21840, n21841, n21842,
    n21843, n21844, n21845, n21846, n21847, n21848,
    n21849, n21850, n21851, n21852, n21853, n21854,
    n21855, n21856, n21857, n21858, n21859, n21860,
    n21861, n21862, n21863, n21864, n21865, n21866,
    n21867, n21868, n21869, n21870, n21871, n21872,
    n21873, n21874, n21875, n21876, n21877, n21878,
    n21879, n21880, n21881, n21882, n21883, n21884,
    n21885, n21886, n21887, n21888, n21889, n21890,
    n21891, n21892, n21893, n21894, n21895, n21896,
    n21897, n21898, n21899, n21900, n21901, n21902,
    n21903, n21904, n21905, n21906, n21907, n21908,
    n21909, n21910, n21911, n21912, n21913, n21914,
    n21915, n21916, n21917, n21918, n21919, n21920,
    n21921, n21922, n21923, n21924, n21925, n21926,
    n21927, n21928, n21929, n21930, n21931, n21932,
    n21933, n21934, n21935, n21936, n21937, n21938,
    n21939, n21940, n21941, n21942, n21943, n21944,
    n21945, n21946, n21947, n21948, n21949, n21950,
    n21951, n21952, n21953, n21954, n21955, n21956,
    n21957, n21958, n21959, n21960, n21961, n21962,
    n21963, n21964, n21965, n21966, n21967, n21968,
    n21969, n21970, n21971, n21972, n21973, n21974,
    n21975, n21976, n21977, n21978, n21979, n21980,
    n21981, n21982, n21983, n21984, n21985, n21986,
    n21987, n21988, n21989, n21990, n21991, n21992,
    n21993, n21994, n21995, n21996, n21997, n21998,
    n21999, n22000, n22001, n22002, n22003, n22004,
    n22005, n22006, n22007, n22008, n22009, n22010,
    n22011, n22012, n22013, n22014, n22015, n22016,
    n22017, n22018, n22019, n22020, n22021, n22022,
    n22023, n22024, n22025, n22026, n22027, n22028,
    n22029, n22030, n22031, n22032, n22033, n22034,
    n22035, n22036, n22037, n22038, n22039, n22040,
    n22041, n22042, n22043, n22044, n22045, n22046,
    n22047, n22048, n22049, n22050, n22051, n22052,
    n22053, n22054, n22055, n22056, n22057, n22058,
    n22059, n22060, n22061, n22062, n22063, n22064,
    n22065, n22066, n22067, n22068, n22069, n22070,
    n22071, n22072, n22073, n22074, n22075, n22076,
    n22077, n22078, n22079, n22080, n22081, n22082,
    n22083, n22084, n22085, n22086, n22087, n22088,
    n22089, n22090, n22091, n22092, n22093, n22094,
    n22095, n22096, n22097, n22098, n22099, n22100,
    n22101, n22102, n22103, n22104, n22105, n22106,
    n22107, n22108, n22109, n22110, n22111, n22112,
    n22113, n22114, n22115, n22116, n22117, n22118,
    n22119, n22120, n22121, n22122, n22123, n22124,
    n22125, n22126, n22127, n22128, n22129, n22130,
    n22131, n22132, n22133, n22134, n22135, n22136,
    n22137, n22138, n22139, n22140, n22141, n22142,
    n22143, n22144, n22145, n22146, n22147, n22148,
    n22149, n22150, n22151, n22152, n22153, n22154,
    n22155, n22156, n22157, n22158, n22159, n22160,
    n22161, n22162, n22163, n22164, n22165, n22166,
    n22167, n22168, n22169, n22170, n22171, n22172,
    n22173, n22174, n22175, n22176, n22177, n22178,
    n22179, n22180, n22181, n22182, n22183, n22184,
    n22185, n22186, n22187, n22188, n22189, n22190,
    n22191, n22192, n22193, n22194, n22195, n22196,
    n22197, n22198, n22199, n22200, n22201, n22202,
    n22203, n22204, n22205, n22206, n22207, n22208,
    n22209, n22210, n22211, n22212, n22213, n22214,
    n22215, n22216, n22217, n22218, n22219, n22220,
    n22221, n22222, n22223, n22224, n22225, n22226,
    n22227, n22228, n22229, n22230, n22231, n22232,
    n22233, n22234, n22235, n22236, n22237, n22238,
    n22239, n22240, n22241, n22242, n22243, n22244,
    n22245, n22246, n22247, n22248, n22249, n22250,
    n22251, n22252, n22253, n22254, n22255, n22256,
    n22257, n22258, n22259, n22260, n22261, n22262,
    n22263, n22264, n22265, n22266, n22267, n22268,
    n22269, n22270, n22271, n22272, n22273, n22274,
    n22275, n22276, n22277, n22278, n22279, n22280,
    n22281, n22282, n22283, n22284, n22285, n22286,
    n22287, n22288, n22289, n22290, n22291, n22292,
    n22293, n22294, n22295, n22296, n22297, n22298,
    n22299, n22300, n22301, n22302, n22303, n22304,
    n22305, n22306, n22307, n22308, n22309, n22310,
    n22311, n22312, n22313, n22314, n22315, n22316,
    n22317, n22318, n22319, n22320, n22321, n22322,
    n22323, n22324, n22325, n22326, n22327, n22328,
    n22329, n22330, n22331, n22332, n22333, n22334,
    n22335, n22336, n22337, n22338, n22339, n22340,
    n22341, n22342, n22343, n22344, n22345, n22346,
    n22347, n22348, n22349, n22350, n22351, n22352,
    n22353, n22354, n22355, n22356, n22357, n22358,
    n22359, n22360, n22361, n22362, n22363, n22364,
    n22365, n22366, n22367, n22368, n22369, n22370,
    n22371, n22372, n22373, n22374, n22375, n22376,
    n22377, n22378, n22379, n22380, n22381, n22382,
    n22383, n22384, n22385, n22386, n22387, n22388,
    n22389, n22390, n22391, n22392, n22393, n22394,
    n22395, n22396, n22397, n22398, n22399, n22400,
    n22401, n22402, n22403, n22404, n22405, n22406,
    n22407, n22408, n22409, n22410, n22411, n22412,
    n22413, n22414, n22415, n22416, n22417, n22418,
    n22419, n22420, n22421, n22422, n22423, n22424,
    n22425, n22426, n22427, n22428, n22429, n22430,
    n22431, n22432, n22433, n22434, n22435, n22436,
    n22437, n22438, n22439, n22440, n22441, n22442,
    n22443, n22444, n22445, n22446, n22447, n22448,
    n22449, n22450, n22451, n22452, n22453, n22454,
    n22455, n22456, n22457, n22458, n22459, n22460,
    n22461, n22462, n22463, n22464, n22465, n22466,
    n22467, n22468, n22469, n22470, n22471, n22472,
    n22473, n22474, n22475, n22476, n22477, n22478,
    n22479, n22480, n22481, n22482, n22483, n22484,
    n22485, n22486, n22487, n22488, n22489, n22490,
    n22491, n22492, n22493, n22494, n22495, n22496,
    n22497, n22498, n22499, n22500, n22501, n22502,
    n22503, n22504, n22505, n22506, n22507, n22508,
    n22509, n22510, n22511, n22512, n22513, n22514,
    n22515, n22516, n22517, n22518, n22519, n22520,
    n22521, n22522, n22523, n22524, n22525, n22526,
    n22527, n22528, n22529, n22530, n22531, n22532,
    n22533, n22534, n22535, n22536, n22537, n22538,
    n22539, n22540, n22541, n22542, n22543, n22544,
    n22545, n22546, n22547, n22548, n22549, n22550,
    n22551, n22552, n22553, n22554, n22555, n22556,
    n22557, n22558, n22559, n22560, n22561, n22562,
    n22563, n22564, n22565, n22566, n22567, n22568,
    n22569, n22570, n22571, n22572, n22573, n22574,
    n22575, n22576, n22577, n22578, n22579, n22580,
    n22581, n22582, n22583, n22584, n22585, n22586,
    n22587, n22588, n22589, n22590, n22591, n22592,
    n22593, n22594, n22595, n22596, n22597, n22598,
    n22599, n22600, n22601, n22602, n22603, n22604,
    n22605, n22606, n22607, n22608, n22609, n22610,
    n22611, n22612, n22613, n22614, n22615, n22616,
    n22617, n22618, n22619, n22620, n22621, n22622,
    n22623, n22624, n22625, n22626, n22627, n22628,
    n22629, n22630, n22631, n22632, n22633, n22634,
    n22635, n22636, n22637, n22638, n22639, n22640,
    n22641, n22642, n22643, n22644, n22645, n22646,
    n22647, n22648, n22649, n22650, n22651, n22652,
    n22653, n22654, n22655, n22656, n22657, n22658,
    n22659, n22660, n22661, n22662, n22663, n22664,
    n22665, n22666, n22667, n22668, n22669, n22670,
    n22671, n22672, n22673, n22674, n22675, n22676,
    n22677, n22678, n22679, n22680, n22681, n22682,
    n22683, n22684, n22685, n22686, n22687, n22688,
    n22689, n22690, n22691, n22692, n22693, n22694,
    n22695, n22696, n22697, n22698, n22699, n22700,
    n22701, n22702, n22703, n22704, n22705, n22706,
    n22707, n22708, n22709, n22710, n22711, n22712,
    n22713, n22714, n22715, n22716, n22717, n22718,
    n22719, n22720, n22721, n22722, n22723, n22724,
    n22725, n22726, n22727, n22728, n22729, n22730,
    n22731, n22732, n22733, n22734, n22735, n22736,
    n22737, n22738, n22739, n22740, n22741, n22742,
    n22743, n22744, n22745, n22746, n22747, n22748,
    n22749, n22750, n22751, n22752, n22753, n22754,
    n22755, n22756, n22757, n22758, n22759, n22760,
    n22761, n22762, n22763, n22764, n22765, n22766,
    n22767, n22768, n22769, n22770, n22771, n22772,
    n22773, n22774, n22775, n22776, n22777, n22778,
    n22779, n22780, n22781, n22782, n22783, n22784,
    n22785, n22786, n22787, n22788, n22789, n22790,
    n22791, n22792, n22793, n22794, n22795, n22796,
    n22797, n22798, n22799, n22800, n22801, n22802,
    n22803, n22804, n22805, n22806, n22807, n22808,
    n22809, n22810, n22811, n22812, n22813, n22814,
    n22815, n22816, n22817, n22818, n22819, n22820,
    n22821, n22822, n22823, n22824, n22825, n22826,
    n22827, n22828, n22829, n22830, n22831, n22832,
    n22833, n22834, n22835, n22836, n22837, n22838,
    n22839, n22840, n22841, n22842, n22843, n22844,
    n22845, n22846, n22847, n22848, n22849, n22850,
    n22851, n22852, n22853, n22854, n22855, n22856,
    n22857, n22858, n22859, n22860, n22861, n22862,
    n22863, n22864, n22865, n22866, n22867, n22868,
    n22869, n22870, n22871, n22872, n22873, n22874,
    n22875, n22876, n22877, n22878, n22879, n22880,
    n22881, n22882, n22883, n22884, n22885, n22886,
    n22887, n22888, n22889, n22890, n22891, n22892,
    n22893, n22894, n22895, n22896, n22897, n22898,
    n22899, n22900, n22901, n22902, n22903, n22904,
    n22905, n22906, n22907, n22908, n22909, n22910,
    n22911, n22912, n22913, n22914, n22915, n22916,
    n22917, n22918, n22919, n22920, n22921, n22922,
    n22923, n22924, n22925, n22926, n22927, n22928,
    n22929, n22930, n22931, n22932, n22933, n22934,
    n22935, n22936, n22937, n22938, n22939, n22940,
    n22941, n22942, n22943, n22944, n22945, n22946,
    n22947, n22948, n22949, n22950, n22951, n22952,
    n22953, n22954, n22955, n22956, n22957, n22958,
    n22959, n22960, n22961, n22962, n22963, n22964,
    n22965, n22966, n22967, n22968, n22969, n22970,
    n22971, n22972, n22973, n22974, n22975, n22976,
    n22977, n22978, n22979, n22980, n22981, n22982,
    n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994,
    n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012,
    n23013, n23014, n23015, n23016, n23017, n23018,
    n23019, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n23028, n23029, n23030,
    n23031, n23032, n23033, n23034, n23035, n23036,
    n23037, n23038, n23039, n23040, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048,
    n23049, n23050, n23051, n23052, n23053, n23054,
    n23055, n23056, n23057, n23058, n23059, n23060,
    n23061, n23062, n23063, n23064, n23065, n23066,
    n23067, n23068, n23069, n23070, n23071, n23072,
    n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084,
    n23085, n23086, n23087, n23088, n23089, n23090,
    n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102,
    n23103, n23104, n23105, n23106, n23107, n23108,
    n23109, n23110, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120,
    n23121, n23122, n23123, n23124, n23125, n23126,
    n23127, n23128, n23129, n23130, n23131, n23132,
    n23133, n23134, n23135, n23136, n23137, n23138,
    n23139, n23140, n23141, n23142, n23143, n23144,
    n23145, n23146, n23147, n23148, n23149, n23150,
    n23151, n23152, n23153, n23154, n23155, n23156,
    n23157, n23158, n23159, n23160, n23161, n23162,
    n23163, n23164, n23165, n23166, n23167, n23168,
    n23169, n23170, n23171, n23172, n23173, n23174,
    n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186,
    n23187, n23188, n23189, n23190, n23191, n23192,
    n23193, n23194, n23195, n23196, n23197, n23198,
    n23199, n23200, n23201, n23202, n23203, n23204,
    n23205, n23206, n23207, n23208, n23209, n23210,
    n23211, n23212, n23213, n23214, n23215, n23216,
    n23217, n23218, n23219, n23220, n23221, n23222,
    n23223, n23224, n23225, n23226, n23227, n23228,
    n23229, n23230, n23231, n23232, n23233, n23234,
    n23235, n23236, n23237, n23238, n23239, n23240,
    n23241, n23242, n23243, n23244, n23245, n23246,
    n23247, n23248, n23249, n23250, n23251, n23252,
    n23253, n23254, n23255, n23256, n23257, n23258,
    n23259, n23260, n23261, n23262, n23263, n23264,
    n23265, n23266, n23267, n23268, n23269, n23270,
    n23271, n23272, n23273, n23274, n23275, n23276,
    n23277, n23278, n23279, n23280, n23281, n23282,
    n23283, n23284, n23285, n23286, n23287, n23288,
    n23289, n23290, n23291, n23292, n23293, n23294,
    n23295, n23296, n23297, n23298, n23299, n23300,
    n23301, n23302, n23303, n23304, n23305, n23306,
    n23307, n23308, n23309, n23310, n23311, n23312,
    n23313, n23314, n23315, n23316, n23317, n23318,
    n23319, n23320, n23321, n23322, n23323, n23324,
    n23325, n23326, n23327, n23328, n23329, n23330,
    n23331, n23332, n23333, n23334, n23335, n23336,
    n23337, n23338, n23339, n23340, n23341, n23342,
    n23343, n23344, n23345, n23346, n23347, n23348,
    n23349, n23350, n23351, n23352, n23353, n23354,
    n23355, n23356, n23357, n23358, n23359, n23360,
    n23361, n23362, n23363, n23364, n23365, n23366,
    n23367, n23368, n23369, n23370, n23371, n23372,
    n23373, n23374, n23375, n23376, n23377, n23378,
    n23379, n23380, n23381, n23382, n23383, n23384,
    n23385, n23386, n23387, n23388, n23389, n23390,
    n23391, n23392, n23393, n23394, n23395, n23396,
    n23397, n23398, n23399, n23400, n23401, n23402,
    n23403, n23404, n23405, n23406, n23407, n23408,
    n23409, n23410, n23411, n23412, n23413, n23414,
    n23415, n23416, n23417, n23418, n23419, n23420,
    n23421, n23422, n23423, n23424, n23425, n23426,
    n23427, n23428, n23429, n23430, n23431, n23432,
    n23433, n23434, n23435, n23436, n23437, n23438,
    n23439, n23440, n23441, n23442, n23443, n23444,
    n23445, n23446, n23447, n23448, n23449, n23450,
    n23451, n23452, n23453, n23454, n23455, n23456,
    n23457, n23458, n23459, n23460, n23461, n23462,
    n23463, n23464, n23465, n23466, n23467, n23468,
    n23469, n23470, n23471, n23472, n23473, n23474,
    n23475, n23476, n23477, n23478, n23479, n23480,
    n23481, n23482, n23483, n23484, n23485, n23486,
    n23487, n23488, n23489, n23490, n23491, n23492,
    n23493, n23494, n23495, n23496, n23497, n23498,
    n23499, n23500, n23501, n23502, n23503, n23504,
    n23505, n23506, n23507, n23508, n23509, n23510,
    n23511, n23512, n23513, n23514, n23515, n23516,
    n23517, n23518, n23519, n23520, n23521, n23522,
    n23523, n23524, n23525, n23526, n23527, n23528,
    n23529, n23530, n23531, n23532, n23533, n23534,
    n23535, n23536, n23537, n23538, n23539, n23540,
    n23541, n23542, n23543, n23544, n23545, n23546,
    n23547, n23548, n23549, n23550, n23551, n23552,
    n23553, n23554, n23555, n23556, n23557, n23558,
    n23559, n23560, n23561, n23562, n23563, n23564,
    n23565, n23566, n23567, n23568, n23569, n23570,
    n23571, n23572, n23573, n23574, n23575, n23576,
    n23577, n23578, n23579, n23580, n23581, n23582,
    n23583, n23584, n23585, n23586, n23587, n23588,
    n23589, n23590, n23591, n23592, n23593, n23594,
    n23595, n23596, n23597, n23598, n23599, n23600,
    n23601, n23602, n23603, n23604, n23605, n23606,
    n23607, n23608, n23609, n23610, n23611, n23612,
    n23613, n23614, n23615, n23616, n23617, n23618,
    n23619, n23620, n23621, n23622, n23623, n23624,
    n23625, n23626, n23627, n23628, n23629, n23630,
    n23631, n23632, n23633, n23634, n23635, n23636,
    n23637, n23638, n23639, n23640, n23641, n23642,
    n23643, n23644, n23645, n23646, n23647, n23648,
    n23649, n23650, n23651, n23652, n23653, n23654,
    n23655, n23656, n23657, n23658, n23659, n23660,
    n23661, n23662, n23663, n23664, n23665, n23666,
    n23667, n23668, n23669, n23670, n23671, n23672,
    n23673, n23674, n23675, n23676, n23677, n23678,
    n23679, n23680, n23681, n23682, n23683, n23684,
    n23685, n23686, n23687, n23688, n23689, n23690,
    n23691, n23692, n23693, n23694, n23695, n23696,
    n23697, n23698, n23699, n23700, n23701, n23702,
    n23703, n23704, n23705, n23706, n23707, n23708,
    n23709, n23710, n23711, n23712, n23713, n23714,
    n23715, n23716, n23717, n23718, n23719, n23720,
    n23721, n23722, n23723, n23724, n23725, n23726,
    n23727, n23728, n23729, n23730, n23731, n23732,
    n23733, n23734, n23735, n23736, n23737, n23738,
    n23739, n23740, n23741, n23742, n23743, n23744,
    n23745, n23746, n23747, n23748, n23749, n23750,
    n23751, n23752, n23753, n23754, n23755, n23756,
    n23757, n23758, n23759, n23760, n23761, n23762,
    n23763, n23764, n23765, n23766, n23767, n23768,
    n23769, n23770, n23771, n23772, n23773, n23774,
    n23775, n23776, n23777, n23778, n23779, n23780,
    n23781, n23782, n23783, n23784, n23785, n23786,
    n23787, n23788, n23789, n23790, n23791, n23792,
    n23793, n23794, n23795, n23796, n23797, n23798,
    n23799, n23800, n23801, n23802, n23803, n23804,
    n23805, n23806, n23807, n23808, n23809, n23810,
    n23811, n23812, n23813, n23814, n23815, n23816,
    n23817, n23818, n23819, n23820, n23821, n23822,
    n23823, n23824, n23825, n23826, n23827, n23828,
    n23829, n23830, n23831, n23832, n23833, n23834,
    n23835, n23836, n23837, n23838, n23839, n23840,
    n23841, n23842, n23843, n23844, n23845, n23846,
    n23847, n23848, n23849, n23850, n23851, n23852,
    n23853, n23854, n23855, n23856, n23857, n23858,
    n23859, n23860, n23861, n23862, n23863, n23864,
    n23865, n23866, n23867, n23868, n23869, n23870,
    n23871, n23872, n23873, n23874, n23875, n23876,
    n23877, n23878, n23879, n23880, n23881, n23882,
    n23883, n23884, n23885, n23886, n23887, n23888,
    n23889, n23890, n23891, n23892, n23893, n23894,
    n23895, n23896, n23897, n23898, n23899, n23900,
    n23901, n23902, n23903, n23904, n23905, n23906,
    n23907, n23908, n23909, n23910, n23911, n23912,
    n23913, n23914, n23915, n23916, n23917, n23918,
    n23919, n23920, n23921, n23922, n23923, n23924,
    n23925, n23926, n23927, n23928, n23929, n23930,
    n23931, n23932, n23933, n23934, n23935, n23936,
    n23937, n23938, n23939, n23940, n23941, n23942,
    n23943, n23944, n23945, n23946, n23947, n23948,
    n23949, n23950, n23951, n23952, n23953, n23954,
    n23955, n23956, n23957, n23958, n23959, n23960,
    n23961, n23962, n23963, n23964, n23965, n23966,
    n23967, n23968, n23969, n23970, n23971, n23972,
    n23973, n23974, n23975, n23976, n23977, n23978,
    n23979, n23980, n23981, n23982, n23983, n23984,
    n23985, n23986, n23987, n23988, n23989, n23990,
    n23991, n23992, n23993, n23994, n23995, n23996,
    n23997, n23998, n23999, n24000, n24001, n24002,
    n24003, n24004, n24005, n24006, n24007, n24008,
    n24009, n24010, n24011, n24012, n24013, n24014,
    n24015, n24016, n24017, n24018, n24019, n24020,
    n24021, n24022, n24023, n24024, n24025, n24026,
    n24027, n24028, n24029, n24030, n24031, n24032,
    n24033, n24034, n24035, n24036, n24037, n24038,
    n24039, n24040, n24041, n24042, n24043, n24044,
    n24045, n24046, n24047, n24048, n24049, n24050,
    n24051, n24052, n24053, n24054, n24055, n24056,
    n24057, n24058, n24059, n24060, n24061, n24062,
    n24063, n24064, n24065, n24066, n24067, n24068,
    n24069, n24070, n24071, n24072, n24073, n24074,
    n24075, n24076, n24077, n24078, n24079, n24080,
    n24081, n24082, n24083, n24084, n24085, n24086,
    n24087, n24088, n24089, n24090, n24091, n24092,
    n24093, n24094, n24095, n24096, n24097, n24098,
    n24099, n24100, n24101, n24102, n24103, n24104,
    n24105, n24106, n24107, n24108, n24109, n24110,
    n24111, n24112, n24113, n24114, n24115, n24116,
    n24117, n24118, n24119, n24120, n24121, n24122,
    n24123, n24124, n24125, n24126, n24127, n24128,
    n24129, n24130, n24131, n24132, n24133, n24134,
    n24135, n24136, n24137, n24138, n24139, n24140,
    n24141, n24142, n24143, n24144, n24145, n24146,
    n24147, n24148, n24149, n24150, n24151, n24152,
    n24153, n24154, n24155, n24156, n24157, n24158,
    n24159, n24160, n24161, n24162, n24163, n24164,
    n24165, n24166, n24167, n24168, n24169, n24170,
    n24171, n24172, n24173, n24174, n24175, n24176,
    n24177, n24178, n24179, n24180, n24181, n24182,
    n24183, n24184, n24185, n24186, n24187, n24188,
    n24189, n24190, n24191, n24192, n24193, n24194,
    n24195, n24196, n24197, n24198, n24199, n24200,
    n24201, n24202, n24203, n24204, n24205, n24206,
    n24207, n24208, n24209, n24210, n24211, n24212,
    n24213, n24214, n24215, n24216, n24217, n24218,
    n24219, n24220, n24221, n24222, n24223, n24224,
    n24225, n24226, n24227, n24228, n24229, n24230,
    n24231, n24232, n24233, n24234, n24235, n24236,
    n24237, n24238, n24239, n24240, n24241, n24242,
    n24243, n24244, n24245, n24246, n24247, n24248,
    n24249, n24250, n24251, n24252, n24253, n24254,
    n24255, n24256, n24257, n24258, n24259, n24260,
    n24261, n24262, n24263, n24264, n24265, n24266,
    n24267, n24268, n24269, n24270, n24271, n24272,
    n24273, n24274, n24275, n24276, n24277, n24278,
    n24279, n24280, n24281, n24282, n24283, n24284,
    n24285, n24286, n24287, n24288, n24289, n24290,
    n24291, n24292, n24293, n24294, n24295, n24296,
    n24297, n24298, n24299, n24300, n24301, n24302,
    n24303, n24304, n24305, n24306, n24307, n24308,
    n24309, n24310, n24311, n24312, n24313, n24314,
    n24315, n24316, n24317, n24318, n24319, n24320,
    n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332,
    n24333, n24334, n24335, n24336, n24337, n24338,
    n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350,
    n24351, n24352, n24353, n24354, n24355, n24356,
    n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368,
    n24369, n24370, n24371, n24372, n24373, n24374,
    n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386,
    n24387, n24388, n24389, n24390, n24391, n24392,
    n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404,
    n24405, n24406, n24407, n24408, n24409, n24410,
    n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422,
    n24423, n24424, n24425, n24426, n24427, n24428,
    n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440,
    n24441, n24442, n24443, n24444, n24445, n24446,
    n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24458,
    n24459, n24460, n24461, n24462, n24463, n24464,
    n24465, n24466, n24467, n24468, n24469, n24470,
    n24471, n24472, n24473, n24474, n24475, n24476,
    n24477, n24478, n24479, n24480, n24481, n24482,
    n24483, n24484, n24485, n24486, n24487, n24488,
    n24489, n24490, n24491, n24492, n24493, n24494,
    n24495, n24496, n24497, n24498, n24499, n24500,
    n24501, n24502, n24503, n24504, n24505, n24506,
    n24507, n24508, n24509, n24510, n24511, n24512,
    n24513, n24514, n24515, n24516, n24517, n24518,
    n24519, n24520, n24521, n24522, n24523, n24524,
    n24525, n24526, n24527, n24528, n24529, n24530,
    n24531, n24532, n24533, n24534, n24535, n24536,
    n24537, n24538, n24539, n24540, n24541, n24542,
    n24543, n24544, n24545, n24546, n24547, n24548,
    n24549, n24550, n24551, n24552, n24553, n24554,
    n24555, n24556, n24558, n24559, n24560, n24561,
    n24562, n24563, n24564, n24565, n24566, n24567,
    n24568, n24569, n24570, n24571, n24572, n24573,
    n24574, n24575, n24576, n24577, n24578, n24579,
    n24580, n24581, n24582, n24583, n24584, n24585,
    n24586, n24587, n24588, n24589, n24590, n24591,
    n24592, n24593, n24594, n24595, n24596, n24597,
    n24598, n24599, n24600, n24601, n24602, n24603,
    n24604, n24605, n24606, n24607, n24608, n24609,
    n24610, n24611, n24612, n24613, n24614, n24615,
    n24616, n24617, n24618, n24619, n24620, n24621,
    n24622, n24623, n24624, n24625, n24626, n24627,
    n24628, n24629, n24630, n24631, n24632, n24633,
    n24634, n24635, n24636, n24637, n24638, n24639,
    n24640, n24641, n24642, n24643, n24644, n24645,
    n24646, n24647, n24648, n24649, n24650, n24651,
    n24652, n24653, n24654, n24655, n24656, n24657,
    n24658, n24659, n24660, n24661, n24662, n24663,
    n24664, n24665, n24666, n24667, n24668, n24669,
    n24670, n24671, n24672, n24673, n24674, n24675,
    n24676, n24677, n24678, n24679, n24680, n24681,
    n24682, n24683, n24684, n24685, n24686, n24687,
    n24688, n24689, n24690, n24691, n24692, n24693,
    n24694, n24695, n24696, n24697, n24698, n24699,
    n24700, n24701, n24702, n24703, n24704, n24705,
    n24706, n24707, n24708, n24709, n24710, n24711,
    n24712, n24713, n24714, n24715, n24716, n24717,
    n24718, n24719, n24720, n24721, n24722, n24723,
    n24724, n24725, n24726, n24727, n24728, n24729,
    n24730, n24731, n24732, n24733, n24734, n24735,
    n24736, n24737, n24738, n24739, n24740, n24741,
    n24742, n24743, n24744, n24745, n24746, n24747,
    n24748, n24749, n24750, n24751, n24752, n24753,
    n24754, n24755, n24756, n24757, n24758, n24759,
    n24760, n24761, n24762, n24763, n24764, n24765,
    n24766, n24767, n24768, n24769, n24770, n24771,
    n24772, n24773, n24774, n24775, n24776, n24777,
    n24778, n24779, n24780, n24781, n24782, n24783,
    n24784, n24785, n24786, n24787, n24788, n24789,
    n24790, n24791, n24792, n24793, n24794, n24795,
    n24796, n24797, n24798, n24799, n24800, n24801,
    n24802, n24803, n24804, n24806, n24807, n24808,
    n24809, n24810, n24811, n24812, n24813, n24814,
    n24815, n24816, n24817, n24818, n24819, n24820,
    n24821, n24822, n24823, n24824, n24825, n24826,
    n24827, n24828, n24829, n24830, n24831, n24832,
    n24833, n24834, n24835, n24836, n24837, n24838,
    n24839, n24840, n24841, n24842, n24843, n24844,
    n24845, n24846, n24847, n24848, n24849, n24850,
    n24851, n24852, n24853, n24854, n24855, n24856,
    n24857, n24858, n24859, n24860, n24861, n24862,
    n24863, n24864, n24865, n24866, n24867, n24868,
    n24869, n24870, n24871, n24872, n24873, n24874,
    n24875, n24876, n24877, n24878, n24879, n24880,
    n24881, n24882, n24883, n24884, n24885, n24886,
    n24887, n24888, n24889, n24890, n24891, n24892,
    n24893, n24894, n24895, n24896, n24897, n24898,
    n24899, n24900, n24901, n24902, n24903, n24904,
    n24905, n24906, n24907, n24908, n24909, n24910,
    n24911, n24912, n24913, n24914, n24915, n24916,
    n24917, n24918, n24919, n24920, n24921, n24922,
    n24923, n24924, n24925, n24926, n24927, n24928,
    n24929, n24930, n24931, n24932, n24933, n24934,
    n24935, n24936, n24937, n24938, n24939, n24940,
    n24941, n24942, n24943, n24944, n24945, n24946,
    n24947, n24948, n24949, n24950, n24951, n24952,
    n24953, n24954, n24955, n24956, n24957, n24958,
    n24959, n24960, n24961, n24962, n24963, n24964,
    n24965, n24966, n24967, n24968, n24969, n24970,
    n24971, n24972, n24973, n24974, n24975, n24976,
    n24977, n24978, n24979, n24980, n24981, n24982,
    n24983, n24984, n24985, n24986, n24987, n24988,
    n24989, n24990, n24991, n24992, n24993, n24994,
    n24995, n24996, n24997, n24998, n24999, n25000,
    n25001, n25002, n25003, n25004, n25005, n25006,
    n25007, n25008, n25009, n25010, n25011, n25012,
    n25013, n25014, n25015, n25016, n25017, n25018,
    n25019, n25020, n25021, n25022, n25023, n25024,
    n25025, n25026, n25027, n25028, n25029, n25030,
    n25031, n25032, n25033, n25034, n25035, n25036,
    n25037, n25038, n25039, n25040, n25041, n25042,
    n25043, n25044, n25045, n25046, n25047, n25049,
    n25050, n25051, n25052, n25053, n25054, n25055,
    n25056, n25057, n25058, n25059, n25060, n25061,
    n25062, n25063, n25064, n25065, n25066, n25067,
    n25068, n25069, n25070, n25071, n25072, n25073,
    n25074, n25075, n25076, n25077, n25078, n25079,
    n25080, n25081, n25082, n25083, n25084, n25085,
    n25086, n25087, n25088, n25089, n25090, n25091,
    n25092, n25093, n25094, n25095, n25096, n25097,
    n25098, n25099, n25100, n25101, n25102, n25103,
    n25104, n25105, n25106, n25107, n25108, n25109,
    n25110, n25111, n25112, n25113, n25114, n25115,
    n25116, n25117, n25118, n25119, n25120, n25121,
    n25122, n25123, n25124, n25125, n25126, n25127,
    n25128, n25129, n25130, n25131, n25132, n25133,
    n25134, n25135, n25136, n25137, n25138, n25139,
    n25140, n25141, n25142, n25143, n25144, n25145,
    n25146, n25147, n25148, n25149, n25150, n25151,
    n25152, n25153, n25154, n25155, n25156, n25157,
    n25158, n25159, n25160, n25161, n25162, n25163,
    n25164, n25165, n25166, n25167, n25168, n25169,
    n25170, n25171, n25172, n25173, n25174, n25175,
    n25176, n25177, n25178, n25179, n25180, n25181,
    n25182, n25183, n25184, n25185, n25186, n25187,
    n25188, n25189, n25190, n25191, n25192, n25193,
    n25194, n25195, n25196, n25197, n25198, n25199,
    n25200, n25201, n25202, n25203, n25204, n25205,
    n25206, n25207, n25208, n25209, n25210, n25211,
    n25212, n25213, n25214, n25215, n25216, n25217,
    n25218, n25219, n25220, n25221, n25222, n25223,
    n25224, n25225, n25226, n25227, n25228, n25229,
    n25230, n25231, n25232, n25233, n25234, n25235,
    n25236, n25237, n25238, n25239, n25240, n25241,
    n25242, n25243, n25244, n25245, n25246, n25247,
    n25248, n25249, n25250, n25251, n25252, n25253,
    n25254, n25255, n25256, n25257, n25258, n25259,
    n25260, n25261, n25262, n25263, n25264, n25265,
    n25266, n25267, n25268, n25269, n25270, n25271,
    n25272, n25273, n25274, n25275, n25276, n25277,
    n25278, n25280, n25281, n25282, n25283, n25284,
    n25285, n25286, n25287, n25288, n25289, n25290,
    n25291, n25292, n25293, n25294, n25295, n25296,
    n25297, n25298, n25299, n25300, n25301, n25302,
    n25303, n25304, n25305, n25306, n25307, n25308,
    n25309, n25310, n25311, n25312, n25313, n25314,
    n25315, n25316, n25317, n25318, n25319, n25320,
    n25321, n25322, n25323, n25324, n25325, n25326,
    n25327, n25328, n25329, n25330, n25331, n25332,
    n25333, n25334, n25335, n25336, n25337, n25338,
    n25339, n25340, n25341, n25342, n25343, n25344,
    n25345, n25346, n25347, n25348, n25349, n25350,
    n25351, n25352, n25353, n25354, n25355, n25356,
    n25357, n25358, n25359, n25360, n25361, n25362,
    n25363, n25364, n25365, n25366, n25367, n25368,
    n25369, n25370, n25371, n25372, n25373, n25374,
    n25375, n25376, n25377, n25378, n25379, n25380,
    n25381, n25382, n25383, n25384, n25385, n25386,
    n25387, n25388, n25389, n25390, n25391, n25392,
    n25393, n25394, n25395, n25396, n25397, n25398,
    n25399, n25400, n25401, n25402, n25403, n25404,
    n25405, n25406, n25407, n25408, n25409, n25410,
    n25411, n25412, n25413, n25414, n25415, n25416,
    n25417, n25418, n25419, n25420, n25421, n25422,
    n25423, n25424, n25425, n25426, n25427, n25428,
    n25429, n25430, n25431, n25432, n25433, n25434,
    n25435, n25436, n25437, n25438, n25439, n25440,
    n25441, n25442, n25443, n25444, n25445, n25446,
    n25447, n25448, n25449, n25450, n25451, n25452,
    n25453, n25454, n25455, n25456, n25457, n25458,
    n25459, n25460, n25461, n25462, n25463, n25464,
    n25465, n25466, n25467, n25468, n25469, n25470,
    n25471, n25472, n25473, n25474, n25475, n25476,
    n25477, n25478, n25479, n25480, n25481, n25482,
    n25483, n25484, n25485, n25486, n25487, n25488,
    n25489, n25490, n25491, n25492, n25493, n25494,
    n25495, n25496, n25497, n25498, n25499, n25500,
    n25501, n25502, n25503, n25504, n25505, n25506,
    n25507, n25508, n25509, n25510, n25511, n25512,
    n25513, n25514, n25515, n25517, n25518, n25519,
    n25520, n25521, n25522, n25523, n25524, n25525,
    n25526, n25527, n25528, n25529, n25530, n25531,
    n25532, n25533, n25534, n25535, n25536, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543,
    n25544, n25545, n25546, n25547, n25548, n25549,
    n25550, n25551, n25552, n25553, n25554, n25555,
    n25556, n25557, n25558, n25559, n25560, n25561,
    n25562, n25563, n25564, n25565, n25566, n25567,
    n25568, n25569, n25570, n25571, n25572, n25573,
    n25574, n25575, n25576, n25577, n25578, n25579,
    n25580, n25581, n25582, n25583, n25584, n25585,
    n25586, n25587, n25588, n25589, n25590, n25591,
    n25592, n25593, n25594, n25595, n25596, n25597,
    n25598, n25599, n25600, n25601, n25602, n25603,
    n25604, n25605, n25606, n25607, n25608, n25609,
    n25610, n25611, n25612, n25613, n25614, n25615,
    n25616, n25617, n25618, n25619, n25620, n25621,
    n25622, n25623, n25624, n25625, n25626, n25627,
    n25628, n25629, n25630, n25631, n25632, n25633,
    n25634, n25635, n25636, n25637, n25638, n25639,
    n25640, n25641, n25642, n25643, n25644, n25645,
    n25646, n25647, n25648, n25649, n25650, n25651,
    n25652, n25653, n25654, n25655, n25656, n25657,
    n25658, n25659, n25660, n25661, n25662, n25663,
    n25664, n25665, n25666, n25667, n25668, n25669,
    n25670, n25671, n25672, n25673, n25674, n25675,
    n25676, n25677, n25678, n25679, n25680, n25681,
    n25682, n25683, n25684, n25685, n25686, n25687,
    n25688, n25689, n25690, n25691, n25692, n25693,
    n25694, n25695, n25696, n25697, n25698, n25699,
    n25700, n25701, n25702, n25703, n25704, n25705,
    n25706, n25707, n25708, n25709, n25710, n25711,
    n25712, n25713, n25714, n25715, n25716, n25717,
    n25718, n25719, n25720, n25721, n25722, n25723,
    n25724, n25725, n25726, n25727, n25728, n25729,
    n25730, n25731, n25732, n25733, n25734, n25736,
    n25737, n25738, n25739, n25740, n25741, n25742,
    n25743, n25744, n25745, n25746, n25747, n25748,
    n25749, n25750, n25751, n25752, n25753, n25754,
    n25755, n25756, n25757, n25758, n25759, n25760,
    n25761, n25762, n25763, n25764, n25765, n25766,
    n25767, n25768, n25769, n25770, n25771, n25772,
    n25773, n25774, n25775, n25776, n25777, n25778,
    n25779, n25780, n25781, n25782, n25783, n25784,
    n25785, n25786, n25787, n25788, n25789, n25790,
    n25791, n25792, n25793, n25794, n25795, n25796,
    n25797, n25798, n25799, n25800, n25801, n25802,
    n25803, n25804, n25805, n25806, n25807, n25808,
    n25809, n25810, n25811, n25812, n25813, n25814,
    n25815, n25816, n25817, n25818, n25819, n25820,
    n25821, n25822, n25823, n25824, n25825, n25826,
    n25827, n25828, n25829, n25830, n25831, n25832,
    n25833, n25834, n25835, n25836, n25837, n25838,
    n25839, n25840, n25841, n25842, n25843, n25844,
    n25845, n25846, n25847, n25848, n25849, n25850,
    n25851, n25852, n25853, n25854, n25855, n25856,
    n25857, n25858, n25859, n25860, n25861, n25862,
    n25863, n25864, n25865, n25866, n25867, n25868,
    n25869, n25870, n25871, n25872, n25873, n25874,
    n25875, n25876, n25877, n25878, n25879, n25880,
    n25881, n25882, n25883, n25884, n25885, n25886,
    n25887, n25888, n25889, n25890, n25891, n25892,
    n25893, n25894, n25895, n25896, n25897, n25898,
    n25899, n25900, n25901, n25902, n25903, n25904,
    n25905, n25906, n25907, n25908, n25909, n25910,
    n25911, n25912, n25913, n25914, n25915, n25916,
    n25917, n25918, n25919, n25920, n25921, n25922,
    n25923, n25924, n25925, n25926, n25927, n25928,
    n25929, n25930, n25931, n25932, n25933, n25934,
    n25935, n25936, n25937, n25938, n25939, n25940,
    n25941, n25942, n25943, n25944, n25946, n25947,
    n25948, n25949, n25950, n25951, n25952, n25953,
    n25954, n25955, n25956, n25957, n25958, n25959,
    n25960, n25961, n25962, n25963, n25964, n25965,
    n25966, n25967, n25968, n25969, n25970, n25971,
    n25972, n25973, n25974, n25975, n25976, n25977,
    n25978, n25979, n25980, n25981, n25982, n25983,
    n25984, n25985, n25986, n25987, n25988, n25989,
    n25990, n25991, n25992, n25993, n25994, n25995,
    n25996, n25997, n25998, n25999, n26000, n26001,
    n26002, n26003, n26004, n26005, n26006, n26007,
    n26008, n26009, n26010, n26011, n26012, n26013,
    n26014, n26015, n26016, n26017, n26018, n26019,
    n26020, n26021, n26022, n26023, n26024, n26025,
    n26026, n26027, n26028, n26029, n26030, n26031,
    n26032, n26033, n26034, n26035, n26036, n26037,
    n26038, n26039, n26040, n26041, n26042, n26043,
    n26044, n26045, n26046, n26047, n26048, n26049,
    n26050, n26051, n26052, n26053, n26054, n26055,
    n26056, n26057, n26058, n26059, n26060, n26061,
    n26062, n26063, n26064, n26065, n26066, n26067,
    n26068, n26069, n26070, n26071, n26072, n26073,
    n26074, n26075, n26076, n26077, n26078, n26079,
    n26080, n26081, n26082, n26083, n26084, n26085,
    n26086, n26087, n26088, n26089, n26090, n26091,
    n26092, n26093, n26094, n26095, n26096, n26097,
    n26098, n26099, n26100, n26101, n26102, n26103,
    n26104, n26105, n26106, n26107, n26108, n26109,
    n26110, n26111, n26112, n26113, n26114, n26115,
    n26116, n26117, n26118, n26119, n26120, n26121,
    n26122, n26123, n26124, n26125, n26126, n26127,
    n26128, n26129, n26130, n26131, n26132, n26133,
    n26134, n26135, n26136, n26137, n26138, n26139,
    n26140, n26142, n26143, n26144, n26145, n26146,
    n26147, n26148, n26149, n26150, n26151, n26152,
    n26153, n26154, n26155, n26156, n26157, n26158,
    n26159, n26160, n26161, n26162, n26163, n26164,
    n26165, n26166, n26167, n26168, n26169, n26170,
    n26171, n26172, n26173, n26174, n26175, n26176,
    n26177, n26178, n26179, n26180, n26181, n26182,
    n26183, n26184, n26185, n26186, n26187, n26188,
    n26189, n26190, n26191, n26192, n26193, n26194,
    n26195, n26196, n26197, n26198, n26199, n26200,
    n26201, n26202, n26203, n26204, n26205, n26206,
    n26207, n26208, n26209, n26210, n26211, n26212,
    n26213, n26214, n26215, n26216, n26217, n26218,
    n26219, n26220, n26221, n26222, n26223, n26224,
    n26225, n26226, n26227, n26228, n26229, n26230,
    n26231, n26232, n26233, n26234, n26235, n26236,
    n26237, n26238, n26239, n26240, n26241, n26242,
    n26243, n26244, n26245, n26246, n26247, n26248,
    n26249, n26250, n26251, n26252, n26253, n26254,
    n26255, n26256, n26257, n26258, n26259, n26260,
    n26261, n26262, n26263, n26264, n26265, n26266,
    n26267, n26268, n26269, n26270, n26271, n26272,
    n26273, n26274, n26275, n26276, n26277, n26278,
    n26279, n26280, n26281, n26282, n26283, n26284,
    n26285, n26286, n26287, n26288, n26289, n26290,
    n26291, n26292, n26293, n26294, n26295, n26296,
    n26297, n26298, n26299, n26300, n26301, n26302,
    n26303, n26304, n26305, n26306, n26307, n26308,
    n26309, n26310, n26311, n26312, n26313, n26314,
    n26315, n26316, n26317, n26318, n26319, n26320,
    n26321, n26322, n26323, n26324, n26325, n26326,
    n26327, n26328, n26329, n26330, n26331, n26332,
    n26333, n26334, n26335, n26336, n26337, n26338,
    n26339, n26340, n26342, n26343, n26344, n26345,
    n26346, n26347, n26348, n26349, n26350, n26351,
    n26352, n26353, n26354, n26355, n26356, n26357,
    n26358, n26359, n26360, n26361, n26362, n26363,
    n26364, n26365, n26366, n26367, n26368, n26369,
    n26370, n26371, n26372, n26373, n26374, n26375,
    n26376, n26377, n26378, n26379, n26380, n26381,
    n26382, n26383, n26384, n26385, n26386, n26387,
    n26388, n26389, n26390, n26391, n26392, n26393,
    n26394, n26395, n26396, n26397, n26398, n26399,
    n26400, n26401, n26402, n26403, n26404, n26405,
    n26406, n26407, n26408, n26409, n26410, n26411,
    n26412, n26413, n26414, n26415, n26416, n26417,
    n26418, n26419, n26420, n26421, n26422, n26423,
    n26424, n26425, n26426, n26427, n26428, n26429,
    n26430, n26431, n26432, n26433, n26434, n26435,
    n26436, n26437, n26438, n26439, n26440, n26441,
    n26442, n26443, n26444, n26445, n26446, n26447,
    n26448, n26449, n26450, n26451, n26452, n26453,
    n26454, n26455, n26456, n26457, n26458, n26459,
    n26460, n26461, n26462, n26463, n26464, n26465,
    n26466, n26467, n26468, n26469, n26470, n26471,
    n26472, n26473, n26474, n26475, n26476, n26477,
    n26478, n26479, n26480, n26481, n26482, n26483,
    n26484, n26485, n26486, n26487, n26488, n26489,
    n26490, n26491, n26492, n26493, n26494, n26495,
    n26496, n26497, n26498, n26499, n26500, n26501,
    n26502, n26503, n26504, n26505, n26506, n26507,
    n26508, n26509, n26510, n26511, n26512, n26513,
    n26514, n26515, n26516, n26517, n26518, n26519,
    n26520, n26521, n26522, n26523, n26524, n26525,
    n26526, n26527, n26528, n26529, n26530, n26532,
    n26533, n26534, n26535, n26536, n26537, n26538,
    n26539, n26540, n26541, n26542, n26543, n26544,
    n26545, n26546, n26547, n26548, n26549, n26550,
    n26551, n26552, n26553, n26554, n26555, n26556,
    n26557, n26558, n26559, n26560, n26561, n26562,
    n26563, n26564, n26565, n26566, n26567, n26568,
    n26569, n26570, n26571, n26572, n26573, n26574,
    n26575, n26576, n26577, n26578, n26579, n26580,
    n26581, n26582, n26583, n26584, n26585, n26586,
    n26587, n26588, n26589, n26590, n26591, n26592,
    n26593, n26594, n26595, n26596, n26597, n26598,
    n26599, n26600, n26601, n26602, n26603, n26604,
    n26605, n26606, n26607, n26608, n26609, n26610,
    n26611, n26612, n26613, n26614, n26615, n26616,
    n26617, n26618, n26619, n26620, n26621, n26622,
    n26623, n26624, n26625, n26626, n26627, n26628,
    n26629, n26630, n26631, n26632, n26633, n26634,
    n26635, n26636, n26637, n26638, n26639, n26640,
    n26641, n26642, n26643, n26644, n26645, n26646,
    n26647, n26648, n26649, n26650, n26651, n26652,
    n26653, n26654, n26655, n26656, n26657, n26658,
    n26659, n26660, n26661, n26662, n26663, n26664,
    n26665, n26666, n26667, n26668, n26669, n26670,
    n26671, n26672, n26673, n26674, n26675, n26676,
    n26677, n26678, n26679, n26680, n26681, n26682,
    n26683, n26684, n26685, n26686, n26687, n26688,
    n26689, n26690, n26691, n26692, n26693, n26694,
    n26695, n26696, n26697, n26698, n26699, n26700,
    n26701, n26702, n26703, n26704, n26705, n26706,
    n26707, n26708, n26709, n26710, n26711, n26712,
    n26713, n26714, n26715, n26717, n26718, n26719,
    n26720, n26721, n26722, n26723, n26724, n26725,
    n26726, n26727, n26728, n26729, n26730, n26731,
    n26732, n26733, n26734, n26735, n26736, n26737,
    n26738, n26739, n26740, n26741, n26742, n26743,
    n26744, n26745, n26746, n26747, n26748, n26749,
    n26750, n26751, n26752, n26753, n26754, n26755,
    n26756, n26757, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767,
    n26768, n26769, n26770, n26771, n26772, n26773,
    n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785,
    n26786, n26787, n26788, n26789, n26790, n26791,
    n26792, n26793, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26802, n26803,
    n26804, n26805, n26806, n26807, n26808, n26809,
    n26810, n26811, n26812, n26813, n26814, n26815,
    n26816, n26817, n26818, n26819, n26820, n26821,
    n26822, n26823, n26824, n26825, n26826, n26827,
    n26828, n26829, n26830, n26831, n26832, n26833,
    n26834, n26835, n26836, n26837, n26838, n26839,
    n26840, n26841, n26842, n26843, n26844, n26845,
    n26846, n26847, n26848, n26849, n26850, n26851,
    n26852, n26853, n26854, n26855, n26856, n26857,
    n26858, n26859, n26860, n26861, n26862, n26863,
    n26864, n26865, n26866, n26867, n26868, n26869,
    n26870, n26871, n26872, n26873, n26874, n26875,
    n26876, n26877, n26878, n26879, n26880, n26881,
    n26882, n26883, n26884, n26885, n26886, n26887,
    n26888, n26889, n26890, n26891, n26892, n26893,
    n26894, n26895, n26896, n26897, n26898, n26899,
    n26900, n26901, n26902, n26903, n26905, n26906,
    n26907, n26908, n26909, n26910, n26911, n26912,
    n26913, n26914, n26915, n26916, n26917, n26918,
    n26919, n26920, n26921, n26922, n26923, n26924,
    n26925, n26926, n26927, n26928, n26929, n26930,
    n26931, n26932, n26933, n26934, n26935, n26936,
    n26937, n26938, n26939, n26940, n26941, n26942,
    n26943, n26944, n26945, n26946, n26947, n26948,
    n26949, n26950, n26951, n26952, n26953, n26954,
    n26955, n26956, n26957, n26958, n26959, n26960,
    n26961, n26962, n26963, n26964, n26965, n26966,
    n26967, n26968, n26969, n26970, n26971, n26972,
    n26973, n26974, n26975, n26976, n26977, n26978,
    n26979, n26980, n26981, n26982, n26983, n26984,
    n26985, n26986, n26987, n26988, n26989, n26990,
    n26991, n26992, n26993, n26994, n26995, n26996,
    n26997, n26998, n26999, n27000, n27001, n27002,
    n27003, n27004, n27005, n27006, n27007, n27008,
    n27009, n27010, n27011, n27012, n27013, n27014,
    n27015, n27016, n27017, n27018, n27019, n27020,
    n27021, n27022, n27023, n27024, n27025, n27026,
    n27027, n27028, n27029, n27030, n27031, n27032,
    n27033, n27034, n27035, n27036, n27037, n27038,
    n27039, n27040, n27041, n27042, n27043, n27044,
    n27045, n27046, n27047, n27048, n27049, n27050,
    n27051, n27052, n27053, n27054, n27055, n27056,
    n27057, n27058, n27059, n27060, n27061, n27062,
    n27063, n27064, n27065, n27066, n27067, n27068,
    n27069, n27070, n27071, n27072, n27073, n27074,
    n27075, n27076, n27077, n27078, n27079, n27080,
    n27081, n27082, n27083, n27084, n27085, n27086,
    n27087, n27088, n27089, n27090, n27092, n27093,
    n27094, n27095, n27096, n27097, n27098, n27099,
    n27100, n27101, n27102, n27103, n27104, n27105,
    n27106, n27107, n27108, n27109, n27110, n27111,
    n27112, n27113, n27114, n27115, n27116, n27117,
    n27118, n27119, n27120, n27121, n27122, n27123,
    n27124, n27125, n27126, n27127, n27128, n27129,
    n27130, n27131, n27132, n27133, n27134, n27135,
    n27136, n27137, n27138, n27139, n27140, n27141,
    n27142, n27143, n27144, n27145, n27146, n27147,
    n27148, n27149, n27150, n27151, n27152, n27153,
    n27154, n27155, n27156, n27157, n27158, n27159,
    n27160, n27161, n27162, n27163, n27164, n27165,
    n27166, n27167, n27168, n27169, n27170, n27171,
    n27172, n27173, n27174, n27175, n27176, n27177,
    n27178, n27179, n27180, n27181, n27182, n27183,
    n27184, n27185, n27186, n27187, n27188, n27189,
    n27190, n27191, n27192, n27193, n27194, n27195,
    n27196, n27197, n27198, n27199, n27200, n27201,
    n27202, n27203, n27204, n27205, n27206, n27207,
    n27208, n27209, n27210, n27211, n27212, n27213,
    n27214, n27215, n27216, n27217, n27218, n27219,
    n27220, n27221, n27222, n27223, n27224, n27225,
    n27226, n27227, n27228, n27229, n27230, n27231,
    n27232, n27233, n27234, n27235, n27236, n27237,
    n27238, n27239, n27240, n27241, n27242, n27243,
    n27244, n27245, n27246, n27247, n27248, n27249,
    n27250, n27251, n27252, n27253, n27254, n27255,
    n27256, n27257, n27259, n27260, n27261, n27262,
    n27263, n27264, n27265, n27266, n27267, n27268,
    n27269, n27270, n27271, n27272, n27273, n27274,
    n27275, n27276, n27277, n27278, n27279, n27280,
    n27281, n27282, n27283, n27284, n27285, n27286,
    n27287, n27288, n27289, n27290, n27291, n27292,
    n27293, n27294, n27295, n27296, n27297, n27298,
    n27299, n27300, n27301, n27302, n27303, n27304,
    n27305, n27306, n27307, n27308, n27309, n27310,
    n27311, n27312, n27313, n27314, n27315, n27316,
    n27317, n27318, n27319, n27320, n27321, n27322,
    n27323, n27324, n27325, n27326, n27327, n27328,
    n27329, n27330, n27331, n27332, n27333, n27334,
    n27335, n27336, n27337, n27338, n27339, n27340,
    n27341, n27342, n27343, n27344, n27345, n27346,
    n27347, n27348, n27349, n27350, n27351, n27352,
    n27353, n27354, n27355, n27356, n27357, n27358,
    n27359, n27360, n27361, n27362, n27363, n27364,
    n27365, n27366, n27367, n27368, n27369, n27370,
    n27371, n27372, n27373, n27374, n27375, n27376,
    n27377, n27378, n27379, n27380, n27381, n27382,
    n27383, n27384, n27385, n27386, n27387, n27388,
    n27389, n27390, n27391, n27392, n27393, n27394,
    n27395, n27396, n27397, n27398, n27399, n27400,
    n27401, n27402, n27403, n27404, n27405, n27406,
    n27407, n27408, n27409, n27410, n27411, n27412,
    n27413, n27414, n27416, n27417, n27418, n27419,
    n27420, n27421, n27422, n27423, n27424, n27425,
    n27426, n27427, n27428, n27429, n27430, n27431,
    n27432, n27433, n27434, n27435, n27436, n27437,
    n27438, n27439, n27440, n27441, n27442, n27443,
    n27444, n27445, n27446, n27447, n27448, n27449,
    n27450, n27451, n27452, n27453, n27454, n27455,
    n27456, n27457, n27458, n27459, n27460, n27461,
    n27462, n27463, n27464, n27465, n27466, n27467,
    n27468, n27469, n27470, n27471, n27472, n27473,
    n27474, n27475, n27476, n27477, n27478, n27479,
    n27480, n27481, n27482, n27483, n27484, n27485,
    n27486, n27487, n27488, n27489, n27490, n27491,
    n27492, n27493, n27494, n27495, n27496, n27497,
    n27498, n27499, n27500, n27501, n27502, n27503,
    n27504, n27505, n27506, n27507, n27508, n27509,
    n27510, n27511, n27512, n27513, n27514, n27515,
    n27516, n27517, n27518, n27519, n27520, n27521,
    n27522, n27523, n27524, n27525, n27526, n27527,
    n27528, n27529, n27530, n27531, n27532, n27533,
    n27534, n27535, n27536, n27537, n27538, n27539,
    n27540, n27541, n27542, n27543, n27544, n27545,
    n27546, n27547, n27548, n27549, n27550, n27551,
    n27552, n27553, n27554, n27555, n27556, n27557,
    n27558, n27559, n27560, n27561, n27562, n27563,
    n27564, n27565, n27566, n27567, n27568, n27569,
    n27570, n27572, n27573, n27574, n27575, n27576,
    n27577, n27578, n27579, n27580, n27581, n27582,
    n27583, n27584, n27585, n27586, n27587, n27588,
    n27589, n27590, n27591, n27592, n27593, n27594,
    n27595, n27596, n27597, n27598, n27599, n27600,
    n27601, n27602, n27603, n27604, n27605, n27606,
    n27607, n27608, n27609, n27610, n27611, n27612,
    n27613, n27614, n27615, n27616, n27617, n27618,
    n27619, n27620, n27621, n27622, n27623, n27624,
    n27625, n27626, n27627, n27628, n27629, n27630,
    n27631, n27632, n27633, n27634, n27635, n27636,
    n27637, n27638, n27639, n27640, n27641, n27642,
    n27643, n27644, n27645, n27646, n27647, n27648,
    n27649, n27650, n27651, n27652, n27653, n27654,
    n27655, n27656, n27657, n27658, n27659, n27660,
    n27661, n27662, n27663, n27664, n27665, n27666,
    n27667, n27668, n27669, n27670, n27671, n27672,
    n27673, n27674, n27675, n27676, n27677, n27678,
    n27679, n27680, n27681, n27682, n27683, n27684,
    n27685, n27686, n27687, n27688, n27689, n27690,
    n27691, n27692, n27693, n27694, n27695, n27696,
    n27697, n27698, n27699, n27700, n27701, n27702,
    n27703, n27704, n27705, n27706, n27707, n27708,
    n27709, n27710, n27711, n27712, n27713, n27714,
    n27715, n27716, n27717, n27718, n27719, n27720,
    n27721, n27723, n27724, n27725, n27726, n27727,
    n27728, n27729, n27730, n27731, n27732, n27733,
    n27734, n27735, n27736, n27737, n27738, n27739,
    n27740, n27741, n27742, n27743, n27744, n27745,
    n27746, n27747, n27748, n27749, n27750, n27751,
    n27752, n27753, n27754, n27755, n27756, n27757,
    n27758, n27759, n27760, n27761, n27762, n27763,
    n27764, n27765, n27766, n27767, n27768, n27769,
    n27770, n27771, n27772, n27773, n27774, n27775,
    n27776, n27777, n27778, n27779, n27780, n27781,
    n27782, n27783, n27784, n27785, n27786, n27787,
    n27788, n27789, n27790, n27791, n27792, n27793,
    n27794, n27795, n27796, n27797, n27798, n27799,
    n27800, n27801, n27802, n27803, n27804, n27805,
    n27806, n27807, n27808, n27809, n27810, n27811,
    n27812, n27813, n27814, n27815, n27816, n27817,
    n27818, n27819, n27820, n27821, n27822, n27823,
    n27824, n27825, n27826, n27827, n27828, n27829,
    n27830, n27831, n27832, n27833, n27834, n27835,
    n27836, n27837, n27838, n27839, n27840, n27841,
    n27842, n27843, n27844, n27845, n27846, n27847,
    n27848, n27849, n27850, n27851, n27852, n27853,
    n27854, n27855, n27856, n27857, n27858, n27859,
    n27860, n27861, n27863, n27864, n27865, n27866,
    n27867, n27868, n27869, n27870, n27871, n27872,
    n27873, n27874, n27875, n27876, n27877, n27878,
    n27879, n27880, n27881, n27882, n27883, n27884,
    n27885, n27886, n27887, n27888, n27889, n27890,
    n27891, n27892, n27893, n27894, n27895, n27896,
    n27897, n27898, n27899, n27900, n27901, n27902,
    n27903, n27904, n27905, n27906, n27907, n27908,
    n27909, n27910, n27911, n27912, n27913, n27914,
    n27915, n27916, n27917, n27918, n27919, n27920,
    n27921, n27922, n27923, n27924, n27925, n27926,
    n27927, n27928, n27929, n27930, n27931, n27932,
    n27933, n27934, n27935, n27936, n27937, n27938,
    n27939, n27940, n27941, n27942, n27943, n27944,
    n27945, n27946, n27947, n27948, n27949, n27950,
    n27951, n27952, n27953, n27954, n27955, n27956,
    n27957, n27958, n27959, n27960, n27961, n27962,
    n27963, n27964, n27965, n27966, n27967, n27968,
    n27969, n27970, n27971, n27972, n27973, n27974,
    n27975, n27976, n27977, n27978, n27979, n27980,
    n27981, n27982, n27983, n27984, n27985, n27986,
    n27987, n27988, n27989, n27990, n27991, n27992,
    n27993, n27994, n27995, n27996, n27997, n27998,
    n27999, n28000, n28001, n28002, n28004, n28005,
    n28006, n28007, n28008, n28009, n28010, n28011,
    n28012, n28013, n28014, n28015, n28016, n28017,
    n28018, n28019, n28020, n28021, n28022, n28023,
    n28024, n28025, n28026, n28027, n28028, n28029,
    n28030, n28031, n28032, n28033, n28034, n28035,
    n28036, n28037, n28038, n28039, n28040, n28041,
    n28042, n28043, n28044, n28045, n28046, n28047,
    n28048, n28049, n28050, n28051, n28052, n28053,
    n28054, n28055, n28056, n28057, n28058, n28059,
    n28060, n28061, n28062, n28063, n28064, n28065,
    n28066, n28067, n28068, n28069, n28070, n28071,
    n28072, n28073, n28074, n28075, n28076, n28077,
    n28078, n28079, n28080, n28081, n28082, n28083,
    n28084, n28085, n28086, n28087, n28088, n28089,
    n28090, n28091, n28092, n28093, n28094, n28095,
    n28096, n28097, n28098, n28099, n28100, n28101,
    n28102, n28103, n28104, n28105, n28106, n28107,
    n28108, n28109, n28110, n28111, n28112, n28113,
    n28114, n28115, n28116, n28117, n28118, n28119,
    n28120, n28121, n28122, n28123, n28124, n28125,
    n28126, n28127, n28128, n28129, n28130, n28131,
    n28132, n28133, n28135, n28136, n28137, n28138,
    n28139, n28140, n28141, n28142, n28143, n28144,
    n28145, n28146, n28147, n28148, n28149, n28150,
    n28151, n28152, n28153, n28154, n28155, n28156,
    n28157, n28158, n28159, n28160, n28161, n28162,
    n28163, n28164, n28165, n28166, n28167, n28168,
    n28169, n28170, n28171, n28172, n28173, n28174,
    n28175, n28176, n28177, n28178, n28179, n28180,
    n28181, n28182, n28183, n28184, n28185, n28186,
    n28187, n28188, n28189, n28190, n28191, n28192,
    n28193, n28194, n28195, n28196, n28197, n28198,
    n28199, n28200, n28201, n28202, n28203, n28204,
    n28205, n28206, n28207, n28208, n28209, n28210,
    n28211, n28212, n28213, n28214, n28215, n28216,
    n28217, n28218, n28219, n28220, n28221, n28222,
    n28223, n28224, n28225, n28226, n28227, n28228,
    n28229, n28230, n28231, n28232, n28233, n28234,
    n28235, n28236, n28237, n28238, n28239, n28240,
    n28241, n28242, n28243, n28244, n28245, n28246,
    n28247, n28248, n28249, n28250, n28251, n28252,
    n28253, n28254, n28255, n28256, n28257, n28258,
    n28260, n28261, n28262, n28263, n28264, n28265,
    n28266, n28267, n28268, n28269, n28270, n28271,
    n28272, n28273, n28274, n28275, n28276, n28277,
    n28278, n28279, n28280, n28281, n28282, n28283,
    n28284, n28285, n28286, n28287, n28288, n28289,
    n28290, n28291, n28292, n28293, n28294, n28295,
    n28296, n28297, n28298, n28299, n28300, n28301,
    n28302, n28303, n28304, n28305, n28306, n28307,
    n28308, n28309, n28310, n28311, n28312, n28313,
    n28314, n28315, n28316, n28317, n28318, n28319,
    n28320, n28321, n28322, n28323, n28324, n28325,
    n28326, n28327, n28328, n28329, n28330, n28331,
    n28332, n28333, n28334, n28335, n28336, n28337,
    n28338, n28339, n28340, n28341, n28342, n28343,
    n28344, n28345, n28346, n28347, n28348, n28349,
    n28350, n28351, n28352, n28353, n28354, n28355,
    n28356, n28357, n28358, n28359, n28360, n28361,
    n28362, n28363, n28364, n28365, n28366, n28367,
    n28368, n28369, n28370, n28371, n28372, n28373,
    n28374, n28375, n28376, n28377, n28378, n28379,
    n28380, n28381, n28383, n28384, n28385, n28386,
    n28387, n28388, n28389, n28390, n28391, n28392,
    n28393, n28394, n28395, n28396, n28397, n28398,
    n28399, n28400, n28401, n28402, n28403, n28404,
    n28405, n28406, n28407, n28408, n28409, n28410,
    n28411, n28412, n28413, n28414, n28415, n28416,
    n28417, n28418, n28419, n28420, n28421, n28422,
    n28423, n28424, n28425, n28426, n28427, n28428,
    n28429, n28430, n28431, n28432, n28433, n28434,
    n28435, n28436, n28437, n28438, n28439, n28440,
    n28441, n28442, n28443, n28444, n28445, n28446,
    n28447, n28448, n28449, n28450, n28451, n28452,
    n28453, n28454, n28455, n28456, n28457, n28458,
    n28459, n28460, n28461, n28462, n28463, n28464,
    n28465, n28466, n28467, n28468, n28469, n28470,
    n28471, n28472, n28473, n28474, n28475, n28476,
    n28477, n28478, n28479, n28480, n28481, n28482,
    n28483, n28484, n28485, n28486, n28487, n28488,
    n28489, n28490, n28491, n28492, n28493, n28494,
    n28495, n28496, n28498, n28499, n28500, n28501,
    n28502, n28503, n28504, n28505, n28506, n28507,
    n28508, n28509, n28510, n28511, n28512, n28513,
    n28514, n28515, n28516, n28517, n28518, n28519,
    n28520, n28521, n28522, n28523, n28524, n28525,
    n28526, n28527, n28528, n28529, n28530, n28531,
    n28532, n28533, n28534, n28535, n28536, n28537,
    n28538, n28539, n28540, n28541, n28542, n28543,
    n28544, n28545, n28546, n28547, n28548, n28549,
    n28550, n28551, n28552, n28553, n28554, n28555,
    n28556, n28557, n28558, n28559, n28560, n28561,
    n28562, n28563, n28564, n28565, n28566, n28567,
    n28568, n28569, n28570, n28571, n28572, n28573,
    n28574, n28575, n28576, n28577, n28578, n28579,
    n28580, n28581, n28582, n28583, n28584, n28585,
    n28586, n28587, n28588, n28589, n28590, n28591,
    n28592, n28593, n28594, n28595, n28596, n28597,
    n28598, n28599, n28600, n28601, n28602, n28603,
    n28604, n28606, n28607, n28608, n28609, n28610,
    n28611, n28612, n28613, n28614, n28615, n28616,
    n28617, n28618, n28619, n28620, n28621, n28622,
    n28623, n28624, n28625, n28626, n28627, n28628,
    n28629, n28630, n28631, n28632, n28633, n28634,
    n28635, n28636, n28637, n28638, n28639, n28640,
    n28641, n28642, n28643, n28644, n28645, n28646,
    n28647, n28648, n28649, n28650, n28651, n28652,
    n28653, n28654, n28655, n28656, n28657, n28658,
    n28659, n28660, n28661, n28662, n28663, n28664,
    n28665, n28666, n28667, n28668, n28669, n28670,
    n28671, n28672, n28673, n28674, n28675, n28676,
    n28677, n28678, n28679, n28680, n28681, n28682,
    n28683, n28684, n28685, n28686, n28687, n28688,
    n28689, n28690, n28691, n28692, n28693, n28694,
    n28695, n28696, n28697, n28698, n28699, n28700,
    n28701, n28702, n28703, n28704, n28705, n28706,
    n28708, n28709, n28710, n28711, n28712, n28713,
    n28714, n28715, n28716, n28717, n28718, n28719,
    n28720, n28721, n28722, n28723, n28724, n28725,
    n28726, n28727, n28728, n28729, n28730, n28731,
    n28732, n28733, n28734, n28735, n28736, n28737,
    n28738, n28739, n28740, n28741, n28742, n28743,
    n28744, n28745, n28746, n28747, n28748, n28749,
    n28750, n28751, n28752, n28753, n28754, n28755,
    n28756, n28757, n28758, n28759, n28760, n28761,
    n28762, n28763, n28764, n28765, n28766, n28767,
    n28768, n28769, n28770, n28771, n28772, n28773,
    n28774, n28775, n28776, n28777, n28778, n28779,
    n28780, n28781, n28782, n28783, n28784, n28785,
    n28786, n28787, n28788, n28789, n28790, n28791,
    n28792, n28793, n28794, n28795, n28796, n28797,
    n28798, n28799, n28800, n28801, n28802, n28803,
    n28804, n28805, n28806, n28807, n28808, n28810,
    n28811, n28812, n28813, n28814, n28815, n28816,
    n28817, n28818, n28819, n28820, n28821, n28822,
    n28823, n28824, n28825, n28826, n28827, n28828,
    n28829, n28830, n28831, n28832, n28833, n28834,
    n28835, n28836, n28837, n28838, n28839, n28840,
    n28841, n28842, n28843, n28844, n28845, n28846,
    n28847, n28848, n28849, n28850, n28851, n28852,
    n28853, n28854, n28855, n28856, n28857, n28858,
    n28859, n28860, n28861, n28862, n28863, n28864,
    n28865, n28866, n28867, n28868, n28869, n28870,
    n28871, n28872, n28873, n28874, n28875, n28876,
    n28877, n28878, n28879, n28880, n28881, n28882,
    n28883, n28884, n28885, n28886, n28887, n28888,
    n28889, n28890, n28891, n28892, n28893, n28894,
    n28895, n28896, n28897, n28898, n28900, n28901,
    n28902, n28903, n28904, n28905, n28906, n28907,
    n28908, n28909, n28910, n28911, n28912, n28913,
    n28914, n28915, n28916, n28917, n28918, n28919,
    n28920, n28921, n28922, n28923, n28924, n28925,
    n28926, n28927, n28928, n28929, n28930, n28931,
    n28932, n28933, n28934, n28935, n28936, n28937,
    n28938, n28939, n28940, n28941, n28942, n28943,
    n28944, n28945, n28946, n28947, n28948, n28949,
    n28950, n28951, n28952, n28953, n28954, n28955,
    n28956, n28957, n28958, n28959, n28960, n28961,
    n28962, n28963, n28964, n28965, n28966, n28967,
    n28968, n28969, n28970, n28971, n28972, n28973,
    n28974, n28975, n28976, n28977, n28978, n28979,
    n28980, n28981, n28982, n28983, n28984, n28985,
    n28986, n28988, n28989, n28990, n28991, n28992,
    n28993, n28994, n28995, n28996, n28997, n28998,
    n28999, n29000, n29001, n29002, n29003, n29004,
    n29005, n29006, n29007, n29008, n29009, n29010,
    n29011, n29012, n29013, n29014, n29015, n29016,
    n29017, n29018, n29019, n29020, n29021, n29022,
    n29023, n29024, n29025, n29026, n29027, n29028,
    n29029, n29030, n29031, n29032, n29033, n29034,
    n29035, n29036, n29037, n29038, n29039, n29040,
    n29041, n29042, n29043, n29044, n29045, n29046,
    n29047, n29048, n29049, n29050, n29051, n29052,
    n29053, n29054, n29055, n29056, n29057, n29058,
    n29059, n29060, n29061, n29062, n29063, n29064,
    n29065, n29066, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077,
    n29078, n29079, n29080, n29081, n29082, n29083,
    n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095,
    n29096, n29097, n29098, n29099, n29100, n29101,
    n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113,
    n29114, n29115, n29116, n29117, n29118, n29119,
    n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131,
    n29132, n29133, n29134, n29135, n29136, n29137,
    n29138, n29139, n29140, n29142, n29143, n29144,
    n29145, n29146, n29147, n29148, n29149, n29150,
    n29151, n29152, n29153, n29154, n29155, n29156,
    n29157, n29158, n29159, n29160, n29161, n29162,
    n29163, n29164, n29165, n29166, n29167, n29168,
    n29169, n29170, n29171, n29172, n29173, n29174,
    n29175, n29176, n29177, n29178, n29179, n29180,
    n29181, n29182, n29183, n29184, n29185, n29186,
    n29187, n29188, n29189, n29190, n29191, n29192,
    n29193, n29194, n29195, n29196, n29197, n29198,
    n29199, n29200, n29201, n29202, n29203, n29205,
    n29206, n29207, n29208, n29209, n29210, n29211,
    n29212, n29213, n29214, n29215, n29216, n29217,
    n29218, n29219, n29220, n29221, n29222, n29223,
    n29224, n29225, n29226, n29227, n29228, n29229,
    n29230, n29231, n29232, n29233, n29234, n29235,
    n29236, n29237, n29238, n29239, n29240, n29241,
    n29242, n29243, n29244, n29245, n29246, n29247,
    n29248, n29249, n29250, n29251, n29252, n29253,
    n29254, n29255, n29256;
  assign n65 = ~pi2  & ~pi3 ;
  assign n66 = pi2  & pi3 ;
  assign n67 = ~n65 & ~n66;
  assign n68 = ~pi4  & ~pi5 ;
  assign n69 = pi4  & pi5 ;
  assign n70 = ~n68 & ~n69;
  assign n71 = n67 & ~n70;
  assign n72 = ~pi20  & ~pi21 ;
  assign n73 = pi20  & pi21 ;
  assign n74 = ~n72 & ~n73;
  assign n75 = ~pi22  & ~pi23 ;
  assign n76 = pi22  & pi23 ;
  assign n77 = ~n75 & ~n76;
  assign n78 = n74 & n77;
  assign n79 = pi27  & pi28 ;
  assign n80 = ~pi29  & pi30 ;
  assign n81 = n79 & n80;
  assign n82 = pi24  & ~pi25 ;
  assign n83 = ~pi23  & pi26 ;
  assign n84 = n82 & n83;
  assign n85 = n81 & n84;
  assign n86 = ~pi27  & pi28 ;
  assign n87 = pi29  & ~pi30 ;
  assign n88 = n86 & n87;
  assign n89 = pi23  & ~pi26 ;
  assign n90 = n82 & n89;
  assign n91 = n88 & n90;
  assign n92 = n81 & n90;
  assign n93 = ~n91 & ~n92;
  assign n94 = n79 & n87;
  assign n95 = ~pi24  & pi25 ;
  assign n96 = ~pi23  & ~pi26 ;
  assign n97 = n95 & n96;
  assign n98 = n94 & n97;
  assign n99 = pi24  & pi25 ;
  assign n100 = n83 & n99;
  assign n101 = pi27  & ~pi28 ;
  assign n102 = n87 & n101;
  assign n103 = n100 & n102;
  assign n104 = ~n98 & ~n103;
  assign n105 = ~pi29  & ~pi30 ;
  assign n106 = ~pi27  & ~pi28 ;
  assign n107 = n105 & n106;
  assign n108 = n89 & n95;
  assign n109 = n107 & n108;
  assign n110 = n86 & n105;
  assign n111 = pi23  & pi26 ;
  assign n112 = n95 & n111;
  assign n113 = n110 & n112;
  assign n114 = ~n109 & ~n113;
  assign n115 = pi29  & pi30 ;
  assign n116 = n86 & n115;
  assign n117 = n83 & n95;
  assign n118 = n116 & n117;
  assign n119 = n79 & n115;
  assign n120 = n100 & n119;
  assign n121 = ~n118 & ~n120;
  assign n122 = n100 & n116;
  assign n123 = ~pi24  & ~pi25 ;
  assign n124 = n111 & n123;
  assign n125 = n119 & n124;
  assign n126 = n112 & n119;
  assign n127 = ~n122 & ~n125;
  assign n128 = ~n126 & n127;
  assign n129 = n121 & n128;
  assign n130 = n101 & n105;
  assign n131 = n100 & n130;
  assign n132 = n89 & n123;
  assign n133 = n110 & n132;
  assign n134 = n94 & n108;
  assign n135 = n89 & n99;
  assign n136 = n94 & n135;
  assign n137 = ~n134 & ~n136;
  assign n138 = n83 & n123;
  assign n139 = n107 & n138;
  assign n140 = n96 & n99;
  assign n141 = n94 & n140;
  assign n142 = ~n139 & ~n141;
  assign n143 = n99 & n111;
  assign n144 = n88 & n143;
  assign n145 = n102 & n132;
  assign n146 = ~n144 & ~n145;
  assign n147 = n84 & n102;
  assign n148 = n88 & n100;
  assign n149 = n88 & n97;
  assign n150 = ~n148 & ~n149;
  assign n151 = n146 & ~n147;
  assign n152 = n150 & n151;
  assign n153 = ~n85 & ~n131;
  assign n154 = ~n133 & n153;
  assign n155 = n93 & n104;
  assign n156 = n114 & n137;
  assign n157 = n142 & n156;
  assign n158 = n154 & n155;
  assign n159 = n157 & n158;
  assign n160 = n129 & n152;
  assign n161 = n159 & n160;
  assign n162 = n88 & n124;
  assign n163 = n102 & n117;
  assign n164 = n102 & n108;
  assign n165 = n102 & n135;
  assign n166 = ~n164 & ~n165;
  assign n167 = n88 & n117;
  assign n168 = n88 & n138;
  assign n169 = ~n167 & ~n168;
  assign n170 = n166 & n169;
  assign n171 = n82 & n96;
  assign n172 = n102 & n171;
  assign n173 = n88 & n171;
  assign n174 = ~n172 & ~n173;
  assign n175 = n102 & n124;
  assign n176 = n96 & n123;
  assign n177 = n94 & n176;
  assign n178 = ~n175 & ~n177;
  assign n179 = n90 & n102;
  assign n180 = n102 & n112;
  assign n181 = n82 & n111;
  assign n182 = n88 & n181;
  assign n183 = n88 & n135;
  assign n184 = ~n162 & ~n163;
  assign n185 = ~n179 & ~n180;
  assign n186 = ~n182 & ~n183;
  assign n187 = n185 & n186;
  assign n188 = n174 & n184;
  assign n189 = n178 & n188;
  assign n190 = n170 & n187;
  assign n191 = n189 & n190;
  assign n192 = n102 & n181;
  assign n193 = n102 & n140;
  assign n194 = ~n192 & ~n193;
  assign n195 = n88 & n108;
  assign n196 = n88 & n112;
  assign n197 = ~n195 & ~n196;
  assign n198 = n194 & n197;
  assign n199 = n119 & n181;
  assign n200 = n119 & n143;
  assign n201 = ~n199 & ~n200;
  assign n202 = n117 & n119;
  assign n203 = n84 & n119;
  assign n204 = ~n202 & ~n203;
  assign n205 = n201 & n204;
  assign n206 = n79 & n105;
  assign n207 = n176 & n206;
  assign n208 = n171 & n206;
  assign n209 = n100 & n110;
  assign n210 = n112 & n130;
  assign n211 = ~n209 & ~n210;
  assign n212 = n110 & n176;
  assign n213 = n130 & n143;
  assign n214 = ~n212 & ~n213;
  assign n215 = n97 & n110;
  assign n216 = n110 & n140;
  assign n217 = ~n215 & ~n216;
  assign n218 = n110 & n124;
  assign n219 = n108 & n110;
  assign n220 = ~n218 & ~n219;
  assign n221 = n110 & n143;
  assign n222 = n110 & n171;
  assign n223 = ~n221 & ~n222;
  assign n224 = n110 & n138;
  assign n225 = n110 & n117;
  assign n226 = ~n224 & ~n225;
  assign n227 = ~n207 & ~n208;
  assign n228 = n211 & n227;
  assign n229 = n214 & n217;
  assign n230 = n220 & n223;
  assign n231 = n226 & n230;
  assign n232 = n228 & n229;
  assign n233 = n231 & n232;
  assign n234 = n110 & n135;
  assign n235 = n90 & n94;
  assign n236 = n119 & n140;
  assign n237 = ~n235 & ~n236;
  assign n238 = n94 & n171;
  assign n239 = n107 & n135;
  assign n240 = n94 & n132;
  assign n241 = ~n239 & ~n240;
  assign n242 = n119 & n132;
  assign n243 = n97 & n119;
  assign n244 = n108 & n119;
  assign n245 = n90 & n119;
  assign n246 = n119 & n138;
  assign n247 = n119 & n135;
  assign n248 = ~n245 & ~n246;
  assign n249 = ~n247 & n248;
  assign n250 = n119 & n171;
  assign n251 = n112 & n116;
  assign n252 = ~n250 & ~n251;
  assign n253 = n116 & n143;
  assign n254 = n119 & n176;
  assign n255 = ~n253 & ~n254;
  assign n256 = ~n242 & ~n243;
  assign n257 = ~n244 & n256;
  assign n258 = n252 & n255;
  assign n259 = n257 & n258;
  assign n260 = n249 & n259;
  assign n261 = ~n234 & ~n238;
  assign n262 = n237 & n261;
  assign n263 = n241 & n262;
  assign n264 = n260 & n263;
  assign n265 = n81 & n100;
  assign n266 = n106 & n115;
  assign n267 = n97 & n266;
  assign n268 = ~n265 & ~n267;
  assign n269 = n108 & n266;
  assign n270 = n81 & n143;
  assign n271 = n81 & n117;
  assign n272 = ~n269 & ~n270;
  assign n273 = ~n271 & n272;
  assign n274 = n268 & n273;
  assign n275 = n101 & n115;
  assign n276 = n100 & n275;
  assign n277 = n116 & n181;
  assign n278 = ~n276 & ~n277;
  assign n279 = n108 & n116;
  assign n280 = n116 & n140;
  assign n281 = ~n279 & ~n280;
  assign n282 = n116 & n132;
  assign n283 = n117 & n275;
  assign n284 = ~n282 & ~n283;
  assign n285 = n116 & n176;
  assign n286 = n90 & n116;
  assign n287 = n116 & n124;
  assign n288 = n143 & n275;
  assign n289 = n97 & n116;
  assign n290 = n116 & n138;
  assign n291 = ~n285 & ~n286;
  assign n292 = ~n287 & ~n288;
  assign n293 = ~n289 & ~n290;
  assign n294 = n292 & n293;
  assign n295 = n291 & n294;
  assign n296 = n84 & n116;
  assign n297 = n116 & n171;
  assign n298 = ~n296 & ~n297;
  assign n299 = n116 & n135;
  assign n300 = n112 & n275;
  assign n301 = ~n299 & ~n300;
  assign n302 = n278 & n301;
  assign n303 = n281 & n284;
  assign n304 = n298 & n303;
  assign n305 = n302 & n304;
  assign n306 = n295 & n305;
  assign n307 = n107 & n171;
  assign n308 = n90 & n107;
  assign n309 = ~n307 & ~n308;
  assign n310 = n107 & n132;
  assign n311 = n107 & n176;
  assign n312 = n124 & n266;
  assign n313 = n132 & n275;
  assign n314 = ~n312 & ~n313;
  assign n315 = n108 & n275;
  assign n316 = n124 & n275;
  assign n317 = ~n315 & ~n316;
  assign n318 = n181 & n266;
  assign n319 = n97 & n275;
  assign n320 = n143 & n266;
  assign n321 = n84 & n266;
  assign n322 = ~n320 & ~n321;
  assign n323 = n171 & n275;
  assign n324 = n100 & n266;
  assign n325 = ~n323 & ~n324;
  assign n326 = n140 & n275;
  assign n327 = n181 & n275;
  assign n328 = ~n326 & ~n327;
  assign n329 = ~n318 & ~n319;
  assign n330 = n317 & n329;
  assign n331 = n322 & n325;
  assign n332 = n328 & n331;
  assign n333 = n330 & n332;
  assign n334 = n117 & n266;
  assign n335 = n90 & n275;
  assign n336 = n176 & n275;
  assign n337 = ~n335 & ~n336;
  assign n338 = n138 & n275;
  assign n339 = n138 & n266;
  assign n340 = n84 & n275;
  assign n341 = ~n339 & ~n340;
  assign n342 = n112 & n266;
  assign n343 = n135 & n275;
  assign n344 = ~n342 & ~n343;
  assign n345 = n341 & n344;
  assign n346 = ~n334 & ~n338;
  assign n347 = n337 & n346;
  assign n348 = n345 & n347;
  assign n349 = ~n310 & ~n311;
  assign n350 = n309 & n349;
  assign n351 = n314 & n350;
  assign n352 = n348 & n351;
  assign n353 = n333 & n352;
  assign n354 = n97 & n107;
  assign n355 = n81 & n181;
  assign n356 = n132 & n266;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~n354 & n357;
  assign n359 = n135 & n266;
  assign n360 = n81 & n112;
  assign n361 = ~n359 & ~n360;
  assign n362 = n171 & n266;
  assign n363 = n90 & n266;
  assign n364 = n176 & n266;
  assign n365 = n140 & n266;
  assign n366 = ~n364 & ~n365;
  assign n367 = ~n362 & ~n363;
  assign n368 = n366 & n367;
  assign n369 = n358 & n361;
  assign n370 = n368 & n369;
  assign n371 = n274 & n370;
  assign n372 = n306 & n371;
  assign n373 = n353 & n372;
  assign n374 = n84 & n88;
  assign n375 = n107 & n140;
  assign n376 = n90 & n110;
  assign n377 = ~n375 & ~n376;
  assign n378 = n132 & n206;
  assign n379 = n97 & n102;
  assign n380 = ~n378 & ~n379;
  assign n381 = n88 & n140;
  assign n382 = n107 & n124;
  assign n383 = ~n381 & ~n382;
  assign n384 = n110 & n181;
  assign n385 = n84 & n110;
  assign n386 = ~n384 & ~n385;
  assign n387 = n94 & n138;
  assign n388 = n81 & n108;
  assign n389 = n102 & n138;
  assign n390 = n88 & n176;
  assign n391 = n88 & n132;
  assign n392 = ~n390 & ~n391;
  assign n393 = ~n389 & n392;
  assign n394 = ~n374 & ~n387;
  assign n395 = ~n388 & n394;
  assign n396 = n377 & n380;
  assign n397 = n383 & n386;
  assign n398 = n396 & n397;
  assign n399 = n393 & n395;
  assign n400 = n398 & n399;
  assign n401 = n81 & n97;
  assign n402 = n102 & n143;
  assign n403 = ~n401 & ~n402;
  assign n404 = n81 & n135;
  assign n405 = n81 & n140;
  assign n406 = n81 & n124;
  assign n407 = n81 & n138;
  assign n408 = ~n406 & ~n407;
  assign n409 = ~n405 & n408;
  assign n410 = n403 & ~n404;
  assign n411 = n198 & n410;
  assign n412 = n205 & n409;
  assign n413 = n411 & n412;
  assign n414 = n191 & n413;
  assign n415 = n233 & n400;
  assign n416 = n414 & n415;
  assign n417 = n161 & n264;
  assign n418 = n416 & n417;
  assign n419 = n373 & n418;
  assign n420 = n138 & n206;
  assign n421 = n117 & n206;
  assign n422 = n84 & n206;
  assign n423 = ~n421 & ~n422;
  assign n424 = n181 & n206;
  assign n425 = n108 & n206;
  assign n426 = n135 & n206;
  assign n427 = n140 & n206;
  assign n428 = ~n426 & ~n427;
  assign n429 = ~n420 & ~n424;
  assign n430 = ~n425 & n429;
  assign n431 = n423 & n428;
  assign n432 = n430 & n431;
  assign n433 = ~n235 & ~n240;
  assign n434 = ~n238 & n433;
  assign n435 = ~n311 & n434;
  assign n436 = ~n98 & ~n387;
  assign n437 = ~n139 & n309;
  assign n438 = n137 & ~n141;
  assign n439 = ~n109 & ~n375;
  assign n440 = ~n354 & n436;
  assign n441 = n439 & n440;
  assign n442 = n437 & n438;
  assign n443 = n441 & n442;
  assign n444 = n87 & n106;
  assign n445 = n171 & n444;
  assign n446 = n100 & n444;
  assign n447 = n102 & n176;
  assign n448 = n84 & n444;
  assign n449 = ~n91 & ~n374;
  assign n450 = ~n103 & ~n379;
  assign n451 = n449 & n450;
  assign n452 = ~n381 & ~n402;
  assign n453 = n198 & n452;
  assign n454 = n393 & n451;
  assign n455 = n453 & n454;
  assign n456 = n152 & n455;
  assign n457 = ~n447 & ~n448;
  assign n458 = n456 & n457;
  assign n459 = n97 & n444;
  assign n460 = n138 & n444;
  assign n461 = ~n459 & ~n460;
  assign n462 = n143 & n444;
  assign n463 = n135 & n444;
  assign n464 = ~n462 & ~n463;
  assign n465 = n108 & n444;
  assign n466 = n124 & n444;
  assign n467 = n90 & n444;
  assign n468 = ~n466 & ~n467;
  assign n469 = n100 & n206;
  assign n470 = n132 & n444;
  assign n471 = ~n469 & ~n470;
  assign n472 = n176 & n444;
  assign n473 = n143 & n206;
  assign n474 = ~n472 & ~n473;
  assign n475 = n464 & ~n465;
  assign n476 = n468 & n471;
  assign n477 = n474 & n476;
  assign n478 = n475 & n477;
  assign n479 = n117 & n444;
  assign n480 = n181 & n444;
  assign n481 = ~n479 & ~n480;
  assign n482 = n140 & n444;
  assign n483 = n112 & n444;
  assign n484 = ~n482 & ~n483;
  assign n485 = n461 & n484;
  assign n486 = n481 & n485;
  assign n487 = n478 & n486;
  assign n488 = ~n445 & ~n446;
  assign n489 = n191 & n488;
  assign n490 = n487 & n489;
  assign n491 = n458 & n490;
  assign n492 = n124 & n206;
  assign n493 = ~n310 & ~n382;
  assign n494 = n112 & n206;
  assign n495 = n97 & n206;
  assign n496 = n90 & n206;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~n239 & ~n492;
  assign n499 = ~n494 & n498;
  assign n500 = n493 & n497;
  assign n501 = n499 & n500;
  assign n502 = n432 & n501;
  assign n503 = n435 & n502;
  assign n504 = n443 & n503;
  assign n505 = n491 & n504;
  assign n506 = n419 & ~n505;
  assign n507 = ~n419 & n505;
  assign n508 = ~n506 & ~n507;
  assign n509 = n108 & n130;
  assign n510 = n124 & n130;
  assign n511 = n130 & n135;
  assign n512 = n130 & n138;
  assign n513 = n84 & n130;
  assign n514 = n130 & n140;
  assign n515 = ~n510 & ~n511;
  assign n516 = ~n512 & ~n513;
  assign n517 = ~n514 & n516;
  assign n518 = n515 & n517;
  assign n519 = ~n509 & n518;
  assign n520 = ~n133 & ~n376;
  assign n521 = n117 & n130;
  assign n522 = n130 & n181;
  assign n523 = ~n521 & ~n522;
  assign n524 = ~n131 & ~n492;
  assign n525 = ~n113 & ~n234;
  assign n526 = ~n378 & n525;
  assign n527 = n386 & n497;
  assign n528 = n520 & n523;
  assign n529 = n524 & n528;
  assign n530 = n526 & n527;
  assign n531 = n529 & n530;
  assign n532 = n432 & n531;
  assign n533 = n233 & n532;
  assign n534 = ~n494 & n533;
  assign n535 = n519 & n534;
  assign n536 = n100 & n107;
  assign n537 = ~n354 & ~n536;
  assign n538 = n130 & n176;
  assign n539 = n130 & n132;
  assign n540 = ~n538 & ~n539;
  assign n541 = n107 & n117;
  assign n542 = n84 & n107;
  assign n543 = n107 & n112;
  assign n544 = n130 & n171;
  assign n545 = n90 & n130;
  assign n546 = n107 & n181;
  assign n547 = ~n544 & ~n545;
  assign n548 = ~n546 & n547;
  assign n549 = ~n541 & ~n542;
  assign n550 = ~n543 & n549;
  assign n551 = n540 & n550;
  assign n552 = n548 & n551;
  assign n553 = n107 & n143;
  assign n554 = n97 & n130;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~n239 & ~n311;
  assign n557 = n439 & n556;
  assign n558 = n493 & n537;
  assign n559 = n555 & n558;
  assign n560 = n437 & n557;
  assign n561 = n559 & n560;
  assign n562 = n552 & n561;
  assign n563 = n535 & n562;
  assign n564 = pi31  & n115;
  assign n565 = ~n80 & ~n87;
  assign n566 = pi31  & ~n565;
  assign n567 = n80 & n101;
  assign n568 = n176 & n567;
  assign n569 = n94 & n181;
  assign n570 = n94 & n112;
  assign n571 = n94 & n117;
  assign n572 = n94 & n100;
  assign n573 = ~n571 & ~n572;
  assign n574 = n84 & n94;
  assign n575 = ~n570 & ~n574;
  assign n576 = n573 & n575;
  assign n577 = n94 & n124;
  assign n578 = n94 & n143;
  assign n579 = n80 & n106;
  assign n580 = n112 & n579;
  assign n581 = ~n578 & ~n580;
  assign n582 = n84 & n579;
  assign n583 = n176 & n579;
  assign n584 = n97 & n579;
  assign n585 = n90 & n579;
  assign n586 = ~n584 & ~n585;
  assign n587 = n181 & n579;
  assign n588 = n143 & n579;
  assign n589 = ~n587 & ~n588;
  assign n590 = n135 & n579;
  assign n591 = n171 & n579;
  assign n592 = ~n590 & ~n591;
  assign n593 = n589 & n592;
  assign n594 = n117 & n579;
  assign n595 = n124 & n579;
  assign n596 = ~n594 & ~n595;
  assign n597 = n108 & n579;
  assign n598 = n140 & n579;
  assign n599 = n132 & n579;
  assign n600 = ~n598 & ~n599;
  assign n601 = n100 & n579;
  assign n602 = n138 & n579;
  assign n603 = ~n601 & ~n602;
  assign n604 = ~n582 & ~n583;
  assign n605 = ~n597 & n604;
  assign n606 = n581 & n586;
  assign n607 = n596 & n600;
  assign n608 = n603 & n607;
  assign n609 = n605 & n606;
  assign n610 = n593 & n609;
  assign n611 = n608 & n610;
  assign n612 = ~n569 & ~n577;
  assign n613 = n576 & n612;
  assign n614 = n611 & n613;
  assign n615 = n434 & n436;
  assign n616 = n438 & n615;
  assign n617 = n614 & n616;
  assign n618 = n491 & n617;
  assign n619 = ~n509 & ~n568;
  assign n620 = n562 & n619;
  assign n621 = n618 & n620;
  assign n622 = ~n219 & ~n448;
  assign n623 = ~n210 & ~n445;
  assign n624 = ~n145 & ~n222;
  assign n625 = ~n131 & ~n133;
  assign n626 = ~n172 & ~n179;
  assign n627 = ~n379 & ~n446;
  assign n628 = ~n447 & n627;
  assign n629 = n625 & n626;
  assign n630 = n214 & n624;
  assign n631 = n629 & n630;
  assign n632 = n628 & n631;
  assign n633 = n217 & ~n376;
  assign n634 = n523 & n622;
  assign n635 = n623 & n634;
  assign n636 = n633 & n635;
  assign n637 = n632 & n636;
  assign n638 = n487 & n637;
  assign n639 = n80 & n86;
  assign n640 = n117 & n639;
  assign n641 = n143 & n639;
  assign n642 = n84 & n639;
  assign n643 = ~n641 & ~n642;
  assign n644 = n112 & n639;
  assign n645 = n181 & n639;
  assign n646 = n140 & n639;
  assign n647 = ~n645 & ~n646;
  assign n648 = n108 & n639;
  assign n649 = n81 & n132;
  assign n650 = n138 & n639;
  assign n651 = n100 & n639;
  assign n652 = ~n644 & ~n648;
  assign n653 = ~n649 & ~n650;
  assign n654 = ~n651 & n653;
  assign n655 = n647 & n652;
  assign n656 = n654 & n655;
  assign n657 = ~n640 & n643;
  assign n658 = n656 & n657;
  assign n659 = n171 & n639;
  assign n660 = ~n404 & ~n659;
  assign n661 = n90 & n639;
  assign n662 = n97 & n639;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~n92 & ~n401;
  assign n665 = n124 & n639;
  assign n666 = n81 & n176;
  assign n667 = n132 & n567;
  assign n668 = ~n666 & ~n667;
  assign n669 = ~n665 & n668;
  assign n670 = n108 & n567;
  assign n671 = n140 & n567;
  assign n672 = ~n670 & ~n671;
  assign n673 = n100 & n567;
  assign n674 = n138 & n567;
  assign n675 = n143 & n567;
  assign n676 = n117 & n567;
  assign n677 = ~n675 & ~n676;
  assign n678 = ~n674 & n677;
  assign n679 = n181 & n567;
  assign n680 = n84 & n567;
  assign n681 = n90 & n567;
  assign n682 = n112 & n567;
  assign n683 = n97 & n567;
  assign n684 = ~n681 & ~n682;
  assign n685 = ~n683 & n684;
  assign n686 = n135 & n567;
  assign n687 = n176 & n639;
  assign n688 = ~n686 & ~n687;
  assign n689 = n132 & n639;
  assign n690 = n124 & n567;
  assign n691 = ~n673 & ~n679;
  assign n692 = ~n680 & ~n689;
  assign n693 = ~n690 & n692;
  assign n694 = n672 & n691;
  assign n695 = n688 & n694;
  assign n696 = n678 & n693;
  assign n697 = n685 & n696;
  assign n698 = n695 & n697;
  assign n699 = ~n388 & n409;
  assign n700 = n81 & n171;
  assign n701 = n135 & n639;
  assign n702 = n171 & n567;
  assign n703 = ~n85 & ~n702;
  assign n704 = ~n700 & ~n701;
  assign n705 = n660 & n704;
  assign n706 = n663 & n664;
  assign n707 = n703 & n706;
  assign n708 = n669 & n705;
  assign n709 = n707 & n708;
  assign n710 = n699 & n709;
  assign n711 = n658 & n710;
  assign n712 = n698 & n711;
  assign n713 = ~n236 & n260;
  assign n714 = ~n239 & n713;
  assign n715 = n373 & n714;
  assign n716 = n712 & n715;
  assign n717 = ~n122 & ~n180;
  assign n718 = n194 & n717;
  assign n719 = ~n118 & ~n147;
  assign n720 = ~n163 & ~n175;
  assign n721 = ~n389 & n720;
  assign n722 = n439 & n719;
  assign n723 = n721 & n722;
  assign n724 = n718 & n723;
  assign n725 = n166 & ~n234;
  assign n726 = n518 & n725;
  assign n727 = n724 & n726;
  assign n728 = n638 & n727;
  assign n729 = n716 & n728;
  assign n730 = ~n621 & ~n729;
  assign n731 = ~n173 & ~n404;
  assign n732 = ~n667 & ~n702;
  assign n733 = ~n310 & ~n536;
  assign n734 = ~n460 & ~n511;
  assign n735 = ~n701 & n734;
  assign n736 = n226 & n735;
  assign n737 = ~n183 & ~n480;
  assign n738 = ~n512 & ~n662;
  assign n739 = ~n91 & ~n381;
  assign n740 = ~n168 & ~n207;
  assign n741 = ~n209 & ~n659;
  assign n742 = ~n182 & ~n459;
  assign n743 = ~n448 & ~n479;
  assign n744 = ~n196 & ~n514;
  assign n745 = ~n120 & ~n221;
  assign n746 = ~n385 & ~n466;
  assign n747 = ~n666 & ~n700;
  assign n748 = n746 & n747;
  assign n749 = n737 & n745;
  assign n750 = n738 & n739;
  assign n751 = n740 & n741;
  assign n752 = n742 & n743;
  assign n753 = n744 & n752;
  assign n754 = n750 & n751;
  assign n755 = n748 & n749;
  assign n756 = n754 & n755;
  assign n757 = n753 & n756;
  assign n758 = ~n374 & ~n665;
  assign n759 = ~n167 & ~n384;
  assign n760 = ~n463 & ~n482;
  assign n761 = ~n378 & ~n465;
  assign n762 = ~n513 & ~n661;
  assign n763 = n761 & n762;
  assign n764 = n760 & n763;
  assign n765 = ~n125 & ~n218;
  assign n766 = ~n162 & ~n195;
  assign n767 = n765 & n766;
  assign n768 = ~n113 & ~n126;
  assign n769 = ~n445 & ~n467;
  assign n770 = ~n510 & n769;
  assign n771 = n150 & n768;
  assign n772 = n758 & n759;
  assign n773 = n771 & n772;
  assign n774 = n205 & n770;
  assign n775 = n767 & n774;
  assign n776 = n736 & n773;
  assign n777 = n764 & n776;
  assign n778 = n658 & n775;
  assign n779 = n777 & n778;
  assign n780 = n757 & n779;
  assign n781 = ~n144 & ~n542;
  assign n782 = ~n541 & ~n546;
  assign n783 = ~n177 & ~n382;
  assign n784 = ~n543 & n783;
  assign n785 = n474 & n781;
  assign n786 = n782 & n785;
  assign n787 = n784 & n786;
  assign n788 = n699 & n787;
  assign n789 = ~n92 & ~n103;
  assign n790 = ~n139 & ~n210;
  assign n791 = n789 & n790;
  assign n792 = n392 & n403;
  assign n793 = n471 & n523;
  assign n794 = n731 & n732;
  assign n795 = n733 & n794;
  assign n796 = n792 & n793;
  assign n797 = n791 & n796;
  assign n798 = n435 & n795;
  assign n799 = n797 & n798;
  assign n800 = n698 & n799;
  assign n801 = n788 & n800;
  assign n802 = n780 & n801;
  assign n803 = ~n729 & ~n802;
  assign n804 = ~n335 & ~n427;
  assign n805 = ~n149 & ~n168;
  assign n806 = ~n195 & ~n425;
  assign n807 = ~n599 & n806;
  assign n808 = n739 & n805;
  assign n809 = n804 & n808;
  assign n810 = n807 & n809;
  assign n811 = ~n360 & ~n473;
  assign n812 = ~n514 & ~n674;
  assign n813 = ~n173 & n314;
  assign n814 = n811 & n812;
  assign n815 = n813 & n814;
  assign n816 = ~n224 & ~n363;
  assign n817 = n436 & ~n679;
  assign n818 = ~n269 & ~n323;
  assign n819 = n573 & n818;
  assign n820 = n816 & n819;
  assign n821 = n817 & n820;
  assign n822 = ~n459 & ~n675;
  assign n823 = n357 & ~n673;
  assign n824 = ~n120 & ~n671;
  assign n825 = ~n334 & ~n390;
  assign n826 = n824 & n825;
  assign n827 = n204 & ~n391;
  assign n828 = ~n445 & ~n542;
  assign n829 = n827 & n828;
  assign n830 = ~n141 & ~n225;
  assign n831 = ~n342 & ~n472;
  assign n832 = ~n689 & n831;
  assign n833 = n822 & n830;
  assign n834 = n832 & n833;
  assign n835 = n823 & n826;
  assign n836 = n834 & n835;
  assign n837 = n815 & n829;
  assign n838 = n836 & n837;
  assign n839 = n821 & n838;
  assign n840 = ~n103 & ~n577;
  assign n841 = ~n320 & ~n687;
  assign n842 = ~n139 & ~n364;
  assign n843 = ~n270 & ~n271;
  assign n844 = ~n402 & ~n583;
  assign n845 = n843 & n844;
  assign n846 = n841 & n842;
  assign n847 = n845 & n846;
  assign n848 = ~n324 & ~n569;
  assign n849 = ~n126 & ~n321;
  assign n850 = ~n265 & ~n382;
  assign n851 = n849 & n850;
  assign n852 = n685 & n851;
  assign n853 = ~n336 & ~n670;
  assign n854 = ~n578 & ~n680;
  assign n855 = ~n200 & ~n267;
  assign n856 = ~n512 & n855;
  assign n857 = ~n318 & ~n574;
  assign n858 = ~n359 & ~n362;
  assign n859 = ~n467 & n858;
  assign n860 = n854 & n857;
  assign n861 = n859 & n860;
  assign n862 = n856 & n861;
  assign n863 = ~n199 & ~n511;
  assign n864 = ~n570 & ~n659;
  assign n865 = ~n676 & n863;
  assign n866 = n864 & n865;
  assign n867 = n862 & n866;
  assign n868 = ~n339 & ~n365;
  assign n869 = ~n510 & ~n686;
  assign n870 = ~n690 & n869;
  assign n871 = n137 & n868;
  assign n872 = n386 & n471;
  assign n873 = n765 & n840;
  assign n874 = n848 & n853;
  assign n875 = n873 & n874;
  assign n876 = n871 & n872;
  assign n877 = n870 & n876;
  assign n878 = n847 & n875;
  assign n879 = n852 & n878;
  assign n880 = n877 & n879;
  assign n881 = n867 & n880;
  assign n882 = ~n483 & ~n538;
  assign n883 = ~n208 & ~n426;
  assign n884 = ~n553 & n883;
  assign n885 = ~n354 & ~n539;
  assign n886 = ~n85 & ~n183;
  assign n887 = ~n319 & ~n462;
  assign n888 = n886 & n887;
  assign n889 = n309 & n497;
  assign n890 = n732 & n882;
  assign n891 = n885 & n890;
  assign n892 = n888 & n889;
  assign n893 = n884 & n892;
  assign n894 = n891 & n893;
  assign n895 = n632 & n810;
  assign n896 = n894 & n895;
  assign n897 = n839 & n896;
  assign n898 = n881 & n897;
  assign n899 = ~n802 & ~n898;
  assign n900 = ~n279 & ~n391;
  assign n901 = ~n648 & n900;
  assign n902 = ~n282 & ~n288;
  assign n903 = ~n308 & n902;
  assign n904 = ~n202 & ~n374;
  assign n905 = ~n209 & ~n289;
  assign n906 = ~n382 & ~n420;
  assign n907 = n905 & n906;
  assign n908 = n663 & n904;
  assign n909 = n907 & n908;
  assign n910 = n901 & n903;
  assign n911 = n909 & n910;
  assign n912 = ~n376 & ~n465;
  assign n913 = ~n196 & ~n492;
  assign n914 = ~n113 & ~n182;
  assign n915 = ~n574 & n914;
  assign n916 = n464 & n912;
  assign n917 = n913 & n916;
  assign n918 = n915 & n917;
  assign n919 = ~n286 & ~n513;
  assign n920 = ~n285 & ~n402;
  assign n921 = ~n422 & ~n446;
  assign n922 = ~n522 & ~n541;
  assign n923 = ~n126 & ~n482;
  assign n924 = ~n340 & ~n514;
  assign n925 = ~n338 & ~n598;
  assign n926 = ~n203 & ~n364;
  assign n927 = ~n387 & ~n602;
  assign n928 = ~n208 & ~n591;
  assign n929 = ~n495 & ~n686;
  assign n930 = ~n356 & ~n375;
  assign n931 = ~n109 & ~n644;
  assign n932 = ~n283 & ~n389;
  assign n933 = ~n553 & ~n640;
  assign n934 = n932 & n933;
  assign n935 = n672 & n930;
  assign n936 = n931 & n935;
  assign n937 = n934 & n936;
  assign n938 = ~n326 & ~n665;
  assign n939 = ~n300 & ~n460;
  assign n940 = ~n343 & ~n597;
  assign n941 = ~n162 & ~n311;
  assign n942 = ~n642 & n941;
  assign n943 = ~n511 & ~n584;
  assign n944 = ~n674 & n882;
  assign n945 = n943 & n944;
  assign n946 = ~n276 & ~n646;
  assign n947 = ~n193 & ~n496;
  assign n948 = n142 & ~n327;
  assign n949 = ~n131 & ~n690;
  assign n950 = n946 & n949;
  assign n951 = n947 & n950;
  assign n952 = n948 & n951;
  assign n953 = ~n355 & ~n362;
  assign n954 = ~n650 & n953;
  assign n955 = n811 & n954;
  assign n956 = ~n98 & ~n136;
  assign n957 = ~n175 & ~n585;
  assign n958 = n956 & n957;
  assign n959 = n816 & n938;
  assign n960 = n939 & n940;
  assign n961 = n959 & n960;
  assign n962 = n942 & n958;
  assign n963 = n961 & n962;
  assign n964 = n945 & n955;
  assign n965 = n963 & n964;
  assign n966 = n952 & n965;
  assign n967 = ~n590 & ~n683;
  assign n968 = ~n645 & n967;
  assign n969 = ~n681 & ~n701;
  assign n970 = n765 & n969;
  assign n971 = ~n134 & ~n472;
  assign n972 = n166 & n971;
  assign n973 = n214 & n317;
  assign n974 = n471 & n924;
  assign n975 = n925 & n926;
  assign n976 = n927 & n928;
  assign n977 = n929 & n976;
  assign n978 = n974 & n975;
  assign n979 = n968 & n973;
  assign n980 = n970 & n972;
  assign n981 = n979 & n980;
  assign n982 = n977 & n978;
  assign n983 = n274 & n982;
  assign n984 = n937 & n981;
  assign n985 = n983 & n984;
  assign n986 = n966 & n985;
  assign n987 = ~n215 & ~n297;
  assign n988 = ~n307 & n987;
  assign n989 = n840 & n988;
  assign n990 = ~n85 & ~n120;
  assign n991 = ~n167 & ~n173;
  assign n992 = ~n390 & ~n447;
  assign n993 = n991 & n992;
  assign n994 = n201 & n990;
  assign n995 = n732 & n919;
  assign n996 = n920 & n921;
  assign n997 = n922 & n923;
  assign n998 = n996 & n997;
  assign n999 = n994 & n995;
  assign n1000 = n548 & n993;
  assign n1001 = n999 & n1000;
  assign n1002 = n989 & n998;
  assign n1003 = n1001 & n1002;
  assign n1004 = n911 & n918;
  assign n1005 = n1003 & n1004;
  assign n1006 = n986 & n1005;
  assign n1007 = ~n898 & ~n1006;
  assign n1008 = ~n271 & ~n492;
  assign n1009 = ~n587 & ~n673;
  assign n1010 = n1008 & n1009;
  assign n1011 = ~n595 & ~n680;
  assign n1012 = ~n164 & ~n338;
  assign n1013 = n1011 & n1012;
  assign n1014 = ~n290 & ~n342;
  assign n1015 = ~n374 & ~n582;
  assign n1016 = ~n307 & ~n514;
  assign n1017 = ~n270 & ~n326;
  assign n1018 = ~n376 & n1017;
  assign n1019 = n1016 & n1018;
  assign n1020 = ~n182 & ~n315;
  assign n1021 = ~n199 & ~n483;
  assign n1022 = ~n648 & n1021;
  assign n1023 = ~n162 & ~n224;
  assign n1024 = ~n445 & ~n543;
  assign n1025 = ~n591 & n1024;
  assign n1026 = n1023 & n1025;
  assign n1027 = ~n280 & ~n402;
  assign n1028 = ~n594 & n1027;
  assign n1029 = n361 & n738;
  assign n1030 = n1014 & n1015;
  assign n1031 = n1020 & n1030;
  assign n1032 = n1028 & n1029;
  assign n1033 = n1022 & n1032;
  assign n1034 = n1019 & n1031;
  assign n1035 = n1026 & n1034;
  assign n1036 = n1033 & n1035;
  assign n1037 = ~n571 & ~n661;
  assign n1038 = ~n682 & ~n700;
  assign n1039 = n1037 & n1038;
  assign n1040 = n555 & n1039;
  assign n1041 = ~n334 & ~n355;
  assign n1042 = ~n195 & ~n265;
  assign n1043 = ~n385 & ~n667;
  assign n1044 = ~n207 & ~n251;
  assign n1045 = ~n365 & n1044;
  assign n1046 = ~n221 & ~n421;
  assign n1047 = ~n469 & ~n521;
  assign n1048 = ~n679 & n1047;
  assign n1049 = n1042 & n1046;
  assign n1050 = n1043 & n1049;
  assign n1051 = n1045 & n1048;
  assign n1052 = n1050 & n1051;
  assign n1053 = n194 & ~n277;
  assign n1054 = ~n203 & ~n425;
  assign n1055 = n622 & n1054;
  assign n1056 = ~n208 & ~n321;
  assign n1057 = ~n327 & ~n339;
  assign n1058 = ~n420 & ~n546;
  assign n1059 = ~n584 & ~n676;
  assign n1060 = ~n702 & n1059;
  assign n1061 = n1057 & n1058;
  assign n1062 = n1041 & n1056;
  assign n1063 = n1061 & n1062;
  assign n1064 = n1053 & n1060;
  assign n1065 = n1055 & n1064;
  assign n1066 = n1040 & n1063;
  assign n1067 = n1065 & n1066;
  assign n1068 = n1052 & n1067;
  assign n1069 = ~n316 & ~n390;
  assign n1070 = ~n482 & ~n651;
  assign n1071 = ~n200 & ~n299;
  assign n1072 = ~n513 & ~n542;
  assign n1073 = ~n544 & ~n650;
  assign n1074 = n1072 & n1073;
  assign n1075 = n969 & n1071;
  assign n1076 = n1074 & n1075;
  assign n1077 = ~n473 & ~n570;
  assign n1078 = ~n465 & ~n649;
  assign n1079 = n468 & ~n666;
  assign n1080 = n1077 & n1078;
  assign n1081 = n1079 & n1080;
  assign n1082 = ~n296 & ~n446;
  assign n1083 = ~n172 & ~n424;
  assign n1084 = ~n569 & n1083;
  assign n1085 = ~n283 & ~n340;
  assign n1086 = ~n202 & ~n646;
  assign n1087 = ~n312 & ~n318;
  assign n1088 = ~n343 & ~n641;
  assign n1089 = n1087 & n1088;
  assign n1090 = n1085 & n1086;
  assign n1091 = n1089 & n1090;
  assign n1092 = n1084 & n1091;
  assign n1093 = ~n177 & ~n287;
  assign n1094 = ~n496 & ~n585;
  assign n1095 = ~n683 & n1094;
  assign n1096 = n1069 & n1093;
  assign n1097 = n1070 & n1082;
  assign n1098 = n1096 & n1097;
  assign n1099 = n1010 & n1095;
  assign n1100 = n1013 & n1099;
  assign n1101 = n1076 & n1098;
  assign n1102 = n1081 & n1101;
  assign n1103 = n1092 & n1100;
  assign n1104 = n1102 & n1103;
  assign n1105 = n161 & n1104;
  assign n1106 = n1036 & n1068;
  assign n1107 = n1105 & n1106;
  assign n1108 = ~n1006 & ~n1107;
  assign n1109 = ~n287 & ~n591;
  assign n1110 = ~n213 & ~n354;
  assign n1111 = n1109 & n1110;
  assign n1112 = ~n445 & ~n544;
  assign n1113 = ~n424 & ~n546;
  assign n1114 = ~n163 & ~n250;
  assign n1115 = ~n253 & ~n702;
  assign n1116 = ~n245 & ~n290;
  assign n1117 = ~n312 & ~n381;
  assign n1118 = ~n365 & ~n651;
  assign n1119 = ~n131 & ~n271;
  assign n1120 = ~n355 & n1119;
  assign n1121 = ~n362 & ~n641;
  assign n1122 = ~n149 & ~n648;
  assign n1123 = n1121 & n1122;
  assign n1124 = ~n543 & ~n679;
  assign n1125 = ~n134 & ~n687;
  assign n1126 = ~n144 & ~n210;
  assign n1127 = ~n296 & ~n402;
  assign n1128 = ~n509 & n1127;
  assign n1129 = n1124 & n1126;
  assign n1130 = n1125 & n1129;
  assign n1131 = n1128 & n1130;
  assign n1132 = ~n202 & ~n388;
  assign n1133 = ~n469 & n1132;
  assign n1134 = n523 & n848;
  assign n1135 = n1112 & n1113;
  assign n1136 = n1114 & n1115;
  assign n1137 = n1116 & n1117;
  assign n1138 = n1118 & n1137;
  assign n1139 = n1135 & n1136;
  assign n1140 = n1133 & n1134;
  assign n1141 = n1111 & n1120;
  assign n1142 = n1123 & n1141;
  assign n1143 = n1139 & n1140;
  assign n1144 = n1138 & n1143;
  assign n1145 = n1131 & n1142;
  assign n1146 = n1144 & n1145;
  assign n1147 = ~n162 & ~n539;
  assign n1148 = ~n179 & ~n199;
  assign n1149 = ~n126 & ~n661;
  assign n1150 = ~n103 & ~n364;
  assign n1151 = ~n420 & n1150;
  assign n1152 = ~n282 & ~n510;
  assign n1153 = n436 & n1152;
  assign n1154 = ~n242 & ~n288;
  assign n1155 = ~n680 & n1154;
  assign n1156 = ~n465 & ~n662;
  assign n1157 = ~n238 & ~n642;
  assign n1158 = n940 & n1016;
  assign n1159 = ~n209 & ~n494;
  assign n1160 = ~n125 & ~n466;
  assign n1161 = ~n164 & ~n300;
  assign n1162 = ~n91 & ~n145;
  assign n1163 = ~n356 & ~n427;
  assign n1164 = ~n675 & n1163;
  assign n1165 = n217 & n1162;
  assign n1166 = n1159 & n1160;
  assign n1167 = n1161 & n1166;
  assign n1168 = n1164 & n1165;
  assign n1169 = n1167 & n1168;
  assign n1170 = ~n165 & ~n665;
  assign n1171 = ~n219 & ~n285;
  assign n1172 = ~n221 & ~n545;
  assign n1173 = ~n167 & ~n339;
  assign n1174 = ~n299 & ~n384;
  assign n1175 = ~n147 & ~n595;
  assign n1176 = ~n315 & ~n401;
  assign n1177 = ~n120 & ~n203;
  assign n1178 = ~n582 & n1177;
  assign n1179 = n464 & n853;
  assign n1180 = n1175 & n1176;
  assign n1181 = n1179 & n1180;
  assign n1182 = n1178 & n1181;
  assign n1183 = ~n359 & ~n601;
  assign n1184 = n241 & n1183;
  assign n1185 = n1157 & n1170;
  assign n1186 = n1171 & n1172;
  assign n1187 = n1173 & n1174;
  assign n1188 = n1186 & n1187;
  assign n1189 = n1184 & n1185;
  assign n1190 = n1158 & n1189;
  assign n1191 = n1188 & n1190;
  assign n1192 = n1169 & n1182;
  assign n1193 = n1191 & n1192;
  assign n1194 = ~n109 & ~n541;
  assign n1195 = ~n666 & n1194;
  assign n1196 = n1043 & n1156;
  assign n1197 = n1195 & n1196;
  assign n1198 = n1153 & n1155;
  assign n1199 = n1197 & n1198;
  assign n1200 = n1193 & n1199;
  assign n1201 = ~n320 & ~n480;
  assign n1202 = n581 & n1201;
  assign n1203 = ~n254 & ~n511;
  assign n1204 = ~n425 & ~n572;
  assign n1205 = n1203 & n1204;
  assign n1206 = ~n208 & ~n513;
  assign n1207 = ~n686 & n1206;
  assign n1208 = ~n472 & ~n483;
  assign n1209 = ~n389 & ~n512;
  assign n1210 = ~n139 & ~n391;
  assign n1211 = ~n671 & n1210;
  assign n1212 = n1208 & n1209;
  assign n1213 = n1211 & n1212;
  assign n1214 = ~n85 & ~n276;
  assign n1215 = ~n310 & ~n326;
  assign n1216 = n1214 & n1215;
  assign n1217 = ~n148 & ~n280;
  assign n1218 = ~n554 & n1217;
  assign n1219 = n925 & n1147;
  assign n1220 = n1148 & n1149;
  assign n1221 = n1219 & n1220;
  assign n1222 = n1151 & n1218;
  assign n1223 = n1202 & n1205;
  assign n1224 = n1207 & n1216;
  assign n1225 = n1223 & n1224;
  assign n1226 = n1221 & n1222;
  assign n1227 = n1213 & n1226;
  assign n1228 = n1225 & n1227;
  assign n1229 = n1146 & n1228;
  assign n1230 = n1200 & n1229;
  assign n1231 = ~n1107 & ~n1230;
  assign n1232 = ~n180 & ~n676;
  assign n1233 = ~n495 & ~n569;
  assign n1234 = ~n379 & ~n597;
  assign n1235 = n1232 & n1234;
  assign n1236 = n1233 & n1235;
  assign n1237 = ~n340 & ~n675;
  assign n1238 = ~n254 & ~n469;
  assign n1239 = n1237 & n1238;
  assign n1240 = ~n163 & ~n318;
  assign n1241 = ~n326 & ~n651;
  assign n1242 = ~n286 & ~n662;
  assign n1243 = ~n85 & ~n210;
  assign n1244 = n383 & n1242;
  assign n1245 = n1243 & n1244;
  assign n1246 = ~n244 & ~n539;
  assign n1247 = ~n580 & ~n665;
  assign n1248 = ~n404 & ~n473;
  assign n1249 = ~n577 & n1248;
  assign n1250 = ~n164 & ~n240;
  assign n1251 = n325 & n1250;
  assign n1252 = n449 & n760;
  assign n1253 = n1172 & n1240;
  assign n1254 = n1241 & n1246;
  assign n1255 = n1247 & n1254;
  assign n1256 = n1252 & n1253;
  assign n1257 = n593 & n1251;
  assign n1258 = n1239 & n1249;
  assign n1259 = n1257 & n1258;
  assign n1260 = n1255 & n1256;
  assign n1261 = n1245 & n1260;
  assign n1262 = n1259 & n1261;
  assign n1263 = ~n242 & ~n300;
  assign n1264 = ~n118 & ~n236;
  assign n1265 = ~n661 & n1264;
  assign n1266 = ~n177 & ~n583;
  assign n1267 = ~n546 & ~n674;
  assign n1268 = ~n203 & ~n235;
  assign n1269 = ~n113 & ~n253;
  assign n1270 = n1268 & n1269;
  assign n1271 = ~n98 & ~n196;
  assign n1272 = ~n218 & ~n267;
  assign n1273 = ~n640 & ~n680;
  assign n1274 = n1272 & n1273;
  assign n1275 = n1266 & n1271;
  assign n1276 = n1267 & n1275;
  assign n1277 = n1270 & n1274;
  assign n1278 = n1276 & n1277;
  assign n1279 = ~n216 & ~n426;
  assign n1280 = ~n183 & ~n459;
  assign n1281 = ~n179 & ~n585;
  assign n1282 = ~n378 & ~n689;
  assign n1283 = ~n165 & ~n376;
  assign n1284 = ~n239 & ~n321;
  assign n1285 = ~n544 & n1284;
  assign n1286 = n1283 & n1285;
  assign n1287 = ~n199 & ~n422;
  assign n1288 = ~n424 & ~n595;
  assign n1289 = ~n646 & ~n670;
  assign n1290 = n1288 & n1289;
  assign n1291 = n1263 & n1287;
  assign n1292 = n1279 & n1280;
  assign n1293 = n1281 & n1282;
  assign n1294 = n1292 & n1293;
  assign n1295 = n1290 & n1291;
  assign n1296 = n1265 & n1295;
  assign n1297 = n1286 & n1294;
  assign n1298 = n1296 & n1297;
  assign n1299 = n1278 & n1298;
  assign n1300 = ~n405 & ~n427;
  assign n1301 = ~n280 & ~n363;
  assign n1302 = ~n172 & ~n465;
  assign n1303 = ~n131 & n537;
  assign n1304 = n1301 & n1302;
  assign n1305 = n1303 & n1304;
  assign n1306 = ~n125 & ~n200;
  assign n1307 = ~n103 & ~n297;
  assign n1308 = n361 & n1307;
  assign n1309 = ~n649 & ~n681;
  assign n1310 = n366 & n1309;
  assign n1311 = ~n310 & ~n391;
  assign n1312 = ~n213 & ~n243;
  assign n1313 = ~n311 & ~n667;
  assign n1314 = ~n141 & ~n460;
  assign n1315 = ~n313 & ~n384;
  assign n1316 = n1314 & n1315;
  assign n1317 = ~n173 & ~n316;
  assign n1318 = n1311 & n1317;
  assign n1319 = n1312 & n1313;
  assign n1320 = n1318 & n1319;
  assign n1321 = n1316 & n1320;
  assign n1322 = ~n148 & ~n193;
  assign n1323 = ~n222 & ~n299;
  assign n1324 = ~n645 & n1323;
  assign n1325 = n278 & n1322;
  assign n1326 = n573 & n1176;
  assign n1327 = n1300 & n1306;
  assign n1328 = n1326 & n1327;
  assign n1329 = n1324 & n1325;
  assign n1330 = n1308 & n1310;
  assign n1331 = n1329 & n1330;
  assign n1332 = n1236 & n1328;
  assign n1333 = n1305 & n1332;
  assign n1334 = n1321 & n1331;
  assign n1335 = n1333 & n1334;
  assign n1336 = n1262 & n1335;
  assign n1337 = n1299 & n1336;
  assign n1338 = ~n1230 & ~n1337;
  assign n1339 = ~n134 & ~n641;
  assign n1340 = ~n165 & ~n308;
  assign n1341 = ~n335 & n1340;
  assign n1342 = ~n239 & ~n465;
  assign n1343 = ~n254 & ~n387;
  assign n1344 = ~n269 & ~n483;
  assign n1345 = n969 & n1344;
  assign n1346 = ~n243 & ~n300;
  assign n1347 = ~n479 & ~n659;
  assign n1348 = ~n480 & n1347;
  assign n1349 = ~n585 & ~n645;
  assign n1350 = ~n364 & ~n376;
  assign n1351 = ~n133 & n1349;
  assign n1352 = n1350 & n1351;
  assign n1353 = n1348 & n1352;
  assign n1354 = ~n310 & ~n582;
  assign n1355 = ~n183 & ~n588;
  assign n1356 = ~n313 & ~n462;
  assign n1357 = ~n167 & ~n509;
  assign n1358 = ~n145 & ~n363;
  assign n1359 = ~n218 & n1069;
  assign n1360 = ~n384 & ~n472;
  assign n1361 = ~n577 & n1360;
  assign n1362 = n930 & n940;
  assign n1363 = n967 & n1086;
  assign n1364 = n1246 & n1282;
  assign n1365 = n1354 & n1355;
  assign n1366 = n1356 & n1357;
  assign n1367 = n1358 & n1366;
  assign n1368 = n1364 & n1365;
  assign n1369 = n1362 & n1363;
  assign n1370 = n1359 & n1361;
  assign n1371 = n1369 & n1370;
  assign n1372 = n1367 & n1368;
  assign n1373 = n1371 & n1372;
  assign n1374 = ~n224 & ~n247;
  assign n1375 = ~n148 & ~n311;
  assign n1376 = ~n297 & ~n598;
  assign n1377 = n596 & n1160;
  assign n1378 = n1376 & n1377;
  assign n1379 = ~n253 & ~n459;
  assign n1380 = ~n91 & ~n289;
  assign n1381 = n104 & n1380;
  assign n1382 = ~n162 & ~n213;
  assign n1383 = ~n568 & ~n602;
  assign n1384 = ~n280 & ~n670;
  assign n1385 = ~n200 & ~n388;
  assign n1386 = n1379 & n1385;
  assign n1387 = n1382 & n1383;
  assign n1388 = n1384 & n1387;
  assign n1389 = n1381 & n1386;
  assign n1390 = n1388 & n1389;
  assign n1391 = ~n147 & ~n651;
  assign n1392 = ~n324 & ~n422;
  assign n1393 = ~n180 & ~n470;
  assign n1394 = ~n315 & ~n447;
  assign n1395 = ~n570 & ~n587;
  assign n1396 = ~n290 & n1395;
  assign n1397 = ~n240 & ~n288;
  assign n1398 = ~n250 & ~n407;
  assign n1399 = ~n580 & ~n671;
  assign n1400 = ~n320 & ~n572;
  assign n1401 = ~n601 & n1400;
  assign n1402 = n922 & n1300;
  assign n1403 = n1391 & n1392;
  assign n1404 = n1393 & n1394;
  assign n1405 = n1397 & n1398;
  assign n1406 = n1399 & n1405;
  assign n1407 = n1403 & n1404;
  assign n1408 = n1401 & n1402;
  assign n1409 = n1396 & n1408;
  assign n1410 = n1406 & n1407;
  assign n1411 = n1409 & n1410;
  assign n1412 = ~n446 & n1339;
  assign n1413 = n1342 & n1343;
  assign n1414 = n1346 & n1374;
  assign n1415 = n1375 & n1414;
  assign n1416 = n1412 & n1413;
  assign n1417 = n1341 & n1345;
  assign n1418 = n1416 & n1417;
  assign n1419 = n1378 & n1415;
  assign n1420 = n1418 & n1419;
  assign n1421 = n1353 & n1390;
  assign n1422 = n1420 & n1421;
  assign n1423 = n1373 & n1411;
  assign n1424 = n1422 & n1423;
  assign n1425 = n1068 & n1424;
  assign n1426 = ~n1337 & ~n1425;
  assign n1427 = ~n283 & ~n287;
  assign n1428 = ~n378 & n1427;
  assign n1429 = n731 & n1428;
  assign n1430 = n767 & n1429;
  assign n1431 = ~n299 & ~n387;
  assign n1432 = ~n401 & ~n585;
  assign n1433 = ~n288 & ~n690;
  assign n1434 = ~n375 & ~n466;
  assign n1435 = n437 & n1434;
  assign n1436 = ~n316 & ~n323;
  assign n1437 = ~n681 & n1436;
  assign n1438 = ~n265 & ~n339;
  assign n1439 = ~n473 & ~n511;
  assign n1440 = ~n541 & n1439;
  assign n1441 = n146 & n1438;
  assign n1442 = n1201 & n1301;
  assign n1443 = n1346 & n1431;
  assign n1444 = n1432 & n1433;
  assign n1445 = n1443 & n1444;
  assign n1446 = n1441 & n1442;
  assign n1447 = n451 & n1440;
  assign n1448 = n1437 & n1447;
  assign n1449 = n1445 & n1446;
  assign n1450 = n1435 & n1449;
  assign n1451 = n1430 & n1448;
  assign n1452 = n1450 & n1451;
  assign n1453 = ~n285 & n1112;
  assign n1454 = ~n382 & n1453;
  assign n1455 = ~n209 & ~n482;
  assign n1456 = ~n570 & ~n682;
  assign n1457 = ~n216 & ~n521;
  assign n1458 = ~n122 & ~n512;
  assign n1459 = ~n343 & ~n405;
  assign n1460 = ~n514 & n1459;
  assign n1461 = n1456 & n1457;
  assign n1462 = n1458 & n1461;
  assign n1463 = n1460 & n1462;
  assign n1464 = ~n539 & ~n597;
  assign n1465 = ~n313 & ~n447;
  assign n1466 = ~n175 & n537;
  assign n1467 = n1464 & n1465;
  assign n1468 = n1466 & n1467;
  assign n1469 = ~n327 & ~n542;
  assign n1470 = ~n113 & ~n648;
  assign n1471 = n166 & n1470;
  assign n1472 = ~n148 & ~n538;
  assign n1473 = ~n141 & ~n192;
  assign n1474 = ~n574 & n1473;
  assign n1475 = n1206 & n1474;
  assign n1476 = ~n335 & ~n495;
  assign n1477 = ~n510 & ~n642;
  assign n1478 = ~n661 & ~n680;
  assign n1479 = ~n683 & n1478;
  assign n1480 = n1476 & n1477;
  assign n1481 = n1117 & n1472;
  assign n1482 = n1480 & n1481;
  assign n1483 = n1479 & n1482;
  assign n1484 = n1475 & n1483;
  assign n1485 = ~n290 & ~n426;
  assign n1486 = ~n238 & ~n472;
  assign n1487 = ~n149 & ~n571;
  assign n1488 = ~n98 & ~n246;
  assign n1489 = ~n671 & n1488;
  assign n1490 = n361 & n622;
  assign n1491 = n1121 & n1469;
  assign n1492 = n1485 & n1486;
  assign n1493 = n1487 & n1492;
  assign n1494 = n1490 & n1491;
  assign n1495 = n1216 & n1489;
  assign n1496 = n1471 & n1495;
  assign n1497 = n1493 & n1494;
  assign n1498 = n1468 & n1497;
  assign n1499 = n1496 & n1498;
  assign n1500 = n1484 & n1499;
  assign n1501 = ~n126 & n555;
  assign n1502 = ~n183 & ~n687;
  assign n1503 = ~n315 & ~n583;
  assign n1504 = n1502 & n1503;
  assign n1505 = ~n131 & ~n168;
  assign n1506 = ~n578 & n1505;
  assign n1507 = ~n245 & ~n644;
  assign n1508 = ~n253 & ~n649;
  assign n1509 = ~n224 & ~n319;
  assign n1510 = ~n340 & n1509;
  assign n1511 = ~n338 & ~n356;
  assign n1512 = ~n365 & ~n459;
  assign n1513 = ~n462 & ~n701;
  assign n1514 = n1512 & n1513;
  assign n1515 = n853 & n1511;
  assign n1516 = n1507 & n1508;
  assign n1517 = n1515 & n1516;
  assign n1518 = n1510 & n1514;
  assign n1519 = n1517 & n1518;
  assign n1520 = ~n202 & ~n225;
  assign n1521 = ~n240 & ~n427;
  assign n1522 = ~n584 & n1521;
  assign n1523 = n1455 & n1520;
  assign n1524 = n1522 & n1523;
  assign n1525 = n1501 & n1504;
  assign n1526 = n1506 & n1525;
  assign n1527 = n1454 & n1524;
  assign n1528 = n1526 & n1527;
  assign n1529 = n1463 & n1519;
  assign n1530 = n1528 & n1529;
  assign n1531 = n1452 & n1530;
  assign n1532 = n1500 & n1531;
  assign n1533 = ~n1425 & ~n1532;
  assign n1534 = ~n243 & ~n405;
  assign n1535 = ~n144 & ~n251;
  assign n1536 = ~n665 & ~n667;
  assign n1537 = ~n267 & ~n285;
  assign n1538 = ~n118 & ~n599;
  assign n1539 = ~n336 & ~n355;
  assign n1540 = n1233 & n1539;
  assign n1541 = ~n402 & ~n446;
  assign n1542 = ~n288 & ~n469;
  assign n1543 = ~n374 & ~n670;
  assign n1544 = ~n676 & n1543;
  assign n1545 = n586 & n1541;
  assign n1546 = n1542 & n1545;
  assign n1547 = n1544 & n1546;
  assign n1548 = n322 & ~n649;
  assign n1549 = n812 & n863;
  assign n1550 = n1534 & n1535;
  assign n1551 = n1536 & n1537;
  assign n1552 = n1538 & n1551;
  assign n1553 = n1549 & n1550;
  assign n1554 = n1540 & n1548;
  assign n1555 = n1553 & n1554;
  assign n1556 = n1552 & n1555;
  assign n1557 = n1547 & n1556;
  assign n1558 = ~n359 & ~n385;
  assign n1559 = ~n276 & ~n578;
  assign n1560 = ~n208 & ~n544;
  assign n1561 = ~n313 & ~n680;
  assign n1562 = ~n179 & ~n536;
  assign n1563 = ~n235 & ~n279;
  assign n1564 = ~n598 & ~n642;
  assign n1565 = n1563 & n1564;
  assign n1566 = n1561 & n1562;
  assign n1567 = n1565 & n1566;
  assign n1568 = ~n173 & ~n270;
  assign n1569 = ~n463 & ~n513;
  assign n1570 = ~n590 & n1569;
  assign n1571 = n1568 & n1570;
  assign n1572 = ~n323 & ~n388;
  assign n1573 = ~n542 & n1572;
  assign n1574 = n493 & n913;
  assign n1575 = n1347 & n1486;
  assign n1576 = n1558 & n1559;
  assign n1577 = n1560 & n1576;
  assign n1578 = n1574 & n1575;
  assign n1579 = n1573 & n1578;
  assign n1580 = n1567 & n1577;
  assign n1581 = n1571 & n1580;
  assign n1582 = n1579 & n1581;
  assign n1583 = ~n407 & n1374;
  assign n1584 = n573 & n1115;
  assign n1585 = ~n113 & ~n139;
  assign n1586 = ~n360 & n1585;
  assign n1587 = ~n318 & ~n425;
  assign n1588 = ~n225 & ~n365;
  assign n1589 = ~n483 & ~n645;
  assign n1590 = n1588 & n1589;
  assign n1591 = n1114 & n1587;
  assign n1592 = n1590 & n1591;
  assign n1593 = ~n420 & ~n671;
  assign n1594 = ~n496 & ~n700;
  assign n1595 = ~n289 & ~n602;
  assign n1596 = ~n200 & ~n234;
  assign n1597 = ~n287 & n1596;
  assign n1598 = n194 & n1149;
  assign n1599 = n1382 & n1593;
  assign n1600 = n1594 & n1595;
  assign n1601 = n1599 & n1600;
  assign n1602 = n1597 & n1598;
  assign n1603 = n1583 & n1584;
  assign n1604 = n1586 & n1603;
  assign n1605 = n1601 & n1602;
  assign n1606 = n1592 & n1605;
  assign n1607 = n1169 & n1604;
  assign n1608 = n1606 & n1607;
  assign n1609 = n1557 & n1608;
  assign n1610 = n1582 & n1609;
  assign n1611 = ~n1532 & ~n1610;
  assign n1612 = ~n463 & ~n674;
  assign n1613 = ~n402 & n1612;
  assign n1614 = ~n582 & ~n676;
  assign n1615 = ~n321 & ~n362;
  assign n1616 = ~n196 & ~n265;
  assign n1617 = ~n599 & n1616;
  assign n1618 = ~n165 & ~n250;
  assign n1619 = ~n427 & ~n578;
  assign n1620 = n1618 & n1619;
  assign n1621 = n919 & n1614;
  assign n1622 = n1615 & n1621;
  assign n1623 = n1613 & n1620;
  assign n1624 = n1617 & n1623;
  assign n1625 = n1622 & n1624;
  assign n1626 = ~n583 & ~n686;
  assign n1627 = ~n509 & ~n542;
  assign n1628 = ~n224 & ~n514;
  assign n1629 = n1627 & n1628;
  assign n1630 = ~n122 & ~n287;
  assign n1631 = ~n200 & ~n690;
  assign n1632 = ~n360 & ~n522;
  assign n1633 = ~n236 & ~n364;
  assign n1634 = n169 & n1632;
  assign n1635 = n1633 & n1634;
  assign n1636 = ~n374 & ~n401;
  assign n1637 = ~n671 & ~n683;
  assign n1638 = n1636 & n1637;
  assign n1639 = n1485 & n1626;
  assign n1640 = n1630 & n1631;
  assign n1641 = n1639 & n1640;
  assign n1642 = n1249 & n1638;
  assign n1643 = n1629 & n1642;
  assign n1644 = n1635 & n1641;
  assign n1645 = n1643 & n1644;
  assign n1646 = n1625 & n1645;
  assign n1647 = ~n666 & n841;
  assign n1648 = ~n598 & ~n665;
  assign n1649 = n1647 & n1648;
  assign n1650 = ~n195 & ~n541;
  assign n1651 = ~n164 & ~n270;
  assign n1652 = ~n238 & ~n338;
  assign n1653 = ~n183 & ~n216;
  assign n1654 = ~n365 & ~n446;
  assign n1655 = n1653 & n1654;
  assign n1656 = n1085 & n1124;
  assign n1657 = n1535 & n1650;
  assign n1658 = n1651 & n1652;
  assign n1659 = n1657 & n1658;
  assign n1660 = n1655 & n1656;
  assign n1661 = n1659 & n1660;
  assign n1662 = ~n163 & ~n239;
  assign n1663 = ~n510 & ~n662;
  assign n1664 = n1662 & n1663;
  assign n1665 = n204 & n1664;
  assign n1666 = ~n225 & ~n354;
  assign n1667 = ~n139 & ~n279;
  assign n1668 = ~n134 & ~n465;
  assign n1669 = ~n173 & ~n207;
  assign n1670 = ~n448 & n1669;
  assign n1671 = ~n288 & ~n316;
  assign n1672 = ~n405 & ~n597;
  assign n1673 = n1671 & n1672;
  assign n1674 = n150 & n1666;
  assign n1675 = n1667 & n1668;
  assign n1676 = n1674 & n1675;
  assign n1677 = n1670 & n1673;
  assign n1678 = n1676 & n1677;
  assign n1679 = ~n326 & ~n339;
  assign n1680 = ~n327 & ~n539;
  assign n1681 = ~n103 & ~n382;
  assign n1682 = ~n247 & ~n334;
  assign n1683 = ~n648 & n1682;
  assign n1684 = ~n209 & ~n595;
  assign n1685 = n1679 & n1684;
  assign n1686 = n1680 & n1681;
  assign n1687 = n1685 & n1686;
  assign n1688 = n1683 & n1687;
  assign n1689 = ~n285 & ~n420;
  assign n1690 = ~n147 & ~n390;
  assign n1691 = n1501 & n1690;
  assign n1692 = ~n85 & ~n335;
  assign n1693 = ~n545 & n1692;
  assign n1694 = n1349 & n1693;
  assign n1695 = ~n242 & ~n277;
  assign n1696 = ~n421 & ~n424;
  assign n1697 = ~n574 & n1696;
  assign n1698 = n471 & n1695;
  assign n1699 = n1394 & n1689;
  assign n1700 = n1698 & n1699;
  assign n1701 = n1120 & n1697;
  assign n1702 = n1700 & n1701;
  assign n1703 = n1665 & n1691;
  assign n1704 = n1694 & n1703;
  assign n1705 = n1678 & n1702;
  assign n1706 = n1688 & n1705;
  assign n1707 = n1704 & n1706;
  assign n1708 = ~n682 & n1344;
  assign n1709 = n1347 & n1708;
  assign n1710 = ~n319 & ~n466;
  assign n1711 = ~n125 & ~n472;
  assign n1712 = ~n568 & ~n588;
  assign n1713 = ~n98 & ~n120;
  assign n1714 = ~n422 & ~n700;
  assign n1715 = ~n246 & ~n311;
  assign n1716 = ~n343 & n1715;
  assign n1717 = n643 & n1710;
  assign n1718 = n1711 & n1712;
  assign n1719 = n1713 & n1714;
  assign n1720 = n1718 & n1719;
  assign n1721 = n1716 & n1717;
  assign n1722 = n1720 & n1721;
  assign n1723 = ~n113 & ~n199;
  assign n1724 = ~n356 & ~n482;
  assign n1725 = ~n546 & ~n571;
  assign n1726 = ~n591 & ~n702;
  assign n1727 = n1725 & n1726;
  assign n1728 = n1723 & n1724;
  assign n1729 = n178 & n1209;
  assign n1730 = n1728 & n1729;
  assign n1731 = n1727 & n1730;
  assign n1732 = n1649 & n1709;
  assign n1733 = n1731 & n1732;
  assign n1734 = n1661 & n1722;
  assign n1735 = n1733 & n1734;
  assign n1736 = n1646 & n1735;
  assign n1737 = n1707 & n1736;
  assign n1738 = ~n1610 & ~n1737;
  assign n1739 = ~n177 & ~n670;
  assign n1740 = ~n405 & n1739;
  assign n1741 = ~n234 & ~n376;
  assign n1742 = ~n569 & ~n661;
  assign n1743 = n1741 & n1742;
  assign n1744 = ~n286 & ~n580;
  assign n1745 = ~n245 & ~n682;
  assign n1746 = ~n276 & ~n420;
  assign n1747 = ~n470 & ~n568;
  assign n1748 = n1746 & n1747;
  assign n1749 = n1744 & n1745;
  assign n1750 = n1748 & n1749;
  assign n1751 = n1045 & n1740;
  assign n1752 = n1743 & n1751;
  assign n1753 = n1750 & n1752;
  assign n1754 = ~n427 & ~n601;
  assign n1755 = ~n448 & n826;
  assign n1756 = ~n212 & ~n381;
  assign n1757 = n537 & ~n546;
  assign n1758 = n1756 & n1757;
  assign n1759 = n1396 & n1758;
  assign n1760 = ~n446 & ~n509;
  assign n1761 = n1508 & n1760;
  assign n1762 = ~n103 & ~n642;
  assign n1763 = n481 & n1431;
  assign n1764 = ~n482 & ~n510;
  assign n1765 = ~n213 & ~n342;
  assign n1766 = ~n209 & ~n594;
  assign n1767 = n1694 & n1766;
  assign n1768 = ~n407 & n1264;
  assign n1769 = n1314 & n1762;
  assign n1770 = n1764 & n1765;
  assign n1771 = n1769 & n1770;
  assign n1772 = n437 & n1768;
  assign n1773 = n1453 & n1761;
  assign n1774 = n1763 & n1773;
  assign n1775 = n1771 & n1772;
  assign n1776 = n1649 & n1775;
  assign n1777 = n862 & n1774;
  assign n1778 = n1767 & n1777;
  assign n1779 = n1776 & n1778;
  assign n1780 = ~n297 & ~n402;
  assign n1781 = ~n590 & n1780;
  assign n1782 = n882 & n1781;
  assign n1783 = ~n145 & ~n651;
  assign n1784 = ~n136 & ~n425;
  assign n1785 = ~n283 & ~n646;
  assign n1786 = ~n242 & ~n388;
  assign n1787 = n822 & n1784;
  assign n1788 = n1785 & n1786;
  assign n1789 = n1787 & n1788;
  assign n1790 = ~n247 & ~n336;
  assign n1791 = ~n514 & ~n595;
  assign n1792 = ~n662 & n1791;
  assign n1793 = n928 & n1790;
  assign n1794 = n1173 & n1469;
  assign n1795 = n1487 & n1754;
  assign n1796 = n1783 & n1795;
  assign n1797 = n1793 & n1794;
  assign n1798 = n1792 & n1797;
  assign n1799 = n1755 & n1796;
  assign n1800 = n1782 & n1789;
  assign n1801 = n1799 & n1800;
  assign n1802 = n1759 & n1798;
  assign n1803 = n1801 & n1802;
  assign n1804 = n1753 & n1803;
  assign n1805 = n1779 & n1804;
  assign n1806 = ~n1737 & ~n1805;
  assign n1807 = ~n355 & ~n384;
  assign n1808 = ~n196 & ~n336;
  assign n1809 = ~n92 & ~n168;
  assign n1810 = ~n212 & ~n312;
  assign n1811 = ~n376 & ~n391;
  assign n1812 = ~n402 & ~n642;
  assign n1813 = n1811 & n1812;
  assign n1814 = n1809 & n1810;
  assign n1815 = n1808 & n1814;
  assign n1816 = n1813 & n1815;
  assign n1817 = ~n601 & ~n700;
  assign n1818 = ~n126 & ~n240;
  assign n1819 = ~n290 & n1818;
  assign n1820 = n1817 & n1819;
  assign n1821 = ~n246 & ~n470;
  assign n1822 = ~n542 & ~n546;
  assign n1823 = ~n659 & ~n680;
  assign n1824 = n1822 & n1823;
  assign n1825 = n204 & n1821;
  assign n1826 = n1232 & n1300;
  assign n1827 = n1807 & n1826;
  assign n1828 = n1824 & n1825;
  assign n1829 = n1207 & n1510;
  assign n1830 = n1828 & n1829;
  assign n1831 = n1820 & n1827;
  assign n1832 = n1830 & n1831;
  assign n1833 = n1816 & n1832;
  assign n1834 = ~n221 & n523;
  assign n1835 = ~n236 & ~n321;
  assign n1836 = ~n665 & n1835;
  assign n1837 = ~n234 & ~n381;
  assign n1838 = ~n165 & ~n277;
  assign n1839 = ~n539 & n1838;
  assign n1840 = ~n207 & ~n210;
  assign n1841 = ~n269 & ~n289;
  assign n1842 = ~n554 & n1841;
  assign n1843 = n765 & n1840;
  assign n1844 = n1842 & n1843;
  assign n1845 = n1839 & n1844;
  assign n1846 = ~n103 & ~n365;
  assign n1847 = ~n469 & ~n479;
  assign n1848 = ~n496 & ~n662;
  assign n1849 = n1847 & n1848;
  assign n1850 = n201 & n1846;
  assign n1851 = n600 & n1121;
  assign n1852 = n1279 & n1356;
  assign n1853 = n1391 & n1394;
  assign n1854 = n1432 & n1837;
  assign n1855 = n1853 & n1854;
  assign n1856 = n1851 & n1852;
  assign n1857 = n1849 & n1850;
  assign n1858 = n1836 & n1857;
  assign n1859 = n1855 & n1856;
  assign n1860 = n1858 & n1859;
  assign n1861 = n1845 & n1860;
  assign n1862 = ~n671 & ~n701;
  assign n1863 = ~n243 & ~n297;
  assign n1864 = ~n342 & ~n422;
  assign n1865 = n1863 & n1864;
  assign n1866 = n931 & n1862;
  assign n1867 = n1865 & n1866;
  assign n1868 = ~n225 & ~n574;
  assign n1869 = ~n390 & ~n583;
  assign n1870 = ~n584 & n668;
  assign n1871 = n1112 & n1869;
  assign n1872 = n1870 & n1871;
  assign n1873 = ~n460 & ~n689;
  assign n1874 = ~n283 & ~n356;
  assign n1875 = ~n379 & ~n421;
  assign n1876 = ~n482 & ~n543;
  assign n1877 = n1875 & n1876;
  assign n1878 = n436 & n1874;
  assign n1879 = n1873 & n1878;
  assign n1880 = n1877 & n1879;
  assign n1881 = ~n219 & ~n299;
  assign n1882 = ~n510 & ~n675;
  assign n1883 = n1881 & n1882;
  assign n1884 = n1535 & n1760;
  assign n1885 = n1868 & n1884;
  assign n1886 = n968 & n1883;
  assign n1887 = n1834 & n1886;
  assign n1888 = n1867 & n1885;
  assign n1889 = n1872 & n1888;
  assign n1890 = n1880 & n1887;
  assign n1891 = n1889 & n1890;
  assign n1892 = n1833 & n1891;
  assign n1893 = n1861 & n1892;
  assign n1894 = ~n1805 & ~n1893;
  assign n1895 = ~n324 & ~n384;
  assign n1896 = ~n522 & n1895;
  assign n1897 = ~n162 & ~n192;
  assign n1898 = ~n208 & ~n319;
  assign n1899 = ~n545 & n1898;
  assign n1900 = n1897 & n1899;
  assign n1901 = n1896 & n1900;
  assign n1902 = ~n239 & ~n316;
  assign n1903 = ~n462 & n1902;
  assign n1904 = ~n113 & ~n553;
  assign n1905 = ~n424 & ~n590;
  assign n1906 = n1904 & n1905;
  assign n1907 = ~n246 & ~n365;
  assign n1908 = n622 & n1112;
  assign n1909 = ~n180 & ~n401;
  assign n1910 = ~n147 & ~n421;
  assign n1911 = ~n334 & ~n640;
  assign n1912 = ~n207 & ~n300;
  assign n1913 = ~n321 & ~n646;
  assign n1914 = ~n674 & n1913;
  assign n1915 = n1909 & n1912;
  assign n1916 = n1910 & n1911;
  assign n1917 = n1915 & n1916;
  assign n1918 = n1914 & n1917;
  assign n1919 = ~n175 & ~n307;
  assign n1920 = ~n682 & n1919;
  assign n1921 = n1627 & n1920;
  assign n1922 = ~n92 & ~n98;
  assign n1923 = ~n359 & n1922;
  assign n1924 = ~n136 & ~n336;
  assign n1925 = ~n521 & ~n649;
  assign n1926 = n1924 & n1925;
  assign n1927 = n1923 & n1926;
  assign n1928 = ~n91 & ~n148;
  assign n1929 = ~n165 & ~n234;
  assign n1930 = ~n282 & ~n375;
  assign n1931 = ~n472 & ~n681;
  assign n1932 = n1930 & n1931;
  assign n1933 = n1928 & n1929;
  assign n1934 = n380 & n1399;
  assign n1935 = n1907 & n1934;
  assign n1936 = n1932 & n1933;
  assign n1937 = n1908 & n1936;
  assign n1938 = n1921 & n1935;
  assign n1939 = n1927 & n1938;
  assign n1940 = n1918 & n1937;
  assign n1941 = n1939 & n1940;
  assign n1942 = ~n271 & ~n667;
  assign n1943 = ~n389 & n1942;
  assign n1944 = ~n426 & ~n673;
  assign n1945 = ~n177 & ~n215;
  assign n1946 = n174 & n1945;
  assign n1947 = ~n85 & ~n296;
  assign n1948 = ~n312 & ~n480;
  assign n1949 = ~n645 & ~n666;
  assign n1950 = n1948 & n1949;
  assign n1951 = n1507 & n1947;
  assign n1952 = n1944 & n1951;
  assign n1953 = n1943 & n1950;
  assign n1954 = n1946 & n1953;
  assign n1955 = n1952 & n1954;
  assign n1956 = ~n133 & ~n235;
  assign n1957 = n600 & n1714;
  assign n1958 = n1956 & n1957;
  assign n1959 = ~n225 & ~n356;
  assign n1960 = ~n492 & ~n680;
  assign n1961 = n1959 & n1960;
  assign n1962 = ~n126 & ~n364;
  assign n1963 = ~n463 & ~n689;
  assign n1964 = n1962 & n1963;
  assign n1965 = ~n313 & ~n425;
  assign n1966 = ~n168 & n1965;
  assign n1967 = ~n299 & ~n583;
  assign n1968 = ~n702 & n1967;
  assign n1969 = ~n141 & ~n648;
  assign n1970 = ~n182 & ~n460;
  assign n1971 = ~n221 & ~n363;
  assign n1972 = n840 & n1971;
  assign n1973 = ~n267 & ~n335;
  assign n1974 = n929 & n1973;
  assign n1975 = n1347 & n1969;
  assign n1976 = n1970 & n1975;
  assign n1977 = n1961 & n1974;
  assign n1978 = n1964 & n1966;
  assign n1979 = n1968 & n1972;
  assign n1980 = n1978 & n1979;
  assign n1981 = n1976 & n1977;
  assign n1982 = n1980 & n1981;
  assign n1983 = n1759 & n1982;
  assign n1984 = ~n122 & ~n578;
  assign n1985 = n392 & n1984;
  assign n1986 = n493 & n882;
  assign n1987 = n938 & n1712;
  assign n1988 = n1764 & n1987;
  assign n1989 = n1985 & n1986;
  assign n1990 = n1903 & n1906;
  assign n1991 = n1989 & n1990;
  assign n1992 = n1958 & n1988;
  assign n1993 = n1991 & n1992;
  assign n1994 = n1901 & n1993;
  assign n1995 = n1955 & n1994;
  assign n1996 = n1941 & n1983;
  assign n1997 = n1995 & n1996;
  assign n1998 = ~n1893 & ~n1997;
  assign n1999 = ~n91 & ~n136;
  assign n2000 = ~n323 & n1999;
  assign n2001 = ~n222 & ~n250;
  assign n2002 = n623 & n2001;
  assign n2003 = n1379 & n2002;
  assign n2004 = n2000 & n2003;
  assign n2005 = ~n215 & ~n701;
  assign n2006 = ~n661 & n882;
  assign n2007 = n1391 & n2006;
  assign n2008 = ~n312 & ~n359;
  assign n2009 = ~n594 & ~n601;
  assign n2010 = ~n139 & ~n207;
  assign n2011 = ~n235 & ~n342;
  assign n2012 = ~n469 & n2011;
  assign n2013 = n392 & n2010;
  assign n2014 = n647 & n927;
  assign n2015 = n1560 & n2005;
  assign n2016 = n2008 & n2009;
  assign n2017 = n2015 & n2016;
  assign n2018 = n2013 & n2014;
  assign n2019 = n2012 & n2018;
  assign n2020 = n1665 & n2017;
  assign n2021 = n2007 & n2020;
  assign n2022 = n1722 & n2019;
  assign n2023 = n2021 & n2022;
  assign n2024 = ~n131 & ~n218;
  assign n2025 = ~n470 & ~n521;
  assign n2026 = n2024 & n2025;
  assign n2027 = ~n279 & ~n542;
  assign n2028 = ~n572 & n2027;
  assign n2029 = ~n234 & ~n671;
  assign n2030 = n1312 & n2029;
  assign n2031 = n1539 & n2030;
  assign n2032 = ~n167 & ~n193;
  assign n2033 = ~n247 & ~n404;
  assign n2034 = ~n494 & n2033;
  assign n2035 = n943 & n2032;
  assign n2036 = n1281 & n2035;
  assign n2037 = n1839 & n2034;
  assign n2038 = n2026 & n2028;
  assign n2039 = n2037 & n2038;
  assign n2040 = n2031 & n2036;
  assign n2041 = n2039 & n2040;
  assign n2042 = n1661 & n2004;
  assign n2043 = n2041 & n2042;
  assign n2044 = n1983 & n2043;
  assign n2045 = n2023 & n2044;
  assign n2046 = ~n1997 & ~n2045;
  assign n2047 = ~n324 & ~n662;
  assign n2048 = ~n164 & ~n219;
  assign n2049 = ~n404 & ~n544;
  assign n2050 = ~n141 & ~n179;
  assign n2051 = n2048 & n2049;
  assign n2052 = n2050 & n2051;
  assign n2053 = ~n245 & ~n354;
  assign n2054 = ~n496 & n2053;
  assign n2055 = ~n213 & ~n650;
  assign n2056 = ~n118 & ~n343;
  assign n2057 = ~n577 & n2056;
  assign n2058 = n2055 & n2057;
  assign n2059 = n2054 & n2058;
  assign n2060 = ~n321 & ~n675;
  assign n2061 = ~n193 & ~n195;
  assign n2062 = ~n356 & n2061;
  assign n2063 = ~n467 & ~n666;
  assign n2064 = ~n147 & n2063;
  assign n2065 = ~n98 & ~n289;
  assign n2066 = ~n225 & ~n338;
  assign n2067 = ~n175 & n2066;
  assign n2068 = ~n327 & ~n388;
  assign n2069 = ~n390 & ~n424;
  assign n2070 = ~n514 & n2069;
  assign n2071 = n1965 & n2068;
  assign n2072 = n2065 & n2071;
  assign n2073 = n2067 & n2070;
  assign n2074 = n2072 & n2073;
  assign n2075 = ~n315 & ~n590;
  assign n2076 = ~n670 & ~n681;
  assign n2077 = n2075 & n2076;
  assign n2078 = n1689 & n2047;
  assign n2079 = n2060 & n2078;
  assign n2080 = n2062 & n2077;
  assign n2081 = n2064 & n2080;
  assign n2082 = n2052 & n2079;
  assign n2083 = n2081 & n2082;
  assign n2084 = n2059 & n2074;
  assign n2085 = n2083 & n2084;
  assign n2086 = ~n269 & ~n594;
  assign n2087 = ~n379 & ~n568;
  assign n2088 = ~n307 & ~n385;
  assign n2089 = ~n210 & ~n446;
  assign n2090 = n1300 & n2089;
  assign n2091 = n2088 & n2090;
  assign n2092 = ~n378 & ~n648;
  assign n2093 = ~n470 & ~n554;
  assign n2094 = ~n492 & n1086;
  assign n2095 = n2093 & n2094;
  assign n2096 = ~n177 & ~n308;
  assign n2097 = ~n148 & ~n473;
  assign n2098 = ~n109 & ~n122;
  assign n2099 = ~n382 & ~n509;
  assign n2100 = n2098 & n2099;
  assign n2101 = n241 & n581;
  assign n2102 = n2096 & n2097;
  assign n2103 = n2101 & n2102;
  assign n2104 = n1613 & n2100;
  assign n2105 = n1670 & n2104;
  assign n2106 = n2103 & n2105;
  assign n2107 = ~n342 & ~n602;
  assign n2108 = n1157 & n2107;
  assign n2109 = ~n212 & ~n406;
  assign n2110 = ~n649 & ~n665;
  assign n2111 = n449 & n2110;
  assign n2112 = ~n287 & ~n355;
  assign n2113 = ~n244 & ~n326;
  assign n2114 = ~n445 & ~n680;
  assign n2115 = ~n682 & n2114;
  assign n2116 = n298 & n2113;
  assign n2117 = n1354 & n1944;
  assign n2118 = n2092 & n2109;
  assign n2119 = n2112 & n2118;
  assign n2120 = n2116 & n2117;
  assign n2121 = n1396 & n2115;
  assign n2122 = n2108 & n2111;
  assign n2123 = n2121 & n2122;
  assign n2124 = n2119 & n2120;
  assign n2125 = n2091 & n2095;
  assign n2126 = n2124 & n2125;
  assign n2127 = n2123 & n2126;
  assign n2128 = n2106 & n2127;
  assign n2129 = ~n387 & ~n401;
  assign n2130 = ~n199 & ~n224;
  assign n2131 = ~n384 & n2130;
  assign n2132 = ~n276 & ~n381;
  assign n2133 = ~n479 & ~n494;
  assign n2134 = ~n553 & ~n569;
  assign n2135 = ~n700 & n2134;
  assign n2136 = n2132 & n2133;
  assign n2137 = n1160 & n1667;
  assign n2138 = n2129 & n2137;
  assign n2139 = n2135 & n2136;
  assign n2140 = n2131 & n2139;
  assign n2141 = n2138 & n2140;
  assign n2142 = ~n247 & ~n316;
  assign n2143 = ~n362 & ~n676;
  assign n2144 = n2142 & n2143;
  assign n2145 = ~n183 & ~n319;
  assign n2146 = ~n495 & ~n512;
  assign n2147 = n2145 & n2146;
  assign n2148 = n573 & n2147;
  assign n2149 = n2144 & n2148;
  assign n2150 = ~n601 & ~n644;
  assign n2151 = ~n113 & n2150;
  assign n2152 = ~n165 & ~n251;
  assign n2153 = ~n267 & ~n542;
  assign n2154 = n2152 & n2153;
  assign n2155 = n337 & n688;
  assign n2156 = n2086 & n2087;
  assign n2157 = n2155 & n2156;
  assign n2158 = n2006 & n2154;
  assign n2159 = n2151 & n2158;
  assign n2160 = n1635 & n2157;
  assign n2161 = n2159 & n2160;
  assign n2162 = n2149 & n2161;
  assign n2163 = n2141 & n2162;
  assign n2164 = n2085 & n2163;
  assign n2165 = n2128 & n2164;
  assign n2166 = ~n2045 & ~n2165;
  assign n2167 = ~n339 & ~n701;
  assign n2168 = ~n145 & ~n297;
  assign n2169 = ~n553 & n2168;
  assign n2170 = ~n316 & ~n522;
  assign n2171 = ~n299 & ~n389;
  assign n2172 = n2170 & n2171;
  assign n2173 = ~n202 & ~n342;
  assign n2174 = n386 & n2173;
  assign n2175 = n2167 & n2174;
  assign n2176 = n2169 & n2172;
  assign n2177 = n2175 & n2176;
  assign n2178 = ~n109 & ~n569;
  assign n2179 = ~n126 & ~n196;
  assign n2180 = ~n200 & ~n239;
  assign n2181 = ~n271 & ~n420;
  assign n2182 = ~n472 & ~n588;
  assign n2183 = n2181 & n2182;
  assign n2184 = n2179 & n2180;
  assign n2185 = n1263 & n1651;
  assign n2186 = n2178 & n2185;
  assign n2187 = n2183 & n2184;
  assign n2188 = n2186 & n2187;
  assign n2189 = n169 & ~n465;
  assign n2190 = ~n282 & ~n597;
  assign n2191 = ~n362 & ~n666;
  assign n2192 = ~n118 & ~n177;
  assign n2193 = ~n122 & ~n421;
  assign n2194 = ~n163 & ~n689;
  assign n2195 = ~n496 & ~n574;
  assign n2196 = n2194 & n2195;
  assign n2197 = ~n243 & ~n323;
  assign n2198 = ~n570 & n2197;
  assign n2199 = n1907 & n2192;
  assign n2200 = n2193 & n2199;
  assign n2201 = n2026 & n2198;
  assign n2202 = n2196 & n2201;
  assign n2203 = n2200 & n2202;
  assign n2204 = ~n236 & ~n245;
  assign n2205 = ~n285 & n2204;
  assign n2206 = ~n207 & ~n250;
  assign n2207 = n217 & n2206;
  assign n2208 = n1764 & n1965;
  assign n2209 = n2150 & n2190;
  assign n2210 = n2191 & n2209;
  assign n2211 = n2207 & n2208;
  assign n2212 = n678 & n1923;
  assign n2213 = n2189 & n2205;
  assign n2214 = n2212 & n2213;
  assign n2215 = n2210 & n2211;
  assign n2216 = n2214 & n2215;
  assign n2217 = n2203 & n2216;
  assign n2218 = ~n199 & n537;
  assign n2219 = n2217 & n2218;
  assign n2220 = ~n447 & ~n494;
  assign n2221 = ~n195 & ~n382;
  assign n2222 = ~n584 & n2221;
  assign n2223 = ~n335 & ~n446;
  assign n2224 = ~n492 & ~n512;
  assign n2225 = n2223 & n2224;
  assign n2226 = ~n379 & ~n650;
  assign n2227 = ~n320 & ~n587;
  assign n2228 = n1281 & n1970;
  assign n2229 = ~n340 & ~n673;
  assign n2230 = ~n193 & n2229;
  assign n2231 = ~n311 & ~n388;
  assign n2232 = ~n543 & ~n686;
  assign n2233 = n2231 & n2232;
  assign n2234 = ~n149 & ~n602;
  assign n2235 = ~n234 & ~n407;
  assign n2236 = ~n509 & ~n594;
  assign n2237 = n2235 & n2236;
  assign n2238 = n2234 & n2237;
  assign n2239 = ~n173 & ~n599;
  assign n2240 = n278 & n2239;
  assign n2241 = ~n85 & ~n402;
  assign n2242 = n214 & n2241;
  assign n2243 = n816 & n2226;
  assign n2244 = n2227 & n2243;
  assign n2245 = n2228 & n2242;
  assign n2246 = n2230 & n2233;
  assign n2247 = n2240 & n2246;
  assign n2248 = n2244 & n2245;
  assign n2249 = n1709 & n2238;
  assign n2250 = n2248 & n2249;
  assign n2251 = n2247 & n2250;
  assign n2252 = ~n120 & ~n133;
  assign n2253 = ~n319 & ~n321;
  assign n2254 = ~n401 & ~n687;
  assign n2255 = n2253 & n2254;
  assign n2256 = n1157 & n2252;
  assign n2257 = n1238 & n2220;
  assign n2258 = n2256 & n2257;
  assign n2259 = n2222 & n2255;
  assign n2260 = n2225 & n2259;
  assign n2261 = n2258 & n2260;
  assign n2262 = n2177 & n2188;
  assign n2263 = n2261 & n2262;
  assign n2264 = n2251 & n2263;
  assign n2265 = n2219 & n2264;
  assign n2266 = ~n2165 & ~n2265;
  assign n2267 = ~n200 & ~n598;
  assign n2268 = n1652 & n2267;
  assign n2269 = n464 & ~n545;
  assign n2270 = n1969 & n2269;
  assign n2271 = ~n320 & ~n578;
  assign n2272 = ~n321 & ~n375;
  assign n2273 = n174 & n2272;
  assign n2274 = ~n122 & ~n327;
  assign n2275 = ~n215 & ~n482;
  assign n2276 = ~n521 & n2275;
  assign n2277 = n2274 & n2276;
  assign n2278 = ~n144 & ~n218;
  assign n2279 = ~n289 & ~n390;
  assign n2280 = ~n511 & n2279;
  assign n2281 = n573 & n2278;
  assign n2282 = n1472 & n1679;
  assign n2283 = n2194 & n2271;
  assign n2284 = n2282 & n2283;
  assign n2285 = n2280 & n2281;
  assign n2286 = n2064 & n2268;
  assign n2287 = n2273 & n2286;
  assign n2288 = n2284 & n2285;
  assign n2289 = n2270 & n2277;
  assign n2290 = n2288 & n2289;
  assign n2291 = n2287 & n2290;
  assign n2292 = n2141 & n2291;
  assign n2293 = ~n310 & ~n642;
  assign n2294 = ~n544 & n2293;
  assign n2295 = ~n574 & n1246;
  assign n2296 = ~n162 & ~n587;
  assign n2297 = ~n85 & ~n472;
  assign n2298 = ~n307 & ~n425;
  assign n2299 = ~n183 & ~n210;
  assign n2300 = ~n378 & ~n687;
  assign n2301 = n194 & ~n354;
  assign n2302 = n967 & n2299;
  assign n2303 = n2300 & n2302;
  assign n2304 = n2301 & n2303;
  assign n2305 = ~n219 & ~n480;
  assign n2306 = ~n92 & ~n300;
  assign n2307 = ~n385 & n2306;
  assign n2308 = ~n167 & ~n312;
  assign n2309 = n1765 & n2308;
  assign n2310 = n2305 & n2309;
  assign n2311 = n2307 & n2310;
  assign n2312 = ~n271 & ~n283;
  assign n2313 = ~n510 & n2312;
  assign n2314 = ~n133 & ~n391;
  assign n2315 = ~n164 & ~n225;
  assign n2316 = ~n242 & ~n448;
  assign n2317 = ~n582 & n2316;
  assign n2318 = n1393 & n2315;
  assign n2319 = n2314 & n2318;
  assign n2320 = n2317 & n2319;
  assign n2321 = n2238 & n2320;
  assign n2322 = ~n207 & ~n675;
  assign n2323 = ~n280 & ~n445;
  assign n2324 = ~n286 & ~n334;
  assign n2325 = ~n179 & ~n577;
  assign n2326 = n433 & n2325;
  assign n2327 = n738 & n2322;
  assign n2328 = n2323 & n2324;
  assign n2329 = n2327 & n2328;
  assign n2330 = n249 & n2326;
  assign n2331 = n2313 & n2330;
  assign n2332 = n2329 & n2331;
  assign n2333 = n2311 & n2332;
  assign n2334 = n2321 & n2333;
  assign n2335 = ~n177 & ~n236;
  assign n2336 = ~n253 & ~n365;
  assign n2337 = ~n422 & ~n591;
  assign n2338 = ~n641 & ~n659;
  assign n2339 = n2337 & n2338;
  assign n2340 = n2335 & n2336;
  assign n2341 = n1358 & n1862;
  assign n2342 = n2340 & n2341;
  assign n2343 = n2339 & n2342;
  assign n2344 = ~n195 & ~n495;
  assign n2345 = n1283 & n2344;
  assign n2346 = n2226 & n2296;
  assign n2347 = n2297 & n2298;
  assign n2348 = n2346 & n2347;
  assign n2349 = n2294 & n2345;
  assign n2350 = n2295 & n2349;
  assign n2351 = n2348 & n2350;
  assign n2352 = n1547 & n2304;
  assign n2353 = n2343 & n2352;
  assign n2354 = n2351 & n2353;
  assign n2355 = n2292 & n2354;
  assign n2356 = n2334 & n2355;
  assign n2357 = ~n2265 & ~n2356;
  assign n2358 = ~n195 & ~n594;
  assign n2359 = ~n246 & ~n308;
  assign n2360 = ~n391 & ~n514;
  assign n2361 = ~n253 & ~n538;
  assign n2362 = ~n267 & ~n406;
  assign n2363 = n2360 & n2362;
  assign n2364 = n2361 & n2363;
  assign n2365 = ~n92 & ~n215;
  assign n2366 = ~n683 & ~n700;
  assign n2367 = ~n243 & ~n336;
  assign n2368 = ~n512 & ~n522;
  assign n2369 = n2367 & n2368;
  assign n2370 = n1356 & n2365;
  assign n2371 = n2366 & n2370;
  assign n2372 = n2369 & n2371;
  assign n2373 = ~n402 & ~n482;
  assign n2374 = ~n494 & ~n701;
  assign n2375 = ~n196 & n2374;
  assign n2376 = ~n98 & ~n210;
  assign n2377 = ~n238 & ~n599;
  assign n2378 = ~n602 & n2377;
  assign n2379 = n2376 & n2378;
  assign n2380 = ~n113 & ~n254;
  assign n2381 = n946 & n2380;
  assign n2382 = n1502 & n2358;
  assign n2383 = n2359 & n2373;
  assign n2384 = n2382 & n2383;
  assign n2385 = n2375 & n2381;
  assign n2386 = n2384 & n2385;
  assign n2387 = n2364 & n2379;
  assign n2388 = n2386 & n2387;
  assign n2389 = n2372 & n2388;
  assign n2390 = ~n385 & ~n568;
  assign n2391 = ~n172 & ~n539;
  assign n2392 = ~n289 & ~n384;
  assign n2393 = ~n389 & ~n642;
  assign n2394 = n2392 & n2393;
  assign n2395 = ~n213 & ~n320;
  assign n2396 = n581 & n2395;
  assign n2397 = n178 & ~n536;
  assign n2398 = ~n363 & ~n446;
  assign n2399 = ~n665 & n2398;
  assign n2400 = n624 & n928;
  assign n2401 = n943 & n2400;
  assign n2402 = n1396 & n2399;
  assign n2403 = n2397 & n2402;
  assign n2404 = n2401 & n2403;
  assign n2405 = ~n192 & ~n378;
  assign n2406 = ~n473 & n2405;
  assign n2407 = ~n244 & ~n667;
  assign n2408 = ~n671 & ~n674;
  assign n2409 = n2407 & n2408;
  assign n2410 = n433 & n1041;
  assign n2411 = n1113 & n1148;
  assign n2412 = n1344 & n1689;
  assign n2413 = n2411 & n2412;
  assign n2414 = n2409 & n2410;
  assign n2415 = n2196 & n2406;
  assign n2416 = n2414 & n2415;
  assign n2417 = n2413 & n2416;
  assign n2418 = n2404 & n2417;
  assign n2419 = ~n495 & ~n650;
  assign n2420 = ~n118 & ~n247;
  assign n2421 = ~n470 & ~n588;
  assign n2422 = n2420 & n2421;
  assign n2423 = n2419 & n2422;
  assign n2424 = ~n120 & ~n250;
  assign n2425 = ~n200 & ~n702;
  assign n2426 = ~n382 & ~n466;
  assign n2427 = ~n544 & n2426;
  assign n2428 = n298 & n1015;
  assign n2429 = n1118 & n1469;
  assign n2430 = n1711 & n2390;
  assign n2431 = n2391 & n2424;
  assign n2432 = n2425 & n2431;
  assign n2433 = n2429 & n2430;
  assign n2434 = n2427 & n2428;
  assign n2435 = n2394 & n2396;
  assign n2436 = n2434 & n2435;
  assign n2437 = n2432 & n2433;
  assign n2438 = n2423 & n2437;
  assign n2439 = n1678 & n2436;
  assign n2440 = n2438 & n2439;
  assign n2441 = n2389 & n2440;
  assign n2442 = n2418 & n2441;
  assign n2443 = ~n2356 & ~n2442;
  assign n2444 = ~n173 & ~n193;
  assign n2445 = ~n536 & n2444;
  assign n2446 = ~n406 & ~n595;
  assign n2447 = ~n659 & n2446;
  assign n2448 = n2131 & n2447;
  assign n2449 = n2445 & n2448;
  assign n2450 = ~n267 & ~n427;
  assign n2451 = ~n382 & ~n667;
  assign n2452 = ~n122 & ~n483;
  assign n2453 = ~n126 & ~n470;
  assign n2454 = n2366 & n2453;
  assign n2455 = ~n598 & ~n640;
  assign n2456 = ~n221 & ~n238;
  assign n2457 = ~n644 & n2456;
  assign n2458 = n2455 & n2457;
  assign n2459 = ~n296 & ~n365;
  assign n2460 = ~n388 & ~n680;
  assign n2461 = n2459 & n2460;
  assign n2462 = n252 & n939;
  assign n2463 = n1394 & n2450;
  assign n2464 = n2451 & n2452;
  assign n2465 = n2463 & n2464;
  assign n2466 = n2461 & n2462;
  assign n2467 = n2172 & n2454;
  assign n2468 = n2466 & n2467;
  assign n2469 = n764 & n2465;
  assign n2470 = n2458 & n2469;
  assign n2471 = n2468 & n2470;
  assign n2472 = ~n139 & ~n426;
  assign n2473 = ~n541 & ~n597;
  assign n2474 = ~n404 & ~n574;
  assign n2475 = ~n133 & ~n240;
  assign n2476 = ~n265 & n1159;
  assign n2477 = n1745 & n2476;
  assign n2478 = ~n141 & ~n216;
  assign n2479 = ~n446 & n2478;
  assign n2480 = ~n85 & ~n254;
  assign n2481 = ~n234 & ~n379;
  assign n2482 = ~n510 & ~n545;
  assign n2483 = ~n570 & ~n701;
  assign n2484 = n2482 & n2483;
  assign n2485 = n1756 & n2481;
  assign n2486 = n2480 & n2485;
  assign n2487 = n1647 & n2484;
  assign n2488 = n2294 & n2479;
  assign n2489 = n2487 & n2488;
  assign n2490 = n2486 & n2489;
  assign n2491 = ~n308 & ~n334;
  assign n2492 = ~n134 & n2491;
  assign n2493 = ~n356 & ~n645;
  assign n2494 = ~n149 & ~n288;
  assign n2495 = n2493 & n2494;
  assign n2496 = ~n91 & ~n244;
  assign n2497 = ~n311 & ~n679;
  assign n2498 = n2496 & n2497;
  assign n2499 = n1713 & n2474;
  assign n2500 = n2475 & n2499;
  assign n2501 = n2492 & n2498;
  assign n2502 = n2495 & n2501;
  assign n2503 = n2477 & n2500;
  assign n2504 = n2502 & n2503;
  assign n2505 = n1092 & n2504;
  assign n2506 = n2490 & n2505;
  assign n2507 = ~n203 & ~n242;
  assign n2508 = ~n327 & ~n448;
  assign n2509 = ~n584 & n2508;
  assign n2510 = n1904 & n2507;
  assign n2511 = n2060 & n2472;
  assign n2512 = n2473 & n2511;
  assign n2513 = n2509 & n2510;
  assign n2514 = n2512 & n2513;
  assign n2515 = n2506 & n2514;
  assign n2516 = ~n271 & ~n290;
  assign n2517 = ~n196 & ~n208;
  assign n2518 = ~n235 & ~n543;
  assign n2519 = n2517 & n2518;
  assign n2520 = n2516 & n2519;
  assign n2521 = ~n136 & ~n648;
  assign n2522 = n497 & ~n601;
  assign n2523 = ~n131 & ~n336;
  assign n2524 = ~n459 & ~n469;
  assign n2525 = ~n473 & ~n585;
  assign n2526 = n2524 & n2525;
  assign n2527 = n573 & n589;
  assign n2528 = n927 & n1593;
  assign n2529 = n1710 & n2521;
  assign n2530 = n2523 & n2529;
  assign n2531 = n2527 & n2528;
  assign n2532 = n2522 & n2526;
  assign n2533 = n2531 & n2532;
  assign n2534 = n2520 & n2530;
  assign n2535 = n2533 & n2534;
  assign n2536 = n2449 & n2535;
  assign n2537 = n2471 & n2536;
  assign n2538 = n2515 & n2537;
  assign n2539 = ~n2442 & ~n2538;
  assign n2540 = ~n378 & ~n645;
  assign n2541 = ~n467 & ~n571;
  assign n2542 = ~n287 & ~n297;
  assign n2543 = ~n134 & ~n283;
  assign n2544 = ~n320 & n2543;
  assign n2545 = n2542 & n2544;
  assign n2546 = ~n118 & ~n538;
  assign n2547 = ~n670 & n2546;
  assign n2548 = ~n362 & ~n509;
  assign n2549 = n555 & n2548;
  assign n2550 = n765 & n1263;
  assign n2551 = n1313 & n1457;
  assign n2552 = n2540 & n2541;
  assign n2553 = n2551 & n2552;
  assign n2554 = n2549 & n2550;
  assign n2555 = n2547 & n2554;
  assign n2556 = n2545 & n2553;
  assign n2557 = n2555 & n2556;
  assign n2558 = n1816 & n2557;
  assign n2559 = ~n149 & ~n335;
  assign n2560 = ~n407 & n2559;
  assign n2561 = ~n277 & ~n316;
  assign n2562 = ~n472 & ~n674;
  assign n2563 = n2561 & n2562;
  assign n2564 = n2521 & n2563;
  assign n2565 = ~n296 & ~n315;
  assign n2566 = ~n120 & ~n426;
  assign n2567 = ~n98 & ~n148;
  assign n2568 = ~n282 & ~n343;
  assign n2569 = ~n379 & ~n445;
  assign n2570 = ~n511 & n2569;
  assign n2571 = n2567 & n2568;
  assign n2572 = n1149 & n2475;
  assign n2573 = n2565 & n2566;
  assign n2574 = n2572 & n2573;
  assign n2575 = n2570 & n2571;
  assign n2576 = n2574 & n2575;
  assign n2577 = ~n215 & ~n359;
  assign n2578 = ~n595 & ~n676;
  assign n2579 = n2577 & n2578;
  assign n2580 = n842 & n931;
  assign n2581 = n2579 & n2580;
  assign n2582 = ~n122 & ~n193;
  assign n2583 = ~n285 & ~n602;
  assign n2584 = ~n666 & ~n686;
  assign n2585 = n2583 & n2584;
  assign n2586 = n731 & n2582;
  assign n2587 = n743 & n1077;
  assign n2588 = n1113 & n1237;
  assign n2589 = n1632 & n2588;
  assign n2590 = n2586 & n2587;
  assign n2591 = n2585 & n2590;
  assign n2592 = n2581 & n2589;
  assign n2593 = n2591 & n2592;
  assign n2594 = n2576 & n2593;
  assign n2595 = ~n199 & ~n514;
  assign n2596 = n2594 & n2595;
  assign n2597 = ~n299 & ~n323;
  assign n2598 = ~n213 & ~n326;
  assign n2599 = ~n163 & ~n682;
  assign n2600 = n223 & ~n496;
  assign n2601 = n1764 & n2516;
  assign n2602 = n2597 & n2598;
  assign n2603 = n2599 & n2602;
  assign n2604 = n2600 & n2601;
  assign n2605 = n823 & n2604;
  assign n2606 = n2603 & n2605;
  assign n2607 = ~n244 & ~n324;
  assign n2608 = ~n470 & ~n584;
  assign n2609 = n2607 & n2608;
  assign n2610 = n237 & n449;
  assign n2611 = n464 & n967;
  assign n2612 = n1508 & n1712;
  assign n2613 = n1869 & n2612;
  assign n2614 = n2610 & n2611;
  assign n2615 = n2560 & n2609;
  assign n2616 = n2614 & n2615;
  assign n2617 = n1305 & n2613;
  assign n2618 = n2564 & n2617;
  assign n2619 = n2616 & n2618;
  assign n2620 = n2606 & n2619;
  assign n2621 = n2558 & n2620;
  assign n2622 = n2596 & n2621;
  assign n2623 = ~n2538 & ~n2622;
  assign n2624 = ~n286 & ~n342;
  assign n2625 = ~n541 & ~n588;
  assign n2626 = n2624 & n2625;
  assign n2627 = ~n120 & ~n310;
  assign n2628 = ~n480 & n2627;
  assign n2629 = n2626 & n2628;
  assign n2630 = ~n270 & ~n683;
  assign n2631 = ~n339 & n1536;
  assign n2632 = n2630 & n2631;
  assign n2633 = ~n389 & ~n649;
  assign n2634 = ~n421 & ~n536;
  assign n2635 = ~n239 & n2092;
  assign n2636 = n2190 & n2633;
  assign n2637 = n2634 & n2636;
  assign n2638 = n2635 & n2637;
  assign n2639 = ~n375 & ~n645;
  assign n2640 = ~n192 & ~n244;
  assign n2641 = n2639 & n2640;
  assign n2642 = ~n448 & ~n462;
  assign n2643 = ~n690 & n2642;
  assign n2644 = ~n242 & ~n359;
  assign n2645 = ~n673 & n2644;
  assign n2646 = n1118 & n1240;
  assign n2647 = n2296 & n2646;
  assign n2648 = n2492 & n2645;
  assign n2649 = n2641 & n2643;
  assign n2650 = n2648 & n2649;
  assign n2651 = n2629 & n2647;
  assign n2652 = n2632 & n2651;
  assign n2653 = n2004 & n2650;
  assign n2654 = n2638 & n2653;
  assign n2655 = n2652 & n2654;
  assign n2656 = n1833 & n2085;
  assign n2657 = n2655 & n2656;
  assign n2658 = ~n2622 & ~n2657;
  assign n2659 = ~n222 & ~n422;
  assign n2660 = ~n269 & ~n543;
  assign n2661 = ~n172 & ~n356;
  assign n2662 = ~n376 & n2661;
  assign n2663 = ~n276 & ~n680;
  assign n2664 = ~n311 & n1300;
  assign n2665 = n2663 & n2664;
  assign n2666 = ~n287 & ~n674;
  assign n2667 = n1280 & n2666;
  assign n2668 = n1783 & n2194;
  assign n2669 = n2297 & n2392;
  assign n2670 = n2668 & n2669;
  assign n2671 = n2667 & n2670;
  assign n2672 = n2665 & n2671;
  assign n2673 = ~n247 & ~n342;
  assign n2674 = ~n646 & n2673;
  assign n2675 = ~n387 & ~n572;
  assign n2676 = n309 & n2675;
  assign n2677 = n1311 & n1837;
  assign n2678 = n1868 & n2659;
  assign n2679 = n2660 & n2678;
  assign n2680 = n2676 & n2677;
  assign n2681 = n1010 & n2662;
  assign n2682 = n2674 & n2681;
  assign n2683 = n2679 & n2680;
  assign n2684 = n2682 & n2683;
  assign n2685 = n2672 & n2684;
  assign n2686 = ~n286 & ~n640;
  assign n2687 = ~n133 & ~n180;
  assign n2688 = ~n202 & ~n390;
  assign n2689 = ~n545 & ~n591;
  assign n2690 = ~n602 & n2689;
  assign n2691 = n2687 & n2688;
  assign n2692 = n2686 & n2691;
  assign n2693 = n2690 & n2692;
  assign n2694 = ~n495 & ~n687;
  assign n2695 = ~n216 & ~n364;
  assign n2696 = n1068 & n2695;
  assign n2697 = n1433 & n2008;
  assign n2698 = ~n144 & ~n245;
  assign n2699 = ~n335 & ~n466;
  assign n2700 = ~n665 & n2699;
  assign n2701 = n178 & n2698;
  assign n2702 = n1764 & n2701;
  assign n2703 = n1022 & n2700;
  assign n2704 = n2697 & n2703;
  assign n2705 = n2702 & n2704;
  assign n2706 = ~n379 & ~n601;
  assign n2707 = n298 & ~n465;
  assign n2708 = n1121 & n2707;
  assign n2709 = ~n246 & ~n462;
  assign n2710 = ~n509 & ~n511;
  assign n2711 = ~n577 & ~n683;
  assign n2712 = n2710 & n2711;
  assign n2713 = n325 & n2709;
  assign n2714 = n765 & n920;
  assign n2715 = n1015 & n1562;
  assign n2716 = n1786 & n2694;
  assign n2717 = n2706 & n2716;
  assign n2718 = n2714 & n2715;
  assign n2719 = n2712 & n2713;
  assign n2720 = n2718 & n2719;
  assign n2721 = n2708 & n2717;
  assign n2722 = n2720 & n2721;
  assign n2723 = n2693 & n2722;
  assign n2724 = n2705 & n2723;
  assign n2725 = n2685 & n2724;
  assign n2726 = n2696 & n2725;
  assign n2727 = ~n2657 & ~n2726;
  assign n2728 = ~n339 & ~n401;
  assign n2729 = ~n148 & ~n595;
  assign n2730 = n2728 & n2729;
  assign n2731 = ~n311 & n600;
  assign n2732 = n1384 & n2731;
  assign n2733 = n93 & ~n354;
  assign n2734 = n174 & n423;
  assign n2735 = n2733 & n2734;
  assign n2736 = ~n381 & ~n554;
  assign n2737 = ~n538 & ~n572;
  assign n2738 = ~n542 & ~n641;
  assign n2739 = ~n165 & ~n203;
  assign n2740 = n2738 & n2739;
  assign n2741 = ~n113 & ~n118;
  assign n2742 = ~n445 & n2741;
  assign n2743 = n1156 & n1172;
  assign n2744 = n1232 & n2060;
  assign n2745 = n2063 & n2480;
  assign n2746 = n2736 & n2737;
  assign n2747 = n2745 & n2746;
  assign n2748 = n2743 & n2744;
  assign n2749 = n1437 & n2742;
  assign n2750 = n2740 & n2749;
  assign n2751 = n2747 & n2748;
  assign n2752 = n2477 & n2751;
  assign n2753 = n2750 & n2752;
  assign n2754 = ~n202 & ~n673;
  assign n2755 = ~n482 & ~n553;
  assign n2756 = ~n234 & ~n644;
  assign n2757 = ~n679 & n2756;
  assign n2758 = ~n182 & ~n296;
  assign n2759 = n1357 & n2758;
  assign n2760 = n1650 & n1784;
  assign n2761 = n2754 & n2755;
  assign n2762 = n2760 & n2761;
  assign n2763 = n2643 & n2759;
  assign n2764 = n2757 & n2763;
  assign n2765 = n2762 & n2764;
  assign n2766 = ~n164 & ~n243;
  assign n2767 = ~n277 & ~n343;
  assign n2768 = ~n578 & ~n582;
  assign n2769 = n2767 & n2768;
  assign n2770 = n471 & n2766;
  assign n2771 = n2008 & n2542;
  assign n2772 = n2694 & n2771;
  assign n2773 = n2769 & n2770;
  assign n2774 = n2730 & n2773;
  assign n2775 = n1019 & n2772;
  assign n2776 = n2732 & n2735;
  assign n2777 = n2775 & n2776;
  assign n2778 = n2774 & n2777;
  assign n2779 = n2765 & n2778;
  assign n2780 = n2418 & n2753;
  assign n2781 = n2779 & n2780;
  assign n2782 = ~n2726 & ~n2781;
  assign n2783 = ~n235 & ~n376;
  assign n2784 = ~n641 & n1969;
  assign n2785 = ~n239 & ~n320;
  assign n2786 = ~n144 & ~n311;
  assign n2787 = ~n299 & ~n521;
  assign n2788 = ~n209 & ~n469;
  assign n2789 = ~n676 & n2788;
  assign n2790 = n1125 & n1267;
  assign n2791 = n2107 & n2785;
  assign n2792 = n2786 & n2787;
  assign n2793 = n2791 & n2792;
  assign n2794 = n2789 & n2790;
  assign n2795 = n2784 & n2794;
  assign n2796 = n2793 & n2795;
  assign n2797 = ~n244 & ~n277;
  assign n2798 = ~n270 & ~n280;
  assign n2799 = ~n385 & ~n407;
  assign n2800 = ~n522 & ~n675;
  assign n2801 = ~n680 & ~n681;
  assign n2802 = n2800 & n2801;
  assign n2803 = n2798 & n2799;
  assign n2804 = n2802 & n2803;
  assign n2805 = ~n327 & ~n640;
  assign n2806 = n1970 & n2805;
  assign n2807 = ~n318 & n1109;
  assign n2808 = n1172 & n1176;
  assign n2809 = n1346 & n1808;
  assign n2810 = n1907 & n2634;
  assign n2811 = n2797 & n2810;
  assign n2812 = n2808 & n2809;
  assign n2813 = n2394 & n2807;
  assign n2814 = n2806 & n2813;
  assign n2815 = n2811 & n2812;
  assign n2816 = n2804 & n2815;
  assign n2817 = n2814 & n2816;
  assign n2818 = ~n323 & ~n402;
  assign n2819 = ~n541 & ~n644;
  assign n2820 = n2818 & n2819;
  assign n2821 = n1681 & n2820;
  assign n2822 = ~n276 & ~n312;
  assign n2823 = ~n338 & n765;
  assign n2824 = ~n172 & ~n288;
  assign n2825 = n268 & n2824;
  assign n2826 = ~n482 & ~n580;
  assign n2827 = ~n597 & n2826;
  assign n2828 = n298 & n2097;
  assign n2829 = n2827 & n2828;
  assign n2830 = ~n584 & ~n700;
  assign n2831 = ~n569 & ~n587;
  assign n2832 = ~n286 & n1667;
  assign n2833 = ~n98 & ~n208;
  assign n2834 = ~n375 & ~n512;
  assign n2835 = n2833 & n2834;
  assign n2836 = n1149 & n2830;
  assign n2837 = n2831 & n2836;
  assign n2838 = n2832 & n2835;
  assign n2839 = n2837 & n2838;
  assign n2840 = ~n359 & ~n494;
  assign n2841 = ~n583 & n2840;
  assign n2842 = n380 & n929;
  assign n2843 = n1054 & n1615;
  assign n2844 = n2842 & n2843;
  assign n2845 = n823 & n2841;
  assign n2846 = n1740 & n2823;
  assign n2847 = n2825 & n2846;
  assign n2848 = n2844 & n2845;
  assign n2849 = n2829 & n2848;
  assign n2850 = n2839 & n2847;
  assign n2851 = n2849 & n2850;
  assign n2852 = ~n404 & ~n445;
  assign n2853 = n93 & n2852;
  assign n2854 = n284 & n596;
  assign n2855 = n1344 & n1487;
  assign n2856 = n2425 & n2491;
  assign n2857 = n2783 & n2822;
  assign n2858 = n2856 & n2857;
  assign n2859 = n2854 & n2855;
  assign n2860 = n2853 & n2859;
  assign n2861 = n2095 & n2858;
  assign n2862 = n2821 & n2861;
  assign n2863 = n2860 & n2862;
  assign n2864 = n2796 & n2863;
  assign n2865 = n2817 & n2851;
  assign n2866 = n2864 & n2865;
  assign n2867 = ~n2781 & ~n2866;
  assign n2868 = ~n269 & ~n640;
  assign n2869 = n268 & n2868;
  assign n2870 = ~n312 & ~n661;
  assign n2871 = ~n406 & ~n546;
  assign n2872 = ~n686 & n1380;
  assign n2873 = n1711 & n1970;
  assign n2874 = n2226 & n2870;
  assign n2875 = n2871 & n2874;
  assign n2876 = n2872 & n2873;
  assign n2877 = n2869 & n2876;
  assign n2878 = n2052 & n2875;
  assign n2879 = n2629 & n2878;
  assign n2880 = n2877 & n2879;
  assign n2881 = n211 & ~n326;
  assign n2882 = n596 & n2881;
  assign n2883 = ~n144 & ~n287;
  assign n2884 = ~n514 & n2883;
  assign n2885 = ~n251 & n1041;
  assign n2886 = n2641 & n2885;
  assign n2887 = n204 & n840;
  assign n2888 = n1714 & n2887;
  assign n2889 = ~n427 & ~n591;
  assign n2890 = n1301 & n2889;
  assign n2891 = n1469 & n2092;
  assign n2892 = n2480 & n2891;
  assign n2893 = n2884 & n2890;
  assign n2894 = n2892 & n2893;
  assign n2895 = n1571 & n1691;
  assign n2896 = n2882 & n2886;
  assign n2897 = n2888 & n2896;
  assign n2898 = n2894 & n2895;
  assign n2899 = n2897 & n2898;
  assign n2900 = n2880 & n2899;
  assign n2901 = n2219 & n2900;
  assign n2902 = ~n2866 & ~n2901;
  assign n2903 = ~n494 & ~n512;
  assign n2904 = ~n125 & ~n584;
  assign n2905 = n2903 & n2904;
  assign n2906 = ~n221 & ~n297;
  assign n2907 = ~n360 & ~n511;
  assign n2908 = n2906 & n2907;
  assign n2909 = ~n362 & ~n682;
  assign n2910 = ~n271 & n520;
  assign n2911 = n1241 & n1666;
  assign n2912 = n2909 & n2911;
  assign n2913 = n2674 & n2910;
  assign n2914 = n2912 & n2913;
  assign n2915 = ~n335 & ~n541;
  assign n2916 = ~n594 & ~n686;
  assign n2917 = n2915 & n2916;
  assign n2918 = n1174 & n1587;
  assign n2919 = n1680 & n2785;
  assign n2920 = n2918 & n2919;
  assign n2921 = n2917 & n2920;
  assign n2922 = n1927 & n2921;
  assign n2923 = ~n131 & ~n300;
  assign n2924 = n278 & n2923;
  assign n2925 = ~n338 & ~n648;
  assign n2926 = ~n288 & ~n313;
  assign n2927 = ~n343 & ~n382;
  assign n2928 = ~n591 & ~n645;
  assign n2929 = ~n674 & n2928;
  assign n2930 = n2926 & n2927;
  assign n2931 = n969 & n2754;
  assign n2932 = n2925 & n2931;
  assign n2933 = n2929 & n2930;
  assign n2934 = n1265 & n1629;
  assign n2935 = n2522 & n2908;
  assign n2936 = n2924 & n2935;
  assign n2937 = n2933 & n2934;
  assign n2938 = n2932 & n2937;
  assign n2939 = n2914 & n2936;
  assign n2940 = n2938 & n2939;
  assign n2941 = n2922 & n2940;
  assign n2942 = ~n364 & ~n700;
  assign n2943 = ~n208 & ~n296;
  assign n2944 = ~n207 & ~n363;
  assign n2945 = ~n219 & ~n689;
  assign n2946 = ~n588 & n1237;
  assign n2947 = n2300 & n2942;
  assign n2948 = n2943 & n2944;
  assign n2949 = n2945 & n2948;
  assign n2950 = n2946 & n2947;
  assign n2951 = n2869 & n2950;
  assign n2952 = n2949 & n2951;
  assign n2953 = ~n324 & ~n574;
  assign n2954 = ~n283 & n1536;
  assign n2955 = n2566 & n2953;
  assign n2956 = n2954 & n2955;
  assign n2957 = ~n285 & ~n583;
  assign n2958 = ~n339 & ~n554;
  assign n2959 = ~n109 & ~n424;
  assign n2960 = ~n250 & ~n545;
  assign n2961 = ~n590 & n2960;
  assign n2962 = n854 & n2957;
  assign n2963 = n2958 & n2959;
  assign n2964 = n2962 & n2963;
  assign n2965 = n2961 & n2964;
  assign n2966 = ~n580 & ~n595;
  assign n2967 = ~n599 & n2966;
  assign n2968 = n1242 & n1339;
  assign n2969 = n1432 & n2968;
  assign n2970 = n2905 & n2967;
  assign n2971 = n2969 & n2970;
  assign n2972 = n2091 & n2956;
  assign n2973 = n2971 & n2972;
  assign n2974 = n478 & n2965;
  assign n2975 = n2973 & n2974;
  assign n2976 = n2952 & n2975;
  assign n2977 = n458 & n2976;
  assign n2978 = n2941 & n2977;
  assign n2979 = ~n2901 & ~n2978;
  assign n2980 = ~n251 & n524;
  assign n2981 = ~n234 & ~n406;
  assign n2982 = ~n149 & ~n222;
  assign n2983 = ~n253 & ~n318;
  assign n2984 = ~n513 & ~n673;
  assign n2985 = n2983 & n2984;
  assign n2986 = n114 & n2982;
  assign n2987 = n939 & n1392;
  assign n2988 = n2419 & n2981;
  assign n2989 = n2987 & n2988;
  assign n2990 = n2985 & n2986;
  assign n2991 = n2980 & n2990;
  assign n2992 = n2989 & n2991;
  assign n2993 = ~n254 & ~n404;
  assign n2994 = ~n546 & n2993;
  assign n2995 = ~n136 & ~n216;
  assign n2996 = ~n339 & ~n466;
  assign n2997 = ~n543 & ~n590;
  assign n2998 = n2996 & n2997;
  assign n2999 = n904 & n2995;
  assign n3000 = n2998 & n2999;
  assign n3001 = n2994 & n3000;
  assign n3002 = ~n343 & ~n666;
  assign n3003 = ~n676 & n3002;
  assign n3004 = n169 & n328;
  assign n3005 = n3003 & n3004;
  assign n3006 = ~n164 & ~n250;
  assign n3007 = ~n307 & n3006;
  assign n3008 = n804 & n3007;
  assign n3009 = ~n662 & n2296;
  assign n3010 = n1968 & n3009;
  assign n3011 = ~n120 & ~n172;
  assign n3012 = ~n215 & ~n244;
  assign n3013 = ~n407 & n3012;
  assign n3014 = n1054 & n3011;
  assign n3015 = n1125 & n1237;
  assign n3016 = n1807 & n3015;
  assign n3017 = n3013 & n3014;
  assign n3018 = n1617 & n2884;
  assign n3019 = n3017 & n3018;
  assign n3020 = n2270 & n3016;
  assign n3021 = n3005 & n3008;
  assign n3022 = n3010 & n3021;
  assign n3023 = n3019 & n3020;
  assign n3024 = n3022 & n3023;
  assign n3025 = ~n180 & ~n213;
  assign n3026 = ~n521 & n3025;
  assign n3027 = ~n98 & ~n270;
  assign n3028 = ~n494 & n3027;
  assign n3029 = ~n125 & ~n179;
  assign n3030 = ~n289 & ~n571;
  assign n3031 = ~n646 & n3030;
  assign n3032 = n1117 & n3029;
  assign n3033 = n3031 & n3032;
  assign n3034 = ~n246 & ~n363;
  assign n3035 = ~n313 & ~n469;
  assign n3036 = ~n554 & ~n594;
  assign n3037 = ~n683 & n3036;
  assign n3038 = n2451 & n3035;
  assign n3039 = n3034 & n3038;
  assign n3040 = n3037 & n3039;
  assign n3041 = ~n182 & ~n334;
  assign n3042 = ~n360 & ~n598;
  assign n3043 = n3041 & n3042;
  assign n3044 = n854 & n1391;
  assign n3045 = n1534 & n1764;
  assign n3046 = n3044 & n3045;
  assign n3047 = n3026 & n3043;
  assign n3048 = n3028 & n3047;
  assign n3049 = n3033 & n3046;
  assign n3050 = n3048 & n3049;
  assign n3051 = n3040 & n3050;
  assign n3052 = ~n445 & ~n568;
  assign n3053 = ~n85 & ~n219;
  assign n3054 = ~n242 & ~n459;
  assign n3055 = ~n467 & ~n570;
  assign n3056 = n3054 & n3055;
  assign n3057 = n842 & n3053;
  assign n3058 = n882 & n1650;
  assign n3059 = n1817 & n2097;
  assign n3060 = n2475 & n3052;
  assign n3061 = n3059 & n3060;
  assign n3062 = n3057 & n3058;
  assign n3063 = n1359 & n3056;
  assign n3064 = n3062 & n3063;
  assign n3065 = n3061 & n3064;
  assign n3066 = n3001 & n3065;
  assign n3067 = n2992 & n3066;
  assign n3068 = n3024 & n3051;
  assign n3069 = n3067 & n3068;
  assign n3070 = ~n2978 & ~n3069;
  assign n3071 = ~n175 & ~n239;
  assign n3072 = ~n402 & ~n591;
  assign n3073 = ~n389 & ~n646;
  assign n3074 = ~n543 & n3073;
  assign n3075 = ~n179 & ~n510;
  assign n3076 = n3074 & n3075;
  assign n3077 = ~n212 & n1041;
  assign n3078 = ~n320 & ~n359;
  assign n3079 = ~n483 & ~n546;
  assign n3080 = ~n164 & ~n673;
  assign n3081 = ~n163 & ~n222;
  assign n3082 = ~n267 & ~n425;
  assign n3083 = n3081 & n3082;
  assign n3084 = n3080 & n3083;
  assign n3085 = ~n339 & ~n472;
  assign n3086 = ~n236 & ~n311;
  assign n3087 = ~n234 & ~n420;
  assign n3088 = n3086 & n3087;
  assign n3089 = n1287 & n2049;
  assign n3090 = n3085 & n3089;
  assign n3091 = n3088 & n3090;
  assign n3092 = ~n238 & ~n376;
  assign n3093 = ~n405 & ~n582;
  assign n3094 = ~n651 & n3093;
  assign n3095 = n2092 & n3092;
  assign n3096 = n3078 & n3079;
  assign n3097 = n3095 & n3096;
  assign n3098 = n903 & n3094;
  assign n3099 = n1968 & n3077;
  assign n3100 = n3098 & n3099;
  assign n3101 = n3084 & n3097;
  assign n3102 = n3100 & n3101;
  assign n3103 = n3091 & n3102;
  assign n3104 = n2295 & n3103;
  assign n3105 = ~n193 & ~n307;
  assign n3106 = ~n120 & ~n145;
  assign n3107 = ~n182 & ~n269;
  assign n3108 = ~n343 & ~n362;
  assign n3109 = ~n659 & ~n690;
  assign n3110 = n3108 & n3109;
  assign n3111 = n3106 & n3107;
  assign n3112 = n497 & n740;
  assign n3113 = n1942 & n2234;
  assign n3114 = n2634 & n3105;
  assign n3115 = n3113 & n3114;
  assign n3116 = n3111 & n3112;
  assign n3117 = n3110 & n3116;
  assign n3118 = n1378 & n3115;
  assign n3119 = n3117 & n3118;
  assign n3120 = ~n103 & ~n219;
  assign n3121 = ~n276 & ~n290;
  assign n3122 = ~n374 & ~n463;
  assign n3123 = n3121 & n3122;
  assign n3124 = n217 & n3120;
  assign n3125 = n493 & n1085;
  assign n3126 = n1508 & n2475;
  assign n3127 = n3071 & n3072;
  assign n3128 = n3126 & n3127;
  assign n3129 = n3124 & n3125;
  assign n3130 = n1316 & n3123;
  assign n3131 = n3129 & n3130;
  assign n3132 = n3076 & n3128;
  assign n3133 = n3131 & n3132;
  assign n3134 = n2839 & n3133;
  assign n3135 = n3119 & n3134;
  assign n3136 = n2753 & n3135;
  assign n3137 = n3104 & n3136;
  assign n3138 = ~n3069 & ~n3137;
  assign n3139 = n1538 & n1764;
  assign n3140 = ~n126 & ~n215;
  assign n3141 = ~n247 & ~n287;
  assign n3142 = n3140 & n3141;
  assign n3143 = ~n177 & ~n364;
  assign n3144 = ~n391 & ~n701;
  assign n3145 = n3143 & n3144;
  assign n3146 = n623 & n930;
  assign n3147 = n1339 & n1760;
  assign n3148 = n2686 & n2706;
  assign n3149 = n3147 & n3148;
  assign n3150 = n3145 & n3146;
  assign n3151 = n3139 & n3142;
  assign n3152 = n3150 & n3151;
  assign n3153 = n3149 & n3152;
  assign n3154 = ~n175 & ~n316;
  assign n3155 = ~n165 & ~n496;
  assign n3156 = ~n144 & ~n235;
  assign n3157 = ~n310 & ~n338;
  assign n3158 = ~n343 & ~n448;
  assign n3159 = n3157 & n3158;
  assign n3160 = n114 & n3156;
  assign n3161 = n555 & n1247;
  assign n3162 = n1279 & n3154;
  assign n3163 = n3155 & n3162;
  assign n3164 = n3160 & n3161;
  assign n3165 = n718 & n3159;
  assign n3166 = n3164 & n3165;
  assign n3167 = n3163 & n3166;
  assign n3168 = n1767 & n3167;
  assign n3169 = ~n167 & ~n315;
  assign n3170 = ~n221 & ~n406;
  assign n3171 = ~n513 & ~n521;
  assign n3172 = ~n179 & ~n326;
  assign n3173 = ~n203 & ~n318;
  assign n3174 = ~n427 & n3173;
  assign n3175 = n197 & n3172;
  assign n3176 = n3174 & n3175;
  assign n3177 = ~n591 & n967;
  assign n3178 = n1395 & n3177;
  assign n3179 = ~n131 & ~n324;
  assign n3180 = ~n462 & ~n538;
  assign n3181 = ~n543 & n3180;
  assign n3182 = n471 & n3179;
  assign n3183 = n2909 & n3169;
  assign n3184 = n3170 & n3171;
  assign n3185 = n3183 & n3184;
  assign n3186 = n3181 & n3182;
  assign n3187 = n3185 & n3186;
  assign n3188 = n815 & n3176;
  assign n3189 = n3178 & n3188;
  assign n3190 = n1390 & n3187;
  assign n3191 = n3189 & n3190;
  assign n3192 = n3153 & n3191;
  assign n3193 = n3103 & n3168;
  assign n3194 = n3192 & n3193;
  assign n3195 = ~n3137 & ~n3194;
  assign n3196 = ~n288 & ~n384;
  assign n3197 = n255 & n3196;
  assign n3198 = ~n109 & ~n180;
  assign n3199 = ~n447 & n3198;
  assign n3200 = n586 & n912;
  assign n3201 = n3199 & n3200;
  assign n3202 = n3197 & n3201;
  assign n3203 = ~n405 & ~n511;
  assign n3204 = ~n318 & ~n649;
  assign n3205 = ~n244 & ~n580;
  assign n3206 = ~n118 & ~n148;
  assign n3207 = ~n570 & n3206;
  assign n3208 = n211 & n220;
  assign n3209 = n3203 & n3204;
  assign n3210 = n3205 & n3209;
  assign n3211 = n3207 & n3208;
  assign n3212 = n3077 & n3211;
  assign n3213 = n3210 & n3212;
  assign n3214 = ~n271 & ~n300;
  assign n3215 = ~n545 & ~n644;
  assign n3216 = n3214 & n3215;
  assign n3217 = n278 & n848;
  assign n3218 = n1537 & n1837;
  assign n3219 = n2226 & n2323;
  assign n3220 = n2634 & n3219;
  assign n3221 = n3217 & n3218;
  assign n3222 = n3216 & n3221;
  assign n3223 = n3220 & n3222;
  assign n3224 = n3202 & n3223;
  assign n3225 = n3213 & n3224;
  assign n3226 = n1646 & n2023;
  assign n3227 = n3225 & n3226;
  assign n3228 = ~n3194 & ~n3227;
  assign n3229 = ~n180 & ~n192;
  assign n3230 = ~n365 & n3229;
  assign n3231 = ~n203 & ~n466;
  assign n3232 = n3230 & n3231;
  assign n3233 = ~n235 & ~n578;
  assign n3234 = ~n147 & ~n243;
  assign n3235 = ~n644 & n3234;
  assign n3236 = n741 & n1614;
  assign n3237 = n1756 & n2450;
  assign n3238 = n2565 & n3171;
  assign n3239 = n3233 & n3238;
  assign n3240 = n3236 & n3237;
  assign n3241 = n2397 & n3235;
  assign n3242 = n3240 & n3241;
  assign n3243 = n3232 & n3239;
  assign n3244 = n3242 & n3243;
  assign n3245 = n2188 & n3244;
  assign n3246 = ~n424 & ~n661;
  assign n3247 = ~n687 & n3246;
  assign n3248 = ~n125 & ~n405;
  assign n3249 = ~n376 & ~n690;
  assign n3250 = n1583 & n3249;
  assign n3251 = ~n389 & n3052;
  assign n3252 = n3248 & n3251;
  assign n3253 = n3247 & n3252;
  assign n3254 = n3250 & n3253;
  assign n3255 = ~n216 & ~n360;
  assign n3256 = n2322 & n3255;
  assign n3257 = ~n250 & ~n671;
  assign n3258 = ~n686 & n3257;
  assign n3259 = n1170 & n2293;
  assign n3260 = n2755 & n3259;
  assign n3261 = n3258 & n3260;
  assign n3262 = ~n323 & n967;
  assign n3263 = n1203 & n3262;
  assign n3264 = ~n144 & ~n265;
  assign n3265 = ~n307 & n3264;
  assign n3266 = ~n276 & ~n473;
  assign n3267 = ~n269 & ~n297;
  assign n3268 = ~n541 & n2659;
  assign n3269 = ~n465 & n928;
  assign n3270 = n1281 & n3269;
  assign n3271 = ~n312 & ~n374;
  assign n3272 = ~n287 & ~n387;
  assign n3273 = ~n447 & ~n681;
  assign n3274 = n3272 & n3273;
  assign n3275 = n842 & n1868;
  assign n3276 = n2981 & n3271;
  assign n3277 = n3275 & n3276;
  assign n3278 = n3268 & n3274;
  assign n3279 = n3277 & n3278;
  assign n3280 = n3270 & n3279;
  assign n3281 = ~n251 & ~n666;
  assign n3282 = ~n113 & ~n649;
  assign n3283 = ~n91 & ~n182;
  assign n3284 = ~n320 & ~n544;
  assign n3285 = n3283 & n3284;
  assign n3286 = n1267 & n3281;
  assign n3287 = n3282 & n3286;
  assign n3288 = n3285 & n3287;
  assign n3289 = ~n492 & ~n495;
  assign n3290 = ~n641 & ~n679;
  assign n3291 = n3289 & n3290;
  assign n3292 = n137 & n403;
  assign n3293 = n1085 & n1587;
  assign n3294 = n2358 & n3266;
  assign n3295 = n3267 & n3294;
  assign n3296 = n3292 & n3293;
  assign n3297 = n2547 & n3291;
  assign n3298 = n3265 & n3297;
  assign n3299 = n3295 & n3296;
  assign n3300 = n3298 & n3299;
  assign n3301 = n3288 & n3300;
  assign n3302 = n3280 & n3301;
  assign n3303 = ~n148 & ~n168;
  assign n3304 = ~n404 & ~n570;
  assign n3305 = ~n571 & ~n640;
  assign n3306 = ~n648 & n3305;
  assign n3307 = n3303 & n3304;
  assign n3308 = n461 & n471;
  assign n3309 = n600 & n622;
  assign n3310 = n2299 & n3309;
  assign n3311 = n3307 & n3308;
  assign n3312 = n3256 & n3306;
  assign n3313 = n3311 & n3312;
  assign n3314 = n3263 & n3310;
  assign n3315 = n3313 & n3314;
  assign n3316 = n3261 & n3315;
  assign n3317 = n3254 & n3316;
  assign n3318 = n3245 & n3317;
  assign n3319 = n3302 & n3318;
  assign n3320 = ~n3227 & ~n3319;
  assign n3321 = n3227 & n3319;
  assign n3322 = ~n3320 & ~n3321;
  assign n3323 = ~n244 & ~n572;
  assign n3324 = ~n681 & n3323;
  assign n3325 = ~n215 & ~n222;
  assign n3326 = ~n379 & n3325;
  assign n3327 = n481 & n3326;
  assign n3328 = n1896 & n3327;
  assign n3329 = ~n265 & ~n338;
  assign n3330 = ~n460 & n3329;
  assign n3331 = n284 & n403;
  assign n3332 = n600 & n740;
  assign n3333 = n927 & n1302;
  assign n3334 = n3332 & n3333;
  assign n3335 = n3330 & n3331;
  assign n3336 = n2233 & n3324;
  assign n3337 = n3335 & n3336;
  assign n3338 = n3334 & n3337;
  assign n3339 = n3040 & n3328;
  assign n3340 = n3338 & n3339;
  assign n3341 = ~n131 & ~n446;
  assign n3342 = ~n580 & n3341;
  assign n3343 = ~n390 & ~n422;
  assign n3344 = ~n473 & ~n595;
  assign n3345 = n3343 & n3344;
  assign n3346 = ~n193 & ~n199;
  assign n3347 = ~n218 & ~n240;
  assign n3348 = ~n354 & n3347;
  assign n3349 = n2599 & n3348;
  assign n3350 = ~n122 & ~n467;
  assign n3351 = ~n136 & ~n494;
  assign n3352 = ~n167 & ~n251;
  assign n3353 = ~n92 & ~n120;
  assign n3354 = ~n225 & ~n269;
  assign n3355 = ~n336 & ~n577;
  assign n3356 = n3354 & n3355;
  assign n3357 = n2419 & n3353;
  assign n3358 = n3170 & n3350;
  assign n3359 = n3351 & n3352;
  assign n3360 = n3358 & n3359;
  assign n3361 = n3356 & n3357;
  assign n3362 = n3360 & n3361;
  assign n3363 = ~n118 & ~n391;
  assign n3364 = n781 & n3363;
  assign n3365 = n882 & n1241;
  assign n3366 = n2008 & n3346;
  assign n3367 = n3365 & n3366;
  assign n3368 = n3342 & n3364;
  assign n3369 = n3345 & n3368;
  assign n3370 = n295 & n3367;
  assign n3371 = n3010 & n3349;
  assign n3372 = n3370 & n3371;
  assign n3373 = n3362 & n3369;
  assign n3374 = n3372 & n3373;
  assign n3375 = n3245 & n3374;
  assign n3376 = n3340 & n3375;
  assign n3377 = ~n183 & ~n469;
  assign n3378 = n268 & n3377;
  assign n3379 = ~n467 & ~n661;
  assign n3380 = ~n311 & ~n462;
  assign n3381 = ~n133 & ~n459;
  assign n3382 = ~n144 & ~n640;
  assign n3383 = n1807 & n3382;
  assign n3384 = n2194 & n2358;
  assign n3385 = n2728 & n2783;
  assign n3386 = n3384 & n3385;
  assign n3387 = n1348 & n3383;
  assign n3388 = n3386 & n3387;
  assign n3389 = ~n136 & ~n595;
  assign n3390 = n1631 & n3389;
  assign n3391 = ~n180 & ~n242;
  assign n3392 = ~n286 & ~n320;
  assign n3393 = ~n538 & ~n585;
  assign n3394 = n3392 & n3393;
  assign n3395 = n281 & n3391;
  assign n3396 = n732 & n1970;
  assign n3397 = n3395 & n3396;
  assign n3398 = n3390 & n3394;
  assign n3399 = n3397 & n3398;
  assign n3400 = ~n336 & n731;
  assign n3401 = ~n584 & ~n665;
  assign n3402 = ~n269 & n2066;
  assign n3403 = n3401 & n3402;
  assign n3404 = ~n356 & ~n544;
  assign n3405 = ~n427 & ~n671;
  assign n3406 = n383 & n3405;
  assign n3407 = n408 & n1203;
  assign n3408 = n1431 & n1457;
  assign n3409 = n2087 & n2096;
  assign n3410 = n3204 & n3404;
  assign n3411 = n3409 & n3410;
  assign n3412 = n3407 & n3408;
  assign n3413 = n3400 & n3406;
  assign n3414 = n3412 & n3413;
  assign n3415 = n3076 & n3411;
  assign n3416 = n3403 & n3415;
  assign n3417 = n3399 & n3414;
  assign n3418 = n3416 & n3417;
  assign n3419 = ~n463 & ~n465;
  assign n3420 = ~n335 & ~n420;
  assign n3421 = ~n680 & n3420;
  assign n3422 = n3419 & n3421;
  assign n3423 = n1506 & n3422;
  assign n3424 = ~n514 & ~n541;
  assign n3425 = n1121 & n3424;
  assign n3426 = ~n246 & ~n424;
  assign n3427 = ~n236 & ~n319;
  assign n3428 = ~n148 & ~n316;
  assign n3429 = ~n92 & ~n196;
  assign n3430 = ~n662 & n3429;
  assign n3431 = n3427 & n3428;
  assign n3432 = n3430 & n3431;
  assign n3433 = n765 & n1233;
  assign n3434 = n1455 & n1534;
  assign n3435 = n2150 & n2754;
  assign n3436 = n3426 & n3435;
  assign n3437 = n3433 & n3434;
  assign n3438 = n1053 & n3425;
  assign n3439 = n3437 & n3438;
  assign n3440 = n3432 & n3436;
  assign n3441 = n3439 & n3440;
  assign n3442 = n3423 & n3441;
  assign n3443 = ~n213 & ~n327;
  assign n3444 = ~n378 & ~n582;
  assign n3445 = n3443 & n3444;
  assign n3446 = n361 & n449;
  assign n3447 = n624 & n920;
  assign n3448 = n1651 & n2472;
  assign n3449 = n2565 & n2903;
  assign n3450 = n3379 & n3380;
  assign n3451 = n3381 & n3450;
  assign n3452 = n3448 & n3449;
  assign n3453 = n3446 & n3447;
  assign n3454 = n3378 & n3445;
  assign n3455 = n3453 & n3454;
  assign n3456 = n3451 & n3452;
  assign n3457 = n3455 & n3456;
  assign n3458 = n3388 & n3457;
  assign n3459 = n3418 & n3458;
  assign n3460 = n3442 & n3459;
  assign n3461 = n3319 & n3460;
  assign n3462 = ~n3376 & ~n3461;
  assign n3463 = n3322 & n3462;
  assign n3464 = ~n3320 & ~n3463;
  assign n3465 = n3194 & n3227;
  assign n3466 = ~n3228 & ~n3465;
  assign n3467 = ~n3464 & n3466;
  assign n3468 = ~n3228 & ~n3467;
  assign n3469 = n3137 & n3194;
  assign n3470 = ~n3195 & ~n3469;
  assign n3471 = ~n3468 & n3470;
  assign n3472 = ~n3195 & ~n3471;
  assign n3473 = n3069 & n3137;
  assign n3474 = ~n3138 & ~n3473;
  assign n3475 = ~n3472 & n3474;
  assign n3476 = ~n3138 & ~n3475;
  assign n3477 = n2978 & n3069;
  assign n3478 = ~n3070 & ~n3477;
  assign n3479 = ~n3476 & n3478;
  assign n3480 = ~n3070 & ~n3479;
  assign n3481 = n2901 & n2978;
  assign n3482 = ~n2979 & ~n3481;
  assign n3483 = ~n3480 & n3482;
  assign n3484 = ~n2979 & ~n3483;
  assign n3485 = n2866 & n2901;
  assign n3486 = ~n2902 & ~n3485;
  assign n3487 = ~n3484 & n3486;
  assign n3488 = ~n2902 & ~n3487;
  assign n3489 = n2781 & n2866;
  assign n3490 = ~n2867 & ~n3489;
  assign n3491 = ~n3488 & n3490;
  assign n3492 = ~n2867 & ~n3491;
  assign n3493 = n2726 & n2781;
  assign n3494 = ~n2782 & ~n3493;
  assign n3495 = ~n3492 & n3494;
  assign n3496 = ~n2782 & ~n3495;
  assign n3497 = n2657 & n2726;
  assign n3498 = ~n2727 & ~n3497;
  assign n3499 = ~n3496 & n3498;
  assign n3500 = ~n2727 & ~n3499;
  assign n3501 = n2622 & n2657;
  assign n3502 = ~n2658 & ~n3501;
  assign n3503 = ~n3500 & n3502;
  assign n3504 = ~n2658 & ~n3503;
  assign n3505 = n2538 & n2622;
  assign n3506 = ~n2623 & ~n3505;
  assign n3507 = ~n3504 & n3506;
  assign n3508 = ~n2623 & ~n3507;
  assign n3509 = n2442 & n2538;
  assign n3510 = ~n2539 & ~n3509;
  assign n3511 = ~n3508 & n3510;
  assign n3512 = ~n2539 & ~n3511;
  assign n3513 = n2356 & n2442;
  assign n3514 = ~n2443 & ~n3513;
  assign n3515 = ~n3512 & n3514;
  assign n3516 = ~n2443 & ~n3515;
  assign n3517 = n2265 & n2356;
  assign n3518 = ~n2357 & ~n3517;
  assign n3519 = ~n3516 & n3518;
  assign n3520 = ~n2357 & ~n3519;
  assign n3521 = n2165 & n2265;
  assign n3522 = ~n2266 & ~n3521;
  assign n3523 = ~n3520 & n3522;
  assign n3524 = ~n2266 & ~n3523;
  assign n3525 = n2045 & n2165;
  assign n3526 = ~n2166 & ~n3525;
  assign n3527 = ~n3524 & n3526;
  assign n3528 = ~n2166 & ~n3527;
  assign n3529 = n1997 & n2045;
  assign n3530 = ~n2046 & ~n3529;
  assign n3531 = ~n3528 & n3530;
  assign n3532 = ~n2046 & ~n3531;
  assign n3533 = n1893 & n1997;
  assign n3534 = ~n1998 & ~n3533;
  assign n3535 = ~n3532 & n3534;
  assign n3536 = ~n1998 & ~n3535;
  assign n3537 = n1805 & n1893;
  assign n3538 = ~n1894 & ~n3537;
  assign n3539 = ~n3536 & n3538;
  assign n3540 = ~n1894 & ~n3539;
  assign n3541 = n1737 & n1805;
  assign n3542 = ~n1806 & ~n3541;
  assign n3543 = ~n3540 & n3542;
  assign n3544 = ~n1806 & ~n3543;
  assign n3545 = n1610 & n1737;
  assign n3546 = ~n1738 & ~n3545;
  assign n3547 = ~n3544 & n3546;
  assign n3548 = ~n1738 & ~n3547;
  assign n3549 = n1532 & n1610;
  assign n3550 = ~n1611 & ~n3549;
  assign n3551 = ~n3548 & n3550;
  assign n3552 = ~n1611 & ~n3551;
  assign n3553 = n1425 & n1532;
  assign n3554 = ~n1533 & ~n3553;
  assign n3555 = ~n3552 & n3554;
  assign n3556 = ~n1533 & ~n3555;
  assign n3557 = n1337 & n1425;
  assign n3558 = ~n1426 & ~n3557;
  assign n3559 = ~n3556 & n3558;
  assign n3560 = ~n1426 & ~n3559;
  assign n3561 = n1230 & n1337;
  assign n3562 = ~n1338 & ~n3561;
  assign n3563 = ~n3560 & n3562;
  assign n3564 = ~n1338 & ~n3563;
  assign n3565 = n1107 & n1230;
  assign n3566 = ~n1231 & ~n3565;
  assign n3567 = ~n3564 & n3566;
  assign n3568 = ~n1231 & ~n3567;
  assign n3569 = n1006 & n1107;
  assign n3570 = ~n1108 & ~n3569;
  assign n3571 = ~n3568 & n3570;
  assign n3572 = ~n1108 & ~n3571;
  assign n3573 = n898 & n1006;
  assign n3574 = ~n1007 & ~n3573;
  assign n3575 = ~n3572 & n3574;
  assign n3576 = ~n1007 & ~n3575;
  assign n3577 = n802 & n898;
  assign n3578 = ~n899 & ~n3577;
  assign n3579 = ~n3576 & n3578;
  assign n3580 = ~n899 & ~n3579;
  assign n3581 = n729 & n802;
  assign n3582 = ~n803 & ~n3581;
  assign n3583 = ~n3580 & n3582;
  assign n3584 = ~n803 & ~n3583;
  assign n3585 = n621 & n729;
  assign n3586 = ~n730 & ~n3585;
  assign n3587 = ~n3584 & n3586;
  assign n3588 = ~n730 & ~n3587;
  assign n3589 = ~n563 & ~n621;
  assign n3590 = n535 & n621;
  assign n3591 = ~n3589 & ~n3590;
  assign n3592 = ~n3588 & n3591;
  assign n3593 = n621 & ~n3592;
  assign n3594 = n566 & ~n3593;
  assign n3595 = ~n564 & ~n3594;
  assign n3596 = ~n563 & ~n3595;
  assign n3597 = n508 & n3596;
  assign n3598 = ~n506 & ~n3597;
  assign n3599 = n129 & n205;
  assign n3600 = ~n139 & ~n382;
  assign n3601 = ~n568 & n3600;
  assign n3602 = n439 & n3601;
  assign n3603 = n3599 & n3602;
  assign n3604 = n614 & n3603;
  assign n3605 = n716 & n3604;
  assign n3606 = n419 & n3605;
  assign n3607 = ~n419 & ~n3605;
  assign n3608 = ~n3606 & ~n3607;
  assign n3609 = ~n3598 & ~n3608;
  assign n3610 = ~n216 & ~n236;
  assign n3611 = n377 & n3610;
  assign n3612 = ~n177 & ~n315;
  assign n3613 = ~n512 & ~n597;
  assign n3614 = n3612 & n3613;
  assign n3615 = n732 & n849;
  assign n3616 = n1541 & n2227;
  assign n3617 = n2305 & n3616;
  assign n3618 = n3614 & n3615;
  assign n3619 = n438 & n3618;
  assign n3620 = n3617 & n3619;
  assign n3621 = ~n421 & ~n448;
  assign n3622 = ~n521 & n3621;
  assign n3623 = n3620 & n3622;
  assign n3624 = ~n313 & ~n378;
  assign n3625 = ~n240 & ~n310;
  assign n3626 = ~n650 & n3625;
  assign n3627 = ~n222 & ~n336;
  assign n3628 = ~n338 & ~n513;
  assign n3629 = ~n173 & ~n340;
  assign n3630 = ~n462 & ~n479;
  assign n3631 = n3629 & n3630;
  assign n3632 = n325 & n2170;
  assign n3633 = n3627 & n3628;
  assign n3634 = n3632 & n3633;
  assign n3635 = n3626 & n3631;
  assign n3636 = n3634 & n3635;
  assign n3637 = ~n144 & ~n196;
  assign n3638 = ~n335 & ~n582;
  assign n3639 = ~n659 & ~n666;
  assign n3640 = n3638 & n3639;
  assign n3641 = n201 & n3637;
  assign n3642 = n1247 & n2097;
  assign n3643 = n2220 & n3204;
  assign n3644 = n3624 & n3643;
  assign n3645 = n3641 & n3642;
  assign n3646 = n1906 & n3640;
  assign n3647 = n3230 & n3611;
  assign n3648 = n3646 & n3647;
  assign n3649 = n3644 & n3645;
  assign n3650 = n2458 & n3649;
  assign n3651 = n1688 & n3648;
  assign n3652 = n3636 & n3651;
  assign n3653 = n3650 & n3652;
  assign n3654 = n2023 & n3623;
  assign n3655 = n3653 & n3654;
  assign n3656 = ~n382 & ~n462;
  assign n3657 = ~n208 & n1760;
  assign n3658 = ~n447 & ~n545;
  assign n3659 = n3657 & n3658;
  assign n3660 = n780 & n3659;
  assign n3661 = ~n144 & n523;
  assign n3662 = n2093 & n2192;
  assign n3663 = n2452 & n3656;
  assign n3664 = n3662 & n3663;
  assign n3665 = n3661 & n3664;
  assign n3666 = n443 & n3665;
  assign n3667 = n264 & n3666;
  assign n3668 = n306 & n698;
  assign n3669 = n3667 & n3668;
  assign n3670 = n3660 & n3669;
  assign n3671 = ~n3655 & ~n3670;
  assign n3672 = n3655 & n3670;
  assign n3673 = ~n3671 & ~n3672;
  assign n3674 = ~pi29  & n3673;
  assign n3675 = ~n3671 & ~n3674;
  assign n3676 = n419 & ~n3675;
  assign n3677 = ~n419 & n3675;
  assign n3678 = ~n3676 & ~n3677;
  assign n3679 = n564 & ~n621;
  assign n3680 = pi30  & ~pi31 ;
  assign n3681 = ~pi30  & pi31 ;
  assign n3682 = ~n3680 & ~n3681;
  assign n3683 = n565 & ~n3682;
  assign n3684 = ~n563 & n3683;
  assign n3685 = n563 & ~n3592;
  assign n3686 = ~n563 & ~n3593;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = n566 & n3687;
  assign n3689 = ~n3679 & ~n3684;
  assign n3690 = ~n3688 & n3689;
  assign n3691 = n3678 & ~n3690;
  assign n3692 = ~n3676 & ~n3691;
  assign n3693 = ~n508 & ~n3596;
  assign n3694 = ~n3597 & ~n3693;
  assign n3695 = ~n3692 & n3694;
  assign n3696 = n3692 & ~n3694;
  assign n3697 = ~n3695 & ~n3696;
  assign n3698 = ~n134 & ~n175;
  assign n3699 = ~n212 & n3698;
  assign n3700 = ~n193 & ~n702;
  assign n3701 = ~n254 & ~n335;
  assign n3702 = ~n362 & ~n568;
  assign n3703 = ~n591 & n3702;
  assign n3704 = n1208 & n3701;
  assign n3705 = n1538 & n1632;
  assign n3706 = n1956 & n3700;
  assign n3707 = n3705 & n3706;
  assign n3708 = n3703 & n3704;
  assign n3709 = n3707 & n3708;
  assign n3710 = ~n420 & ~n469;
  assign n3711 = ~n139 & n3710;
  assign n3712 = ~n277 & ~n374;
  assign n3713 = ~n543 & n3712;
  assign n3714 = ~n136 & ~n182;
  assign n3715 = ~n651 & n3714;
  assign n3716 = ~n270 & ~n389;
  assign n3717 = ~n645 & ~n673;
  assign n3718 = ~n682 & n3717;
  assign n3719 = n1394 & n3716;
  assign n3720 = n1630 & n3628;
  assign n3721 = n3719 & n3720;
  assign n3722 = n1761 & n3718;
  assign n3723 = n3713 & n3715;
  assign n3724 = n3722 & n3723;
  assign n3725 = n2821 & n3721;
  assign n3726 = n3005 & n3725;
  assign n3727 = n3724 & n3726;
  assign n3728 = n2952 & n3727;
  assign n3729 = ~n271 & ~n319;
  assign n3730 = ~n245 & ~n482;
  assign n3731 = ~n536 & n3730;
  assign n3732 = ~n109 & ~n162;
  assign n3733 = ~n426 & ~n465;
  assign n3734 = ~n511 & ~n594;
  assign n3735 = n3733 & n3734;
  assign n3736 = n166 & n3732;
  assign n3737 = n252 & n643;
  assign n3738 = n1246 & n1869;
  assign n3739 = n3729 & n3738;
  assign n3740 = n3736 & n3737;
  assign n3741 = n1961 & n3735;
  assign n3742 = n3731 & n3741;
  assign n3743 = n3739 & n3740;
  assign n3744 = n3742 & n3743;
  assign n3745 = ~n242 & ~n354;
  assign n3746 = ~n385 & ~n473;
  assign n3747 = ~n514 & ~n544;
  assign n3748 = ~n601 & n3747;
  assign n3749 = n3745 & n3746;
  assign n3750 = n464 & n581;
  assign n3751 = n586 & n1457;
  assign n3752 = n3750 & n3751;
  assign n3753 = n3748 & n3749;
  assign n3754 = n817 & n3699;
  assign n3755 = n3711 & n3754;
  assign n3756 = n3752 & n3753;
  assign n3757 = n3755 & n3756;
  assign n3758 = n1321 & n3709;
  assign n3759 = n3757 & n3758;
  assign n3760 = n3744 & n3759;
  assign n3761 = n3728 & n3760;
  assign n3762 = n3655 & ~n3761;
  assign n3763 = ~n335 & ~n670;
  assign n3764 = ~n179 & ~n225;
  assign n3765 = ~n296 & ~n359;
  assign n3766 = ~n661 & ~n686;
  assign n3767 = n3765 & n3766;
  assign n3768 = n1042 & n3764;
  assign n3769 = n3767 & n3768;
  assign n3770 = ~n360 & ~n362;
  assign n3771 = ~n427 & ~n554;
  assign n3772 = n3770 & n3771;
  assign n3773 = n1152 & n1485;
  assign n3774 = n2360 & n2523;
  assign n3775 = n3426 & n3774;
  assign n3776 = n3772 & n3773;
  assign n3777 = n3775 & n3776;
  assign n3778 = ~n250 & ~n645;
  assign n3779 = ~n363 & ~n690;
  assign n3780 = n3778 & n3779;
  assign n3781 = n3699 & n3780;
  assign n3782 = ~n480 & ~n513;
  assign n3783 = ~n641 & n3782;
  assign n3784 = ~n277 & ~n568;
  assign n3785 = ~n590 & n3784;
  assign n3786 = ~n109 & ~n244;
  assign n3787 = ~n342 & ~n405;
  assign n3788 = ~n446 & ~n448;
  assign n3789 = ~n679 & n3788;
  assign n3790 = n3786 & n3787;
  assign n3791 = n3789 & n3790;
  assign n3792 = n3783 & n3785;
  assign n3793 = n3791 & n3792;
  assign n3794 = ~n675 & ~n682;
  assign n3795 = ~n702 & n3794;
  assign n3796 = ~n182 & ~n208;
  assign n3797 = ~n599 & n3796;
  assign n3798 = n1342 & n1394;
  assign n3799 = n2150 & n2597;
  assign n3800 = n2695 & n3401;
  assign n3801 = n3799 & n3800;
  assign n3802 = n3797 & n3798;
  assign n3803 = n3795 & n3802;
  assign n3804 = n3781 & n3801;
  assign n3805 = n3803 & n3804;
  assign n3806 = n3793 & n3805;
  assign n3807 = ~n209 & ~n587;
  assign n3808 = ~n192 & n3807;
  assign n3809 = ~n183 & ~n242;
  assign n3810 = ~n243 & ~n355;
  assign n3811 = ~n577 & n3810;
  assign n3812 = n461 & n3809;
  assign n3813 = n596 & n624;
  assign n3814 = n904 & n2634;
  assign n3815 = n3170 & n3763;
  assign n3816 = n3814 & n3815;
  assign n3817 = n3812 & n3813;
  assign n3818 = n1345 & n3811;
  assign n3819 = n3808 & n3818;
  assign n3820 = n3816 & n3817;
  assign n3821 = n3769 & n3820;
  assign n3822 = n3777 & n3819;
  assign n3823 = n3821 & n3822;
  assign n3824 = n3806 & n3823;
  assign n3825 = n2292 & n3824;
  assign n3826 = ~n240 & ~n363;
  assign n3827 = ~n109 & ~n425;
  assign n3828 = n3826 & n3827;
  assign n3829 = ~n218 & ~n343;
  assign n3830 = ~n536 & n3829;
  assign n3831 = n524 & n3830;
  assign n3832 = ~n208 & ~n238;
  assign n3833 = ~n297 & ~n459;
  assign n3834 = n3832 & n3833;
  assign n3835 = n1077 & n1121;
  assign n3836 = n3834 & n3835;
  assign n3837 = n3828 & n3836;
  assign n3838 = n3831 & n3837;
  assign n3839 = ~n141 & ~n165;
  assign n3840 = ~n479 & n3839;
  assign n3841 = n573 & n3840;
  assign n3842 = ~n289 & ~n687;
  assign n3843 = ~n602 & ~n686;
  assign n3844 = ~n126 & ~n244;
  assign n3845 = ~n522 & ~n651;
  assign n3846 = ~n267 & ~n316;
  assign n3847 = ~n324 & ~n376;
  assign n3848 = ~n391 & ~n700;
  assign n3849 = n3847 & n3848;
  assign n3850 = n2194 & n3846;
  assign n3851 = n2424 & n3850;
  assign n3852 = n3849 & n3851;
  assign n3853 = ~n327 & ~n480;
  assign n3854 = ~n591 & n3853;
  assign n3855 = ~n167 & ~n245;
  assign n3856 = ~n463 & ~n554;
  assign n3857 = ~n650 & ~n673;
  assign n3858 = n3856 & n3857;
  assign n3859 = n1014 & n1237;
  assign n3860 = n1354 & n2220;
  assign n3861 = n3842 & n3843;
  assign n3862 = n3844 & n3845;
  assign n3863 = n3855 & n3862;
  assign n3864 = n3860 & n3861;
  assign n3865 = n3858 & n3859;
  assign n3866 = n3854 & n3865;
  assign n3867 = n3863 & n3864;
  assign n3868 = n3866 & n3867;
  assign n3869 = n3852 & n3868;
  assign n3870 = ~n243 & ~n462;
  assign n3871 = n2005 & n3870;
  assign n3872 = ~n133 & ~n221;
  assign n3873 = ~n253 & ~n420;
  assign n3874 = ~n421 & ~n587;
  assign n3875 = n3873 & n3874;
  assign n3876 = n1041 & n1267;
  assign n3877 = n1355 & n2063;
  assign n3878 = n2297 & n3071;
  assign n3879 = n3872 & n3878;
  assign n3880 = n3876 & n3877;
  assign n3881 = n3871 & n3875;
  assign n3882 = n3880 & n3881;
  assign n3883 = n3841 & n3879;
  assign n3884 = n3882 & n3883;
  assign n3885 = n3838 & n3884;
  assign n3886 = n3418 & n3885;
  assign n3887 = n3869 & n3886;
  assign n3888 = ~n3825 & ~n3887;
  assign n3889 = n3825 & n3887;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = ~pi26  & n3890;
  assign n3892 = ~n3888 & ~n3891;
  assign n3893 = n3761 & ~n3892;
  assign n3894 = ~n3761 & n3892;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = ~pi31  & ~n565;
  assign n3897 = ~n729 & n3896;
  assign n3898 = ~n802 & n3683;
  assign n3899 = n564 & ~n898;
  assign n3900 = n3580 & ~n3582;
  assign n3901 = ~n3583 & ~n3900;
  assign n3902 = n566 & n3901;
  assign n3903 = ~n3898 & ~n3899;
  assign n3904 = ~n3897 & n3903;
  assign n3905 = ~n3902 & n3904;
  assign n3906 = n3895 & ~n3905;
  assign n3907 = ~n3893 & ~n3906;
  assign n3908 = ~n3655 & n3761;
  assign n3909 = ~n3762 & ~n3908;
  assign n3910 = ~n3907 & n3909;
  assign n3911 = ~n3762 & ~n3910;
  assign n3912 = pi29  & ~n3673;
  assign n3913 = ~n3674 & ~n3912;
  assign n3914 = ~n3911 & n3913;
  assign n3915 = n3911 & ~n3913;
  assign n3916 = ~n3914 & ~n3915;
  assign n3917 = n564 & ~n729;
  assign n3918 = ~n621 & n3683;
  assign n3919 = ~n563 & n3896;
  assign n3920 = n3588 & ~n3591;
  assign n3921 = ~n3592 & ~n3920;
  assign n3922 = n566 & n3921;
  assign n3923 = ~n3918 & ~n3919;
  assign n3924 = ~n3917 & n3923;
  assign n3925 = ~n3922 & n3924;
  assign n3926 = n3916 & ~n3925;
  assign n3927 = ~n3914 & ~n3926;
  assign n3928 = ~n3678 & n3690;
  assign n3929 = ~n3691 & ~n3928;
  assign n3930 = ~n3927 & n3929;
  assign n3931 = n3927 & ~n3929;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = ~n3916 & n3925;
  assign n3934 = ~n3926 & ~n3933;
  assign n3935 = ~pi28  & ~pi29 ;
  assign n3936 = pi28  & pi29 ;
  assign n3937 = ~n3935 & ~n3936;
  assign n3938 = ~n79 & ~n106;
  assign n3939 = ~pi26  & ~pi27 ;
  assign n3940 = pi26  & pi27 ;
  assign n3941 = ~n3939 & ~n3940;
  assign n3942 = ~n3938 & ~n3941;
  assign n3943 = n3937 & n3942;
  assign n3944 = n3937 & n3941;
  assign n3945 = ~n3593 & n3944;
  assign n3946 = ~n3943 & ~n3945;
  assign n3947 = ~n563 & ~n3946;
  assign n3948 = ~pi29  & n3947;
  assign n3949 = pi29  & ~n3947;
  assign n3950 = ~n3948 & ~n3949;
  assign n3951 = ~n621 & n3896;
  assign n3952 = ~n729 & n3683;
  assign n3953 = n564 & ~n802;
  assign n3954 = n3584 & ~n3586;
  assign n3955 = ~n3587 & ~n3954;
  assign n3956 = n566 & n3955;
  assign n3957 = ~n3951 & ~n3953;
  assign n3958 = ~n3952 & n3957;
  assign n3959 = ~n3956 & n3958;
  assign n3960 = n3950 & n3959;
  assign n3961 = n3907 & ~n3909;
  assign n3962 = ~n3910 & ~n3961;
  assign n3963 = ~n3950 & ~n3959;
  assign n3964 = ~n3960 & ~n3963;
  assign n3965 = ~n3962 & n3964;
  assign n3966 = ~n3960 & ~n3965;
  assign n3967 = n3934 & n3966;
  assign n3968 = n3962 & ~n3964;
  assign n3969 = ~n3965 & ~n3968;
  assign n3970 = ~n180 & ~n280;
  assign n3971 = ~n312 & n3970;
  assign n3972 = ~n224 & ~n390;
  assign n3973 = ~n690 & n3972;
  assign n3974 = ~n195 & ~n290;
  assign n3975 = ~n644 & ~n650;
  assign n3976 = ~n682 & n3975;
  assign n3977 = n2868 & n3974;
  assign n3978 = n3976 & n3977;
  assign n3979 = n3973 & n3978;
  assign n3980 = ~n238 & ~n388;
  assign n3981 = ~n572 & n3980;
  assign n3982 = ~n172 & ~n203;
  assign n3983 = ~n379 & ~n492;
  assign n3984 = n3982 & n3983;
  assign n3985 = n211 & n436;
  assign n3986 = n967 & n2092;
  assign n3987 = n2296 & n3986;
  assign n3988 = n3984 & n3985;
  assign n3989 = n1504 & n3981;
  assign n3990 = n3988 & n3989;
  assign n3991 = n3987 & n3990;
  assign n3992 = ~n299 & ~n340;
  assign n3993 = ~n494 & n3992;
  assign n3994 = ~n173 & ~n427;
  assign n3995 = ~n282 & ~n479;
  assign n3996 = ~n175 & ~n270;
  assign n3997 = n703 & n3996;
  assign n3998 = n3995 & n3997;
  assign n3999 = ~n202 & ~n319;
  assign n4000 = ~n472 & n3999;
  assign n4001 = n194 & n2942;
  assign n4002 = n2953 & n3205;
  assign n4003 = n3994 & n4002;
  assign n4004 = n4000 & n4001;
  assign n4005 = n3993 & n4004;
  assign n4006 = n2277 & n4003;
  assign n4007 = n3998 & n4006;
  assign n4008 = n3979 & n4005;
  assign n4009 = n4007 & n4008;
  assign n4010 = n3991 & n4009;
  assign n4011 = ~n316 & ~n424;
  assign n4012 = ~n601 & n4011;
  assign n4013 = ~n212 & ~n326;
  assign n4014 = ~n384 & ~n389;
  assign n4015 = ~n447 & ~n570;
  assign n4016 = ~n689 & n4015;
  assign n4017 = n4013 & n4014;
  assign n4018 = n137 & n461;
  assign n4019 = n4017 & n4018;
  assign n4020 = n4012 & n4016;
  assign n4021 = n4019 & n4020;
  assign n4022 = n1557 & n4021;
  assign n4023 = ~n149 & ~n536;
  assign n4024 = ~n553 & ~n582;
  assign n4025 = n4023 & n4024;
  assign n4026 = n540 & n738;
  assign n4027 = n2475 & n3855;
  assign n4028 = n4026 & n4027;
  assign n4029 = n1908 & n4025;
  assign n4030 = n3971 & n4029;
  assign n4031 = n4028 & n4030;
  assign n4032 = n4010 & n4031;
  assign n4033 = n4022 & n4032;
  assign n4034 = n3825 & ~n4033;
  assign n4035 = ~n3825 & n4033;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = ~n898 & n3896;
  assign n4038 = ~n1006 & n3683;
  assign n4039 = n564 & ~n1107;
  assign n4040 = n3572 & ~n3574;
  assign n4041 = ~n3575 & ~n4040;
  assign n4042 = n566 & n4041;
  assign n4043 = ~n4037 & ~n4038;
  assign n4044 = ~n4039 & n4043;
  assign n4045 = ~n4042 & n4044;
  assign n4046 = n4036 & ~n4045;
  assign n4047 = ~n4034 & ~n4046;
  assign n4048 = pi26  & ~n3890;
  assign n4049 = ~n3891 & ~n4048;
  assign n4050 = ~n4047 & n4049;
  assign n4051 = n4047 & ~n4049;
  assign n4052 = ~n4050 & ~n4051;
  assign n4053 = ~n802 & n3896;
  assign n4054 = ~n898 & n3683;
  assign n4055 = n564 & ~n1006;
  assign n4056 = n3576 & ~n3578;
  assign n4057 = ~n3579 & ~n4056;
  assign n4058 = n566 & n4057;
  assign n4059 = ~n4053 & ~n4054;
  assign n4060 = ~n4055 & n4059;
  assign n4061 = ~n4058 & n4060;
  assign n4062 = n4052 & ~n4061;
  assign n4063 = ~n4050 & ~n4062;
  assign n4064 = ~n3895 & n3905;
  assign n4065 = ~n3906 & ~n4064;
  assign n4066 = n4063 & ~n4065;
  assign n4067 = ~n4063 & n4065;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = ~n621 & n3943;
  assign n4070 = n3938 & ~n3941;
  assign n4071 = ~n563 & n4070;
  assign n4072 = n3687 & n3944;
  assign n4073 = ~n4069 & ~n4071;
  assign n4074 = ~n4072 & n4073;
  assign n4075 = pi29  & n4074;
  assign n4076 = ~pi29  & ~n4074;
  assign n4077 = ~n4075 & ~n4076;
  assign n4078 = n4068 & n4077;
  assign n4079 = ~n4066 & ~n4078;
  assign n4080 = ~n3969 & n4079;
  assign n4081 = ~n4068 & ~n4077;
  assign n4082 = ~n4078 & ~n4081;
  assign n4083 = ~n145 & ~n218;
  assign n4084 = ~n473 & ~n572;
  assign n4085 = ~n674 & n4084;
  assign n4086 = n4083 & n4085;
  assign n4087 = ~n180 & ~n222;
  assign n4088 = ~n276 & ~n407;
  assign n4089 = ~n640 & n4088;
  assign n4090 = n3034 & n4087;
  assign n4091 = n4089 & n4090;
  assign n4092 = ~n118 & n464;
  assign n4093 = ~n207 & ~n315;
  assign n4094 = ~n125 & ~n247;
  assign n4095 = ~n308 & ~n356;
  assign n4096 = ~n667 & n4095;
  assign n4097 = n1078 & n4094;
  assign n4098 = n1263 & n2831;
  assign n4099 = n4093 & n4098;
  assign n4100 = n4096 & n4097;
  assign n4101 = n1111 & n2222;
  assign n4102 = n4100 & n4101;
  assign n4103 = n4099 & n4102;
  assign n4104 = ~n335 & ~n690;
  assign n4105 = ~n279 & ~n282;
  assign n4106 = ~n321 & ~n541;
  assign n4107 = n4105 & n4106;
  assign n4108 = n1116 & n2129;
  assign n4109 = n4104 & n4108;
  assign n4110 = n4107 & n4109;
  assign n4111 = ~n251 & ~n427;
  assign n4112 = ~n445 & ~n583;
  assign n4113 = ~n598 & n4112;
  assign n4114 = n194 & n4111;
  assign n4115 = n3872 & n4114;
  assign n4116 = n4113 & n4115;
  assign n4117 = ~n103 & ~n235;
  assign n4118 = ~n426 & ~n510;
  assign n4119 = ~n542 & n4118;
  assign n4120 = n1392 & n4117;
  assign n4121 = n2540 & n4120;
  assign n4122 = n4092 & n4119;
  assign n4123 = n4121 & n4122;
  assign n4124 = n3261 & n4123;
  assign n4125 = n4110 & n4116;
  assign n4126 = n4124 & n4125;
  assign n4127 = n4103 & n4126;
  assign n4128 = ~n216 & ~n391;
  assign n4129 = n2234 & n4128;
  assign n4130 = ~n203 & ~n265;
  assign n4131 = ~n269 & ~n536;
  assign n4132 = ~n666 & ~n702;
  assign n4133 = n4131 & n4132;
  assign n4134 = n523 & n4130;
  assign n4135 = n1679 & n2220;
  assign n4136 = n2706 & n4135;
  assign n4137 = n4133 & n4134;
  assign n4138 = n3077 & n4129;
  assign n4139 = n4137 & n4138;
  assign n4140 = n4086 & n4136;
  assign n4141 = n4091 & n4140;
  assign n4142 = n2074 & n4139;
  assign n4143 = n4141 & n4142;
  assign n4144 = n4127 & n4143;
  assign n4145 = n864 & n1246;
  assign n4146 = n2903 & n4145;
  assign n4147 = ~n122 & ~n335;
  assign n4148 = ~n425 & n4147;
  assign n4149 = n1301 & n4148;
  assign n4150 = ~n221 & ~n364;
  assign n4151 = ~n667 & n4150;
  assign n4152 = n137 & n3282;
  assign n4153 = n4151 & n4152;
  assign n4154 = n4146 & n4153;
  assign n4155 = n4149 & n4154;
  assign n4156 = ~n510 & ~n679;
  assign n4157 = ~n277 & ~n661;
  assign n4158 = n341 & n4157;
  assign n4159 = n449 & n1910;
  assign n4160 = n4158 & n4159;
  assign n4161 = ~n238 & ~n251;
  assign n4162 = ~n215 & ~n542;
  assign n4163 = ~n195 & ~n379;
  assign n4164 = ~n390 & ~n572;
  assign n4165 = n4163 & n4164;
  assign n4166 = ~n460 & ~n545;
  assign n4167 = n268 & n4166;
  assign n4168 = n408 & n743;
  assign n4169 = n928 & n1485;
  assign n4170 = n1666 & n1712;
  assign n4171 = n4161 & n4162;
  assign n4172 = n4170 & n4171;
  assign n4173 = n4168 & n4169;
  assign n4174 = n3795 & n4167;
  assign n4175 = n4165 & n4174;
  assign n4176 = n4172 & n4173;
  assign n4177 = n1019 & n4176;
  assign n4178 = n4175 & n4177;
  assign n4179 = ~n175 & ~n495;
  assign n4180 = ~n595 & ~n666;
  assign n4181 = ~n689 & n4180;
  assign n4182 = n1343 & n4179;
  assign n4183 = n1614 & n1710;
  assign n4184 = n1760 & n2096;
  assign n4185 = n2424 & n2754;
  assign n4186 = n4184 & n4185;
  assign n4187 = n4182 & n4183;
  assign n4188 = n4181 & n4187;
  assign n4189 = n1245 & n4186;
  assign n4190 = n3831 & n4160;
  assign n4191 = n4189 & n4190;
  assign n4192 = n2311 & n4188;
  assign n4193 = n4191 & n4192;
  assign n4194 = n4178 & n4193;
  assign n4195 = ~n164 & ~n472;
  assign n4196 = ~n212 & ~n597;
  assign n4197 = ~n680 & ~n701;
  assign n4198 = n4196 & n4197;
  assign n4199 = n2300 & n3627;
  assign n4200 = n4195 & n4199;
  assign n4201 = n4198 & n4200;
  assign n4202 = ~n168 & ~n546;
  assign n4203 = ~n569 & ~n646;
  assign n4204 = n4202 & n4203;
  assign n4205 = ~n125 & ~n148;
  assign n4206 = ~n279 & ~n285;
  assign n4207 = ~n445 & ~n483;
  assign n4208 = ~n574 & ~n587;
  assign n4209 = ~n650 & n4208;
  assign n4210 = n4206 & n4207;
  assign n4211 = n1393 & n4205;
  assign n4212 = n4156 & n4211;
  assign n4213 = n4209 & n4210;
  assign n4214 = n1683 & n4204;
  assign n4215 = n4213 & n4214;
  assign n4216 = n1958 & n4212;
  assign n4217 = n4215 & n4216;
  assign n4218 = n4201 & n4217;
  assign n4219 = n4155 & n4218;
  assign n4220 = n4194 & n4219;
  assign n4221 = ~n4144 & ~n4220;
  assign n4222 = n4144 & n4220;
  assign n4223 = ~n4221 & ~n4222;
  assign n4224 = ~pi23  & n4223;
  assign n4225 = ~n4221 & ~n4224;
  assign n4226 = n3825 & ~n4225;
  assign n4227 = ~n3825 & n4225;
  assign n4228 = ~n4226 & ~n4227;
  assign n4229 = ~n1107 & n3683;
  assign n4230 = ~n1006 & n3896;
  assign n4231 = n564 & ~n1230;
  assign n4232 = n3568 & ~n3570;
  assign n4233 = ~n3571 & ~n4232;
  assign n4234 = n566 & n4233;
  assign n4235 = ~n4229 & ~n4230;
  assign n4236 = ~n4231 & n4235;
  assign n4237 = ~n4234 & n4236;
  assign n4238 = n4228 & ~n4237;
  assign n4239 = ~n4226 & ~n4238;
  assign n4240 = ~n4036 & n4045;
  assign n4241 = ~n4046 & ~n4240;
  assign n4242 = ~n4239 & n4241;
  assign n4243 = n4239 & ~n4241;
  assign n4244 = ~n4242 & ~n4243;
  assign n4245 = pi23  & ~n4223;
  assign n4246 = ~n4224 & ~n4245;
  assign n4247 = ~n1230 & n3683;
  assign n4248 = n564 & ~n1337;
  assign n4249 = ~n1107 & n3896;
  assign n4250 = n3564 & ~n3566;
  assign n4251 = ~n3567 & ~n4250;
  assign n4252 = n566 & n4251;
  assign n4253 = ~n4247 & ~n4248;
  assign n4254 = ~n4249 & n4253;
  assign n4255 = ~n4252 & n4254;
  assign n4256 = n4246 & ~n4255;
  assign n4257 = ~n267 & ~n271;
  assign n4258 = ~n674 & n4257;
  assign n4259 = ~n126 & ~n391;
  assign n4260 = ~n644 & ~n689;
  assign n4261 = n4259 & n4260;
  assign n4262 = n2061 & n4261;
  assign n4263 = n4258 & n4262;
  assign n4264 = ~n148 & ~n598;
  assign n4265 = ~n277 & ~n311;
  assign n4266 = ~n323 & ~n700;
  assign n4267 = ~n125 & ~n363;
  assign n4268 = ~n541 & n2373;
  assign n4269 = n3624 & n4267;
  assign n4270 = n4268 & n4269;
  assign n4271 = n3403 & n4270;
  assign n4272 = ~n336 & ~n553;
  assign n4273 = ~n591 & n4272;
  assign n4274 = ~n279 & ~n571;
  assign n4275 = ~n131 & ~n270;
  assign n4276 = ~n401 & n4275;
  assign n4277 = n742 & n840;
  assign n4278 = n885 & n1354;
  assign n4279 = n4266 & n4274;
  assign n4280 = n4278 & n4279;
  assign n4281 = n2610 & n4277;
  assign n4282 = n4273 & n4276;
  assign n4283 = n4281 & n4282;
  assign n4284 = n4280 & n4283;
  assign n4285 = n4271 & n4284;
  assign n4286 = ~n406 & ~n578;
  assign n4287 = ~n585 & n4286;
  assign n4288 = n741 & n4287;
  assign n4289 = ~n422 & ~n642;
  assign n4290 = ~n673 & n4289;
  assign n4291 = n1203 & n1457;
  assign n4292 = n1631 & n2190;
  assign n4293 = n4264 & n4265;
  assign n4294 = n4292 & n4293;
  assign n4295 = n4290 & n4291;
  assign n4296 = n4294 & n4295;
  assign n4297 = n1454 & n4288;
  assign n4298 = n4296 & n4297;
  assign n4299 = n4263 & n4298;
  assign n4300 = n1753 & n4299;
  assign n4301 = n3024 & n4285;
  assign n4302 = n4300 & n4301;
  assign n4303 = n4144 & ~n4302;
  assign n4304 = ~n109 & ~n343;
  assign n4305 = ~n466 & ~n568;
  assign n4306 = ~n585 & n4305;
  assign n4307 = n1115 & n4304;
  assign n4308 = n1679 & n2871;
  assign n4309 = n4307 & n4308;
  assign n4310 = n3713 & n4306;
  assign n4311 = n4309 & n4310;
  assign n4312 = ~n244 & ~n269;
  assign n4313 = ~n365 & ~n385;
  assign n4314 = ~n463 & ~n511;
  assign n4315 = n4313 & n4314;
  assign n4316 = n461 & n4312;
  assign n4317 = n781 & n1458;
  assign n4318 = n2566 & n3778;
  assign n4319 = n4317 & n4318;
  assign n4320 = n4315 & n4316;
  assign n4321 = n4258 & n4320;
  assign n4322 = n4319 & n4321;
  assign n4323 = n2638 & n4311;
  assign n4324 = n4322 & n4323;
  assign n4325 = n1380 & n1472;
  assign n4326 = ~n363 & n2980;
  assign n4327 = ~n85 & ~n207;
  assign n4328 = ~n222 & n4327;
  assign n4329 = n592 & n2945;
  assign n4330 = n4328 & n4329;
  assign n4331 = ~n405 & ~n480;
  assign n4332 = ~n553 & n4331;
  assign n4333 = n237 & n298;
  assign n4334 = n920 & n929;
  assign n4335 = n2220 & n4334;
  assign n4336 = n4332 & n4333;
  assign n4337 = n817 & n2062;
  assign n4338 = n3345 & n4337;
  assign n4339 = n4335 & n4336;
  assign n4340 = n4326 & n4330;
  assign n4341 = n4339 & n4340;
  assign n4342 = n4338 & n4341;
  assign n4343 = ~n221 & ~n276;
  assign n4344 = ~n472 & ~n650;
  assign n4345 = n4343 & n4344;
  assign n4346 = n924 & n1125;
  assign n4347 = n1433 & n1594;
  assign n4348 = n1762 & n2150;
  assign n4349 = n2754 & n4348;
  assign n4350 = n4346 & n4347;
  assign n4351 = n669 & n4345;
  assign n4352 = n4325 & n4351;
  assign n4353 = n4349 & n4350;
  assign n4354 = n4352 & n4353;
  assign n4355 = n1901 & n4354;
  assign n4356 = n2321 & n4355;
  assign n4357 = n4324 & n4342;
  assign n4358 = n4356 & n4357;
  assign n4359 = ~n92 & n1431;
  assign n4360 = ~n388 & ~n584;
  assign n4361 = ~n689 & n4360;
  assign n4362 = ~n147 & ~n221;
  assign n4363 = ~n277 & ~n308;
  assign n4364 = ~n447 & ~n577;
  assign n4365 = ~n701 & n4364;
  assign n4366 = n4362 & n4363;
  assign n4367 = n555 & n759;
  assign n4368 = n853 & n1432;
  assign n4369 = n4367 & n4368;
  assign n4370 = n4365 & n4366;
  assign n4371 = n4369 & n4370;
  assign n4372 = ~n239 & ~n253;
  assign n4373 = ~n287 & ~n546;
  assign n4374 = n4372 & n4373;
  assign n4375 = n1689 & n2097;
  assign n4376 = n4374 & n4375;
  assign n4377 = n1239 & n4359;
  assign n4378 = n4361 & n4377;
  assign n4379 = n4376 & n4378;
  assign n4380 = n2304 & n4371;
  assign n4381 = n4379 & n4380;
  assign n4382 = ~n389 & n827;
  assign n4383 = ~n279 & ~n362;
  assign n4384 = ~n459 & ~n686;
  assign n4385 = ~n149 & ~n572;
  assign n4386 = n4156 & n4385;
  assign n4387 = ~n319 & ~n326;
  assign n4388 = ~n375 & n4387;
  assign n4389 = n1785 & n3379;
  assign n4390 = n4388 & n4389;
  assign n4391 = ~n580 & ~n645;
  assign n4392 = n493 & n4391;
  assign n4393 = n741 & n919;
  assign n4394 = n1380 & n1631;
  assign n4395 = n1907 & n1965;
  assign n4396 = n2981 & n4383;
  assign n4397 = n4384 & n4396;
  assign n4398 = n4394 & n4395;
  assign n4399 = n4392 & n4393;
  assign n4400 = n4386 & n4399;
  assign n4401 = n4397 & n4398;
  assign n4402 = n4382 & n4390;
  assign n4403 = n4401 & n4402;
  assign n4404 = n4400 & n4403;
  assign n4405 = ~n271 & ~n296;
  assign n4406 = ~n103 & ~n163;
  assign n4407 = ~n236 & ~n243;
  assign n4408 = ~n288 & ~n360;
  assign n4409 = ~n521 & ~n543;
  assign n4410 = ~n571 & ~n651;
  assign n4411 = ~n665 & n4410;
  assign n4412 = n4408 & n4409;
  assign n4413 = n4406 & n4407;
  assign n4414 = n603 & n4405;
  assign n4415 = n4413 & n4414;
  assign n4416 = n4411 & n4412;
  assign n4417 = n4415 & n4416;
  assign n4418 = ~n426 & ~n470;
  assign n4419 = ~n85 & ~n280;
  assign n4420 = ~n379 & n4419;
  assign n4421 = ~n134 & ~n173;
  assign n4422 = ~n511 & n4421;
  assign n4423 = n481 & n3154;
  assign n4424 = n4418 & n4423;
  assign n4425 = n4420 & n4422;
  assign n4426 = n4424 & n4425;
  assign n4427 = ~n240 & ~n448;
  assign n4428 = ~n466 & ~n591;
  assign n4429 = n4427 & n4428;
  assign n4430 = n1015 & n1116;
  assign n4431 = n1344 & n1538;
  assign n4432 = n4430 & n4431;
  assign n4433 = n3028 & n4429;
  assign n4434 = n4432 & n4433;
  assign n4435 = n918 & n4434;
  assign n4436 = n4417 & n4426;
  assign n4437 = n4435 & n4436;
  assign n4438 = n4381 & n4437;
  assign n4439 = n4404 & n4438;
  assign n4440 = ~n4358 & ~n4439;
  assign n4441 = n4358 & n4439;
  assign n4442 = ~n4440 & ~n4441;
  assign n4443 = ~pi20  & n4442;
  assign n4444 = ~n4440 & ~n4443;
  assign n4445 = n4302 & ~n4444;
  assign n4446 = ~n4302 & n4444;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = n564 & ~n1532;
  assign n4449 = ~n1425 & n3683;
  assign n4450 = ~n1337 & n3896;
  assign n4451 = n3556 & ~n3558;
  assign n4452 = ~n3559 & ~n4451;
  assign n4453 = n566 & n4452;
  assign n4454 = ~n4448 & ~n4449;
  assign n4455 = ~n4450 & n4454;
  assign n4456 = ~n4453 & n4455;
  assign n4457 = n4447 & ~n4456;
  assign n4458 = ~n4445 & ~n4457;
  assign n4459 = ~n4144 & n4302;
  assign n4460 = ~n4303 & ~n4459;
  assign n4461 = ~n4458 & n4460;
  assign n4462 = ~n4303 & ~n4461;
  assign n4463 = ~n4246 & n4255;
  assign n4464 = ~n4256 & ~n4463;
  assign n4465 = ~n4462 & n4464;
  assign n4466 = ~n4256 & ~n4465;
  assign n4467 = ~n4228 & n4237;
  assign n4468 = ~n4238 & ~n4467;
  assign n4469 = ~n4466 & n4468;
  assign n4470 = n4466 & ~n4468;
  assign n4471 = ~n4469 & ~n4470;
  assign n4472 = ~n3937 & n3941;
  assign n4473 = ~n729 & n4472;
  assign n4474 = ~n802 & n4070;
  assign n4475 = ~n898 & n3943;
  assign n4476 = n3901 & n3944;
  assign n4477 = ~n4474 & ~n4475;
  assign n4478 = ~n4473 & n4477;
  assign n4479 = ~n4476 & n4478;
  assign n4480 = pi29  & n4479;
  assign n4481 = ~pi29  & ~n4479;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = n4471 & ~n4482;
  assign n4484 = ~n4469 & ~n4483;
  assign n4485 = n4244 & ~n4484;
  assign n4486 = ~n4242 & ~n4485;
  assign n4487 = ~n4052 & n4061;
  assign n4488 = ~n4062 & ~n4487;
  assign n4489 = ~n4486 & n4488;
  assign n4490 = ~n729 & n3943;
  assign n4491 = ~n621 & n4070;
  assign n4492 = ~n563 & n4472;
  assign n4493 = n3921 & n3944;
  assign n4494 = ~n4491 & ~n4492;
  assign n4495 = ~n4490 & n4494;
  assign n4496 = ~n4493 & n4495;
  assign n4497 = pi29  & n4496;
  assign n4498 = ~pi29  & ~n4496;
  assign n4499 = ~n4497 & ~n4498;
  assign n4500 = n4486 & ~n4488;
  assign n4501 = ~n4489 & ~n4500;
  assign n4502 = ~n4499 & n4501;
  assign n4503 = ~n4489 & ~n4502;
  assign n4504 = ~n4082 & ~n4503;
  assign n4505 = n4082 & n4503;
  assign n4506 = ~n4504 & ~n4505;
  assign n4507 = ~pi25  & pi26 ;
  assign n4508 = pi25  & ~pi26 ;
  assign n4509 = ~n4507 & ~n4508;
  assign n4510 = pi23  & ~pi24 ;
  assign n4511 = ~pi23  & pi24 ;
  assign n4512 = ~n4510 & ~n4511;
  assign n4513 = ~n99 & ~n123;
  assign n4514 = n4512 & ~n4513;
  assign n4515 = ~n4509 & n4514;
  assign n4516 = ~n4509 & ~n4512;
  assign n4517 = ~n3593 & n4516;
  assign n4518 = ~n4515 & ~n4517;
  assign n4519 = ~n563 & ~n4518;
  assign n4520 = ~pi26  & n4519;
  assign n4521 = pi26  & ~n4519;
  assign n4522 = ~n4520 & ~n4521;
  assign n4523 = ~n621 & n4472;
  assign n4524 = ~n729 & n4070;
  assign n4525 = ~n802 & n3943;
  assign n4526 = n3944 & n3955;
  assign n4527 = ~n4523 & ~n4525;
  assign n4528 = ~n4524 & n4527;
  assign n4529 = ~n4526 & n4528;
  assign n4530 = pi29  & n4529;
  assign n4531 = ~pi29  & ~n4529;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = ~n4522 & ~n4532;
  assign n4534 = ~n4244 & n4484;
  assign n4535 = ~n4485 & ~n4534;
  assign n4536 = n4522 & n4532;
  assign n4537 = ~n4533 & ~n4536;
  assign n4538 = n4535 & n4537;
  assign n4539 = ~n4533 & ~n4538;
  assign n4540 = n4499 & ~n4501;
  assign n4541 = ~n4502 & ~n4540;
  assign n4542 = ~n4539 & n4541;
  assign n4543 = n4458 & ~n4460;
  assign n4544 = ~n4461 & ~n4543;
  assign n4545 = ~n1337 & n3683;
  assign n4546 = n564 & ~n1425;
  assign n4547 = ~n1230 & n3896;
  assign n4548 = n3560 & ~n3562;
  assign n4549 = ~n3563 & ~n4548;
  assign n4550 = n566 & n4549;
  assign n4551 = ~n4545 & ~n4546;
  assign n4552 = ~n4547 & n4551;
  assign n4553 = ~n4550 & n4552;
  assign n4554 = n4544 & ~n4553;
  assign n4555 = n1469 & n1689;
  assign n4556 = ~n109 & ~n212;
  assign n4557 = ~n242 & ~n379;
  assign n4558 = ~n546 & ~n683;
  assign n4559 = n4557 & n4558;
  assign n4560 = n471 & n4556;
  assign n4561 = n4559 & n4560;
  assign n4562 = ~n280 & ~n323;
  assign n4563 = ~n144 & ~n199;
  assign n4564 = ~n356 & ~n406;
  assign n4565 = ~n577 & n4564;
  assign n4566 = n1626 & n4563;
  assign n4567 = n4562 & n4566;
  assign n4568 = n4565 & n4567;
  assign n4569 = ~n175 & ~n209;
  assign n4570 = ~n570 & n4569;
  assign n4571 = n738 & n2272;
  assign n4572 = n4570 & n4571;
  assign n4573 = n1205 & n1763;
  assign n4574 = n3731 & n4555;
  assign n4575 = n4573 & n4574;
  assign n4576 = n4561 & n4572;
  assign n4577 = n4575 & n4576;
  assign n4578 = n4568 & n4577;
  assign n4579 = ~n447 & n1907;
  assign n4580 = n1970 & n4579;
  assign n4581 = ~n384 & ~n580;
  assign n4582 = n2230 & n4581;
  assign n4583 = ~n463 & n2009;
  assign n4584 = n437 & n4583;
  assign n4585 = ~n267 & ~n279;
  assign n4586 = ~n355 & ~n543;
  assign n4587 = ~n554 & ~n590;
  assign n4588 = ~n649 & n4587;
  assign n4589 = n4585 & n4586;
  assign n4590 = n3352 & n4589;
  assign n4591 = n4588 & n4590;
  assign n4592 = ~n131 & ~n569;
  assign n4593 = ~n571 & ~n674;
  assign n4594 = n4592 & n4593;
  assign n4595 = n940 & n1376;
  assign n4596 = n1714 & n1808;
  assign n4597 = n4595 & n4596;
  assign n4598 = n972 & n4594;
  assign n4599 = n1270 & n4598;
  assign n4600 = n4580 & n4597;
  assign n4601 = n4582 & n4584;
  assign n4602 = n4600 & n4601;
  assign n4603 = n4591 & n4599;
  assign n4604 = n4602 & n4603;
  assign n4605 = ~n312 & ~n538;
  assign n4606 = ~n644 & n4605;
  assign n4607 = ~n290 & ~n318;
  assign n4608 = n1112 & n4607;
  assign n4609 = n1631 & n1910;
  assign n4610 = n4093 & n4609;
  assign n4611 = n4606 & n4608;
  assign n4612 = n4610 & n4611;
  assign n4613 = n1755 & n2665;
  assign n4614 = n4612 & n4613;
  assign n4615 = n1430 & n2914;
  assign n4616 = n4614 & n4615;
  assign n4617 = n4578 & n4616;
  assign n4618 = n4604 & n4617;
  assign n4619 = n4358 & ~n4618;
  assign n4620 = ~n4358 & n4618;
  assign n4621 = ~n4619 & ~n4620;
  assign n4622 = n564 & ~n1737;
  assign n4623 = ~n1610 & n3683;
  assign n4624 = ~n1532 & n3896;
  assign n4625 = n3548 & ~n3550;
  assign n4626 = ~n3551 & ~n4625;
  assign n4627 = n566 & n4626;
  assign n4628 = ~n4622 & ~n4623;
  assign n4629 = ~n4624 & n4628;
  assign n4630 = ~n4627 & n4629;
  assign n4631 = n4621 & ~n4630;
  assign n4632 = ~n4619 & ~n4631;
  assign n4633 = pi20  & ~n4442;
  assign n4634 = ~n4443 & ~n4633;
  assign n4635 = ~n4632 & n4634;
  assign n4636 = n4632 & ~n4634;
  assign n4637 = ~n4635 & ~n4636;
  assign n4638 = n564 & ~n1610;
  assign n4639 = ~n1532 & n3683;
  assign n4640 = ~n1425 & n3896;
  assign n4641 = n3552 & ~n3554;
  assign n4642 = ~n3555 & ~n4641;
  assign n4643 = n566 & n4642;
  assign n4644 = ~n4638 & ~n4639;
  assign n4645 = ~n4640 & n4644;
  assign n4646 = ~n4643 & n4645;
  assign n4647 = n4637 & ~n4646;
  assign n4648 = ~n4635 & ~n4647;
  assign n4649 = ~n4447 & n4456;
  assign n4650 = ~n4457 & ~n4649;
  assign n4651 = ~n4648 & n4650;
  assign n4652 = n4648 & ~n4650;
  assign n4653 = ~n4651 & ~n4652;
  assign n4654 = ~n1107 & n4070;
  assign n4655 = ~n1006 & n4472;
  assign n4656 = ~n1230 & n3943;
  assign n4657 = n3944 & n4233;
  assign n4658 = ~n4654 & ~n4655;
  assign n4659 = ~n4656 & n4658;
  assign n4660 = ~n4657 & n4659;
  assign n4661 = pi29  & n4660;
  assign n4662 = ~pi29  & ~n4660;
  assign n4663 = ~n4661 & ~n4662;
  assign n4664 = n4653 & ~n4663;
  assign n4665 = ~n4651 & ~n4664;
  assign n4666 = ~n4544 & n4553;
  assign n4667 = ~n4554 & ~n4666;
  assign n4668 = ~n4665 & n4667;
  assign n4669 = ~n4554 & ~n4668;
  assign n4670 = n4462 & ~n4464;
  assign n4671 = ~n4465 & ~n4670;
  assign n4672 = ~n4669 & n4671;
  assign n4673 = n4669 & ~n4671;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = ~n802 & n4472;
  assign n4676 = ~n898 & n4070;
  assign n4677 = ~n1006 & n3943;
  assign n4678 = n3944 & n4057;
  assign n4679 = ~n4675 & ~n4676;
  assign n4680 = ~n4677 & n4679;
  assign n4681 = ~n4678 & n4680;
  assign n4682 = pi29  & n4681;
  assign n4683 = ~pi29  & ~n4681;
  assign n4684 = ~n4682 & ~n4683;
  assign n4685 = n4674 & ~n4684;
  assign n4686 = ~n4672 & ~n4685;
  assign n4687 = ~n4471 & n4482;
  assign n4688 = ~n4483 & ~n4687;
  assign n4689 = ~n4686 & n4688;
  assign n4690 = ~n621 & n4515;
  assign n4691 = n4512 & n4513;
  assign n4692 = ~n563 & n4691;
  assign n4693 = n3687 & n4516;
  assign n4694 = ~n4690 & ~n4692;
  assign n4695 = ~n4693 & n4694;
  assign n4696 = ~pi26  & ~n4695;
  assign n4697 = pi26  & n4695;
  assign n4698 = ~n4696 & ~n4697;
  assign n4699 = n4686 & ~n4688;
  assign n4700 = ~n4689 & ~n4699;
  assign n4701 = ~n4698 & n4700;
  assign n4702 = ~n4689 & ~n4701;
  assign n4703 = ~n4535 & ~n4537;
  assign n4704 = ~n4538 & ~n4703;
  assign n4705 = ~n4702 & n4704;
  assign n4706 = ~n898 & n4472;
  assign n4707 = ~n1006 & n4070;
  assign n4708 = ~n1107 & n3943;
  assign n4709 = n3944 & n4041;
  assign n4710 = ~n4706 & ~n4707;
  assign n4711 = ~n4708 & n4710;
  assign n4712 = ~n4709 & n4711;
  assign n4713 = pi29  & n4712;
  assign n4714 = ~pi29  & ~n4712;
  assign n4715 = ~n4713 & ~n4714;
  assign n4716 = n4665 & ~n4667;
  assign n4717 = ~n4668 & ~n4716;
  assign n4718 = ~n4715 & n4717;
  assign n4719 = n4715 & ~n4717;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = n4509 & ~n4512;
  assign n4722 = ~n621 & n4721;
  assign n4723 = ~n729 & n4691;
  assign n4724 = ~n802 & n4515;
  assign n4725 = n3955 & n4516;
  assign n4726 = ~n4722 & ~n4724;
  assign n4727 = ~n4723 & n4726;
  assign n4728 = ~n4725 & n4727;
  assign n4729 = pi26  & n4728;
  assign n4730 = ~pi26  & ~n4728;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = n4720 & ~n4731;
  assign n4733 = ~n4718 & ~n4732;
  assign n4734 = ~n729 & n4515;
  assign n4735 = ~n621 & n4691;
  assign n4736 = ~n563 & n4721;
  assign n4737 = n3921 & n4516;
  assign n4738 = ~n4735 & ~n4736;
  assign n4739 = ~n4734 & n4738;
  assign n4740 = ~n4737 & n4739;
  assign n4741 = pi26  & n4740;
  assign n4742 = ~pi26  & ~n4740;
  assign n4743 = ~n4741 & ~n4742;
  assign n4744 = ~n4733 & ~n4743;
  assign n4745 = ~n4674 & n4684;
  assign n4746 = ~n4685 & ~n4745;
  assign n4747 = n4733 & n4743;
  assign n4748 = ~n4744 & ~n4747;
  assign n4749 = n4746 & n4748;
  assign n4750 = ~n4744 & ~n4749;
  assign n4751 = n4698 & ~n4700;
  assign n4752 = ~n4701 & ~n4751;
  assign n4753 = ~n4750 & n4752;
  assign n4754 = ~n1337 & n3943;
  assign n4755 = ~n1230 & n4070;
  assign n4756 = ~n1107 & n4472;
  assign n4757 = n3944 & n4251;
  assign n4758 = ~n4754 & ~n4755;
  assign n4759 = ~n4756 & n4758;
  assign n4760 = ~n4757 & n4759;
  assign n4761 = ~pi29  & ~n4760;
  assign n4762 = pi29  & n4760;
  assign n4763 = ~n4761 & ~n4762;
  assign n4764 = ~n4637 & n4646;
  assign n4765 = ~n4647 & ~n4764;
  assign n4766 = ~n4763 & n4765;
  assign n4767 = ~n245 & ~n318;
  assign n4768 = ~n365 & ~n594;
  assign n4769 = ~n92 & ~n335;
  assign n4770 = n4768 & n4769;
  assign n4771 = ~n253 & ~n313;
  assign n4772 = n589 & n4771;
  assign n4773 = n1124 & n1397;
  assign n4774 = n1431 & n1786;
  assign n4775 = n2008 & n2391;
  assign n4776 = n2943 & n4767;
  assign n4777 = n4775 & n4776;
  assign n4778 = n4773 & n4774;
  assign n4779 = n4770 & n4772;
  assign n4780 = n4778 & n4779;
  assign n4781 = n1286 & n4777;
  assign n4782 = n4780 & n4781;
  assign n4783 = n2965 & n4782;
  assign n4784 = n757 & n3153;
  assign n4785 = n4783 & n4784;
  assign n4786 = n966 & n4785;
  assign n4787 = ~n246 & ~n319;
  assign n4788 = n943 & n4787;
  assign n4789 = ~n245 & ~n446;
  assign n4790 = ~n210 & ~n212;
  assign n4791 = ~n224 & ~n421;
  assign n4792 = n4790 & n4791;
  assign n4793 = n1911 & n4789;
  assign n4794 = n4792 & n4793;
  assign n4795 = ~n172 & ~n296;
  assign n4796 = ~n405 & ~n578;
  assign n4797 = n237 & n4796;
  assign n4798 = n1965 & n4797;
  assign n4799 = ~n318 & ~n659;
  assign n4800 = n840 & n4799;
  assign n4801 = n923 & n947;
  assign n4802 = n1615 & n2474;
  assign n4803 = n4562 & n4795;
  assign n4804 = n4802 & n4803;
  assign n4805 = n4800 & n4801;
  assign n4806 = n968 & n4788;
  assign n4807 = n4805 & n4806;
  assign n4808 = n2095 & n4804;
  assign n4809 = n4794 & n4798;
  assign n4810 = n4808 & n4809;
  assign n4811 = n4807 & n4810;
  assign n4812 = ~n225 & ~n234;
  assign n4813 = n1355 & n4812;
  assign n4814 = ~n222 & ~n679;
  assign n4815 = n2541 & n4814;
  assign n4816 = ~n192 & ~n200;
  assign n4817 = ~n594 & ~n644;
  assign n4818 = n4816 & n4817;
  assign n4819 = n537 & n1714;
  assign n4820 = n1869 & n2229;
  assign n4821 = n2274 & n2361;
  assign n4822 = n3052 & n4821;
  assign n4823 = n4819 & n4820;
  assign n4824 = n1396 & n4818;
  assign n4825 = n4813 & n4815;
  assign n4826 = n4824 & n4825;
  assign n4827 = n4822 & n4823;
  assign n4828 = n274 & n4827;
  assign n4829 = n4826 & n4828;
  assign n4830 = n4811 & n4829;
  assign n4831 = n1200 & n4830;
  assign n4832 = ~n4786 & ~n4831;
  assign n4833 = n4786 & n4831;
  assign n4834 = ~n4832 & ~n4833;
  assign n4835 = ~pi17  & n4834;
  assign n4836 = ~n4832 & ~n4835;
  assign n4837 = n4358 & ~n4836;
  assign n4838 = ~n4358 & n4836;
  assign n4839 = ~n4837 & ~n4838;
  assign n4840 = n564 & ~n1805;
  assign n4841 = ~n1737 & n3683;
  assign n4842 = ~n1610 & n3896;
  assign n4843 = n3544 & ~n3546;
  assign n4844 = ~n3547 & ~n4843;
  assign n4845 = n566 & n4844;
  assign n4846 = ~n4840 & ~n4841;
  assign n4847 = ~n4842 & n4846;
  assign n4848 = ~n4845 & n4847;
  assign n4849 = n4839 & ~n4848;
  assign n4850 = ~n4837 & ~n4849;
  assign n4851 = ~n4621 & n4630;
  assign n4852 = ~n4631 & ~n4851;
  assign n4853 = ~n4850 & n4852;
  assign n4854 = n4850 & ~n4852;
  assign n4855 = ~n4853 & ~n4854;
  assign n4856 = pi17  & ~n4834;
  assign n4857 = ~n4835 & ~n4856;
  assign n4858 = ~n1805 & n3683;
  assign n4859 = n564 & ~n1893;
  assign n4860 = ~n1737 & n3896;
  assign n4861 = n3540 & ~n3542;
  assign n4862 = ~n3543 & ~n4861;
  assign n4863 = n566 & n4862;
  assign n4864 = ~n4858 & ~n4859;
  assign n4865 = ~n4860 & n4864;
  assign n4866 = ~n4863 & n4865;
  assign n4867 = n4857 & ~n4866;
  assign n4868 = n114 & ~n238;
  assign n4869 = n1267 & n1668;
  assign n4870 = n1868 & n4869;
  assign n4871 = n4868 & n4870;
  assign n4872 = n3178 & n4871;
  assign n4873 = ~n460 & ~n512;
  assign n4874 = n3155 & n4873;
  assign n4875 = ~n199 & ~n218;
  assign n4876 = ~n239 & ~n290;
  assign n4877 = ~n510 & ~n598;
  assign n4878 = ~n659 & ~n681;
  assign n4879 = n4877 & n4878;
  assign n4880 = n4875 & n4876;
  assign n4881 = n540 & n732;
  assign n4882 = n1041 & n1713;
  assign n4883 = n4881 & n4882;
  assign n4884 = n4879 & n4880;
  assign n4885 = n4874 & n4884;
  assign n4886 = n2735 & n4883;
  assign n4887 = n4885 & n4886;
  assign n4888 = ~n177 & ~n200;
  assign n4889 = ~n245 & ~n250;
  assign n4890 = ~n276 & ~n390;
  assign n4891 = ~n424 & ~n463;
  assign n4892 = ~n467 & ~n642;
  assign n4893 = n4891 & n4892;
  assign n4894 = n4889 & n4890;
  assign n4895 = n237 & n4888;
  assign n4896 = n2923 & n3170;
  assign n4897 = n4895 & n4896;
  assign n4898 = n4893 & n4894;
  assign n4899 = n3230 & n4898;
  assign n4900 = n1435 & n4897;
  assign n4901 = n3033 & n4900;
  assign n4902 = n3328 & n4899;
  assign n4903 = n4901 & n4902;
  assign n4904 = n4872 & n4887;
  assign n4905 = n4903 & n4904;
  assign n4906 = n3728 & n4905;
  assign n4907 = n4786 & ~n4906;
  assign n4908 = ~n340 & ~n495;
  assign n4909 = n1558 & n4908;
  assign n4910 = n1873 & n4909;
  assign n4911 = ~n334 & ~n676;
  assign n4912 = ~n141 & ~n513;
  assign n4913 = n1397 & n4912;
  assign n4914 = n3729 & n4911;
  assign n4915 = n4913 & n4914;
  assign n4916 = ~n193 & ~n212;
  assign n4917 = ~n243 & ~n327;
  assign n4918 = ~n588 & n4917;
  assign n4919 = n920 & n4916;
  assign n4920 = n1714 & n2150;
  assign n4921 = n3428 & n4920;
  assign n4922 = n4918 & n4919;
  assign n4923 = n2662 & n3324;
  assign n4924 = n4922 & n4923;
  assign n4925 = n4910 & n4921;
  assign n4926 = n4915 & n4925;
  assign n4927 = n4924 & n4926;
  assign n4928 = n4872 & n4927;
  assign n4929 = ~n91 & ~n401;
  assign n4930 = ~n554 & n4929;
  assign n4931 = ~n183 & ~n496;
  assign n4932 = ~n242 & ~n290;
  assign n4933 = ~n247 & ~n289;
  assign n4934 = ~n103 & n4933;
  assign n4935 = ~n239 & ~n388;
  assign n4936 = n2048 & n4935;
  assign n4937 = ~n168 & ~n321;
  assign n4938 = ~n323 & ~n384;
  assign n4939 = ~n473 & ~n659;
  assign n4940 = ~n687 & n4939;
  assign n4941 = n4937 & n4938;
  assign n4942 = n408 & n4941;
  assign n4943 = n1834 & n4940;
  assign n4944 = n3715 & n4934;
  assign n4945 = n4936 & n4944;
  assign n4946 = n4942 & n4943;
  assign n4947 = n1213 & n3232;
  assign n4948 = n4946 & n4947;
  assign n4949 = n4945 & n4948;
  assign n4950 = ~n378 & ~n569;
  assign n4951 = ~n680 & n4950;
  assign n4952 = ~n179 & ~n279;
  assign n4953 = ~n690 & n4952;
  assign n4954 = n268 & n3052;
  assign n4955 = n4953 & n4954;
  assign n4956 = n4951 & n4955;
  assign n4957 = ~n585 & n733;
  assign n4958 = ~n200 & ~n318;
  assign n4959 = ~n338 & ~n355;
  assign n4960 = ~n364 & ~n375;
  assign n4961 = ~n510 & ~n543;
  assign n4962 = n4960 & n4961;
  assign n4963 = n4958 & n4959;
  assign n4964 = n121 & n1173;
  assign n4965 = n2358 & n4964;
  assign n4966 = n4962 & n4963;
  assign n4967 = n4957 & n4966;
  assign n4968 = n4965 & n4967;
  assign n4969 = ~n196 & ~n269;
  assign n4970 = ~n446 & ~n571;
  assign n4971 = n4969 & n4970;
  assign n4972 = n732 & n923;
  assign n4973 = n927 & n4931;
  assign n4974 = n4932 & n4973;
  assign n4975 = n4971 & n4972;
  assign n4976 = n2884 & n4930;
  assign n4977 = n4975 & n4976;
  assign n4978 = n4326 & n4974;
  assign n4979 = n4977 & n4978;
  assign n4980 = n4956 & n4979;
  assign n4981 = n4968 & n4980;
  assign n4982 = n4949 & n4981;
  assign n4983 = n4928 & n4982;
  assign n4984 = ~n103 & ~n270;
  assign n4985 = n169 & ~n200;
  assign n4986 = ~n584 & ~n595;
  assign n4987 = ~n199 & ~n215;
  assign n4988 = ~n267 & ~n300;
  assign n4989 = ~n318 & ~n494;
  assign n4990 = ~n690 & n4989;
  assign n4991 = n4987 & n4988;
  assign n4992 = n1650 & n2063;
  assign n4993 = n4984 & n4986;
  assign n4994 = n4992 & n4993;
  assign n4995 = n4990 & n4991;
  assign n4996 = n1584 & n4985;
  assign n4997 = n4995 & n4996;
  assign n4998 = n3008 & n4994;
  assign n4999 = n4561 & n4998;
  assign n5000 = n4997 & n4999;
  assign n5001 = n1710 & n2086;
  assign n5002 = ~n210 & ~n360;
  assign n5003 = ~n265 & ~n312;
  assign n5004 = ~n700 & n5003;
  assign n5005 = n93 & n1785;
  assign n5006 = n2958 & n3381;
  assign n5007 = n3870 & n5006;
  assign n5008 = n5004 & n5005;
  assign n5009 = n4813 & n5008;
  assign n5010 = n5007 & n5009;
  assign n5011 = ~n192 & ~n240;
  assign n5012 = ~n327 & ~n472;
  assign n5013 = ~n509 & ~n642;
  assign n5014 = n5012 & n5013;
  assign n5015 = n1472 & n5011;
  assign n5016 = n2112 & n2300;
  assign n5017 = n5002 & n5016;
  assign n5018 = n5014 & n5015;
  assign n5019 = n4874 & n5018;
  assign n5020 = n5017 & n5019;
  assign n5021 = n911 & n5020;
  assign n5022 = n5010 & n5021;
  assign n5023 = ~n492 & ~n650;
  assign n5024 = ~n324 & ~n587;
  assign n5025 = n1744 & n5024;
  assign n5026 = n1869 & n4265;
  assign n5027 = n5023 & n5026;
  assign n5028 = n1964 & n5025;
  assign n5029 = n3026 & n5028;
  assign n5030 = n5027 & n5029;
  assign n5031 = ~n134 & ~n406;
  assign n5032 = ~n597 & n5031;
  assign n5033 = n1559 & n5032;
  assign n5034 = n2479 & n5033;
  assign n5035 = ~n131 & ~n644;
  assign n5036 = ~n670 & n5035;
  assign n5037 = n223 & n423;
  assign n5038 = n781 & n1070;
  assign n5039 = n1354 & n5038;
  assign n5040 = n5036 & n5037;
  assign n5041 = n970 & n1836;
  assign n5042 = n5001 & n5041;
  assign n5043 = n5039 & n5040;
  assign n5044 = n5042 & n5043;
  assign n5045 = n5034 & n5044;
  assign n5046 = n5030 & n5045;
  assign n5047 = n5000 & n5046;
  assign n5048 = n5022 & n5047;
  assign n5049 = ~n4983 & ~n5048;
  assign n5050 = n4983 & n5048;
  assign n5051 = ~n5049 & ~n5050;
  assign n5052 = ~pi14  & n5051;
  assign n5053 = ~n5049 & ~n5052;
  assign n5054 = n4906 & ~n5053;
  assign n5055 = ~n4906 & n5053;
  assign n5056 = ~n5054 & ~n5055;
  assign n5057 = n564 & ~n2045;
  assign n5058 = ~n1997 & n3683;
  assign n5059 = ~n1893 & n3896;
  assign n5060 = n3532 & ~n3534;
  assign n5061 = ~n3535 & ~n5060;
  assign n5062 = n566 & n5061;
  assign n5063 = ~n5057 & ~n5058;
  assign n5064 = ~n5059 & n5063;
  assign n5065 = ~n5062 & n5064;
  assign n5066 = n5056 & ~n5065;
  assign n5067 = ~n5054 & ~n5066;
  assign n5068 = ~n4786 & n4906;
  assign n5069 = ~n4907 & ~n5068;
  assign n5070 = ~n5067 & n5069;
  assign n5071 = ~n4907 & ~n5070;
  assign n5072 = ~n4857 & n4866;
  assign n5073 = ~n4867 & ~n5072;
  assign n5074 = ~n5071 & n5073;
  assign n5075 = ~n4867 & ~n5074;
  assign n5076 = ~n4839 & n4848;
  assign n5077 = ~n4849 & ~n5076;
  assign n5078 = ~n5075 & n5077;
  assign n5079 = n5075 & ~n5077;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = ~n1532 & n3943;
  assign n5082 = ~n1425 & n4070;
  assign n5083 = ~n1337 & n4472;
  assign n5084 = n3944 & n4452;
  assign n5085 = ~n5081 & ~n5082;
  assign n5086 = ~n5083 & n5085;
  assign n5087 = ~n5084 & n5086;
  assign n5088 = pi29  & n5087;
  assign n5089 = ~pi29  & ~n5087;
  assign n5090 = ~n5088 & ~n5089;
  assign n5091 = n5080 & ~n5090;
  assign n5092 = ~n5078 & ~n5091;
  assign n5093 = n4855 & ~n5092;
  assign n5094 = ~n4853 & ~n5093;
  assign n5095 = n4763 & ~n4765;
  assign n5096 = ~n4766 & ~n5095;
  assign n5097 = ~n5094 & n5096;
  assign n5098 = ~n4766 & ~n5097;
  assign n5099 = ~n4653 & n4663;
  assign n5100 = ~n4664 & ~n5099;
  assign n5101 = ~n5098 & n5100;
  assign n5102 = ~n729 & n4721;
  assign n5103 = ~n802 & n4691;
  assign n5104 = ~n898 & n4515;
  assign n5105 = n3901 & n4516;
  assign n5106 = ~n5103 & ~n5104;
  assign n5107 = ~n5102 & n5106;
  assign n5108 = ~n5105 & n5107;
  assign n5109 = ~pi26  & ~n5108;
  assign n5110 = pi26  & n5108;
  assign n5111 = ~n5109 & ~n5110;
  assign n5112 = n5098 & ~n5100;
  assign n5113 = ~n5101 & ~n5112;
  assign n5114 = ~n5111 & n5113;
  assign n5115 = ~n5101 & ~n5114;
  assign n5116 = n78 & ~n3593;
  assign n5117 = ~pi21  & ~pi22 ;
  assign n5118 = pi21  & pi22 ;
  assign n5119 = ~n5117 & ~n5118;
  assign n5120 = ~n74 & n77;
  assign n5121 = ~n5119 & n5120;
  assign n5122 = ~n5116 & ~n5121;
  assign n5123 = ~n563 & ~n5122;
  assign n5124 = pi23  & ~n5123;
  assign n5125 = ~pi23  & n5123;
  assign n5126 = ~n5124 & ~n5125;
  assign n5127 = ~n5115 & ~n5126;
  assign n5128 = n5115 & n5126;
  assign n5129 = ~n5127 & ~n5128;
  assign n5130 = ~n4720 & n4731;
  assign n5131 = ~n4732 & ~n5130;
  assign n5132 = n5129 & n5131;
  assign n5133 = ~n5127 & ~n5132;
  assign n5134 = ~n4746 & ~n4748;
  assign n5135 = ~n4749 & ~n5134;
  assign n5136 = ~n5133 & n5135;
  assign n5137 = n5094 & ~n5096;
  assign n5138 = ~n5097 & ~n5137;
  assign n5139 = ~n802 & n4721;
  assign n5140 = ~n898 & n4691;
  assign n5141 = ~n1006 & n4515;
  assign n5142 = n4057 & n4516;
  assign n5143 = ~n5139 & ~n5140;
  assign n5144 = ~n5141 & n5143;
  assign n5145 = ~n5142 & n5144;
  assign n5146 = pi26  & n5145;
  assign n5147 = ~pi26  & ~n5145;
  assign n5148 = ~n5146 & ~n5147;
  assign n5149 = n5138 & ~n5148;
  assign n5150 = ~n4855 & n5092;
  assign n5151 = ~n5093 & ~n5150;
  assign n5152 = ~n1425 & n3943;
  assign n5153 = ~n1337 & n4070;
  assign n5154 = ~n1230 & n4472;
  assign n5155 = n3944 & n4549;
  assign n5156 = ~n5152 & ~n5153;
  assign n5157 = ~n5154 & n5156;
  assign n5158 = ~n5155 & n5157;
  assign n5159 = pi29  & n5158;
  assign n5160 = ~pi29  & ~n5158;
  assign n5161 = ~n5159 & ~n5160;
  assign n5162 = n5151 & ~n5161;
  assign n5163 = ~n898 & n4721;
  assign n5164 = ~n1006 & n4691;
  assign n5165 = ~n1107 & n4515;
  assign n5166 = n4041 & n4516;
  assign n5167 = ~n5163 & ~n5164;
  assign n5168 = ~n5165 & n5167;
  assign n5169 = ~n5166 & n5168;
  assign n5170 = pi26  & n5169;
  assign n5171 = ~pi26  & ~n5169;
  assign n5172 = ~n5170 & ~n5171;
  assign n5173 = ~n5151 & n5161;
  assign n5174 = ~n5162 & ~n5173;
  assign n5175 = ~n5172 & n5174;
  assign n5176 = ~n5162 & ~n5175;
  assign n5177 = ~n5138 & n5148;
  assign n5178 = ~n5149 & ~n5177;
  assign n5179 = ~n5176 & n5178;
  assign n5180 = ~n5149 & ~n5179;
  assign n5181 = n5111 & ~n5113;
  assign n5182 = ~n5114 & ~n5181;
  assign n5183 = ~n5180 & n5182;
  assign n5184 = ~n621 & n5121;
  assign n5185 = ~n74 & n5119;
  assign n5186 = ~n563 & n5185;
  assign n5187 = n78 & n3687;
  assign n5188 = ~n5184 & ~n5186;
  assign n5189 = ~n5187 & n5188;
  assign n5190 = ~pi23  & ~n5189;
  assign n5191 = pi23  & n5189;
  assign n5192 = ~n5190 & ~n5191;
  assign n5193 = n5180 & ~n5182;
  assign n5194 = ~n5183 & ~n5193;
  assign n5195 = ~n5192 & n5194;
  assign n5196 = ~n5183 & ~n5195;
  assign n5197 = ~n5129 & ~n5131;
  assign n5198 = ~n5132 & ~n5197;
  assign n5199 = ~n5196 & n5198;
  assign n5200 = n5196 & ~n5198;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = n5172 & ~n5174;
  assign n5203 = ~n5175 & ~n5202;
  assign n5204 = ~n5080 & n5090;
  assign n5205 = ~n5091 & ~n5204;
  assign n5206 = n5067 & ~n5069;
  assign n5207 = ~n5070 & ~n5206;
  assign n5208 = ~n1893 & n3683;
  assign n5209 = n564 & ~n1997;
  assign n5210 = ~n1805 & n3896;
  assign n5211 = n3536 & ~n3538;
  assign n5212 = ~n3539 & ~n5211;
  assign n5213 = n566 & n5212;
  assign n5214 = ~n5208 & ~n5209;
  assign n5215 = ~n5210 & n5214;
  assign n5216 = ~n5213 & n5215;
  assign n5217 = n5207 & ~n5216;
  assign n5218 = ~n1737 & n3943;
  assign n5219 = ~n1610 & n4070;
  assign n5220 = ~n1532 & n4472;
  assign n5221 = n3944 & n4626;
  assign n5222 = ~n5218 & ~n5219;
  assign n5223 = ~n5220 & n5222;
  assign n5224 = ~n5221 & n5223;
  assign n5225 = ~pi29  & ~n5224;
  assign n5226 = pi29  & n5224;
  assign n5227 = ~n5225 & ~n5226;
  assign n5228 = ~n5207 & n5216;
  assign n5229 = ~n5217 & ~n5228;
  assign n5230 = ~n5227 & n5229;
  assign n5231 = ~n5217 & ~n5230;
  assign n5232 = n5071 & ~n5073;
  assign n5233 = ~n5074 & ~n5232;
  assign n5234 = n5231 & ~n5233;
  assign n5235 = ~n1610 & n3943;
  assign n5236 = ~n1532 & n4070;
  assign n5237 = ~n1425 & n4472;
  assign n5238 = n3944 & n4642;
  assign n5239 = ~n5235 & ~n5236;
  assign n5240 = ~n5237 & n5239;
  assign n5241 = ~n5238 & n5240;
  assign n5242 = pi29  & n5241;
  assign n5243 = ~pi29  & ~n5241;
  assign n5244 = ~n5242 & ~n5243;
  assign n5245 = ~n5231 & n5233;
  assign n5246 = ~n5234 & ~n5245;
  assign n5247 = n5244 & n5246;
  assign n5248 = ~n5234 & ~n5247;
  assign n5249 = ~n5205 & ~n5248;
  assign n5250 = n5205 & n5248;
  assign n5251 = ~n5249 & ~n5250;
  assign n5252 = ~n1107 & n4691;
  assign n5253 = ~n1006 & n4721;
  assign n5254 = ~n1230 & n4515;
  assign n5255 = n4233 & n4516;
  assign n5256 = ~n5252 & ~n5253;
  assign n5257 = ~n5254 & n5256;
  assign n5258 = ~n5255 & n5257;
  assign n5259 = pi26  & n5258;
  assign n5260 = ~pi26  & ~n5258;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = n5251 & n5261;
  assign n5263 = ~n5249 & ~n5262;
  assign n5264 = n5203 & n5263;
  assign n5265 = ~n5203 & ~n5263;
  assign n5266 = ~n5264 & ~n5265;
  assign n5267 = n74 & ~n77;
  assign n5268 = ~n621 & n5267;
  assign n5269 = ~n729 & n5185;
  assign n5270 = ~n802 & n5121;
  assign n5271 = n78 & n3955;
  assign n5272 = ~n5268 & ~n5270;
  assign n5273 = ~n5269 & n5272;
  assign n5274 = ~n5271 & n5273;
  assign n5275 = pi23  & n5274;
  assign n5276 = ~pi23  & ~n5274;
  assign n5277 = ~n5275 & ~n5276;
  assign n5278 = n5266 & ~n5277;
  assign n5279 = ~n5264 & ~n5278;
  assign n5280 = ~n729 & n5121;
  assign n5281 = ~n621 & n5185;
  assign n5282 = ~n563 & n5267;
  assign n5283 = n78 & n3921;
  assign n5284 = ~n5281 & ~n5282;
  assign n5285 = ~n5280 & n5284;
  assign n5286 = ~n5283 & n5285;
  assign n5287 = pi23  & n5286;
  assign n5288 = ~pi23  & ~n5286;
  assign n5289 = ~n5287 & ~n5288;
  assign n5290 = ~n5279 & ~n5289;
  assign n5291 = n5279 & n5289;
  assign n5292 = ~n5290 & ~n5291;
  assign n5293 = n5176 & ~n5178;
  assign n5294 = ~n5179 & ~n5293;
  assign n5295 = n5292 & n5294;
  assign n5296 = ~n5290 & ~n5295;
  assign n5297 = n5192 & ~n5194;
  assign n5298 = ~n5195 & ~n5297;
  assign n5299 = ~n5296 & n5298;
  assign n5300 = ~pi19  & ~pi20 ;
  assign n5301 = pi19  & pi20 ;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = ~pi17  & ~pi18 ;
  assign n5304 = pi17  & pi18 ;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = n5302 & n5305;
  assign n5307 = ~n3593 & n5306;
  assign n5308 = ~pi18  & ~pi19 ;
  assign n5309 = pi18  & pi19 ;
  assign n5310 = ~n5308 & ~n5309;
  assign n5311 = n5302 & ~n5305;
  assign n5312 = ~n5310 & n5311;
  assign n5313 = ~n5307 & ~n5312;
  assign n5314 = ~n563 & ~n5313;
  assign n5315 = pi20  & ~n5314;
  assign n5316 = ~pi20  & n5314;
  assign n5317 = ~n5315 & ~n5316;
  assign n5318 = ~n5251 & ~n5261;
  assign n5319 = ~n5262 & ~n5318;
  assign n5320 = ~n5244 & ~n5246;
  assign n5321 = ~n5247 & ~n5320;
  assign n5322 = ~n1337 & n4515;
  assign n5323 = ~n1230 & n4691;
  assign n5324 = ~n1107 & n4721;
  assign n5325 = n4251 & n4516;
  assign n5326 = ~n5322 & ~n5323;
  assign n5327 = ~n5324 & n5326;
  assign n5328 = ~n5325 & n5327;
  assign n5329 = pi26  & n5328;
  assign n5330 = ~pi26  & ~n5328;
  assign n5331 = ~n5329 & ~n5330;
  assign n5332 = ~n5321 & ~n5331;
  assign n5333 = ~n225 & ~n355;
  assign n5334 = ~n568 & ~n665;
  assign n5335 = n5333 & n5334;
  assign n5336 = n1612 & n4266;
  assign n5337 = n5335 & n5336;
  assign n5338 = ~n254 & ~n270;
  assign n5339 = ~n168 & ~n467;
  assign n5340 = n1171 & n5339;
  assign n5341 = ~n238 & n278;
  assign n5342 = n1382 & n5341;
  assign n5343 = ~n265 & ~n539;
  assign n5344 = ~n180 & ~n234;
  assign n5345 = n403 & n5344;
  assign n5346 = n436 & n904;
  assign n5347 = n943 & n1783;
  assign n5348 = n2566 & n4093;
  assign n5349 = n4767 & n5343;
  assign n5350 = n5348 & n5349;
  assign n5351 = n5346 & n5347;
  assign n5352 = n5340 & n5345;
  assign n5353 = n5351 & n5352;
  assign n5354 = n5342 & n5350;
  assign n5355 = n5353 & n5354;
  assign n5356 = n1353 & n5355;
  assign n5357 = ~n196 & ~n469;
  assign n5358 = ~n687 & n5357;
  assign n5359 = n3105 & n5358;
  assign n5360 = ~n92 & ~n209;
  assign n5361 = ~n343 & ~n522;
  assign n5362 = n5360 & n5361;
  assign n5363 = n252 & n1112;
  assign n5364 = n3282 & n5363;
  assign n5365 = n3342 & n5362;
  assign n5366 = n5364 & n5365;
  assign n5367 = n5359 & n5366;
  assign n5368 = ~n342 & ~n512;
  assign n5369 = ~n246 & ~n543;
  assign n5370 = ~n242 & n497;
  assign n5371 = n3870 & n5370;
  assign n5372 = ~n167 & ~n689;
  assign n5373 = ~n509 & ~n553;
  assign n5374 = ~n583 & ~n648;
  assign n5375 = n5373 & n5374;
  assign n5376 = n677 & n1756;
  assign n5377 = n3763 & n5369;
  assign n5378 = n5372 & n5377;
  assign n5379 = n5375 & n5376;
  assign n5380 = n1265 & n3828;
  assign n5381 = n4325 & n5380;
  assign n5382 = n5378 & n5379;
  assign n5383 = n5371 & n5382;
  assign n5384 = n3979 & n5381;
  assign n5385 = n5383 & n5384;
  assign n5386 = ~n139 & ~n147;
  assign n5387 = ~n310 & ~n427;
  assign n5388 = ~n472 & n5387;
  assign n5389 = n1113 & n5386;
  assign n5390 = n1469 & n3154;
  assign n5391 = n5338 & n5368;
  assign n5392 = n5390 & n5391;
  assign n5393 = n5388 & n5389;
  assign n5394 = n1010 & n5393;
  assign n5395 = n2708 & n5392;
  assign n5396 = n5337 & n5395;
  assign n5397 = n5394 & n5396;
  assign n5398 = n5367 & n5397;
  assign n5399 = n5356 & n5385;
  assign n5400 = n5398 & n5399;
  assign n5401 = n4983 & ~n5400;
  assign n5402 = ~n4983 & n5400;
  assign n5403 = ~n5401 & ~n5402;
  assign n5404 = ~n2165 & n3683;
  assign n5405 = n564 & ~n2265;
  assign n5406 = ~n2045 & n3896;
  assign n5407 = n3524 & ~n3526;
  assign n5408 = ~n3527 & ~n5407;
  assign n5409 = n566 & n5408;
  assign n5410 = ~n5405 & ~n5406;
  assign n5411 = ~n5404 & n5410;
  assign n5412 = ~n5409 & n5411;
  assign n5413 = n5403 & ~n5412;
  assign n5414 = ~n5401 & ~n5413;
  assign n5415 = pi14  & ~n5051;
  assign n5416 = ~n5052 & ~n5415;
  assign n5417 = ~n5414 & n5416;
  assign n5418 = n5414 & ~n5416;
  assign n5419 = ~n5417 & ~n5418;
  assign n5420 = n564 & ~n2165;
  assign n5421 = ~n2045 & n3683;
  assign n5422 = ~n1997 & n3896;
  assign n5423 = n3528 & ~n3530;
  assign n5424 = ~n3531 & ~n5423;
  assign n5425 = n566 & n5424;
  assign n5426 = ~n5421 & ~n5422;
  assign n5427 = ~n5420 & n5426;
  assign n5428 = ~n5425 & n5427;
  assign n5429 = n5419 & ~n5428;
  assign n5430 = ~n5417 & ~n5429;
  assign n5431 = ~n5056 & n5065;
  assign n5432 = ~n5066 & ~n5431;
  assign n5433 = ~n5430 & n5432;
  assign n5434 = n5430 & ~n5432;
  assign n5435 = ~n5433 & ~n5434;
  assign n5436 = ~n1805 & n3943;
  assign n5437 = ~n1737 & n4070;
  assign n5438 = ~n1610 & n4472;
  assign n5439 = n3944 & n4844;
  assign n5440 = ~n5436 & ~n5437;
  assign n5441 = ~n5438 & n5440;
  assign n5442 = ~n5439 & n5441;
  assign n5443 = pi29  & n5442;
  assign n5444 = ~pi29  & ~n5442;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = n5435 & ~n5445;
  assign n5447 = ~n5433 & ~n5446;
  assign n5448 = n5227 & ~n5229;
  assign n5449 = ~n5230 & ~n5448;
  assign n5450 = ~n5447 & n5449;
  assign n5451 = n5447 & ~n5449;
  assign n5452 = ~n5450 & ~n5451;
  assign n5453 = ~n1425 & n4515;
  assign n5454 = ~n1337 & n4691;
  assign n5455 = ~n1230 & n4721;
  assign n5456 = n4516 & n4549;
  assign n5457 = ~n5453 & ~n5454;
  assign n5458 = ~n5455 & n5457;
  assign n5459 = ~n5456 & n5458;
  assign n5460 = pi26  & n5459;
  assign n5461 = ~pi26  & ~n5459;
  assign n5462 = ~n5460 & ~n5461;
  assign n5463 = n5452 & ~n5462;
  assign n5464 = ~n5450 & ~n5463;
  assign n5465 = n5321 & n5331;
  assign n5466 = ~n5332 & ~n5465;
  assign n5467 = ~n5464 & n5466;
  assign n5468 = ~n5332 & ~n5467;
  assign n5469 = n5319 & n5468;
  assign n5470 = ~n5319 & ~n5468;
  assign n5471 = ~n5469 & ~n5470;
  assign n5472 = ~n729 & n5267;
  assign n5473 = ~n802 & n5185;
  assign n5474 = ~n898 & n5121;
  assign n5475 = n78 & n3901;
  assign n5476 = ~n5473 & ~n5474;
  assign n5477 = ~n5472 & n5476;
  assign n5478 = ~n5475 & n5477;
  assign n5479 = pi23  & n5478;
  assign n5480 = ~pi23  & ~n5478;
  assign n5481 = ~n5479 & ~n5480;
  assign n5482 = n5471 & n5481;
  assign n5483 = ~n5469 & ~n5482;
  assign n5484 = ~n5317 & n5483;
  assign n5485 = n5317 & ~n5483;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = ~n5266 & n5277;
  assign n5488 = ~n5278 & ~n5487;
  assign n5489 = n5486 & n5488;
  assign n5490 = ~n5484 & ~n5489;
  assign n5491 = ~n5292 & ~n5294;
  assign n5492 = ~n5295 & ~n5491;
  assign n5493 = ~n5490 & n5492;
  assign n5494 = n5490 & ~n5492;
  assign n5495 = ~n5493 & ~n5494;
  assign n5496 = ~n5471 & ~n5481;
  assign n5497 = ~n5482 & ~n5496;
  assign n5498 = ~n802 & n5267;
  assign n5499 = ~n898 & n5185;
  assign n5500 = ~n1006 & n5121;
  assign n5501 = n78 & n4057;
  assign n5502 = ~n5498 & ~n5499;
  assign n5503 = ~n5500 & n5502;
  assign n5504 = ~n5501 & n5503;
  assign n5505 = ~pi23  & ~n5504;
  assign n5506 = pi23  & n5504;
  assign n5507 = ~n5505 & ~n5506;
  assign n5508 = n5464 & ~n5466;
  assign n5509 = ~n5467 & ~n5508;
  assign n5510 = ~n5507 & n5509;
  assign n5511 = ~n5452 & n5462;
  assign n5512 = ~n5463 & ~n5511;
  assign n5513 = ~n1893 & n3943;
  assign n5514 = ~n1805 & n4070;
  assign n5515 = ~n1737 & n4472;
  assign n5516 = n3944 & n4862;
  assign n5517 = ~n5513 & ~n5514;
  assign n5518 = ~n5515 & n5517;
  assign n5519 = ~n5516 & n5518;
  assign n5520 = ~pi29  & ~n5519;
  assign n5521 = pi29  & n5519;
  assign n5522 = ~n5520 & ~n5521;
  assign n5523 = ~n5419 & n5428;
  assign n5524 = ~n5429 & ~n5523;
  assign n5525 = ~n5522 & n5524;
  assign n5526 = ~n247 & ~n319;
  assign n5527 = ~n173 & ~n236;
  assign n5528 = ~n385 & n5527;
  assign n5529 = ~n448 & ~n459;
  assign n5530 = n1350 & n2472;
  assign n5531 = n2738 & n5529;
  assign n5532 = n5530 & n5531;
  assign n5533 = ~n343 & ~n355;
  assign n5534 = ~n570 & ~n673;
  assign n5535 = n1094 & n5534;
  assign n5536 = n1614 & n5533;
  assign n5537 = n4156 & n5526;
  assign n5538 = n5536 & n5537;
  assign n5539 = n2064 & n5535;
  assign n5540 = n2560 & n5528;
  assign n5541 = n5539 & n5540;
  assign n5542 = n5532 & n5538;
  assign n5543 = n5541 & n5542;
  assign n5544 = ~n283 & ~n390;
  assign n5545 = ~n470 & n5544;
  assign n5546 = ~n289 & ~n310;
  assign n5547 = ~n649 & n5546;
  assign n5548 = n600 & ~n640;
  assign n5549 = n3071 & n5548;
  assign n5550 = ~n225 & ~n282;
  assign n5551 = n737 & n5023;
  assign n5552 = ~n202 & ~n219;
  assign n5553 = ~n234 & ~n316;
  assign n5554 = ~n460 & n5553;
  assign n5555 = n361 & n5552;
  assign n5556 = n921 & n3203;
  assign n5557 = n5550 & n5556;
  assign n5558 = n5554 & n5555;
  assign n5559 = n2151 & n5551;
  assign n5560 = n5558 & n5559;
  assign n5561 = n5557 & n5560;
  assign n5562 = ~n192 & ~n578;
  assign n5563 = n1615 & n5562;
  assign n5564 = n3628 & n4405;
  assign n5565 = n5563 & n5564;
  assign n5566 = n5545 & n5547;
  assign n5567 = n5565 & n5566;
  assign n5568 = n5549 & n5567;
  assign n5569 = n2372 & n4956;
  assign n5570 = n5568 & n5569;
  assign n5571 = n5543 & n5561;
  assign n5572 = n5570 & n5571;
  assign n5573 = n1262 & n5572;
  assign n5574 = ~n224 & ~n448;
  assign n5575 = ~n310 & ~n578;
  assign n5576 = ~n662 & ~n690;
  assign n5577 = n5575 & n5576;
  assign n5578 = ~n208 & ~n246;
  assign n5579 = ~n340 & n5578;
  assign n5580 = n3266 & n4266;
  assign n5581 = n5579 & n5580;
  assign n5582 = n3139 & n5577;
  assign n5583 = n5581 & n5582;
  assign n5584 = ~n319 & ~n666;
  assign n5585 = ~n683 & n5584;
  assign n5586 = ~n222 & ~n265;
  assign n5587 = ~n665 & ~n670;
  assign n5588 = n5586 & n5587;
  assign n5589 = n596 & n1869;
  assign n5590 = n2093 & n2475;
  assign n5591 = n2480 & n3658;
  assign n5592 = n3843 & n5574;
  assign n5593 = n5591 & n5592;
  assign n5594 = n5589 & n5590;
  assign n5595 = n5585 & n5588;
  assign n5596 = n5594 & n5595;
  assign n5597 = n1567 & n5593;
  assign n5598 = n5596 & n5597;
  assign n5599 = n5583 & n5598;
  assign n5600 = ~n91 & ~n98;
  assign n5601 = ~n212 & ~n299;
  assign n5602 = ~n495 & ~n539;
  assign n5603 = ~n588 & n5602;
  assign n5604 = n5600 & n5601;
  assign n5605 = n211 & n857;
  assign n5606 = n969 & n1121;
  assign n5607 = n1301 & n1614;
  assign n5608 = n1651 & n1808;
  assign n5609 = n5607 & n5608;
  assign n5610 = n5605 & n5606;
  assign n5611 = n5603 & n5604;
  assign n5612 = n1946 & n3611;
  assign n5613 = n5611 & n5612;
  assign n5614 = n5609 & n5610;
  assign n5615 = n5613 & n5614;
  assign n5616 = n4311 & n5615;
  assign n5617 = n4103 & n5561;
  assign n5618 = n5616 & n5617;
  assign n5619 = n5599 & n5618;
  assign n5620 = ~n5573 & ~n5619;
  assign n5621 = n5573 & n5619;
  assign n5622 = ~n5620 & ~n5621;
  assign n5623 = ~pi11  & n5622;
  assign n5624 = ~n5620 & ~n5623;
  assign n5625 = n4983 & ~n5624;
  assign n5626 = ~n4983 & n5624;
  assign n5627 = ~n5625 & ~n5626;
  assign n5628 = n564 & ~n2356;
  assign n5629 = ~n2265 & n3683;
  assign n5630 = ~n2165 & n3896;
  assign n5631 = n3520 & ~n3522;
  assign n5632 = ~n3523 & ~n5631;
  assign n5633 = n566 & n5632;
  assign n5634 = ~n5628 & ~n5629;
  assign n5635 = ~n5630 & n5634;
  assign n5636 = ~n5633 & n5635;
  assign n5637 = n5627 & ~n5636;
  assign n5638 = ~n5625 & ~n5637;
  assign n5639 = ~n5403 & n5412;
  assign n5640 = ~n5413 & ~n5639;
  assign n5641 = ~n5638 & n5640;
  assign n5642 = n5638 & ~n5640;
  assign n5643 = ~n5641 & ~n5642;
  assign n5644 = pi11  & ~n5622;
  assign n5645 = ~n5623 & ~n5644;
  assign n5646 = ~n2356 & n3683;
  assign n5647 = n564 & ~n2442;
  assign n5648 = ~n2265 & n3896;
  assign n5649 = n3516 & ~n3518;
  assign n5650 = ~n3519 & ~n5649;
  assign n5651 = n566 & n5650;
  assign n5652 = ~n5647 & ~n5648;
  assign n5653 = ~n5646 & n5652;
  assign n5654 = ~n5651 & n5653;
  assign n5655 = n5645 & ~n5654;
  assign n5656 = ~n180 & ~n679;
  assign n5657 = n2063 & n5656;
  assign n5658 = ~n141 & ~n577;
  assign n5659 = n2272 & n5658;
  assign n5660 = ~n168 & ~n300;
  assign n5661 = ~n425 & ~n681;
  assign n5662 = n2008 & n5661;
  assign n5663 = n5660 & n5662;
  assign n5664 = ~n236 & ~n287;
  assign n5665 = ~n307 & ~n343;
  assign n5666 = ~n459 & ~n492;
  assign n5667 = ~n640 & n5666;
  assign n5668 = n5664 & n5665;
  assign n5669 = n2706 & n3171;
  assign n5670 = n5668 & n5669;
  assign n5671 = n1743 & n5667;
  assign n5672 = n5657 & n5659;
  assign n5673 = n5671 & n5672;
  assign n5674 = n5663 & n5670;
  assign n5675 = n5673 & n5674;
  assign n5676 = n4116 & n5675;
  assign n5677 = n2404 & n5676;
  assign n5678 = n2389 & n5677;
  assign n5679 = n1707 & n5678;
  assign n5680 = n5573 & ~n5679;
  assign n5681 = ~n574 & ~n675;
  assign n5682 = ~n356 & ~n580;
  assign n5683 = ~n323 & ~n448;
  assign n5684 = ~n587 & n5683;
  assign n5685 = n284 & n2455;
  assign n5686 = n5682 & n5685;
  assign n5687 = n5684 & n5686;
  assign n5688 = ~n235 & ~n311;
  assign n5689 = ~n354 & ~n407;
  assign n5690 = ~n427 & ~n538;
  assign n5691 = ~n651 & ~n662;
  assign n5692 = ~n676 & n5691;
  assign n5693 = n5689 & n5690;
  assign n5694 = n4161 & n5688;
  assign n5695 = n5693 & n5694;
  assign n5696 = n5692 & n5695;
  assign n5697 = ~n109 & ~n165;
  assign n5698 = ~n200 & ~n215;
  assign n5699 = ~n467 & ~n492;
  assign n5700 = n5698 & n5699;
  assign n5701 = n5697 & n5700;
  assign n5702 = n2908 & n5701;
  assign n5703 = ~n149 & ~n172;
  assign n5704 = ~n207 & ~n362;
  assign n5705 = ~n402 & ~n445;
  assign n5706 = ~n521 & ~n599;
  assign n5707 = ~n701 & n5706;
  assign n5708 = n5704 & n5705;
  assign n5709 = n328 & n5703;
  assign n5710 = n1114 & n5709;
  assign n5711 = n5707 & n5708;
  assign n5712 = n1968 & n4957;
  assign n5713 = n5711 & n5712;
  assign n5714 = n1820 & n5710;
  assign n5715 = n5713 & n5714;
  assign n5716 = n5696 & n5702;
  assign n5717 = n5715 & n5716;
  assign n5718 = ~n85 & n5343;
  assign n5719 = ~n92 & ~n253;
  assign n5720 = n3079 & n5719;
  assign n5721 = n5718 & n5720;
  assign n5722 = ~n296 & ~n591;
  assign n5723 = ~n244 & ~n568;
  assign n5724 = n1970 & n5723;
  assign n5725 = ~n145 & ~n210;
  assign n5726 = ~n285 & ~n338;
  assign n5727 = n5725 & n5726;
  assign n5728 = n596 & n1347;
  assign n5729 = n1433 & n1762;
  assign n5730 = n3169 & n3346;
  assign n5731 = n4156 & n5730;
  assign n5732 = n5728 & n5729;
  assign n5733 = n2905 & n5727;
  assign n5734 = n5724 & n5733;
  assign n5735 = n5731 & n5732;
  assign n5736 = n5734 & n5735;
  assign n5737 = n5034 & n5736;
  assign n5738 = ~n192 & ~n420;
  assign n5739 = ~n463 & n5738;
  assign n5740 = n2065 & n5681;
  assign n5741 = n5722 & n5740;
  assign n5742 = n1540 & n5739;
  assign n5743 = n5585 & n5742;
  assign n5744 = n2564 & n5741;
  assign n5745 = n5721 & n5744;
  assign n5746 = n400 & n5743;
  assign n5747 = n5687 & n5746;
  assign n5748 = n5745 & n5747;
  assign n5749 = n5717 & n5737;
  assign n5750 = n5748 & n5749;
  assign n5751 = ~n234 & ~n588;
  assign n5752 = ~n168 & ~n355;
  assign n5753 = ~n389 & ~n466;
  assign n5754 = n5752 & n5753;
  assign n5755 = n298 & n4984;
  assign n5756 = n5751 & n5755;
  assign n5757 = n5754 & n5756;
  assign n5758 = ~n141 & n194;
  assign n5759 = ~n283 & n5758;
  assign n5760 = ~n238 & ~n342;
  assign n5761 = ~n172 & ~n553;
  assign n5762 = ~n641 & ~n681;
  assign n5763 = n5761 & n5762;
  assign n5764 = n885 & n1172;
  assign n5765 = n3078 & n4986;
  assign n5766 = n5760 & n5765;
  assign n5767 = n5763 & n5764;
  assign n5768 = n5766 & n5767;
  assign n5769 = ~n422 & ~n571;
  assign n5770 = n882 & n5769;
  assign n5771 = n1233 & n3826;
  assign n5772 = n5770 & n5771;
  assign n5773 = ~n173 & ~n510;
  assign n5774 = ~n582 & ~n650;
  assign n5775 = n5773 & n5774;
  assign n5776 = n220 & n524;
  assign n5777 = n928 & n1114;
  assign n5778 = n1538 & n2390;
  assign n5779 = n5777 & n5778;
  assign n5780 = n5775 & n5776;
  assign n5781 = n826 & n5780;
  assign n5782 = n4580 & n5779;
  assign n5783 = n5759 & n5772;
  assign n5784 = n5782 & n5783;
  assign n5785 = n5768 & n5781;
  assign n5786 = n5784 & n5785;
  assign n5787 = ~n183 & ~n224;
  assign n5788 = ~n300 & ~n316;
  assign n5789 = ~n659 & n5788;
  assign n5790 = n493 & n5787;
  assign n5791 = n811 & n1944;
  assign n5792 = n2365 & n3844;
  assign n5793 = n5791 & n5792;
  assign n5794 = n5789 & n5790;
  assign n5795 = n5793 & n5794;
  assign n5796 = ~n509 & ~n554;
  assign n5797 = ~n574 & ~n670;
  assign n5798 = n5796 & n5797;
  assign n5799 = n581 & n624;
  assign n5800 = n922 & n1115;
  assign n5801 = n1342 & n3427;
  assign n5802 = n5800 & n5801;
  assign n5803 = n5798 & n5799;
  assign n5804 = n3247 & n5803;
  assign n5805 = n4584 & n5802;
  assign n5806 = n5804 & n5805;
  assign n5807 = n5757 & n5795;
  assign n5808 = n5806 & n5807;
  assign n5809 = n4578 & n5808;
  assign n5810 = n5786 & n5809;
  assign n5811 = ~n5750 & ~n5810;
  assign n5812 = n5750 & n5810;
  assign n5813 = ~n5811 & ~n5812;
  assign n5814 = ~pi8  & n5813;
  assign n5815 = ~n5811 & ~n5814;
  assign n5816 = n5573 & ~n5815;
  assign n5817 = ~n5573 & n5815;
  assign n5818 = ~n5816 & ~n5817;
  assign n5819 = n564 & ~n2622;
  assign n5820 = ~n2538 & n3683;
  assign n5821 = ~n2442 & n3896;
  assign n5822 = n3508 & ~n3510;
  assign n5823 = ~n3511 & ~n5822;
  assign n5824 = n566 & n5823;
  assign n5825 = ~n5819 & ~n5821;
  assign n5826 = ~n5820 & n5825;
  assign n5827 = ~n5824 & n5826;
  assign n5828 = n5818 & ~n5827;
  assign n5829 = ~n5816 & ~n5828;
  assign n5830 = ~n5573 & n5679;
  assign n5831 = ~n5680 & ~n5830;
  assign n5832 = ~n5829 & n5831;
  assign n5833 = ~n5680 & ~n5832;
  assign n5834 = ~n5645 & n5654;
  assign n5835 = ~n5655 & ~n5834;
  assign n5836 = ~n5833 & n5835;
  assign n5837 = ~n5655 & ~n5836;
  assign n5838 = ~n5627 & n5636;
  assign n5839 = ~n5637 & ~n5838;
  assign n5840 = ~n5837 & n5839;
  assign n5841 = n5837 & ~n5839;
  assign n5842 = ~n5840 & ~n5841;
  assign n5843 = ~n2045 & n3943;
  assign n5844 = ~n1997 & n4070;
  assign n5845 = ~n1893 & n4472;
  assign n5846 = n3944 & n5061;
  assign n5847 = ~n5843 & ~n5844;
  assign n5848 = ~n5845 & n5847;
  assign n5849 = ~n5846 & n5848;
  assign n5850 = pi29  & n5849;
  assign n5851 = ~pi29  & ~n5849;
  assign n5852 = ~n5850 & ~n5851;
  assign n5853 = n5842 & ~n5852;
  assign n5854 = ~n5840 & ~n5853;
  assign n5855 = n5643 & ~n5854;
  assign n5856 = ~n5641 & ~n5855;
  assign n5857 = n5522 & ~n5524;
  assign n5858 = ~n5525 & ~n5857;
  assign n5859 = ~n5856 & n5858;
  assign n5860 = ~n5525 & ~n5859;
  assign n5861 = ~n5435 & n5445;
  assign n5862 = ~n5446 & ~n5861;
  assign n5863 = n5860 & ~n5862;
  assign n5864 = ~n5860 & n5862;
  assign n5865 = ~n5863 & ~n5864;
  assign n5866 = ~n1532 & n4515;
  assign n5867 = ~n1425 & n4691;
  assign n5868 = ~n1337 & n4721;
  assign n5869 = n4452 & n4516;
  assign n5870 = ~n5866 & ~n5867;
  assign n5871 = ~n5868 & n5870;
  assign n5872 = ~n5869 & n5871;
  assign n5873 = pi26  & n5872;
  assign n5874 = ~pi26  & ~n5872;
  assign n5875 = ~n5873 & ~n5874;
  assign n5876 = n5865 & n5875;
  assign n5877 = ~n5863 & ~n5876;
  assign n5878 = n5512 & n5877;
  assign n5879 = ~n5512 & ~n5877;
  assign n5880 = ~n5878 & ~n5879;
  assign n5881 = ~n898 & n5267;
  assign n5882 = ~n1006 & n5185;
  assign n5883 = ~n1107 & n5121;
  assign n5884 = n78 & n4041;
  assign n5885 = ~n5881 & ~n5882;
  assign n5886 = ~n5883 & n5885;
  assign n5887 = ~n5884 & n5886;
  assign n5888 = pi23  & n5887;
  assign n5889 = ~pi23  & ~n5887;
  assign n5890 = ~n5888 & ~n5889;
  assign n5891 = n5880 & ~n5890;
  assign n5892 = ~n5878 & ~n5891;
  assign n5893 = n5507 & ~n5509;
  assign n5894 = ~n5510 & ~n5893;
  assign n5895 = ~n5892 & n5894;
  assign n5896 = ~n5510 & ~n5895;
  assign n5897 = ~n5497 & ~n5896;
  assign n5898 = n5497 & n5896;
  assign n5899 = ~n5897 & ~n5898;
  assign n5900 = ~n621 & n5312;
  assign n5901 = ~n5305 & n5310;
  assign n5902 = ~n563 & n5901;
  assign n5903 = n3687 & n5306;
  assign n5904 = ~n5900 & ~n5902;
  assign n5905 = ~n5903 & n5904;
  assign n5906 = pi20  & n5905;
  assign n5907 = ~pi20  & ~n5905;
  assign n5908 = ~n5906 & ~n5907;
  assign n5909 = n5899 & ~n5908;
  assign n5910 = ~n5897 & ~n5909;
  assign n5911 = ~n5486 & ~n5488;
  assign n5912 = ~n5489 & ~n5911;
  assign n5913 = ~n5910 & n5912;
  assign n5914 = n5910 & ~n5912;
  assign n5915 = ~n5913 & ~n5914;
  assign n5916 = ~n5880 & n5890;
  assign n5917 = ~n5891 & ~n5916;
  assign n5918 = ~n5865 & ~n5875;
  assign n5919 = ~n5876 & ~n5918;
  assign n5920 = n5856 & ~n5858;
  assign n5921 = ~n5859 & ~n5920;
  assign n5922 = ~n1610 & n4515;
  assign n5923 = ~n1532 & n4691;
  assign n5924 = ~n1425 & n4721;
  assign n5925 = n4516 & n4642;
  assign n5926 = ~n5922 & ~n5923;
  assign n5927 = ~n5924 & n5926;
  assign n5928 = ~n5925 & n5927;
  assign n5929 = pi26  & n5928;
  assign n5930 = ~pi26  & ~n5928;
  assign n5931 = ~n5929 & ~n5930;
  assign n5932 = n5921 & ~n5931;
  assign n5933 = ~n5643 & n5854;
  assign n5934 = ~n5855 & ~n5933;
  assign n5935 = ~n1997 & n3943;
  assign n5936 = ~n1893 & n4070;
  assign n5937 = ~n1805 & n4472;
  assign n5938 = n3944 & n5212;
  assign n5939 = ~n5935 & ~n5936;
  assign n5940 = ~n5937 & n5939;
  assign n5941 = ~n5938 & n5940;
  assign n5942 = pi29  & n5941;
  assign n5943 = ~pi29  & ~n5941;
  assign n5944 = ~n5942 & ~n5943;
  assign n5945 = n5934 & ~n5944;
  assign n5946 = ~n1737 & n4515;
  assign n5947 = ~n1610 & n4691;
  assign n5948 = ~n1532 & n4721;
  assign n5949 = n4516 & n4626;
  assign n5950 = ~n5946 & ~n5947;
  assign n5951 = ~n5948 & n5950;
  assign n5952 = ~n5949 & n5951;
  assign n5953 = pi26  & n5952;
  assign n5954 = ~pi26  & ~n5952;
  assign n5955 = ~n5953 & ~n5954;
  assign n5956 = ~n5934 & n5944;
  assign n5957 = ~n5945 & ~n5956;
  assign n5958 = ~n5955 & n5957;
  assign n5959 = ~n5945 & ~n5958;
  assign n5960 = ~n5921 & n5931;
  assign n5961 = ~n5932 & ~n5960;
  assign n5962 = ~n5959 & n5961;
  assign n5963 = ~n5932 & ~n5962;
  assign n5964 = n5919 & n5963;
  assign n5965 = ~n5919 & ~n5963;
  assign n5966 = ~n5964 & ~n5965;
  assign n5967 = ~n1107 & n5185;
  assign n5968 = ~n1006 & n5267;
  assign n5969 = ~n1230 & n5121;
  assign n5970 = n78 & n4233;
  assign n5971 = ~n5967 & ~n5968;
  assign n5972 = ~n5969 & n5971;
  assign n5973 = ~n5970 & n5972;
  assign n5974 = pi23  & n5973;
  assign n5975 = ~pi23  & ~n5973;
  assign n5976 = ~n5974 & ~n5975;
  assign n5977 = n5966 & n5976;
  assign n5978 = ~n5964 & ~n5977;
  assign n5979 = n5917 & n5978;
  assign n5980 = ~n5917 & ~n5978;
  assign n5981 = ~n5979 & ~n5980;
  assign n5982 = ~n5302 & n5305;
  assign n5983 = ~n621 & n5982;
  assign n5984 = ~n729 & n5901;
  assign n5985 = ~n802 & n5312;
  assign n5986 = n3955 & n5306;
  assign n5987 = ~n5983 & ~n5985;
  assign n5988 = ~n5984 & n5987;
  assign n5989 = ~n5986 & n5988;
  assign n5990 = pi20  & n5989;
  assign n5991 = ~pi20  & ~n5989;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = n5981 & ~n5992;
  assign n5994 = ~n5979 & ~n5993;
  assign n5995 = ~n729 & n5312;
  assign n5996 = ~n621 & n5901;
  assign n5997 = ~n563 & n5982;
  assign n5998 = n3921 & n5306;
  assign n5999 = ~n5996 & ~n5997;
  assign n6000 = ~n5995 & n5999;
  assign n6001 = ~n5998 & n6000;
  assign n6002 = pi20  & n6001;
  assign n6003 = ~pi20  & ~n6001;
  assign n6004 = ~n6002 & ~n6003;
  assign n6005 = ~n5994 & ~n6004;
  assign n6006 = n5892 & ~n5894;
  assign n6007 = ~n5895 & ~n6006;
  assign n6008 = n5994 & n6004;
  assign n6009 = ~n6005 & ~n6008;
  assign n6010 = n6007 & n6009;
  assign n6011 = ~n6005 & ~n6010;
  assign n6012 = ~n5899 & n5908;
  assign n6013 = ~n5909 & ~n6012;
  assign n6014 = ~n6011 & n6013;
  assign n6015 = n6011 & ~n6013;
  assign n6016 = ~n6014 & ~n6015;
  assign n6017 = ~n5966 & ~n5976;
  assign n6018 = ~n5977 & ~n6017;
  assign n6019 = ~n1337 & n5121;
  assign n6020 = ~n1230 & n5185;
  assign n6021 = ~n1107 & n5267;
  assign n6022 = n78 & n4251;
  assign n6023 = ~n6019 & ~n6020;
  assign n6024 = ~n6021 & n6023;
  assign n6025 = ~n6022 & n6024;
  assign n6026 = ~pi23  & ~n6025;
  assign n6027 = pi23  & n6025;
  assign n6028 = ~n6026 & ~n6027;
  assign n6029 = n5959 & ~n5961;
  assign n6030 = ~n5962 & ~n6029;
  assign n6031 = ~n6028 & n6030;
  assign n6032 = n5955 & ~n5957;
  assign n6033 = ~n5958 & ~n6032;
  assign n6034 = ~n5842 & n5852;
  assign n6035 = ~n5853 & ~n6034;
  assign n6036 = n5829 & ~n5831;
  assign n6037 = ~n5832 & ~n6036;
  assign n6038 = ~n2356 & n3896;
  assign n6039 = n564 & ~n2538;
  assign n6040 = ~n2442 & n3683;
  assign n6041 = n3512 & ~n3514;
  assign n6042 = ~n3515 & ~n6041;
  assign n6043 = n566 & n6042;
  assign n6044 = ~n6038 & ~n6040;
  assign n6045 = ~n6039 & n6044;
  assign n6046 = ~n6043 & n6045;
  assign n6047 = n6037 & ~n6046;
  assign n6048 = ~n2165 & n4070;
  assign n6049 = ~n2265 & n3943;
  assign n6050 = ~n2045 & n4472;
  assign n6051 = n3944 & n5408;
  assign n6052 = ~n6049 & ~n6050;
  assign n6053 = ~n6048 & n6052;
  assign n6054 = ~n6051 & n6053;
  assign n6055 = ~pi29  & ~n6054;
  assign n6056 = pi29  & n6054;
  assign n6057 = ~n6055 & ~n6056;
  assign n6058 = ~n6037 & n6046;
  assign n6059 = ~n6047 & ~n6058;
  assign n6060 = ~n6057 & n6059;
  assign n6061 = ~n6047 & ~n6060;
  assign n6062 = n5833 & ~n5835;
  assign n6063 = ~n5836 & ~n6062;
  assign n6064 = n6061 & ~n6063;
  assign n6065 = ~n2165 & n3943;
  assign n6066 = ~n2045 & n4070;
  assign n6067 = ~n1997 & n4472;
  assign n6068 = n3944 & n5424;
  assign n6069 = ~n6066 & ~n6067;
  assign n6070 = ~n6065 & n6069;
  assign n6071 = ~n6068 & n6070;
  assign n6072 = pi29  & n6071;
  assign n6073 = ~pi29  & ~n6071;
  assign n6074 = ~n6072 & ~n6073;
  assign n6075 = ~n6061 & n6063;
  assign n6076 = ~n6064 & ~n6075;
  assign n6077 = n6074 & n6076;
  assign n6078 = ~n6064 & ~n6077;
  assign n6079 = ~n6035 & ~n6078;
  assign n6080 = n6035 & n6078;
  assign n6081 = ~n6079 & ~n6080;
  assign n6082 = ~n1805 & n4515;
  assign n6083 = ~n1737 & n4691;
  assign n6084 = ~n1610 & n4721;
  assign n6085 = n4516 & n4844;
  assign n6086 = ~n6082 & ~n6083;
  assign n6087 = ~n6084 & n6086;
  assign n6088 = ~n6085 & n6087;
  assign n6089 = pi26  & n6088;
  assign n6090 = ~pi26  & ~n6088;
  assign n6091 = ~n6089 & ~n6090;
  assign n6092 = n6081 & n6091;
  assign n6093 = ~n6079 & ~n6092;
  assign n6094 = n6033 & n6093;
  assign n6095 = ~n6033 & ~n6093;
  assign n6096 = ~n6094 & ~n6095;
  assign n6097 = ~n1425 & n5121;
  assign n6098 = ~n1337 & n5185;
  assign n6099 = ~n1230 & n5267;
  assign n6100 = n78 & n4549;
  assign n6101 = ~n6097 & ~n6098;
  assign n6102 = ~n6099 & n6101;
  assign n6103 = ~n6100 & n6102;
  assign n6104 = pi23  & n6103;
  assign n6105 = ~pi23  & ~n6103;
  assign n6106 = ~n6104 & ~n6105;
  assign n6107 = n6096 & ~n6106;
  assign n6108 = ~n6094 & ~n6107;
  assign n6109 = n6028 & ~n6030;
  assign n6110 = ~n6031 & ~n6109;
  assign n6111 = ~n6108 & n6110;
  assign n6112 = ~n6031 & ~n6111;
  assign n6113 = ~n6018 & ~n6112;
  assign n6114 = n6018 & n6112;
  assign n6115 = ~n6113 & ~n6114;
  assign n6116 = ~n729 & n5982;
  assign n6117 = ~n802 & n5901;
  assign n6118 = ~n898 & n5312;
  assign n6119 = n3901 & n5306;
  assign n6120 = ~n6117 & ~n6118;
  assign n6121 = ~n6116 & n6120;
  assign n6122 = ~n6119 & n6121;
  assign n6123 = pi20  & n6122;
  assign n6124 = ~pi20  & ~n6122;
  assign n6125 = ~n6123 & ~n6124;
  assign n6126 = n6115 & ~n6125;
  assign n6127 = ~n6113 & ~n6126;
  assign n6128 = ~pi14  & ~pi15 ;
  assign n6129 = pi14  & pi15 ;
  assign n6130 = ~n6128 & ~n6129;
  assign n6131 = ~pi16  & ~pi17 ;
  assign n6132 = pi16  & pi17 ;
  assign n6133 = ~n6131 & ~n6132;
  assign n6134 = n6130 & n6133;
  assign n6135 = ~n3593 & n6134;
  assign n6136 = ~pi15  & ~pi16 ;
  assign n6137 = pi15  & pi16 ;
  assign n6138 = ~n6136 & ~n6137;
  assign n6139 = ~n6130 & n6133;
  assign n6140 = ~n6138 & n6139;
  assign n6141 = ~n6135 & ~n6140;
  assign n6142 = ~n563 & ~n6141;
  assign n6143 = pi17  & ~n6142;
  assign n6144 = ~pi17  & n6142;
  assign n6145 = ~n6143 & ~n6144;
  assign n6146 = ~n6127 & ~n6145;
  assign n6147 = n6127 & n6145;
  assign n6148 = ~n6146 & ~n6147;
  assign n6149 = ~n5981 & n5992;
  assign n6150 = ~n5993 & ~n6149;
  assign n6151 = n6148 & n6150;
  assign n6152 = ~n6146 & ~n6151;
  assign n6153 = ~n6007 & ~n6009;
  assign n6154 = ~n6010 & ~n6153;
  assign n6155 = ~n6152 & n6154;
  assign n6156 = ~n6148 & ~n6150;
  assign n6157 = ~n6151 & ~n6156;
  assign n6158 = n6108 & ~n6110;
  assign n6159 = ~n6111 & ~n6158;
  assign n6160 = ~n802 & n5982;
  assign n6161 = ~n898 & n5901;
  assign n6162 = ~n1006 & n5312;
  assign n6163 = n4057 & n5306;
  assign n6164 = ~n6160 & ~n6161;
  assign n6165 = ~n6162 & n6164;
  assign n6166 = ~n6163 & n6165;
  assign n6167 = pi20  & n6166;
  assign n6168 = ~pi20  & ~n6166;
  assign n6169 = ~n6167 & ~n6168;
  assign n6170 = n6159 & ~n6169;
  assign n6171 = ~n6096 & n6106;
  assign n6172 = ~n6107 & ~n6171;
  assign n6173 = ~n6081 & ~n6091;
  assign n6174 = ~n6092 & ~n6173;
  assign n6175 = ~n6074 & ~n6076;
  assign n6176 = ~n6077 & ~n6175;
  assign n6177 = ~n1893 & n4515;
  assign n6178 = ~n1805 & n4691;
  assign n6179 = ~n1737 & n4721;
  assign n6180 = n4516 & n4862;
  assign n6181 = ~n6177 & ~n6178;
  assign n6182 = ~n6179 & n6181;
  assign n6183 = ~n6180 & n6182;
  assign n6184 = pi26  & n6183;
  assign n6185 = ~pi26  & ~n6183;
  assign n6186 = ~n6184 & ~n6185;
  assign n6187 = ~n6176 & ~n6186;
  assign n6188 = ~n244 & ~n597;
  assign n6189 = ~n641 & n6188;
  assign n6190 = n449 & ~n509;
  assign n6191 = n1149 & n6190;
  assign n6192 = ~n222 & ~n235;
  assign n6193 = ~n307 & ~n648;
  assign n6194 = n6192 & n6193;
  assign n6195 = n1868 & n2193;
  assign n6196 = n2390 & n4384;
  assign n6197 = n5760 & n6196;
  assign n6198 = n6194 & n6195;
  assign n6199 = n1013 & n4129;
  assign n6200 = n6198 & n6199;
  assign n6201 = n6191 & n6197;
  assign n6202 = n6200 & n6201;
  assign n6203 = ~n125 & ~n131;
  assign n6204 = ~n207 & ~n310;
  assign n6205 = ~n494 & ~n681;
  assign n6206 = n6204 & n6205;
  assign n6207 = n741 & n6203;
  assign n6208 = n1112 & n1346;
  assign n6209 = n1562 & n4768;
  assign n6210 = n6208 & n6209;
  assign n6211 = n6206 & n6207;
  assign n6212 = n6189 & n6211;
  assign n6213 = n5772 & n6210;
  assign n6214 = n6212 & n6213;
  assign n6215 = n5687 & n6214;
  assign n6216 = n1625 & n6202;
  assign n6217 = n6215 & n6216;
  assign n6218 = n4381 & n6217;
  assign n6219 = n5750 & ~n6218;
  assign n6220 = ~n387 & ~n570;
  assign n6221 = ~n463 & ~n473;
  assign n6222 = ~n651 & n6221;
  assign n6223 = n1147 & n2298;
  assign n6224 = n2324 & n6223;
  assign n6225 = n6222 & n6224;
  assign n6226 = ~n522 & n668;
  assign n6227 = n731 & n1203;
  assign n6228 = n2598 & n3072;
  assign n6229 = n6220 & n6228;
  assign n6230 = n6226 & n6227;
  assign n6231 = n1583 & n3981;
  assign n6232 = n6230 & n6231;
  assign n6233 = n1236 & n6229;
  assign n6234 = n6232 & n6233;
  assign n6235 = n1278 & n6225;
  assign n6236 = n6234 & n6235;
  assign n6237 = n3806 & n6236;
  assign n6238 = n5022 & n6237;
  assign n6239 = ~pi2  & ~n6238;
  assign n6240 = pi2  & n6238;
  assign n6241 = ~n6239 & ~n6240;
  assign n6242 = ~pi5  & n6241;
  assign n6243 = ~n6239 & ~n6242;
  assign n6244 = n5750 & ~n6243;
  assign n6245 = ~n5750 & n6243;
  assign n6246 = ~n6244 & ~n6245;
  assign n6247 = ~n2657 & n3896;
  assign n6248 = ~n2726 & n3683;
  assign n6249 = n564 & ~n2781;
  assign n6250 = n3496 & ~n3498;
  assign n6251 = ~n3499 & ~n6250;
  assign n6252 = n566 & n6251;
  assign n6253 = ~n6247 & ~n6249;
  assign n6254 = ~n6248 & n6253;
  assign n6255 = ~n6252 & n6254;
  assign n6256 = n6246 & ~n6255;
  assign n6257 = ~n6244 & ~n6256;
  assign n6258 = ~n5750 & n6218;
  assign n6259 = ~n6219 & ~n6258;
  assign n6260 = ~n6257 & n6259;
  assign n6261 = ~n6219 & ~n6260;
  assign n6262 = pi8  & ~n5813;
  assign n6263 = ~n5814 & ~n6262;
  assign n6264 = ~n6261 & n6263;
  assign n6265 = n6261 & ~n6263;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = ~n2538 & n3896;
  assign n6268 = ~n2622 & n3683;
  assign n6269 = n564 & ~n2657;
  assign n6270 = n3504 & ~n3506;
  assign n6271 = ~n3507 & ~n6270;
  assign n6272 = n566 & n6271;
  assign n6273 = ~n6267 & ~n6269;
  assign n6274 = ~n6268 & n6273;
  assign n6275 = ~n6272 & n6274;
  assign n6276 = n6266 & ~n6275;
  assign n6277 = ~n6264 & ~n6276;
  assign n6278 = ~n5818 & n5827;
  assign n6279 = ~n5828 & ~n6278;
  assign n6280 = ~n6277 & n6279;
  assign n6281 = n6277 & ~n6279;
  assign n6282 = ~n6280 & ~n6281;
  assign n6283 = ~n2356 & n3943;
  assign n6284 = ~n2265 & n4070;
  assign n6285 = ~n2165 & n4472;
  assign n6286 = n3944 & n5632;
  assign n6287 = ~n6283 & ~n6284;
  assign n6288 = ~n6285 & n6287;
  assign n6289 = ~n6286 & n6288;
  assign n6290 = pi29  & n6289;
  assign n6291 = ~pi29  & ~n6289;
  assign n6292 = ~n6290 & ~n6291;
  assign n6293 = n6282 & ~n6292;
  assign n6294 = ~n6280 & ~n6293;
  assign n6295 = n6057 & ~n6059;
  assign n6296 = ~n6060 & ~n6295;
  assign n6297 = ~n6294 & n6296;
  assign n6298 = n6294 & ~n6296;
  assign n6299 = ~n6297 & ~n6298;
  assign n6300 = ~n1997 & n4515;
  assign n6301 = ~n1893 & n4691;
  assign n6302 = ~n1805 & n4721;
  assign n6303 = n4516 & n5212;
  assign n6304 = ~n6300 & ~n6301;
  assign n6305 = ~n6302 & n6304;
  assign n6306 = ~n6303 & n6305;
  assign n6307 = pi26  & n6306;
  assign n6308 = ~pi26  & ~n6306;
  assign n6309 = ~n6307 & ~n6308;
  assign n6310 = n6299 & ~n6309;
  assign n6311 = ~n6297 & ~n6310;
  assign n6312 = n6176 & n6186;
  assign n6313 = ~n6187 & ~n6312;
  assign n6314 = ~n6311 & n6313;
  assign n6315 = ~n6187 & ~n6314;
  assign n6316 = n6174 & n6315;
  assign n6317 = ~n6174 & ~n6315;
  assign n6318 = ~n6316 & ~n6317;
  assign n6319 = ~n1532 & n5121;
  assign n6320 = ~n1425 & n5185;
  assign n6321 = ~n1337 & n5267;
  assign n6322 = n78 & n4452;
  assign n6323 = ~n6319 & ~n6320;
  assign n6324 = ~n6321 & n6323;
  assign n6325 = ~n6322 & n6324;
  assign n6326 = pi23  & n6325;
  assign n6327 = ~pi23  & ~n6325;
  assign n6328 = ~n6326 & ~n6327;
  assign n6329 = n6318 & n6328;
  assign n6330 = ~n6316 & ~n6329;
  assign n6331 = n6172 & n6330;
  assign n6332 = ~n6172 & ~n6330;
  assign n6333 = ~n6331 & ~n6332;
  assign n6334 = ~n898 & n5982;
  assign n6335 = ~n1006 & n5901;
  assign n6336 = ~n1107 & n5312;
  assign n6337 = n4041 & n5306;
  assign n6338 = ~n6334 & ~n6335;
  assign n6339 = ~n6336 & n6338;
  assign n6340 = ~n6337 & n6339;
  assign n6341 = pi20  & n6340;
  assign n6342 = ~pi20  & ~n6340;
  assign n6343 = ~n6341 & ~n6342;
  assign n6344 = n6333 & ~n6343;
  assign n6345 = ~n6331 & ~n6344;
  assign n6346 = ~n6159 & n6169;
  assign n6347 = ~n6170 & ~n6346;
  assign n6348 = ~n6345 & n6347;
  assign n6349 = ~n6170 & ~n6348;
  assign n6350 = ~n6115 & n6125;
  assign n6351 = ~n6126 & ~n6350;
  assign n6352 = n6349 & ~n6351;
  assign n6353 = ~n6349 & n6351;
  assign n6354 = ~n6352 & ~n6353;
  assign n6355 = ~n621 & n6140;
  assign n6356 = ~n6130 & n6138;
  assign n6357 = ~n563 & n6356;
  assign n6358 = n3687 & n6134;
  assign n6359 = ~n6355 & ~n6357;
  assign n6360 = ~n6358 & n6359;
  assign n6361 = pi17  & n6360;
  assign n6362 = ~pi17  & ~n6360;
  assign n6363 = ~n6361 & ~n6362;
  assign n6364 = n6354 & n6363;
  assign n6365 = ~n6352 & ~n6364;
  assign n6366 = n6157 & n6365;
  assign n6367 = ~n6157 & ~n6365;
  assign n6368 = ~n6366 & ~n6367;
  assign n6369 = ~n6354 & ~n6363;
  assign n6370 = ~n6364 & ~n6369;
  assign n6371 = ~n6318 & ~n6328;
  assign n6372 = ~n6329 & ~n6371;
  assign n6373 = ~n1610 & n5121;
  assign n6374 = ~n1532 & n5185;
  assign n6375 = ~n1425 & n5267;
  assign n6376 = n78 & n4642;
  assign n6377 = ~n6373 & ~n6374;
  assign n6378 = ~n6375 & n6377;
  assign n6379 = ~n6376 & n6378;
  assign n6380 = ~pi23  & ~n6379;
  assign n6381 = pi23  & n6379;
  assign n6382 = ~n6380 & ~n6381;
  assign n6383 = n6311 & ~n6313;
  assign n6384 = ~n6314 & ~n6383;
  assign n6385 = ~n6382 & n6384;
  assign n6386 = ~n6299 & n6309;
  assign n6387 = ~n6310 & ~n6386;
  assign n6388 = ~n2356 & n4070;
  assign n6389 = ~n2442 & n3943;
  assign n6390 = ~n2265 & n4472;
  assign n6391 = n3944 & n5650;
  assign n6392 = ~n6389 & ~n6390;
  assign n6393 = ~n6388 & n6392;
  assign n6394 = ~n6391 & n6393;
  assign n6395 = ~pi29  & ~n6394;
  assign n6396 = pi29  & n6394;
  assign n6397 = ~n6395 & ~n6396;
  assign n6398 = ~n6266 & n6275;
  assign n6399 = ~n6276 & ~n6398;
  assign n6400 = ~n6397 & n6399;
  assign n6401 = n6257 & ~n6259;
  assign n6402 = ~n6260 & ~n6401;
  assign n6403 = ~n2622 & n3896;
  assign n6404 = n564 & ~n2726;
  assign n6405 = ~n2657 & n3683;
  assign n6406 = n3500 & ~n3502;
  assign n6407 = ~n3503 & ~n6406;
  assign n6408 = n566 & n6407;
  assign n6409 = ~n6403 & ~n6405;
  assign n6410 = ~n6404 & n6409;
  assign n6411 = ~n6408 & n6410;
  assign n6412 = n6402 & ~n6411;
  assign n6413 = ~n225 & ~n597;
  assign n6414 = ~n599 & n6413;
  assign n6415 = n987 & n2830;
  assign n6416 = n6414 & n6415;
  assign n6417 = ~n388 & ~n426;
  assign n6418 = ~n577 & n6417;
  assign n6419 = n848 & n1083;
  assign n6420 = n3352 & n3419;
  assign n6421 = n6419 & n6420;
  assign n6422 = n6418 & n6421;
  assign n6423 = ~n387 & ~n480;
  assign n6424 = n1536 & n6423;
  assign n6425 = n3763 & n3994;
  assign n6426 = n4932 & n6425;
  assign n6427 = n1207 & n6424;
  assign n6428 = n5577 & n5657;
  assign n6429 = n6427 & n6428;
  assign n6430 = n1921 & n6426;
  assign n6431 = n6416 & n6430;
  assign n6432 = n6422 & n6429;
  assign n6433 = n6431 & n6432;
  assign n6434 = n161 & n6433;
  assign n6435 = n2817 & n3103;
  assign n6436 = n6434 & n6435;
  assign n6437 = pi2  & ~n6436;
  assign n6438 = n1536 & n1594;
  assign n6439 = n4093 & n6438;
  assign n6440 = ~n467 & ~n543;
  assign n6441 = ~n163 & ~n238;
  assign n6442 = ~n321 & ~n522;
  assign n6443 = n6441 & n6442;
  assign n6444 = n217 & n537;
  assign n6445 = n2226 & n5368;
  assign n6446 = n6440 & n6445;
  assign n6447 = n6443 & n6444;
  assign n6448 = n1053 & n4555;
  assign n6449 = n6447 & n6448;
  assign n6450 = n1245 & n6446;
  assign n6451 = n4915 & n6439;
  assign n6452 = n6450 & n6451;
  assign n6453 = n3777 & n6449;
  assign n6454 = n6452 & n6453;
  assign n6455 = n1373 & n6454;
  assign n6456 = n3302 & n6455;
  assign n6457 = pi2  & ~n6456;
  assign n6458 = ~n175 & ~n271;
  assign n6459 = ~n315 & ~n363;
  assign n6460 = ~n601 & n6459;
  assign n6461 = n537 & n6458;
  assign n6462 = n600 & n1118;
  assign n6463 = n2190 & n3855;
  assign n6464 = n6462 & n6463;
  assign n6465 = n6460 & n6461;
  assign n6466 = n1207 & n3268;
  assign n6467 = n5659 & n6466;
  assign n6468 = n6464 & n6465;
  assign n6469 = n5721 & n6468;
  assign n6470 = n6467 & n6469;
  assign n6471 = ~n149 & ~n203;
  assign n6472 = ~n424 & ~n496;
  assign n6473 = ~n640 & n6472;
  assign n6474 = n573 & n6471;
  assign n6475 = n6473 & n6474;
  assign n6476 = ~n192 & ~n482;
  assign n6477 = n1382 & n6476;
  assign n6478 = n2923 & n3381;
  assign n6479 = n3763 & n4911;
  assign n6480 = n5339 & n6479;
  assign n6481 = n6477 & n6478;
  assign n6482 = n3871 & n6481;
  assign n6483 = n6475 & n6480;
  assign n6484 = n6482 & n6483;
  assign n6485 = n3399 & n3852;
  assign n6486 = n6484 & n6485;
  assign n6487 = n6470 & n6486;
  assign n6488 = n2128 & n6487;
  assign n6489 = pi2  & ~n6488;
  assign n6490 = ~pi2  & n6488;
  assign n6491 = ~n6489 & ~n6490;
  assign n6492 = ~n2901 & n3896;
  assign n6493 = ~n2978 & n3683;
  assign n6494 = n564 & ~n3069;
  assign n6495 = n3480 & ~n3482;
  assign n6496 = ~n3483 & ~n6495;
  assign n6497 = n566 & n6496;
  assign n6498 = ~n6492 & ~n6494;
  assign n6499 = ~n6493 & n6498;
  assign n6500 = ~n6497 & n6499;
  assign n6501 = n6491 & ~n6500;
  assign n6502 = ~n6489 & ~n6501;
  assign n6503 = ~pi2  & n6456;
  assign n6504 = ~n6457 & ~n6503;
  assign n6505 = ~n6502 & n6504;
  assign n6506 = ~n6457 & ~n6505;
  assign n6507 = ~pi2  & n6436;
  assign n6508 = ~n6437 & ~n6507;
  assign n6509 = ~n6506 & n6508;
  assign n6510 = ~n6437 & ~n6509;
  assign n6511 = pi5  & ~n6241;
  assign n6512 = ~n6242 & ~n6511;
  assign n6513 = ~n6510 & n6512;
  assign n6514 = n6510 & ~n6512;
  assign n6515 = ~n6513 & ~n6514;
  assign n6516 = n564 & ~n2866;
  assign n6517 = ~n2726 & n3896;
  assign n6518 = ~n2781 & n3683;
  assign n6519 = n3492 & ~n3494;
  assign n6520 = ~n3495 & ~n6519;
  assign n6521 = n566 & n6520;
  assign n6522 = ~n6516 & ~n6518;
  assign n6523 = ~n6517 & n6522;
  assign n6524 = ~n6521 & n6523;
  assign n6525 = n6515 & ~n6524;
  assign n6526 = ~n6513 & ~n6525;
  assign n6527 = ~n6246 & n6255;
  assign n6528 = ~n6256 & ~n6527;
  assign n6529 = ~n6526 & n6528;
  assign n6530 = n6526 & ~n6528;
  assign n6531 = ~n6529 & ~n6530;
  assign n6532 = ~n2622 & n3943;
  assign n6533 = ~n2538 & n4070;
  assign n6534 = ~n2442 & n4472;
  assign n6535 = n3944 & n5823;
  assign n6536 = ~n6532 & ~n6534;
  assign n6537 = ~n6533 & n6536;
  assign n6538 = ~n6535 & n6537;
  assign n6539 = pi29  & n6538;
  assign n6540 = ~pi29  & ~n6538;
  assign n6541 = ~n6539 & ~n6540;
  assign n6542 = n6531 & ~n6541;
  assign n6543 = ~n6529 & ~n6542;
  assign n6544 = ~n6402 & n6411;
  assign n6545 = ~n6412 & ~n6544;
  assign n6546 = ~n6543 & n6545;
  assign n6547 = ~n6412 & ~n6546;
  assign n6548 = n6397 & ~n6399;
  assign n6549 = ~n6400 & ~n6548;
  assign n6550 = ~n6547 & n6549;
  assign n6551 = ~n6400 & ~n6550;
  assign n6552 = ~n6282 & n6292;
  assign n6553 = ~n6293 & ~n6552;
  assign n6554 = n6551 & ~n6553;
  assign n6555 = ~n6551 & n6553;
  assign n6556 = ~n6554 & ~n6555;
  assign n6557 = ~n2045 & n4515;
  assign n6558 = ~n1997 & n4691;
  assign n6559 = ~n1893 & n4721;
  assign n6560 = n4516 & n5061;
  assign n6561 = ~n6557 & ~n6558;
  assign n6562 = ~n6559 & n6561;
  assign n6563 = ~n6560 & n6562;
  assign n6564 = pi26  & n6563;
  assign n6565 = ~pi26  & ~n6563;
  assign n6566 = ~n6564 & ~n6565;
  assign n6567 = n6556 & n6566;
  assign n6568 = ~n6554 & ~n6567;
  assign n6569 = n6387 & n6568;
  assign n6570 = ~n6387 & ~n6568;
  assign n6571 = ~n6569 & ~n6570;
  assign n6572 = ~n1737 & n5121;
  assign n6573 = ~n1610 & n5185;
  assign n6574 = ~n1532 & n5267;
  assign n6575 = n78 & n4626;
  assign n6576 = ~n6572 & ~n6573;
  assign n6577 = ~n6574 & n6576;
  assign n6578 = ~n6575 & n6577;
  assign n6579 = pi23  & n6578;
  assign n6580 = ~pi23  & ~n6578;
  assign n6581 = ~n6579 & ~n6580;
  assign n6582 = n6571 & ~n6581;
  assign n6583 = ~n6569 & ~n6582;
  assign n6584 = n6382 & ~n6384;
  assign n6585 = ~n6385 & ~n6584;
  assign n6586 = ~n6583 & n6585;
  assign n6587 = ~n6385 & ~n6586;
  assign n6588 = ~n6372 & ~n6587;
  assign n6589 = n6372 & n6587;
  assign n6590 = ~n6588 & ~n6589;
  assign n6591 = ~n1107 & n5901;
  assign n6592 = ~n1006 & n5982;
  assign n6593 = ~n1230 & n5312;
  assign n6594 = n4233 & n5306;
  assign n6595 = ~n6591 & ~n6592;
  assign n6596 = ~n6593 & n6595;
  assign n6597 = ~n6594 & n6596;
  assign n6598 = pi20  & n6597;
  assign n6599 = ~pi20  & ~n6597;
  assign n6600 = ~n6598 & ~n6599;
  assign n6601 = n6590 & ~n6600;
  assign n6602 = ~n6588 & ~n6601;
  assign n6603 = ~n6333 & n6343;
  assign n6604 = ~n6344 & ~n6603;
  assign n6605 = ~n6602 & n6604;
  assign n6606 = n6602 & ~n6604;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = n6130 & ~n6133;
  assign n6609 = ~n621 & n6608;
  assign n6610 = ~n729 & n6356;
  assign n6611 = ~n802 & n6140;
  assign n6612 = n3955 & n6134;
  assign n6613 = ~n6609 & ~n6611;
  assign n6614 = ~n6610 & n6613;
  assign n6615 = ~n6612 & n6614;
  assign n6616 = pi17  & n6615;
  assign n6617 = ~pi17  & ~n6615;
  assign n6618 = ~n6616 & ~n6617;
  assign n6619 = n6607 & ~n6618;
  assign n6620 = ~n6605 & ~n6619;
  assign n6621 = ~n729 & n6140;
  assign n6622 = ~n621 & n6356;
  assign n6623 = ~n563 & n6608;
  assign n6624 = n3921 & n6134;
  assign n6625 = ~n6622 & ~n6623;
  assign n6626 = ~n6621 & n6625;
  assign n6627 = ~n6624 & n6626;
  assign n6628 = pi17  & n6627;
  assign n6629 = ~pi17  & ~n6627;
  assign n6630 = ~n6628 & ~n6629;
  assign n6631 = ~n6620 & ~n6630;
  assign n6632 = n6620 & n6630;
  assign n6633 = ~n6631 & ~n6632;
  assign n6634 = n6345 & ~n6347;
  assign n6635 = ~n6348 & ~n6634;
  assign n6636 = n6633 & n6635;
  assign n6637 = ~n6631 & ~n6636;
  assign n6638 = ~n6370 & ~n6637;
  assign n6639 = n6370 & n6637;
  assign n6640 = ~n6638 & ~n6639;
  assign n6641 = ~pi11  & ~pi12 ;
  assign n6642 = pi11  & pi12 ;
  assign n6643 = ~n6641 & ~n6642;
  assign n6644 = ~pi13  & ~pi14 ;
  assign n6645 = pi13  & pi14 ;
  assign n6646 = ~n6644 & ~n6645;
  assign n6647 = n6643 & n6646;
  assign n6648 = ~n3593 & n6647;
  assign n6649 = ~pi12  & ~pi13 ;
  assign n6650 = pi12  & pi13 ;
  assign n6651 = ~n6649 & ~n6650;
  assign n6652 = ~n6643 & n6646;
  assign n6653 = ~n6651 & n6652;
  assign n6654 = ~n6648 & ~n6653;
  assign n6655 = ~n563 & ~n6654;
  assign n6656 = pi14  & ~n6655;
  assign n6657 = ~pi14  & n6655;
  assign n6658 = ~n6656 & ~n6657;
  assign n6659 = n6583 & ~n6585;
  assign n6660 = ~n6586 & ~n6659;
  assign n6661 = ~n1337 & n5312;
  assign n6662 = ~n1230 & n5901;
  assign n6663 = ~n1107 & n5982;
  assign n6664 = n4251 & n5306;
  assign n6665 = ~n6661 & ~n6662;
  assign n6666 = ~n6663 & n6665;
  assign n6667 = ~n6664 & n6666;
  assign n6668 = pi20  & n6667;
  assign n6669 = ~pi20  & ~n6667;
  assign n6670 = ~n6668 & ~n6669;
  assign n6671 = n6660 & ~n6670;
  assign n6672 = ~n6571 & n6581;
  assign n6673 = ~n6582 & ~n6672;
  assign n6674 = ~n6556 & ~n6566;
  assign n6675 = ~n6567 & ~n6674;
  assign n6676 = n6547 & ~n6549;
  assign n6677 = ~n6550 & ~n6676;
  assign n6678 = ~n2165 & n4515;
  assign n6679 = ~n2045 & n4691;
  assign n6680 = ~n1997 & n4721;
  assign n6681 = n4516 & n5424;
  assign n6682 = ~n6679 & ~n6680;
  assign n6683 = ~n6678 & n6682;
  assign n6684 = ~n6681 & n6683;
  assign n6685 = pi26  & n6684;
  assign n6686 = ~pi26  & ~n6684;
  assign n6687 = ~n6685 & ~n6686;
  assign n6688 = n6677 & ~n6687;
  assign n6689 = ~n2356 & n4472;
  assign n6690 = ~n2538 & n3943;
  assign n6691 = ~n2442 & n4070;
  assign n6692 = n3944 & n6042;
  assign n6693 = ~n6689 & ~n6691;
  assign n6694 = ~n6690 & n6693;
  assign n6695 = ~n6692 & n6694;
  assign n6696 = pi29  & n6695;
  assign n6697 = ~pi29  & ~n6695;
  assign n6698 = ~n6696 & ~n6697;
  assign n6699 = n6543 & ~n6545;
  assign n6700 = ~n6546 & ~n6699;
  assign n6701 = ~n6698 & n6700;
  assign n6702 = n6698 & ~n6700;
  assign n6703 = ~n6701 & ~n6702;
  assign n6704 = ~n2165 & n4691;
  assign n6705 = ~n2265 & n4515;
  assign n6706 = ~n2045 & n4721;
  assign n6707 = n4516 & n5408;
  assign n6708 = ~n6705 & ~n6706;
  assign n6709 = ~n6704 & n6708;
  assign n6710 = ~n6707 & n6709;
  assign n6711 = pi26  & n6710;
  assign n6712 = ~pi26  & ~n6710;
  assign n6713 = ~n6711 & ~n6712;
  assign n6714 = n6703 & ~n6713;
  assign n6715 = ~n6701 & ~n6714;
  assign n6716 = ~n6677 & n6687;
  assign n6717 = ~n6688 & ~n6716;
  assign n6718 = ~n6715 & n6717;
  assign n6719 = ~n6688 & ~n6718;
  assign n6720 = n6675 & n6719;
  assign n6721 = ~n6675 & ~n6719;
  assign n6722 = ~n6720 & ~n6721;
  assign n6723 = ~n1805 & n5121;
  assign n6724 = ~n1737 & n5185;
  assign n6725 = ~n1610 & n5267;
  assign n6726 = n78 & n4844;
  assign n6727 = ~n6723 & ~n6724;
  assign n6728 = ~n6725 & n6727;
  assign n6729 = ~n6726 & n6728;
  assign n6730 = pi23  & n6729;
  assign n6731 = ~pi23  & ~n6729;
  assign n6732 = ~n6730 & ~n6731;
  assign n6733 = n6722 & n6732;
  assign n6734 = ~n6720 & ~n6733;
  assign n6735 = n6673 & n6734;
  assign n6736 = ~n6673 & ~n6734;
  assign n6737 = ~n6735 & ~n6736;
  assign n6738 = ~n1425 & n5312;
  assign n6739 = ~n1337 & n5901;
  assign n6740 = ~n1230 & n5982;
  assign n6741 = n4549 & n5306;
  assign n6742 = ~n6738 & ~n6739;
  assign n6743 = ~n6740 & n6742;
  assign n6744 = ~n6741 & n6743;
  assign n6745 = pi20  & n6744;
  assign n6746 = ~pi20  & ~n6744;
  assign n6747 = ~n6745 & ~n6746;
  assign n6748 = n6737 & ~n6747;
  assign n6749 = ~n6735 & ~n6748;
  assign n6750 = ~n6660 & n6670;
  assign n6751 = ~n6671 & ~n6750;
  assign n6752 = ~n6749 & n6751;
  assign n6753 = ~n6671 & ~n6752;
  assign n6754 = ~n6590 & n6600;
  assign n6755 = ~n6601 & ~n6754;
  assign n6756 = n6753 & ~n6755;
  assign n6757 = ~n6753 & n6755;
  assign n6758 = ~n6756 & ~n6757;
  assign n6759 = ~n729 & n6608;
  assign n6760 = ~n802 & n6356;
  assign n6761 = ~n898 & n6140;
  assign n6762 = n3901 & n6134;
  assign n6763 = ~n6760 & ~n6761;
  assign n6764 = ~n6759 & n6763;
  assign n6765 = ~n6762 & n6764;
  assign n6766 = pi17  & n6765;
  assign n6767 = ~pi17  & ~n6765;
  assign n6768 = ~n6766 & ~n6767;
  assign n6769 = n6758 & n6768;
  assign n6770 = ~n6756 & ~n6769;
  assign n6771 = ~n6658 & n6770;
  assign n6772 = n6658 & ~n6770;
  assign n6773 = ~n6771 & ~n6772;
  assign n6774 = ~n6607 & n6618;
  assign n6775 = ~n6619 & ~n6774;
  assign n6776 = n6773 & n6775;
  assign n6777 = ~n6771 & ~n6776;
  assign n6778 = ~n6633 & ~n6635;
  assign n6779 = ~n6636 & ~n6778;
  assign n6780 = ~n6777 & n6779;
  assign n6781 = n6777 & ~n6779;
  assign n6782 = ~n6780 & ~n6781;
  assign n6783 = ~n802 & n6608;
  assign n6784 = ~n898 & n6356;
  assign n6785 = ~n1006 & n6140;
  assign n6786 = n4057 & n6134;
  assign n6787 = ~n6783 & ~n6784;
  assign n6788 = ~n6785 & n6787;
  assign n6789 = ~n6786 & n6788;
  assign n6790 = ~pi17  & ~n6789;
  assign n6791 = pi17  & n6789;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = n6749 & ~n6751;
  assign n6794 = ~n6752 & ~n6793;
  assign n6795 = ~n6792 & n6794;
  assign n6796 = ~n6722 & ~n6732;
  assign n6797 = ~n6733 & ~n6796;
  assign n6798 = ~n1893 & n5121;
  assign n6799 = ~n1805 & n5185;
  assign n6800 = ~n1737 & n5267;
  assign n6801 = n78 & n4862;
  assign n6802 = ~n6798 & ~n6799;
  assign n6803 = ~n6800 & n6802;
  assign n6804 = ~n6801 & n6803;
  assign n6805 = ~pi23  & ~n6804;
  assign n6806 = pi23  & n6804;
  assign n6807 = ~n6805 & ~n6806;
  assign n6808 = n6715 & ~n6717;
  assign n6809 = ~n6718 & ~n6808;
  assign n6810 = ~n6807 & n6809;
  assign n6811 = ~n6703 & n6713;
  assign n6812 = ~n6714 & ~n6811;
  assign n6813 = n6506 & ~n6508;
  assign n6814 = ~n6509 & ~n6813;
  assign n6815 = ~n2866 & n3683;
  assign n6816 = n564 & ~n2901;
  assign n6817 = ~n2781 & n3896;
  assign n6818 = n3488 & ~n3490;
  assign n6819 = ~n3491 & ~n6818;
  assign n6820 = n566 & n6819;
  assign n6821 = ~n6815 & ~n6816;
  assign n6822 = ~n6817 & n6821;
  assign n6823 = ~n6820 & n6822;
  assign n6824 = n6814 & ~n6823;
  assign n6825 = n6502 & ~n6504;
  assign n6826 = ~n6505 & ~n6825;
  assign n6827 = ~n2866 & n3896;
  assign n6828 = n564 & ~n2978;
  assign n6829 = ~n2901 & n3683;
  assign n6830 = n3484 & ~n3486;
  assign n6831 = ~n3487 & ~n6830;
  assign n6832 = n566 & n6831;
  assign n6833 = ~n6827 & ~n6829;
  assign n6834 = ~n6828 & n6833;
  assign n6835 = ~n6832 & n6834;
  assign n6836 = n6826 & ~n6835;
  assign n6837 = ~n251 & n1268;
  assign n6838 = n5722 & n6837;
  assign n6839 = ~n219 & ~n577;
  assign n6840 = n660 & n6839;
  assign n6841 = ~n286 & ~n308;
  assign n6842 = ~n543 & ~n665;
  assign n6843 = ~n671 & n6842;
  assign n6844 = n366 & n6841;
  assign n6845 = n688 & n969;
  assign n6846 = n1783 & n1965;
  assign n6847 = n3266 & n5023;
  assign n6848 = n5368 & n6847;
  assign n6849 = n6845 & n6846;
  assign n6850 = n6843 & n6844;
  assign n6851 = n6849 & n6850;
  assign n6852 = n4910 & n6848;
  assign n6853 = n6851 & n6852;
  assign n6854 = n2606 & n6853;
  assign n6855 = ~n381 & n537;
  assign n6856 = n1147 & n1595;
  assign n6857 = n1689 & n2472;
  assign n6858 = n2639 & n3196;
  assign n6859 = n6857 & n6858;
  assign n6860 = n6855 & n6856;
  assign n6861 = n249 & n3783;
  assign n6862 = n6840 & n6861;
  assign n6863 = n6859 & n6860;
  assign n6864 = n6838 & n6863;
  assign n6865 = n6862 & n6864;
  assign n6866 = n5010 & n6865;
  assign n6867 = n5000 & n6854;
  assign n6868 = n6866 & n6867;
  assign n6869 = ~n2978 & n3896;
  assign n6870 = n564 & ~n3137;
  assign n6871 = ~n3069 & n3683;
  assign n6872 = n3476 & ~n3478;
  assign n6873 = ~n3479 & ~n6872;
  assign n6874 = n566 & n6873;
  assign n6875 = ~n6869 & ~n6871;
  assign n6876 = ~n6870 & n6875;
  assign n6877 = ~n6874 & n6876;
  assign n6878 = ~n6868 & ~n6877;
  assign n6879 = ~n326 & ~n582;
  assign n6880 = n1970 & n6879;
  assign n6881 = ~n338 & ~n374;
  assign n6882 = ~n588 & n6881;
  assign n6883 = ~n120 & ~n270;
  assign n6884 = ~n387 & ~n674;
  assign n6885 = ~n682 & n6884;
  assign n6886 = n223 & n6883;
  assign n6887 = n403 & n1148;
  assign n6888 = n1342 & n5660;
  assign n6889 = n6887 & n6888;
  assign n6890 = n6885 & n6886;
  assign n6891 = n5528 & n6882;
  assign n6892 = n6890 & n6891;
  assign n6893 = n4794 & n6889;
  assign n6894 = n6892 & n6893;
  assign n6895 = ~n144 & ~n282;
  assign n6896 = ~n342 & ~n375;
  assign n6897 = n6895 & n6896;
  assign n6898 = n1469 & n6897;
  assign n6899 = ~n216 & ~n661;
  assign n6900 = n497 & n6899;
  assign n6901 = n1174 & n1486;
  assign n6902 = n1786 & n2452;
  assign n6903 = n2472 & n2474;
  assign n6904 = n2944 & n3700;
  assign n6905 = n3870 & n6904;
  assign n6906 = n6902 & n6903;
  assign n6907 = n6900 & n6901;
  assign n6908 = n970 & n6880;
  assign n6909 = n6907 & n6908;
  assign n6910 = n6905 & n6906;
  assign n6911 = n6898 & n6910;
  assign n6912 = n5583 & n6909;
  assign n6913 = n6911 & n6912;
  assign n6914 = n1411 & n6894;
  assign n6915 = n6913 & n6914;
  assign n6916 = ~n3069 & n3896;
  assign n6917 = ~n3137 & n3683;
  assign n6918 = n564 & ~n3194;
  assign n6919 = n3472 & ~n3474;
  assign n6920 = ~n3475 & ~n6919;
  assign n6921 = n566 & n6920;
  assign n6922 = ~n6916 & ~n6918;
  assign n6923 = ~n6917 & n6922;
  assign n6924 = ~n6921 & n6923;
  assign n6925 = ~n6915 & ~n6924;
  assign n6926 = ~n196 & ~n426;
  assign n6927 = ~n522 & ~n597;
  assign n6928 = ~n686 & n6927;
  assign n6929 = n1342 & n6926;
  assign n6930 = n1355 & n2945;
  assign n6931 = n6929 & n6930;
  assign n6932 = n1740 & n6928;
  assign n6933 = n6931 & n6932;
  assign n6934 = ~n113 & ~n568;
  assign n6935 = n2823 & n6934;
  assign n6936 = ~n271 & ~n482;
  assign n6937 = ~n545 & n6936;
  assign n6938 = n743 & n6937;
  assign n6939 = ~n212 & ~n584;
  assign n6940 = ~n594 & n6939;
  assign n6941 = n471 & n3106;
  assign n6942 = n1233 & n2193;
  assign n6943 = n2359 & n2633;
  assign n6944 = n6942 & n6943;
  assign n6945 = n6940 & n6941;
  assign n6946 = n2406 & n6945;
  assign n6947 = n5663 & n6944;
  assign n6948 = n6935 & n6938;
  assign n6949 = n6947 & n6948;
  assign n6950 = n6946 & n6949;
  assign n6951 = ~n253 & n3842;
  assign n6952 = n2884 & n6951;
  assign n6953 = ~n236 & ~n335;
  assign n6954 = ~n381 & ~n447;
  assign n6955 = ~n553 & ~n598;
  assign n6956 = n6954 & n6955;
  assign n6957 = n1043 & n6953;
  assign n6958 = n2324 & n6957;
  assign n6959 = n6956 & n6958;
  assign n6960 = n6952 & n6959;
  assign n6961 = n821 & n3001;
  assign n6962 = n6933 & n6961;
  assign n6963 = n6960 & n6962;
  assign n6964 = n5717 & n6950;
  assign n6965 = n6963 & n6964;
  assign n6966 = ~n3137 & n3896;
  assign n6967 = n564 & ~n3227;
  assign n6968 = ~n3194 & n3683;
  assign n6969 = n3468 & ~n3470;
  assign n6970 = ~n3471 & ~n6969;
  assign n6971 = n566 & n6970;
  assign n6972 = ~n6967 & ~n6968;
  assign n6973 = ~n6966 & n6972;
  assign n6974 = ~n6971 & n6973;
  assign n6975 = ~n6965 & ~n6974;
  assign n6976 = ~n218 & ~n448;
  assign n6977 = ~n141 & ~n404;
  assign n6978 = ~n466 & n6977;
  assign n6979 = n169 & n6976;
  assign n6980 = n6978 & n6979;
  assign n6981 = ~n91 & ~n319;
  assign n6982 = ~n513 & ~n642;
  assign n6983 = ~n659 & n6982;
  assign n6984 = n672 & n6981;
  assign n6985 = n1020 & n1383;
  assign n6986 = n6984 & n6985;
  assign n6987 = n2273 & n6983;
  assign n6988 = n4606 & n6987;
  assign n6989 = n6986 & n6988;
  assign n6990 = ~n162 & ~n683;
  assign n6991 = n217 & n6990;
  assign n6992 = ~n126 & ~n402;
  assign n6993 = ~n469 & ~n598;
  assign n6994 = n6992 & n6993;
  assign n6995 = n201 & n461;
  assign n6996 = n464 & n840;
  assign n6997 = n1630 & n1904;
  assign n6998 = n3404 & n4911;
  assign n6999 = n6997 & n6998;
  assign n7000 = n6995 & n6996;
  assign n7001 = n2397 & n6994;
  assign n7002 = n4165 & n6991;
  assign n7003 = n7001 & n7002;
  assign n7004 = n6999 & n7000;
  assign n7005 = n6980 & n7004;
  assign n7006 = n7003 & n7005;
  assign n7007 = n6989 & n7006;
  assign n7008 = n2941 & n7007;
  assign n7009 = n564 & ~n3319;
  assign n7010 = ~n3227 & n3683;
  assign n7011 = ~n3194 & n3896;
  assign n7012 = n3464 & ~n3466;
  assign n7013 = ~n3467 & ~n7012;
  assign n7014 = n566 & n7013;
  assign n7015 = ~n7010 & ~n7011;
  assign n7016 = ~n7009 & n7015;
  assign n7017 = ~n7014 & n7016;
  assign n7018 = ~n7008 & ~n7017;
  assign n7019 = ~n513 & n2832;
  assign n7020 = ~n182 & ~n569;
  assign n7021 = n4092 & n7020;
  assign n7022 = ~n131 & ~n148;
  assign n7023 = ~n247 & ~n701;
  assign n7024 = n7022 & n7023;
  assign n7025 = n930 & n2055;
  assign n7026 = n3351 & n7025;
  assign n7027 = n7024 & n7026;
  assign n7028 = n824 & n1148;
  assign n7029 = n1247 & n1432;
  assign n7030 = n1464 & n1754;
  assign n7031 = n2480 & n2797;
  assign n7032 = n3845 & n4104;
  assign n7033 = n7031 & n7032;
  assign n7034 = n7029 & n7030;
  assign n7035 = n7028 & n7034;
  assign n7036 = n7019 & n7033;
  assign n7037 = n7021 & n7036;
  assign n7038 = n7027 & n7035;
  assign n7039 = n7037 & n7038;
  assign n7040 = n2796 & n7039;
  assign n7041 = n4178 & n4811;
  assign n7042 = n7040 & n7041;
  assign n7043 = ~n3376 & n3683;
  assign n7044 = ~n3319 & n3896;
  assign n7045 = n564 & ~n3460;
  assign n7046 = ~n3376 & n3460;
  assign n7047 = n3319 & ~n7046;
  assign n7048 = ~n3319 & n7046;
  assign n7049 = ~n7047 & ~n7048;
  assign n7050 = n566 & n7049;
  assign n7051 = ~n7043 & ~n7045;
  assign n7052 = ~n7044 & n7051;
  assign n7053 = ~n7050 & n7052;
  assign n7054 = ~n7042 & ~n7053;
  assign n7055 = ~n290 & n3657;
  assign n7056 = ~n200 & ~n646;
  assign n7057 = ~n673 & n7056;
  assign n7058 = n930 & n2797;
  assign n7059 = n7057 & n7058;
  assign n7060 = ~n583 & n2784;
  assign n7061 = ~n165 & ~n242;
  assign n7062 = ~n311 & ~n569;
  assign n7063 = n7061 & n7062;
  assign n7064 = n737 & n741;
  assign n7065 = n925 & n7064;
  assign n7066 = n2375 & n7063;
  assign n7067 = n7065 & n7066;
  assign n7068 = ~n133 & ~n192;
  assign n7069 = n1011 & n7068;
  assign n7070 = ~n149 & ~n212;
  assign n7071 = ~n296 & ~n374;
  assign n7072 = ~n404 & ~n554;
  assign n7073 = n7071 & n7072;
  assign n7074 = n464 & n7070;
  assign n7075 = n493 & n1394;
  assign n7076 = n1632 & n1762;
  assign n7077 = n2296 & n3079;
  assign n7078 = n7076 & n7077;
  assign n7079 = n7074 & n7075;
  assign n7080 = n7069 & n7073;
  assign n7081 = n7079 & n7080;
  assign n7082 = n7060 & n7078;
  assign n7083 = n7081 & n7082;
  assign n7084 = n7067 & n7083;
  assign n7085 = ~n145 & ~n172;
  assign n7086 = ~n175 & ~n213;
  assign n7087 = n7085 & n7086;
  assign n7088 = n1172 & n3233;
  assign n7089 = n7087 & n7088;
  assign n7090 = n2028 & n3711;
  assign n7091 = n7089 & n7090;
  assign n7092 = n2364 & n7055;
  assign n7093 = n7059 & n7092;
  assign n7094 = n7091 & n7093;
  assign n7095 = n3254 & n7094;
  assign n7096 = n2217 & n7084;
  assign n7097 = n7095 & n7096;
  assign n7098 = n7054 & ~n7097;
  assign n7099 = ~n7054 & n7097;
  assign n7100 = ~n7098 & ~n7099;
  assign n7101 = ~n3319 & n3683;
  assign n7102 = n564 & ~n3376;
  assign n7103 = ~n3227 & n3896;
  assign n7104 = ~n3322 & ~n3462;
  assign n7105 = ~n3463 & ~n7104;
  assign n7106 = n566 & n7105;
  assign n7107 = ~n7102 & ~n7103;
  assign n7108 = ~n7101 & n7107;
  assign n7109 = ~n7106 & n7108;
  assign n7110 = n7100 & ~n7109;
  assign n7111 = ~n7098 & ~n7110;
  assign n7112 = n7008 & n7017;
  assign n7113 = ~n7018 & ~n7112;
  assign n7114 = ~n7111 & n7113;
  assign n7115 = ~n7018 & ~n7114;
  assign n7116 = n6965 & n6974;
  assign n7117 = ~n6975 & ~n7116;
  assign n7118 = ~n7115 & n7117;
  assign n7119 = ~n6975 & ~n7118;
  assign n7120 = n6915 & n6924;
  assign n7121 = ~n6925 & ~n7120;
  assign n7122 = ~n7119 & n7121;
  assign n7123 = ~n6925 & ~n7122;
  assign n7124 = n6868 & n6877;
  assign n7125 = ~n6878 & ~n7124;
  assign n7126 = ~n7123 & n7125;
  assign n7127 = ~n6878 & ~n7126;
  assign n7128 = ~n6491 & n6500;
  assign n7129 = ~n6501 & ~n7128;
  assign n7130 = ~n7127 & n7129;
  assign n7131 = n7127 & ~n7129;
  assign n7132 = ~n7130 & ~n7131;
  assign n7133 = ~n2866 & n3943;
  assign n7134 = ~n2726 & n4472;
  assign n7135 = ~n2781 & n4070;
  assign n7136 = n3944 & n6520;
  assign n7137 = ~n7133 & ~n7135;
  assign n7138 = ~n7134 & n7137;
  assign n7139 = ~n7136 & n7138;
  assign n7140 = pi29  & n7139;
  assign n7141 = ~pi29  & ~n7139;
  assign n7142 = ~n7140 & ~n7141;
  assign n7143 = n7132 & ~n7142;
  assign n7144 = ~n7130 & ~n7143;
  assign n7145 = ~n6826 & n6835;
  assign n7146 = ~n6836 & ~n7145;
  assign n7147 = ~n7144 & n7146;
  assign n7148 = ~n6836 & ~n7147;
  assign n7149 = ~n6814 & n6823;
  assign n7150 = ~n6824 & ~n7149;
  assign n7151 = ~n7148 & n7150;
  assign n7152 = ~n6824 & ~n7151;
  assign n7153 = ~n6515 & n6524;
  assign n7154 = ~n6525 & ~n7153;
  assign n7155 = ~n7152 & n7154;
  assign n7156 = n7152 & ~n7154;
  assign n7157 = ~n7155 & ~n7156;
  assign n7158 = ~n2538 & n4472;
  assign n7159 = ~n2622 & n4070;
  assign n7160 = ~n2657 & n3943;
  assign n7161 = n3944 & n6271;
  assign n7162 = ~n7158 & ~n7160;
  assign n7163 = ~n7159 & n7162;
  assign n7164 = ~n7161 & n7163;
  assign n7165 = pi29  & n7164;
  assign n7166 = ~pi29  & ~n7164;
  assign n7167 = ~n7165 & ~n7166;
  assign n7168 = n7157 & ~n7167;
  assign n7169 = ~n7155 & ~n7168;
  assign n7170 = ~n6531 & n6541;
  assign n7171 = ~n6542 & ~n7170;
  assign n7172 = n7169 & ~n7171;
  assign n7173 = ~n7169 & n7171;
  assign n7174 = ~n7172 & ~n7173;
  assign n7175 = ~n2356 & n4515;
  assign n7176 = ~n2265 & n4691;
  assign n7177 = ~n2165 & n4721;
  assign n7178 = n4516 & n5632;
  assign n7179 = ~n7175 & ~n7176;
  assign n7180 = ~n7177 & n7179;
  assign n7181 = ~n7178 & n7180;
  assign n7182 = pi26  & n7181;
  assign n7183 = ~pi26  & ~n7181;
  assign n7184 = ~n7182 & ~n7183;
  assign n7185 = n7174 & n7184;
  assign n7186 = ~n7172 & ~n7185;
  assign n7187 = n6812 & n7186;
  assign n7188 = ~n6812 & ~n7186;
  assign n7189 = ~n7187 & ~n7188;
  assign n7190 = ~n1997 & n5121;
  assign n7191 = ~n1893 & n5185;
  assign n7192 = ~n1805 & n5267;
  assign n7193 = n78 & n5212;
  assign n7194 = ~n7190 & ~n7191;
  assign n7195 = ~n7192 & n7194;
  assign n7196 = ~n7193 & n7195;
  assign n7197 = pi23  & n7196;
  assign n7198 = ~pi23  & ~n7196;
  assign n7199 = ~n7197 & ~n7198;
  assign n7200 = n7189 & ~n7199;
  assign n7201 = ~n7187 & ~n7200;
  assign n7202 = n6807 & ~n6809;
  assign n7203 = ~n6810 & ~n7202;
  assign n7204 = ~n7201 & n7203;
  assign n7205 = ~n6810 & ~n7204;
  assign n7206 = ~n6797 & ~n7205;
  assign n7207 = n6797 & n7205;
  assign n7208 = ~n7206 & ~n7207;
  assign n7209 = ~n1532 & n5312;
  assign n7210 = ~n1425 & n5901;
  assign n7211 = ~n1337 & n5982;
  assign n7212 = n4452 & n5306;
  assign n7213 = ~n7209 & ~n7210;
  assign n7214 = ~n7211 & n7213;
  assign n7215 = ~n7212 & n7214;
  assign n7216 = pi20  & n7215;
  assign n7217 = ~pi20  & ~n7215;
  assign n7218 = ~n7216 & ~n7217;
  assign n7219 = n7208 & ~n7218;
  assign n7220 = ~n7206 & ~n7219;
  assign n7221 = ~n6737 & n6747;
  assign n7222 = ~n6748 & ~n7221;
  assign n7223 = ~n7220 & n7222;
  assign n7224 = n7220 & ~n7222;
  assign n7225 = ~n7223 & ~n7224;
  assign n7226 = ~n898 & n6608;
  assign n7227 = ~n1006 & n6356;
  assign n7228 = ~n1107 & n6140;
  assign n7229 = n4041 & n6134;
  assign n7230 = ~n7226 & ~n7227;
  assign n7231 = ~n7228 & n7230;
  assign n7232 = ~n7229 & n7231;
  assign n7233 = pi17  & n7232;
  assign n7234 = ~pi17  & ~n7232;
  assign n7235 = ~n7233 & ~n7234;
  assign n7236 = n7225 & ~n7235;
  assign n7237 = ~n7223 & ~n7236;
  assign n7238 = n6792 & ~n6794;
  assign n7239 = ~n6795 & ~n7238;
  assign n7240 = ~n7237 & n7239;
  assign n7241 = ~n6795 & ~n7240;
  assign n7242 = ~n621 & n6653;
  assign n7243 = ~n6643 & n6651;
  assign n7244 = ~n563 & n7243;
  assign n7245 = n3687 & n6647;
  assign n7246 = ~n7242 & ~n7244;
  assign n7247 = ~n7245 & n7246;
  assign n7248 = pi14  & n7247;
  assign n7249 = ~pi14  & ~n7247;
  assign n7250 = ~n7248 & ~n7249;
  assign n7251 = ~n7241 & ~n7250;
  assign n7252 = ~n6758 & ~n6768;
  assign n7253 = ~n6769 & ~n7252;
  assign n7254 = n7241 & n7250;
  assign n7255 = ~n7251 & ~n7254;
  assign n7256 = ~n7253 & n7255;
  assign n7257 = ~n7251 & ~n7256;
  assign n7258 = ~n6773 & ~n6775;
  assign n7259 = ~n6776 & ~n7258;
  assign n7260 = ~n7257 & n7259;
  assign n7261 = n7257 & ~n7259;
  assign n7262 = ~n7260 & ~n7261;
  assign n7263 = ~n7225 & n7235;
  assign n7264 = ~n7236 & ~n7263;
  assign n7265 = n7201 & ~n7203;
  assign n7266 = ~n7204 & ~n7265;
  assign n7267 = ~n1610 & n5312;
  assign n7268 = ~n1532 & n5901;
  assign n7269 = ~n1425 & n5982;
  assign n7270 = n4642 & n5306;
  assign n7271 = ~n7267 & ~n7268;
  assign n7272 = ~n7269 & n7271;
  assign n7273 = ~n7270 & n7272;
  assign n7274 = pi20  & n7273;
  assign n7275 = ~pi20  & ~n7273;
  assign n7276 = ~n7274 & ~n7275;
  assign n7277 = n7266 & ~n7276;
  assign n7278 = ~n7189 & n7199;
  assign n7279 = ~n7200 & ~n7278;
  assign n7280 = ~n7174 & ~n7184;
  assign n7281 = ~n7185 & ~n7280;
  assign n7282 = ~n2356 & n4691;
  assign n7283 = ~n2442 & n4515;
  assign n7284 = ~n2265 & n4721;
  assign n7285 = n4516 & n5650;
  assign n7286 = ~n7283 & ~n7284;
  assign n7287 = ~n7282 & n7286;
  assign n7288 = ~n7285 & n7287;
  assign n7289 = pi26  & n7288;
  assign n7290 = ~pi26  & ~n7288;
  assign n7291 = ~n7289 & ~n7290;
  assign n7292 = ~n7157 & n7167;
  assign n7293 = ~n7168 & ~n7292;
  assign n7294 = ~n7291 & n7293;
  assign n7295 = ~n2622 & n4472;
  assign n7296 = ~n2726 & n3943;
  assign n7297 = ~n2657 & n4070;
  assign n7298 = n3944 & n6407;
  assign n7299 = ~n7295 & ~n7297;
  assign n7300 = ~n7296 & n7299;
  assign n7301 = ~n7298 & n7300;
  assign n7302 = pi29  & n7301;
  assign n7303 = ~pi29  & ~n7301;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = n7148 & ~n7150;
  assign n7306 = ~n7151 & ~n7305;
  assign n7307 = ~n7304 & n7306;
  assign n7308 = n7304 & ~n7306;
  assign n7309 = ~n7307 & ~n7308;
  assign n7310 = ~n2356 & n4721;
  assign n7311 = ~n2538 & n4515;
  assign n7312 = ~n2442 & n4691;
  assign n7313 = n4516 & n6042;
  assign n7314 = ~n7310 & ~n7312;
  assign n7315 = ~n7311 & n7314;
  assign n7316 = ~n7313 & n7315;
  assign n7317 = pi26  & n7316;
  assign n7318 = ~pi26  & ~n7316;
  assign n7319 = ~n7317 & ~n7318;
  assign n7320 = n7309 & ~n7319;
  assign n7321 = ~n7307 & ~n7320;
  assign n7322 = n7291 & ~n7293;
  assign n7323 = ~n7294 & ~n7322;
  assign n7324 = ~n7321 & n7323;
  assign n7325 = ~n7294 & ~n7324;
  assign n7326 = n7281 & n7325;
  assign n7327 = ~n7281 & ~n7325;
  assign n7328 = ~n7326 & ~n7327;
  assign n7329 = ~n2045 & n5121;
  assign n7330 = ~n1997 & n5185;
  assign n7331 = ~n1893 & n5267;
  assign n7332 = n78 & n5061;
  assign n7333 = ~n7329 & ~n7330;
  assign n7334 = ~n7331 & n7333;
  assign n7335 = ~n7332 & n7334;
  assign n7336 = pi23  & n7335;
  assign n7337 = ~pi23  & ~n7335;
  assign n7338 = ~n7336 & ~n7337;
  assign n7339 = n7328 & n7338;
  assign n7340 = ~n7326 & ~n7339;
  assign n7341 = n7279 & n7340;
  assign n7342 = ~n7279 & ~n7340;
  assign n7343 = ~n7341 & ~n7342;
  assign n7344 = ~n1737 & n5312;
  assign n7345 = ~n1610 & n5901;
  assign n7346 = ~n1532 & n5982;
  assign n7347 = n4626 & n5306;
  assign n7348 = ~n7344 & ~n7345;
  assign n7349 = ~n7346 & n7348;
  assign n7350 = ~n7347 & n7349;
  assign n7351 = pi20  & n7350;
  assign n7352 = ~pi20  & ~n7350;
  assign n7353 = ~n7351 & ~n7352;
  assign n7354 = n7343 & ~n7353;
  assign n7355 = ~n7341 & ~n7354;
  assign n7356 = ~n7266 & n7276;
  assign n7357 = ~n7277 & ~n7356;
  assign n7358 = ~n7355 & n7357;
  assign n7359 = ~n7277 & ~n7358;
  assign n7360 = ~n7208 & n7218;
  assign n7361 = ~n7219 & ~n7360;
  assign n7362 = n7359 & ~n7361;
  assign n7363 = ~n7359 & n7361;
  assign n7364 = ~n7362 & ~n7363;
  assign n7365 = ~n1107 & n6356;
  assign n7366 = ~n1006 & n6608;
  assign n7367 = ~n1230 & n6140;
  assign n7368 = n4233 & n6134;
  assign n7369 = ~n7365 & ~n7366;
  assign n7370 = ~n7367 & n7369;
  assign n7371 = ~n7368 & n7370;
  assign n7372 = pi17  & n7371;
  assign n7373 = ~pi17  & ~n7371;
  assign n7374 = ~n7372 & ~n7373;
  assign n7375 = n7364 & n7374;
  assign n7376 = ~n7362 & ~n7375;
  assign n7377 = n7264 & n7376;
  assign n7378 = ~n7264 & ~n7376;
  assign n7379 = ~n7377 & ~n7378;
  assign n7380 = n6643 & ~n6646;
  assign n7381 = ~n621 & n7380;
  assign n7382 = ~n729 & n7243;
  assign n7383 = ~n802 & n6653;
  assign n7384 = n3955 & n6647;
  assign n7385 = ~n7381 & ~n7383;
  assign n7386 = ~n7382 & n7385;
  assign n7387 = ~n7384 & n7386;
  assign n7388 = pi14  & n7387;
  assign n7389 = ~pi14  & ~n7387;
  assign n7390 = ~n7388 & ~n7389;
  assign n7391 = n7379 & ~n7390;
  assign n7392 = ~n7377 & ~n7391;
  assign n7393 = ~n729 & n6653;
  assign n7394 = ~n621 & n7243;
  assign n7395 = ~n563 & n7380;
  assign n7396 = n3921 & n6647;
  assign n7397 = ~n7394 & ~n7395;
  assign n7398 = ~n7393 & n7397;
  assign n7399 = ~n7396 & n7398;
  assign n7400 = pi14  & n7399;
  assign n7401 = ~pi14  & ~n7399;
  assign n7402 = ~n7400 & ~n7401;
  assign n7403 = ~n7392 & ~n7402;
  assign n7404 = n7237 & ~n7239;
  assign n7405 = ~n7240 & ~n7404;
  assign n7406 = n7392 & n7402;
  assign n7407 = ~n7403 & ~n7406;
  assign n7408 = n7405 & n7407;
  assign n7409 = ~n7403 & ~n7408;
  assign n7410 = n7253 & ~n7255;
  assign n7411 = ~n7256 & ~n7410;
  assign n7412 = ~n7409 & n7411;
  assign n7413 = ~n7364 & ~n7374;
  assign n7414 = ~n7375 & ~n7413;
  assign n7415 = ~n1337 & n6140;
  assign n7416 = ~n1230 & n6356;
  assign n7417 = ~n1107 & n6608;
  assign n7418 = n4251 & n6134;
  assign n7419 = ~n7415 & ~n7416;
  assign n7420 = ~n7417 & n7419;
  assign n7421 = ~n7418 & n7420;
  assign n7422 = ~pi17  & ~n7421;
  assign n7423 = pi17  & n7421;
  assign n7424 = ~n7422 & ~n7423;
  assign n7425 = n7355 & ~n7357;
  assign n7426 = ~n7358 & ~n7425;
  assign n7427 = ~n7424 & n7426;
  assign n7428 = ~n7328 & ~n7338;
  assign n7429 = ~n7339 & ~n7428;
  assign n7430 = ~n2165 & n5121;
  assign n7431 = ~n2045 & n5185;
  assign n7432 = ~n1997 & n5267;
  assign n7433 = n78 & n5424;
  assign n7434 = ~n7431 & ~n7432;
  assign n7435 = ~n7430 & n7434;
  assign n7436 = ~n7433 & n7435;
  assign n7437 = ~pi23  & ~n7436;
  assign n7438 = pi23  & n7436;
  assign n7439 = ~n7437 & ~n7438;
  assign n7440 = n7321 & ~n7323;
  assign n7441 = ~n7324 & ~n7440;
  assign n7442 = ~n7439 & n7441;
  assign n7443 = ~n2657 & n4472;
  assign n7444 = ~n2726 & n4070;
  assign n7445 = ~n2781 & n3943;
  assign n7446 = n3944 & n6251;
  assign n7447 = ~n7443 & ~n7445;
  assign n7448 = ~n7444 & n7447;
  assign n7449 = ~n7446 & n7448;
  assign n7450 = pi29  & n7449;
  assign n7451 = ~pi29  & ~n7449;
  assign n7452 = ~n7450 & ~n7451;
  assign n7453 = n7144 & ~n7146;
  assign n7454 = ~n7147 & ~n7453;
  assign n7455 = ~n7452 & n7454;
  assign n7456 = n7452 & ~n7454;
  assign n7457 = ~n7455 & ~n7456;
  assign n7458 = ~n2622 & n4515;
  assign n7459 = ~n2538 & n4691;
  assign n7460 = ~n2442 & n4721;
  assign n7461 = n4516 & n5823;
  assign n7462 = ~n7458 & ~n7460;
  assign n7463 = ~n7459 & n7462;
  assign n7464 = ~n7461 & n7463;
  assign n7465 = pi26  & n7464;
  assign n7466 = ~pi26  & ~n7464;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = n7457 & ~n7467;
  assign n7469 = ~n7455 & ~n7468;
  assign n7470 = ~n7309 & n7319;
  assign n7471 = ~n7320 & ~n7470;
  assign n7472 = ~n7469 & n7471;
  assign n7473 = n7469 & ~n7471;
  assign n7474 = ~n7472 & ~n7473;
  assign n7475 = ~n2165 & n5185;
  assign n7476 = ~n2265 & n5121;
  assign n7477 = ~n2045 & n5267;
  assign n7478 = n78 & n5408;
  assign n7479 = ~n7476 & ~n7477;
  assign n7480 = ~n7475 & n7479;
  assign n7481 = ~n7478 & n7480;
  assign n7482 = pi23  & n7481;
  assign n7483 = ~pi23  & ~n7481;
  assign n7484 = ~n7482 & ~n7483;
  assign n7485 = n7474 & ~n7484;
  assign n7486 = ~n7472 & ~n7485;
  assign n7487 = n7439 & ~n7441;
  assign n7488 = ~n7442 & ~n7487;
  assign n7489 = ~n7486 & n7488;
  assign n7490 = ~n7442 & ~n7489;
  assign n7491 = ~n7429 & ~n7490;
  assign n7492 = n7429 & n7490;
  assign n7493 = ~n7491 & ~n7492;
  assign n7494 = ~n1805 & n5312;
  assign n7495 = ~n1737 & n5901;
  assign n7496 = ~n1610 & n5982;
  assign n7497 = n4844 & n5306;
  assign n7498 = ~n7494 & ~n7495;
  assign n7499 = ~n7496 & n7498;
  assign n7500 = ~n7497 & n7499;
  assign n7501 = pi20  & n7500;
  assign n7502 = ~pi20  & ~n7500;
  assign n7503 = ~n7501 & ~n7502;
  assign n7504 = n7493 & ~n7503;
  assign n7505 = ~n7491 & ~n7504;
  assign n7506 = ~n7343 & n7353;
  assign n7507 = ~n7354 & ~n7506;
  assign n7508 = ~n7505 & n7507;
  assign n7509 = n7505 & ~n7507;
  assign n7510 = ~n7508 & ~n7509;
  assign n7511 = ~n1425 & n6140;
  assign n7512 = ~n1337 & n6356;
  assign n7513 = ~n1230 & n6608;
  assign n7514 = n4549 & n6134;
  assign n7515 = ~n7511 & ~n7512;
  assign n7516 = ~n7513 & n7515;
  assign n7517 = ~n7514 & n7516;
  assign n7518 = pi17  & n7517;
  assign n7519 = ~pi17  & ~n7517;
  assign n7520 = ~n7518 & ~n7519;
  assign n7521 = n7510 & ~n7520;
  assign n7522 = ~n7508 & ~n7521;
  assign n7523 = n7424 & ~n7426;
  assign n7524 = ~n7427 & ~n7523;
  assign n7525 = ~n7522 & n7524;
  assign n7526 = ~n7427 & ~n7525;
  assign n7527 = ~n7414 & ~n7526;
  assign n7528 = n7414 & n7526;
  assign n7529 = ~n7527 & ~n7528;
  assign n7530 = ~n729 & n7380;
  assign n7531 = ~n802 & n7243;
  assign n7532 = ~n898 & n6653;
  assign n7533 = n3901 & n6647;
  assign n7534 = ~n7531 & ~n7532;
  assign n7535 = ~n7530 & n7534;
  assign n7536 = ~n7533 & n7535;
  assign n7537 = pi14  & n7536;
  assign n7538 = ~pi14  & ~n7536;
  assign n7539 = ~n7537 & ~n7538;
  assign n7540 = n7529 & ~n7539;
  assign n7541 = ~n7527 & ~n7540;
  assign n7542 = ~pi10  & ~pi11 ;
  assign n7543 = pi10  & pi11 ;
  assign n7544 = ~n7542 & ~n7543;
  assign n7545 = ~pi8  & ~pi9 ;
  assign n7546 = pi8  & pi9 ;
  assign n7547 = ~n7545 & ~n7546;
  assign n7548 = n7544 & n7547;
  assign n7549 = ~n3593 & n7548;
  assign n7550 = ~pi9  & ~pi10 ;
  assign n7551 = pi9  & pi10 ;
  assign n7552 = ~n7550 & ~n7551;
  assign n7553 = n7544 & ~n7547;
  assign n7554 = ~n7552 & n7553;
  assign n7555 = ~n7549 & ~n7554;
  assign n7556 = ~n563 & ~n7555;
  assign n7557 = pi11  & ~n7556;
  assign n7558 = ~pi11  & n7556;
  assign n7559 = ~n7557 & ~n7558;
  assign n7560 = ~n7541 & ~n7559;
  assign n7561 = n7541 & n7559;
  assign n7562 = ~n7560 & ~n7561;
  assign n7563 = ~n7379 & n7390;
  assign n7564 = ~n7391 & ~n7563;
  assign n7565 = n7562 & n7564;
  assign n7566 = ~n7560 & ~n7565;
  assign n7567 = ~n7405 & ~n7407;
  assign n7568 = ~n7408 & ~n7567;
  assign n7569 = ~n7566 & n7568;
  assign n7570 = n7522 & ~n7524;
  assign n7571 = ~n7525 & ~n7570;
  assign n7572 = ~n802 & n7380;
  assign n7573 = ~n898 & n7243;
  assign n7574 = ~n1006 & n6653;
  assign n7575 = n4057 & n6647;
  assign n7576 = ~n7572 & ~n7573;
  assign n7577 = ~n7574 & n7576;
  assign n7578 = ~n7575 & n7577;
  assign n7579 = pi14  & n7578;
  assign n7580 = ~pi14  & ~n7578;
  assign n7581 = ~n7579 & ~n7580;
  assign n7582 = n7571 & ~n7581;
  assign n7583 = ~n7510 & n7520;
  assign n7584 = ~n7521 & ~n7583;
  assign n7585 = n7486 & ~n7488;
  assign n7586 = ~n7489 & ~n7585;
  assign n7587 = ~n1893 & n5312;
  assign n7588 = ~n1805 & n5901;
  assign n7589 = ~n1737 & n5982;
  assign n7590 = n4862 & n5306;
  assign n7591 = ~n7587 & ~n7588;
  assign n7592 = ~n7589 & n7591;
  assign n7593 = ~n7590 & n7592;
  assign n7594 = pi20  & n7593;
  assign n7595 = ~pi20  & ~n7593;
  assign n7596 = ~n7594 & ~n7595;
  assign n7597 = n7586 & ~n7596;
  assign n7598 = ~n2866 & n4070;
  assign n7599 = ~n2781 & n4472;
  assign n7600 = ~n2901 & n3943;
  assign n7601 = n3944 & n6819;
  assign n7602 = ~n7598 & ~n7599;
  assign n7603 = ~n7600 & n7602;
  assign n7604 = ~n7601 & n7603;
  assign n7605 = pi29  & n7604;
  assign n7606 = ~pi29  & ~n7604;
  assign n7607 = ~n7605 & ~n7606;
  assign n7608 = n7123 & ~n7125;
  assign n7609 = ~n7126 & ~n7608;
  assign n7610 = ~n7607 & n7609;
  assign n7611 = ~n2866 & n4472;
  assign n7612 = ~n2978 & n3943;
  assign n7613 = ~n2901 & n4070;
  assign n7614 = n3944 & n6831;
  assign n7615 = ~n7611 & ~n7613;
  assign n7616 = ~n7612 & n7615;
  assign n7617 = ~n7614 & n7616;
  assign n7618 = pi29  & n7617;
  assign n7619 = ~pi29  & ~n7617;
  assign n7620 = ~n7618 & ~n7619;
  assign n7621 = n7119 & ~n7121;
  assign n7622 = ~n7122 & ~n7621;
  assign n7623 = ~n7620 & n7622;
  assign n7624 = ~n2901 & n4472;
  assign n7625 = ~n2978 & n4070;
  assign n7626 = ~n3069 & n3943;
  assign n7627 = n3944 & n6496;
  assign n7628 = ~n7624 & ~n7626;
  assign n7629 = ~n7625 & n7628;
  assign n7630 = ~n7627 & n7629;
  assign n7631 = ~pi29  & ~n7630;
  assign n7632 = pi29  & n7630;
  assign n7633 = ~n7631 & ~n7632;
  assign n7634 = n7115 & ~n7117;
  assign n7635 = ~n7118 & ~n7634;
  assign n7636 = ~n7633 & n7635;
  assign n7637 = ~n2978 & n4472;
  assign n7638 = ~n3137 & n3943;
  assign n7639 = ~n3069 & n4070;
  assign n7640 = n3944 & n6873;
  assign n7641 = ~n7637 & ~n7639;
  assign n7642 = ~n7638 & n7641;
  assign n7643 = ~n7640 & n7642;
  assign n7644 = ~pi29  & ~n7643;
  assign n7645 = pi29  & n7643;
  assign n7646 = ~n7644 & ~n7645;
  assign n7647 = n7111 & ~n7113;
  assign n7648 = ~n7114 & ~n7647;
  assign n7649 = ~n7646 & n7648;
  assign n7650 = ~n3069 & n4472;
  assign n7651 = ~n3137 & n4070;
  assign n7652 = ~n3194 & n3943;
  assign n7653 = n3944 & n6920;
  assign n7654 = ~n7650 & ~n7652;
  assign n7655 = ~n7651 & n7654;
  assign n7656 = ~n7653 & n7655;
  assign n7657 = ~pi29  & ~n7656;
  assign n7658 = pi29  & n7656;
  assign n7659 = ~n7657 & ~n7658;
  assign n7660 = ~n7100 & n7109;
  assign n7661 = ~n7110 & ~n7660;
  assign n7662 = ~n7659 & n7661;
  assign n7663 = ~n3137 & n4472;
  assign n7664 = ~n3194 & n4070;
  assign n7665 = ~n3227 & n3943;
  assign n7666 = n3944 & n6970;
  assign n7667 = ~n7664 & ~n7665;
  assign n7668 = ~n7663 & n7667;
  assign n7669 = ~n7666 & n7668;
  assign n7670 = ~pi29  & ~n7669;
  assign n7671 = pi29  & n7669;
  assign n7672 = ~n7670 & ~n7671;
  assign n7673 = n7042 & n7053;
  assign n7674 = ~n7054 & ~n7673;
  assign n7675 = ~n7672 & n7674;
  assign n7676 = ~n3319 & n3943;
  assign n7677 = ~n3227 & n4070;
  assign n7678 = ~n3194 & n4472;
  assign n7679 = n3944 & n7013;
  assign n7680 = ~n7677 & ~n7678;
  assign n7681 = ~n7676 & n7680;
  assign n7682 = ~n7679 & n7681;
  assign n7683 = ~pi29  & ~n7682;
  assign n7684 = pi29  & n7682;
  assign n7685 = ~n7683 & ~n7684;
  assign n7686 = ~n3376 & n3896;
  assign n7687 = ~n3460 & n3683;
  assign n7688 = n3376 & ~n3460;
  assign n7689 = ~n7046 & ~n7688;
  assign n7690 = n566 & ~n7689;
  assign n7691 = ~n7686 & ~n7687;
  assign n7692 = ~n7690 & n7691;
  assign n7693 = ~n7685 & ~n7692;
  assign n7694 = ~n565 & ~n3460;
  assign n7695 = ~n3460 & n3941;
  assign n7696 = pi29  & n7695;
  assign n7697 = ~n3376 & n4472;
  assign n7698 = ~n3460 & n4070;
  assign n7699 = n3944 & ~n7689;
  assign n7700 = ~n7697 & ~n7698;
  assign n7701 = ~n7699 & n7700;
  assign n7702 = ~n7696 & n7701;
  assign n7703 = ~n3460 & n3943;
  assign n7704 = ~n3319 & n4472;
  assign n7705 = ~n3376 & n4070;
  assign n7706 = n3944 & n7049;
  assign n7707 = ~n7703 & ~n7705;
  assign n7708 = ~n7704 & n7707;
  assign n7709 = ~n7706 & n7708;
  assign n7710 = pi29  & n7702;
  assign n7711 = n7709 & n7710;
  assign n7712 = n7694 & n7711;
  assign n7713 = ~n3319 & n4070;
  assign n7714 = ~n3376 & n3943;
  assign n7715 = ~n3227 & n4472;
  assign n7716 = n3944 & n7105;
  assign n7717 = ~n7714 & ~n7715;
  assign n7718 = ~n7713 & n7717;
  assign n7719 = ~n7716 & n7718;
  assign n7720 = ~pi29  & ~n7719;
  assign n7721 = pi29  & n7719;
  assign n7722 = ~n7720 & ~n7721;
  assign n7723 = ~n7694 & ~n7711;
  assign n7724 = ~n7712 & ~n7723;
  assign n7725 = ~n7722 & n7724;
  assign n7726 = ~n7712 & ~n7725;
  assign n7727 = n7685 & n7692;
  assign n7728 = ~n7693 & ~n7727;
  assign n7729 = ~n7726 & n7728;
  assign n7730 = ~n7693 & ~n7729;
  assign n7731 = n7672 & ~n7674;
  assign n7732 = ~n7675 & ~n7731;
  assign n7733 = ~n7730 & n7732;
  assign n7734 = ~n7675 & ~n7733;
  assign n7735 = n7659 & ~n7661;
  assign n7736 = ~n7662 & ~n7735;
  assign n7737 = ~n7734 & n7736;
  assign n7738 = ~n7662 & ~n7737;
  assign n7739 = n7646 & ~n7648;
  assign n7740 = ~n7649 & ~n7739;
  assign n7741 = ~n7738 & n7740;
  assign n7742 = ~n7649 & ~n7741;
  assign n7743 = n7633 & ~n7635;
  assign n7744 = ~n7636 & ~n7743;
  assign n7745 = ~n7742 & n7744;
  assign n7746 = ~n7636 & ~n7745;
  assign n7747 = n7620 & ~n7622;
  assign n7748 = ~n7623 & ~n7747;
  assign n7749 = ~n7746 & n7748;
  assign n7750 = ~n7623 & ~n7749;
  assign n7751 = n7607 & ~n7609;
  assign n7752 = ~n7610 & ~n7751;
  assign n7753 = ~n7750 & n7752;
  assign n7754 = ~n7610 & ~n7753;
  assign n7755 = ~n7132 & n7142;
  assign n7756 = ~n7143 & ~n7755;
  assign n7757 = ~n7754 & n7756;
  assign n7758 = ~n2538 & n4721;
  assign n7759 = ~n2622 & n4691;
  assign n7760 = ~n2657 & n4515;
  assign n7761 = n4516 & n6271;
  assign n7762 = ~n7758 & ~n7760;
  assign n7763 = ~n7759 & n7762;
  assign n7764 = ~n7761 & n7763;
  assign n7765 = ~pi26  & ~n7764;
  assign n7766 = pi26  & n7764;
  assign n7767 = ~n7765 & ~n7766;
  assign n7768 = n7754 & ~n7756;
  assign n7769 = ~n7757 & ~n7768;
  assign n7770 = ~n7767 & n7769;
  assign n7771 = ~n7757 & ~n7770;
  assign n7772 = ~n7457 & n7467;
  assign n7773 = ~n7468 & ~n7772;
  assign n7774 = ~n7771 & n7773;
  assign n7775 = n7771 & ~n7773;
  assign n7776 = ~n7774 & ~n7775;
  assign n7777 = ~n2356 & n5121;
  assign n7778 = ~n2265 & n5185;
  assign n7779 = ~n2165 & n5267;
  assign n7780 = n78 & n5632;
  assign n7781 = ~n7777 & ~n7778;
  assign n7782 = ~n7779 & n7781;
  assign n7783 = ~n7780 & n7782;
  assign n7784 = pi23  & n7783;
  assign n7785 = ~pi23  & ~n7783;
  assign n7786 = ~n7784 & ~n7785;
  assign n7787 = n7776 & ~n7786;
  assign n7788 = ~n7774 & ~n7787;
  assign n7789 = ~n7474 & n7484;
  assign n7790 = ~n7485 & ~n7789;
  assign n7791 = ~n7788 & n7790;
  assign n7792 = n7788 & ~n7790;
  assign n7793 = ~n7791 & ~n7792;
  assign n7794 = ~n1997 & n5312;
  assign n7795 = ~n1893 & n5901;
  assign n7796 = ~n1805 & n5982;
  assign n7797 = n5212 & n5306;
  assign n7798 = ~n7794 & ~n7795;
  assign n7799 = ~n7796 & n7798;
  assign n7800 = ~n7797 & n7799;
  assign n7801 = pi20  & n7800;
  assign n7802 = ~pi20  & ~n7800;
  assign n7803 = ~n7801 & ~n7802;
  assign n7804 = n7793 & ~n7803;
  assign n7805 = ~n7791 & ~n7804;
  assign n7806 = ~n7586 & n7596;
  assign n7807 = ~n7597 & ~n7806;
  assign n7808 = ~n7805 & n7807;
  assign n7809 = ~n7597 & ~n7808;
  assign n7810 = ~n7493 & n7503;
  assign n7811 = ~n7504 & ~n7810;
  assign n7812 = n7809 & ~n7811;
  assign n7813 = ~n7809 & n7811;
  assign n7814 = ~n7812 & ~n7813;
  assign n7815 = ~n1532 & n6140;
  assign n7816 = ~n1425 & n6356;
  assign n7817 = ~n1337 & n6608;
  assign n7818 = n4452 & n6134;
  assign n7819 = ~n7815 & ~n7816;
  assign n7820 = ~n7817 & n7819;
  assign n7821 = ~n7818 & n7820;
  assign n7822 = pi17  & n7821;
  assign n7823 = ~pi17  & ~n7821;
  assign n7824 = ~n7822 & ~n7823;
  assign n7825 = n7814 & n7824;
  assign n7826 = ~n7812 & ~n7825;
  assign n7827 = n7584 & n7826;
  assign n7828 = ~n7584 & ~n7826;
  assign n7829 = ~n7827 & ~n7828;
  assign n7830 = ~n898 & n7380;
  assign n7831 = ~n1006 & n7243;
  assign n7832 = ~n1107 & n6653;
  assign n7833 = n4041 & n6647;
  assign n7834 = ~n7830 & ~n7831;
  assign n7835 = ~n7832 & n7834;
  assign n7836 = ~n7833 & n7835;
  assign n7837 = pi14  & n7836;
  assign n7838 = ~pi14  & ~n7836;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = n7829 & ~n7839;
  assign n7841 = ~n7827 & ~n7840;
  assign n7842 = ~n7571 & n7581;
  assign n7843 = ~n7582 & ~n7842;
  assign n7844 = ~n7841 & n7843;
  assign n7845 = ~n7582 & ~n7844;
  assign n7846 = ~n621 & n7554;
  assign n7847 = ~n7547 & n7552;
  assign n7848 = ~n563 & n7847;
  assign n7849 = n3687 & n7548;
  assign n7850 = ~n7846 & ~n7848;
  assign n7851 = ~n7849 & n7850;
  assign n7852 = pi11  & n7851;
  assign n7853 = ~pi11  & ~n7851;
  assign n7854 = ~n7852 & ~n7853;
  assign n7855 = ~n7845 & ~n7854;
  assign n7856 = n7845 & n7854;
  assign n7857 = ~n7855 & ~n7856;
  assign n7858 = ~n7529 & n7539;
  assign n7859 = ~n7540 & ~n7858;
  assign n7860 = n7857 & n7859;
  assign n7861 = ~n7855 & ~n7860;
  assign n7862 = ~n7562 & ~n7564;
  assign n7863 = ~n7565 & ~n7862;
  assign n7864 = ~n7861 & n7863;
  assign n7865 = n7861 & ~n7863;
  assign n7866 = ~n7864 & ~n7865;
  assign n7867 = ~n7814 & ~n7824;
  assign n7868 = ~n7825 & ~n7867;
  assign n7869 = ~n1610 & n6140;
  assign n7870 = ~n1532 & n6356;
  assign n7871 = ~n1425 & n6608;
  assign n7872 = n4642 & n6134;
  assign n7873 = ~n7869 & ~n7870;
  assign n7874 = ~n7871 & n7873;
  assign n7875 = ~n7872 & n7874;
  assign n7876 = ~pi17  & ~n7875;
  assign n7877 = pi17  & n7875;
  assign n7878 = ~n7876 & ~n7877;
  assign n7879 = n7805 & ~n7807;
  assign n7880 = ~n7808 & ~n7879;
  assign n7881 = ~n7878 & n7880;
  assign n7882 = n7750 & ~n7752;
  assign n7883 = ~n7753 & ~n7882;
  assign n7884 = ~n2622 & n4721;
  assign n7885 = ~n2726 & n4515;
  assign n7886 = ~n2657 & n4691;
  assign n7887 = n4516 & n6407;
  assign n7888 = ~n7884 & ~n7886;
  assign n7889 = ~n7885 & n7888;
  assign n7890 = ~n7887 & n7889;
  assign n7891 = pi26  & n7890;
  assign n7892 = ~pi26  & ~n7890;
  assign n7893 = ~n7891 & ~n7892;
  assign n7894 = n7883 & ~n7893;
  assign n7895 = n7746 & ~n7748;
  assign n7896 = ~n7749 & ~n7895;
  assign n7897 = ~n2657 & n4721;
  assign n7898 = ~n2726 & n4691;
  assign n7899 = ~n2781 & n4515;
  assign n7900 = n4516 & n6251;
  assign n7901 = ~n7897 & ~n7899;
  assign n7902 = ~n7898 & n7901;
  assign n7903 = ~n7900 & n7902;
  assign n7904 = pi26  & n7903;
  assign n7905 = ~pi26  & ~n7903;
  assign n7906 = ~n7904 & ~n7905;
  assign n7907 = n7896 & ~n7906;
  assign n7908 = n7742 & ~n7744;
  assign n7909 = ~n7745 & ~n7908;
  assign n7910 = ~n2866 & n4515;
  assign n7911 = ~n2726 & n4721;
  assign n7912 = ~n2781 & n4691;
  assign n7913 = n4516 & n6520;
  assign n7914 = ~n7910 & ~n7912;
  assign n7915 = ~n7911 & n7914;
  assign n7916 = ~n7913 & n7915;
  assign n7917 = pi26  & n7916;
  assign n7918 = ~pi26  & ~n7916;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = n7909 & ~n7919;
  assign n7921 = n7738 & ~n7740;
  assign n7922 = ~n7741 & ~n7921;
  assign n7923 = ~n2866 & n4691;
  assign n7924 = ~n2781 & n4721;
  assign n7925 = ~n2901 & n4515;
  assign n7926 = n4516 & n6819;
  assign n7927 = ~n7923 & ~n7924;
  assign n7928 = ~n7925 & n7927;
  assign n7929 = ~n7926 & n7928;
  assign n7930 = pi26  & n7929;
  assign n7931 = ~pi26  & ~n7929;
  assign n7932 = ~n7930 & ~n7931;
  assign n7933 = n7922 & ~n7932;
  assign n7934 = n7734 & ~n7736;
  assign n7935 = ~n7737 & ~n7934;
  assign n7936 = ~n2866 & n4721;
  assign n7937 = ~n2978 & n4515;
  assign n7938 = ~n2901 & n4691;
  assign n7939 = n4516 & n6831;
  assign n7940 = ~n7936 & ~n7938;
  assign n7941 = ~n7937 & n7940;
  assign n7942 = ~n7939 & n7941;
  assign n7943 = pi26  & n7942;
  assign n7944 = ~pi26  & ~n7942;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = n7935 & ~n7945;
  assign n7947 = n7730 & ~n7732;
  assign n7948 = ~n7733 & ~n7947;
  assign n7949 = ~n2901 & n4721;
  assign n7950 = ~n2978 & n4691;
  assign n7951 = ~n3069 & n4515;
  assign n7952 = n4516 & n6496;
  assign n7953 = ~n7949 & ~n7951;
  assign n7954 = ~n7950 & n7953;
  assign n7955 = ~n7952 & n7954;
  assign n7956 = pi26  & n7955;
  assign n7957 = ~pi26  & ~n7955;
  assign n7958 = ~n7956 & ~n7957;
  assign n7959 = n7948 & ~n7958;
  assign n7960 = ~n2978 & n4721;
  assign n7961 = ~n3137 & n4515;
  assign n7962 = ~n3069 & n4691;
  assign n7963 = n4516 & n6873;
  assign n7964 = ~n7960 & ~n7962;
  assign n7965 = ~n7961 & n7964;
  assign n7966 = ~n7963 & n7965;
  assign n7967 = pi26  & n7966;
  assign n7968 = ~pi26  & ~n7966;
  assign n7969 = ~n7967 & ~n7968;
  assign n7970 = n7726 & ~n7728;
  assign n7971 = ~n7729 & ~n7970;
  assign n7972 = ~n7969 & n7971;
  assign n7973 = ~n3069 & n4721;
  assign n7974 = ~n3137 & n4691;
  assign n7975 = ~n3194 & n4515;
  assign n7976 = n4516 & n6920;
  assign n7977 = ~n7973 & ~n7975;
  assign n7978 = ~n7974 & n7977;
  assign n7979 = ~n7976 & n7978;
  assign n7980 = ~pi26  & ~n7979;
  assign n7981 = pi26  & n7979;
  assign n7982 = ~n7980 & ~n7981;
  assign n7983 = n7722 & ~n7724;
  assign n7984 = ~n7725 & ~n7983;
  assign n7985 = ~n7982 & n7984;
  assign n7986 = ~n3137 & n4721;
  assign n7987 = ~n3194 & n4691;
  assign n7988 = ~n3227 & n4515;
  assign n7989 = n4516 & n6970;
  assign n7990 = ~n7987 & ~n7988;
  assign n7991 = ~n7986 & n7990;
  assign n7992 = ~n7989 & n7991;
  assign n7993 = ~pi26  & ~n7992;
  assign n7994 = pi26  & n7992;
  assign n7995 = ~n7993 & ~n7994;
  assign n7996 = pi29  & ~n7702;
  assign n7997 = n7709 & ~n7996;
  assign n7998 = ~n7709 & n7996;
  assign n7999 = ~n7997 & ~n7998;
  assign n8000 = ~n7995 & n7999;
  assign n8001 = ~n3319 & n4515;
  assign n8002 = ~n3227 & n4691;
  assign n8003 = ~n3194 & n4721;
  assign n8004 = n4516 & n7013;
  assign n8005 = ~n8002 & ~n8003;
  assign n8006 = ~n8001 & n8005;
  assign n8007 = ~n8004 & n8006;
  assign n8008 = pi26  & n8007;
  assign n8009 = ~pi26  & ~n8007;
  assign n8010 = ~n8008 & ~n8009;
  assign n8011 = n7696 & ~n7701;
  assign n8012 = ~n7702 & ~n8011;
  assign n8013 = ~n8010 & n8012;
  assign n8014 = ~n3460 & ~n4512;
  assign n8015 = pi26  & n8014;
  assign n8016 = ~n3376 & n4721;
  assign n8017 = ~n3460 & n4691;
  assign n8018 = n4516 & ~n7689;
  assign n8019 = ~n8016 & ~n8017;
  assign n8020 = ~n8018 & n8019;
  assign n8021 = ~n8015 & n8020;
  assign n8022 = ~n3460 & n4515;
  assign n8023 = ~n3319 & n4721;
  assign n8024 = ~n3376 & n4691;
  assign n8025 = n4516 & n7049;
  assign n8026 = ~n8022 & ~n8024;
  assign n8027 = ~n8023 & n8026;
  assign n8028 = ~n8025 & n8027;
  assign n8029 = pi26  & n8021;
  assign n8030 = n8028 & n8029;
  assign n8031 = n7695 & n8030;
  assign n8032 = ~n3319 & n4691;
  assign n8033 = ~n3376 & n4515;
  assign n8034 = ~n3227 & n4721;
  assign n8035 = n4516 & n7105;
  assign n8036 = ~n8033 & ~n8034;
  assign n8037 = ~n8032 & n8036;
  assign n8038 = ~n8035 & n8037;
  assign n8039 = pi26  & n8038;
  assign n8040 = ~pi26  & ~n8038;
  assign n8041 = ~n8039 & ~n8040;
  assign n8042 = ~n7695 & ~n8030;
  assign n8043 = ~n8031 & ~n8042;
  assign n8044 = ~n8041 & n8043;
  assign n8045 = ~n8031 & ~n8044;
  assign n8046 = n8010 & ~n8012;
  assign n8047 = ~n8013 & ~n8046;
  assign n8048 = ~n8045 & n8047;
  assign n8049 = ~n8013 & ~n8048;
  assign n8050 = n7995 & ~n7999;
  assign n8051 = ~n8000 & ~n8050;
  assign n8052 = ~n8049 & n8051;
  assign n8053 = ~n8000 & ~n8052;
  assign n8054 = n7982 & ~n7984;
  assign n8055 = ~n7985 & ~n8054;
  assign n8056 = ~n8053 & n8055;
  assign n8057 = ~n7985 & ~n8056;
  assign n8058 = n7969 & ~n7971;
  assign n8059 = ~n7972 & ~n8058;
  assign n8060 = ~n8057 & n8059;
  assign n8061 = ~n7972 & ~n8060;
  assign n8062 = ~n7948 & n7958;
  assign n8063 = ~n7959 & ~n8062;
  assign n8064 = ~n8061 & n8063;
  assign n8065 = ~n7959 & ~n8064;
  assign n8066 = ~n7935 & n7945;
  assign n8067 = ~n7946 & ~n8066;
  assign n8068 = ~n8065 & n8067;
  assign n8069 = ~n7946 & ~n8068;
  assign n8070 = ~n7922 & n7932;
  assign n8071 = ~n7933 & ~n8070;
  assign n8072 = ~n8069 & n8071;
  assign n8073 = ~n7933 & ~n8072;
  assign n8074 = ~n7909 & n7919;
  assign n8075 = ~n7920 & ~n8074;
  assign n8076 = ~n8073 & n8075;
  assign n8077 = ~n7920 & ~n8076;
  assign n8078 = ~n7896 & n7906;
  assign n8079 = ~n7907 & ~n8078;
  assign n8080 = ~n8077 & n8079;
  assign n8081 = ~n7907 & ~n8080;
  assign n8082 = ~n7883 & n7893;
  assign n8083 = ~n7894 & ~n8082;
  assign n8084 = ~n8081 & n8083;
  assign n8085 = ~n7894 & ~n8084;
  assign n8086 = n7767 & ~n7769;
  assign n8087 = ~n7770 & ~n8086;
  assign n8088 = ~n8085 & n8087;
  assign n8089 = ~n2356 & n5185;
  assign n8090 = ~n2442 & n5121;
  assign n8091 = ~n2265 & n5267;
  assign n8092 = n78 & n5650;
  assign n8093 = ~n8090 & ~n8091;
  assign n8094 = ~n8089 & n8093;
  assign n8095 = ~n8092 & n8094;
  assign n8096 = ~pi23  & ~n8095;
  assign n8097 = pi23  & n8095;
  assign n8098 = ~n8096 & ~n8097;
  assign n8099 = n8085 & ~n8087;
  assign n8100 = ~n8088 & ~n8099;
  assign n8101 = ~n8098 & n8100;
  assign n8102 = ~n8088 & ~n8101;
  assign n8103 = ~n7776 & n7786;
  assign n8104 = ~n7787 & ~n8103;
  assign n8105 = ~n8102 & n8104;
  assign n8106 = n8102 & ~n8104;
  assign n8107 = ~n8105 & ~n8106;
  assign n8108 = ~n2045 & n5312;
  assign n8109 = ~n1997 & n5901;
  assign n8110 = ~n1893 & n5982;
  assign n8111 = n5061 & n5306;
  assign n8112 = ~n8108 & ~n8109;
  assign n8113 = ~n8110 & n8112;
  assign n8114 = ~n8111 & n8113;
  assign n8115 = pi20  & n8114;
  assign n8116 = ~pi20  & ~n8114;
  assign n8117 = ~n8115 & ~n8116;
  assign n8118 = n8107 & ~n8117;
  assign n8119 = ~n8105 & ~n8118;
  assign n8120 = ~n7793 & n7803;
  assign n8121 = ~n7804 & ~n8120;
  assign n8122 = ~n8119 & n8121;
  assign n8123 = n8119 & ~n8121;
  assign n8124 = ~n8122 & ~n8123;
  assign n8125 = ~n1737 & n6140;
  assign n8126 = ~n1610 & n6356;
  assign n8127 = ~n1532 & n6608;
  assign n8128 = n4626 & n6134;
  assign n8129 = ~n8125 & ~n8126;
  assign n8130 = ~n8127 & n8129;
  assign n8131 = ~n8128 & n8130;
  assign n8132 = pi17  & n8131;
  assign n8133 = ~pi17  & ~n8131;
  assign n8134 = ~n8132 & ~n8133;
  assign n8135 = n8124 & ~n8134;
  assign n8136 = ~n8122 & ~n8135;
  assign n8137 = n7878 & ~n7880;
  assign n8138 = ~n7881 & ~n8137;
  assign n8139 = ~n8136 & n8138;
  assign n8140 = ~n7881 & ~n8139;
  assign n8141 = ~n7868 & ~n8140;
  assign n8142 = n7868 & n8140;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = ~n1107 & n7243;
  assign n8145 = ~n1006 & n7380;
  assign n8146 = ~n1230 & n6653;
  assign n8147 = n4233 & n6647;
  assign n8148 = ~n8144 & ~n8145;
  assign n8149 = ~n8146 & n8148;
  assign n8150 = ~n8147 & n8149;
  assign n8151 = pi14  & n8150;
  assign n8152 = ~pi14  & ~n8150;
  assign n8153 = ~n8151 & ~n8152;
  assign n8154 = n8143 & ~n8153;
  assign n8155 = ~n8141 & ~n8154;
  assign n8156 = ~n7829 & n7839;
  assign n8157 = ~n7840 & ~n8156;
  assign n8158 = ~n8155 & n8157;
  assign n8159 = n8155 & ~n8157;
  assign n8160 = ~n8158 & ~n8159;
  assign n8161 = ~n7544 & n7547;
  assign n8162 = ~n621 & n8161;
  assign n8163 = ~n729 & n7847;
  assign n8164 = ~n802 & n7554;
  assign n8165 = n3955 & n7548;
  assign n8166 = ~n8162 & ~n8164;
  assign n8167 = ~n8163 & n8166;
  assign n8168 = ~n8165 & n8167;
  assign n8169 = pi11  & n8168;
  assign n8170 = ~pi11  & ~n8168;
  assign n8171 = ~n8169 & ~n8170;
  assign n8172 = n8160 & ~n8171;
  assign n8173 = ~n8158 & ~n8172;
  assign n8174 = ~n729 & n7554;
  assign n8175 = ~n621 & n7847;
  assign n8176 = ~n563 & n8161;
  assign n8177 = n3921 & n7548;
  assign n8178 = ~n8175 & ~n8176;
  assign n8179 = ~n8174 & n8178;
  assign n8180 = ~n8177 & n8179;
  assign n8181 = pi11  & n8180;
  assign n8182 = ~pi11  & ~n8180;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = ~n8173 & ~n8183;
  assign n8185 = n8173 & n8183;
  assign n8186 = ~n8184 & ~n8185;
  assign n8187 = n7841 & ~n7843;
  assign n8188 = ~n7844 & ~n8187;
  assign n8189 = n8186 & n8188;
  assign n8190 = ~n8184 & ~n8189;
  assign n8191 = ~n7857 & ~n7859;
  assign n8192 = ~n7860 & ~n8191;
  assign n8193 = ~n8190 & n8192;
  assign n8194 = ~pi7  & ~pi8 ;
  assign n8195 = pi7  & pi8 ;
  assign n8196 = ~n8194 & ~n8195;
  assign n8197 = ~pi5  & ~pi6 ;
  assign n8198 = pi5  & pi6 ;
  assign n8199 = ~n8197 & ~n8198;
  assign n8200 = n8196 & n8199;
  assign n8201 = ~n3593 & n8200;
  assign n8202 = ~pi6  & ~pi7 ;
  assign n8203 = pi6  & pi7 ;
  assign n8204 = ~n8202 & ~n8203;
  assign n8205 = n8196 & ~n8199;
  assign n8206 = ~n8204 & n8205;
  assign n8207 = ~n8201 & ~n8206;
  assign n8208 = ~n563 & ~n8207;
  assign n8209 = pi8  & ~n8208;
  assign n8210 = ~pi8  & n8208;
  assign n8211 = ~n8209 & ~n8210;
  assign n8212 = n8136 & ~n8138;
  assign n8213 = ~n8139 & ~n8212;
  assign n8214 = ~n1337 & n6653;
  assign n8215 = ~n1230 & n7243;
  assign n8216 = ~n1107 & n7380;
  assign n8217 = n4251 & n6647;
  assign n8218 = ~n8214 & ~n8215;
  assign n8219 = ~n8216 & n8218;
  assign n8220 = ~n8217 & n8219;
  assign n8221 = pi14  & n8220;
  assign n8222 = ~pi14  & ~n8220;
  assign n8223 = ~n8221 & ~n8222;
  assign n8224 = n8213 & ~n8223;
  assign n8225 = ~n2356 & n5267;
  assign n8226 = ~n2538 & n5121;
  assign n8227 = ~n2442 & n5185;
  assign n8228 = n78 & n6042;
  assign n8229 = ~n8225 & ~n8227;
  assign n8230 = ~n8226 & n8229;
  assign n8231 = ~n8228 & n8230;
  assign n8232 = ~pi23  & ~n8231;
  assign n8233 = pi23  & n8231;
  assign n8234 = ~n8232 & ~n8233;
  assign n8235 = n8081 & ~n8083;
  assign n8236 = ~n8084 & ~n8235;
  assign n8237 = ~n8234 & n8236;
  assign n8238 = ~n2622 & n5121;
  assign n8239 = ~n2538 & n5185;
  assign n8240 = ~n2442 & n5267;
  assign n8241 = n78 & n5823;
  assign n8242 = ~n8238 & ~n8240;
  assign n8243 = ~n8239 & n8242;
  assign n8244 = ~n8241 & n8243;
  assign n8245 = ~pi23  & ~n8244;
  assign n8246 = pi23  & n8244;
  assign n8247 = ~n8245 & ~n8246;
  assign n8248 = n8077 & ~n8079;
  assign n8249 = ~n8080 & ~n8248;
  assign n8250 = ~n8247 & n8249;
  assign n8251 = ~n2538 & n5267;
  assign n8252 = ~n2622 & n5185;
  assign n8253 = ~n2657 & n5121;
  assign n8254 = n78 & n6271;
  assign n8255 = ~n8251 & ~n8253;
  assign n8256 = ~n8252 & n8255;
  assign n8257 = ~n8254 & n8256;
  assign n8258 = ~pi23  & ~n8257;
  assign n8259 = pi23  & n8257;
  assign n8260 = ~n8258 & ~n8259;
  assign n8261 = n8073 & ~n8075;
  assign n8262 = ~n8076 & ~n8261;
  assign n8263 = ~n8260 & n8262;
  assign n8264 = ~n2622 & n5267;
  assign n8265 = ~n2726 & n5121;
  assign n8266 = ~n2657 & n5185;
  assign n8267 = n78 & n6407;
  assign n8268 = ~n8264 & ~n8266;
  assign n8269 = ~n8265 & n8268;
  assign n8270 = ~n8267 & n8269;
  assign n8271 = ~pi23  & ~n8270;
  assign n8272 = pi23  & n8270;
  assign n8273 = ~n8271 & ~n8272;
  assign n8274 = n8069 & ~n8071;
  assign n8275 = ~n8072 & ~n8274;
  assign n8276 = ~n8273 & n8275;
  assign n8277 = ~n2657 & n5267;
  assign n8278 = ~n2726 & n5185;
  assign n8279 = ~n2781 & n5121;
  assign n8280 = n78 & n6251;
  assign n8281 = ~n8277 & ~n8279;
  assign n8282 = ~n8278 & n8281;
  assign n8283 = ~n8280 & n8282;
  assign n8284 = ~pi23  & ~n8283;
  assign n8285 = pi23  & n8283;
  assign n8286 = ~n8284 & ~n8285;
  assign n8287 = n8065 & ~n8067;
  assign n8288 = ~n8068 & ~n8287;
  assign n8289 = ~n8286 & n8288;
  assign n8290 = ~n2866 & n5121;
  assign n8291 = ~n2726 & n5267;
  assign n8292 = ~n2781 & n5185;
  assign n8293 = n78 & n6520;
  assign n8294 = ~n8290 & ~n8292;
  assign n8295 = ~n8291 & n8294;
  assign n8296 = ~n8293 & n8295;
  assign n8297 = ~pi23  & ~n8296;
  assign n8298 = pi23  & n8296;
  assign n8299 = ~n8297 & ~n8298;
  assign n8300 = n8061 & ~n8063;
  assign n8301 = ~n8064 & ~n8300;
  assign n8302 = ~n8299 & n8301;
  assign n8303 = ~n2866 & n5185;
  assign n8304 = ~n2781 & n5267;
  assign n8305 = ~n2901 & n5121;
  assign n8306 = n78 & n6819;
  assign n8307 = ~n8303 & ~n8304;
  assign n8308 = ~n8305 & n8307;
  assign n8309 = ~n8306 & n8308;
  assign n8310 = ~pi23  & ~n8309;
  assign n8311 = pi23  & n8309;
  assign n8312 = ~n8310 & ~n8311;
  assign n8313 = n8057 & ~n8059;
  assign n8314 = ~n8060 & ~n8313;
  assign n8315 = ~n8312 & n8314;
  assign n8316 = n8053 & ~n8055;
  assign n8317 = ~n8056 & ~n8316;
  assign n8318 = ~n2866 & n5267;
  assign n8319 = ~n2978 & n5121;
  assign n8320 = ~n2901 & n5185;
  assign n8321 = n78 & n6831;
  assign n8322 = ~n8318 & ~n8320;
  assign n8323 = ~n8319 & n8322;
  assign n8324 = ~n8321 & n8323;
  assign n8325 = pi23  & n8324;
  assign n8326 = ~pi23  & ~n8324;
  assign n8327 = ~n8325 & ~n8326;
  assign n8328 = n8317 & ~n8327;
  assign n8329 = n8049 & ~n8051;
  assign n8330 = ~n8052 & ~n8329;
  assign n8331 = ~n2901 & n5267;
  assign n8332 = ~n2978 & n5185;
  assign n8333 = ~n3069 & n5121;
  assign n8334 = n78 & n6496;
  assign n8335 = ~n8331 & ~n8333;
  assign n8336 = ~n8332 & n8335;
  assign n8337 = ~n8334 & n8336;
  assign n8338 = pi23  & n8337;
  assign n8339 = ~pi23  & ~n8337;
  assign n8340 = ~n8338 & ~n8339;
  assign n8341 = n8330 & ~n8340;
  assign n8342 = ~n2978 & n5267;
  assign n8343 = ~n3137 & n5121;
  assign n8344 = ~n3069 & n5185;
  assign n8345 = n78 & n6873;
  assign n8346 = ~n8342 & ~n8344;
  assign n8347 = ~n8343 & n8346;
  assign n8348 = ~n8345 & n8347;
  assign n8349 = ~pi23  & ~n8348;
  assign n8350 = pi23  & n8348;
  assign n8351 = ~n8349 & ~n8350;
  assign n8352 = n8045 & ~n8047;
  assign n8353 = ~n8048 & ~n8352;
  assign n8354 = ~n8351 & n8353;
  assign n8355 = ~n3069 & n5267;
  assign n8356 = ~n3137 & n5185;
  assign n8357 = ~n3194 & n5121;
  assign n8358 = n78 & n6920;
  assign n8359 = ~n8355 & ~n8357;
  assign n8360 = ~n8356 & n8359;
  assign n8361 = ~n8358 & n8360;
  assign n8362 = pi23  & n8361;
  assign n8363 = ~pi23  & ~n8361;
  assign n8364 = ~n8362 & ~n8363;
  assign n8365 = n8041 & ~n8043;
  assign n8366 = ~n8044 & ~n8365;
  assign n8367 = ~n8364 & n8366;
  assign n8368 = ~n3137 & n5267;
  assign n8369 = ~n3194 & n5185;
  assign n8370 = ~n3227 & n5121;
  assign n8371 = n78 & n6970;
  assign n8372 = ~n8369 & ~n8370;
  assign n8373 = ~n8368 & n8372;
  assign n8374 = ~n8371 & n8373;
  assign n8375 = ~pi23  & ~n8374;
  assign n8376 = pi23  & n8374;
  assign n8377 = ~n8375 & ~n8376;
  assign n8378 = pi26  & ~n8021;
  assign n8379 = n8028 & ~n8378;
  assign n8380 = ~n8028 & n8378;
  assign n8381 = ~n8379 & ~n8380;
  assign n8382 = ~n8377 & n8381;
  assign n8383 = ~n3319 & n5121;
  assign n8384 = ~n3227 & n5185;
  assign n8385 = ~n3194 & n5267;
  assign n8386 = n78 & n7013;
  assign n8387 = ~n8384 & ~n8385;
  assign n8388 = ~n8383 & n8387;
  assign n8389 = ~n8386 & n8388;
  assign n8390 = pi23  & n8389;
  assign n8391 = ~pi23  & ~n8389;
  assign n8392 = ~n8390 & ~n8391;
  assign n8393 = n8015 & ~n8020;
  assign n8394 = ~n8021 & ~n8393;
  assign n8395 = ~n8392 & n8394;
  assign n8396 = n74 & ~n3460;
  assign n8397 = pi23  & n8396;
  assign n8398 = ~n3376 & n5267;
  assign n8399 = ~n3460 & n5185;
  assign n8400 = n78 & ~n7689;
  assign n8401 = ~n8398 & ~n8399;
  assign n8402 = ~n8400 & n8401;
  assign n8403 = ~n8397 & n8402;
  assign n8404 = ~n3460 & n5121;
  assign n8405 = ~n3319 & n5267;
  assign n8406 = ~n3376 & n5185;
  assign n8407 = n78 & n7049;
  assign n8408 = ~n8404 & ~n8406;
  assign n8409 = ~n8405 & n8408;
  assign n8410 = ~n8407 & n8409;
  assign n8411 = pi23  & n8403;
  assign n8412 = n8410 & n8411;
  assign n8413 = n8014 & n8412;
  assign n8414 = ~n3319 & n5185;
  assign n8415 = ~n3376 & n5121;
  assign n8416 = ~n3227 & n5267;
  assign n8417 = n78 & n7105;
  assign n8418 = ~n8415 & ~n8416;
  assign n8419 = ~n8414 & n8418;
  assign n8420 = ~n8417 & n8419;
  assign n8421 = pi23  & n8420;
  assign n8422 = ~pi23  & ~n8420;
  assign n8423 = ~n8421 & ~n8422;
  assign n8424 = ~n8014 & ~n8412;
  assign n8425 = ~n8413 & ~n8424;
  assign n8426 = ~n8423 & n8425;
  assign n8427 = ~n8413 & ~n8426;
  assign n8428 = n8392 & ~n8394;
  assign n8429 = ~n8395 & ~n8428;
  assign n8430 = ~n8427 & n8429;
  assign n8431 = ~n8395 & ~n8430;
  assign n8432 = n8377 & ~n8381;
  assign n8433 = ~n8382 & ~n8432;
  assign n8434 = ~n8431 & n8433;
  assign n8435 = ~n8382 & ~n8434;
  assign n8436 = n8364 & ~n8366;
  assign n8437 = ~n8367 & ~n8436;
  assign n8438 = ~n8435 & n8437;
  assign n8439 = ~n8367 & ~n8438;
  assign n8440 = n8351 & ~n8353;
  assign n8441 = ~n8354 & ~n8440;
  assign n8442 = ~n8439 & n8441;
  assign n8443 = ~n8354 & ~n8442;
  assign n8444 = ~n8330 & n8340;
  assign n8445 = ~n8341 & ~n8444;
  assign n8446 = ~n8443 & n8445;
  assign n8447 = ~n8341 & ~n8446;
  assign n8448 = ~n8317 & n8327;
  assign n8449 = ~n8328 & ~n8448;
  assign n8450 = ~n8447 & n8449;
  assign n8451 = ~n8328 & ~n8450;
  assign n8452 = n8312 & ~n8314;
  assign n8453 = ~n8315 & ~n8452;
  assign n8454 = ~n8451 & n8453;
  assign n8455 = ~n8315 & ~n8454;
  assign n8456 = n8299 & ~n8301;
  assign n8457 = ~n8302 & ~n8456;
  assign n8458 = ~n8455 & n8457;
  assign n8459 = ~n8302 & ~n8458;
  assign n8460 = n8286 & ~n8288;
  assign n8461 = ~n8289 & ~n8460;
  assign n8462 = ~n8459 & n8461;
  assign n8463 = ~n8289 & ~n8462;
  assign n8464 = n8273 & ~n8275;
  assign n8465 = ~n8276 & ~n8464;
  assign n8466 = ~n8463 & n8465;
  assign n8467 = ~n8276 & ~n8466;
  assign n8468 = n8260 & ~n8262;
  assign n8469 = ~n8263 & ~n8468;
  assign n8470 = ~n8467 & n8469;
  assign n8471 = ~n8263 & ~n8470;
  assign n8472 = n8247 & ~n8249;
  assign n8473 = ~n8250 & ~n8472;
  assign n8474 = ~n8471 & n8473;
  assign n8475 = ~n8250 & ~n8474;
  assign n8476 = n8234 & ~n8236;
  assign n8477 = ~n8237 & ~n8476;
  assign n8478 = ~n8475 & n8477;
  assign n8479 = ~n8237 & ~n8478;
  assign n8480 = n8098 & ~n8100;
  assign n8481 = ~n8101 & ~n8480;
  assign n8482 = ~n8479 & n8481;
  assign n8483 = ~n2165 & n5312;
  assign n8484 = ~n2045 & n5901;
  assign n8485 = ~n1997 & n5982;
  assign n8486 = n5306 & n5424;
  assign n8487 = ~n8484 & ~n8485;
  assign n8488 = ~n8483 & n8487;
  assign n8489 = ~n8486 & n8488;
  assign n8490 = ~pi20  & ~n8489;
  assign n8491 = pi20  & n8489;
  assign n8492 = ~n8490 & ~n8491;
  assign n8493 = n8479 & ~n8481;
  assign n8494 = ~n8482 & ~n8493;
  assign n8495 = ~n8492 & n8494;
  assign n8496 = ~n8482 & ~n8495;
  assign n8497 = ~n8107 & n8117;
  assign n8498 = ~n8118 & ~n8497;
  assign n8499 = ~n8496 & n8498;
  assign n8500 = n8496 & ~n8498;
  assign n8501 = ~n8499 & ~n8500;
  assign n8502 = ~n1805 & n6140;
  assign n8503 = ~n1737 & n6356;
  assign n8504 = ~n1610 & n6608;
  assign n8505 = n4844 & n6134;
  assign n8506 = ~n8502 & ~n8503;
  assign n8507 = ~n8504 & n8506;
  assign n8508 = ~n8505 & n8507;
  assign n8509 = pi17  & n8508;
  assign n8510 = ~pi17  & ~n8508;
  assign n8511 = ~n8509 & ~n8510;
  assign n8512 = n8501 & ~n8511;
  assign n8513 = ~n8499 & ~n8512;
  assign n8514 = ~n8124 & n8134;
  assign n8515 = ~n8135 & ~n8514;
  assign n8516 = ~n8513 & n8515;
  assign n8517 = n8513 & ~n8515;
  assign n8518 = ~n8516 & ~n8517;
  assign n8519 = ~n1425 & n6653;
  assign n8520 = ~n1337 & n7243;
  assign n8521 = ~n1230 & n7380;
  assign n8522 = n4549 & n6647;
  assign n8523 = ~n8519 & ~n8520;
  assign n8524 = ~n8521 & n8523;
  assign n8525 = ~n8522 & n8524;
  assign n8526 = pi14  & n8525;
  assign n8527 = ~pi14  & ~n8525;
  assign n8528 = ~n8526 & ~n8527;
  assign n8529 = n8518 & ~n8528;
  assign n8530 = ~n8516 & ~n8529;
  assign n8531 = ~n8213 & n8223;
  assign n8532 = ~n8224 & ~n8531;
  assign n8533 = ~n8530 & n8532;
  assign n8534 = ~n8224 & ~n8533;
  assign n8535 = ~n8143 & n8153;
  assign n8536 = ~n8154 & ~n8535;
  assign n8537 = n8534 & ~n8536;
  assign n8538 = ~n8534 & n8536;
  assign n8539 = ~n8537 & ~n8538;
  assign n8540 = ~n729 & n8161;
  assign n8541 = ~n802 & n7847;
  assign n8542 = ~n898 & n7554;
  assign n8543 = n3901 & n7548;
  assign n8544 = ~n8541 & ~n8542;
  assign n8545 = ~n8540 & n8544;
  assign n8546 = ~n8543 & n8545;
  assign n8547 = pi11  & n8546;
  assign n8548 = ~pi11  & ~n8546;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = n8539 & n8549;
  assign n8551 = ~n8537 & ~n8550;
  assign n8552 = ~n8211 & n8551;
  assign n8553 = n8211 & ~n8551;
  assign n8554 = ~n8552 & ~n8553;
  assign n8555 = ~n8160 & n8171;
  assign n8556 = ~n8172 & ~n8555;
  assign n8557 = n8554 & n8556;
  assign n8558 = ~n8552 & ~n8557;
  assign n8559 = ~n8186 & ~n8188;
  assign n8560 = ~n8189 & ~n8559;
  assign n8561 = ~n8558 & n8560;
  assign n8562 = n8558 & ~n8560;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = n8475 & ~n8477;
  assign n8565 = ~n8478 & ~n8564;
  assign n8566 = ~n2165 & n5901;
  assign n8567 = ~n2265 & n5312;
  assign n8568 = ~n2045 & n5982;
  assign n8569 = n5306 & n5408;
  assign n8570 = ~n8567 & ~n8568;
  assign n8571 = ~n8566 & n8570;
  assign n8572 = ~n8569 & n8571;
  assign n8573 = pi20  & n8572;
  assign n8574 = ~pi20  & ~n8572;
  assign n8575 = ~n8573 & ~n8574;
  assign n8576 = n8565 & ~n8575;
  assign n8577 = n8471 & ~n8473;
  assign n8578 = ~n8474 & ~n8577;
  assign n8579 = ~n2356 & n5312;
  assign n8580 = ~n2265 & n5901;
  assign n8581 = ~n2165 & n5982;
  assign n8582 = n5306 & n5632;
  assign n8583 = ~n8579 & ~n8580;
  assign n8584 = ~n8581 & n8583;
  assign n8585 = ~n8582 & n8584;
  assign n8586 = pi20  & n8585;
  assign n8587 = ~pi20  & ~n8585;
  assign n8588 = ~n8586 & ~n8587;
  assign n8589 = n8578 & ~n8588;
  assign n8590 = n8467 & ~n8469;
  assign n8591 = ~n8470 & ~n8590;
  assign n8592 = ~n2356 & n5901;
  assign n8593 = ~n2442 & n5312;
  assign n8594 = ~n2265 & n5982;
  assign n8595 = n5306 & n5650;
  assign n8596 = ~n8593 & ~n8594;
  assign n8597 = ~n8592 & n8596;
  assign n8598 = ~n8595 & n8597;
  assign n8599 = pi20  & n8598;
  assign n8600 = ~pi20  & ~n8598;
  assign n8601 = ~n8599 & ~n8600;
  assign n8602 = n8591 & ~n8601;
  assign n8603 = n8463 & ~n8465;
  assign n8604 = ~n8466 & ~n8603;
  assign n8605 = ~n2356 & n5982;
  assign n8606 = ~n2538 & n5312;
  assign n8607 = ~n2442 & n5901;
  assign n8608 = n5306 & n6042;
  assign n8609 = ~n8605 & ~n8607;
  assign n8610 = ~n8606 & n8609;
  assign n8611 = ~n8608 & n8610;
  assign n8612 = pi20  & n8611;
  assign n8613 = ~pi20  & ~n8611;
  assign n8614 = ~n8612 & ~n8613;
  assign n8615 = n8604 & ~n8614;
  assign n8616 = n8459 & ~n8461;
  assign n8617 = ~n8462 & ~n8616;
  assign n8618 = ~n2622 & n5312;
  assign n8619 = ~n2538 & n5901;
  assign n8620 = ~n2442 & n5982;
  assign n8621 = n5306 & n5823;
  assign n8622 = ~n8618 & ~n8620;
  assign n8623 = ~n8619 & n8622;
  assign n8624 = ~n8621 & n8623;
  assign n8625 = pi20  & n8624;
  assign n8626 = ~pi20  & ~n8624;
  assign n8627 = ~n8625 & ~n8626;
  assign n8628 = n8617 & ~n8627;
  assign n8629 = n8455 & ~n8457;
  assign n8630 = ~n8458 & ~n8629;
  assign n8631 = ~n2538 & n5982;
  assign n8632 = ~n2622 & n5901;
  assign n8633 = ~n2657 & n5312;
  assign n8634 = n5306 & n6271;
  assign n8635 = ~n8631 & ~n8633;
  assign n8636 = ~n8632 & n8635;
  assign n8637 = ~n8634 & n8636;
  assign n8638 = pi20  & n8637;
  assign n8639 = ~pi20  & ~n8637;
  assign n8640 = ~n8638 & ~n8639;
  assign n8641 = n8630 & ~n8640;
  assign n8642 = n8451 & ~n8453;
  assign n8643 = ~n8454 & ~n8642;
  assign n8644 = ~n2622 & n5982;
  assign n8645 = ~n2726 & n5312;
  assign n8646 = ~n2657 & n5901;
  assign n8647 = n5306 & n6407;
  assign n8648 = ~n8644 & ~n8646;
  assign n8649 = ~n8645 & n8648;
  assign n8650 = ~n8647 & n8649;
  assign n8651 = pi20  & n8650;
  assign n8652 = ~pi20  & ~n8650;
  assign n8653 = ~n8651 & ~n8652;
  assign n8654 = n8643 & ~n8653;
  assign n8655 = ~n2657 & n5982;
  assign n8656 = ~n2726 & n5901;
  assign n8657 = ~n2781 & n5312;
  assign n8658 = n5306 & n6251;
  assign n8659 = ~n8655 & ~n8657;
  assign n8660 = ~n8656 & n8659;
  assign n8661 = ~n8658 & n8660;
  assign n8662 = ~pi20  & ~n8661;
  assign n8663 = pi20  & n8661;
  assign n8664 = ~n8662 & ~n8663;
  assign n8665 = n8447 & ~n8449;
  assign n8666 = ~n8450 & ~n8665;
  assign n8667 = ~n8664 & n8666;
  assign n8668 = ~n2866 & n5312;
  assign n8669 = ~n2726 & n5982;
  assign n8670 = ~n2781 & n5901;
  assign n8671 = n5306 & n6520;
  assign n8672 = ~n8668 & ~n8670;
  assign n8673 = ~n8669 & n8672;
  assign n8674 = ~n8671 & n8673;
  assign n8675 = ~pi20  & ~n8674;
  assign n8676 = pi20  & n8674;
  assign n8677 = ~n8675 & ~n8676;
  assign n8678 = n8443 & ~n8445;
  assign n8679 = ~n8446 & ~n8678;
  assign n8680 = ~n8677 & n8679;
  assign n8681 = n8439 & ~n8441;
  assign n8682 = ~n8442 & ~n8681;
  assign n8683 = ~n2866 & n5901;
  assign n8684 = ~n2781 & n5982;
  assign n8685 = ~n2901 & n5312;
  assign n8686 = n5306 & n6819;
  assign n8687 = ~n8683 & ~n8684;
  assign n8688 = ~n8685 & n8687;
  assign n8689 = ~n8686 & n8688;
  assign n8690 = pi20  & n8689;
  assign n8691 = ~pi20  & ~n8689;
  assign n8692 = ~n8690 & ~n8691;
  assign n8693 = n8682 & ~n8692;
  assign n8694 = n8435 & ~n8437;
  assign n8695 = ~n8438 & ~n8694;
  assign n8696 = ~n2866 & n5982;
  assign n8697 = ~n2978 & n5312;
  assign n8698 = ~n2901 & n5901;
  assign n8699 = n5306 & n6831;
  assign n8700 = ~n8696 & ~n8698;
  assign n8701 = ~n8697 & n8700;
  assign n8702 = ~n8699 & n8701;
  assign n8703 = pi20  & n8702;
  assign n8704 = ~pi20  & ~n8702;
  assign n8705 = ~n8703 & ~n8704;
  assign n8706 = n8695 & ~n8705;
  assign n8707 = n8431 & ~n8433;
  assign n8708 = ~n8434 & ~n8707;
  assign n8709 = ~n2901 & n5982;
  assign n8710 = ~n2978 & n5901;
  assign n8711 = ~n3069 & n5312;
  assign n8712 = n5306 & n6496;
  assign n8713 = ~n8709 & ~n8711;
  assign n8714 = ~n8710 & n8713;
  assign n8715 = ~n8712 & n8714;
  assign n8716 = pi20  & n8715;
  assign n8717 = ~pi20  & ~n8715;
  assign n8718 = ~n8716 & ~n8717;
  assign n8719 = n8708 & ~n8718;
  assign n8720 = ~n2978 & n5982;
  assign n8721 = ~n3137 & n5312;
  assign n8722 = ~n3069 & n5901;
  assign n8723 = n5306 & n6873;
  assign n8724 = ~n8720 & ~n8722;
  assign n8725 = ~n8721 & n8724;
  assign n8726 = ~n8723 & n8725;
  assign n8727 = ~pi20  & ~n8726;
  assign n8728 = pi20  & n8726;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = n8427 & ~n8429;
  assign n8731 = ~n8430 & ~n8730;
  assign n8732 = ~n8729 & n8731;
  assign n8733 = ~n3069 & n5982;
  assign n8734 = ~n3137 & n5901;
  assign n8735 = ~n3194 & n5312;
  assign n8736 = n5306 & n6920;
  assign n8737 = ~n8733 & ~n8735;
  assign n8738 = ~n8734 & n8737;
  assign n8739 = ~n8736 & n8738;
  assign n8740 = pi20  & n8739;
  assign n8741 = ~pi20  & ~n8739;
  assign n8742 = ~n8740 & ~n8741;
  assign n8743 = n8423 & ~n8425;
  assign n8744 = ~n8426 & ~n8743;
  assign n8745 = ~n8742 & n8744;
  assign n8746 = ~n3137 & n5982;
  assign n8747 = ~n3194 & n5901;
  assign n8748 = ~n3227 & n5312;
  assign n8749 = n5306 & n6970;
  assign n8750 = ~n8747 & ~n8748;
  assign n8751 = ~n8746 & n8750;
  assign n8752 = ~n8749 & n8751;
  assign n8753 = ~pi20  & ~n8752;
  assign n8754 = pi20  & n8752;
  assign n8755 = ~n8753 & ~n8754;
  assign n8756 = pi23  & ~n8403;
  assign n8757 = n8410 & ~n8756;
  assign n8758 = ~n8410 & n8756;
  assign n8759 = ~n8757 & ~n8758;
  assign n8760 = ~n8755 & n8759;
  assign n8761 = ~n3319 & n5312;
  assign n8762 = ~n3227 & n5901;
  assign n8763 = ~n3194 & n5982;
  assign n8764 = n5306 & n7013;
  assign n8765 = ~n8762 & ~n8763;
  assign n8766 = ~n8761 & n8765;
  assign n8767 = ~n8764 & n8766;
  assign n8768 = pi20  & n8767;
  assign n8769 = ~pi20  & ~n8767;
  assign n8770 = ~n8768 & ~n8769;
  assign n8771 = n8397 & ~n8402;
  assign n8772 = ~n8403 & ~n8771;
  assign n8773 = ~n8770 & n8772;
  assign n8774 = ~n3460 & n5305;
  assign n8775 = pi20  & n8774;
  assign n8776 = ~n3376 & n5982;
  assign n8777 = ~n3460 & n5901;
  assign n8778 = n5306 & ~n7689;
  assign n8779 = ~n8776 & ~n8777;
  assign n8780 = ~n8778 & n8779;
  assign n8781 = ~n8775 & n8780;
  assign n8782 = ~n3460 & n5312;
  assign n8783 = ~n3319 & n5982;
  assign n8784 = ~n3376 & n5901;
  assign n8785 = n5306 & n7049;
  assign n8786 = ~n8782 & ~n8784;
  assign n8787 = ~n8783 & n8786;
  assign n8788 = ~n8785 & n8787;
  assign n8789 = pi20  & n8781;
  assign n8790 = n8788 & n8789;
  assign n8791 = n8396 & n8790;
  assign n8792 = ~n3319 & n5901;
  assign n8793 = ~n3376 & n5312;
  assign n8794 = ~n3227 & n5982;
  assign n8795 = n5306 & n7105;
  assign n8796 = ~n8793 & ~n8794;
  assign n8797 = ~n8792 & n8796;
  assign n8798 = ~n8795 & n8797;
  assign n8799 = pi20  & n8798;
  assign n8800 = ~pi20  & ~n8798;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = ~n8396 & ~n8790;
  assign n8803 = ~n8791 & ~n8802;
  assign n8804 = ~n8801 & n8803;
  assign n8805 = ~n8791 & ~n8804;
  assign n8806 = n8770 & ~n8772;
  assign n8807 = ~n8773 & ~n8806;
  assign n8808 = ~n8805 & n8807;
  assign n8809 = ~n8773 & ~n8808;
  assign n8810 = n8755 & ~n8759;
  assign n8811 = ~n8760 & ~n8810;
  assign n8812 = ~n8809 & n8811;
  assign n8813 = ~n8760 & ~n8812;
  assign n8814 = n8742 & ~n8744;
  assign n8815 = ~n8745 & ~n8814;
  assign n8816 = ~n8813 & n8815;
  assign n8817 = ~n8745 & ~n8816;
  assign n8818 = n8729 & ~n8731;
  assign n8819 = ~n8732 & ~n8818;
  assign n8820 = ~n8817 & n8819;
  assign n8821 = ~n8732 & ~n8820;
  assign n8822 = ~n8708 & n8718;
  assign n8823 = ~n8719 & ~n8822;
  assign n8824 = ~n8821 & n8823;
  assign n8825 = ~n8719 & ~n8824;
  assign n8826 = ~n8695 & n8705;
  assign n8827 = ~n8706 & ~n8826;
  assign n8828 = ~n8825 & n8827;
  assign n8829 = ~n8706 & ~n8828;
  assign n8830 = ~n8682 & n8692;
  assign n8831 = ~n8693 & ~n8830;
  assign n8832 = ~n8829 & n8831;
  assign n8833 = ~n8693 & ~n8832;
  assign n8834 = n8677 & ~n8679;
  assign n8835 = ~n8680 & ~n8834;
  assign n8836 = ~n8833 & n8835;
  assign n8837 = ~n8680 & ~n8836;
  assign n8838 = n8664 & ~n8666;
  assign n8839 = ~n8667 & ~n8838;
  assign n8840 = ~n8837 & n8839;
  assign n8841 = ~n8667 & ~n8840;
  assign n8842 = ~n8643 & n8653;
  assign n8843 = ~n8654 & ~n8842;
  assign n8844 = ~n8841 & n8843;
  assign n8845 = ~n8654 & ~n8844;
  assign n8846 = ~n8630 & n8640;
  assign n8847 = ~n8641 & ~n8846;
  assign n8848 = ~n8845 & n8847;
  assign n8849 = ~n8641 & ~n8848;
  assign n8850 = ~n8617 & n8627;
  assign n8851 = ~n8628 & ~n8850;
  assign n8852 = ~n8849 & n8851;
  assign n8853 = ~n8628 & ~n8852;
  assign n8854 = ~n8604 & n8614;
  assign n8855 = ~n8615 & ~n8854;
  assign n8856 = ~n8853 & n8855;
  assign n8857 = ~n8615 & ~n8856;
  assign n8858 = ~n8591 & n8601;
  assign n8859 = ~n8602 & ~n8858;
  assign n8860 = ~n8857 & n8859;
  assign n8861 = ~n8602 & ~n8860;
  assign n8862 = ~n8578 & n8588;
  assign n8863 = ~n8589 & ~n8862;
  assign n8864 = ~n8861 & n8863;
  assign n8865 = ~n8589 & ~n8864;
  assign n8866 = ~n8565 & n8575;
  assign n8867 = ~n8576 & ~n8866;
  assign n8868 = ~n8865 & n8867;
  assign n8869 = ~n8576 & ~n8868;
  assign n8870 = n8492 & ~n8494;
  assign n8871 = ~n8495 & ~n8870;
  assign n8872 = ~n8869 & n8871;
  assign n8873 = ~n1893 & n6140;
  assign n8874 = ~n1805 & n6356;
  assign n8875 = ~n1737 & n6608;
  assign n8876 = n4862 & n6134;
  assign n8877 = ~n8873 & ~n8874;
  assign n8878 = ~n8875 & n8877;
  assign n8879 = ~n8876 & n8878;
  assign n8880 = ~pi17  & ~n8879;
  assign n8881 = pi17  & n8879;
  assign n8882 = ~n8880 & ~n8881;
  assign n8883 = n8869 & ~n8871;
  assign n8884 = ~n8872 & ~n8883;
  assign n8885 = ~n8882 & n8884;
  assign n8886 = ~n8872 & ~n8885;
  assign n8887 = ~n8501 & n8511;
  assign n8888 = ~n8512 & ~n8887;
  assign n8889 = ~n8886 & n8888;
  assign n8890 = n8886 & ~n8888;
  assign n8891 = ~n8889 & ~n8890;
  assign n8892 = ~n1532 & n6653;
  assign n8893 = ~n1425 & n7243;
  assign n8894 = ~n1337 & n7380;
  assign n8895 = n4452 & n6647;
  assign n8896 = ~n8892 & ~n8893;
  assign n8897 = ~n8894 & n8896;
  assign n8898 = ~n8895 & n8897;
  assign n8899 = pi14  & n8898;
  assign n8900 = ~pi14  & ~n8898;
  assign n8901 = ~n8899 & ~n8900;
  assign n8902 = n8891 & ~n8901;
  assign n8903 = ~n8889 & ~n8902;
  assign n8904 = ~n8518 & n8528;
  assign n8905 = ~n8529 & ~n8904;
  assign n8906 = ~n8903 & n8905;
  assign n8907 = n8903 & ~n8905;
  assign n8908 = ~n8906 & ~n8907;
  assign n8909 = ~n898 & n8161;
  assign n8910 = ~n1006 & n7847;
  assign n8911 = ~n1107 & n7554;
  assign n8912 = n4041 & n7548;
  assign n8913 = ~n8909 & ~n8910;
  assign n8914 = ~n8911 & n8913;
  assign n8915 = ~n8912 & n8914;
  assign n8916 = pi11  & n8915;
  assign n8917 = ~pi11  & ~n8915;
  assign n8918 = ~n8916 & ~n8917;
  assign n8919 = n8908 & ~n8918;
  assign n8920 = ~n8906 & ~n8919;
  assign n8921 = ~n802 & n8161;
  assign n8922 = ~n898 & n7847;
  assign n8923 = ~n1006 & n7554;
  assign n8924 = n4057 & n7548;
  assign n8925 = ~n8921 & ~n8922;
  assign n8926 = ~n8923 & n8925;
  assign n8927 = ~n8924 & n8926;
  assign n8928 = pi11  & n8927;
  assign n8929 = ~pi11  & ~n8927;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 = ~n8920 & ~n8930;
  assign n8932 = n8920 & n8930;
  assign n8933 = ~n8931 & ~n8932;
  assign n8934 = n8530 & ~n8532;
  assign n8935 = ~n8533 & ~n8934;
  assign n8936 = n8933 & n8935;
  assign n8937 = ~n8931 & ~n8936;
  assign n8938 = ~n621 & n8206;
  assign n8939 = ~n8199 & n8204;
  assign n8940 = ~n563 & n8939;
  assign n8941 = n3687 & n8200;
  assign n8942 = ~n8938 & ~n8940;
  assign n8943 = ~n8941 & n8942;
  assign n8944 = pi8  & n8943;
  assign n8945 = ~pi8  & ~n8943;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = ~n8937 & ~n8946;
  assign n8948 = ~n8539 & ~n8549;
  assign n8949 = ~n8550 & ~n8948;
  assign n8950 = n8937 & n8946;
  assign n8951 = ~n8947 & ~n8950;
  assign n8952 = ~n8949 & n8951;
  assign n8953 = ~n8947 & ~n8952;
  assign n8954 = ~n8554 & ~n8556;
  assign n8955 = ~n8557 & ~n8954;
  assign n8956 = ~n8953 & n8955;
  assign n8957 = n8953 & ~n8955;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = ~n1997 & n6140;
  assign n8960 = ~n1893 & n6356;
  assign n8961 = ~n1805 & n6608;
  assign n8962 = n5212 & n6134;
  assign n8963 = ~n8959 & ~n8960;
  assign n8964 = ~n8961 & n8963;
  assign n8965 = ~n8962 & n8964;
  assign n8966 = ~pi17  & ~n8965;
  assign n8967 = pi17  & n8965;
  assign n8968 = ~n8966 & ~n8967;
  assign n8969 = n8865 & ~n8867;
  assign n8970 = ~n8868 & ~n8969;
  assign n8971 = ~n8968 & n8970;
  assign n8972 = ~n2045 & n6140;
  assign n8973 = ~n1997 & n6356;
  assign n8974 = ~n1893 & n6608;
  assign n8975 = n5061 & n6134;
  assign n8976 = ~n8972 & ~n8973;
  assign n8977 = ~n8974 & n8976;
  assign n8978 = ~n8975 & n8977;
  assign n8979 = ~pi17  & ~n8978;
  assign n8980 = pi17  & n8978;
  assign n8981 = ~n8979 & ~n8980;
  assign n8982 = n8861 & ~n8863;
  assign n8983 = ~n8864 & ~n8982;
  assign n8984 = ~n8981 & n8983;
  assign n8985 = ~n2165 & n6140;
  assign n8986 = ~n2045 & n6356;
  assign n8987 = ~n1997 & n6608;
  assign n8988 = n5424 & n6134;
  assign n8989 = ~n8986 & ~n8987;
  assign n8990 = ~n8985 & n8989;
  assign n8991 = ~n8988 & n8990;
  assign n8992 = ~pi17  & ~n8991;
  assign n8993 = pi17  & n8991;
  assign n8994 = ~n8992 & ~n8993;
  assign n8995 = n8857 & ~n8859;
  assign n8996 = ~n8860 & ~n8995;
  assign n8997 = ~n8994 & n8996;
  assign n8998 = ~n2165 & n6356;
  assign n8999 = ~n2265 & n6140;
  assign n9000 = ~n2045 & n6608;
  assign n9001 = n5408 & n6134;
  assign n9002 = ~n8999 & ~n9000;
  assign n9003 = ~n8998 & n9002;
  assign n9004 = ~n9001 & n9003;
  assign n9005 = ~pi17  & ~n9004;
  assign n9006 = pi17  & n9004;
  assign n9007 = ~n9005 & ~n9006;
  assign n9008 = n8853 & ~n8855;
  assign n9009 = ~n8856 & ~n9008;
  assign n9010 = ~n9007 & n9009;
  assign n9011 = ~n2356 & n6140;
  assign n9012 = ~n2265 & n6356;
  assign n9013 = ~n2165 & n6608;
  assign n9014 = n5632 & n6134;
  assign n9015 = ~n9011 & ~n9012;
  assign n9016 = ~n9013 & n9015;
  assign n9017 = ~n9014 & n9016;
  assign n9018 = ~pi17  & ~n9017;
  assign n9019 = pi17  & n9017;
  assign n9020 = ~n9018 & ~n9019;
  assign n9021 = n8849 & ~n8851;
  assign n9022 = ~n8852 & ~n9021;
  assign n9023 = ~n9020 & n9022;
  assign n9024 = ~n2356 & n6356;
  assign n9025 = ~n2442 & n6140;
  assign n9026 = ~n2265 & n6608;
  assign n9027 = n5650 & n6134;
  assign n9028 = ~n9025 & ~n9026;
  assign n9029 = ~n9024 & n9028;
  assign n9030 = ~n9027 & n9029;
  assign n9031 = ~pi17  & ~n9030;
  assign n9032 = pi17  & n9030;
  assign n9033 = ~n9031 & ~n9032;
  assign n9034 = n8845 & ~n8847;
  assign n9035 = ~n8848 & ~n9034;
  assign n9036 = ~n9033 & n9035;
  assign n9037 = ~n2356 & n6608;
  assign n9038 = ~n2538 & n6140;
  assign n9039 = ~n2442 & n6356;
  assign n9040 = n6042 & n6134;
  assign n9041 = ~n9037 & ~n9039;
  assign n9042 = ~n9038 & n9041;
  assign n9043 = ~n9040 & n9042;
  assign n9044 = ~pi17  & ~n9043;
  assign n9045 = pi17  & n9043;
  assign n9046 = ~n9044 & ~n9045;
  assign n9047 = n8841 & ~n8843;
  assign n9048 = ~n8844 & ~n9047;
  assign n9049 = ~n9046 & n9048;
  assign n9050 = n8837 & ~n8839;
  assign n9051 = ~n8840 & ~n9050;
  assign n9052 = ~n2622 & n6140;
  assign n9053 = ~n2538 & n6356;
  assign n9054 = ~n2442 & n6608;
  assign n9055 = n5823 & n6134;
  assign n9056 = ~n9052 & ~n9054;
  assign n9057 = ~n9053 & n9056;
  assign n9058 = ~n9055 & n9057;
  assign n9059 = pi17  & n9058;
  assign n9060 = ~pi17  & ~n9058;
  assign n9061 = ~n9059 & ~n9060;
  assign n9062 = n9051 & ~n9061;
  assign n9063 = n8833 & ~n8835;
  assign n9064 = ~n8836 & ~n9063;
  assign n9065 = ~n2538 & n6608;
  assign n9066 = ~n2622 & n6356;
  assign n9067 = ~n2657 & n6140;
  assign n9068 = n6134 & n6271;
  assign n9069 = ~n9065 & ~n9067;
  assign n9070 = ~n9066 & n9069;
  assign n9071 = ~n9068 & n9070;
  assign n9072 = pi17  & n9071;
  assign n9073 = ~pi17  & ~n9071;
  assign n9074 = ~n9072 & ~n9073;
  assign n9075 = n9064 & ~n9074;
  assign n9076 = ~n2622 & n6608;
  assign n9077 = ~n2726 & n6140;
  assign n9078 = ~n2657 & n6356;
  assign n9079 = n6134 & n6407;
  assign n9080 = ~n9076 & ~n9078;
  assign n9081 = ~n9077 & n9080;
  assign n9082 = ~n9079 & n9081;
  assign n9083 = ~pi17  & ~n9082;
  assign n9084 = pi17  & n9082;
  assign n9085 = ~n9083 & ~n9084;
  assign n9086 = n8829 & ~n8831;
  assign n9087 = ~n8832 & ~n9086;
  assign n9088 = ~n9085 & n9087;
  assign n9089 = ~n2657 & n6608;
  assign n9090 = ~n2726 & n6356;
  assign n9091 = ~n2781 & n6140;
  assign n9092 = n6134 & n6251;
  assign n9093 = ~n9089 & ~n9091;
  assign n9094 = ~n9090 & n9093;
  assign n9095 = ~n9092 & n9094;
  assign n9096 = ~pi17  & ~n9095;
  assign n9097 = pi17  & n9095;
  assign n9098 = ~n9096 & ~n9097;
  assign n9099 = n8825 & ~n8827;
  assign n9100 = ~n8828 & ~n9099;
  assign n9101 = ~n9098 & n9100;
  assign n9102 = ~n2866 & n6140;
  assign n9103 = ~n2726 & n6608;
  assign n9104 = ~n2781 & n6356;
  assign n9105 = n6134 & n6520;
  assign n9106 = ~n9102 & ~n9104;
  assign n9107 = ~n9103 & n9106;
  assign n9108 = ~n9105 & n9107;
  assign n9109 = ~pi17  & ~n9108;
  assign n9110 = pi17  & n9108;
  assign n9111 = ~n9109 & ~n9110;
  assign n9112 = n8821 & ~n8823;
  assign n9113 = ~n8824 & ~n9112;
  assign n9114 = ~n9111 & n9113;
  assign n9115 = n8817 & ~n8819;
  assign n9116 = ~n8820 & ~n9115;
  assign n9117 = ~n2866 & n6356;
  assign n9118 = ~n2781 & n6608;
  assign n9119 = ~n2901 & n6140;
  assign n9120 = n6134 & n6819;
  assign n9121 = ~n9117 & ~n9118;
  assign n9122 = ~n9119 & n9121;
  assign n9123 = ~n9120 & n9122;
  assign n9124 = pi17  & n9123;
  assign n9125 = ~pi17  & ~n9123;
  assign n9126 = ~n9124 & ~n9125;
  assign n9127 = n9116 & ~n9126;
  assign n9128 = n8813 & ~n8815;
  assign n9129 = ~n8816 & ~n9128;
  assign n9130 = ~n2866 & n6608;
  assign n9131 = ~n2978 & n6140;
  assign n9132 = ~n2901 & n6356;
  assign n9133 = n6134 & n6831;
  assign n9134 = ~n9130 & ~n9132;
  assign n9135 = ~n9131 & n9134;
  assign n9136 = ~n9133 & n9135;
  assign n9137 = pi17  & n9136;
  assign n9138 = ~pi17  & ~n9136;
  assign n9139 = ~n9137 & ~n9138;
  assign n9140 = n9129 & ~n9139;
  assign n9141 = n8809 & ~n8811;
  assign n9142 = ~n8812 & ~n9141;
  assign n9143 = ~n2901 & n6608;
  assign n9144 = ~n2978 & n6356;
  assign n9145 = ~n3069 & n6140;
  assign n9146 = n6134 & n6496;
  assign n9147 = ~n9143 & ~n9145;
  assign n9148 = ~n9144 & n9147;
  assign n9149 = ~n9146 & n9148;
  assign n9150 = pi17  & n9149;
  assign n9151 = ~pi17  & ~n9149;
  assign n9152 = ~n9150 & ~n9151;
  assign n9153 = n9142 & ~n9152;
  assign n9154 = ~n2978 & n6608;
  assign n9155 = ~n3137 & n6140;
  assign n9156 = ~n3069 & n6356;
  assign n9157 = n6134 & n6873;
  assign n9158 = ~n9154 & ~n9156;
  assign n9159 = ~n9155 & n9158;
  assign n9160 = ~n9157 & n9159;
  assign n9161 = ~pi17  & ~n9160;
  assign n9162 = pi17  & n9160;
  assign n9163 = ~n9161 & ~n9162;
  assign n9164 = n8805 & ~n8807;
  assign n9165 = ~n8808 & ~n9164;
  assign n9166 = ~n9163 & n9165;
  assign n9167 = ~n3069 & n6608;
  assign n9168 = ~n3137 & n6356;
  assign n9169 = ~n3194 & n6140;
  assign n9170 = n6134 & n6920;
  assign n9171 = ~n9167 & ~n9169;
  assign n9172 = ~n9168 & n9171;
  assign n9173 = ~n9170 & n9172;
  assign n9174 = pi17  & n9173;
  assign n9175 = ~pi17  & ~n9173;
  assign n9176 = ~n9174 & ~n9175;
  assign n9177 = n8801 & ~n8803;
  assign n9178 = ~n8804 & ~n9177;
  assign n9179 = ~n9176 & n9178;
  assign n9180 = ~n3137 & n6608;
  assign n9181 = ~n3194 & n6356;
  assign n9182 = ~n3227 & n6140;
  assign n9183 = n6134 & n6970;
  assign n9184 = ~n9181 & ~n9182;
  assign n9185 = ~n9180 & n9184;
  assign n9186 = ~n9183 & n9185;
  assign n9187 = ~pi17  & ~n9186;
  assign n9188 = pi17  & n9186;
  assign n9189 = ~n9187 & ~n9188;
  assign n9190 = pi20  & ~n8781;
  assign n9191 = n8788 & ~n9190;
  assign n9192 = ~n8788 & n9190;
  assign n9193 = ~n9191 & ~n9192;
  assign n9194 = ~n9189 & n9193;
  assign n9195 = ~n3319 & n6140;
  assign n9196 = ~n3227 & n6356;
  assign n9197 = ~n3194 & n6608;
  assign n9198 = n6134 & n7013;
  assign n9199 = ~n9196 & ~n9197;
  assign n9200 = ~n9195 & n9199;
  assign n9201 = ~n9198 & n9200;
  assign n9202 = pi17  & n9201;
  assign n9203 = ~pi17  & ~n9201;
  assign n9204 = ~n9202 & ~n9203;
  assign n9205 = n8775 & ~n8780;
  assign n9206 = ~n8781 & ~n9205;
  assign n9207 = ~n9204 & n9206;
  assign n9208 = ~n3460 & n6130;
  assign n9209 = pi17  & n9208;
  assign n9210 = ~n3376 & n6608;
  assign n9211 = ~n3460 & n6356;
  assign n9212 = n6134 & ~n7689;
  assign n9213 = ~n9210 & ~n9211;
  assign n9214 = ~n9212 & n9213;
  assign n9215 = ~n9209 & n9214;
  assign n9216 = ~n3460 & n6140;
  assign n9217 = ~n3319 & n6608;
  assign n9218 = ~n3376 & n6356;
  assign n9219 = n6134 & n7049;
  assign n9220 = ~n9216 & ~n9218;
  assign n9221 = ~n9217 & n9220;
  assign n9222 = ~n9219 & n9221;
  assign n9223 = pi17  & n9215;
  assign n9224 = n9222 & n9223;
  assign n9225 = n8774 & n9224;
  assign n9226 = ~n3319 & n6356;
  assign n9227 = ~n3376 & n6140;
  assign n9228 = ~n3227 & n6608;
  assign n9229 = n6134 & n7105;
  assign n9230 = ~n9227 & ~n9228;
  assign n9231 = ~n9226 & n9230;
  assign n9232 = ~n9229 & n9231;
  assign n9233 = pi17  & n9232;
  assign n9234 = ~pi17  & ~n9232;
  assign n9235 = ~n9233 & ~n9234;
  assign n9236 = ~n8774 & ~n9224;
  assign n9237 = ~n9225 & ~n9236;
  assign n9238 = ~n9235 & n9237;
  assign n9239 = ~n9225 & ~n9238;
  assign n9240 = n9204 & ~n9206;
  assign n9241 = ~n9207 & ~n9240;
  assign n9242 = ~n9239 & n9241;
  assign n9243 = ~n9207 & ~n9242;
  assign n9244 = n9189 & ~n9193;
  assign n9245 = ~n9194 & ~n9244;
  assign n9246 = ~n9243 & n9245;
  assign n9247 = ~n9194 & ~n9246;
  assign n9248 = n9176 & ~n9178;
  assign n9249 = ~n9179 & ~n9248;
  assign n9250 = ~n9247 & n9249;
  assign n9251 = ~n9179 & ~n9250;
  assign n9252 = n9163 & ~n9165;
  assign n9253 = ~n9166 & ~n9252;
  assign n9254 = ~n9251 & n9253;
  assign n9255 = ~n9166 & ~n9254;
  assign n9256 = ~n9142 & n9152;
  assign n9257 = ~n9153 & ~n9256;
  assign n9258 = ~n9255 & n9257;
  assign n9259 = ~n9153 & ~n9258;
  assign n9260 = ~n9129 & n9139;
  assign n9261 = ~n9140 & ~n9260;
  assign n9262 = ~n9259 & n9261;
  assign n9263 = ~n9140 & ~n9262;
  assign n9264 = ~n9116 & n9126;
  assign n9265 = ~n9127 & ~n9264;
  assign n9266 = ~n9263 & n9265;
  assign n9267 = ~n9127 & ~n9266;
  assign n9268 = n9111 & ~n9113;
  assign n9269 = ~n9114 & ~n9268;
  assign n9270 = ~n9267 & n9269;
  assign n9271 = ~n9114 & ~n9270;
  assign n9272 = n9098 & ~n9100;
  assign n9273 = ~n9101 & ~n9272;
  assign n9274 = ~n9271 & n9273;
  assign n9275 = ~n9101 & ~n9274;
  assign n9276 = n9085 & ~n9087;
  assign n9277 = ~n9088 & ~n9276;
  assign n9278 = ~n9275 & n9277;
  assign n9279 = ~n9088 & ~n9278;
  assign n9280 = ~n9064 & n9074;
  assign n9281 = ~n9075 & ~n9280;
  assign n9282 = ~n9279 & n9281;
  assign n9283 = ~n9075 & ~n9282;
  assign n9284 = ~n9051 & n9061;
  assign n9285 = ~n9062 & ~n9284;
  assign n9286 = ~n9283 & n9285;
  assign n9287 = ~n9062 & ~n9286;
  assign n9288 = n9046 & ~n9048;
  assign n9289 = ~n9049 & ~n9288;
  assign n9290 = ~n9287 & n9289;
  assign n9291 = ~n9049 & ~n9290;
  assign n9292 = n9033 & ~n9035;
  assign n9293 = ~n9036 & ~n9292;
  assign n9294 = ~n9291 & n9293;
  assign n9295 = ~n9036 & ~n9294;
  assign n9296 = n9020 & ~n9022;
  assign n9297 = ~n9023 & ~n9296;
  assign n9298 = ~n9295 & n9297;
  assign n9299 = ~n9023 & ~n9298;
  assign n9300 = n9007 & ~n9009;
  assign n9301 = ~n9010 & ~n9300;
  assign n9302 = ~n9299 & n9301;
  assign n9303 = ~n9010 & ~n9302;
  assign n9304 = n8994 & ~n8996;
  assign n9305 = ~n8997 & ~n9304;
  assign n9306 = ~n9303 & n9305;
  assign n9307 = ~n8997 & ~n9306;
  assign n9308 = n8981 & ~n8983;
  assign n9309 = ~n8984 & ~n9308;
  assign n9310 = ~n9307 & n9309;
  assign n9311 = ~n8984 & ~n9310;
  assign n9312 = n8968 & ~n8970;
  assign n9313 = ~n8971 & ~n9312;
  assign n9314 = ~n9311 & n9313;
  assign n9315 = ~n8971 & ~n9314;
  assign n9316 = n8882 & ~n8884;
  assign n9317 = ~n8885 & ~n9316;
  assign n9318 = ~n9315 & n9317;
  assign n9319 = ~n1610 & n6653;
  assign n9320 = ~n1532 & n7243;
  assign n9321 = ~n1425 & n7380;
  assign n9322 = n4642 & n6647;
  assign n9323 = ~n9319 & ~n9320;
  assign n9324 = ~n9321 & n9323;
  assign n9325 = ~n9322 & n9324;
  assign n9326 = ~pi14  & ~n9325;
  assign n9327 = pi14  & n9325;
  assign n9328 = ~n9326 & ~n9327;
  assign n9329 = n9315 & ~n9317;
  assign n9330 = ~n9318 & ~n9329;
  assign n9331 = ~n9328 & n9330;
  assign n9332 = ~n9318 & ~n9331;
  assign n9333 = ~n8891 & n8901;
  assign n9334 = ~n8902 & ~n9333;
  assign n9335 = ~n9332 & n9334;
  assign n9336 = n9332 & ~n9334;
  assign n9337 = ~n9335 & ~n9336;
  assign n9338 = ~n1107 & n7847;
  assign n9339 = ~n1006 & n8161;
  assign n9340 = ~n1230 & n7554;
  assign n9341 = n4233 & n7548;
  assign n9342 = ~n9338 & ~n9339;
  assign n9343 = ~n9340 & n9342;
  assign n9344 = ~n9341 & n9343;
  assign n9345 = pi11  & n9344;
  assign n9346 = ~pi11  & ~n9344;
  assign n9347 = ~n9345 & ~n9346;
  assign n9348 = n9337 & ~n9347;
  assign n9349 = ~n9335 & ~n9348;
  assign n9350 = ~n8908 & n8918;
  assign n9351 = ~n8919 & ~n9350;
  assign n9352 = ~n9349 & n9351;
  assign n9353 = n9349 & ~n9351;
  assign n9354 = ~n9352 & ~n9353;
  assign n9355 = ~n8196 & n8199;
  assign n9356 = ~n621 & n9355;
  assign n9357 = ~n729 & n8939;
  assign n9358 = ~n802 & n8206;
  assign n9359 = n3955 & n8200;
  assign n9360 = ~n9356 & ~n9358;
  assign n9361 = ~n9357 & n9360;
  assign n9362 = ~n9359 & n9361;
  assign n9363 = pi8  & n9362;
  assign n9364 = ~pi8  & ~n9362;
  assign n9365 = ~n9363 & ~n9364;
  assign n9366 = n9354 & ~n9365;
  assign n9367 = ~n9352 & ~n9366;
  assign n9368 = ~n729 & n8206;
  assign n9369 = ~n621 & n8939;
  assign n9370 = ~n563 & n9355;
  assign n9371 = n3921 & n8200;
  assign n9372 = ~n9369 & ~n9370;
  assign n9373 = ~n9368 & n9372;
  assign n9374 = ~n9371 & n9373;
  assign n9375 = pi8  & n9374;
  assign n9376 = ~pi8  & ~n9374;
  assign n9377 = ~n9375 & ~n9376;
  assign n9378 = ~n9367 & ~n9377;
  assign n9379 = ~n8933 & ~n8935;
  assign n9380 = ~n8936 & ~n9379;
  assign n9381 = n9367 & n9377;
  assign n9382 = ~n9378 & ~n9381;
  assign n9383 = n9380 & n9382;
  assign n9384 = ~n9378 & ~n9383;
  assign n9385 = n8949 & ~n8951;
  assign n9386 = ~n8952 & ~n9385;
  assign n9387 = ~n9384 & n9386;
  assign n9388 = n9311 & ~n9313;
  assign n9389 = ~n9314 & ~n9388;
  assign n9390 = ~n1737 & n6653;
  assign n9391 = ~n1610 & n7243;
  assign n9392 = ~n1532 & n7380;
  assign n9393 = n4626 & n6647;
  assign n9394 = ~n9390 & ~n9391;
  assign n9395 = ~n9392 & n9394;
  assign n9396 = ~n9393 & n9395;
  assign n9397 = pi14  & n9396;
  assign n9398 = ~pi14  & ~n9396;
  assign n9399 = ~n9397 & ~n9398;
  assign n9400 = n9389 & ~n9399;
  assign n9401 = n9307 & ~n9309;
  assign n9402 = ~n9310 & ~n9401;
  assign n9403 = ~n1805 & n6653;
  assign n9404 = ~n1737 & n7243;
  assign n9405 = ~n1610 & n7380;
  assign n9406 = n4844 & n6647;
  assign n9407 = ~n9403 & ~n9404;
  assign n9408 = ~n9405 & n9407;
  assign n9409 = ~n9406 & n9408;
  assign n9410 = pi14  & n9409;
  assign n9411 = ~pi14  & ~n9409;
  assign n9412 = ~n9410 & ~n9411;
  assign n9413 = n9402 & ~n9412;
  assign n9414 = n9303 & ~n9305;
  assign n9415 = ~n9306 & ~n9414;
  assign n9416 = ~n1893 & n6653;
  assign n9417 = ~n1805 & n7243;
  assign n9418 = ~n1737 & n7380;
  assign n9419 = n4862 & n6647;
  assign n9420 = ~n9416 & ~n9417;
  assign n9421 = ~n9418 & n9420;
  assign n9422 = ~n9419 & n9421;
  assign n9423 = pi14  & n9422;
  assign n9424 = ~pi14  & ~n9422;
  assign n9425 = ~n9423 & ~n9424;
  assign n9426 = n9415 & ~n9425;
  assign n9427 = n9299 & ~n9301;
  assign n9428 = ~n9302 & ~n9427;
  assign n9429 = ~n1997 & n6653;
  assign n9430 = ~n1893 & n7243;
  assign n9431 = ~n1805 & n7380;
  assign n9432 = n5212 & n6647;
  assign n9433 = ~n9429 & ~n9430;
  assign n9434 = ~n9431 & n9433;
  assign n9435 = ~n9432 & n9434;
  assign n9436 = pi14  & n9435;
  assign n9437 = ~pi14  & ~n9435;
  assign n9438 = ~n9436 & ~n9437;
  assign n9439 = n9428 & ~n9438;
  assign n9440 = n9295 & ~n9297;
  assign n9441 = ~n9298 & ~n9440;
  assign n9442 = ~n2045 & n6653;
  assign n9443 = ~n1997 & n7243;
  assign n9444 = ~n1893 & n7380;
  assign n9445 = n5061 & n6647;
  assign n9446 = ~n9442 & ~n9443;
  assign n9447 = ~n9444 & n9446;
  assign n9448 = ~n9445 & n9447;
  assign n9449 = pi14  & n9448;
  assign n9450 = ~pi14  & ~n9448;
  assign n9451 = ~n9449 & ~n9450;
  assign n9452 = n9441 & ~n9451;
  assign n9453 = n9291 & ~n9293;
  assign n9454 = ~n9294 & ~n9453;
  assign n9455 = ~n2165 & n6653;
  assign n9456 = ~n2045 & n7243;
  assign n9457 = ~n1997 & n7380;
  assign n9458 = n5424 & n6647;
  assign n9459 = ~n9456 & ~n9457;
  assign n9460 = ~n9455 & n9459;
  assign n9461 = ~n9458 & n9460;
  assign n9462 = pi14  & n9461;
  assign n9463 = ~pi14  & ~n9461;
  assign n9464 = ~n9462 & ~n9463;
  assign n9465 = n9454 & ~n9464;
  assign n9466 = n9287 & ~n9289;
  assign n9467 = ~n9290 & ~n9466;
  assign n9468 = ~n2165 & n7243;
  assign n9469 = ~n2265 & n6653;
  assign n9470 = ~n2045 & n7380;
  assign n9471 = n5408 & n6647;
  assign n9472 = ~n9469 & ~n9470;
  assign n9473 = ~n9468 & n9472;
  assign n9474 = ~n9471 & n9473;
  assign n9475 = pi14  & n9474;
  assign n9476 = ~pi14  & ~n9474;
  assign n9477 = ~n9475 & ~n9476;
  assign n9478 = n9467 & ~n9477;
  assign n9479 = ~n2356 & n6653;
  assign n9480 = ~n2265 & n7243;
  assign n9481 = ~n2165 & n7380;
  assign n9482 = n5632 & n6647;
  assign n9483 = ~n9479 & ~n9480;
  assign n9484 = ~n9481 & n9483;
  assign n9485 = ~n9482 & n9484;
  assign n9486 = ~pi14  & ~n9485;
  assign n9487 = pi14  & n9485;
  assign n9488 = ~n9486 & ~n9487;
  assign n9489 = n9283 & ~n9285;
  assign n9490 = ~n9286 & ~n9489;
  assign n9491 = ~n9488 & n9490;
  assign n9492 = ~n2356 & n7243;
  assign n9493 = ~n2442 & n6653;
  assign n9494 = ~n2265 & n7380;
  assign n9495 = n5650 & n6647;
  assign n9496 = ~n9493 & ~n9494;
  assign n9497 = ~n9492 & n9496;
  assign n9498 = ~n9495 & n9497;
  assign n9499 = ~pi14  & ~n9498;
  assign n9500 = pi14  & n9498;
  assign n9501 = ~n9499 & ~n9500;
  assign n9502 = n9279 & ~n9281;
  assign n9503 = ~n9282 & ~n9502;
  assign n9504 = ~n9501 & n9503;
  assign n9505 = n9275 & ~n9277;
  assign n9506 = ~n9278 & ~n9505;
  assign n9507 = ~n2356 & n7380;
  assign n9508 = ~n2538 & n6653;
  assign n9509 = ~n2442 & n7243;
  assign n9510 = n6042 & n6647;
  assign n9511 = ~n9507 & ~n9509;
  assign n9512 = ~n9508 & n9511;
  assign n9513 = ~n9510 & n9512;
  assign n9514 = pi14  & n9513;
  assign n9515 = ~pi14  & ~n9513;
  assign n9516 = ~n9514 & ~n9515;
  assign n9517 = n9506 & ~n9516;
  assign n9518 = n9271 & ~n9273;
  assign n9519 = ~n9274 & ~n9518;
  assign n9520 = ~n2622 & n6653;
  assign n9521 = ~n2538 & n7243;
  assign n9522 = ~n2442 & n7380;
  assign n9523 = n5823 & n6647;
  assign n9524 = ~n9520 & ~n9522;
  assign n9525 = ~n9521 & n9524;
  assign n9526 = ~n9523 & n9525;
  assign n9527 = pi14  & n9526;
  assign n9528 = ~pi14  & ~n9526;
  assign n9529 = ~n9527 & ~n9528;
  assign n9530 = n9519 & ~n9529;
  assign n9531 = n9267 & ~n9269;
  assign n9532 = ~n9270 & ~n9531;
  assign n9533 = ~n2538 & n7380;
  assign n9534 = ~n2622 & n7243;
  assign n9535 = ~n2657 & n6653;
  assign n9536 = n6271 & n6647;
  assign n9537 = ~n9533 & ~n9535;
  assign n9538 = ~n9534 & n9537;
  assign n9539 = ~n9536 & n9538;
  assign n9540 = pi14  & n9539;
  assign n9541 = ~pi14  & ~n9539;
  assign n9542 = ~n9540 & ~n9541;
  assign n9543 = n9532 & ~n9542;
  assign n9544 = ~n2622 & n7380;
  assign n9545 = ~n2726 & n6653;
  assign n9546 = ~n2657 & n7243;
  assign n9547 = n6407 & n6647;
  assign n9548 = ~n9544 & ~n9546;
  assign n9549 = ~n9545 & n9548;
  assign n9550 = ~n9547 & n9549;
  assign n9551 = ~pi14  & ~n9550;
  assign n9552 = pi14  & n9550;
  assign n9553 = ~n9551 & ~n9552;
  assign n9554 = n9263 & ~n9265;
  assign n9555 = ~n9266 & ~n9554;
  assign n9556 = ~n9553 & n9555;
  assign n9557 = ~n2657 & n7380;
  assign n9558 = ~n2726 & n7243;
  assign n9559 = ~n2781 & n6653;
  assign n9560 = n6251 & n6647;
  assign n9561 = ~n9557 & ~n9559;
  assign n9562 = ~n9558 & n9561;
  assign n9563 = ~n9560 & n9562;
  assign n9564 = ~pi14  & ~n9563;
  assign n9565 = pi14  & n9563;
  assign n9566 = ~n9564 & ~n9565;
  assign n9567 = n9259 & ~n9261;
  assign n9568 = ~n9262 & ~n9567;
  assign n9569 = ~n9566 & n9568;
  assign n9570 = ~n2866 & n6653;
  assign n9571 = ~n2726 & n7380;
  assign n9572 = ~n2781 & n7243;
  assign n9573 = n6520 & n6647;
  assign n9574 = ~n9570 & ~n9572;
  assign n9575 = ~n9571 & n9574;
  assign n9576 = ~n9573 & n9575;
  assign n9577 = ~pi14  & ~n9576;
  assign n9578 = pi14  & n9576;
  assign n9579 = ~n9577 & ~n9578;
  assign n9580 = n9255 & ~n9257;
  assign n9581 = ~n9258 & ~n9580;
  assign n9582 = ~n9579 & n9581;
  assign n9583 = n9251 & ~n9253;
  assign n9584 = ~n9254 & ~n9583;
  assign n9585 = ~n2866 & n7243;
  assign n9586 = ~n2781 & n7380;
  assign n9587 = ~n2901 & n6653;
  assign n9588 = n6647 & n6819;
  assign n9589 = ~n9585 & ~n9586;
  assign n9590 = ~n9587 & n9589;
  assign n9591 = ~n9588 & n9590;
  assign n9592 = pi14  & n9591;
  assign n9593 = ~pi14  & ~n9591;
  assign n9594 = ~n9592 & ~n9593;
  assign n9595 = n9584 & ~n9594;
  assign n9596 = n9247 & ~n9249;
  assign n9597 = ~n9250 & ~n9596;
  assign n9598 = ~n2866 & n7380;
  assign n9599 = ~n2978 & n6653;
  assign n9600 = ~n2901 & n7243;
  assign n9601 = n6647 & n6831;
  assign n9602 = ~n9598 & ~n9600;
  assign n9603 = ~n9599 & n9602;
  assign n9604 = ~n9601 & n9603;
  assign n9605 = pi14  & n9604;
  assign n9606 = ~pi14  & ~n9604;
  assign n9607 = ~n9605 & ~n9606;
  assign n9608 = n9597 & ~n9607;
  assign n9609 = n9243 & ~n9245;
  assign n9610 = ~n9246 & ~n9609;
  assign n9611 = ~n2901 & n7380;
  assign n9612 = ~n2978 & n7243;
  assign n9613 = ~n3069 & n6653;
  assign n9614 = n6496 & n6647;
  assign n9615 = ~n9611 & ~n9613;
  assign n9616 = ~n9612 & n9615;
  assign n9617 = ~n9614 & n9616;
  assign n9618 = pi14  & n9617;
  assign n9619 = ~pi14  & ~n9617;
  assign n9620 = ~n9618 & ~n9619;
  assign n9621 = n9610 & ~n9620;
  assign n9622 = ~n2978 & n7380;
  assign n9623 = ~n3137 & n6653;
  assign n9624 = ~n3069 & n7243;
  assign n9625 = n6647 & n6873;
  assign n9626 = ~n9622 & ~n9624;
  assign n9627 = ~n9623 & n9626;
  assign n9628 = ~n9625 & n9627;
  assign n9629 = ~pi14  & ~n9628;
  assign n9630 = pi14  & n9628;
  assign n9631 = ~n9629 & ~n9630;
  assign n9632 = n9239 & ~n9241;
  assign n9633 = ~n9242 & ~n9632;
  assign n9634 = ~n9631 & n9633;
  assign n9635 = ~n3069 & n7380;
  assign n9636 = ~n3137 & n7243;
  assign n9637 = ~n3194 & n6653;
  assign n9638 = n6647 & n6920;
  assign n9639 = ~n9635 & ~n9637;
  assign n9640 = ~n9636 & n9639;
  assign n9641 = ~n9638 & n9640;
  assign n9642 = pi14  & n9641;
  assign n9643 = ~pi14  & ~n9641;
  assign n9644 = ~n9642 & ~n9643;
  assign n9645 = n9235 & ~n9237;
  assign n9646 = ~n9238 & ~n9645;
  assign n9647 = ~n9644 & n9646;
  assign n9648 = ~n3137 & n7380;
  assign n9649 = ~n3194 & n7243;
  assign n9650 = ~n3227 & n6653;
  assign n9651 = n6647 & n6970;
  assign n9652 = ~n9649 & ~n9650;
  assign n9653 = ~n9648 & n9652;
  assign n9654 = ~n9651 & n9653;
  assign n9655 = ~pi14  & ~n9654;
  assign n9656 = pi14  & n9654;
  assign n9657 = ~n9655 & ~n9656;
  assign n9658 = pi17  & ~n9215;
  assign n9659 = n9222 & ~n9658;
  assign n9660 = ~n9222 & n9658;
  assign n9661 = ~n9659 & ~n9660;
  assign n9662 = ~n9657 & n9661;
  assign n9663 = ~n3319 & n6653;
  assign n9664 = ~n3227 & n7243;
  assign n9665 = ~n3194 & n7380;
  assign n9666 = n6647 & n7013;
  assign n9667 = ~n9664 & ~n9665;
  assign n9668 = ~n9663 & n9667;
  assign n9669 = ~n9666 & n9668;
  assign n9670 = pi14  & n9669;
  assign n9671 = ~pi14  & ~n9669;
  assign n9672 = ~n9670 & ~n9671;
  assign n9673 = n9209 & ~n9214;
  assign n9674 = ~n9215 & ~n9673;
  assign n9675 = ~n9672 & n9674;
  assign n9676 = ~n3460 & n6643;
  assign n9677 = pi14  & n9676;
  assign n9678 = ~n3376 & n7380;
  assign n9679 = ~n3460 & n7243;
  assign n9680 = n6647 & ~n7689;
  assign n9681 = ~n9678 & ~n9679;
  assign n9682 = ~n9680 & n9681;
  assign n9683 = ~n9677 & n9682;
  assign n9684 = ~n3460 & n6653;
  assign n9685 = ~n3319 & n7380;
  assign n9686 = ~n3376 & n7243;
  assign n9687 = n6647 & n7049;
  assign n9688 = ~n9684 & ~n9686;
  assign n9689 = ~n9685 & n9688;
  assign n9690 = ~n9687 & n9689;
  assign n9691 = pi14  & n9683;
  assign n9692 = n9690 & n9691;
  assign n9693 = n9208 & n9692;
  assign n9694 = ~n3319 & n7243;
  assign n9695 = ~n3376 & n6653;
  assign n9696 = ~n3227 & n7380;
  assign n9697 = n6647 & n7105;
  assign n9698 = ~n9695 & ~n9696;
  assign n9699 = ~n9694 & n9698;
  assign n9700 = ~n9697 & n9699;
  assign n9701 = pi14  & n9700;
  assign n9702 = ~pi14  & ~n9700;
  assign n9703 = ~n9701 & ~n9702;
  assign n9704 = ~n9208 & ~n9692;
  assign n9705 = ~n9693 & ~n9704;
  assign n9706 = ~n9703 & n9705;
  assign n9707 = ~n9693 & ~n9706;
  assign n9708 = n9672 & ~n9674;
  assign n9709 = ~n9675 & ~n9708;
  assign n9710 = ~n9707 & n9709;
  assign n9711 = ~n9675 & ~n9710;
  assign n9712 = n9657 & ~n9661;
  assign n9713 = ~n9662 & ~n9712;
  assign n9714 = ~n9711 & n9713;
  assign n9715 = ~n9662 & ~n9714;
  assign n9716 = n9644 & ~n9646;
  assign n9717 = ~n9647 & ~n9716;
  assign n9718 = ~n9715 & n9717;
  assign n9719 = ~n9647 & ~n9718;
  assign n9720 = n9631 & ~n9633;
  assign n9721 = ~n9634 & ~n9720;
  assign n9722 = ~n9719 & n9721;
  assign n9723 = ~n9634 & ~n9722;
  assign n9724 = ~n9610 & n9620;
  assign n9725 = ~n9621 & ~n9724;
  assign n9726 = ~n9723 & n9725;
  assign n9727 = ~n9621 & ~n9726;
  assign n9728 = ~n9597 & n9607;
  assign n9729 = ~n9608 & ~n9728;
  assign n9730 = ~n9727 & n9729;
  assign n9731 = ~n9608 & ~n9730;
  assign n9732 = ~n9584 & n9594;
  assign n9733 = ~n9595 & ~n9732;
  assign n9734 = ~n9731 & n9733;
  assign n9735 = ~n9595 & ~n9734;
  assign n9736 = n9579 & ~n9581;
  assign n9737 = ~n9582 & ~n9736;
  assign n9738 = ~n9735 & n9737;
  assign n9739 = ~n9582 & ~n9738;
  assign n9740 = n9566 & ~n9568;
  assign n9741 = ~n9569 & ~n9740;
  assign n9742 = ~n9739 & n9741;
  assign n9743 = ~n9569 & ~n9742;
  assign n9744 = n9553 & ~n9555;
  assign n9745 = ~n9556 & ~n9744;
  assign n9746 = ~n9743 & n9745;
  assign n9747 = ~n9556 & ~n9746;
  assign n9748 = ~n9532 & n9542;
  assign n9749 = ~n9543 & ~n9748;
  assign n9750 = ~n9747 & n9749;
  assign n9751 = ~n9543 & ~n9750;
  assign n9752 = ~n9519 & n9529;
  assign n9753 = ~n9530 & ~n9752;
  assign n9754 = ~n9751 & n9753;
  assign n9755 = ~n9530 & ~n9754;
  assign n9756 = ~n9506 & n9516;
  assign n9757 = ~n9517 & ~n9756;
  assign n9758 = ~n9755 & n9757;
  assign n9759 = ~n9517 & ~n9758;
  assign n9760 = n9501 & ~n9503;
  assign n9761 = ~n9504 & ~n9760;
  assign n9762 = ~n9759 & n9761;
  assign n9763 = ~n9504 & ~n9762;
  assign n9764 = n9488 & ~n9490;
  assign n9765 = ~n9491 & ~n9764;
  assign n9766 = ~n9763 & n9765;
  assign n9767 = ~n9491 & ~n9766;
  assign n9768 = ~n9467 & n9477;
  assign n9769 = ~n9478 & ~n9768;
  assign n9770 = ~n9767 & n9769;
  assign n9771 = ~n9478 & ~n9770;
  assign n9772 = ~n9454 & n9464;
  assign n9773 = ~n9465 & ~n9772;
  assign n9774 = ~n9771 & n9773;
  assign n9775 = ~n9465 & ~n9774;
  assign n9776 = ~n9441 & n9451;
  assign n9777 = ~n9452 & ~n9776;
  assign n9778 = ~n9775 & n9777;
  assign n9779 = ~n9452 & ~n9778;
  assign n9780 = ~n9428 & n9438;
  assign n9781 = ~n9439 & ~n9780;
  assign n9782 = ~n9779 & n9781;
  assign n9783 = ~n9439 & ~n9782;
  assign n9784 = ~n9415 & n9425;
  assign n9785 = ~n9426 & ~n9784;
  assign n9786 = ~n9783 & n9785;
  assign n9787 = ~n9426 & ~n9786;
  assign n9788 = ~n9402 & n9412;
  assign n9789 = ~n9413 & ~n9788;
  assign n9790 = ~n9787 & n9789;
  assign n9791 = ~n9413 & ~n9790;
  assign n9792 = ~n9389 & n9399;
  assign n9793 = ~n9400 & ~n9792;
  assign n9794 = ~n9791 & n9793;
  assign n9795 = ~n9400 & ~n9794;
  assign n9796 = n9328 & ~n9330;
  assign n9797 = ~n9331 & ~n9796;
  assign n9798 = ~n9795 & n9797;
  assign n9799 = ~n1337 & n7554;
  assign n9800 = ~n1230 & n7847;
  assign n9801 = ~n1107 & n8161;
  assign n9802 = n4251 & n7548;
  assign n9803 = ~n9799 & ~n9800;
  assign n9804 = ~n9801 & n9803;
  assign n9805 = ~n9802 & n9804;
  assign n9806 = ~pi11  & ~n9805;
  assign n9807 = pi11  & n9805;
  assign n9808 = ~n9806 & ~n9807;
  assign n9809 = n9795 & ~n9797;
  assign n9810 = ~n9798 & ~n9809;
  assign n9811 = ~n9808 & n9810;
  assign n9812 = ~n9798 & ~n9811;
  assign n9813 = ~n9337 & n9347;
  assign n9814 = ~n9348 & ~n9813;
  assign n9815 = ~n9812 & n9814;
  assign n9816 = n9812 & ~n9814;
  assign n9817 = ~n9815 & ~n9816;
  assign n9818 = ~n729 & n9355;
  assign n9819 = ~n802 & n8939;
  assign n9820 = ~n898 & n8206;
  assign n9821 = n3901 & n8200;
  assign n9822 = ~n9819 & ~n9820;
  assign n9823 = ~n9818 & n9822;
  assign n9824 = ~n9821 & n9823;
  assign n9825 = pi8  & n9824;
  assign n9826 = ~pi8  & ~n9824;
  assign n9827 = ~n9825 & ~n9826;
  assign n9828 = n9817 & ~n9827;
  assign n9829 = ~n9815 & ~n9828;
  assign n9830 = n67 & n70;
  assign n9831 = ~n3593 & n9830;
  assign n9832 = ~pi3  & ~pi4 ;
  assign n9833 = pi3  & pi4 ;
  assign n9834 = ~n9832 & ~n9833;
  assign n9835 = ~n67 & n70;
  assign n9836 = ~n9834 & n9835;
  assign n9837 = ~n9831 & ~n9836;
  assign n9838 = ~n563 & ~n9837;
  assign n9839 = pi5  & ~n9838;
  assign n9840 = ~pi5  & n9838;
  assign n9841 = ~n9839 & ~n9840;
  assign n9842 = ~n9829 & ~n9841;
  assign n9843 = n9829 & n9841;
  assign n9844 = ~n9842 & ~n9843;
  assign n9845 = ~n9354 & n9365;
  assign n9846 = ~n9366 & ~n9845;
  assign n9847 = n9844 & n9846;
  assign n9848 = ~n9842 & ~n9847;
  assign n9849 = ~n9380 & ~n9382;
  assign n9850 = ~n9383 & ~n9849;
  assign n9851 = ~n9848 & n9850;
  assign n9852 = ~n1425 & n7554;
  assign n9853 = ~n1337 & n7847;
  assign n9854 = ~n1230 & n8161;
  assign n9855 = n4549 & n7548;
  assign n9856 = ~n9852 & ~n9853;
  assign n9857 = ~n9854 & n9856;
  assign n9858 = ~n9855 & n9857;
  assign n9859 = ~pi11  & ~n9858;
  assign n9860 = pi11  & n9858;
  assign n9861 = ~n9859 & ~n9860;
  assign n9862 = n9791 & ~n9793;
  assign n9863 = ~n9794 & ~n9862;
  assign n9864 = ~n9861 & n9863;
  assign n9865 = ~n1532 & n7554;
  assign n9866 = ~n1425 & n7847;
  assign n9867 = ~n1337 & n8161;
  assign n9868 = n4452 & n7548;
  assign n9869 = ~n9865 & ~n9866;
  assign n9870 = ~n9867 & n9869;
  assign n9871 = ~n9868 & n9870;
  assign n9872 = ~pi11  & ~n9871;
  assign n9873 = pi11  & n9871;
  assign n9874 = ~n9872 & ~n9873;
  assign n9875 = n9787 & ~n9789;
  assign n9876 = ~n9790 & ~n9875;
  assign n9877 = ~n9874 & n9876;
  assign n9878 = ~n1610 & n7554;
  assign n9879 = ~n1532 & n7847;
  assign n9880 = ~n1425 & n8161;
  assign n9881 = n4642 & n7548;
  assign n9882 = ~n9878 & ~n9879;
  assign n9883 = ~n9880 & n9882;
  assign n9884 = ~n9881 & n9883;
  assign n9885 = ~pi11  & ~n9884;
  assign n9886 = pi11  & n9884;
  assign n9887 = ~n9885 & ~n9886;
  assign n9888 = n9783 & ~n9785;
  assign n9889 = ~n9786 & ~n9888;
  assign n9890 = ~n9887 & n9889;
  assign n9891 = ~n1737 & n7554;
  assign n9892 = ~n1610 & n7847;
  assign n9893 = ~n1532 & n8161;
  assign n9894 = n4626 & n7548;
  assign n9895 = ~n9891 & ~n9892;
  assign n9896 = ~n9893 & n9895;
  assign n9897 = ~n9894 & n9896;
  assign n9898 = ~pi11  & ~n9897;
  assign n9899 = pi11  & n9897;
  assign n9900 = ~n9898 & ~n9899;
  assign n9901 = n9779 & ~n9781;
  assign n9902 = ~n9782 & ~n9901;
  assign n9903 = ~n9900 & n9902;
  assign n9904 = ~n1805 & n7554;
  assign n9905 = ~n1737 & n7847;
  assign n9906 = ~n1610 & n8161;
  assign n9907 = n4844 & n7548;
  assign n9908 = ~n9904 & ~n9905;
  assign n9909 = ~n9906 & n9908;
  assign n9910 = ~n9907 & n9909;
  assign n9911 = ~pi11  & ~n9910;
  assign n9912 = pi11  & n9910;
  assign n9913 = ~n9911 & ~n9912;
  assign n9914 = n9775 & ~n9777;
  assign n9915 = ~n9778 & ~n9914;
  assign n9916 = ~n9913 & n9915;
  assign n9917 = ~n1893 & n7554;
  assign n9918 = ~n1805 & n7847;
  assign n9919 = ~n1737 & n8161;
  assign n9920 = n4862 & n7548;
  assign n9921 = ~n9917 & ~n9918;
  assign n9922 = ~n9919 & n9921;
  assign n9923 = ~n9920 & n9922;
  assign n9924 = ~pi11  & ~n9923;
  assign n9925 = pi11  & n9923;
  assign n9926 = ~n9924 & ~n9925;
  assign n9927 = n9771 & ~n9773;
  assign n9928 = ~n9774 & ~n9927;
  assign n9929 = ~n9926 & n9928;
  assign n9930 = ~n1997 & n7554;
  assign n9931 = ~n1893 & n7847;
  assign n9932 = ~n1805 & n8161;
  assign n9933 = n5212 & n7548;
  assign n9934 = ~n9930 & ~n9931;
  assign n9935 = ~n9932 & n9934;
  assign n9936 = ~n9933 & n9935;
  assign n9937 = ~pi11  & ~n9936;
  assign n9938 = pi11  & n9936;
  assign n9939 = ~n9937 & ~n9938;
  assign n9940 = n9767 & ~n9769;
  assign n9941 = ~n9770 & ~n9940;
  assign n9942 = ~n9939 & n9941;
  assign n9943 = n9763 & ~n9765;
  assign n9944 = ~n9766 & ~n9943;
  assign n9945 = ~n2045 & n7554;
  assign n9946 = ~n1997 & n7847;
  assign n9947 = ~n1893 & n8161;
  assign n9948 = n5061 & n7548;
  assign n9949 = ~n9945 & ~n9946;
  assign n9950 = ~n9947 & n9949;
  assign n9951 = ~n9948 & n9950;
  assign n9952 = pi11  & n9951;
  assign n9953 = ~pi11  & ~n9951;
  assign n9954 = ~n9952 & ~n9953;
  assign n9955 = n9944 & ~n9954;
  assign n9956 = n9759 & ~n9761;
  assign n9957 = ~n9762 & ~n9956;
  assign n9958 = ~n2165 & n7554;
  assign n9959 = ~n2045 & n7847;
  assign n9960 = ~n1997 & n8161;
  assign n9961 = n5424 & n7548;
  assign n9962 = ~n9959 & ~n9960;
  assign n9963 = ~n9958 & n9962;
  assign n9964 = ~n9961 & n9963;
  assign n9965 = pi11  & n9964;
  assign n9966 = ~pi11  & ~n9964;
  assign n9967 = ~n9965 & ~n9966;
  assign n9968 = n9957 & ~n9967;
  assign n9969 = ~n2165 & n7847;
  assign n9970 = ~n2265 & n7554;
  assign n9971 = ~n2045 & n8161;
  assign n9972 = n5408 & n7548;
  assign n9973 = ~n9970 & ~n9971;
  assign n9974 = ~n9969 & n9973;
  assign n9975 = ~n9972 & n9974;
  assign n9976 = ~pi11  & ~n9975;
  assign n9977 = pi11  & n9975;
  assign n9978 = ~n9976 & ~n9977;
  assign n9979 = n9755 & ~n9757;
  assign n9980 = ~n9758 & ~n9979;
  assign n9981 = ~n9978 & n9980;
  assign n9982 = ~n2356 & n7554;
  assign n9983 = ~n2265 & n7847;
  assign n9984 = ~n2165 & n8161;
  assign n9985 = n5632 & n7548;
  assign n9986 = ~n9982 & ~n9983;
  assign n9987 = ~n9984 & n9986;
  assign n9988 = ~n9985 & n9987;
  assign n9989 = ~pi11  & ~n9988;
  assign n9990 = pi11  & n9988;
  assign n9991 = ~n9989 & ~n9990;
  assign n9992 = n9751 & ~n9753;
  assign n9993 = ~n9754 & ~n9992;
  assign n9994 = ~n9991 & n9993;
  assign n9995 = ~n2356 & n7847;
  assign n9996 = ~n2442 & n7554;
  assign n9997 = ~n2265 & n8161;
  assign n9998 = n5650 & n7548;
  assign n9999 = ~n9996 & ~n9997;
  assign n10000 = ~n9995 & n9999;
  assign n10001 = ~n9998 & n10000;
  assign n10002 = ~pi11  & ~n10001;
  assign n10003 = pi11  & n10001;
  assign n10004 = ~n10002 & ~n10003;
  assign n10005 = n9747 & ~n9749;
  assign n10006 = ~n9750 & ~n10005;
  assign n10007 = ~n10004 & n10006;
  assign n10008 = n9743 & ~n9745;
  assign n10009 = ~n9746 & ~n10008;
  assign n10010 = ~n2356 & n8161;
  assign n10011 = ~n2538 & n7554;
  assign n10012 = ~n2442 & n7847;
  assign n10013 = n6042 & n7548;
  assign n10014 = ~n10010 & ~n10012;
  assign n10015 = ~n10011 & n10014;
  assign n10016 = ~n10013 & n10015;
  assign n10017 = pi11  & n10016;
  assign n10018 = ~pi11  & ~n10016;
  assign n10019 = ~n10017 & ~n10018;
  assign n10020 = n10009 & ~n10019;
  assign n10021 = n9739 & ~n9741;
  assign n10022 = ~n9742 & ~n10021;
  assign n10023 = ~n2622 & n7554;
  assign n10024 = ~n2538 & n7847;
  assign n10025 = ~n2442 & n8161;
  assign n10026 = n5823 & n7548;
  assign n10027 = ~n10023 & ~n10025;
  assign n10028 = ~n10024 & n10027;
  assign n10029 = ~n10026 & n10028;
  assign n10030 = pi11  & n10029;
  assign n10031 = ~pi11  & ~n10029;
  assign n10032 = ~n10030 & ~n10031;
  assign n10033 = n10022 & ~n10032;
  assign n10034 = n9735 & ~n9737;
  assign n10035 = ~n9738 & ~n10034;
  assign n10036 = ~n2538 & n8161;
  assign n10037 = ~n2622 & n7847;
  assign n10038 = ~n2657 & n7554;
  assign n10039 = n6271 & n7548;
  assign n10040 = ~n10036 & ~n10038;
  assign n10041 = ~n10037 & n10040;
  assign n10042 = ~n10039 & n10041;
  assign n10043 = pi11  & n10042;
  assign n10044 = ~pi11  & ~n10042;
  assign n10045 = ~n10043 & ~n10044;
  assign n10046 = n10035 & ~n10045;
  assign n10047 = ~n2622 & n8161;
  assign n10048 = ~n2726 & n7554;
  assign n10049 = ~n2657 & n7847;
  assign n10050 = n6407 & n7548;
  assign n10051 = ~n10047 & ~n10049;
  assign n10052 = ~n10048 & n10051;
  assign n10053 = ~n10050 & n10052;
  assign n10054 = ~pi11  & ~n10053;
  assign n10055 = pi11  & n10053;
  assign n10056 = ~n10054 & ~n10055;
  assign n10057 = n9731 & ~n9733;
  assign n10058 = ~n9734 & ~n10057;
  assign n10059 = ~n10056 & n10058;
  assign n10060 = ~n2657 & n8161;
  assign n10061 = ~n2726 & n7847;
  assign n10062 = ~n2781 & n7554;
  assign n10063 = n6251 & n7548;
  assign n10064 = ~n10060 & ~n10062;
  assign n10065 = ~n10061 & n10064;
  assign n10066 = ~n10063 & n10065;
  assign n10067 = ~pi11  & ~n10066;
  assign n10068 = pi11  & n10066;
  assign n10069 = ~n10067 & ~n10068;
  assign n10070 = n9727 & ~n9729;
  assign n10071 = ~n9730 & ~n10070;
  assign n10072 = ~n10069 & n10071;
  assign n10073 = ~n2866 & n7554;
  assign n10074 = ~n2726 & n8161;
  assign n10075 = ~n2781 & n7847;
  assign n10076 = n6520 & n7548;
  assign n10077 = ~n10073 & ~n10075;
  assign n10078 = ~n10074 & n10077;
  assign n10079 = ~n10076 & n10078;
  assign n10080 = ~pi11  & ~n10079;
  assign n10081 = pi11  & n10079;
  assign n10082 = ~n10080 & ~n10081;
  assign n10083 = n9723 & ~n9725;
  assign n10084 = ~n9726 & ~n10083;
  assign n10085 = ~n10082 & n10084;
  assign n10086 = n9719 & ~n9721;
  assign n10087 = ~n9722 & ~n10086;
  assign n10088 = ~n2866 & n7847;
  assign n10089 = ~n2781 & n8161;
  assign n10090 = ~n2901 & n7554;
  assign n10091 = n6819 & n7548;
  assign n10092 = ~n10088 & ~n10089;
  assign n10093 = ~n10090 & n10092;
  assign n10094 = ~n10091 & n10093;
  assign n10095 = pi11  & n10094;
  assign n10096 = ~pi11  & ~n10094;
  assign n10097 = ~n10095 & ~n10096;
  assign n10098 = n10087 & ~n10097;
  assign n10099 = n9715 & ~n9717;
  assign n10100 = ~n9718 & ~n10099;
  assign n10101 = ~n2866 & n8161;
  assign n10102 = ~n2978 & n7554;
  assign n10103 = ~n2901 & n7847;
  assign n10104 = n6831 & n7548;
  assign n10105 = ~n10101 & ~n10103;
  assign n10106 = ~n10102 & n10105;
  assign n10107 = ~n10104 & n10106;
  assign n10108 = pi11  & n10107;
  assign n10109 = ~pi11  & ~n10107;
  assign n10110 = ~n10108 & ~n10109;
  assign n10111 = n10100 & ~n10110;
  assign n10112 = n9711 & ~n9713;
  assign n10113 = ~n9714 & ~n10112;
  assign n10114 = ~n2901 & n8161;
  assign n10115 = ~n2978 & n7847;
  assign n10116 = ~n3069 & n7554;
  assign n10117 = n6496 & n7548;
  assign n10118 = ~n10114 & ~n10116;
  assign n10119 = ~n10115 & n10118;
  assign n10120 = ~n10117 & n10119;
  assign n10121 = pi11  & n10120;
  assign n10122 = ~pi11  & ~n10120;
  assign n10123 = ~n10121 & ~n10122;
  assign n10124 = n10113 & ~n10123;
  assign n10125 = ~n2978 & n8161;
  assign n10126 = ~n3137 & n7554;
  assign n10127 = ~n3069 & n7847;
  assign n10128 = n6873 & n7548;
  assign n10129 = ~n10125 & ~n10127;
  assign n10130 = ~n10126 & n10129;
  assign n10131 = ~n10128 & n10130;
  assign n10132 = ~pi11  & ~n10131;
  assign n10133 = pi11  & n10131;
  assign n10134 = ~n10132 & ~n10133;
  assign n10135 = n9707 & ~n9709;
  assign n10136 = ~n9710 & ~n10135;
  assign n10137 = ~n10134 & n10136;
  assign n10138 = ~n3069 & n8161;
  assign n10139 = ~n3137 & n7847;
  assign n10140 = ~n3194 & n7554;
  assign n10141 = n6920 & n7548;
  assign n10142 = ~n10138 & ~n10140;
  assign n10143 = ~n10139 & n10142;
  assign n10144 = ~n10141 & n10143;
  assign n10145 = pi11  & n10144;
  assign n10146 = ~pi11  & ~n10144;
  assign n10147 = ~n10145 & ~n10146;
  assign n10148 = n9703 & ~n9705;
  assign n10149 = ~n9706 & ~n10148;
  assign n10150 = ~n10147 & n10149;
  assign n10151 = ~n3137 & n8161;
  assign n10152 = ~n3194 & n7847;
  assign n10153 = ~n3227 & n7554;
  assign n10154 = n6970 & n7548;
  assign n10155 = ~n10152 & ~n10153;
  assign n10156 = ~n10151 & n10155;
  assign n10157 = ~n10154 & n10156;
  assign n10158 = ~pi11  & ~n10157;
  assign n10159 = pi11  & n10157;
  assign n10160 = ~n10158 & ~n10159;
  assign n10161 = pi14  & ~n9683;
  assign n10162 = n9690 & ~n10161;
  assign n10163 = ~n9690 & n10161;
  assign n10164 = ~n10162 & ~n10163;
  assign n10165 = ~n10160 & n10164;
  assign n10166 = ~n3319 & n7554;
  assign n10167 = ~n3227 & n7847;
  assign n10168 = ~n3194 & n8161;
  assign n10169 = n7013 & n7548;
  assign n10170 = ~n10167 & ~n10168;
  assign n10171 = ~n10166 & n10170;
  assign n10172 = ~n10169 & n10171;
  assign n10173 = pi11  & n10172;
  assign n10174 = ~pi11  & ~n10172;
  assign n10175 = ~n10173 & ~n10174;
  assign n10176 = n9677 & ~n9682;
  assign n10177 = ~n9683 & ~n10176;
  assign n10178 = ~n10175 & n10177;
  assign n10179 = ~n3460 & n7547;
  assign n10180 = pi11  & n10179;
  assign n10181 = ~n3376 & n8161;
  assign n10182 = ~n3460 & n7847;
  assign n10183 = n7548 & ~n7689;
  assign n10184 = ~n10181 & ~n10182;
  assign n10185 = ~n10183 & n10184;
  assign n10186 = ~n10180 & n10185;
  assign n10187 = ~n3460 & n7554;
  assign n10188 = ~n3319 & n8161;
  assign n10189 = ~n3376 & n7847;
  assign n10190 = n7049 & n7548;
  assign n10191 = ~n10187 & ~n10189;
  assign n10192 = ~n10188 & n10191;
  assign n10193 = ~n10190 & n10192;
  assign n10194 = pi11  & n10186;
  assign n10195 = n10193 & n10194;
  assign n10196 = n9676 & n10195;
  assign n10197 = ~n3319 & n7847;
  assign n10198 = ~n3376 & n7554;
  assign n10199 = ~n3227 & n8161;
  assign n10200 = n7105 & n7548;
  assign n10201 = ~n10198 & ~n10199;
  assign n10202 = ~n10197 & n10201;
  assign n10203 = ~n10200 & n10202;
  assign n10204 = pi11  & n10203;
  assign n10205 = ~pi11  & ~n10203;
  assign n10206 = ~n10204 & ~n10205;
  assign n10207 = ~n9676 & ~n10195;
  assign n10208 = ~n10196 & ~n10207;
  assign n10209 = ~n10206 & n10208;
  assign n10210 = ~n10196 & ~n10209;
  assign n10211 = n10175 & ~n10177;
  assign n10212 = ~n10178 & ~n10211;
  assign n10213 = ~n10210 & n10212;
  assign n10214 = ~n10178 & ~n10213;
  assign n10215 = n10160 & ~n10164;
  assign n10216 = ~n10165 & ~n10215;
  assign n10217 = ~n10214 & n10216;
  assign n10218 = ~n10165 & ~n10217;
  assign n10219 = n10147 & ~n10149;
  assign n10220 = ~n10150 & ~n10219;
  assign n10221 = ~n10218 & n10220;
  assign n10222 = ~n10150 & ~n10221;
  assign n10223 = n10134 & ~n10136;
  assign n10224 = ~n10137 & ~n10223;
  assign n10225 = ~n10222 & n10224;
  assign n10226 = ~n10137 & ~n10225;
  assign n10227 = ~n10113 & n10123;
  assign n10228 = ~n10124 & ~n10227;
  assign n10229 = ~n10226 & n10228;
  assign n10230 = ~n10124 & ~n10229;
  assign n10231 = ~n10100 & n10110;
  assign n10232 = ~n10111 & ~n10231;
  assign n10233 = ~n10230 & n10232;
  assign n10234 = ~n10111 & ~n10233;
  assign n10235 = ~n10087 & n10097;
  assign n10236 = ~n10098 & ~n10235;
  assign n10237 = ~n10234 & n10236;
  assign n10238 = ~n10098 & ~n10237;
  assign n10239 = n10082 & ~n10084;
  assign n10240 = ~n10085 & ~n10239;
  assign n10241 = ~n10238 & n10240;
  assign n10242 = ~n10085 & ~n10241;
  assign n10243 = n10069 & ~n10071;
  assign n10244 = ~n10072 & ~n10243;
  assign n10245 = ~n10242 & n10244;
  assign n10246 = ~n10072 & ~n10245;
  assign n10247 = n10056 & ~n10058;
  assign n10248 = ~n10059 & ~n10247;
  assign n10249 = ~n10246 & n10248;
  assign n10250 = ~n10059 & ~n10249;
  assign n10251 = ~n10035 & n10045;
  assign n10252 = ~n10046 & ~n10251;
  assign n10253 = ~n10250 & n10252;
  assign n10254 = ~n10046 & ~n10253;
  assign n10255 = ~n10022 & n10032;
  assign n10256 = ~n10033 & ~n10255;
  assign n10257 = ~n10254 & n10256;
  assign n10258 = ~n10033 & ~n10257;
  assign n10259 = ~n10009 & n10019;
  assign n10260 = ~n10020 & ~n10259;
  assign n10261 = ~n10258 & n10260;
  assign n10262 = ~n10020 & ~n10261;
  assign n10263 = n10004 & ~n10006;
  assign n10264 = ~n10007 & ~n10263;
  assign n10265 = ~n10262 & n10264;
  assign n10266 = ~n10007 & ~n10265;
  assign n10267 = n9991 & ~n9993;
  assign n10268 = ~n9994 & ~n10267;
  assign n10269 = ~n10266 & n10268;
  assign n10270 = ~n9994 & ~n10269;
  assign n10271 = n9978 & ~n9980;
  assign n10272 = ~n9981 & ~n10271;
  assign n10273 = ~n10270 & n10272;
  assign n10274 = ~n9981 & ~n10273;
  assign n10275 = ~n9957 & n9967;
  assign n10276 = ~n9968 & ~n10275;
  assign n10277 = ~n10274 & n10276;
  assign n10278 = ~n9968 & ~n10277;
  assign n10279 = ~n9944 & n9954;
  assign n10280 = ~n9955 & ~n10279;
  assign n10281 = ~n10278 & n10280;
  assign n10282 = ~n9955 & ~n10281;
  assign n10283 = n9939 & ~n9941;
  assign n10284 = ~n9942 & ~n10283;
  assign n10285 = ~n10282 & n10284;
  assign n10286 = ~n9942 & ~n10285;
  assign n10287 = n9926 & ~n9928;
  assign n10288 = ~n9929 & ~n10287;
  assign n10289 = ~n10286 & n10288;
  assign n10290 = ~n9929 & ~n10289;
  assign n10291 = n9913 & ~n9915;
  assign n10292 = ~n9916 & ~n10291;
  assign n10293 = ~n10290 & n10292;
  assign n10294 = ~n9916 & ~n10293;
  assign n10295 = n9900 & ~n9902;
  assign n10296 = ~n9903 & ~n10295;
  assign n10297 = ~n10294 & n10296;
  assign n10298 = ~n9903 & ~n10297;
  assign n10299 = n9887 & ~n9889;
  assign n10300 = ~n9890 & ~n10299;
  assign n10301 = ~n10298 & n10300;
  assign n10302 = ~n9890 & ~n10301;
  assign n10303 = n9874 & ~n9876;
  assign n10304 = ~n9877 & ~n10303;
  assign n10305 = ~n10302 & n10304;
  assign n10306 = ~n9877 & ~n10305;
  assign n10307 = n9861 & ~n9863;
  assign n10308 = ~n9864 & ~n10307;
  assign n10309 = ~n10306 & n10308;
  assign n10310 = ~n9864 & ~n10309;
  assign n10311 = n9808 & ~n9810;
  assign n10312 = ~n9811 & ~n10311;
  assign n10313 = ~n10310 & n10312;
  assign n10314 = ~n802 & n9355;
  assign n10315 = ~n898 & n8939;
  assign n10316 = ~n1006 & n8206;
  assign n10317 = n4057 & n8200;
  assign n10318 = ~n10314 & ~n10315;
  assign n10319 = ~n10316 & n10318;
  assign n10320 = ~n10317 & n10319;
  assign n10321 = ~pi8  & ~n10320;
  assign n10322 = pi8  & n10320;
  assign n10323 = ~n10321 & ~n10322;
  assign n10324 = n10310 & ~n10312;
  assign n10325 = ~n10313 & ~n10324;
  assign n10326 = ~n10323 & n10325;
  assign n10327 = ~n10313 & ~n10326;
  assign n10328 = ~n621 & n9836;
  assign n10329 = ~n67 & n9834;
  assign n10330 = ~n563 & n10329;
  assign n10331 = n3687 & n9830;
  assign n10332 = ~n10328 & ~n10330;
  assign n10333 = ~n10331 & n10332;
  assign n10334 = pi5  & n10333;
  assign n10335 = ~pi5  & ~n10333;
  assign n10336 = ~n10334 & ~n10335;
  assign n10337 = ~n10327 & ~n10336;
  assign n10338 = n10327 & n10336;
  assign n10339 = ~n10337 & ~n10338;
  assign n10340 = ~n9817 & n9827;
  assign n10341 = ~n9828 & ~n10340;
  assign n10342 = n10339 & n10341;
  assign n10343 = ~n10337 & ~n10342;
  assign n10344 = ~n9844 & ~n9846;
  assign n10345 = ~n9847 & ~n10344;
  assign n10346 = ~n10343 & n10345;
  assign n10347 = n10343 & ~n10345;
  assign n10348 = ~n10346 & ~n10347;
  assign n10349 = n10306 & ~n10308;
  assign n10350 = ~n10309 & ~n10349;
  assign n10351 = ~n898 & n9355;
  assign n10352 = ~n1006 & n8939;
  assign n10353 = ~n1107 & n8206;
  assign n10354 = n4041 & n8200;
  assign n10355 = ~n10351 & ~n10352;
  assign n10356 = ~n10353 & n10355;
  assign n10357 = ~n10354 & n10356;
  assign n10358 = pi8  & n10357;
  assign n10359 = ~pi8  & ~n10357;
  assign n10360 = ~n10358 & ~n10359;
  assign n10361 = n10350 & ~n10360;
  assign n10362 = n10302 & ~n10304;
  assign n10363 = ~n10305 & ~n10362;
  assign n10364 = ~n1107 & n8939;
  assign n10365 = ~n1006 & n9355;
  assign n10366 = ~n1230 & n8206;
  assign n10367 = n4233 & n8200;
  assign n10368 = ~n10364 & ~n10365;
  assign n10369 = ~n10366 & n10368;
  assign n10370 = ~n10367 & n10369;
  assign n10371 = pi8  & n10370;
  assign n10372 = ~pi8  & ~n10370;
  assign n10373 = ~n10371 & ~n10372;
  assign n10374 = n10363 & ~n10373;
  assign n10375 = n10298 & ~n10300;
  assign n10376 = ~n10301 & ~n10375;
  assign n10377 = ~n1337 & n8206;
  assign n10378 = ~n1230 & n8939;
  assign n10379 = ~n1107 & n9355;
  assign n10380 = n4251 & n8200;
  assign n10381 = ~n10377 & ~n10378;
  assign n10382 = ~n10379 & n10381;
  assign n10383 = ~n10380 & n10382;
  assign n10384 = pi8  & n10383;
  assign n10385 = ~pi8  & ~n10383;
  assign n10386 = ~n10384 & ~n10385;
  assign n10387 = n10376 & ~n10386;
  assign n10388 = n10294 & ~n10296;
  assign n10389 = ~n10297 & ~n10388;
  assign n10390 = ~n1425 & n8206;
  assign n10391 = ~n1337 & n8939;
  assign n10392 = ~n1230 & n9355;
  assign n10393 = n4549 & n8200;
  assign n10394 = ~n10390 & ~n10391;
  assign n10395 = ~n10392 & n10394;
  assign n10396 = ~n10393 & n10395;
  assign n10397 = pi8  & n10396;
  assign n10398 = ~pi8  & ~n10396;
  assign n10399 = ~n10397 & ~n10398;
  assign n10400 = n10389 & ~n10399;
  assign n10401 = n10290 & ~n10292;
  assign n10402 = ~n10293 & ~n10401;
  assign n10403 = ~n1532 & n8206;
  assign n10404 = ~n1425 & n8939;
  assign n10405 = ~n1337 & n9355;
  assign n10406 = n4452 & n8200;
  assign n10407 = ~n10403 & ~n10404;
  assign n10408 = ~n10405 & n10407;
  assign n10409 = ~n10406 & n10408;
  assign n10410 = pi8  & n10409;
  assign n10411 = ~pi8  & ~n10409;
  assign n10412 = ~n10410 & ~n10411;
  assign n10413 = n10402 & ~n10412;
  assign n10414 = n10286 & ~n10288;
  assign n10415 = ~n10289 & ~n10414;
  assign n10416 = ~n1610 & n8206;
  assign n10417 = ~n1532 & n8939;
  assign n10418 = ~n1425 & n9355;
  assign n10419 = n4642 & n8200;
  assign n10420 = ~n10416 & ~n10417;
  assign n10421 = ~n10418 & n10420;
  assign n10422 = ~n10419 & n10421;
  assign n10423 = pi8  & n10422;
  assign n10424 = ~pi8  & ~n10422;
  assign n10425 = ~n10423 & ~n10424;
  assign n10426 = n10415 & ~n10425;
  assign n10427 = n10282 & ~n10284;
  assign n10428 = ~n10285 & ~n10427;
  assign n10429 = ~n1737 & n8206;
  assign n10430 = ~n1610 & n8939;
  assign n10431 = ~n1532 & n9355;
  assign n10432 = n4626 & n8200;
  assign n10433 = ~n10429 & ~n10430;
  assign n10434 = ~n10431 & n10433;
  assign n10435 = ~n10432 & n10434;
  assign n10436 = pi8  & n10435;
  assign n10437 = ~pi8  & ~n10435;
  assign n10438 = ~n10436 & ~n10437;
  assign n10439 = n10428 & ~n10438;
  assign n10440 = ~n1805 & n8206;
  assign n10441 = ~n1737 & n8939;
  assign n10442 = ~n1610 & n9355;
  assign n10443 = n4844 & n8200;
  assign n10444 = ~n10440 & ~n10441;
  assign n10445 = ~n10442 & n10444;
  assign n10446 = ~n10443 & n10445;
  assign n10447 = ~pi8  & ~n10446;
  assign n10448 = pi8  & n10446;
  assign n10449 = ~n10447 & ~n10448;
  assign n10450 = n10278 & ~n10280;
  assign n10451 = ~n10281 & ~n10450;
  assign n10452 = ~n10449 & n10451;
  assign n10453 = ~n1893 & n8206;
  assign n10454 = ~n1805 & n8939;
  assign n10455 = ~n1737 & n9355;
  assign n10456 = n4862 & n8200;
  assign n10457 = ~n10453 & ~n10454;
  assign n10458 = ~n10455 & n10457;
  assign n10459 = ~n10456 & n10458;
  assign n10460 = ~pi8  & ~n10459;
  assign n10461 = pi8  & n10459;
  assign n10462 = ~n10460 & ~n10461;
  assign n10463 = n10274 & ~n10276;
  assign n10464 = ~n10277 & ~n10463;
  assign n10465 = ~n10462 & n10464;
  assign n10466 = n10270 & ~n10272;
  assign n10467 = ~n10273 & ~n10466;
  assign n10468 = ~n1997 & n8206;
  assign n10469 = ~n1893 & n8939;
  assign n10470 = ~n1805 & n9355;
  assign n10471 = n5212 & n8200;
  assign n10472 = ~n10468 & ~n10469;
  assign n10473 = ~n10470 & n10472;
  assign n10474 = ~n10471 & n10473;
  assign n10475 = pi8  & n10474;
  assign n10476 = ~pi8  & ~n10474;
  assign n10477 = ~n10475 & ~n10476;
  assign n10478 = n10467 & ~n10477;
  assign n10479 = n10266 & ~n10268;
  assign n10480 = ~n10269 & ~n10479;
  assign n10481 = ~n2045 & n8206;
  assign n10482 = ~n1997 & n8939;
  assign n10483 = ~n1893 & n9355;
  assign n10484 = n5061 & n8200;
  assign n10485 = ~n10481 & ~n10482;
  assign n10486 = ~n10483 & n10485;
  assign n10487 = ~n10484 & n10486;
  assign n10488 = pi8  & n10487;
  assign n10489 = ~pi8  & ~n10487;
  assign n10490 = ~n10488 & ~n10489;
  assign n10491 = n10480 & ~n10490;
  assign n10492 = n10262 & ~n10264;
  assign n10493 = ~n10265 & ~n10492;
  assign n10494 = ~n2165 & n8206;
  assign n10495 = ~n2045 & n8939;
  assign n10496 = ~n1997 & n9355;
  assign n10497 = n5424 & n8200;
  assign n10498 = ~n10495 & ~n10496;
  assign n10499 = ~n10494 & n10498;
  assign n10500 = ~n10497 & n10499;
  assign n10501 = pi8  & n10500;
  assign n10502 = ~pi8  & ~n10500;
  assign n10503 = ~n10501 & ~n10502;
  assign n10504 = n10493 & ~n10503;
  assign n10505 = ~n2165 & n8939;
  assign n10506 = ~n2265 & n8206;
  assign n10507 = ~n2045 & n9355;
  assign n10508 = n5408 & n8200;
  assign n10509 = ~n10506 & ~n10507;
  assign n10510 = ~n10505 & n10509;
  assign n10511 = ~n10508 & n10510;
  assign n10512 = ~pi8  & ~n10511;
  assign n10513 = pi8  & n10511;
  assign n10514 = ~n10512 & ~n10513;
  assign n10515 = n10258 & ~n10260;
  assign n10516 = ~n10261 & ~n10515;
  assign n10517 = ~n10514 & n10516;
  assign n10518 = ~n2356 & n8206;
  assign n10519 = ~n2265 & n8939;
  assign n10520 = ~n2165 & n9355;
  assign n10521 = n5632 & n8200;
  assign n10522 = ~n10518 & ~n10519;
  assign n10523 = ~n10520 & n10522;
  assign n10524 = ~n10521 & n10523;
  assign n10525 = ~pi8  & ~n10524;
  assign n10526 = pi8  & n10524;
  assign n10527 = ~n10525 & ~n10526;
  assign n10528 = n10254 & ~n10256;
  assign n10529 = ~n10257 & ~n10528;
  assign n10530 = ~n10527 & n10529;
  assign n10531 = ~n2356 & n8939;
  assign n10532 = ~n2442 & n8206;
  assign n10533 = ~n2265 & n9355;
  assign n10534 = n5650 & n8200;
  assign n10535 = ~n10532 & ~n10533;
  assign n10536 = ~n10531 & n10535;
  assign n10537 = ~n10534 & n10536;
  assign n10538 = ~pi8  & ~n10537;
  assign n10539 = pi8  & n10537;
  assign n10540 = ~n10538 & ~n10539;
  assign n10541 = n10250 & ~n10252;
  assign n10542 = ~n10253 & ~n10541;
  assign n10543 = ~n10540 & n10542;
  assign n10544 = n10246 & ~n10248;
  assign n10545 = ~n10249 & ~n10544;
  assign n10546 = ~n2356 & n9355;
  assign n10547 = ~n2538 & n8206;
  assign n10548 = ~n2442 & n8939;
  assign n10549 = n6042 & n8200;
  assign n10550 = ~n10546 & ~n10548;
  assign n10551 = ~n10547 & n10550;
  assign n10552 = ~n10549 & n10551;
  assign n10553 = pi8  & n10552;
  assign n10554 = ~pi8  & ~n10552;
  assign n10555 = ~n10553 & ~n10554;
  assign n10556 = n10545 & ~n10555;
  assign n10557 = n10242 & ~n10244;
  assign n10558 = ~n10245 & ~n10557;
  assign n10559 = ~n2622 & n8206;
  assign n10560 = ~n2538 & n8939;
  assign n10561 = ~n2442 & n9355;
  assign n10562 = n5823 & n8200;
  assign n10563 = ~n10559 & ~n10561;
  assign n10564 = ~n10560 & n10563;
  assign n10565 = ~n10562 & n10564;
  assign n10566 = pi8  & n10565;
  assign n10567 = ~pi8  & ~n10565;
  assign n10568 = ~n10566 & ~n10567;
  assign n10569 = n10558 & ~n10568;
  assign n10570 = n10238 & ~n10240;
  assign n10571 = ~n10241 & ~n10570;
  assign n10572 = ~n2538 & n9355;
  assign n10573 = ~n2622 & n8939;
  assign n10574 = ~n2657 & n8206;
  assign n10575 = n6271 & n8200;
  assign n10576 = ~n10572 & ~n10574;
  assign n10577 = ~n10573 & n10576;
  assign n10578 = ~n10575 & n10577;
  assign n10579 = pi8  & n10578;
  assign n10580 = ~pi8  & ~n10578;
  assign n10581 = ~n10579 & ~n10580;
  assign n10582 = n10571 & ~n10581;
  assign n10583 = ~n2622 & n9355;
  assign n10584 = ~n2726 & n8206;
  assign n10585 = ~n2657 & n8939;
  assign n10586 = n6407 & n8200;
  assign n10587 = ~n10583 & ~n10585;
  assign n10588 = ~n10584 & n10587;
  assign n10589 = ~n10586 & n10588;
  assign n10590 = ~pi8  & ~n10589;
  assign n10591 = pi8  & n10589;
  assign n10592 = ~n10590 & ~n10591;
  assign n10593 = n10234 & ~n10236;
  assign n10594 = ~n10237 & ~n10593;
  assign n10595 = ~n10592 & n10594;
  assign n10596 = ~n2657 & n9355;
  assign n10597 = ~n2726 & n8939;
  assign n10598 = ~n2781 & n8206;
  assign n10599 = n6251 & n8200;
  assign n10600 = ~n10596 & ~n10598;
  assign n10601 = ~n10597 & n10600;
  assign n10602 = ~n10599 & n10601;
  assign n10603 = ~pi8  & ~n10602;
  assign n10604 = pi8  & n10602;
  assign n10605 = ~n10603 & ~n10604;
  assign n10606 = n10230 & ~n10232;
  assign n10607 = ~n10233 & ~n10606;
  assign n10608 = ~n10605 & n10607;
  assign n10609 = ~n2866 & n8206;
  assign n10610 = ~n2726 & n9355;
  assign n10611 = ~n2781 & n8939;
  assign n10612 = n6520 & n8200;
  assign n10613 = ~n10609 & ~n10611;
  assign n10614 = ~n10610 & n10613;
  assign n10615 = ~n10612 & n10614;
  assign n10616 = ~pi8  & ~n10615;
  assign n10617 = pi8  & n10615;
  assign n10618 = ~n10616 & ~n10617;
  assign n10619 = n10226 & ~n10228;
  assign n10620 = ~n10229 & ~n10619;
  assign n10621 = ~n10618 & n10620;
  assign n10622 = n10222 & ~n10224;
  assign n10623 = ~n10225 & ~n10622;
  assign n10624 = ~n2866 & n8939;
  assign n10625 = ~n2781 & n9355;
  assign n10626 = ~n2901 & n8206;
  assign n10627 = n6819 & n8200;
  assign n10628 = ~n10624 & ~n10625;
  assign n10629 = ~n10626 & n10628;
  assign n10630 = ~n10627 & n10629;
  assign n10631 = pi8  & n10630;
  assign n10632 = ~pi8  & ~n10630;
  assign n10633 = ~n10631 & ~n10632;
  assign n10634 = n10623 & ~n10633;
  assign n10635 = n10218 & ~n10220;
  assign n10636 = ~n10221 & ~n10635;
  assign n10637 = ~n2866 & n9355;
  assign n10638 = ~n2978 & n8206;
  assign n10639 = ~n2901 & n8939;
  assign n10640 = n6831 & n8200;
  assign n10641 = ~n10637 & ~n10639;
  assign n10642 = ~n10638 & n10641;
  assign n10643 = ~n10640 & n10642;
  assign n10644 = pi8  & n10643;
  assign n10645 = ~pi8  & ~n10643;
  assign n10646 = ~n10644 & ~n10645;
  assign n10647 = n10636 & ~n10646;
  assign n10648 = n10214 & ~n10216;
  assign n10649 = ~n10217 & ~n10648;
  assign n10650 = ~n2901 & n9355;
  assign n10651 = ~n2978 & n8939;
  assign n10652 = ~n3069 & n8206;
  assign n10653 = n6496 & n8200;
  assign n10654 = ~n10650 & ~n10652;
  assign n10655 = ~n10651 & n10654;
  assign n10656 = ~n10653 & n10655;
  assign n10657 = pi8  & n10656;
  assign n10658 = ~pi8  & ~n10656;
  assign n10659 = ~n10657 & ~n10658;
  assign n10660 = n10649 & ~n10659;
  assign n10661 = ~n2978 & n9355;
  assign n10662 = ~n3137 & n8206;
  assign n10663 = ~n3069 & n8939;
  assign n10664 = n6873 & n8200;
  assign n10665 = ~n10661 & ~n10663;
  assign n10666 = ~n10662 & n10665;
  assign n10667 = ~n10664 & n10666;
  assign n10668 = ~pi8  & ~n10667;
  assign n10669 = pi8  & n10667;
  assign n10670 = ~n10668 & ~n10669;
  assign n10671 = n10210 & ~n10212;
  assign n10672 = ~n10213 & ~n10671;
  assign n10673 = ~n10670 & n10672;
  assign n10674 = ~n3069 & n9355;
  assign n10675 = ~n3137 & n8939;
  assign n10676 = ~n3194 & n8206;
  assign n10677 = n6920 & n8200;
  assign n10678 = ~n10674 & ~n10676;
  assign n10679 = ~n10675 & n10678;
  assign n10680 = ~n10677 & n10679;
  assign n10681 = pi8  & n10680;
  assign n10682 = ~pi8  & ~n10680;
  assign n10683 = ~n10681 & ~n10682;
  assign n10684 = n10206 & ~n10208;
  assign n10685 = ~n10209 & ~n10684;
  assign n10686 = ~n10683 & n10685;
  assign n10687 = ~n3137 & n9355;
  assign n10688 = ~n3194 & n8939;
  assign n10689 = ~n3227 & n8206;
  assign n10690 = n6970 & n8200;
  assign n10691 = ~n10688 & ~n10689;
  assign n10692 = ~n10687 & n10691;
  assign n10693 = ~n10690 & n10692;
  assign n10694 = ~pi8  & ~n10693;
  assign n10695 = pi8  & n10693;
  assign n10696 = ~n10694 & ~n10695;
  assign n10697 = pi11  & ~n10186;
  assign n10698 = n10193 & ~n10697;
  assign n10699 = ~n10193 & n10697;
  assign n10700 = ~n10698 & ~n10699;
  assign n10701 = ~n10696 & n10700;
  assign n10702 = ~n3319 & n8206;
  assign n10703 = ~n3227 & n8939;
  assign n10704 = ~n3194 & n9355;
  assign n10705 = n7013 & n8200;
  assign n10706 = ~n10703 & ~n10704;
  assign n10707 = ~n10702 & n10706;
  assign n10708 = ~n10705 & n10707;
  assign n10709 = pi8  & n10708;
  assign n10710 = ~pi8  & ~n10708;
  assign n10711 = ~n10709 & ~n10710;
  assign n10712 = n10180 & ~n10185;
  assign n10713 = ~n10186 & ~n10712;
  assign n10714 = ~n10711 & n10713;
  assign n10715 = ~n3460 & n8199;
  assign n10716 = pi8  & n10715;
  assign n10717 = ~n3376 & n9355;
  assign n10718 = ~n3460 & n8939;
  assign n10719 = ~n7689 & n8200;
  assign n10720 = ~n10717 & ~n10718;
  assign n10721 = ~n10719 & n10720;
  assign n10722 = ~n10716 & n10721;
  assign n10723 = ~n3460 & n8206;
  assign n10724 = ~n3319 & n9355;
  assign n10725 = ~n3376 & n8939;
  assign n10726 = n7049 & n8200;
  assign n10727 = ~n10723 & ~n10725;
  assign n10728 = ~n10724 & n10727;
  assign n10729 = ~n10726 & n10728;
  assign n10730 = pi8  & n10722;
  assign n10731 = n10729 & n10730;
  assign n10732 = n10179 & n10731;
  assign n10733 = ~n3319 & n8939;
  assign n10734 = ~n3376 & n8206;
  assign n10735 = ~n3227 & n9355;
  assign n10736 = n7105 & n8200;
  assign n10737 = ~n10734 & ~n10735;
  assign n10738 = ~n10733 & n10737;
  assign n10739 = ~n10736 & n10738;
  assign n10740 = pi8  & n10739;
  assign n10741 = ~pi8  & ~n10739;
  assign n10742 = ~n10740 & ~n10741;
  assign n10743 = ~n10179 & ~n10731;
  assign n10744 = ~n10732 & ~n10743;
  assign n10745 = ~n10742 & n10744;
  assign n10746 = ~n10732 & ~n10745;
  assign n10747 = n10711 & ~n10713;
  assign n10748 = ~n10714 & ~n10747;
  assign n10749 = ~n10746 & n10748;
  assign n10750 = ~n10714 & ~n10749;
  assign n10751 = n10696 & ~n10700;
  assign n10752 = ~n10701 & ~n10751;
  assign n10753 = ~n10750 & n10752;
  assign n10754 = ~n10701 & ~n10753;
  assign n10755 = n10683 & ~n10685;
  assign n10756 = ~n10686 & ~n10755;
  assign n10757 = ~n10754 & n10756;
  assign n10758 = ~n10686 & ~n10757;
  assign n10759 = n10670 & ~n10672;
  assign n10760 = ~n10673 & ~n10759;
  assign n10761 = ~n10758 & n10760;
  assign n10762 = ~n10673 & ~n10761;
  assign n10763 = ~n10649 & n10659;
  assign n10764 = ~n10660 & ~n10763;
  assign n10765 = ~n10762 & n10764;
  assign n10766 = ~n10660 & ~n10765;
  assign n10767 = ~n10636 & n10646;
  assign n10768 = ~n10647 & ~n10767;
  assign n10769 = ~n10766 & n10768;
  assign n10770 = ~n10647 & ~n10769;
  assign n10771 = ~n10623 & n10633;
  assign n10772 = ~n10634 & ~n10771;
  assign n10773 = ~n10770 & n10772;
  assign n10774 = ~n10634 & ~n10773;
  assign n10775 = n10618 & ~n10620;
  assign n10776 = ~n10621 & ~n10775;
  assign n10777 = ~n10774 & n10776;
  assign n10778 = ~n10621 & ~n10777;
  assign n10779 = n10605 & ~n10607;
  assign n10780 = ~n10608 & ~n10779;
  assign n10781 = ~n10778 & n10780;
  assign n10782 = ~n10608 & ~n10781;
  assign n10783 = n10592 & ~n10594;
  assign n10784 = ~n10595 & ~n10783;
  assign n10785 = ~n10782 & n10784;
  assign n10786 = ~n10595 & ~n10785;
  assign n10787 = ~n10571 & n10581;
  assign n10788 = ~n10582 & ~n10787;
  assign n10789 = ~n10786 & n10788;
  assign n10790 = ~n10582 & ~n10789;
  assign n10791 = ~n10558 & n10568;
  assign n10792 = ~n10569 & ~n10791;
  assign n10793 = ~n10790 & n10792;
  assign n10794 = ~n10569 & ~n10793;
  assign n10795 = ~n10545 & n10555;
  assign n10796 = ~n10556 & ~n10795;
  assign n10797 = ~n10794 & n10796;
  assign n10798 = ~n10556 & ~n10797;
  assign n10799 = n10540 & ~n10542;
  assign n10800 = ~n10543 & ~n10799;
  assign n10801 = ~n10798 & n10800;
  assign n10802 = ~n10543 & ~n10801;
  assign n10803 = n10527 & ~n10529;
  assign n10804 = ~n10530 & ~n10803;
  assign n10805 = ~n10802 & n10804;
  assign n10806 = ~n10530 & ~n10805;
  assign n10807 = n10514 & ~n10516;
  assign n10808 = ~n10517 & ~n10807;
  assign n10809 = ~n10806 & n10808;
  assign n10810 = ~n10517 & ~n10809;
  assign n10811 = ~n10493 & n10503;
  assign n10812 = ~n10504 & ~n10811;
  assign n10813 = ~n10810 & n10812;
  assign n10814 = ~n10504 & ~n10813;
  assign n10815 = ~n10480 & n10490;
  assign n10816 = ~n10491 & ~n10815;
  assign n10817 = ~n10814 & n10816;
  assign n10818 = ~n10491 & ~n10817;
  assign n10819 = ~n10467 & n10477;
  assign n10820 = ~n10478 & ~n10819;
  assign n10821 = ~n10818 & n10820;
  assign n10822 = ~n10478 & ~n10821;
  assign n10823 = n10462 & ~n10464;
  assign n10824 = ~n10465 & ~n10823;
  assign n10825 = ~n10822 & n10824;
  assign n10826 = ~n10465 & ~n10825;
  assign n10827 = n10449 & ~n10451;
  assign n10828 = ~n10452 & ~n10827;
  assign n10829 = ~n10826 & n10828;
  assign n10830 = ~n10452 & ~n10829;
  assign n10831 = ~n10428 & n10438;
  assign n10832 = ~n10439 & ~n10831;
  assign n10833 = ~n10830 & n10832;
  assign n10834 = ~n10439 & ~n10833;
  assign n10835 = ~n10415 & n10425;
  assign n10836 = ~n10426 & ~n10835;
  assign n10837 = ~n10834 & n10836;
  assign n10838 = ~n10426 & ~n10837;
  assign n10839 = ~n10402 & n10412;
  assign n10840 = ~n10413 & ~n10839;
  assign n10841 = ~n10838 & n10840;
  assign n10842 = ~n10413 & ~n10841;
  assign n10843 = ~n10389 & n10399;
  assign n10844 = ~n10400 & ~n10843;
  assign n10845 = ~n10842 & n10844;
  assign n10846 = ~n10400 & ~n10845;
  assign n10847 = ~n10376 & n10386;
  assign n10848 = ~n10387 & ~n10847;
  assign n10849 = ~n10846 & n10848;
  assign n10850 = ~n10387 & ~n10849;
  assign n10851 = ~n10363 & n10373;
  assign n10852 = ~n10374 & ~n10851;
  assign n10853 = ~n10850 & n10852;
  assign n10854 = ~n10374 & ~n10853;
  assign n10855 = ~n10350 & n10360;
  assign n10856 = ~n10361 & ~n10855;
  assign n10857 = ~n10854 & n10856;
  assign n10858 = ~n10361 & ~n10857;
  assign n10859 = n10323 & ~n10325;
  assign n10860 = ~n10326 & ~n10859;
  assign n10861 = ~n10858 & n10860;
  assign n10862 = ~n729 & n9836;
  assign n10863 = ~n621 & n10329;
  assign n10864 = n71 & ~n563;
  assign n10865 = n3921 & n9830;
  assign n10866 = ~n10863 & ~n10864;
  assign n10867 = ~n10862 & n10866;
  assign n10868 = ~n10865 & n10867;
  assign n10869 = ~pi5  & ~n10868;
  assign n10870 = pi5  & n10868;
  assign n10871 = ~n10869 & ~n10870;
  assign n10872 = n10858 & ~n10860;
  assign n10873 = ~n10861 & ~n10872;
  assign n10874 = ~n10871 & n10873;
  assign n10875 = ~n10861 & ~n10874;
  assign n10876 = ~n10339 & ~n10341;
  assign n10877 = ~n10342 & ~n10876;
  assign n10878 = ~n10875 & n10877;
  assign n10879 = ~pi0  & ~pi1 ;
  assign n10880 = ~pi1  & ~pi2 ;
  assign n10881 = pi1  & pi2 ;
  assign n10882 = ~n10880 & ~n10881;
  assign n10883 = n10879 & n10882;
  assign n10884 = pi0  & n10882;
  assign n10885 = ~n3593 & n10884;
  assign n10886 = ~n10883 & ~n10885;
  assign n10887 = ~n563 & ~n10886;
  assign n10888 = ~pi2  & n10887;
  assign n10889 = pi2  & ~n10887;
  assign n10890 = ~n10888 & ~n10889;
  assign n10891 = n71 & ~n621;
  assign n10892 = ~n729 & n10329;
  assign n10893 = ~n802 & n9836;
  assign n10894 = n3955 & n9830;
  assign n10895 = ~n10891 & ~n10893;
  assign n10896 = ~n10892 & n10895;
  assign n10897 = ~n10894 & n10896;
  assign n10898 = pi5  & n10897;
  assign n10899 = ~pi5  & ~n10897;
  assign n10900 = ~n10898 & ~n10899;
  assign n10901 = ~n10890 & ~n10900;
  assign n10902 = n10890 & n10900;
  assign n10903 = ~n10901 & ~n10902;
  assign n10904 = n10854 & ~n10856;
  assign n10905 = ~n10857 & ~n10904;
  assign n10906 = n10903 & n10905;
  assign n10907 = ~n10901 & ~n10906;
  assign n10908 = n10871 & ~n10873;
  assign n10909 = ~n10874 & ~n10908;
  assign n10910 = ~n10907 & n10909;
  assign n10911 = n71 & ~n729;
  assign n10912 = ~n802 & n10329;
  assign n10913 = ~n898 & n9836;
  assign n10914 = n3901 & n9830;
  assign n10915 = ~n10912 & ~n10913;
  assign n10916 = ~n10911 & n10915;
  assign n10917 = ~n10914 & n10916;
  assign n10918 = ~pi5  & ~n10917;
  assign n10919 = pi5  & n10917;
  assign n10920 = ~n10918 & ~n10919;
  assign n10921 = n10850 & ~n10852;
  assign n10922 = ~n10853 & ~n10921;
  assign n10923 = ~n10920 & n10922;
  assign n10924 = n71 & ~n802;
  assign n10925 = ~n898 & n10329;
  assign n10926 = ~n1006 & n9836;
  assign n10927 = n4057 & n9830;
  assign n10928 = ~n10924 & ~n10925;
  assign n10929 = ~n10926 & n10928;
  assign n10930 = ~n10927 & n10929;
  assign n10931 = ~pi5  & ~n10930;
  assign n10932 = pi5  & n10930;
  assign n10933 = ~n10931 & ~n10932;
  assign n10934 = n10846 & ~n10848;
  assign n10935 = ~n10849 & ~n10934;
  assign n10936 = ~n10933 & n10935;
  assign n10937 = n71 & ~n898;
  assign n10938 = ~n1006 & n10329;
  assign n10939 = ~n1107 & n9836;
  assign n10940 = n4041 & n9830;
  assign n10941 = ~n10937 & ~n10938;
  assign n10942 = ~n10939 & n10941;
  assign n10943 = ~n10940 & n10942;
  assign n10944 = ~pi5  & ~n10943;
  assign n10945 = pi5  & n10943;
  assign n10946 = ~n10944 & ~n10945;
  assign n10947 = n10842 & ~n10844;
  assign n10948 = ~n10845 & ~n10947;
  assign n10949 = ~n10946 & n10948;
  assign n10950 = ~n1107 & n10329;
  assign n10951 = n71 & ~n1006;
  assign n10952 = ~n1230 & n9836;
  assign n10953 = n4233 & n9830;
  assign n10954 = ~n10950 & ~n10951;
  assign n10955 = ~n10952 & n10954;
  assign n10956 = ~n10953 & n10955;
  assign n10957 = ~pi5  & ~n10956;
  assign n10958 = pi5  & n10956;
  assign n10959 = ~n10957 & ~n10958;
  assign n10960 = n10838 & ~n10840;
  assign n10961 = ~n10841 & ~n10960;
  assign n10962 = ~n10959 & n10961;
  assign n10963 = ~n1337 & n9836;
  assign n10964 = ~n1230 & n10329;
  assign n10965 = n71 & ~n1107;
  assign n10966 = n4251 & n9830;
  assign n10967 = ~n10963 & ~n10964;
  assign n10968 = ~n10965 & n10967;
  assign n10969 = ~n10966 & n10968;
  assign n10970 = ~pi5  & ~n10969;
  assign n10971 = pi5  & n10969;
  assign n10972 = ~n10970 & ~n10971;
  assign n10973 = n10834 & ~n10836;
  assign n10974 = ~n10837 & ~n10973;
  assign n10975 = ~n10972 & n10974;
  assign n10976 = ~n1425 & n9836;
  assign n10977 = ~n1337 & n10329;
  assign n10978 = n71 & ~n1230;
  assign n10979 = n4549 & n9830;
  assign n10980 = ~n10976 & ~n10977;
  assign n10981 = ~n10978 & n10980;
  assign n10982 = ~n10979 & n10981;
  assign n10983 = ~pi5  & ~n10982;
  assign n10984 = pi5  & n10982;
  assign n10985 = ~n10983 & ~n10984;
  assign n10986 = n10830 & ~n10832;
  assign n10987 = ~n10833 & ~n10986;
  assign n10988 = ~n10985 & n10987;
  assign n10989 = n10826 & ~n10828;
  assign n10990 = ~n10829 & ~n10989;
  assign n10991 = ~n1532 & n9836;
  assign n10992 = ~n1425 & n10329;
  assign n10993 = n71 & ~n1337;
  assign n10994 = n4452 & n9830;
  assign n10995 = ~n10991 & ~n10992;
  assign n10996 = ~n10993 & n10995;
  assign n10997 = ~n10994 & n10996;
  assign n10998 = pi5  & n10997;
  assign n10999 = ~pi5  & ~n10997;
  assign n11000 = ~n10998 & ~n10999;
  assign n11001 = n10990 & ~n11000;
  assign n11002 = n10822 & ~n10824;
  assign n11003 = ~n10825 & ~n11002;
  assign n11004 = ~n1610 & n9836;
  assign n11005 = ~n1532 & n10329;
  assign n11006 = n71 & ~n1425;
  assign n11007 = n4642 & n9830;
  assign n11008 = ~n11004 & ~n11005;
  assign n11009 = ~n11006 & n11008;
  assign n11010 = ~n11007 & n11009;
  assign n11011 = pi5  & n11010;
  assign n11012 = ~pi5  & ~n11010;
  assign n11013 = ~n11011 & ~n11012;
  assign n11014 = n11003 & ~n11013;
  assign n11015 = ~n1737 & n9836;
  assign n11016 = ~n1610 & n10329;
  assign n11017 = n71 & ~n1532;
  assign n11018 = n4626 & n9830;
  assign n11019 = ~n11015 & ~n11016;
  assign n11020 = ~n11017 & n11019;
  assign n11021 = ~n11018 & n11020;
  assign n11022 = ~pi5  & ~n11021;
  assign n11023 = pi5  & n11021;
  assign n11024 = ~n11022 & ~n11023;
  assign n11025 = n10818 & ~n10820;
  assign n11026 = ~n10821 & ~n11025;
  assign n11027 = ~n11024 & n11026;
  assign n11028 = ~n1805 & n9836;
  assign n11029 = ~n1737 & n10329;
  assign n11030 = n71 & ~n1610;
  assign n11031 = n4844 & n9830;
  assign n11032 = ~n11028 & ~n11029;
  assign n11033 = ~n11030 & n11032;
  assign n11034 = ~n11031 & n11033;
  assign n11035 = ~pi5  & ~n11034;
  assign n11036 = pi5  & n11034;
  assign n11037 = ~n11035 & ~n11036;
  assign n11038 = n10814 & ~n10816;
  assign n11039 = ~n10817 & ~n11038;
  assign n11040 = ~n11037 & n11039;
  assign n11041 = ~n1893 & n9836;
  assign n11042 = ~n1805 & n10329;
  assign n11043 = n71 & ~n1737;
  assign n11044 = n4862 & n9830;
  assign n11045 = ~n11041 & ~n11042;
  assign n11046 = ~n11043 & n11045;
  assign n11047 = ~n11044 & n11046;
  assign n11048 = ~pi5  & ~n11047;
  assign n11049 = pi5  & n11047;
  assign n11050 = ~n11048 & ~n11049;
  assign n11051 = n10810 & ~n10812;
  assign n11052 = ~n10813 & ~n11051;
  assign n11053 = ~n11050 & n11052;
  assign n11054 = n10806 & ~n10808;
  assign n11055 = ~n10809 & ~n11054;
  assign n11056 = ~n1997 & n9836;
  assign n11057 = ~n1893 & n10329;
  assign n11058 = n71 & ~n1805;
  assign n11059 = n5212 & n9830;
  assign n11060 = ~n11056 & ~n11057;
  assign n11061 = ~n11058 & n11060;
  assign n11062 = ~n11059 & n11061;
  assign n11063 = pi5  & n11062;
  assign n11064 = ~pi5  & ~n11062;
  assign n11065 = ~n11063 & ~n11064;
  assign n11066 = n11055 & ~n11065;
  assign n11067 = n10802 & ~n10804;
  assign n11068 = ~n10805 & ~n11067;
  assign n11069 = ~n2045 & n9836;
  assign n11070 = ~n1997 & n10329;
  assign n11071 = n71 & ~n1893;
  assign n11072 = n5061 & n9830;
  assign n11073 = ~n11069 & ~n11070;
  assign n11074 = ~n11071 & n11073;
  assign n11075 = ~n11072 & n11074;
  assign n11076 = pi5  & n11075;
  assign n11077 = ~pi5  & ~n11075;
  assign n11078 = ~n11076 & ~n11077;
  assign n11079 = n11068 & ~n11078;
  assign n11080 = n10798 & ~n10800;
  assign n11081 = ~n10801 & ~n11080;
  assign n11082 = ~n2165 & n9836;
  assign n11083 = ~n2045 & n10329;
  assign n11084 = n71 & ~n1997;
  assign n11085 = n5424 & n9830;
  assign n11086 = ~n11083 & ~n11084;
  assign n11087 = ~n11082 & n11086;
  assign n11088 = ~n11085 & n11087;
  assign n11089 = pi5  & n11088;
  assign n11090 = ~pi5  & ~n11088;
  assign n11091 = ~n11089 & ~n11090;
  assign n11092 = n11081 & ~n11091;
  assign n11093 = ~n2165 & n10329;
  assign n11094 = ~n2265 & n9836;
  assign n11095 = n71 & ~n2045;
  assign n11096 = n5408 & n9830;
  assign n11097 = ~n11094 & ~n11095;
  assign n11098 = ~n11093 & n11097;
  assign n11099 = ~n11096 & n11098;
  assign n11100 = ~pi5  & ~n11099;
  assign n11101 = pi5  & n11099;
  assign n11102 = ~n11100 & ~n11101;
  assign n11103 = n10794 & ~n10796;
  assign n11104 = ~n10797 & ~n11103;
  assign n11105 = ~n11102 & n11104;
  assign n11106 = ~n2356 & n9836;
  assign n11107 = ~n2265 & n10329;
  assign n11108 = n71 & ~n2165;
  assign n11109 = n5632 & n9830;
  assign n11110 = ~n11106 & ~n11107;
  assign n11111 = ~n11108 & n11110;
  assign n11112 = ~n11109 & n11111;
  assign n11113 = ~pi5  & ~n11112;
  assign n11114 = pi5  & n11112;
  assign n11115 = ~n11113 & ~n11114;
  assign n11116 = n10790 & ~n10792;
  assign n11117 = ~n10793 & ~n11116;
  assign n11118 = ~n11115 & n11117;
  assign n11119 = ~n2356 & n10329;
  assign n11120 = ~n2442 & n9836;
  assign n11121 = n71 & ~n2265;
  assign n11122 = n5650 & n9830;
  assign n11123 = ~n11120 & ~n11121;
  assign n11124 = ~n11119 & n11123;
  assign n11125 = ~n11122 & n11124;
  assign n11126 = ~pi5  & ~n11125;
  assign n11127 = pi5  & n11125;
  assign n11128 = ~n11126 & ~n11127;
  assign n11129 = n10786 & ~n10788;
  assign n11130 = ~n10789 & ~n11129;
  assign n11131 = ~n11128 & n11130;
  assign n11132 = n10782 & ~n10784;
  assign n11133 = ~n10785 & ~n11132;
  assign n11134 = n71 & ~n2356;
  assign n11135 = ~n2538 & n9836;
  assign n11136 = ~n2442 & n10329;
  assign n11137 = n6042 & n9830;
  assign n11138 = ~n11134 & ~n11136;
  assign n11139 = ~n11135 & n11138;
  assign n11140 = ~n11137 & n11139;
  assign n11141 = pi5  & n11140;
  assign n11142 = ~pi5  & ~n11140;
  assign n11143 = ~n11141 & ~n11142;
  assign n11144 = n11133 & ~n11143;
  assign n11145 = n10778 & ~n10780;
  assign n11146 = ~n10781 & ~n11145;
  assign n11147 = ~n2622 & n9836;
  assign n11148 = ~n2538 & n10329;
  assign n11149 = n71 & ~n2442;
  assign n11150 = n5823 & n9830;
  assign n11151 = ~n11147 & ~n11149;
  assign n11152 = ~n11148 & n11151;
  assign n11153 = ~n11150 & n11152;
  assign n11154 = pi5  & n11153;
  assign n11155 = ~pi5  & ~n11153;
  assign n11156 = ~n11154 & ~n11155;
  assign n11157 = n11146 & ~n11156;
  assign n11158 = n10774 & ~n10776;
  assign n11159 = ~n10777 & ~n11158;
  assign n11160 = n71 & ~n2538;
  assign n11161 = ~n2622 & n10329;
  assign n11162 = ~n2657 & n9836;
  assign n11163 = n6271 & n9830;
  assign n11164 = ~n11160 & ~n11162;
  assign n11165 = ~n11161 & n11164;
  assign n11166 = ~n11163 & n11165;
  assign n11167 = pi5  & n11166;
  assign n11168 = ~pi5  & ~n11166;
  assign n11169 = ~n11167 & ~n11168;
  assign n11170 = n11159 & ~n11169;
  assign n11171 = n71 & ~n2622;
  assign n11172 = ~n2726 & n9836;
  assign n11173 = ~n2657 & n10329;
  assign n11174 = n6407 & n9830;
  assign n11175 = ~n11171 & ~n11173;
  assign n11176 = ~n11172 & n11175;
  assign n11177 = ~n11174 & n11176;
  assign n11178 = ~pi5  & ~n11177;
  assign n11179 = pi5  & n11177;
  assign n11180 = ~n11178 & ~n11179;
  assign n11181 = n10770 & ~n10772;
  assign n11182 = ~n10773 & ~n11181;
  assign n11183 = ~n11180 & n11182;
  assign n11184 = n71 & ~n2657;
  assign n11185 = ~n2726 & n10329;
  assign n11186 = ~n2781 & n9836;
  assign n11187 = n6251 & n9830;
  assign n11188 = ~n11184 & ~n11186;
  assign n11189 = ~n11185 & n11188;
  assign n11190 = ~n11187 & n11189;
  assign n11191 = ~pi5  & ~n11190;
  assign n11192 = pi5  & n11190;
  assign n11193 = ~n11191 & ~n11192;
  assign n11194 = n10766 & ~n10768;
  assign n11195 = ~n10769 & ~n11194;
  assign n11196 = ~n11193 & n11195;
  assign n11197 = ~n2866 & n9836;
  assign n11198 = n71 & ~n2726;
  assign n11199 = ~n2781 & n10329;
  assign n11200 = n6520 & n9830;
  assign n11201 = ~n11197 & ~n11199;
  assign n11202 = ~n11198 & n11201;
  assign n11203 = ~n11200 & n11202;
  assign n11204 = ~pi5  & ~n11203;
  assign n11205 = pi5  & n11203;
  assign n11206 = ~n11204 & ~n11205;
  assign n11207 = n10762 & ~n10764;
  assign n11208 = ~n10765 & ~n11207;
  assign n11209 = ~n11206 & n11208;
  assign n11210 = n10758 & ~n10760;
  assign n11211 = ~n10761 & ~n11210;
  assign n11212 = ~n2866 & n10329;
  assign n11213 = n71 & ~n2781;
  assign n11214 = ~n2901 & n9836;
  assign n11215 = n6819 & n9830;
  assign n11216 = ~n11212 & ~n11213;
  assign n11217 = ~n11214 & n11216;
  assign n11218 = ~n11215 & n11217;
  assign n11219 = pi5  & n11218;
  assign n11220 = ~pi5  & ~n11218;
  assign n11221 = ~n11219 & ~n11220;
  assign n11222 = n11211 & ~n11221;
  assign n11223 = n10754 & ~n10756;
  assign n11224 = ~n10757 & ~n11223;
  assign n11225 = n71 & ~n2866;
  assign n11226 = ~n2978 & n9836;
  assign n11227 = ~n2901 & n10329;
  assign n11228 = n6831 & n9830;
  assign n11229 = ~n11225 & ~n11227;
  assign n11230 = ~n11226 & n11229;
  assign n11231 = ~n11228 & n11230;
  assign n11232 = pi5  & n11231;
  assign n11233 = ~pi5  & ~n11231;
  assign n11234 = ~n11232 & ~n11233;
  assign n11235 = n11224 & ~n11234;
  assign n11236 = n10750 & ~n10752;
  assign n11237 = ~n10753 & ~n11236;
  assign n11238 = n71 & ~n2901;
  assign n11239 = ~n2978 & n10329;
  assign n11240 = ~n3069 & n9836;
  assign n11241 = n6496 & n9830;
  assign n11242 = ~n11238 & ~n11240;
  assign n11243 = ~n11239 & n11242;
  assign n11244 = ~n11241 & n11243;
  assign n11245 = pi5  & n11244;
  assign n11246 = ~pi5  & ~n11244;
  assign n11247 = ~n11245 & ~n11246;
  assign n11248 = n11237 & ~n11247;
  assign n11249 = n71 & ~n2978;
  assign n11250 = ~n3137 & n9836;
  assign n11251 = ~n3069 & n10329;
  assign n11252 = n6873 & n9830;
  assign n11253 = ~n11249 & ~n11251;
  assign n11254 = ~n11250 & n11253;
  assign n11255 = ~n11252 & n11254;
  assign n11256 = ~pi5  & ~n11255;
  assign n11257 = pi5  & n11255;
  assign n11258 = ~n11256 & ~n11257;
  assign n11259 = n10746 & ~n10748;
  assign n11260 = ~n10749 & ~n11259;
  assign n11261 = ~n11258 & n11260;
  assign n11262 = n71 & ~n3069;
  assign n11263 = ~n3137 & n10329;
  assign n11264 = ~n3194 & n9836;
  assign n11265 = n6920 & n9830;
  assign n11266 = ~n11262 & ~n11264;
  assign n11267 = ~n11263 & n11266;
  assign n11268 = ~n11265 & n11267;
  assign n11269 = pi5  & n11268;
  assign n11270 = ~pi5  & ~n11268;
  assign n11271 = ~n11269 & ~n11270;
  assign n11272 = n10742 & ~n10744;
  assign n11273 = ~n10745 & ~n11272;
  assign n11274 = ~n11271 & n11273;
  assign n11275 = n71 & ~n3137;
  assign n11276 = ~n3194 & n10329;
  assign n11277 = ~n3227 & n9836;
  assign n11278 = n6970 & n9830;
  assign n11279 = ~n11276 & ~n11277;
  assign n11280 = ~n11275 & n11279;
  assign n11281 = ~n11278 & n11280;
  assign n11282 = ~pi5  & ~n11281;
  assign n11283 = pi5  & n11281;
  assign n11284 = ~n11282 & ~n11283;
  assign n11285 = pi8  & ~n10722;
  assign n11286 = n10729 & ~n11285;
  assign n11287 = ~n10729 & n11285;
  assign n11288 = ~n11286 & ~n11287;
  assign n11289 = ~n11284 & n11288;
  assign n11290 = ~n3319 & n9836;
  assign n11291 = ~n3227 & n10329;
  assign n11292 = n71 & ~n3194;
  assign n11293 = n7013 & n9830;
  assign n11294 = ~n11291 & ~n11292;
  assign n11295 = ~n11290 & n11294;
  assign n11296 = ~n11293 & n11295;
  assign n11297 = pi5  & n11296;
  assign n11298 = ~pi5  & ~n11296;
  assign n11299 = ~n11297 & ~n11298;
  assign n11300 = n10716 & ~n10721;
  assign n11301 = ~n10722 & ~n11300;
  assign n11302 = ~n11299 & n11301;
  assign n11303 = n67 & ~n3460;
  assign n11304 = pi5  & n11303;
  assign n11305 = n71 & ~n3376;
  assign n11306 = ~n3460 & n10329;
  assign n11307 = ~n7689 & n9830;
  assign n11308 = ~n11305 & ~n11306;
  assign n11309 = ~n11307 & n11308;
  assign n11310 = ~n11304 & n11309;
  assign n11311 = ~n3460 & n9836;
  assign n11312 = n71 & ~n3319;
  assign n11313 = ~n3376 & n10329;
  assign n11314 = n7049 & n9830;
  assign n11315 = ~n11311 & ~n11313;
  assign n11316 = ~n11312 & n11315;
  assign n11317 = ~n11314 & n11316;
  assign n11318 = pi5  & n11310;
  assign n11319 = n11317 & n11318;
  assign n11320 = n10715 & n11319;
  assign n11321 = ~n3319 & n10329;
  assign n11322 = ~n3376 & n9836;
  assign n11323 = n71 & ~n3227;
  assign n11324 = n7105 & n9830;
  assign n11325 = ~n11322 & ~n11323;
  assign n11326 = ~n11321 & n11325;
  assign n11327 = ~n11324 & n11326;
  assign n11328 = pi5  & n11327;
  assign n11329 = ~pi5  & ~n11327;
  assign n11330 = ~n11328 & ~n11329;
  assign n11331 = ~n10715 & ~n11319;
  assign n11332 = ~n11320 & ~n11331;
  assign n11333 = ~n11330 & n11332;
  assign n11334 = ~n11320 & ~n11333;
  assign n11335 = n11299 & ~n11301;
  assign n11336 = ~n11302 & ~n11335;
  assign n11337 = ~n11334 & n11336;
  assign n11338 = ~n11302 & ~n11337;
  assign n11339 = n11284 & ~n11288;
  assign n11340 = ~n11289 & ~n11339;
  assign n11341 = ~n11338 & n11340;
  assign n11342 = ~n11289 & ~n11341;
  assign n11343 = n11271 & ~n11273;
  assign n11344 = ~n11274 & ~n11343;
  assign n11345 = ~n11342 & n11344;
  assign n11346 = ~n11274 & ~n11345;
  assign n11347 = n11258 & ~n11260;
  assign n11348 = ~n11261 & ~n11347;
  assign n11349 = ~n11346 & n11348;
  assign n11350 = ~n11261 & ~n11349;
  assign n11351 = ~n11237 & n11247;
  assign n11352 = ~n11248 & ~n11351;
  assign n11353 = ~n11350 & n11352;
  assign n11354 = ~n11248 & ~n11353;
  assign n11355 = ~n11224 & n11234;
  assign n11356 = ~n11235 & ~n11355;
  assign n11357 = ~n11354 & n11356;
  assign n11358 = ~n11235 & ~n11357;
  assign n11359 = ~n11211 & n11221;
  assign n11360 = ~n11222 & ~n11359;
  assign n11361 = ~n11358 & n11360;
  assign n11362 = ~n11222 & ~n11361;
  assign n11363 = n11206 & ~n11208;
  assign n11364 = ~n11209 & ~n11363;
  assign n11365 = ~n11362 & n11364;
  assign n11366 = ~n11209 & ~n11365;
  assign n11367 = n11193 & ~n11195;
  assign n11368 = ~n11196 & ~n11367;
  assign n11369 = ~n11366 & n11368;
  assign n11370 = ~n11196 & ~n11369;
  assign n11371 = n11180 & ~n11182;
  assign n11372 = ~n11183 & ~n11371;
  assign n11373 = ~n11370 & n11372;
  assign n11374 = ~n11183 & ~n11373;
  assign n11375 = ~n11159 & n11169;
  assign n11376 = ~n11170 & ~n11375;
  assign n11377 = ~n11374 & n11376;
  assign n11378 = ~n11170 & ~n11377;
  assign n11379 = ~n11146 & n11156;
  assign n11380 = ~n11157 & ~n11379;
  assign n11381 = ~n11378 & n11380;
  assign n11382 = ~n11157 & ~n11381;
  assign n11383 = ~n11133 & n11143;
  assign n11384 = ~n11144 & ~n11383;
  assign n11385 = ~n11382 & n11384;
  assign n11386 = ~n11144 & ~n11385;
  assign n11387 = n11128 & ~n11130;
  assign n11388 = ~n11131 & ~n11387;
  assign n11389 = ~n11386 & n11388;
  assign n11390 = ~n11131 & ~n11389;
  assign n11391 = n11115 & ~n11117;
  assign n11392 = ~n11118 & ~n11391;
  assign n11393 = ~n11390 & n11392;
  assign n11394 = ~n11118 & ~n11393;
  assign n11395 = n11102 & ~n11104;
  assign n11396 = ~n11105 & ~n11395;
  assign n11397 = ~n11394 & n11396;
  assign n11398 = ~n11105 & ~n11397;
  assign n11399 = ~n11081 & n11091;
  assign n11400 = ~n11092 & ~n11399;
  assign n11401 = ~n11398 & n11400;
  assign n11402 = ~n11092 & ~n11401;
  assign n11403 = ~n11068 & n11078;
  assign n11404 = ~n11079 & ~n11403;
  assign n11405 = ~n11402 & n11404;
  assign n11406 = ~n11079 & ~n11405;
  assign n11407 = ~n11055 & n11065;
  assign n11408 = ~n11066 & ~n11407;
  assign n11409 = ~n11406 & n11408;
  assign n11410 = ~n11066 & ~n11409;
  assign n11411 = n11050 & ~n11052;
  assign n11412 = ~n11053 & ~n11411;
  assign n11413 = ~n11410 & n11412;
  assign n11414 = ~n11053 & ~n11413;
  assign n11415 = n11037 & ~n11039;
  assign n11416 = ~n11040 & ~n11415;
  assign n11417 = ~n11414 & n11416;
  assign n11418 = ~n11040 & ~n11417;
  assign n11419 = n11024 & ~n11026;
  assign n11420 = ~n11027 & ~n11419;
  assign n11421 = ~n11418 & n11420;
  assign n11422 = ~n11027 & ~n11421;
  assign n11423 = ~n11003 & n11013;
  assign n11424 = ~n11014 & ~n11423;
  assign n11425 = ~n11422 & n11424;
  assign n11426 = ~n11014 & ~n11425;
  assign n11427 = ~n10990 & n11000;
  assign n11428 = ~n11001 & ~n11427;
  assign n11429 = ~n11426 & n11428;
  assign n11430 = ~n11001 & ~n11429;
  assign n11431 = n10985 & ~n10987;
  assign n11432 = ~n10988 & ~n11431;
  assign n11433 = ~n11430 & n11432;
  assign n11434 = ~n10988 & ~n11433;
  assign n11435 = n10972 & ~n10974;
  assign n11436 = ~n10975 & ~n11435;
  assign n11437 = ~n11434 & n11436;
  assign n11438 = ~n10975 & ~n11437;
  assign n11439 = n10959 & ~n10961;
  assign n11440 = ~n10962 & ~n11439;
  assign n11441 = ~n11438 & n11440;
  assign n11442 = ~n10962 & ~n11441;
  assign n11443 = n10946 & ~n10948;
  assign n11444 = ~n10949 & ~n11443;
  assign n11445 = ~n11442 & n11444;
  assign n11446 = ~n10949 & ~n11445;
  assign n11447 = n10933 & ~n10935;
  assign n11448 = ~n10936 & ~n11447;
  assign n11449 = ~n11446 & n11448;
  assign n11450 = ~n10936 & ~n11449;
  assign n11451 = n10920 & ~n10922;
  assign n11452 = ~n10923 & ~n11451;
  assign n11453 = ~n11450 & n11452;
  assign n11454 = ~n10923 & ~n11453;
  assign n11455 = ~n10903 & ~n10905;
  assign n11456 = ~n10906 & ~n11455;
  assign n11457 = ~n11454 & n11456;
  assign n11458 = n11454 & ~n11456;
  assign n11459 = ~n11457 & ~n11458;
  assign n11460 = n11450 & ~n11452;
  assign n11461 = ~n11453 & ~n11460;
  assign n11462 = ~n621 & n10883;
  assign n11463 = ~pi0  & pi1 ;
  assign n11464 = ~n563 & n11463;
  assign n11465 = n3687 & n10884;
  assign n11466 = ~n11462 & ~n11464;
  assign n11467 = ~n11465 & n11466;
  assign n11468 = pi2  & n11467;
  assign n11469 = ~pi2  & ~n11467;
  assign n11470 = ~n11468 & ~n11469;
  assign n11471 = n11461 & ~n11470;
  assign n11472 = n11446 & ~n11448;
  assign n11473 = ~n11449 & ~n11472;
  assign n11474 = ~n729 & n10883;
  assign n11475 = ~n621 & n11463;
  assign n11476 = pi0  & ~n10882;
  assign n11477 = ~n563 & n11476;
  assign n11478 = n3921 & n10884;
  assign n11479 = ~n11475 & ~n11477;
  assign n11480 = ~n11474 & n11479;
  assign n11481 = ~n11478 & n11480;
  assign n11482 = pi2  & n11481;
  assign n11483 = ~pi2  & ~n11481;
  assign n11484 = ~n11482 & ~n11483;
  assign n11485 = n11473 & ~n11484;
  assign n11486 = n11442 & ~n11444;
  assign n11487 = ~n11445 & ~n11486;
  assign n11488 = ~n621 & n11476;
  assign n11489 = ~n729 & n11463;
  assign n11490 = ~n802 & n10883;
  assign n11491 = n3955 & n10884;
  assign n11492 = ~n11488 & ~n11490;
  assign n11493 = ~n11489 & n11492;
  assign n11494 = ~n11491 & n11493;
  assign n11495 = pi2  & n11494;
  assign n11496 = ~pi2  & ~n11494;
  assign n11497 = ~n11495 & ~n11496;
  assign n11498 = n11487 & ~n11497;
  assign n11499 = n11438 & ~n11440;
  assign n11500 = ~n11441 & ~n11499;
  assign n11501 = ~n729 & n11476;
  assign n11502 = ~n802 & n11463;
  assign n11503 = ~n898 & n10883;
  assign n11504 = n3901 & n10884;
  assign n11505 = ~n11502 & ~n11503;
  assign n11506 = ~n11501 & n11505;
  assign n11507 = ~n11504 & n11506;
  assign n11508 = pi2  & n11507;
  assign n11509 = ~pi2  & ~n11507;
  assign n11510 = ~n11508 & ~n11509;
  assign n11511 = n11500 & ~n11510;
  assign n11512 = n11434 & ~n11436;
  assign n11513 = ~n11437 & ~n11512;
  assign n11514 = ~n802 & n11476;
  assign n11515 = ~n898 & n11463;
  assign n11516 = ~n1006 & n10883;
  assign n11517 = n4057 & n10884;
  assign n11518 = ~n11514 & ~n11515;
  assign n11519 = ~n11516 & n11518;
  assign n11520 = ~n11517 & n11519;
  assign n11521 = pi2  & n11520;
  assign n11522 = ~pi2  & ~n11520;
  assign n11523 = ~n11521 & ~n11522;
  assign n11524 = n11513 & ~n11523;
  assign n11525 = ~n11513 & n11523;
  assign n11526 = ~n11524 & ~n11525;
  assign n11527 = n11426 & ~n11428;
  assign n11528 = ~n11429 & ~n11527;
  assign n11529 = n11422 & ~n11424;
  assign n11530 = ~n11425 & ~n11529;
  assign n11531 = ~n1425 & n10883;
  assign n11532 = ~n1337 & n11463;
  assign n11533 = ~n1230 & n11476;
  assign n11534 = n4549 & n10884;
  assign n11535 = ~n11531 & ~n11532;
  assign n11536 = ~n11533 & n11535;
  assign n11537 = ~n11534 & n11536;
  assign n11538 = pi2  & n11537;
  assign n11539 = ~pi2  & ~n11537;
  assign n11540 = n11418 & ~n11420;
  assign n11541 = ~n11421 & ~n11540;
  assign n11542 = ~n1532 & n10883;
  assign n11543 = ~n1425 & n11463;
  assign n11544 = ~n1337 & n11476;
  assign n11545 = n4452 & n10884;
  assign n11546 = ~n11542 & ~n11543;
  assign n11547 = ~n11544 & n11546;
  assign n11548 = ~n11545 & n11547;
  assign n11549 = pi2  & n11548;
  assign n11550 = ~pi2  & ~n11548;
  assign n11551 = n11414 & ~n11416;
  assign n11552 = ~n11417 & ~n11551;
  assign n11553 = n11406 & ~n11408;
  assign n11554 = ~n11409 & ~n11553;
  assign n11555 = n11402 & ~n11404;
  assign n11556 = ~n11405 & ~n11555;
  assign n11557 = n11398 & ~n11400;
  assign n11558 = ~n11401 & ~n11557;
  assign n11559 = ~n1997 & n10883;
  assign n11560 = ~n1893 & n11463;
  assign n11561 = ~n1805 & n11476;
  assign n11562 = n5212 & n10884;
  assign n11563 = ~n11559 & ~n11560;
  assign n11564 = ~n11561 & n11563;
  assign n11565 = ~n11562 & n11564;
  assign n11566 = pi2  & n11565;
  assign n11567 = ~pi2  & ~n11565;
  assign n11568 = n11394 & ~n11396;
  assign n11569 = ~n11397 & ~n11568;
  assign n11570 = ~n2045 & n10883;
  assign n11571 = ~n1997 & n11463;
  assign n11572 = ~n1893 & n11476;
  assign n11573 = n5061 & n10884;
  assign n11574 = ~n11570 & ~n11571;
  assign n11575 = ~n11572 & n11574;
  assign n11576 = ~n11573 & n11575;
  assign n11577 = pi2  & n11576;
  assign n11578 = ~pi2  & ~n11576;
  assign n11579 = n11390 & ~n11392;
  assign n11580 = ~n11393 & ~n11579;
  assign n11581 = n11382 & ~n11384;
  assign n11582 = ~n11385 & ~n11581;
  assign n11583 = n11378 & ~n11380;
  assign n11584 = ~n11381 & ~n11583;
  assign n11585 = n11374 & ~n11376;
  assign n11586 = ~n11377 & ~n11585;
  assign n11587 = ~n2356 & n11476;
  assign n11588 = ~n2538 & n10883;
  assign n11589 = ~n2442 & n11463;
  assign n11590 = n6042 & n10884;
  assign n11591 = ~n11587 & ~n11589;
  assign n11592 = ~n11588 & n11591;
  assign n11593 = ~n11590 & n11592;
  assign n11594 = pi2  & n11593;
  assign n11595 = ~pi2  & ~n11593;
  assign n11596 = n11370 & ~n11372;
  assign n11597 = ~n11373 & ~n11596;
  assign n11598 = ~n2622 & n10883;
  assign n11599 = ~n2538 & n11463;
  assign n11600 = ~n2442 & n11476;
  assign n11601 = n5823 & n10884;
  assign n11602 = ~n11598 & ~n11600;
  assign n11603 = ~n11599 & n11602;
  assign n11604 = ~n11601 & n11603;
  assign n11605 = pi2  & n11604;
  assign n11606 = ~pi2  & ~n11604;
  assign n11607 = n11366 & ~n11368;
  assign n11608 = ~n11369 & ~n11607;
  assign n11609 = n11358 & ~n11360;
  assign n11610 = ~n11361 & ~n11609;
  assign n11611 = n11354 & ~n11356;
  assign n11612 = ~n11357 & ~n11611;
  assign n11613 = n11350 & ~n11352;
  assign n11614 = ~n11353 & ~n11613;
  assign n11615 = ~n2866 & n11463;
  assign n11616 = ~n2781 & n11476;
  assign n11617 = ~n2901 & n10883;
  assign n11618 = n6819 & n10884;
  assign n11619 = ~n11615 & ~n11616;
  assign n11620 = ~n11617 & n11619;
  assign n11621 = ~n11618 & n11620;
  assign n11622 = pi2  & n11621;
  assign n11623 = ~pi2  & ~n11621;
  assign n11624 = n11346 & ~n11348;
  assign n11625 = ~n11349 & ~n11624;
  assign n11626 = ~n2866 & n11476;
  assign n11627 = ~n2978 & n10883;
  assign n11628 = ~n2901 & n11463;
  assign n11629 = n6831 & n10884;
  assign n11630 = ~n11626 & ~n11628;
  assign n11631 = ~n11627 & n11630;
  assign n11632 = ~n11629 & n11631;
  assign n11633 = pi2  & n11632;
  assign n11634 = ~pi2  & ~n11632;
  assign n11635 = n11342 & ~n11344;
  assign n11636 = ~n11345 & ~n11635;
  assign n11637 = n11334 & ~n11336;
  assign n11638 = ~n11337 & ~n11637;
  assign n11639 = pi5  & ~n11310;
  assign n11640 = n11317 & ~n11639;
  assign n11641 = ~n11317 & n11639;
  assign n11642 = ~n11640 & ~n11641;
  assign n11643 = n7013 & n10884;
  assign n11644 = ~n3194 & n11476;
  assign n11645 = ~n3227 & n11463;
  assign n11646 = ~n3319 & n10883;
  assign n11647 = ~n11644 & ~n11645;
  assign n11648 = ~n11646 & n11647;
  assign n11649 = ~n11643 & n11648;
  assign n11650 = pi2  & n11649;
  assign n11651 = ~pi2  & ~n11649;
  assign n11652 = ~n11650 & ~n11651;
  assign n11653 = n7049 & n10884;
  assign n11654 = pi1  & ~n3376;
  assign n11655 = n3460 & ~n11654;
  assign n11656 = ~n10880 & ~n11655;
  assign n11657 = ~pi0  & ~n11656;
  assign n11658 = ~n3319 & ~n10882;
  assign n11659 = n3376 & n3460;
  assign n11660 = ~n11658 & n11659;
  assign n11661 = ~n11657 & ~n11660;
  assign n11662 = pi2  & ~n11653;
  assign n11663 = ~n11661 & n11662;
  assign n11664 = ~n11303 & ~n11663;
  assign n11665 = ~n3376 & n10883;
  assign n11666 = n7105 & n10884;
  assign n11667 = ~n3227 & n11476;
  assign n11668 = ~n3319 & n11463;
  assign n11669 = ~n11665 & ~n11667;
  assign n11670 = ~n11668 & n11669;
  assign n11671 = ~n11666 & n11670;
  assign n11672 = ~pi2  & ~n11671;
  assign n11673 = pi2  & n11671;
  assign n11674 = ~n11672 & ~n11673;
  assign n11675 = ~n11664 & ~n11674;
  assign n11676 = n11652 & ~n11675;
  assign n11677 = ~n11652 & n11675;
  assign n11678 = n11304 & ~n11309;
  assign n11679 = ~n11310 & ~n11678;
  assign n11680 = ~n11677 & ~n11679;
  assign n11681 = ~n11676 & ~n11680;
  assign n11682 = n11642 & n11681;
  assign n11683 = ~n11642 & ~n11681;
  assign n11684 = ~n3137 & n11476;
  assign n11685 = ~n3194 & n11463;
  assign n11686 = ~n3227 & n10883;
  assign n11687 = n6970 & n10884;
  assign n11688 = ~n11685 & ~n11686;
  assign n11689 = ~n11684 & n11688;
  assign n11690 = ~n11687 & n11689;
  assign n11691 = pi2  & ~n11690;
  assign n11692 = ~pi2  & n11690;
  assign n11693 = ~n11691 & ~n11692;
  assign n11694 = ~n11683 & n11693;
  assign n11695 = ~n3069 & n11476;
  assign n11696 = ~n3137 & n11463;
  assign n11697 = ~n3194 & n10883;
  assign n11698 = n6920 & n10884;
  assign n11699 = ~n11695 & ~n11697;
  assign n11700 = ~n11696 & n11699;
  assign n11701 = ~n11698 & n11700;
  assign n11702 = pi2  & n11701;
  assign n11703 = ~pi2  & ~n11701;
  assign n11704 = ~n11702 & ~n11703;
  assign n11705 = n11330 & ~n11332;
  assign n11706 = ~n11333 & ~n11705;
  assign n11707 = ~n11704 & n11706;
  assign n11708 = ~n11682 & ~n11694;
  assign n11709 = ~n11707 & n11708;
  assign n11710 = n11704 & ~n11706;
  assign n11711 = ~n11709 & ~n11710;
  assign n11712 = n11638 & n11711;
  assign n11713 = ~n11638 & ~n11711;
  assign n11714 = ~n2978 & n11476;
  assign n11715 = ~n3137 & n10883;
  assign n11716 = ~n3069 & n11463;
  assign n11717 = n6873 & n10884;
  assign n11718 = ~n11714 & ~n11716;
  assign n11719 = ~n11715 & n11718;
  assign n11720 = ~n11717 & n11719;
  assign n11721 = pi2  & ~n11720;
  assign n11722 = ~pi2  & n11720;
  assign n11723 = ~n11721 & ~n11722;
  assign n11724 = ~n11713 & n11723;
  assign n11725 = ~n2901 & n11476;
  assign n11726 = ~n2978 & n11463;
  assign n11727 = ~n3069 & n10883;
  assign n11728 = n6496 & n10884;
  assign n11729 = ~n11725 & ~n11727;
  assign n11730 = ~n11726 & n11729;
  assign n11731 = ~n11728 & n11730;
  assign n11732 = pi2  & n11731;
  assign n11733 = ~pi2  & ~n11731;
  assign n11734 = ~n11732 & ~n11733;
  assign n11735 = n11338 & ~n11340;
  assign n11736 = ~n11341 & ~n11735;
  assign n11737 = ~n11734 & n11736;
  assign n11738 = ~n11712 & ~n11737;
  assign n11739 = ~n11724 & n11738;
  assign n11740 = n11734 & ~n11736;
  assign n11741 = ~n11739 & ~n11740;
  assign n11742 = n11636 & n11741;
  assign n11743 = ~n11633 & ~n11634;
  assign n11744 = ~n11742 & n11743;
  assign n11745 = ~n11636 & ~n11741;
  assign n11746 = ~n11744 & ~n11745;
  assign n11747 = n11625 & n11746;
  assign n11748 = ~n11622 & ~n11623;
  assign n11749 = ~n11747 & n11748;
  assign n11750 = ~n11625 & ~n11746;
  assign n11751 = ~n11749 & ~n11750;
  assign n11752 = n11614 & n11751;
  assign n11753 = ~n11614 & ~n11751;
  assign n11754 = ~n2866 & n10883;
  assign n11755 = ~n2726 & n11476;
  assign n11756 = ~n2781 & n11463;
  assign n11757 = n6520 & n10884;
  assign n11758 = ~n11754 & ~n11756;
  assign n11759 = ~n11755 & n11758;
  assign n11760 = ~n11757 & n11759;
  assign n11761 = pi2  & ~n11760;
  assign n11762 = ~pi2  & n11760;
  assign n11763 = ~n11761 & ~n11762;
  assign n11764 = ~n11753 & n11763;
  assign n11765 = ~n11752 & ~n11764;
  assign n11766 = n11612 & ~n11765;
  assign n11767 = ~n11612 & n11765;
  assign n11768 = ~n2657 & n11476;
  assign n11769 = ~n2726 & n11463;
  assign n11770 = ~n2781 & n10883;
  assign n11771 = n6251 & n10884;
  assign n11772 = ~n11768 & ~n11770;
  assign n11773 = ~n11769 & n11772;
  assign n11774 = ~n11771 & n11773;
  assign n11775 = pi2  & ~n11774;
  assign n11776 = ~pi2  & n11774;
  assign n11777 = ~n11775 & ~n11776;
  assign n11778 = ~n11767 & n11777;
  assign n11779 = ~n11766 & ~n11778;
  assign n11780 = n11610 & ~n11779;
  assign n11781 = ~n11610 & n11779;
  assign n11782 = ~n2622 & n11476;
  assign n11783 = ~n2726 & n10883;
  assign n11784 = ~n2657 & n11463;
  assign n11785 = n6407 & n10884;
  assign n11786 = ~n11782 & ~n11784;
  assign n11787 = ~n11783 & n11786;
  assign n11788 = ~n11785 & n11787;
  assign n11789 = pi2  & ~n11788;
  assign n11790 = ~pi2  & n11788;
  assign n11791 = ~n11789 & ~n11790;
  assign n11792 = ~n11781 & n11791;
  assign n11793 = ~n2538 & n11476;
  assign n11794 = ~n2622 & n11463;
  assign n11795 = ~n2657 & n10883;
  assign n11796 = n6271 & n10884;
  assign n11797 = ~n11793 & ~n11795;
  assign n11798 = ~n11794 & n11797;
  assign n11799 = ~n11796 & n11798;
  assign n11800 = pi2  & n11799;
  assign n11801 = ~pi2  & ~n11799;
  assign n11802 = ~n11800 & ~n11801;
  assign n11803 = n11362 & ~n11364;
  assign n11804 = ~n11365 & ~n11803;
  assign n11805 = ~n11802 & n11804;
  assign n11806 = ~n11780 & ~n11805;
  assign n11807 = ~n11792 & n11806;
  assign n11808 = n11802 & ~n11804;
  assign n11809 = ~n11807 & ~n11808;
  assign n11810 = n11608 & n11809;
  assign n11811 = ~n11605 & ~n11606;
  assign n11812 = ~n11810 & n11811;
  assign n11813 = ~n11608 & ~n11809;
  assign n11814 = ~n11812 & ~n11813;
  assign n11815 = n11597 & n11814;
  assign n11816 = ~n11594 & ~n11595;
  assign n11817 = ~n11815 & n11816;
  assign n11818 = ~n11597 & ~n11814;
  assign n11819 = ~n11817 & ~n11818;
  assign n11820 = n11586 & n11819;
  assign n11821 = ~n11586 & ~n11819;
  assign n11822 = ~n2356 & n11463;
  assign n11823 = ~n2442 & n10883;
  assign n11824 = ~n2265 & n11476;
  assign n11825 = n5650 & n10884;
  assign n11826 = ~n11823 & ~n11824;
  assign n11827 = ~n11822 & n11826;
  assign n11828 = ~n11825 & n11827;
  assign n11829 = pi2  & ~n11828;
  assign n11830 = ~pi2  & n11828;
  assign n11831 = ~n11829 & ~n11830;
  assign n11832 = ~n11821 & n11831;
  assign n11833 = ~n11820 & ~n11832;
  assign n11834 = n11584 & ~n11833;
  assign n11835 = ~n11584 & n11833;
  assign n11836 = ~n2356 & n10883;
  assign n11837 = ~n2265 & n11463;
  assign n11838 = ~n2165 & n11476;
  assign n11839 = n5632 & n10884;
  assign n11840 = ~n11836 & ~n11837;
  assign n11841 = ~n11838 & n11840;
  assign n11842 = ~n11839 & n11841;
  assign n11843 = pi2  & ~n11842;
  assign n11844 = ~pi2  & n11842;
  assign n11845 = ~n11843 & ~n11844;
  assign n11846 = ~n11835 & n11845;
  assign n11847 = ~n11834 & ~n11846;
  assign n11848 = n11582 & ~n11847;
  assign n11849 = ~n11582 & n11847;
  assign n11850 = ~n2165 & n11463;
  assign n11851 = ~n2265 & n10883;
  assign n11852 = ~n2045 & n11476;
  assign n11853 = n5408 & n10884;
  assign n11854 = ~n11851 & ~n11852;
  assign n11855 = ~n11850 & n11854;
  assign n11856 = ~n11853 & n11855;
  assign n11857 = pi2  & ~n11856;
  assign n11858 = ~pi2  & n11856;
  assign n11859 = ~n11857 & ~n11858;
  assign n11860 = ~n11849 & n11859;
  assign n11861 = ~n2165 & n10883;
  assign n11862 = ~n2045 & n11463;
  assign n11863 = ~n1997 & n11476;
  assign n11864 = n5424 & n10884;
  assign n11865 = ~n11862 & ~n11863;
  assign n11866 = ~n11861 & n11865;
  assign n11867 = ~n11864 & n11866;
  assign n11868 = pi2  & n11867;
  assign n11869 = ~pi2  & ~n11867;
  assign n11870 = ~n11868 & ~n11869;
  assign n11871 = n11386 & ~n11388;
  assign n11872 = ~n11389 & ~n11871;
  assign n11873 = ~n11870 & n11872;
  assign n11874 = ~n11848 & ~n11873;
  assign n11875 = ~n11860 & n11874;
  assign n11876 = n11870 & ~n11872;
  assign n11877 = ~n11875 & ~n11876;
  assign n11878 = n11580 & n11877;
  assign n11879 = ~n11577 & ~n11578;
  assign n11880 = ~n11878 & n11879;
  assign n11881 = ~n11580 & ~n11877;
  assign n11882 = ~n11880 & ~n11881;
  assign n11883 = n11569 & n11882;
  assign n11884 = ~n11566 & ~n11567;
  assign n11885 = ~n11883 & n11884;
  assign n11886 = ~n11569 & ~n11882;
  assign n11887 = ~n11885 & ~n11886;
  assign n11888 = n11558 & n11887;
  assign n11889 = ~n11558 & ~n11887;
  assign n11890 = ~n1893 & n10883;
  assign n11891 = ~n1805 & n11463;
  assign n11892 = ~n1737 & n11476;
  assign n11893 = n4862 & n10884;
  assign n11894 = ~n11890 & ~n11891;
  assign n11895 = ~n11892 & n11894;
  assign n11896 = ~n11893 & n11895;
  assign n11897 = pi2  & ~n11896;
  assign n11898 = ~pi2  & n11896;
  assign n11899 = ~n11897 & ~n11898;
  assign n11900 = ~n11889 & n11899;
  assign n11901 = ~n11888 & ~n11900;
  assign n11902 = n11556 & ~n11901;
  assign n11903 = ~n11556 & n11901;
  assign n11904 = ~n1805 & n10883;
  assign n11905 = ~n1737 & n11463;
  assign n11906 = ~n1610 & n11476;
  assign n11907 = n4844 & n10884;
  assign n11908 = ~n11904 & ~n11905;
  assign n11909 = ~n11906 & n11908;
  assign n11910 = ~n11907 & n11909;
  assign n11911 = pi2  & ~n11910;
  assign n11912 = ~pi2  & n11910;
  assign n11913 = ~n11911 & ~n11912;
  assign n11914 = ~n11903 & n11913;
  assign n11915 = ~n11902 & ~n11914;
  assign n11916 = n11554 & ~n11915;
  assign n11917 = ~n11554 & n11915;
  assign n11918 = ~n1737 & n10883;
  assign n11919 = ~n1610 & n11463;
  assign n11920 = ~n1532 & n11476;
  assign n11921 = n4626 & n10884;
  assign n11922 = ~n11918 & ~n11919;
  assign n11923 = ~n11920 & n11922;
  assign n11924 = ~n11921 & n11923;
  assign n11925 = pi2  & ~n11924;
  assign n11926 = ~pi2  & n11924;
  assign n11927 = ~n11925 & ~n11926;
  assign n11928 = ~n11917 & n11927;
  assign n11929 = ~n1610 & n10883;
  assign n11930 = ~n1532 & n11463;
  assign n11931 = ~n1425 & n11476;
  assign n11932 = n4642 & n10884;
  assign n11933 = ~n11929 & ~n11930;
  assign n11934 = ~n11931 & n11933;
  assign n11935 = ~n11932 & n11934;
  assign n11936 = pi2  & n11935;
  assign n11937 = ~pi2  & ~n11935;
  assign n11938 = ~n11936 & ~n11937;
  assign n11939 = n11410 & ~n11412;
  assign n11940 = ~n11413 & ~n11939;
  assign n11941 = ~n11938 & n11940;
  assign n11942 = ~n11916 & ~n11941;
  assign n11943 = ~n11928 & n11942;
  assign n11944 = n11938 & ~n11940;
  assign n11945 = ~n11943 & ~n11944;
  assign n11946 = n11552 & n11945;
  assign n11947 = ~n11549 & ~n11550;
  assign n11948 = ~n11946 & n11947;
  assign n11949 = ~n11552 & ~n11945;
  assign n11950 = ~n11948 & ~n11949;
  assign n11951 = n11541 & n11950;
  assign n11952 = ~n11538 & ~n11539;
  assign n11953 = ~n11951 & n11952;
  assign n11954 = ~n11541 & ~n11950;
  assign n11955 = ~n11953 & ~n11954;
  assign n11956 = n11530 & n11955;
  assign n11957 = ~n11530 & ~n11955;
  assign n11958 = ~n1337 & n10883;
  assign n11959 = ~n1230 & n11463;
  assign n11960 = ~n1107 & n11476;
  assign n11961 = n4251 & n10884;
  assign n11962 = ~n11958 & ~n11959;
  assign n11963 = ~n11960 & n11962;
  assign n11964 = ~n11961 & n11963;
  assign n11965 = pi2  & ~n11964;
  assign n11966 = ~pi2  & n11964;
  assign n11967 = ~n11965 & ~n11966;
  assign n11968 = ~n11957 & n11967;
  assign n11969 = ~n11956 & ~n11968;
  assign n11970 = n11528 & ~n11969;
  assign n11971 = ~n11528 & n11969;
  assign n11972 = ~n1107 & n11463;
  assign n11973 = ~n1006 & n11476;
  assign n11974 = ~n1230 & n10883;
  assign n11975 = n4233 & n10884;
  assign n11976 = ~n11972 & ~n11973;
  assign n11977 = ~n11974 & n11976;
  assign n11978 = ~n11975 & n11977;
  assign n11979 = pi2  & ~n11978;
  assign n11980 = ~pi2  & n11978;
  assign n11981 = ~n11979 & ~n11980;
  assign n11982 = ~n11971 & n11981;
  assign n11983 = ~n898 & n11476;
  assign n11984 = ~n1006 & n11463;
  assign n11985 = ~n1107 & n10883;
  assign n11986 = n4041 & n10884;
  assign n11987 = ~n11983 & ~n11984;
  assign n11988 = ~n11985 & n11987;
  assign n11989 = ~n11986 & n11988;
  assign n11990 = pi2  & n11989;
  assign n11991 = ~pi2  & ~n11989;
  assign n11992 = ~n11990 & ~n11991;
  assign n11993 = n11430 & ~n11432;
  assign n11994 = ~n11433 & ~n11993;
  assign n11995 = ~n11992 & n11994;
  assign n11996 = ~n11970 & ~n11995;
  assign n11997 = ~n11982 & n11996;
  assign n11998 = n11992 & ~n11994;
  assign n11999 = ~n11997 & ~n11998;
  assign n12000 = n11526 & n11999;
  assign n12001 = ~n11524 & ~n12000;
  assign n12002 = ~n11500 & n11510;
  assign n12003 = ~n11511 & ~n12002;
  assign n12004 = ~n12001 & n12003;
  assign n12005 = ~n11511 & ~n12004;
  assign n12006 = ~n11487 & n11497;
  assign n12007 = ~n11498 & ~n12006;
  assign n12008 = ~n12005 & n12007;
  assign n12009 = ~n11498 & ~n12008;
  assign n12010 = ~n11473 & n11484;
  assign n12011 = ~n11485 & ~n12010;
  assign n12012 = ~n12009 & n12011;
  assign n12013 = ~n11485 & ~n12012;
  assign n12014 = ~n11461 & n11470;
  assign n12015 = ~n11471 & ~n12014;
  assign n12016 = ~n12013 & n12015;
  assign n12017 = ~n11471 & ~n12016;
  assign n12018 = n11459 & ~n12017;
  assign n12019 = ~n11457 & ~n12018;
  assign n12020 = n10907 & ~n10909;
  assign n12021 = ~n10910 & ~n12020;
  assign n12022 = ~n12019 & n12021;
  assign n12023 = ~n10910 & ~n12022;
  assign n12024 = n10875 & ~n10877;
  assign n12025 = ~n10878 & ~n12024;
  assign n12026 = ~n12023 & n12025;
  assign n12027 = ~n10878 & ~n12026;
  assign n12028 = n10348 & ~n12027;
  assign n12029 = ~n10346 & ~n12028;
  assign n12030 = n9848 & ~n9850;
  assign n12031 = ~n9851 & ~n12030;
  assign n12032 = ~n12029 & n12031;
  assign n12033 = ~n9851 & ~n12032;
  assign n12034 = n9384 & ~n9386;
  assign n12035 = ~n9387 & ~n12034;
  assign n12036 = ~n12033 & n12035;
  assign n12037 = ~n9387 & ~n12036;
  assign n12038 = n8958 & ~n12037;
  assign n12039 = ~n8956 & ~n12038;
  assign n12040 = n8563 & ~n12039;
  assign n12041 = ~n8561 & ~n12040;
  assign n12042 = n8190 & ~n8192;
  assign n12043 = ~n8193 & ~n12042;
  assign n12044 = ~n12041 & n12043;
  assign n12045 = ~n8193 & ~n12044;
  assign n12046 = n7866 & ~n12045;
  assign n12047 = ~n7864 & ~n12046;
  assign n12048 = n7566 & ~n7568;
  assign n12049 = ~n7569 & ~n12048;
  assign n12050 = ~n12047 & n12049;
  assign n12051 = ~n7569 & ~n12050;
  assign n12052 = n7409 & ~n7411;
  assign n12053 = ~n7412 & ~n12052;
  assign n12054 = ~n12051 & n12053;
  assign n12055 = ~n7412 & ~n12054;
  assign n12056 = n7262 & ~n12055;
  assign n12057 = ~n7260 & ~n12056;
  assign n12058 = n6782 & ~n12057;
  assign n12059 = ~n6780 & ~n12058;
  assign n12060 = n6640 & ~n12059;
  assign n12061 = ~n6638 & ~n12060;
  assign n12062 = n6368 & ~n12061;
  assign n12063 = ~n6366 & ~n12062;
  assign n12064 = n6152 & ~n6154;
  assign n12065 = ~n6155 & ~n12064;
  assign n12066 = ~n12063 & n12065;
  assign n12067 = ~n6155 & ~n12066;
  assign n12068 = n6016 & ~n12067;
  assign n12069 = ~n6014 & ~n12068;
  assign n12070 = n5915 & ~n12069;
  assign n12071 = ~n5913 & ~n12070;
  assign n12072 = n5495 & ~n12071;
  assign n12073 = ~n5493 & ~n12072;
  assign n12074 = n5296 & ~n5298;
  assign n12075 = ~n5299 & ~n12074;
  assign n12076 = ~n12073 & n12075;
  assign n12077 = ~n5299 & ~n12076;
  assign n12078 = n5201 & ~n12077;
  assign n12079 = ~n5199 & ~n12078;
  assign n12080 = n5133 & ~n5135;
  assign n12081 = ~n5136 & ~n12080;
  assign n12082 = ~n12079 & n12081;
  assign n12083 = ~n5136 & ~n12082;
  assign n12084 = n4750 & ~n4752;
  assign n12085 = ~n4753 & ~n12084;
  assign n12086 = ~n12083 & n12085;
  assign n12087 = ~n4753 & ~n12086;
  assign n12088 = n4702 & ~n4704;
  assign n12089 = ~n4705 & ~n12088;
  assign n12090 = ~n12087 & n12089;
  assign n12091 = ~n4705 & ~n12090;
  assign n12092 = n4539 & ~n4541;
  assign n12093 = ~n4542 & ~n12092;
  assign n12094 = ~n12091 & n12093;
  assign n12095 = ~n4542 & ~n12094;
  assign n12096 = n4506 & ~n12095;
  assign n12097 = ~n4504 & ~n12096;
  assign n12098 = n3969 & ~n4079;
  assign n12099 = ~n4080 & ~n12098;
  assign n12100 = ~n12097 & n12099;
  assign n12101 = ~n4080 & ~n12100;
  assign n12102 = ~n3934 & ~n3966;
  assign n12103 = ~n3967 & ~n12102;
  assign n12104 = ~n12101 & n12103;
  assign n12105 = ~n3967 & ~n12104;
  assign n12106 = n3932 & ~n12105;
  assign n12107 = ~n3930 & ~n12106;
  assign n12108 = n3697 & ~n12107;
  assign n12109 = ~n3695 & ~n12108;
  assign n12110 = n3598 & n3608;
  assign n12111 = ~n3609 & ~n12110;
  assign n12112 = ~n12109 & n12111;
  assign n12113 = ~n3609 & ~n12112;
  assign n12114 = ~n196 & ~n318;
  assign n12115 = ~n323 & ~n421;
  assign n12116 = ~n462 & n12115;
  assign n12117 = n1149 & n12114;
  assign n12118 = n1283 & n1762;
  assign n12119 = n4383 & n12118;
  assign n12120 = n12116 & n12117;
  assign n12121 = n4815 & n12120;
  assign n12122 = n12119 & n12121;
  assign n12123 = ~n265 & ~n287;
  assign n12124 = ~n483 & n12123;
  assign n12125 = n1391 & n12124;
  assign n12126 = ~n666 & n2267;
  assign n12127 = ~n216 & ~n359;
  assign n12128 = ~n496 & n12127;
  assign n12129 = ~n254 & ~n381;
  assign n12130 = ~n473 & ~n588;
  assign n12131 = ~n646 & ~n681;
  assign n12132 = n12130 & n12131;
  assign n12133 = n298 & n12129;
  assign n12134 = n2493 & n2566;
  assign n12135 = n3170 & n12134;
  assign n12136 = n12132 & n12133;
  assign n12137 = n12126 & n12128;
  assign n12138 = n12136 & n12137;
  assign n12139 = n12125 & n12135;
  assign n12140 = n12138 & n12139;
  assign n12141 = n3423 & n12140;
  assign n12142 = n2334 & n12141;
  assign n12143 = n4022 & n12142;
  assign n12144 = ~n182 & ~n673;
  assign n12145 = n278 & n12144;
  assign n12146 = n940 & n1114;
  assign n12147 = n1380 & n1632;
  assign n12148 = n1965 & n12147;
  assign n12149 = n12145 & n12146;
  assign n12150 = n1207 & n2730;
  assign n12151 = n6978 & n12150;
  assign n12152 = n12148 & n12149;
  assign n12153 = n6935 & n12152;
  assign n12154 = n2343 & n12151;
  assign n12155 = n12153 & n12154;
  assign n12156 = n12122 & n12155;
  assign n12157 = n4010 & n12156;
  assign n12158 = n12143 & n12157;
  assign n12159 = ~n536 & n555;
  assign n12160 = n552 & n12159;
  assign n12161 = n12158 & n12160;
  assign n12162 = ~n3606 & ~n12161;
  assign n12163 = ~n12113 & n12162;
  assign n12164 = n3606 & n12161;
  assign n12165 = n12113 & n12164;
  assign n12166 = ~n12163 & ~n12165;
  assign n12167 = n12109 & ~n12111;
  assign n12168 = ~n12112 & ~n12167;
  assign n12169 = ~n12162 & ~n12164;
  assign n12170 = ~n12113 & ~n12169;
  assign n12171 = n12113 & n12169;
  assign n12172 = ~n12170 & ~n12171;
  assign n12173 = n12168 & n12172;
  assign n12174 = ~n3697 & n12107;
  assign n12175 = ~n12108 & ~n12174;
  assign n12176 = n12168 & n12175;
  assign n12177 = ~n3932 & n12105;
  assign n12178 = ~n12106 & ~n12177;
  assign n12179 = n12175 & n12178;
  assign n12180 = n12101 & ~n12103;
  assign n12181 = ~n12104 & ~n12180;
  assign n12182 = n12178 & n12181;
  assign n12183 = n12097 & ~n12099;
  assign n12184 = ~n12100 & ~n12183;
  assign n12185 = n12181 & n12184;
  assign n12186 = ~n4506 & n12095;
  assign n12187 = ~n12096 & ~n12186;
  assign n12188 = n12184 & n12187;
  assign n12189 = n12091 & ~n12093;
  assign n12190 = ~n12094 & ~n12189;
  assign n12191 = n12187 & n12190;
  assign n12192 = n12087 & ~n12089;
  assign n12193 = ~n12090 & ~n12192;
  assign n12194 = n12190 & n12193;
  assign n12195 = n12083 & ~n12085;
  assign n12196 = ~n12086 & ~n12195;
  assign n12197 = n12193 & n12196;
  assign n12198 = n12079 & ~n12081;
  assign n12199 = ~n12082 & ~n12198;
  assign n12200 = n12196 & n12199;
  assign n12201 = ~n5201 & n12077;
  assign n12202 = ~n12078 & ~n12201;
  assign n12203 = n12199 & n12202;
  assign n12204 = n12073 & ~n12075;
  assign n12205 = ~n12076 & ~n12204;
  assign n12206 = n12202 & n12205;
  assign n12207 = ~n5495 & n12071;
  assign n12208 = ~n12072 & ~n12207;
  assign n12209 = n12205 & n12208;
  assign n12210 = ~n5915 & n12069;
  assign n12211 = ~n12070 & ~n12210;
  assign n12212 = n12208 & n12211;
  assign n12213 = ~n6016 & n12067;
  assign n12214 = ~n12068 & ~n12213;
  assign n12215 = n12211 & n12214;
  assign n12216 = n12063 & ~n12065;
  assign n12217 = ~n12066 & ~n12216;
  assign n12218 = n12214 & n12217;
  assign n12219 = ~n6368 & n12061;
  assign n12220 = ~n12062 & ~n12219;
  assign n12221 = n12217 & n12220;
  assign n12222 = ~n6640 & n12059;
  assign n12223 = ~n12060 & ~n12222;
  assign n12224 = n12220 & n12223;
  assign n12225 = ~n6782 & n12057;
  assign n12226 = ~n12058 & ~n12225;
  assign n12227 = n12223 & n12226;
  assign n12228 = ~n7262 & n12055;
  assign n12229 = ~n12056 & ~n12228;
  assign n12230 = n12226 & n12229;
  assign n12231 = n12051 & ~n12053;
  assign n12232 = ~n12054 & ~n12231;
  assign n12233 = n12229 & n12232;
  assign n12234 = n12047 & ~n12049;
  assign n12235 = ~n12050 & ~n12234;
  assign n12236 = n12232 & n12235;
  assign n12237 = ~n7866 & n12045;
  assign n12238 = ~n12046 & ~n12237;
  assign n12239 = n12235 & n12238;
  assign n12240 = n12041 & ~n12043;
  assign n12241 = ~n12044 & ~n12240;
  assign n12242 = n12238 & n12241;
  assign n12243 = ~n8563 & n12039;
  assign n12244 = ~n12040 & ~n12243;
  assign n12245 = n12241 & n12244;
  assign n12246 = ~n8958 & n12037;
  assign n12247 = ~n12038 & ~n12246;
  assign n12248 = n12244 & n12247;
  assign n12249 = n12033 & ~n12035;
  assign n12250 = ~n12036 & ~n12249;
  assign n12251 = n12247 & n12250;
  assign n12252 = n12029 & ~n12031;
  assign n12253 = ~n12032 & ~n12252;
  assign n12254 = n12250 & n12253;
  assign n12255 = ~n10348 & n12027;
  assign n12256 = ~n12028 & ~n12255;
  assign n12257 = n12253 & n12256;
  assign n12258 = n12023 & ~n12025;
  assign n12259 = ~n12026 & ~n12258;
  assign n12260 = n12256 & n12259;
  assign n12261 = n12019 & ~n12021;
  assign n12262 = ~n12022 & ~n12261;
  assign n12263 = n12259 & n12262;
  assign n12264 = ~n11459 & n12017;
  assign n12265 = ~n12018 & ~n12264;
  assign n12266 = n12262 & n12265;
  assign n12267 = n12013 & ~n12015;
  assign n12268 = ~n12016 & ~n12267;
  assign n12269 = n12265 & n12268;
  assign n12270 = n12009 & ~n12011;
  assign n12271 = ~n12012 & ~n12270;
  assign n12272 = n12268 & n12271;
  assign n12273 = n12005 & ~n12007;
  assign n12274 = ~n12008 & ~n12273;
  assign n12275 = n12271 & n12274;
  assign n12276 = ~n12271 & ~n12274;
  assign n12277 = ~n12275 & ~n12276;
  assign n12278 = n12001 & ~n12003;
  assign n12279 = ~n12004 & ~n12278;
  assign n12280 = ~n11526 & ~n11999;
  assign n12281 = ~n12000 & ~n12280;
  assign n12282 = n12279 & ~n12281;
  assign n12283 = ~n12274 & n12282;
  assign n12284 = n12279 & ~n12283;
  assign n12285 = n12277 & n12284;
  assign n12286 = ~n12275 & ~n12285;
  assign n12287 = ~n12268 & ~n12271;
  assign n12288 = ~n12272 & ~n12287;
  assign n12289 = ~n12286 & n12288;
  assign n12290 = ~n12272 & ~n12289;
  assign n12291 = ~n12265 & ~n12268;
  assign n12292 = ~n12269 & ~n12291;
  assign n12293 = ~n12290 & n12292;
  assign n12294 = ~n12269 & ~n12293;
  assign n12295 = ~n12262 & ~n12265;
  assign n12296 = ~n12266 & ~n12295;
  assign n12297 = ~n12294 & n12296;
  assign n12298 = ~n12266 & ~n12297;
  assign n12299 = ~n12259 & ~n12262;
  assign n12300 = ~n12263 & ~n12299;
  assign n12301 = ~n12298 & n12300;
  assign n12302 = ~n12263 & ~n12301;
  assign n12303 = ~n12256 & ~n12259;
  assign n12304 = ~n12260 & ~n12303;
  assign n12305 = ~n12302 & n12304;
  assign n12306 = ~n12260 & ~n12305;
  assign n12307 = ~n12253 & ~n12256;
  assign n12308 = ~n12257 & ~n12307;
  assign n12309 = ~n12306 & n12308;
  assign n12310 = ~n12257 & ~n12309;
  assign n12311 = ~n12250 & ~n12253;
  assign n12312 = ~n12254 & ~n12311;
  assign n12313 = ~n12310 & n12312;
  assign n12314 = ~n12254 & ~n12313;
  assign n12315 = ~n12247 & ~n12250;
  assign n12316 = ~n12251 & ~n12315;
  assign n12317 = ~n12314 & n12316;
  assign n12318 = ~n12251 & ~n12317;
  assign n12319 = ~n12244 & ~n12247;
  assign n12320 = ~n12248 & ~n12319;
  assign n12321 = ~n12318 & n12320;
  assign n12322 = ~n12248 & ~n12321;
  assign n12323 = ~n12241 & ~n12244;
  assign n12324 = ~n12245 & ~n12323;
  assign n12325 = ~n12322 & n12324;
  assign n12326 = ~n12245 & ~n12325;
  assign n12327 = ~n12238 & ~n12241;
  assign n12328 = ~n12242 & ~n12327;
  assign n12329 = ~n12326 & n12328;
  assign n12330 = ~n12242 & ~n12329;
  assign n12331 = ~n12235 & ~n12238;
  assign n12332 = ~n12239 & ~n12331;
  assign n12333 = ~n12330 & n12332;
  assign n12334 = ~n12239 & ~n12333;
  assign n12335 = ~n12232 & ~n12235;
  assign n12336 = ~n12236 & ~n12335;
  assign n12337 = ~n12334 & n12336;
  assign n12338 = ~n12236 & ~n12337;
  assign n12339 = ~n12229 & ~n12232;
  assign n12340 = ~n12233 & ~n12339;
  assign n12341 = ~n12338 & n12340;
  assign n12342 = ~n12233 & ~n12341;
  assign n12343 = ~n12226 & ~n12229;
  assign n12344 = ~n12230 & ~n12343;
  assign n12345 = ~n12342 & n12344;
  assign n12346 = ~n12230 & ~n12345;
  assign n12347 = ~n12223 & ~n12226;
  assign n12348 = ~n12227 & ~n12347;
  assign n12349 = ~n12346 & n12348;
  assign n12350 = ~n12227 & ~n12349;
  assign n12351 = ~n12220 & ~n12223;
  assign n12352 = ~n12224 & ~n12351;
  assign n12353 = ~n12350 & n12352;
  assign n12354 = ~n12224 & ~n12353;
  assign n12355 = ~n12217 & ~n12220;
  assign n12356 = ~n12221 & ~n12355;
  assign n12357 = ~n12354 & n12356;
  assign n12358 = ~n12221 & ~n12357;
  assign n12359 = ~n12214 & ~n12217;
  assign n12360 = ~n12218 & ~n12359;
  assign n12361 = ~n12358 & n12360;
  assign n12362 = ~n12218 & ~n12361;
  assign n12363 = ~n12211 & ~n12214;
  assign n12364 = ~n12215 & ~n12363;
  assign n12365 = ~n12362 & n12364;
  assign n12366 = ~n12215 & ~n12365;
  assign n12367 = ~n12208 & ~n12211;
  assign n12368 = ~n12212 & ~n12367;
  assign n12369 = ~n12366 & n12368;
  assign n12370 = ~n12212 & ~n12369;
  assign n12371 = ~n12205 & ~n12208;
  assign n12372 = ~n12209 & ~n12371;
  assign n12373 = ~n12370 & n12372;
  assign n12374 = ~n12209 & ~n12373;
  assign n12375 = ~n12202 & ~n12205;
  assign n12376 = ~n12206 & ~n12375;
  assign n12377 = ~n12374 & n12376;
  assign n12378 = ~n12206 & ~n12377;
  assign n12379 = ~n12199 & ~n12202;
  assign n12380 = ~n12203 & ~n12379;
  assign n12381 = ~n12378 & n12380;
  assign n12382 = ~n12203 & ~n12381;
  assign n12383 = ~n12196 & ~n12199;
  assign n12384 = ~n12200 & ~n12383;
  assign n12385 = ~n12382 & n12384;
  assign n12386 = ~n12200 & ~n12385;
  assign n12387 = ~n12193 & ~n12196;
  assign n12388 = ~n12197 & ~n12387;
  assign n12389 = ~n12386 & n12388;
  assign n12390 = ~n12197 & ~n12389;
  assign n12391 = ~n12190 & ~n12193;
  assign n12392 = ~n12194 & ~n12391;
  assign n12393 = ~n12390 & n12392;
  assign n12394 = ~n12194 & ~n12393;
  assign n12395 = ~n12187 & ~n12190;
  assign n12396 = ~n12191 & ~n12395;
  assign n12397 = ~n12394 & n12396;
  assign n12398 = ~n12191 & ~n12397;
  assign n12399 = ~n12184 & ~n12187;
  assign n12400 = ~n12188 & ~n12399;
  assign n12401 = ~n12398 & n12400;
  assign n12402 = ~n12188 & ~n12401;
  assign n12403 = ~n12181 & ~n12184;
  assign n12404 = ~n12185 & ~n12403;
  assign n12405 = ~n12402 & n12404;
  assign n12406 = ~n12185 & ~n12405;
  assign n12407 = ~n12178 & ~n12181;
  assign n12408 = ~n12182 & ~n12407;
  assign n12409 = ~n12406 & n12408;
  assign n12410 = ~n12182 & ~n12409;
  assign n12411 = ~n12175 & ~n12178;
  assign n12412 = ~n12179 & ~n12411;
  assign n12413 = ~n12410 & n12412;
  assign n12414 = ~n12179 & ~n12413;
  assign n12415 = ~n12168 & ~n12175;
  assign n12416 = ~n12176 & ~n12415;
  assign n12417 = ~n12414 & n12416;
  assign n12418 = ~n12176 & ~n12417;
  assign n12419 = ~n12168 & ~n12172;
  assign n12420 = ~n12173 & ~n12419;
  assign n12421 = ~n12418 & n12420;
  assign n12422 = ~n12173 & ~n12421;
  assign n12423 = n12165 & ~n12422;
  assign n12424 = ~n12166 & ~n12423;
  assign n12425 = n78 & ~n12424;
  assign n12426 = ~n5185 & ~n5267;
  assign n12427 = n5121 & ~n12165;
  assign n12428 = n12426 & ~n12427;
  assign n12429 = ~n12163 & ~n12428;
  assign n12430 = ~n12425 & ~n12429;
  assign n12431 = pi23  & n12430;
  assign n12432 = ~pi23  & ~n12430;
  assign n12433 = ~n12431 & ~n12432;
  assign n12434 = ~n236 & ~n324;
  assign n12435 = ~n494 & n12434;
  assign n12436 = n2787 & n3656;
  assign n12437 = n12435 & n12436;
  assign n12438 = ~n253 & ~n405;
  assign n12439 = n2167 & n12438;
  assign n12440 = n2599 & n2754;
  assign n12441 = n4789 & n12440;
  assign n12442 = n6840 & n12439;
  assign n12443 = n12441 & n12442;
  assign n12444 = n468 & ~n645;
  assign n12445 = n863 & n12444;
  assign n12446 = n3074 & n12445;
  assign n12447 = n5549 & n12437;
  assign n12448 = n12446 & n12447;
  assign n12449 = n12443 & n12448;
  assign n12450 = ~n296 & ~n542;
  assign n12451 = ~n133 & ~n270;
  assign n12452 = ~n338 & ~n354;
  assign n12453 = ~n689 & ~n700;
  assign n12454 = n12452 & n12453;
  assign n12455 = n12450 & n12451;
  assign n12456 = n12454 & n12455;
  assign n12457 = n1398 & n4083;
  assign n12458 = ~n98 & ~n460;
  assign n12459 = ~n172 & ~n319;
  assign n12460 = ~n334 & ~n571;
  assign n12461 = n12459 & n12460;
  assign n12462 = n2360 & n12458;
  assign n12463 = n12461 & n12462;
  assign n12464 = n4951 & n12457;
  assign n12465 = n12463 & n12464;
  assign n12466 = ~n92 & ~n595;
  assign n12467 = ~n667 & n12466;
  assign n12468 = ~n168 & n1375;
  assign n12469 = n2150 & n12468;
  assign n12470 = n12467 & n12469;
  assign n12471 = ~n254 & ~n313;
  assign n12472 = ~n388 & ~n671;
  assign n12473 = n12471 & n12472;
  assign n12474 = n1241 & n1537;
  assign n12475 = n1969 & n2093;
  assign n12476 = n3155 & n12475;
  assign n12477 = n12473 & n12474;
  assign n12478 = n4934 & n12477;
  assign n12479 = n12456 & n12476;
  assign n12480 = n12478 & n12479;
  assign n12481 = n12465 & n12470;
  assign n12482 = n12480 & n12481;
  assign n12483 = n12449 & n12482;
  assign n12484 = n3302 & n12483;
  assign n12485 = ~n389 & ~n407;
  assign n12486 = n1392 & n2097;
  assign n12487 = ~n587 & n2768;
  assign n12488 = n1356 & n1384;
  assign n12489 = n2630 & n5550;
  assign n12490 = n12485 & n12489;
  assign n12491 = n12487 & n12488;
  assign n12492 = n12486 & n12491;
  assign n12493 = n989 & n12490;
  assign n12494 = n3270 & n12493;
  assign n12495 = n2149 & n12492;
  assign n12496 = n12494 & n12495;
  assign n12497 = ~n136 & ~n180;
  assign n12498 = ~n445 & ~n460;
  assign n12499 = ~n580 & n12498;
  assign n12500 = n1266 & n12497;
  assign n12501 = n1486 & n1538;
  assign n12502 = n1593 & n1630;
  assign n12503 = n1754 & n12502;
  assign n12504 = n12500 & n12501;
  assign n12505 = n4359 & n12499;
  assign n12506 = n12504 & n12505;
  assign n12507 = n12503 & n12506;
  assign n12508 = n1845 & n3388;
  assign n12509 = n12507 & n12508;
  assign n12510 = n12496 & n12509;
  assign n12511 = n2506 & n12510;
  assign n12512 = ~n12484 & ~n12511;
  assign n12513 = ~n5901 & ~n5982;
  assign n12514 = ~n5302 & n12513;
  assign n12515 = ~n12163 & ~n12514;
  assign n12516 = pi20  & ~n12515;
  assign n12517 = ~pi20  & n12515;
  assign n12518 = ~n12516 & ~n12517;
  assign n12519 = n12484 & n12511;
  assign n12520 = ~n12512 & ~n12519;
  assign n12521 = n12518 & n12520;
  assign n12522 = ~n12512 & ~n12521;
  assign n12523 = n12143 & ~n12522;
  assign n12524 = ~n12143 & n12522;
  assign n12525 = ~n12523 & ~n12524;
  assign n12526 = n3896 & n12190;
  assign n12527 = n564 & n12196;
  assign n12528 = n3683 & n12193;
  assign n12529 = n12390 & ~n12392;
  assign n12530 = ~n12393 & ~n12529;
  assign n12531 = n566 & n12530;
  assign n12532 = ~n12527 & ~n12528;
  assign n12533 = ~n12526 & n12532;
  assign n12534 = ~n12531 & n12533;
  assign n12535 = n12525 & ~n12534;
  assign n12536 = ~n12525 & n12534;
  assign n12537 = ~n12535 & ~n12536;
  assign n12538 = ~n590 & n1456;
  assign n12539 = n2663 & n12538;
  assign n12540 = ~n118 & ~n162;
  assign n12541 = ~n210 & ~n225;
  assign n12542 = ~n267 & ~n334;
  assign n12543 = ~n447 & ~n666;
  assign n12544 = n12542 & n12543;
  assign n12545 = n12540 & n12541;
  assign n12546 = n921 & n1651;
  assign n12547 = n1904 & n2566;
  assign n12548 = n12546 & n12547;
  assign n12549 = n12544 & n12545;
  assign n12550 = n1202 & n3324;
  assign n12551 = n12549 & n12550;
  assign n12552 = n12548 & n12551;
  assign n12553 = n2693 & n12552;
  assign n12554 = ~n122 & ~n168;
  assign n12555 = ~n224 & ~n405;
  assign n12556 = ~n522 & n12555;
  assign n12557 = n344 & n12554;
  assign n12558 = n741 & n1175;
  assign n12559 = n1237 & n2097;
  assign n12560 = n2272 & n3710;
  assign n12561 = n12559 & n12560;
  assign n12562 = n12557 & n12558;
  assign n12563 = n4930 & n12556;
  assign n12564 = n12562 & n12563;
  assign n12565 = n2031 & n12561;
  assign n12566 = n12539 & n12565;
  assign n12567 = n12564 & n12566;
  assign n12568 = n2705 & n12567;
  assign n12569 = n5717 & n12553;
  assign n12570 = n12568 & n12569;
  assign n12571 = n12484 & ~n12570;
  assign n12572 = ~n12484 & n12570;
  assign n12573 = ~n12571 & ~n12572;
  assign n12574 = n3896 & n12196;
  assign n12575 = n3683 & n12199;
  assign n12576 = n564 & n12202;
  assign n12577 = n12382 & ~n12384;
  assign n12578 = ~n12385 & ~n12577;
  assign n12579 = n566 & n12578;
  assign n12580 = ~n12575 & ~n12576;
  assign n12581 = ~n12574 & n12580;
  assign n12582 = ~n12579 & n12581;
  assign n12583 = n12573 & ~n12582;
  assign n12584 = ~n12571 & ~n12583;
  assign n12585 = ~n12518 & ~n12520;
  assign n12586 = ~n12521 & ~n12585;
  assign n12587 = n12584 & ~n12586;
  assign n12588 = ~n12584 & n12586;
  assign n12589 = ~n12587 & ~n12588;
  assign n12590 = n3896 & n12193;
  assign n12591 = n3683 & n12196;
  assign n12592 = n564 & n12199;
  assign n12593 = n12386 & ~n12388;
  assign n12594 = ~n12389 & ~n12593;
  assign n12595 = n566 & n12594;
  assign n12596 = ~n12591 & ~n12592;
  assign n12597 = ~n12590 & n12596;
  assign n12598 = ~n12595 & n12597;
  assign n12599 = n12589 & n12598;
  assign n12600 = ~n12587 & ~n12599;
  assign n12601 = n12537 & n12600;
  assign n12602 = ~n12537 & ~n12600;
  assign n12603 = ~n12601 & ~n12602;
  assign n12604 = n4472 & n12181;
  assign n12605 = n4070 & n12184;
  assign n12606 = n3943 & n12187;
  assign n12607 = n12402 & ~n12404;
  assign n12608 = ~n12405 & ~n12607;
  assign n12609 = n3944 & n12608;
  assign n12610 = ~n12605 & ~n12606;
  assign n12611 = ~n12604 & n12610;
  assign n12612 = ~n12609 & n12611;
  assign n12613 = pi29  & n12612;
  assign n12614 = ~pi29  & ~n12612;
  assign n12615 = ~n12613 & ~n12614;
  assign n12616 = n12603 & ~n12615;
  assign n12617 = ~n12603 & n12615;
  assign n12618 = ~n12616 & ~n12617;
  assign n12619 = ~n12589 & ~n12598;
  assign n12620 = ~n12599 & ~n12619;
  assign n12621 = ~n425 & ~n544;
  assign n12622 = ~n583 & ~n640;
  assign n12623 = n12621 & n12622;
  assign n12624 = n2191 & n3380;
  assign n12625 = n12623 & n12624;
  assign n12626 = ~n192 & ~n682;
  assign n12627 = ~n297 & ~n388;
  assign n12628 = ~n164 & ~n279;
  assign n12629 = ~n446 & ~n514;
  assign n12630 = n12628 & n12629;
  assign n12631 = n178 & n403;
  assign n12632 = n743 & n1174;
  assign n12633 = n1247 & n3763;
  assign n12634 = n12626 & n12627;
  assign n12635 = n12633 & n12634;
  assign n12636 = n12631 & n12632;
  assign n12637 = n2205 & n12630;
  assign n12638 = n3142 & n12637;
  assign n12639 = n12635 & n12636;
  assign n12640 = n12625 & n12639;
  assign n12641 = n5768 & n12638;
  assign n12642 = n12640 & n12641;
  assign n12643 = n3051 & n12642;
  assign n12644 = n4324 & n12643;
  assign n12645 = ~n163 & ~n199;
  assign n12646 = n361 & n12645;
  assign n12647 = ~n279 & ~n286;
  assign n12648 = ~n420 & ~n482;
  assign n12649 = n12647 & n12648;
  assign n12650 = ~n209 & ~n253;
  assign n12651 = ~n577 & ~n645;
  assign n12652 = n12650 & n12651;
  assign n12653 = n194 & n2234;
  assign n12654 = n2390 & n3071;
  assign n12655 = n12653 & n12654;
  assign n12656 = n3400 & n12652;
  assign n12657 = n6991 & n12646;
  assign n12658 = n12649 & n12657;
  assign n12659 = n12655 & n12656;
  assign n12660 = n12658 & n12659;
  assign n12661 = n12465 & n12660;
  assign n12662 = n3280 & n12661;
  assign n12663 = n3623 & n5385;
  assign n12664 = n12662 & n12663;
  assign n12665 = ~n12644 & ~n12664;
  assign n12666 = ~n6356 & ~n6608;
  assign n12667 = ~n6133 & n12666;
  assign n12668 = ~n12163 & ~n12667;
  assign n12669 = pi17  & ~n12668;
  assign n12670 = ~pi17  & n12668;
  assign n12671 = ~n12669 & ~n12670;
  assign n12672 = n12644 & n12664;
  assign n12673 = ~n12665 & ~n12672;
  assign n12674 = n12671 & n12673;
  assign n12675 = ~n12665 & ~n12674;
  assign n12676 = n12484 & ~n12675;
  assign n12677 = ~n12484 & n12675;
  assign n12678 = ~n12676 & ~n12677;
  assign n12679 = n3896 & n12199;
  assign n12680 = n564 & n12205;
  assign n12681 = n3683 & n12202;
  assign n12682 = n12378 & ~n12380;
  assign n12683 = ~n12381 & ~n12682;
  assign n12684 = n566 & n12683;
  assign n12685 = ~n12680 & ~n12681;
  assign n12686 = ~n12679 & n12685;
  assign n12687 = ~n12684 & n12686;
  assign n12688 = n12678 & ~n12687;
  assign n12689 = ~n12676 & ~n12688;
  assign n12690 = ~n12573 & n12582;
  assign n12691 = ~n12583 & ~n12690;
  assign n12692 = ~n12689 & n12691;
  assign n12693 = n12689 & ~n12691;
  assign n12694 = ~n12692 & ~n12693;
  assign n12695 = ~n12671 & ~n12673;
  assign n12696 = ~n12674 & ~n12695;
  assign n12697 = n3896 & n12202;
  assign n12698 = n3683 & n12205;
  assign n12699 = n564 & n12208;
  assign n12700 = n12374 & ~n12376;
  assign n12701 = ~n12377 & ~n12700;
  assign n12702 = n566 & n12701;
  assign n12703 = ~n12698 & ~n12699;
  assign n12704 = ~n12697 & n12703;
  assign n12705 = ~n12702 & n12704;
  assign n12706 = n12696 & ~n12705;
  assign n12707 = ~n324 & ~n446;
  assign n12708 = ~n642 & ~n670;
  assign n12709 = ~n683 & n12708;
  assign n12710 = n281 & n12707;
  assign n12711 = n1267 & n1391;
  assign n12712 = n2096 & n3172;
  assign n12713 = n12711 & n12712;
  assign n12714 = n12709 & n12710;
  assign n12715 = n12713 & n12714;
  assign n12716 = ~n208 & ~n376;
  assign n12717 = ~n271 & ~n539;
  assign n12718 = ~n650 & ~n675;
  assign n12719 = n12717 & n12718;
  assign n12720 = n758 & n12719;
  assign n12721 = ~n145 & ~n288;
  assign n12722 = ~n312 & ~n587;
  assign n12723 = n12721 & n12722;
  assign n12724 = n2220 & n3350;
  assign n12725 = n4384 & n5338;
  assign n12726 = n12716 & n12725;
  assign n12727 = n12723 & n12724;
  assign n12728 = n12726 & n12727;
  assign n12729 = n6416 & n12720;
  assign n12730 = n12728 & n12729;
  assign n12731 = n4968 & n12730;
  assign n12732 = ~n679 & n3323;
  assign n12733 = n12731 & n12732;
  assign n12734 = n2390 & n3171;
  assign n12735 = ~n199 & ~n382;
  assign n12736 = ~n390 & ~n598;
  assign n12737 = ~n602 & n12736;
  assign n12738 = n622 & n12735;
  assign n12739 = n1904 & n12485;
  assign n12740 = n12738 & n12739;
  assign n12741 = n2054 & n12737;
  assign n12742 = n2674 & n12734;
  assign n12743 = n12741 & n12742;
  assign n12744 = n3781 & n12740;
  assign n12745 = n12743 & n12744;
  assign n12746 = n12715 & n12745;
  assign n12747 = n3442 & n12746;
  assign n12748 = n12733 & n12747;
  assign n12749 = n12644 & ~n12748;
  assign n12750 = ~n342 & ~n645;
  assign n12751 = n5599 & n12750;
  assign n12752 = ~n404 & ~n492;
  assign n12753 = ~n479 & ~n675;
  assign n12754 = ~n168 & ~n327;
  assign n12755 = n742 & n12754;
  assign n12756 = n855 & n3870;
  assign n12757 = n12752 & n12753;
  assign n12758 = n12756 & n12757;
  assign n12759 = n12755 & n12758;
  assign n12760 = n5759 & n12759;
  assign n12761 = n1918 & n3362;
  assign n12762 = n12760 & n12761;
  assign n12763 = n1146 & n12762;
  assign n12764 = n12751 & n12763;
  assign n12765 = n925 & n1714;
  assign n12766 = ~n167 & ~n375;
  assign n12767 = ~n224 & ~n702;
  assign n12768 = ~n307 & ~n572;
  assign n12769 = n1469 & n12768;
  assign n12770 = n2220 & n12767;
  assign n12771 = n12769 & n12770;
  assign n12772 = ~n202 & ~n250;
  assign n12773 = ~n267 & ~n480;
  assign n12774 = ~n587 & n12773;
  assign n12775 = n12766 & n12772;
  assign n12776 = n12774 & n12775;
  assign n12777 = n4936 & n5001;
  assign n12778 = n12765 & n12777;
  assign n12779 = n1475 & n12776;
  assign n12780 = n4288 & n12771;
  assign n12781 = n12779 & n12780;
  assign n12782 = n2576 & n12778;
  assign n12783 = n12781 & n12782;
  assign n12784 = n2558 & n12783;
  assign n12785 = n6854 & n12784;
  assign n12786 = ~n12764 & ~n12785;
  assign n12787 = ~n7243 & ~n7380;
  assign n12788 = ~n6646 & n12787;
  assign n12789 = ~n12163 & ~n12788;
  assign n12790 = pi14  & ~n12789;
  assign n12791 = ~pi14  & n12789;
  assign n12792 = ~n12790 & ~n12791;
  assign n12793 = n12764 & n12785;
  assign n12794 = ~n12786 & ~n12793;
  assign n12795 = n12792 & n12794;
  assign n12796 = ~n12786 & ~n12795;
  assign n12797 = n12748 & ~n12796;
  assign n12798 = ~n12748 & n12796;
  assign n12799 = ~n12797 & ~n12798;
  assign n12800 = n3896 & n12208;
  assign n12801 = n564 & n12214;
  assign n12802 = n3683 & n12211;
  assign n12803 = n12366 & ~n12368;
  assign n12804 = ~n12369 & ~n12803;
  assign n12805 = n566 & n12804;
  assign n12806 = ~n12801 & ~n12802;
  assign n12807 = ~n12800 & n12806;
  assign n12808 = ~n12805 & n12807;
  assign n12809 = n12799 & ~n12808;
  assign n12810 = ~n12797 & ~n12809;
  assign n12811 = ~n12644 & n12748;
  assign n12812 = ~n12749 & ~n12811;
  assign n12813 = ~n12810 & n12812;
  assign n12814 = ~n12749 & ~n12813;
  assign n12815 = ~n12696 & n12705;
  assign n12816 = ~n12706 & ~n12815;
  assign n12817 = ~n12814 & n12816;
  assign n12818 = ~n12706 & ~n12817;
  assign n12819 = ~n12678 & n12687;
  assign n12820 = ~n12688 & ~n12819;
  assign n12821 = ~n12818 & n12820;
  assign n12822 = n12818 & ~n12820;
  assign n12823 = ~n12821 & ~n12822;
  assign n12824 = n4472 & n12190;
  assign n12825 = n4070 & n12193;
  assign n12826 = n3943 & n12196;
  assign n12827 = n3944 & n12530;
  assign n12828 = ~n12825 & ~n12826;
  assign n12829 = ~n12824 & n12828;
  assign n12830 = ~n12827 & n12829;
  assign n12831 = pi29  & n12830;
  assign n12832 = ~pi29  & ~n12830;
  assign n12833 = ~n12831 & ~n12832;
  assign n12834 = n12823 & ~n12833;
  assign n12835 = ~n12821 & ~n12834;
  assign n12836 = n12694 & ~n12835;
  assign n12837 = ~n12692 & ~n12836;
  assign n12838 = n12620 & n12837;
  assign n12839 = ~n12620 & ~n12837;
  assign n12840 = ~n12838 & ~n12839;
  assign n12841 = n4472 & n12184;
  assign n12842 = n4070 & n12187;
  assign n12843 = n3943 & n12190;
  assign n12844 = n12398 & ~n12400;
  assign n12845 = ~n12401 & ~n12844;
  assign n12846 = n3944 & n12845;
  assign n12847 = ~n12842 & ~n12843;
  assign n12848 = ~n12841 & n12847;
  assign n12849 = ~n12846 & n12848;
  assign n12850 = pi29  & n12849;
  assign n12851 = ~pi29  & ~n12849;
  assign n12852 = ~n12850 & ~n12851;
  assign n12853 = n12840 & n12852;
  assign n12854 = ~n12838 & ~n12853;
  assign n12855 = ~n12618 & ~n12854;
  assign n12856 = n12618 & n12854;
  assign n12857 = ~n12855 & ~n12856;
  assign n12858 = n4721 & n12168;
  assign n12859 = n4691 & n12175;
  assign n12860 = n4515 & n12178;
  assign n12861 = n12414 & ~n12416;
  assign n12862 = ~n12417 & ~n12861;
  assign n12863 = n4516 & n12862;
  assign n12864 = ~n12859 & ~n12860;
  assign n12865 = ~n12858 & n12864;
  assign n12866 = ~n12863 & n12865;
  assign n12867 = pi26  & n12866;
  assign n12868 = ~pi26  & ~n12866;
  assign n12869 = ~n12867 & ~n12868;
  assign n12870 = n12857 & n12869;
  assign n12871 = ~n12855 & ~n12870;
  assign n12872 = ~n12433 & n12871;
  assign n12873 = n12433 & ~n12871;
  assign n12874 = ~n12872 & ~n12873;
  assign n12875 = ~n12601 & ~n12616;
  assign n12876 = n4472 & n12178;
  assign n12877 = n4070 & n12181;
  assign n12878 = n3943 & n12184;
  assign n12879 = n12406 & ~n12408;
  assign n12880 = ~n12409 & ~n12879;
  assign n12881 = n3944 & n12880;
  assign n12882 = ~n12877 & ~n12878;
  assign n12883 = ~n12876 & n12882;
  assign n12884 = ~n12881 & n12883;
  assign n12885 = pi29  & n12884;
  assign n12886 = ~pi29  & ~n12884;
  assign n12887 = ~n12885 & ~n12886;
  assign n12888 = ~n12523 & ~n12535;
  assign n12889 = ~n118 & ~n649;
  assign n12890 = n1014 & n12889;
  assign n12891 = n1354 & n1837;
  assign n12892 = n3052 & n3995;
  assign n12893 = n4195 & n12892;
  assign n12894 = n12890 & n12891;
  assign n12895 = n884 & n3973;
  assign n12896 = n12894 & n12895;
  assign n12897 = n12893 & n12896;
  assign n12898 = ~n131 & ~n308;
  assign n12899 = ~n539 & n12898;
  assign n12900 = n737 & n1020;
  assign n12901 = n1172 & n1764;
  assign n12902 = n3281 & n12901;
  assign n12903 = n12899 & n12900;
  assign n12904 = n12902 & n12903;
  assign n12905 = n955 & n4149;
  assign n12906 = n6191 & n12905;
  assign n12907 = n12904 & n12906;
  assign n12908 = n12897 & n12907;
  assign n12909 = n12449 & n12908;
  assign n12910 = n4928 & n12909;
  assign n12911 = ~n12143 & n12910;
  assign n12912 = n12143 & ~n12910;
  assign n12913 = ~n12911 & ~n12912;
  assign n12914 = ~n12888 & n12913;
  assign n12915 = n12888 & ~n12913;
  assign n12916 = ~n12914 & ~n12915;
  assign n12917 = n3896 & n12187;
  assign n12918 = n3683 & n12190;
  assign n12919 = n564 & n12193;
  assign n12920 = n12394 & ~n12396;
  assign n12921 = ~n12397 & ~n12920;
  assign n12922 = n566 & n12921;
  assign n12923 = ~n12918 & ~n12919;
  assign n12924 = ~n12917 & n12923;
  assign n12925 = ~n12922 & n12924;
  assign n12926 = n12916 & ~n12925;
  assign n12927 = ~n12916 & n12925;
  assign n12928 = ~n12926 & ~n12927;
  assign n12929 = ~n12887 & n12928;
  assign n12930 = n12887 & ~n12928;
  assign n12931 = ~n12929 & ~n12930;
  assign n12932 = ~n12875 & n12931;
  assign n12933 = n12875 & ~n12931;
  assign n12934 = ~n12932 & ~n12933;
  assign n12935 = n4721 & n12172;
  assign n12936 = n4691 & n12168;
  assign n12937 = n4515 & n12175;
  assign n12938 = n12418 & ~n12420;
  assign n12939 = ~n12421 & ~n12938;
  assign n12940 = n4516 & n12939;
  assign n12941 = ~n12936 & ~n12937;
  assign n12942 = ~n12935 & n12941;
  assign n12943 = ~n12940 & n12942;
  assign n12944 = pi26  & n12943;
  assign n12945 = ~pi26  & ~n12943;
  assign n12946 = ~n12944 & ~n12945;
  assign n12947 = n12934 & ~n12946;
  assign n12948 = ~n12934 & n12946;
  assign n12949 = ~n12947 & ~n12948;
  assign n12950 = n12874 & n12949;
  assign n12951 = ~n12874 & ~n12949;
  assign n12952 = ~n12950 & ~n12951;
  assign n12953 = ~n12857 & ~n12869;
  assign n12954 = ~n12870 & ~n12953;
  assign n12955 = ~n12840 & ~n12852;
  assign n12956 = ~n12853 & ~n12955;
  assign n12957 = n4721 & n12175;
  assign n12958 = n4691 & n12178;
  assign n12959 = n4515 & n12181;
  assign n12960 = n12410 & ~n12412;
  assign n12961 = ~n12413 & ~n12960;
  assign n12962 = n4516 & n12961;
  assign n12963 = ~n12958 & ~n12959;
  assign n12964 = ~n12957 & n12963;
  assign n12965 = ~n12962 & n12964;
  assign n12966 = pi26  & n12965;
  assign n12967 = ~pi26  & ~n12965;
  assign n12968 = ~n12966 & ~n12967;
  assign n12969 = ~n12956 & ~n12968;
  assign n12970 = ~n12694 & n12835;
  assign n12971 = ~n12836 & ~n12970;
  assign n12972 = n4472 & n12187;
  assign n12973 = n4070 & n12190;
  assign n12974 = n3943 & n12193;
  assign n12975 = n3944 & n12921;
  assign n12976 = ~n12973 & ~n12974;
  assign n12977 = ~n12972 & n12976;
  assign n12978 = ~n12975 & n12977;
  assign n12979 = pi29  & n12978;
  assign n12980 = ~pi29  & ~n12978;
  assign n12981 = ~n12979 & ~n12980;
  assign n12982 = n12971 & ~n12981;
  assign n12983 = n4721 & n12178;
  assign n12984 = n4691 & n12181;
  assign n12985 = n4515 & n12184;
  assign n12986 = n4516 & n12880;
  assign n12987 = ~n12984 & ~n12985;
  assign n12988 = ~n12983 & n12987;
  assign n12989 = ~n12986 & n12988;
  assign n12990 = pi26  & n12989;
  assign n12991 = ~pi26  & ~n12989;
  assign n12992 = ~n12990 & ~n12991;
  assign n12993 = ~n12971 & n12981;
  assign n12994 = ~n12982 & ~n12993;
  assign n12995 = ~n12992 & n12994;
  assign n12996 = ~n12982 & ~n12995;
  assign n12997 = n12956 & n12968;
  assign n12998 = ~n12969 & ~n12997;
  assign n12999 = ~n12996 & n12998;
  assign n13000 = ~n12969 & ~n12999;
  assign n13001 = n12954 & n13000;
  assign n13002 = ~n12954 & ~n13000;
  assign n13003 = ~n13001 & ~n13002;
  assign n13004 = ~n12164 & ~n12171;
  assign n13005 = ~n12422 & ~n13004;
  assign n13006 = ~n12172 & ~n13005;
  assign n13007 = ~n12423 & ~n13006;
  assign n13008 = n78 & n13007;
  assign n13009 = n5121 & n12172;
  assign n13010 = ~n5267 & n12165;
  assign n13011 = ~n12163 & ~n12426;
  assign n13012 = ~n13010 & n13011;
  assign n13013 = ~n13009 & ~n13012;
  assign n13014 = ~n13008 & n13013;
  assign n13015 = pi23  & n13014;
  assign n13016 = ~pi23  & ~n13014;
  assign n13017 = ~n13015 & ~n13016;
  assign n13018 = n13003 & n13017;
  assign n13019 = ~n13001 & ~n13018;
  assign n13020 = n12952 & n13019;
  assign n13021 = ~n12952 & ~n13019;
  assign n13022 = ~n13020 & ~n13021;
  assign n13023 = ~n13003 & ~n13017;
  assign n13024 = ~n13018 & ~n13023;
  assign n13025 = n12810 & ~n12812;
  assign n13026 = ~n12813 & ~n13025;
  assign n13027 = n3896 & n12205;
  assign n13028 = n3683 & n12208;
  assign n13029 = n564 & n12211;
  assign n13030 = n12370 & ~n12372;
  assign n13031 = ~n12373 & ~n13030;
  assign n13032 = n566 & n13031;
  assign n13033 = ~n13028 & ~n13029;
  assign n13034 = ~n13027 & n13033;
  assign n13035 = ~n13032 & n13034;
  assign n13036 = n13026 & ~n13035;
  assign n13037 = n4472 & n12196;
  assign n13038 = n4070 & n12199;
  assign n13039 = n3943 & n12202;
  assign n13040 = n3944 & n12578;
  assign n13041 = ~n13038 & ~n13039;
  assign n13042 = ~n13037 & n13041;
  assign n13043 = ~n13040 & n13042;
  assign n13044 = pi29  & n13043;
  assign n13045 = ~pi29  & ~n13043;
  assign n13046 = ~n13044 & ~n13045;
  assign n13047 = ~n13026 & n13035;
  assign n13048 = ~n13036 & ~n13047;
  assign n13049 = ~n13046 & n13048;
  assign n13050 = ~n13036 & ~n13049;
  assign n13051 = n12814 & ~n12816;
  assign n13052 = ~n12817 & ~n13051;
  assign n13053 = ~n13050 & n13052;
  assign n13054 = n4472 & n12193;
  assign n13055 = n4070 & n12196;
  assign n13056 = n3943 & n12199;
  assign n13057 = n3944 & n12594;
  assign n13058 = ~n13055 & ~n13056;
  assign n13059 = ~n13054 & n13058;
  assign n13060 = ~n13057 & n13059;
  assign n13061 = pi29  & n13060;
  assign n13062 = ~pi29  & ~n13060;
  assign n13063 = ~n13061 & ~n13062;
  assign n13064 = n13050 & ~n13052;
  assign n13065 = ~n13053 & ~n13064;
  assign n13066 = ~n13063 & n13065;
  assign n13067 = ~n13053 & ~n13066;
  assign n13068 = ~n12823 & n12833;
  assign n13069 = ~n12834 & ~n13068;
  assign n13070 = ~n13067 & n13069;
  assign n13071 = n13067 & ~n13069;
  assign n13072 = ~n13070 & ~n13071;
  assign n13073 = n4721 & n12181;
  assign n13074 = n4691 & n12184;
  assign n13075 = n4515 & n12187;
  assign n13076 = n4516 & n12608;
  assign n13077 = ~n13074 & ~n13075;
  assign n13078 = ~n13073 & n13077;
  assign n13079 = ~n13076 & n13078;
  assign n13080 = pi26  & n13079;
  assign n13081 = ~pi26  & ~n13079;
  assign n13082 = ~n13080 & ~n13081;
  assign n13083 = n13072 & ~n13082;
  assign n13084 = ~n13070 & ~n13083;
  assign n13085 = n12992 & ~n12994;
  assign n13086 = ~n12995 & ~n13085;
  assign n13087 = ~n13084 & n13086;
  assign n13088 = n13084 & ~n13086;
  assign n13089 = ~n13087 & ~n13088;
  assign n13090 = n5267 & n12172;
  assign n13091 = n5185 & n12168;
  assign n13092 = n5121 & n12175;
  assign n13093 = n78 & n12939;
  assign n13094 = ~n13091 & ~n13092;
  assign n13095 = ~n13090 & n13094;
  assign n13096 = ~n13093 & n13095;
  assign n13097 = pi23  & n13096;
  assign n13098 = ~pi23  & ~n13096;
  assign n13099 = ~n13097 & ~n13098;
  assign n13100 = n13089 & ~n13099;
  assign n13101 = ~n13087 & ~n13100;
  assign n13102 = n5267 & n12166;
  assign n13103 = n5185 & n12172;
  assign n13104 = n5121 & n12168;
  assign n13105 = n12422 & n13004;
  assign n13106 = ~n13005 & ~n13105;
  assign n13107 = n78 & n13106;
  assign n13108 = ~n13102 & ~n13104;
  assign n13109 = ~n13103 & n13108;
  assign n13110 = ~n13107 & n13109;
  assign n13111 = pi23  & n13110;
  assign n13112 = ~pi23  & ~n13110;
  assign n13113 = ~n13111 & ~n13112;
  assign n13114 = ~n13101 & ~n13113;
  assign n13115 = n12996 & ~n12998;
  assign n13116 = ~n12999 & ~n13115;
  assign n13117 = n13101 & n13113;
  assign n13118 = ~n13114 & ~n13117;
  assign n13119 = n13116 & n13118;
  assign n13120 = ~n13114 & ~n13119;
  assign n13121 = ~n13024 & ~n13120;
  assign n13122 = n4721 & n12184;
  assign n13123 = n4691 & n12187;
  assign n13124 = n4515 & n12190;
  assign n13125 = n4516 & n12845;
  assign n13126 = ~n13123 & ~n13124;
  assign n13127 = ~n13122 & n13126;
  assign n13128 = ~n13125 & n13127;
  assign n13129 = pi26  & n13128;
  assign n13130 = ~pi26  & ~n13128;
  assign n13131 = ~n13129 & ~n13130;
  assign n13132 = n13063 & ~n13065;
  assign n13133 = ~n13066 & ~n13132;
  assign n13134 = ~n13131 & n13133;
  assign n13135 = ~n12799 & n12808;
  assign n13136 = ~n12809 & ~n13135;
  assign n13137 = n596 & n1535;
  assign n13138 = ~n162 & ~n299;
  assign n13139 = ~n376 & ~n546;
  assign n13140 = n13138 & n13139;
  assign n13141 = n4162 & n13140;
  assign n13142 = ~n195 & ~n235;
  assign n13143 = ~n340 & ~n650;
  assign n13144 = n13142 & n13143;
  assign n13145 = n1156 & n1710;
  assign n13146 = n1783 & n13145;
  assign n13147 = n826 & n13144;
  assign n13148 = n1151 & n1943;
  assign n13149 = n3785 & n13137;
  assign n13150 = n13148 & n13149;
  assign n13151 = n13146 & n13147;
  assign n13152 = n13141 & n13151;
  assign n13153 = n13150 & n13152;
  assign n13154 = ~n92 & ~n133;
  assign n13155 = ~n213 & ~n666;
  assign n13156 = n13154 & n13155;
  assign n13157 = n740 & n812;
  assign n13158 = n1837 & n2599;
  assign n13159 = n13157 & n13158;
  assign n13160 = n4386 & n13156;
  assign n13161 = n13159 & n13160;
  assign n13162 = ~n179 & ~n192;
  assign n13163 = ~n202 & ~n282;
  assign n13164 = ~n448 & ~n513;
  assign n13165 = ~n554 & ~n645;
  assign n13166 = n13164 & n13165;
  assign n13167 = n13162 & n13163;
  assign n13168 = n523 & n882;
  assign n13169 = n1486 & n2271;
  assign n13170 = n4767 & n13169;
  assign n13171 = n13167 & n13168;
  assign n13172 = n1437 & n13166;
  assign n13173 = n13171 & n13172;
  assign n13174 = n3008 & n13170;
  assign n13175 = n4091 & n13174;
  assign n13176 = n13161 & n13173;
  assign n13177 = n13175 & n13176;
  assign n13178 = n2851 & n13177;
  assign n13179 = n13153 & n13178;
  assign n13180 = n12764 & ~n13179;
  assign n13181 = ~n12764 & n13179;
  assign n13182 = ~n13180 & ~n13181;
  assign n13183 = n3896 & n12214;
  assign n13184 = n3683 & n12217;
  assign n13185 = n564 & n12220;
  assign n13186 = n12358 & ~n12360;
  assign n13187 = ~n12361 & ~n13186;
  assign n13188 = n566 & n13187;
  assign n13189 = ~n13184 & ~n13185;
  assign n13190 = ~n13183 & n13189;
  assign n13191 = ~n13188 & n13190;
  assign n13192 = n13182 & ~n13191;
  assign n13193 = ~n13180 & ~n13192;
  assign n13194 = ~n12792 & ~n12794;
  assign n13195 = ~n12795 & ~n13194;
  assign n13196 = n13193 & ~n13195;
  assign n13197 = ~n13193 & n13195;
  assign n13198 = ~n13196 & ~n13197;
  assign n13199 = n3896 & n12211;
  assign n13200 = n3683 & n12214;
  assign n13201 = n564 & n12217;
  assign n13202 = n12362 & ~n12364;
  assign n13203 = ~n12365 & ~n13202;
  assign n13204 = n566 & n13203;
  assign n13205 = ~n13200 & ~n13201;
  assign n13206 = ~n13199 & n13205;
  assign n13207 = ~n13204 & n13206;
  assign n13208 = n13198 & n13207;
  assign n13209 = ~n13196 & ~n13208;
  assign n13210 = n13136 & n13209;
  assign n13211 = ~n13136 & ~n13209;
  assign n13212 = ~n13210 & ~n13211;
  assign n13213 = n4472 & n12199;
  assign n13214 = n4070 & n12202;
  assign n13215 = n3943 & n12205;
  assign n13216 = n3944 & n12683;
  assign n13217 = ~n13214 & ~n13215;
  assign n13218 = ~n13213 & n13217;
  assign n13219 = ~n13216 & n13218;
  assign n13220 = pi29  & n13219;
  assign n13221 = ~pi29  & ~n13219;
  assign n13222 = ~n13220 & ~n13221;
  assign n13223 = n13212 & ~n13222;
  assign n13224 = ~n13210 & ~n13223;
  assign n13225 = n13046 & ~n13048;
  assign n13226 = ~n13049 & ~n13225;
  assign n13227 = ~n13224 & n13226;
  assign n13228 = n13224 & ~n13226;
  assign n13229 = ~n13227 & ~n13228;
  assign n13230 = n4721 & n12187;
  assign n13231 = n4691 & n12190;
  assign n13232 = n4515 & n12193;
  assign n13233 = n4516 & n12921;
  assign n13234 = ~n13231 & ~n13232;
  assign n13235 = ~n13230 & n13234;
  assign n13236 = ~n13233 & n13235;
  assign n13237 = pi26  & n13236;
  assign n13238 = ~pi26  & ~n13236;
  assign n13239 = ~n13237 & ~n13238;
  assign n13240 = n13229 & ~n13239;
  assign n13241 = ~n13227 & ~n13240;
  assign n13242 = n13131 & ~n13133;
  assign n13243 = ~n13134 & ~n13242;
  assign n13244 = ~n13241 & n13243;
  assign n13245 = ~n13134 & ~n13244;
  assign n13246 = ~n13072 & n13082;
  assign n13247 = ~n13083 & ~n13246;
  assign n13248 = ~n13245 & n13247;
  assign n13249 = n13245 & ~n13247;
  assign n13250 = ~n13248 & ~n13249;
  assign n13251 = n5267 & n12168;
  assign n13252 = n5185 & n12175;
  assign n13253 = n5121 & n12178;
  assign n13254 = n78 & n12862;
  assign n13255 = ~n13252 & ~n13253;
  assign n13256 = ~n13251 & n13255;
  assign n13257 = ~n13254 & n13256;
  assign n13258 = pi23  & n13257;
  assign n13259 = ~pi23  & ~n13257;
  assign n13260 = ~n13258 & ~n13259;
  assign n13261 = n13250 & ~n13260;
  assign n13262 = ~n13248 & ~n13261;
  assign n13263 = n5306 & ~n12424;
  assign n13264 = n5311 & ~n12165;
  assign n13265 = n12513 & ~n13264;
  assign n13266 = ~n12163 & ~n13265;
  assign n13267 = ~n13263 & ~n13266;
  assign n13268 = pi20  & n13267;
  assign n13269 = ~pi20  & ~n13267;
  assign n13270 = ~n13268 & ~n13269;
  assign n13271 = ~n13262 & ~n13270;
  assign n13272 = n13262 & n13270;
  assign n13273 = ~n13271 & ~n13272;
  assign n13274 = ~n13089 & n13099;
  assign n13275 = ~n13100 & ~n13274;
  assign n13276 = n13273 & n13275;
  assign n13277 = ~n13271 & ~n13276;
  assign n13278 = ~n13116 & ~n13118;
  assign n13279 = ~n13119 & ~n13278;
  assign n13280 = ~n13277 & n13279;
  assign n13281 = n13241 & ~n13243;
  assign n13282 = ~n13244 & ~n13281;
  assign n13283 = n5267 & n12175;
  assign n13284 = n5185 & n12178;
  assign n13285 = n5121 & n12181;
  assign n13286 = n78 & n12961;
  assign n13287 = ~n13284 & ~n13285;
  assign n13288 = ~n13283 & n13287;
  assign n13289 = ~n13286 & n13288;
  assign n13290 = pi23  & n13289;
  assign n13291 = ~pi23  & ~n13289;
  assign n13292 = ~n13290 & ~n13291;
  assign n13293 = n13282 & ~n13292;
  assign n13294 = ~n13198 & ~n13207;
  assign n13295 = ~n13208 & ~n13294;
  assign n13296 = n4472 & n12202;
  assign n13297 = n4070 & n12205;
  assign n13298 = n3943 & n12208;
  assign n13299 = n3944 & n12701;
  assign n13300 = ~n13297 & ~n13298;
  assign n13301 = ~n13296 & n13300;
  assign n13302 = ~n13299 & n13301;
  assign n13303 = pi29  & n13302;
  assign n13304 = ~pi29  & ~n13302;
  assign n13305 = ~n13303 & ~n13304;
  assign n13306 = ~n13295 & ~n13305;
  assign n13307 = ~n165 & ~n340;
  assign n13308 = ~n588 & n13307;
  assign n13309 = n1542 & n3658;
  assign n13310 = n13308 & n13309;
  assign n13311 = n278 & n1156;
  assign n13312 = ~n126 & ~n202;
  assign n13313 = ~n283 & ~n311;
  assign n13314 = ~n553 & ~n659;
  assign n13315 = n13313 & n13314;
  assign n13316 = n781 & n13312;
  assign n13317 = n2358 & n2957;
  assign n13318 = n13316 & n13317;
  assign n13319 = n2108 & n13315;
  assign n13320 = n13318 & n13319;
  assign n13321 = ~n145 & ~n148;
  assign n13322 = ~n196 & ~n209;
  assign n13323 = ~n360 & ~n590;
  assign n13324 = n13322 & n13323;
  assign n13325 = n386 & n13321;
  assign n13326 = n403 & n4933;
  assign n13327 = n13325 & n13326;
  assign n13328 = n2757 & n13324;
  assign n13329 = n3626 & n13311;
  assign n13330 = n13328 & n13329;
  assign n13331 = n4798 & n13327;
  assign n13332 = n13310 & n13331;
  assign n13333 = n13320 & n13330;
  assign n13334 = n13332 & n13333;
  assign n13335 = n3418 & n13334;
  assign n13336 = n6470 & n13335;
  assign n13337 = ~n203 & ~n336;
  assign n13338 = ~n118 & ~n219;
  assign n13339 = ~n479 & n2958;
  assign n13340 = n13338 & n13339;
  assign n13341 = n1966 & n13340;
  assign n13342 = ~n420 & ~n679;
  assign n13343 = n380 & n13342;
  assign n13344 = n1756 & n3204;
  assign n13345 = n13337 & n13344;
  assign n13346 = n856 & n13343;
  assign n13347 = n1111 & n2994;
  assign n13348 = n4934 & n13347;
  assign n13349 = n13345 & n13346;
  assign n13350 = n13348 & n13349;
  assign n13351 = n13341 & n13350;
  assign n13352 = n1411 & n1955;
  assign n13353 = n6202 & n13352;
  assign n13354 = n966 & n13351;
  assign n13355 = n13353 & n13354;
  assign n13356 = ~n13336 & ~n13355;
  assign n13357 = ~n7847 & ~n8161;
  assign n13358 = ~n7544 & n13357;
  assign n13359 = ~n12163 & ~n13358;
  assign n13360 = pi11  & ~n13359;
  assign n13361 = ~pi11  & n13359;
  assign n13362 = ~n13360 & ~n13361;
  assign n13363 = n13336 & n13355;
  assign n13364 = ~n13356 & ~n13363;
  assign n13365 = n13362 & n13364;
  assign n13366 = ~n13356 & ~n13365;
  assign n13367 = n12764 & ~n13366;
  assign n13368 = ~n12764 & n13366;
  assign n13369 = ~n13367 & ~n13368;
  assign n13370 = n3896 & n12217;
  assign n13371 = n564 & n12223;
  assign n13372 = n3683 & n12220;
  assign n13373 = n12354 & ~n12356;
  assign n13374 = ~n12357 & ~n13373;
  assign n13375 = n566 & n13374;
  assign n13376 = ~n13371 & ~n13372;
  assign n13377 = ~n13370 & n13376;
  assign n13378 = ~n13375 & n13377;
  assign n13379 = n13369 & ~n13378;
  assign n13380 = ~n13367 & ~n13379;
  assign n13381 = ~n13182 & n13191;
  assign n13382 = ~n13192 & ~n13381;
  assign n13383 = ~n13380 & n13382;
  assign n13384 = n13380 & ~n13382;
  assign n13385 = ~n13383 & ~n13384;
  assign n13386 = ~n13362 & ~n13364;
  assign n13387 = ~n13365 & ~n13386;
  assign n13388 = n3896 & n12220;
  assign n13389 = n3683 & n12223;
  assign n13390 = n564 & n12226;
  assign n13391 = n12350 & ~n12352;
  assign n13392 = ~n12353 & ~n13391;
  assign n13393 = n566 & n13392;
  assign n13394 = ~n13389 & ~n13390;
  assign n13395 = ~n13388 & n13394;
  assign n13396 = ~n13393 & n13395;
  assign n13397 = n13387 & ~n13396;
  assign n13398 = ~n126 & ~n133;
  assign n13399 = ~n265 & ~n270;
  assign n13400 = ~n665 & n13399;
  assign n13401 = n493 & n13398;
  assign n13402 = n623 & n2868;
  assign n13403 = n5526 & n13402;
  assign n13404 = n13400 & n13401;
  assign n13405 = n13403 & n13404;
  assign n13406 = ~n288 & ~n407;
  assign n13407 = ~n286 & ~n495;
  assign n13408 = ~n544 & n13407;
  assign n13409 = n1432 & n13408;
  assign n13410 = ~n296 & ~n470;
  assign n13411 = ~n494 & ~n577;
  assign n13412 = n13410 & n13411;
  assign n13413 = ~n406 & ~n479;
  assign n13414 = ~n588 & ~n644;
  assign n13415 = n13413 & n13414;
  assign n13416 = n688 & n1020;
  assign n13417 = n1157 & n2063;
  assign n13418 = n2192 & n2234;
  assign n13419 = n13417 & n13418;
  assign n13420 = n13415 & n13416;
  assign n13421 = n2189 & n13412;
  assign n13422 = n13420 & n13421;
  assign n13423 = n1040 & n13419;
  assign n13424 = n3263 & n13409;
  assign n13425 = n13423 & n13424;
  assign n13426 = n13422 & n13425;
  assign n13427 = n2672 & n13426;
  assign n13428 = ~n147 & ~n246;
  assign n13429 = ~n483 & ~n599;
  assign n13430 = n13428 & n13429;
  assign n13431 = n281 & n344;
  assign n13432 = n913 & n13406;
  assign n13433 = n13431 & n13432;
  assign n13434 = n1055 & n13430;
  assign n13435 = n2396 & n13137;
  assign n13436 = n13434 & n13435;
  assign n13437 = n13433 & n13436;
  assign n13438 = n13405 & n13437;
  assign n13439 = n4887 & n13438;
  assign n13440 = n13427 & n13439;
  assign n13441 = n13336 & ~n13440;
  assign n13442 = ~n149 & ~n213;
  assign n13443 = ~n282 & ~n286;
  assign n13444 = ~n492 & ~n496;
  assign n13445 = n13443 & n13444;
  assign n13446 = n672 & n13442;
  assign n13447 = n1909 & n13446;
  assign n13448 = n1381 & n13445;
  assign n13449 = n12646 & n13448;
  assign n13450 = n13447 & n13449;
  assign n13451 = ~n269 & ~n421;
  assign n13452 = n537 & n13451;
  assign n13453 = ~n285 & ~n318;
  assign n13454 = ~n577 & n13453;
  assign n13455 = n114 & n1113;
  assign n13456 = n2314 & n13455;
  assign n13457 = n13452 & n13454;
  assign n13458 = n13456 & n13457;
  assign n13459 = ~n147 & ~n218;
  assign n13460 = ~n686 & n13459;
  assign n13461 = n1394 & n1458;
  assign n13462 = n1486 & n2822;
  assign n13463 = n2943 & n13462;
  assign n13464 = n13460 & n13461;
  assign n13465 = n2067 & n4788;
  assign n13466 = n13464 & n13465;
  assign n13467 = n13463 & n13466;
  assign n13468 = ~n280 & ~n479;
  assign n13469 = ~n661 & n13468;
  assign n13470 = n471 & n596;
  assign n13471 = n741 & n1281;
  assign n13472 = n2737 & n13471;
  assign n13473 = n13469 & n13470;
  assign n13474 = n1155 & n1310;
  assign n13475 = n3074 & n13474;
  assign n13476 = n13472 & n13473;
  assign n13477 = n4330 & n13476;
  assign n13478 = n13458 & n13475;
  assign n13479 = n13477 & n13478;
  assign n13480 = n13450 & n13467;
  assign n13481 = n13479 & n13480;
  assign n13482 = n3024 & n13481;
  assign n13483 = ~n145 & ~n512;
  assign n13484 = ~n539 & ~n702;
  assign n13485 = n13483 & n13484;
  assign n13486 = n919 & n2358;
  assign n13487 = n13485 & n13486;
  assign n13488 = n2495 & n13487;
  assign n13489 = n2732 & n13488;
  assign n13490 = ~n192 & ~n406;
  assign n13491 = ~n597 & n13490;
  assign n13492 = ~n213 & ~n318;
  assign n13493 = ~n545 & n13492;
  assign n13494 = ~n323 & n13491;
  assign n13495 = n13493 & n13494;
  assign n13496 = ~n203 & ~n216;
  assign n13497 = ~n385 & ~n511;
  assign n13498 = ~n642 & ~n644;
  assign n13499 = n13497 & n13498;
  assign n13500 = n804 & n13496;
  assign n13501 = n1160 & n1344;
  assign n13502 = n2474 & n13501;
  assign n13503 = n13499 & n13500;
  assign n13504 = n1586 & n5545;
  assign n13505 = n13503 & n13504;
  assign n13506 = n2632 & n13502;
  assign n13507 = n13505 & n13506;
  assign n13508 = n13495 & n13507;
  assign n13509 = n13489 & n13508;
  assign n13510 = n1941 & n3869;
  assign n13511 = n13509 & n13510;
  assign n13512 = ~n13482 & ~n13511;
  assign n13513 = ~n8939 & ~n9355;
  assign n13514 = ~n8196 & n13513;
  assign n13515 = ~n12163 & ~n13514;
  assign n13516 = pi8  & ~n13515;
  assign n13517 = ~pi8  & n13515;
  assign n13518 = ~n13516 & ~n13517;
  assign n13519 = n13482 & n13511;
  assign n13520 = ~n13512 & ~n13519;
  assign n13521 = n13518 & n13520;
  assign n13522 = ~n13512 & ~n13521;
  assign n13523 = n13336 & ~n13522;
  assign n13524 = ~n13336 & n13522;
  assign n13525 = ~n13523 & ~n13524;
  assign n13526 = n3896 & n12226;
  assign n13527 = n564 & n12232;
  assign n13528 = n3683 & n12229;
  assign n13529 = n12342 & ~n12344;
  assign n13530 = ~n12345 & ~n13529;
  assign n13531 = n566 & n13530;
  assign n13532 = ~n13527 & ~n13528;
  assign n13533 = ~n13526 & n13532;
  assign n13534 = ~n13531 & n13533;
  assign n13535 = n13525 & ~n13534;
  assign n13536 = ~n13523 & ~n13535;
  assign n13537 = ~n13336 & n13440;
  assign n13538 = ~n13441 & ~n13537;
  assign n13539 = ~n13536 & n13538;
  assign n13540 = ~n13441 & ~n13539;
  assign n13541 = ~n13387 & n13396;
  assign n13542 = ~n13397 & ~n13541;
  assign n13543 = ~n13540 & n13542;
  assign n13544 = ~n13397 & ~n13543;
  assign n13545 = ~n13369 & n13378;
  assign n13546 = ~n13379 & ~n13545;
  assign n13547 = ~n13544 & n13546;
  assign n13548 = n13544 & ~n13546;
  assign n13549 = ~n13547 & ~n13548;
  assign n13550 = n4472 & n12208;
  assign n13551 = n4070 & n12211;
  assign n13552 = n3943 & n12214;
  assign n13553 = n3944 & n12804;
  assign n13554 = ~n13551 & ~n13552;
  assign n13555 = ~n13550 & n13554;
  assign n13556 = ~n13553 & n13555;
  assign n13557 = pi29  & n13556;
  assign n13558 = ~pi29  & ~n13556;
  assign n13559 = ~n13557 & ~n13558;
  assign n13560 = n13549 & ~n13559;
  assign n13561 = ~n13547 & ~n13560;
  assign n13562 = n13385 & ~n13561;
  assign n13563 = ~n13383 & ~n13562;
  assign n13564 = n13295 & n13305;
  assign n13565 = ~n13306 & ~n13564;
  assign n13566 = ~n13563 & n13565;
  assign n13567 = ~n13306 & ~n13566;
  assign n13568 = ~n13212 & n13222;
  assign n13569 = ~n13223 & ~n13568;
  assign n13570 = ~n13567 & n13569;
  assign n13571 = n13567 & ~n13569;
  assign n13572 = ~n13570 & ~n13571;
  assign n13573 = n4721 & n12190;
  assign n13574 = n4691 & n12193;
  assign n13575 = n4515 & n12196;
  assign n13576 = n4516 & n12530;
  assign n13577 = ~n13574 & ~n13575;
  assign n13578 = ~n13573 & n13577;
  assign n13579 = ~n13576 & n13578;
  assign n13580 = pi26  & n13579;
  assign n13581 = ~pi26  & ~n13579;
  assign n13582 = ~n13580 & ~n13581;
  assign n13583 = n13572 & ~n13582;
  assign n13584 = ~n13570 & ~n13583;
  assign n13585 = ~n13229 & n13239;
  assign n13586 = ~n13240 & ~n13585;
  assign n13587 = ~n13584 & n13586;
  assign n13588 = n13584 & ~n13586;
  assign n13589 = ~n13587 & ~n13588;
  assign n13590 = n5267 & n12178;
  assign n13591 = n5185 & n12181;
  assign n13592 = n5121 & n12184;
  assign n13593 = n78 & n12880;
  assign n13594 = ~n13591 & ~n13592;
  assign n13595 = ~n13590 & n13594;
  assign n13596 = ~n13593 & n13595;
  assign n13597 = pi23  & n13596;
  assign n13598 = ~pi23  & ~n13596;
  assign n13599 = ~n13597 & ~n13598;
  assign n13600 = n13589 & ~n13599;
  assign n13601 = ~n13587 & ~n13600;
  assign n13602 = ~n13282 & n13292;
  assign n13603 = ~n13293 & ~n13602;
  assign n13604 = ~n13601 & n13603;
  assign n13605 = ~n13293 & ~n13604;
  assign n13606 = ~n13250 & n13260;
  assign n13607 = ~n13261 & ~n13606;
  assign n13608 = ~n13605 & n13607;
  assign n13609 = n13605 & ~n13607;
  assign n13610 = ~n13608 & ~n13609;
  assign n13611 = n5306 & n13007;
  assign n13612 = n5312 & n12172;
  assign n13613 = ~n5982 & n12165;
  assign n13614 = ~n12163 & ~n12513;
  assign n13615 = ~n13613 & n13614;
  assign n13616 = ~n13612 & ~n13615;
  assign n13617 = ~n13611 & n13616;
  assign n13618 = pi20  & n13617;
  assign n13619 = ~pi20  & ~n13617;
  assign n13620 = ~n13618 & ~n13619;
  assign n13621 = n13610 & ~n13620;
  assign n13622 = ~n13608 & ~n13621;
  assign n13623 = ~n13273 & ~n13275;
  assign n13624 = ~n13276 & ~n13623;
  assign n13625 = ~n13622 & n13624;
  assign n13626 = n13622 & ~n13624;
  assign n13627 = ~n13625 & ~n13626;
  assign n13628 = n13563 & ~n13565;
  assign n13629 = ~n13566 & ~n13628;
  assign n13630 = n4721 & n12193;
  assign n13631 = n4691 & n12196;
  assign n13632 = n4515 & n12199;
  assign n13633 = n4516 & n12594;
  assign n13634 = ~n13631 & ~n13632;
  assign n13635 = ~n13630 & n13634;
  assign n13636 = ~n13633 & n13635;
  assign n13637 = pi26  & n13636;
  assign n13638 = ~pi26  & ~n13636;
  assign n13639 = ~n13637 & ~n13638;
  assign n13640 = n13629 & ~n13639;
  assign n13641 = ~n13385 & n13561;
  assign n13642 = ~n13562 & ~n13641;
  assign n13643 = n4472 & n12205;
  assign n13644 = n4070 & n12208;
  assign n13645 = n3943 & n12211;
  assign n13646 = n3944 & n13031;
  assign n13647 = ~n13644 & ~n13645;
  assign n13648 = ~n13643 & n13647;
  assign n13649 = ~n13646 & n13648;
  assign n13650 = pi29  & n13649;
  assign n13651 = ~pi29  & ~n13649;
  assign n13652 = ~n13650 & ~n13651;
  assign n13653 = n13642 & ~n13652;
  assign n13654 = n4721 & n12196;
  assign n13655 = n4691 & n12199;
  assign n13656 = n4515 & n12202;
  assign n13657 = n4516 & n12578;
  assign n13658 = ~n13655 & ~n13656;
  assign n13659 = ~n13654 & n13658;
  assign n13660 = ~n13657 & n13659;
  assign n13661 = pi26  & n13660;
  assign n13662 = ~pi26  & ~n13660;
  assign n13663 = ~n13661 & ~n13662;
  assign n13664 = ~n13642 & n13652;
  assign n13665 = ~n13653 & ~n13664;
  assign n13666 = ~n13663 & n13665;
  assign n13667 = ~n13653 & ~n13666;
  assign n13668 = ~n13629 & n13639;
  assign n13669 = ~n13640 & ~n13668;
  assign n13670 = ~n13667 & n13669;
  assign n13671 = ~n13640 & ~n13670;
  assign n13672 = ~n13572 & n13582;
  assign n13673 = ~n13583 & ~n13672;
  assign n13674 = ~n13671 & n13673;
  assign n13675 = n13671 & ~n13673;
  assign n13676 = ~n13674 & ~n13675;
  assign n13677 = n5267 & n12181;
  assign n13678 = n5185 & n12184;
  assign n13679 = n5121 & n12187;
  assign n13680 = n78 & n12608;
  assign n13681 = ~n13678 & ~n13679;
  assign n13682 = ~n13677 & n13681;
  assign n13683 = ~n13680 & n13682;
  assign n13684 = pi23  & n13683;
  assign n13685 = ~pi23  & ~n13683;
  assign n13686 = ~n13684 & ~n13685;
  assign n13687 = n13676 & ~n13686;
  assign n13688 = ~n13674 & ~n13687;
  assign n13689 = ~n13589 & n13599;
  assign n13690 = ~n13600 & ~n13689;
  assign n13691 = ~n13688 & n13690;
  assign n13692 = n13688 & ~n13690;
  assign n13693 = ~n13691 & ~n13692;
  assign n13694 = n5982 & n12172;
  assign n13695 = n5901 & n12168;
  assign n13696 = n5312 & n12175;
  assign n13697 = n5306 & n12939;
  assign n13698 = ~n13695 & ~n13696;
  assign n13699 = ~n13694 & n13698;
  assign n13700 = ~n13697 & n13699;
  assign n13701 = pi20  & n13700;
  assign n13702 = ~pi20  & ~n13700;
  assign n13703 = ~n13701 & ~n13702;
  assign n13704 = n13693 & ~n13703;
  assign n13705 = ~n13691 & ~n13704;
  assign n13706 = n5982 & n12166;
  assign n13707 = n5901 & n12172;
  assign n13708 = n5312 & n12168;
  assign n13709 = n5306 & n13106;
  assign n13710 = ~n13706 & ~n13708;
  assign n13711 = ~n13707 & n13710;
  assign n13712 = ~n13709 & n13711;
  assign n13713 = pi20  & n13712;
  assign n13714 = ~pi20  & ~n13712;
  assign n13715 = ~n13713 & ~n13714;
  assign n13716 = ~n13705 & ~n13715;
  assign n13717 = n13601 & ~n13603;
  assign n13718 = ~n13604 & ~n13717;
  assign n13719 = n13705 & n13715;
  assign n13720 = ~n13716 & ~n13719;
  assign n13721 = n13718 & n13720;
  assign n13722 = ~n13716 & ~n13721;
  assign n13723 = ~n13610 & n13620;
  assign n13724 = ~n13621 & ~n13723;
  assign n13725 = ~n13722 & n13724;
  assign n13726 = n13667 & ~n13669;
  assign n13727 = ~n13670 & ~n13726;
  assign n13728 = n5267 & n12184;
  assign n13729 = n5185 & n12187;
  assign n13730 = n5121 & n12190;
  assign n13731 = n78 & n12845;
  assign n13732 = ~n13729 & ~n13730;
  assign n13733 = ~n13728 & n13732;
  assign n13734 = ~n13731 & n13733;
  assign n13735 = pi23  & n13734;
  assign n13736 = ~pi23  & ~n13734;
  assign n13737 = ~n13735 & ~n13736;
  assign n13738 = n13727 & ~n13737;
  assign n13739 = n13536 & ~n13538;
  assign n13740 = ~n13539 & ~n13739;
  assign n13741 = n3896 & n12223;
  assign n13742 = n3683 & n12226;
  assign n13743 = n564 & n12229;
  assign n13744 = n12346 & ~n12348;
  assign n13745 = ~n12349 & ~n13744;
  assign n13746 = n566 & n13745;
  assign n13747 = ~n13742 & ~n13743;
  assign n13748 = ~n13741 & n13747;
  assign n13749 = ~n13746 & n13748;
  assign n13750 = n13740 & ~n13749;
  assign n13751 = n4472 & n12214;
  assign n13752 = n4070 & n12217;
  assign n13753 = n3943 & n12220;
  assign n13754 = n3944 & n13187;
  assign n13755 = ~n13752 & ~n13753;
  assign n13756 = ~n13751 & n13755;
  assign n13757 = ~n13754 & n13756;
  assign n13758 = pi29  & n13757;
  assign n13759 = ~pi29  & ~n13757;
  assign n13760 = ~n13758 & ~n13759;
  assign n13761 = ~n13740 & n13749;
  assign n13762 = ~n13750 & ~n13761;
  assign n13763 = ~n13760 & n13762;
  assign n13764 = ~n13750 & ~n13763;
  assign n13765 = n13540 & ~n13542;
  assign n13766 = ~n13543 & ~n13765;
  assign n13767 = ~n13764 & n13766;
  assign n13768 = n4472 & n12211;
  assign n13769 = n4070 & n12214;
  assign n13770 = n3943 & n12217;
  assign n13771 = n3944 & n13203;
  assign n13772 = ~n13769 & ~n13770;
  assign n13773 = ~n13768 & n13772;
  assign n13774 = ~n13771 & n13773;
  assign n13775 = pi29  & n13774;
  assign n13776 = ~pi29  & ~n13774;
  assign n13777 = ~n13775 & ~n13776;
  assign n13778 = n13764 & ~n13766;
  assign n13779 = ~n13767 & ~n13778;
  assign n13780 = ~n13777 & n13779;
  assign n13781 = ~n13767 & ~n13780;
  assign n13782 = ~n13549 & n13559;
  assign n13783 = ~n13560 & ~n13782;
  assign n13784 = ~n13781 & n13783;
  assign n13785 = n13781 & ~n13783;
  assign n13786 = ~n13784 & ~n13785;
  assign n13787 = n4721 & n12199;
  assign n13788 = n4691 & n12202;
  assign n13789 = n4515 & n12205;
  assign n13790 = n4516 & n12683;
  assign n13791 = ~n13788 & ~n13789;
  assign n13792 = ~n13787 & n13791;
  assign n13793 = ~n13790 & n13792;
  assign n13794 = pi26  & n13793;
  assign n13795 = ~pi26  & ~n13793;
  assign n13796 = ~n13794 & ~n13795;
  assign n13797 = n13786 & ~n13796;
  assign n13798 = ~n13784 & ~n13797;
  assign n13799 = n13663 & ~n13665;
  assign n13800 = ~n13666 & ~n13799;
  assign n13801 = ~n13798 & n13800;
  assign n13802 = n13798 & ~n13800;
  assign n13803 = ~n13801 & ~n13802;
  assign n13804 = n5267 & n12187;
  assign n13805 = n5185 & n12190;
  assign n13806 = n5121 & n12193;
  assign n13807 = n78 & n12921;
  assign n13808 = ~n13805 & ~n13806;
  assign n13809 = ~n13804 & n13808;
  assign n13810 = ~n13807 & n13809;
  assign n13811 = pi23  & n13810;
  assign n13812 = ~pi23  & ~n13810;
  assign n13813 = ~n13811 & ~n13812;
  assign n13814 = n13803 & ~n13813;
  assign n13815 = ~n13801 & ~n13814;
  assign n13816 = ~n13727 & n13737;
  assign n13817 = ~n13738 & ~n13816;
  assign n13818 = ~n13815 & n13817;
  assign n13819 = ~n13738 & ~n13818;
  assign n13820 = ~n13676 & n13686;
  assign n13821 = ~n13687 & ~n13820;
  assign n13822 = ~n13819 & n13821;
  assign n13823 = n13819 & ~n13821;
  assign n13824 = ~n13822 & ~n13823;
  assign n13825 = n5982 & n12168;
  assign n13826 = n5901 & n12175;
  assign n13827 = n5312 & n12178;
  assign n13828 = n5306 & n12862;
  assign n13829 = ~n13826 & ~n13827;
  assign n13830 = ~n13825 & n13829;
  assign n13831 = ~n13828 & n13830;
  assign n13832 = pi20  & n13831;
  assign n13833 = ~pi20  & ~n13831;
  assign n13834 = ~n13832 & ~n13833;
  assign n13835 = n13824 & ~n13834;
  assign n13836 = ~n13822 & ~n13835;
  assign n13837 = n6134 & ~n12424;
  assign n13838 = n6140 & ~n12165;
  assign n13839 = n12666 & ~n13838;
  assign n13840 = ~n12163 & ~n13839;
  assign n13841 = ~n13837 & ~n13840;
  assign n13842 = pi17  & n13841;
  assign n13843 = ~pi17  & ~n13841;
  assign n13844 = ~n13842 & ~n13843;
  assign n13845 = ~n13836 & ~n13844;
  assign n13846 = n13836 & n13844;
  assign n13847 = ~n13845 & ~n13846;
  assign n13848 = ~n13693 & n13703;
  assign n13849 = ~n13704 & ~n13848;
  assign n13850 = n13847 & n13849;
  assign n13851 = ~n13845 & ~n13850;
  assign n13852 = ~n13718 & ~n13720;
  assign n13853 = ~n13721 & ~n13852;
  assign n13854 = ~n13851 & n13853;
  assign n13855 = n13815 & ~n13817;
  assign n13856 = ~n13818 & ~n13855;
  assign n13857 = n5982 & n12175;
  assign n13858 = n5901 & n12178;
  assign n13859 = n5312 & n12181;
  assign n13860 = n5306 & n12961;
  assign n13861 = ~n13858 & ~n13859;
  assign n13862 = ~n13857 & n13861;
  assign n13863 = ~n13860 & n13862;
  assign n13864 = pi20  & n13863;
  assign n13865 = ~pi20  & ~n13863;
  assign n13866 = ~n13864 & ~n13865;
  assign n13867 = n13856 & ~n13866;
  assign n13868 = n4721 & n12202;
  assign n13869 = n4691 & n12205;
  assign n13870 = n4515 & n12208;
  assign n13871 = n4516 & n12701;
  assign n13872 = ~n13869 & ~n13870;
  assign n13873 = ~n13868 & n13872;
  assign n13874 = ~n13871 & n13873;
  assign n13875 = pi26  & n13874;
  assign n13876 = ~pi26  & ~n13874;
  assign n13877 = ~n13875 & ~n13876;
  assign n13878 = n13777 & ~n13779;
  assign n13879 = ~n13780 & ~n13878;
  assign n13880 = ~n13877 & n13879;
  assign n13881 = ~n270 & n1965;
  assign n13882 = ~n467 & n13881;
  assign n13883 = ~n147 & ~n407;
  assign n13884 = ~n583 & ~n590;
  assign n13885 = ~n642 & n13884;
  assign n13886 = n166 & n13883;
  assign n13887 = n211 & n1399;
  assign n13888 = n2785 & n13887;
  assign n13889 = n13885 & n13886;
  assign n13890 = n5724 & n13491;
  assign n13891 = n13889 & n13890;
  assign n13892 = n1076 & n13888;
  assign n13893 = n13882 & n13892;
  assign n13894 = n1052 & n13891;
  assign n13895 = n13893 & n13894;
  assign n13896 = n2594 & n13895;
  assign n13897 = n2685 & n13896;
  assign n13898 = n13482 & ~n13897;
  assign n13899 = n10879 & ~n10882;
  assign n13900 = ~pi2  & ~n13899;
  assign n13901 = ~n12163 & n13900;
  assign n13902 = pi2  & n12163;
  assign n13903 = ~n13901 & ~n13902;
  assign n13904 = ~n109 & ~n177;
  assign n13905 = ~n319 & ~n385;
  assign n13906 = ~n391 & ~n482;
  assign n13907 = ~n679 & n13906;
  assign n13908 = n13904 & n13905;
  assign n13909 = n1301 & n1472;
  assign n13910 = n1909 & n2450;
  assign n13911 = n3872 & n13910;
  assign n13912 = n13908 & n13909;
  assign n13913 = n13907 & n13912;
  assign n13914 = n1026 & n13911;
  assign n13915 = n13913 & n13914;
  assign n13916 = ~n407 & ~n646;
  assign n13917 = n1203 & n13916;
  assign n13918 = n13412 & n13917;
  assign n13919 = n237 & ~n362;
  assign n13920 = n1356 & n13919;
  assign n13921 = n1341 & n2924;
  assign n13922 = n4361 & n12765;
  assign n13923 = n13921 & n13922;
  assign n13924 = n3998 & n13920;
  assign n13925 = n13918 & n13924;
  assign n13926 = n3288 & n13923;
  assign n13927 = n13925 & n13926;
  assign n13928 = n13915 & n13927;
  assign n13929 = ~n374 & ~n599;
  assign n13930 = n922 & n13929;
  assign n13931 = n1349 & n2272;
  assign n13932 = n3267 & n4093;
  assign n13933 = n13931 & n13932;
  assign n13934 = n4359 & n13930;
  assign n13935 = n13933 & n13934;
  assign n13936 = n6475 & n6980;
  assign n13937 = n13935 & n13936;
  assign n13938 = n4201 & n13320;
  assign n13939 = n13937 & n13938;
  assign n13940 = n13928 & n13939;
  assign n13941 = n13903 & ~n13940;
  assign n13942 = ~n71 & ~n10329;
  assign n13943 = ~n70 & n13942;
  assign n13944 = ~n12163 & ~n13943;
  assign n13945 = ~pi5  & n13944;
  assign n13946 = pi5  & ~n13944;
  assign n13947 = ~n13945 & ~n13946;
  assign n13948 = ~n13903 & n13940;
  assign n13949 = ~n13941 & ~n13948;
  assign n13950 = n13947 & n13949;
  assign n13951 = ~n13941 & ~n13950;
  assign n13952 = n13482 & ~n13951;
  assign n13953 = ~n13482 & n13951;
  assign n13954 = ~n13952 & ~n13953;
  assign n13955 = n3896 & n12235;
  assign n13956 = n564 & n12241;
  assign n13957 = n3683 & n12238;
  assign n13958 = n12330 & ~n12332;
  assign n13959 = ~n12333 & ~n13958;
  assign n13960 = n566 & n13959;
  assign n13961 = ~n13956 & ~n13957;
  assign n13962 = ~n13955 & n13961;
  assign n13963 = ~n13960 & n13962;
  assign n13964 = n13954 & ~n13963;
  assign n13965 = ~n13952 & ~n13964;
  assign n13966 = ~n13482 & n13897;
  assign n13967 = ~n13898 & ~n13966;
  assign n13968 = ~n13965 & n13967;
  assign n13969 = ~n13898 & ~n13968;
  assign n13970 = ~n13518 & ~n13520;
  assign n13971 = ~n13521 & ~n13970;
  assign n13972 = ~n13969 & n13971;
  assign n13973 = n13969 & ~n13971;
  assign n13974 = ~n13972 & ~n13973;
  assign n13975 = n3896 & n12229;
  assign n13976 = n3683 & n12232;
  assign n13977 = n564 & n12235;
  assign n13978 = n12338 & ~n12340;
  assign n13979 = ~n12341 & ~n13978;
  assign n13980 = n566 & n13979;
  assign n13981 = ~n13976 & ~n13977;
  assign n13982 = ~n13975 & n13981;
  assign n13983 = ~n13980 & n13982;
  assign n13984 = n13974 & ~n13983;
  assign n13985 = ~n13972 & ~n13984;
  assign n13986 = ~n13525 & n13534;
  assign n13987 = ~n13535 & ~n13986;
  assign n13988 = ~n13985 & n13987;
  assign n13989 = n13985 & ~n13987;
  assign n13990 = ~n13988 & ~n13989;
  assign n13991 = n4472 & n12217;
  assign n13992 = n4070 & n12220;
  assign n13993 = n3943 & n12223;
  assign n13994 = n3944 & n13374;
  assign n13995 = ~n13992 & ~n13993;
  assign n13996 = ~n13991 & n13995;
  assign n13997 = ~n13994 & n13996;
  assign n13998 = pi29  & n13997;
  assign n13999 = ~pi29  & ~n13997;
  assign n14000 = ~n13998 & ~n13999;
  assign n14001 = n13990 & ~n14000;
  assign n14002 = ~n13988 & ~n14001;
  assign n14003 = n13760 & ~n13762;
  assign n14004 = ~n13763 & ~n14003;
  assign n14005 = ~n14002 & n14004;
  assign n14006 = n14002 & ~n14004;
  assign n14007 = ~n14005 & ~n14006;
  assign n14008 = n4721 & n12205;
  assign n14009 = n4691 & n12208;
  assign n14010 = n4515 & n12211;
  assign n14011 = n4516 & n13031;
  assign n14012 = ~n14009 & ~n14010;
  assign n14013 = ~n14008 & n14012;
  assign n14014 = ~n14011 & n14013;
  assign n14015 = pi26  & n14014;
  assign n14016 = ~pi26  & ~n14014;
  assign n14017 = ~n14015 & ~n14016;
  assign n14018 = n14007 & ~n14017;
  assign n14019 = ~n14005 & ~n14018;
  assign n14020 = n13877 & ~n13879;
  assign n14021 = ~n13880 & ~n14020;
  assign n14022 = ~n14019 & n14021;
  assign n14023 = ~n13880 & ~n14022;
  assign n14024 = ~n13786 & n13796;
  assign n14025 = ~n13797 & ~n14024;
  assign n14026 = ~n14023 & n14025;
  assign n14027 = n14023 & ~n14025;
  assign n14028 = ~n14026 & ~n14027;
  assign n14029 = n5267 & n12190;
  assign n14030 = n5185 & n12193;
  assign n14031 = n5121 & n12196;
  assign n14032 = n78 & n12530;
  assign n14033 = ~n14030 & ~n14031;
  assign n14034 = ~n14029 & n14033;
  assign n14035 = ~n14032 & n14034;
  assign n14036 = pi23  & n14035;
  assign n14037 = ~pi23  & ~n14035;
  assign n14038 = ~n14036 & ~n14037;
  assign n14039 = n14028 & ~n14038;
  assign n14040 = ~n14026 & ~n14039;
  assign n14041 = ~n13803 & n13813;
  assign n14042 = ~n13814 & ~n14041;
  assign n14043 = ~n14040 & n14042;
  assign n14044 = n14040 & ~n14042;
  assign n14045 = ~n14043 & ~n14044;
  assign n14046 = n5982 & n12178;
  assign n14047 = n5901 & n12181;
  assign n14048 = n5312 & n12184;
  assign n14049 = n5306 & n12880;
  assign n14050 = ~n14047 & ~n14048;
  assign n14051 = ~n14046 & n14050;
  assign n14052 = ~n14049 & n14051;
  assign n14053 = pi20  & n14052;
  assign n14054 = ~pi20  & ~n14052;
  assign n14055 = ~n14053 & ~n14054;
  assign n14056 = n14045 & ~n14055;
  assign n14057 = ~n14043 & ~n14056;
  assign n14058 = ~n13856 & n13866;
  assign n14059 = ~n13867 & ~n14058;
  assign n14060 = ~n14057 & n14059;
  assign n14061 = ~n13867 & ~n14060;
  assign n14062 = ~n13824 & n13834;
  assign n14063 = ~n13835 & ~n14062;
  assign n14064 = ~n14061 & n14063;
  assign n14065 = n14061 & ~n14063;
  assign n14066 = ~n14064 & ~n14065;
  assign n14067 = n6134 & n13007;
  assign n14068 = n6140 & n12172;
  assign n14069 = ~n6608 & n12165;
  assign n14070 = ~n12163 & ~n12666;
  assign n14071 = ~n14069 & n14070;
  assign n14072 = ~n14068 & ~n14071;
  assign n14073 = ~n14067 & n14072;
  assign n14074 = pi17  & n14073;
  assign n14075 = ~pi17  & ~n14073;
  assign n14076 = ~n14074 & ~n14075;
  assign n14077 = n14066 & ~n14076;
  assign n14078 = ~n14064 & ~n14077;
  assign n14079 = ~n13847 & ~n13849;
  assign n14080 = ~n13850 & ~n14079;
  assign n14081 = ~n14078 & n14080;
  assign n14082 = n14078 & ~n14080;
  assign n14083 = ~n14081 & ~n14082;
  assign n14084 = n14019 & ~n14021;
  assign n14085 = ~n14022 & ~n14084;
  assign n14086 = n5267 & n12193;
  assign n14087 = n5185 & n12196;
  assign n14088 = n5121 & n12199;
  assign n14089 = n78 & n12594;
  assign n14090 = ~n14087 & ~n14088;
  assign n14091 = ~n14086 & n14090;
  assign n14092 = ~n14089 & n14091;
  assign n14093 = pi23  & n14092;
  assign n14094 = ~pi23  & ~n14092;
  assign n14095 = ~n14093 & ~n14094;
  assign n14096 = n14085 & ~n14095;
  assign n14097 = n4472 & n12220;
  assign n14098 = n4070 & n12223;
  assign n14099 = n3943 & n12226;
  assign n14100 = n3944 & n13392;
  assign n14101 = ~n14098 & ~n14099;
  assign n14102 = ~n14097 & n14101;
  assign n14103 = ~n14100 & n14102;
  assign n14104 = pi29  & n14103;
  assign n14105 = ~pi29  & ~n14103;
  assign n14106 = ~n14104 & ~n14105;
  assign n14107 = ~n13974 & n13983;
  assign n14108 = ~n13984 & ~n14107;
  assign n14109 = ~n14106 & n14108;
  assign n14110 = n13965 & ~n13967;
  assign n14111 = ~n13968 & ~n14110;
  assign n14112 = n3896 & n12232;
  assign n14113 = n3683 & n12235;
  assign n14114 = n564 & n12238;
  assign n14115 = n12334 & ~n12336;
  assign n14116 = ~n12337 & ~n14115;
  assign n14117 = n566 & n14116;
  assign n14118 = ~n14113 & ~n14114;
  assign n14119 = ~n14112 & n14118;
  assign n14120 = ~n14117 & n14119;
  assign n14121 = n14111 & ~n14120;
  assign n14122 = ~n163 & ~n219;
  assign n14123 = ~n283 & ~n648;
  assign n14124 = n14122 & n14123;
  assign n14125 = n1281 & n2630;
  assign n14126 = n2786 & n2981;
  assign n14127 = n4795 & n12766;
  assign n14128 = n14126 & n14127;
  assign n14129 = n14124 & n14125;
  assign n14130 = n14128 & n14129;
  assign n14131 = n2007 & n3432;
  assign n14132 = n14130 & n14131;
  assign n14133 = n3793 & n14132;
  assign n14134 = n867 & n14133;
  assign n14135 = n4127 & n14134;
  assign n14136 = ~n13903 & ~n14135;
  assign n14137 = ~n568 & n1233;
  assign n14138 = n12716 & n14137;
  assign n14139 = ~n467 & ~n554;
  assign n14140 = n194 & n14139;
  assign n14141 = n1354 & n2047;
  assign n14142 = n2472 & n2706;
  assign n14143 = n4767 & n12458;
  assign n14144 = n14142 & n14143;
  assign n14145 = n14140 & n14141;
  assign n14146 = n358 & n2697;
  assign n14147 = n14145 & n14146;
  assign n14148 = n12125 & n14144;
  assign n14149 = n14138 & n14148;
  assign n14150 = n1463 & n14147;
  assign n14151 = n1688 & n14150;
  assign n14152 = n14149 & n14151;
  assign n14153 = n13928 & n14152;
  assign n14154 = ~n13903 & ~n14153;
  assign n14155 = n13903 & n14153;
  assign n14156 = ~n14154 & ~n14155;
  assign n14157 = ~n277 & ~n541;
  assign n14158 = ~n587 & ~n650;
  assign n14159 = ~n662 & n14158;
  assign n14160 = n6939 & n14157;
  assign n14161 = n14159 & n14160;
  assign n14162 = n948 & n14161;
  assign n14163 = ~n312 & ~n360;
  assign n14164 = ~n445 & n14163;
  assign n14165 = n2297 & n2959;
  assign n14166 = n5751 & n14165;
  assign n14167 = n14164 & n14166;
  assign n14168 = ~n222 & ~n363;
  assign n14169 = ~n402 & ~n538;
  assign n14170 = ~n702 & n14169;
  assign n14171 = n524 & n14168;
  assign n14172 = n1339 & n2060;
  assign n14173 = n3155 & n14172;
  assign n14174 = n14170 & n14171;
  assign n14175 = n3611 & n4204;
  assign n14176 = n14174 & n14175;
  assign n14177 = n14173 & n14176;
  assign n14178 = n2449 & n14167;
  assign n14179 = n14177 & n14178;
  assign n14180 = ~n172 & ~n374;
  assign n14181 = ~n679 & n2236;
  assign n14182 = n2474 & n14180;
  assign n14183 = n14181 & n14182;
  assign n14184 = n14179 & n14183;
  assign n14185 = ~n539 & ~n676;
  assign n14186 = ~n163 & ~n269;
  assign n14187 = ~n285 & ~n300;
  assign n14188 = ~n701 & n14187;
  assign n14189 = n1487 & n14186;
  assign n14190 = n2150 & n3380;
  assign n14191 = n14185 & n14190;
  assign n14192 = n14188 & n14189;
  assign n14193 = n2268 & n13412;
  assign n14194 = n14192 & n14193;
  assign n14195 = n2520 & n14191;
  assign n14196 = n14194 & n14195;
  assign n14197 = n14162 & n14196;
  assign n14198 = n12553 & n14197;
  assign n14199 = n14184 & n14198;
  assign n14200 = n13903 & n14199;
  assign n14201 = ~n13903 & ~n14199;
  assign n14202 = ~n14200 & ~n14201;
  assign n14203 = n3896 & n12247;
  assign n14204 = n3683 & n12250;
  assign n14205 = n564 & n12253;
  assign n14206 = n12314 & ~n12316;
  assign n14207 = ~n12317 & ~n14206;
  assign n14208 = n566 & n14207;
  assign n14209 = ~n14204 & ~n14205;
  assign n14210 = ~n14203 & n14209;
  assign n14211 = ~n14208 & n14210;
  assign n14212 = n14202 & n14211;
  assign n14213 = ~n14200 & ~n14212;
  assign n14214 = n14156 & n14213;
  assign n14215 = ~n14154 & ~n14214;
  assign n14216 = n13903 & n14135;
  assign n14217 = ~n14136 & ~n14216;
  assign n14218 = ~n14215 & n14217;
  assign n14219 = ~n14136 & ~n14218;
  assign n14220 = ~n13947 & ~n13949;
  assign n14221 = ~n13950 & ~n14220;
  assign n14222 = ~n14219 & n14221;
  assign n14223 = n14219 & ~n14221;
  assign n14224 = ~n14222 & ~n14223;
  assign n14225 = n3896 & n12238;
  assign n14226 = n3683 & n12241;
  assign n14227 = n564 & n12244;
  assign n14228 = n12326 & ~n12328;
  assign n14229 = ~n12329 & ~n14228;
  assign n14230 = n566 & n14229;
  assign n14231 = ~n14226 & ~n14227;
  assign n14232 = ~n14225 & n14231;
  assign n14233 = ~n14230 & n14232;
  assign n14234 = n14224 & ~n14233;
  assign n14235 = ~n14222 & ~n14234;
  assign n14236 = ~n13954 & n13963;
  assign n14237 = ~n13964 & ~n14236;
  assign n14238 = ~n14235 & n14237;
  assign n14239 = n14235 & ~n14237;
  assign n14240 = ~n14238 & ~n14239;
  assign n14241 = n4472 & n12226;
  assign n14242 = n4070 & n12229;
  assign n14243 = n3943 & n12232;
  assign n14244 = n3944 & n13530;
  assign n14245 = ~n14242 & ~n14243;
  assign n14246 = ~n14241 & n14245;
  assign n14247 = ~n14244 & n14246;
  assign n14248 = pi29  & n14247;
  assign n14249 = ~pi29  & ~n14247;
  assign n14250 = ~n14248 & ~n14249;
  assign n14251 = n14240 & ~n14250;
  assign n14252 = ~n14238 & ~n14251;
  assign n14253 = ~n14111 & n14120;
  assign n14254 = ~n14121 & ~n14253;
  assign n14255 = ~n14252 & n14254;
  assign n14256 = ~n14121 & ~n14255;
  assign n14257 = n14106 & ~n14108;
  assign n14258 = ~n14109 & ~n14257;
  assign n14259 = ~n14256 & n14258;
  assign n14260 = ~n14109 & ~n14259;
  assign n14261 = ~n13990 & n14000;
  assign n14262 = ~n14001 & ~n14261;
  assign n14263 = ~n14260 & n14262;
  assign n14264 = n14260 & ~n14262;
  assign n14265 = ~n14263 & ~n14264;
  assign n14266 = n4721 & n12208;
  assign n14267 = n4691 & n12211;
  assign n14268 = n4515 & n12214;
  assign n14269 = n4516 & n12804;
  assign n14270 = ~n14267 & ~n14268;
  assign n14271 = ~n14266 & n14270;
  assign n14272 = ~n14269 & n14271;
  assign n14273 = pi26  & n14272;
  assign n14274 = ~pi26  & ~n14272;
  assign n14275 = ~n14273 & ~n14274;
  assign n14276 = n14265 & ~n14275;
  assign n14277 = ~n14263 & ~n14276;
  assign n14278 = ~n14007 & n14017;
  assign n14279 = ~n14018 & ~n14278;
  assign n14280 = ~n14277 & n14279;
  assign n14281 = n14277 & ~n14279;
  assign n14282 = ~n14280 & ~n14281;
  assign n14283 = n5267 & n12196;
  assign n14284 = n5185 & n12199;
  assign n14285 = n5121 & n12202;
  assign n14286 = n78 & n12578;
  assign n14287 = ~n14284 & ~n14285;
  assign n14288 = ~n14283 & n14287;
  assign n14289 = ~n14286 & n14288;
  assign n14290 = pi23  & n14289;
  assign n14291 = ~pi23  & ~n14289;
  assign n14292 = ~n14290 & ~n14291;
  assign n14293 = n14282 & ~n14292;
  assign n14294 = ~n14280 & ~n14293;
  assign n14295 = ~n14085 & n14095;
  assign n14296 = ~n14096 & ~n14295;
  assign n14297 = ~n14294 & n14296;
  assign n14298 = ~n14096 & ~n14297;
  assign n14299 = ~n14028 & n14038;
  assign n14300 = ~n14039 & ~n14299;
  assign n14301 = ~n14298 & n14300;
  assign n14302 = n14298 & ~n14300;
  assign n14303 = ~n14301 & ~n14302;
  assign n14304 = n5982 & n12181;
  assign n14305 = n5901 & n12184;
  assign n14306 = n5312 & n12187;
  assign n14307 = n5306 & n12608;
  assign n14308 = ~n14305 & ~n14306;
  assign n14309 = ~n14304 & n14308;
  assign n14310 = ~n14307 & n14309;
  assign n14311 = pi20  & n14310;
  assign n14312 = ~pi20  & ~n14310;
  assign n14313 = ~n14311 & ~n14312;
  assign n14314 = n14303 & ~n14313;
  assign n14315 = ~n14301 & ~n14314;
  assign n14316 = ~n14045 & n14055;
  assign n14317 = ~n14056 & ~n14316;
  assign n14318 = ~n14315 & n14317;
  assign n14319 = n14315 & ~n14317;
  assign n14320 = ~n14318 & ~n14319;
  assign n14321 = n6608 & n12172;
  assign n14322 = n6356 & n12168;
  assign n14323 = n6140 & n12175;
  assign n14324 = n6134 & n12939;
  assign n14325 = ~n14322 & ~n14323;
  assign n14326 = ~n14321 & n14325;
  assign n14327 = ~n14324 & n14326;
  assign n14328 = pi17  & n14327;
  assign n14329 = ~pi17  & ~n14327;
  assign n14330 = ~n14328 & ~n14329;
  assign n14331 = n14320 & ~n14330;
  assign n14332 = ~n14318 & ~n14331;
  assign n14333 = n6608 & n12166;
  assign n14334 = n6356 & n12172;
  assign n14335 = n6140 & n12168;
  assign n14336 = n6134 & n13106;
  assign n14337 = ~n14333 & ~n14335;
  assign n14338 = ~n14334 & n14337;
  assign n14339 = ~n14336 & n14338;
  assign n14340 = pi17  & n14339;
  assign n14341 = ~pi17  & ~n14339;
  assign n14342 = ~n14340 & ~n14341;
  assign n14343 = ~n14332 & ~n14342;
  assign n14344 = n14057 & ~n14059;
  assign n14345 = ~n14060 & ~n14344;
  assign n14346 = n14332 & n14342;
  assign n14347 = ~n14343 & ~n14346;
  assign n14348 = n14345 & n14347;
  assign n14349 = ~n14343 & ~n14348;
  assign n14350 = ~n14066 & n14076;
  assign n14351 = ~n14077 & ~n14350;
  assign n14352 = ~n14349 & n14351;
  assign n14353 = n14294 & ~n14296;
  assign n14354 = ~n14297 & ~n14353;
  assign n14355 = n5982 & n12184;
  assign n14356 = n5901 & n12187;
  assign n14357 = n5312 & n12190;
  assign n14358 = n5306 & n12845;
  assign n14359 = ~n14356 & ~n14357;
  assign n14360 = ~n14355 & n14359;
  assign n14361 = ~n14358 & n14360;
  assign n14362 = pi20  & n14361;
  assign n14363 = ~pi20  & ~n14361;
  assign n14364 = ~n14362 & ~n14363;
  assign n14365 = n14354 & ~n14364;
  assign n14366 = n14256 & ~n14258;
  assign n14367 = ~n14259 & ~n14366;
  assign n14368 = n4721 & n12211;
  assign n14369 = n4691 & n12214;
  assign n14370 = n4515 & n12217;
  assign n14371 = n4516 & n13203;
  assign n14372 = ~n14369 & ~n14370;
  assign n14373 = ~n14368 & n14372;
  assign n14374 = ~n14371 & n14373;
  assign n14375 = pi26  & n14374;
  assign n14376 = ~pi26  & ~n14374;
  assign n14377 = ~n14375 & ~n14376;
  assign n14378 = n14367 & ~n14377;
  assign n14379 = n14252 & ~n14254;
  assign n14380 = ~n14255 & ~n14379;
  assign n14381 = n4472 & n12223;
  assign n14382 = n4070 & n12226;
  assign n14383 = n3943 & n12229;
  assign n14384 = n3944 & n13745;
  assign n14385 = ~n14382 & ~n14383;
  assign n14386 = ~n14381 & n14385;
  assign n14387 = ~n14384 & n14386;
  assign n14388 = pi29  & n14387;
  assign n14389 = ~pi29  & ~n14387;
  assign n14390 = ~n14388 & ~n14389;
  assign n14391 = n14380 & ~n14390;
  assign n14392 = n4721 & n12214;
  assign n14393 = n4691 & n12217;
  assign n14394 = n4515 & n12220;
  assign n14395 = n4516 & n13187;
  assign n14396 = ~n14393 & ~n14394;
  assign n14397 = ~n14392 & n14396;
  assign n14398 = ~n14395 & n14397;
  assign n14399 = pi26  & n14398;
  assign n14400 = ~pi26  & ~n14398;
  assign n14401 = ~n14399 & ~n14400;
  assign n14402 = ~n14380 & n14390;
  assign n14403 = ~n14391 & ~n14402;
  assign n14404 = ~n14401 & n14403;
  assign n14405 = ~n14391 & ~n14404;
  assign n14406 = ~n14367 & n14377;
  assign n14407 = ~n14378 & ~n14406;
  assign n14408 = ~n14405 & n14407;
  assign n14409 = ~n14378 & ~n14408;
  assign n14410 = ~n14265 & n14275;
  assign n14411 = ~n14276 & ~n14410;
  assign n14412 = ~n14409 & n14411;
  assign n14413 = n14409 & ~n14411;
  assign n14414 = ~n14412 & ~n14413;
  assign n14415 = n5267 & n12199;
  assign n14416 = n5185 & n12202;
  assign n14417 = n5121 & n12205;
  assign n14418 = n78 & n12683;
  assign n14419 = ~n14416 & ~n14417;
  assign n14420 = ~n14415 & n14419;
  assign n14421 = ~n14418 & n14420;
  assign n14422 = pi23  & n14421;
  assign n14423 = ~pi23  & ~n14421;
  assign n14424 = ~n14422 & ~n14423;
  assign n14425 = n14414 & ~n14424;
  assign n14426 = ~n14412 & ~n14425;
  assign n14427 = ~n14282 & n14292;
  assign n14428 = ~n14293 & ~n14427;
  assign n14429 = ~n14426 & n14428;
  assign n14430 = n14426 & ~n14428;
  assign n14431 = ~n14429 & ~n14430;
  assign n14432 = n5982 & n12187;
  assign n14433 = n5901 & n12190;
  assign n14434 = n5312 & n12193;
  assign n14435 = n5306 & n12921;
  assign n14436 = ~n14433 & ~n14434;
  assign n14437 = ~n14432 & n14436;
  assign n14438 = ~n14435 & n14437;
  assign n14439 = pi20  & n14438;
  assign n14440 = ~pi20  & ~n14438;
  assign n14441 = ~n14439 & ~n14440;
  assign n14442 = n14431 & ~n14441;
  assign n14443 = ~n14429 & ~n14442;
  assign n14444 = ~n14354 & n14364;
  assign n14445 = ~n14365 & ~n14444;
  assign n14446 = ~n14443 & n14445;
  assign n14447 = ~n14365 & ~n14446;
  assign n14448 = ~n14303 & n14313;
  assign n14449 = ~n14314 & ~n14448;
  assign n14450 = ~n14447 & n14449;
  assign n14451 = n14447 & ~n14449;
  assign n14452 = ~n14450 & ~n14451;
  assign n14453 = n6608 & n12168;
  assign n14454 = n6356 & n12175;
  assign n14455 = n6140 & n12178;
  assign n14456 = n6134 & n12862;
  assign n14457 = ~n14454 & ~n14455;
  assign n14458 = ~n14453 & n14457;
  assign n14459 = ~n14456 & n14458;
  assign n14460 = pi17  & n14459;
  assign n14461 = ~pi17  & ~n14459;
  assign n14462 = ~n14460 & ~n14461;
  assign n14463 = n14452 & ~n14462;
  assign n14464 = ~n14450 & ~n14463;
  assign n14465 = n6647 & ~n12424;
  assign n14466 = n6652 & ~n12165;
  assign n14467 = n12787 & ~n14466;
  assign n14468 = ~n12163 & ~n14467;
  assign n14469 = ~n14465 & ~n14468;
  assign n14470 = pi14  & n14469;
  assign n14471 = ~pi14  & ~n14469;
  assign n14472 = ~n14470 & ~n14471;
  assign n14473 = ~n14464 & ~n14472;
  assign n14474 = n14464 & n14472;
  assign n14475 = ~n14473 & ~n14474;
  assign n14476 = ~n14320 & n14330;
  assign n14477 = ~n14331 & ~n14476;
  assign n14478 = n14475 & n14477;
  assign n14479 = ~n14473 & ~n14478;
  assign n14480 = ~n14345 & ~n14347;
  assign n14481 = ~n14348 & ~n14480;
  assign n14482 = ~n14479 & n14481;
  assign n14483 = n14443 & ~n14445;
  assign n14484 = ~n14446 & ~n14483;
  assign n14485 = n6608 & n12175;
  assign n14486 = n6356 & n12178;
  assign n14487 = n6140 & n12181;
  assign n14488 = n6134 & n12961;
  assign n14489 = ~n14486 & ~n14487;
  assign n14490 = ~n14485 & n14489;
  assign n14491 = ~n14488 & n14490;
  assign n14492 = pi17  & n14491;
  assign n14493 = ~pi17  & ~n14491;
  assign n14494 = ~n14492 & ~n14493;
  assign n14495 = n14484 & ~n14494;
  assign n14496 = n14405 & ~n14407;
  assign n14497 = ~n14408 & ~n14496;
  assign n14498 = n5267 & n12202;
  assign n14499 = n5185 & n12205;
  assign n14500 = n5121 & n12208;
  assign n14501 = n78 & n12701;
  assign n14502 = ~n14499 & ~n14500;
  assign n14503 = ~n14498 & n14502;
  assign n14504 = ~n14501 & n14503;
  assign n14505 = pi23  & n14504;
  assign n14506 = ~pi23  & ~n14504;
  assign n14507 = ~n14505 & ~n14506;
  assign n14508 = n14497 & ~n14507;
  assign n14509 = n14215 & ~n14217;
  assign n14510 = ~n14218 & ~n14509;
  assign n14511 = n3896 & n12241;
  assign n14512 = n3683 & n12244;
  assign n14513 = n564 & n12247;
  assign n14514 = n12322 & ~n12324;
  assign n14515 = ~n12325 & ~n14514;
  assign n14516 = n566 & n14515;
  assign n14517 = ~n14512 & ~n14513;
  assign n14518 = ~n14511 & n14517;
  assign n14519 = ~n14516 & n14518;
  assign n14520 = n14510 & ~n14519;
  assign n14521 = ~n14156 & ~n14213;
  assign n14522 = ~n14214 & ~n14521;
  assign n14523 = n3896 & n12244;
  assign n14524 = n3683 & n12247;
  assign n14525 = n564 & n12250;
  assign n14526 = n12318 & ~n12320;
  assign n14527 = ~n12321 & ~n14526;
  assign n14528 = n566 & n14527;
  assign n14529 = ~n14524 & ~n14525;
  assign n14530 = ~n14523 & n14529;
  assign n14531 = ~n14528 & n14530;
  assign n14532 = n14522 & ~n14531;
  assign n14533 = ~n14202 & ~n14211;
  assign n14534 = ~n14212 & ~n14533;
  assign n14535 = ~n207 & ~n218;
  assign n14536 = ~n245 & ~n577;
  assign n14537 = ~n597 & n14536;
  assign n14538 = n14535 & n14537;
  assign n14539 = n3971 & n14538;
  assign n14540 = ~n338 & ~n521;
  assign n14541 = ~n594 & n14540;
  assign n14542 = n969 & n1284;
  assign n14543 = n1125 & n1175;
  assign n14544 = n1246 & n3381;
  assign n14545 = n14543 & n14544;
  assign n14546 = n14541 & n14542;
  assign n14547 = n3425 & n14546;
  assign n14548 = n2956 & n14545;
  assign n14549 = n4382 & n13310;
  assign n14550 = n14548 & n14549;
  assign n14551 = n14539 & n14547;
  assign n14552 = n14550 & n14551;
  assign n14553 = n1582 & n14552;
  assign n14554 = n5385 & n14553;
  assign n14555 = n3896 & n12250;
  assign n14556 = n564 & n12256;
  assign n14557 = n3683 & n12253;
  assign n14558 = n12310 & ~n12312;
  assign n14559 = ~n12313 & ~n14558;
  assign n14560 = n566 & n14559;
  assign n14561 = ~n14556 & ~n14557;
  assign n14562 = ~n14555 & n14561;
  assign n14563 = ~n14560 & n14562;
  assign n14564 = ~n14554 & ~n14563;
  assign n14565 = ~n239 & ~n545;
  assign n14566 = ~n574 & ~n646;
  assign n14567 = n14565 & n14566;
  assign n14568 = n537 & n1082;
  assign n14569 = n1398 & n1911;
  assign n14570 = n3351 & n3379;
  assign n14571 = n4274 & n14570;
  assign n14572 = n14568 & n14569;
  assign n14573 = n14567 & n14572;
  assign n14574 = n3084 & n14571;
  assign n14575 = n14573 & n14574;
  assign n14576 = n3709 & n6422;
  assign n14577 = n14575 & n14576;
  assign n14578 = n1452 & n14577;
  assign n14579 = n1833 & n14578;
  assign n14580 = n3896 & n12253;
  assign n14581 = n564 & n12259;
  assign n14582 = n3683 & n12256;
  assign n14583 = n12306 & ~n12308;
  assign n14584 = ~n12309 & ~n14583;
  assign n14585 = n566 & n14584;
  assign n14586 = ~n14581 & ~n14582;
  assign n14587 = ~n14580 & n14586;
  assign n14588 = ~n14585 & n14587;
  assign n14589 = ~n14579 & ~n14588;
  assign n14590 = ~n177 & ~n179;
  assign n14591 = ~n385 & ~n590;
  assign n14592 = ~n674 & n14591;
  assign n14593 = n1783 & n14590;
  assign n14594 = n1869 & n2365;
  assign n14595 = n14593 & n14594;
  assign n14596 = n345 & n14592;
  assign n14597 = n2294 & n3265;
  assign n14598 = n4934 & n14597;
  assign n14599 = n14595 & n14596;
  assign n14600 = n14598 & n14599;
  assign n14601 = n3213 & n14600;
  assign n14602 = n2471 & n14601;
  assign n14603 = n14184 & n14602;
  assign n14604 = n3896 & n12256;
  assign n14605 = n564 & n12262;
  assign n14606 = n3683 & n12259;
  assign n14607 = n12302 & ~n12304;
  assign n14608 = ~n12305 & ~n14607;
  assign n14609 = n566 & n14608;
  assign n14610 = ~n14605 & ~n14606;
  assign n14611 = ~n14604 & n14610;
  assign n14612 = ~n14609 & n14611;
  assign n14613 = ~n14603 & ~n14612;
  assign n14614 = ~n216 & ~n289;
  assign n14615 = ~n447 & ~n641;
  assign n14616 = n14614 & n14615;
  assign n14617 = n194 & n1786;
  assign n14618 = n14616 & n14617;
  assign n14619 = ~n239 & ~n276;
  assign n14620 = ~n297 & ~n401;
  assign n14621 = n14619 & n14620;
  assign n14622 = n325 & n464;
  assign n14623 = n1148 & n2112;
  assign n14624 = n4931 & n14623;
  assign n14625 = n14621 & n14622;
  assign n14626 = n2294 & n3711;
  assign n14627 = n14625 & n14626;
  assign n14628 = n14618 & n14624;
  assign n14629 = n14627 & n14628;
  assign n14630 = n937 & n4417;
  assign n14631 = n14629 & n14630;
  assign n14632 = n4194 & n14631;
  assign n14633 = n3896 & n12259;
  assign n14634 = n564 & n12265;
  assign n14635 = n3683 & n12262;
  assign n14636 = n12298 & ~n12300;
  assign n14637 = ~n12301 & ~n14636;
  assign n14638 = n566 & n14637;
  assign n14639 = ~n14634 & ~n14635;
  assign n14640 = ~n14633 & n14639;
  assign n14641 = ~n14638 & n14640;
  assign n14642 = ~n14632 & ~n14641;
  assign n14643 = ~n120 & ~n387;
  assign n14644 = n3807 & n14643;
  assign n14645 = ~n222 & ~n247;
  assign n14646 = ~n511 & n14645;
  assign n14647 = ~n103 & ~n167;
  assign n14648 = ~n240 & ~n242;
  assign n14649 = ~n324 & ~n521;
  assign n14650 = ~n675 & n14649;
  assign n14651 = n14647 & n14648;
  assign n14652 = n1594 & n2271;
  assign n14653 = n4767 & n14652;
  assign n14654 = n14650 & n14651;
  assign n14655 = n2240 & n14646;
  assign n14656 = n14654 & n14655;
  assign n14657 = n4390 & n14653;
  assign n14658 = n14656 & n14657;
  assign n14659 = n6933 & n14658;
  assign n14660 = ~n466 & ~n480;
  assign n14661 = n461 & n14660;
  assign n14662 = n555 & n882;
  assign n14663 = n1112 & n2959;
  assign n14664 = n12752 & n14663;
  assign n14665 = n14661 & n14662;
  assign n14666 = n368 & n3711;
  assign n14667 = n5718 & n13452;
  assign n14668 = n14666 & n14667;
  assign n14669 = n14664 & n14665;
  assign n14670 = n348 & n14669;
  assign n14671 = n14668 & n14670;
  assign n14672 = ~n122 & ~n172;
  assign n14673 = ~n648 & n14672;
  assign n14674 = n403 & n2706;
  assign n14675 = n4264 & n12767;
  assign n14676 = n14674 & n14675;
  assign n14677 = n2111 & n14673;
  assign n14678 = n3390 & n5758;
  assign n14679 = n14644 & n14678;
  assign n14680 = n14676 & n14677;
  assign n14681 = n295 & n6838;
  assign n14682 = n14680 & n14681;
  assign n14683 = n13161 & n14679;
  assign n14684 = n14682 & n14683;
  assign n14685 = n14659 & n14684;
  assign n14686 = n14671 & n14685;
  assign n14687 = n3896 & n12262;
  assign n14688 = n564 & n12268;
  assign n14689 = n3683 & n12265;
  assign n14690 = n12294 & ~n12296;
  assign n14691 = ~n12297 & ~n14690;
  assign n14692 = n566 & n14691;
  assign n14693 = ~n14688 & ~n14689;
  assign n14694 = ~n14687 & n14693;
  assign n14695 = ~n14692 & n14694;
  assign n14696 = ~n14686 & ~n14695;
  assign n14697 = ~n225 & ~n496;
  assign n14698 = ~n543 & ~n595;
  assign n14699 = n14697 & n14698;
  assign n14700 = n237 & n922;
  assign n14701 = n1233 & n1535;
  assign n14702 = n1907 & n2008;
  assign n14703 = n3154 & n14702;
  assign n14704 = n14700 & n14701;
  assign n14705 = n3854 & n14699;
  assign n14706 = n3993 & n14705;
  assign n14707 = n14703 & n14704;
  assign n14708 = n14706 & n14707;
  assign n14709 = n2106 & n14708;
  assign n14710 = n13489 & n14709;
  assign n14711 = ~n406 & ~n675;
  assign n14712 = ~n336 & ~n554;
  assign n14713 = ~n651 & n14712;
  assign n14714 = n201 & n1156;
  assign n14715 = n1689 & n2088;
  assign n14716 = n3073 & n14711;
  assign n14717 = n14715 & n14716;
  assign n14718 = n14713 & n14714;
  assign n14719 = n14717 & n14718;
  assign n14720 = n2545 & n14719;
  assign n14721 = n3991 & n14720;
  assign n14722 = n12122 & n14721;
  assign n14723 = n14710 & n14722;
  assign n14724 = n3896 & n12265;
  assign n14725 = n564 & n12271;
  assign n14726 = n3683 & n12268;
  assign n14727 = n12290 & ~n12292;
  assign n14728 = ~n12293 & ~n14727;
  assign n14729 = n566 & n14728;
  assign n14730 = ~n14725 & ~n14726;
  assign n14731 = ~n14724 & n14730;
  assign n14732 = ~n14729 & n14731;
  assign n14733 = ~n14723 & ~n14732;
  assign n14734 = ~n92 & ~n514;
  assign n14735 = ~n679 & n14734;
  assign n14736 = n4384 & n14735;
  assign n14737 = n942 & n14736;
  assign n14738 = ~n207 & n1633;
  assign n14739 = n12627 & n14738;
  assign n14740 = ~n134 & ~n202;
  assign n14741 = ~n267 & ~n355;
  assign n14742 = ~n378 & ~n402;
  assign n14743 = ~n426 & ~n662;
  assign n14744 = n14742 & n14743;
  assign n14745 = n14740 & n14741;
  assign n14746 = n1232 & n14745;
  assign n14747 = n170 & n14744;
  assign n14748 = n3074 & n14747;
  assign n14749 = n14739 & n14746;
  assign n14750 = n14748 & n14749;
  assign n14751 = n13405 & n14737;
  assign n14752 = n14750 & n14751;
  assign n14753 = ~n585 & n2096;
  assign n14754 = ~n362 & ~n424;
  assign n14755 = ~n512 & ~n674;
  assign n14756 = n14754 & n14755;
  assign n14757 = n214 & n2493;
  assign n14758 = n2943 & n14757;
  assign n14759 = n1968 & n14756;
  assign n14760 = n14753 & n14759;
  assign n14761 = n1468 & n14758;
  assign n14762 = n5359 & n14761;
  assign n14763 = n14760 & n14762;
  assign n14764 = n2992 & n14763;
  assign n14765 = n14752 & n14764;
  assign n14766 = n2292 & n14765;
  assign n14767 = n3896 & n12268;
  assign n14768 = n564 & n12274;
  assign n14769 = n3683 & n12271;
  assign n14770 = n12286 & ~n12288;
  assign n14771 = ~n12289 & ~n14770;
  assign n14772 = n566 & n14771;
  assign n14773 = ~n14768 & ~n14769;
  assign n14774 = ~n14767 & n14773;
  assign n14775 = ~n14772 & n14774;
  assign n14776 = ~n14766 & ~n14775;
  assign n14777 = ~n113 & ~n131;
  assign n14778 = ~n545 & ~n676;
  assign n14779 = n14777 & n14778;
  assign n14780 = n268 & n325;
  assign n14781 = n1587 & n14780;
  assign n14782 = n4420 & n14779;
  assign n14783 = n14781 & n14782;
  assign n14784 = n656 & n3250;
  assign n14785 = n6898 & n14784;
  assign n14786 = n5757 & n14783;
  assign n14787 = n14785 & n14786;
  assign n14788 = n3620 & n3744;
  assign n14789 = n14787 & n14788;
  assign n14790 = n4381 & n14789;
  assign n14791 = n3896 & n12271;
  assign n14792 = n564 & n12279;
  assign n14793 = n3683 & n12274;
  assign n14794 = ~n12277 & ~n12284;
  assign n14795 = ~n12285 & ~n14794;
  assign n14796 = n566 & n14795;
  assign n14797 = ~n14792 & ~n14793;
  assign n14798 = ~n14791 & n14797;
  assign n14799 = ~n14796 & n14798;
  assign n14800 = ~n14790 & ~n14799;
  assign n14801 = ~n195 & ~n327;
  assign n14802 = ~n271 & ~n324;
  assign n14803 = ~n536 & n14802;
  assign n14804 = n2945 & n14801;
  assign n14805 = n14803 & n14804;
  assign n14806 = n1903 & n14805;
  assign n14807 = ~n300 & n967;
  assign n14808 = n1016 & n1085;
  assign n14809 = n6220 & n14808;
  assign n14810 = n669 & n14807;
  assign n14811 = n4985 & n14810;
  assign n14812 = n736 & n14809;
  assign n14813 = n3841 & n14618;
  assign n14814 = n14812 & n14813;
  assign n14815 = n14806 & n14811;
  assign n14816 = n14814 & n14815;
  assign n14817 = ~n207 & ~n662;
  assign n14818 = ~n313 & n524;
  assign n14819 = n2178 & n2424;
  assign n14820 = n2736 & n14817;
  assign n14821 = n14819 & n14820;
  assign n14822 = n14818 & n14821;
  assign n14823 = n829 & n2804;
  assign n14824 = n2829 & n2882;
  assign n14825 = n14823 & n14824;
  assign n14826 = n14822 & n14825;
  assign n14827 = n6989 & n14826;
  assign n14828 = n14816 & n14827;
  assign n14829 = n3104 & n14828;
  assign n14830 = n3896 & n12279;
  assign n14831 = n3683 & n12281;
  assign n14832 = ~n12279 & n12281;
  assign n14833 = ~n12282 & ~n14832;
  assign n14834 = n566 & ~n14833;
  assign n14835 = ~n14830 & ~n14831;
  assign n14836 = ~n14834 & n14835;
  assign n14837 = ~n14829 & ~n14836;
  assign n14838 = ~n234 & ~n591;
  assign n14839 = ~n676 & n14838;
  assign n14840 = ~n253 & ~n462;
  assign n14841 = ~n513 & ~n574;
  assign n14842 = ~n701 & n14841;
  assign n14843 = n433 & n14840;
  assign n14844 = n1689 & n1786;
  assign n14845 = n1944 & n2178;
  assign n14846 = n14844 & n14845;
  assign n14847 = n14842 & n14843;
  assign n14848 = n1629 & n14839;
  assign n14849 = n14847 & n14848;
  assign n14850 = n14846 & n14849;
  assign n14851 = ~n245 & ~n283;
  assign n14852 = ~n313 & ~n339;
  assign n14853 = ~n381 & ~n545;
  assign n14854 = ~n568 & ~n572;
  assign n14855 = ~n690 & n14854;
  assign n14856 = n14852 & n14853;
  assign n14857 = n672 & n14851;
  assign n14858 = n1121 & n1562;
  assign n14859 = n2092 & n14858;
  assign n14860 = n14856 & n14857;
  assign n14861 = n1308 & n14855;
  assign n14862 = n3611 & n4012;
  assign n14863 = n14861 & n14862;
  assign n14864 = n14859 & n14860;
  assign n14865 = n14863 & n14864;
  assign n14866 = n14162 & n14865;
  assign n14867 = n14850 & n14866;
  assign n14868 = n13427 & n14867;
  assign n14869 = n14837 & ~n14868;
  assign n14870 = ~n14837 & n14868;
  assign n14871 = ~n14869 & ~n14870;
  assign n14872 = n3896 & n12274;
  assign n14873 = n3683 & n12279;
  assign n14874 = n564 & n12281;
  assign n14875 = n12274 & ~n12282;
  assign n14876 = ~n12283 & ~n14875;
  assign n14877 = n566 & ~n14876;
  assign n14878 = ~n14873 & ~n14874;
  assign n14879 = ~n14872 & n14878;
  assign n14880 = ~n14877 & n14879;
  assign n14881 = n14871 & ~n14880;
  assign n14882 = ~n14869 & ~n14881;
  assign n14883 = n14790 & n14799;
  assign n14884 = ~n14800 & ~n14883;
  assign n14885 = ~n14882 & n14884;
  assign n14886 = ~n14800 & ~n14885;
  assign n14887 = n14766 & n14775;
  assign n14888 = ~n14776 & ~n14887;
  assign n14889 = ~n14886 & n14888;
  assign n14890 = ~n14776 & ~n14889;
  assign n14891 = n14723 & n14732;
  assign n14892 = ~n14733 & ~n14891;
  assign n14893 = ~n14890 & n14892;
  assign n14894 = ~n14733 & ~n14893;
  assign n14895 = n14686 & n14695;
  assign n14896 = ~n14696 & ~n14895;
  assign n14897 = ~n14894 & n14896;
  assign n14898 = ~n14696 & ~n14897;
  assign n14899 = n14632 & n14641;
  assign n14900 = ~n14642 & ~n14899;
  assign n14901 = ~n14898 & n14900;
  assign n14902 = ~n14642 & ~n14901;
  assign n14903 = n14603 & n14612;
  assign n14904 = ~n14613 & ~n14903;
  assign n14905 = ~n14902 & n14904;
  assign n14906 = ~n14613 & ~n14905;
  assign n14907 = n14579 & n14588;
  assign n14908 = ~n14589 & ~n14907;
  assign n14909 = ~n14906 & n14908;
  assign n14910 = ~n14589 & ~n14909;
  assign n14911 = n14554 & n14563;
  assign n14912 = ~n14564 & ~n14911;
  assign n14913 = ~n14910 & n14912;
  assign n14914 = ~n14564 & ~n14913;
  assign n14915 = ~n14534 & ~n14914;
  assign n14916 = n14534 & n14914;
  assign n14917 = ~n14915 & ~n14916;
  assign n14918 = n4472 & n12238;
  assign n14919 = n4070 & n12241;
  assign n14920 = n3943 & n12244;
  assign n14921 = n3944 & n14229;
  assign n14922 = ~n14919 & ~n14920;
  assign n14923 = ~n14918 & n14922;
  assign n14924 = ~n14921 & n14923;
  assign n14925 = pi29  & n14924;
  assign n14926 = ~pi29  & ~n14924;
  assign n14927 = ~n14925 & ~n14926;
  assign n14928 = n14917 & ~n14927;
  assign n14929 = ~n14915 & ~n14928;
  assign n14930 = ~n14522 & n14531;
  assign n14931 = ~n14532 & ~n14930;
  assign n14932 = ~n14929 & n14931;
  assign n14933 = ~n14532 & ~n14932;
  assign n14934 = ~n14510 & n14519;
  assign n14935 = ~n14520 & ~n14934;
  assign n14936 = ~n14933 & n14935;
  assign n14937 = ~n14520 & ~n14936;
  assign n14938 = ~n14224 & n14233;
  assign n14939 = ~n14234 & ~n14938;
  assign n14940 = ~n14937 & n14939;
  assign n14941 = n14937 & ~n14939;
  assign n14942 = ~n14940 & ~n14941;
  assign n14943 = n4472 & n12229;
  assign n14944 = n4070 & n12232;
  assign n14945 = n3943 & n12235;
  assign n14946 = n3944 & n13979;
  assign n14947 = ~n14944 & ~n14945;
  assign n14948 = ~n14943 & n14947;
  assign n14949 = ~n14946 & n14948;
  assign n14950 = pi29  & n14949;
  assign n14951 = ~pi29  & ~n14949;
  assign n14952 = ~n14950 & ~n14951;
  assign n14953 = n14942 & ~n14952;
  assign n14954 = ~n14940 & ~n14953;
  assign n14955 = ~n14240 & n14250;
  assign n14956 = ~n14251 & ~n14955;
  assign n14957 = ~n14954 & n14956;
  assign n14958 = n14954 & ~n14956;
  assign n14959 = ~n14957 & ~n14958;
  assign n14960 = n4721 & n12217;
  assign n14961 = n4691 & n12220;
  assign n14962 = n4515 & n12223;
  assign n14963 = n4516 & n13374;
  assign n14964 = ~n14961 & ~n14962;
  assign n14965 = ~n14960 & n14964;
  assign n14966 = ~n14963 & n14965;
  assign n14967 = pi26  & n14966;
  assign n14968 = ~pi26  & ~n14966;
  assign n14969 = ~n14967 & ~n14968;
  assign n14970 = n14959 & ~n14969;
  assign n14971 = ~n14957 & ~n14970;
  assign n14972 = n14401 & ~n14403;
  assign n14973 = ~n14404 & ~n14972;
  assign n14974 = ~n14971 & n14973;
  assign n14975 = n14971 & ~n14973;
  assign n14976 = ~n14974 & ~n14975;
  assign n14977 = n5267 & n12205;
  assign n14978 = n5185 & n12208;
  assign n14979 = n5121 & n12211;
  assign n14980 = n78 & n13031;
  assign n14981 = ~n14978 & ~n14979;
  assign n14982 = ~n14977 & n14981;
  assign n14983 = ~n14980 & n14982;
  assign n14984 = pi23  & n14983;
  assign n14985 = ~pi23  & ~n14983;
  assign n14986 = ~n14984 & ~n14985;
  assign n14987 = n14976 & ~n14986;
  assign n14988 = ~n14974 & ~n14987;
  assign n14989 = ~n14497 & n14507;
  assign n14990 = ~n14508 & ~n14989;
  assign n14991 = ~n14988 & n14990;
  assign n14992 = ~n14508 & ~n14991;
  assign n14993 = ~n14414 & n14424;
  assign n14994 = ~n14425 & ~n14993;
  assign n14995 = ~n14992 & n14994;
  assign n14996 = n14992 & ~n14994;
  assign n14997 = ~n14995 & ~n14996;
  assign n14998 = n5982 & n12190;
  assign n14999 = n5901 & n12193;
  assign n15000 = n5312 & n12196;
  assign n15001 = n5306 & n12530;
  assign n15002 = ~n14999 & ~n15000;
  assign n15003 = ~n14998 & n15002;
  assign n15004 = ~n15001 & n15003;
  assign n15005 = pi20  & n15004;
  assign n15006 = ~pi20  & ~n15004;
  assign n15007 = ~n15005 & ~n15006;
  assign n15008 = n14997 & ~n15007;
  assign n15009 = ~n14995 & ~n15008;
  assign n15010 = ~n14431 & n14441;
  assign n15011 = ~n14442 & ~n15010;
  assign n15012 = ~n15009 & n15011;
  assign n15013 = n15009 & ~n15011;
  assign n15014 = ~n15012 & ~n15013;
  assign n15015 = n6608 & n12178;
  assign n15016 = n6356 & n12181;
  assign n15017 = n6140 & n12184;
  assign n15018 = n6134 & n12880;
  assign n15019 = ~n15016 & ~n15017;
  assign n15020 = ~n15015 & n15019;
  assign n15021 = ~n15018 & n15020;
  assign n15022 = pi17  & n15021;
  assign n15023 = ~pi17  & ~n15021;
  assign n15024 = ~n15022 & ~n15023;
  assign n15025 = n15014 & ~n15024;
  assign n15026 = ~n15012 & ~n15025;
  assign n15027 = ~n14484 & n14494;
  assign n15028 = ~n14495 & ~n15027;
  assign n15029 = ~n15026 & n15028;
  assign n15030 = ~n14495 & ~n15029;
  assign n15031 = ~n14452 & n14462;
  assign n15032 = ~n14463 & ~n15031;
  assign n15033 = ~n15030 & n15032;
  assign n15034 = n15030 & ~n15032;
  assign n15035 = ~n15033 & ~n15034;
  assign n15036 = n6647 & n13007;
  assign n15037 = n6653 & n12172;
  assign n15038 = ~n7380 & n12165;
  assign n15039 = ~n12163 & ~n12787;
  assign n15040 = ~n15038 & n15039;
  assign n15041 = ~n15037 & ~n15040;
  assign n15042 = ~n15036 & n15041;
  assign n15043 = pi14  & n15042;
  assign n15044 = ~pi14  & ~n15042;
  assign n15045 = ~n15043 & ~n15044;
  assign n15046 = n15035 & ~n15045;
  assign n15047 = ~n15033 & ~n15046;
  assign n15048 = ~n14475 & ~n14477;
  assign n15049 = ~n14478 & ~n15048;
  assign n15050 = ~n15047 & n15049;
  assign n15051 = n15047 & ~n15049;
  assign n15052 = ~n15050 & ~n15051;
  assign n15053 = n14988 & ~n14990;
  assign n15054 = ~n14991 & ~n15053;
  assign n15055 = n5982 & n12193;
  assign n15056 = n5901 & n12196;
  assign n15057 = n5312 & n12199;
  assign n15058 = n5306 & n12594;
  assign n15059 = ~n15056 & ~n15057;
  assign n15060 = ~n15055 & n15059;
  assign n15061 = ~n15058 & n15060;
  assign n15062 = pi20  & n15061;
  assign n15063 = ~pi20  & ~n15061;
  assign n15064 = ~n15062 & ~n15063;
  assign n15065 = n15054 & ~n15064;
  assign n15066 = n4721 & n12220;
  assign n15067 = n4691 & n12223;
  assign n15068 = n4515 & n12226;
  assign n15069 = n4516 & n13392;
  assign n15070 = ~n15067 & ~n15068;
  assign n15071 = ~n15066 & n15070;
  assign n15072 = ~n15069 & n15071;
  assign n15073 = pi26  & n15072;
  assign n15074 = ~pi26  & ~n15072;
  assign n15075 = ~n15073 & ~n15074;
  assign n15076 = ~n14942 & n14952;
  assign n15077 = ~n14953 & ~n15076;
  assign n15078 = ~n15075 & n15077;
  assign n15079 = n14933 & ~n14935;
  assign n15080 = ~n14936 & ~n15079;
  assign n15081 = n4472 & n12232;
  assign n15082 = n4070 & n12235;
  assign n15083 = n3943 & n12238;
  assign n15084 = n3944 & n14116;
  assign n15085 = ~n15082 & ~n15083;
  assign n15086 = ~n15081 & n15085;
  assign n15087 = ~n15084 & n15086;
  assign n15088 = pi29  & n15087;
  assign n15089 = ~pi29  & ~n15087;
  assign n15090 = ~n15088 & ~n15089;
  assign n15091 = n15080 & ~n15090;
  assign n15092 = n4721 & n12223;
  assign n15093 = n4691 & n12226;
  assign n15094 = n4515 & n12229;
  assign n15095 = n4516 & n13745;
  assign n15096 = ~n15093 & ~n15094;
  assign n15097 = ~n15092 & n15096;
  assign n15098 = ~n15095 & n15097;
  assign n15099 = pi26  & n15098;
  assign n15100 = ~pi26  & ~n15098;
  assign n15101 = ~n15099 & ~n15100;
  assign n15102 = ~n15080 & n15090;
  assign n15103 = ~n15091 & ~n15102;
  assign n15104 = ~n15101 & n15103;
  assign n15105 = ~n15091 & ~n15104;
  assign n15106 = n15075 & ~n15077;
  assign n15107 = ~n15078 & ~n15106;
  assign n15108 = ~n15105 & n15107;
  assign n15109 = ~n15078 & ~n15108;
  assign n15110 = ~n14959 & n14969;
  assign n15111 = ~n14970 & ~n15110;
  assign n15112 = ~n15109 & n15111;
  assign n15113 = n15109 & ~n15111;
  assign n15114 = ~n15112 & ~n15113;
  assign n15115 = n5267 & n12208;
  assign n15116 = n5185 & n12211;
  assign n15117 = n5121 & n12214;
  assign n15118 = n78 & n12804;
  assign n15119 = ~n15116 & ~n15117;
  assign n15120 = ~n15115 & n15119;
  assign n15121 = ~n15118 & n15120;
  assign n15122 = pi23  & n15121;
  assign n15123 = ~pi23  & ~n15121;
  assign n15124 = ~n15122 & ~n15123;
  assign n15125 = n15114 & ~n15124;
  assign n15126 = ~n15112 & ~n15125;
  assign n15127 = ~n14976 & n14986;
  assign n15128 = ~n14987 & ~n15127;
  assign n15129 = ~n15126 & n15128;
  assign n15130 = n15126 & ~n15128;
  assign n15131 = ~n15129 & ~n15130;
  assign n15132 = n5982 & n12196;
  assign n15133 = n5901 & n12199;
  assign n15134 = n5312 & n12202;
  assign n15135 = n5306 & n12578;
  assign n15136 = ~n15133 & ~n15134;
  assign n15137 = ~n15132 & n15136;
  assign n15138 = ~n15135 & n15137;
  assign n15139 = pi20  & n15138;
  assign n15140 = ~pi20  & ~n15138;
  assign n15141 = ~n15139 & ~n15140;
  assign n15142 = n15131 & ~n15141;
  assign n15143 = ~n15129 & ~n15142;
  assign n15144 = ~n15054 & n15064;
  assign n15145 = ~n15065 & ~n15144;
  assign n15146 = ~n15143 & n15145;
  assign n15147 = ~n15065 & ~n15146;
  assign n15148 = ~n14997 & n15007;
  assign n15149 = ~n15008 & ~n15148;
  assign n15150 = ~n15147 & n15149;
  assign n15151 = n15147 & ~n15149;
  assign n15152 = ~n15150 & ~n15151;
  assign n15153 = n6608 & n12181;
  assign n15154 = n6356 & n12184;
  assign n15155 = n6140 & n12187;
  assign n15156 = n6134 & n12608;
  assign n15157 = ~n15154 & ~n15155;
  assign n15158 = ~n15153 & n15157;
  assign n15159 = ~n15156 & n15158;
  assign n15160 = pi17  & n15159;
  assign n15161 = ~pi17  & ~n15159;
  assign n15162 = ~n15160 & ~n15161;
  assign n15163 = n15152 & ~n15162;
  assign n15164 = ~n15150 & ~n15163;
  assign n15165 = ~n15014 & n15024;
  assign n15166 = ~n15025 & ~n15165;
  assign n15167 = ~n15164 & n15166;
  assign n15168 = n15164 & ~n15166;
  assign n15169 = ~n15167 & ~n15168;
  assign n15170 = n7380 & n12172;
  assign n15171 = n7243 & n12168;
  assign n15172 = n6653 & n12175;
  assign n15173 = n6647 & n12939;
  assign n15174 = ~n15171 & ~n15172;
  assign n15175 = ~n15170 & n15174;
  assign n15176 = ~n15173 & n15175;
  assign n15177 = pi14  & n15176;
  assign n15178 = ~pi14  & ~n15176;
  assign n15179 = ~n15177 & ~n15178;
  assign n15180 = n15169 & ~n15179;
  assign n15181 = ~n15167 & ~n15180;
  assign n15182 = n7380 & n12166;
  assign n15183 = n7243 & n12172;
  assign n15184 = n6653 & n12168;
  assign n15185 = n6647 & n13106;
  assign n15186 = ~n15182 & ~n15184;
  assign n15187 = ~n15183 & n15186;
  assign n15188 = ~n15185 & n15187;
  assign n15189 = pi14  & n15188;
  assign n15190 = ~pi14  & ~n15188;
  assign n15191 = ~n15189 & ~n15190;
  assign n15192 = ~n15181 & ~n15191;
  assign n15193 = n15026 & ~n15028;
  assign n15194 = ~n15029 & ~n15193;
  assign n15195 = n15181 & n15191;
  assign n15196 = ~n15192 & ~n15195;
  assign n15197 = n15194 & n15196;
  assign n15198 = ~n15192 & ~n15197;
  assign n15199 = ~n15035 & n15045;
  assign n15200 = ~n15046 & ~n15199;
  assign n15201 = ~n15198 & n15200;
  assign n15202 = n15143 & ~n15145;
  assign n15203 = ~n15146 & ~n15202;
  assign n15204 = n6608 & n12184;
  assign n15205 = n6356 & n12187;
  assign n15206 = n6140 & n12190;
  assign n15207 = n6134 & n12845;
  assign n15208 = ~n15205 & ~n15206;
  assign n15209 = ~n15204 & n15208;
  assign n15210 = ~n15207 & n15209;
  assign n15211 = pi17  & n15210;
  assign n15212 = ~pi17  & ~n15210;
  assign n15213 = ~n15211 & ~n15212;
  assign n15214 = n15203 & ~n15213;
  assign n15215 = n15105 & ~n15107;
  assign n15216 = ~n15108 & ~n15215;
  assign n15217 = n5267 & n12211;
  assign n15218 = n5185 & n12214;
  assign n15219 = n5121 & n12217;
  assign n15220 = n78 & n13203;
  assign n15221 = ~n15218 & ~n15219;
  assign n15222 = ~n15217 & n15221;
  assign n15223 = ~n15220 & n15222;
  assign n15224 = pi23  & n15223;
  assign n15225 = ~pi23  & ~n15223;
  assign n15226 = ~n15224 & ~n15225;
  assign n15227 = n15216 & ~n15226;
  assign n15228 = n14929 & ~n14931;
  assign n15229 = ~n14932 & ~n15228;
  assign n15230 = n4472 & n12235;
  assign n15231 = n4070 & n12238;
  assign n15232 = n3943 & n12241;
  assign n15233 = n3944 & n13959;
  assign n15234 = ~n15231 & ~n15232;
  assign n15235 = ~n15230 & n15234;
  assign n15236 = ~n15233 & n15235;
  assign n15237 = pi29  & n15236;
  assign n15238 = ~pi29  & ~n15236;
  assign n15239 = ~n15237 & ~n15238;
  assign n15240 = n15229 & ~n15239;
  assign n15241 = n4721 & n12226;
  assign n15242 = n4515 & n12232;
  assign n15243 = n4691 & n12229;
  assign n15244 = n4516 & n13530;
  assign n15245 = ~n15242 & ~n15243;
  assign n15246 = ~n15241 & n15245;
  assign n15247 = ~n15244 & n15246;
  assign n15248 = pi26  & n15247;
  assign n15249 = ~pi26  & ~n15247;
  assign n15250 = ~n15248 & ~n15249;
  assign n15251 = ~n15229 & n15239;
  assign n15252 = ~n15240 & ~n15251;
  assign n15253 = ~n15250 & n15252;
  assign n15254 = ~n15240 & ~n15253;
  assign n15255 = n15101 & ~n15103;
  assign n15256 = ~n15104 & ~n15255;
  assign n15257 = ~n15254 & n15256;
  assign n15258 = n15254 & ~n15256;
  assign n15259 = ~n15257 & ~n15258;
  assign n15260 = n5267 & n12214;
  assign n15261 = n5185 & n12217;
  assign n15262 = n5121 & n12220;
  assign n15263 = n78 & n13187;
  assign n15264 = ~n15261 & ~n15262;
  assign n15265 = ~n15260 & n15264;
  assign n15266 = ~n15263 & n15265;
  assign n15267 = pi23  & n15266;
  assign n15268 = ~pi23  & ~n15266;
  assign n15269 = ~n15267 & ~n15268;
  assign n15270 = n15259 & ~n15269;
  assign n15271 = ~n15257 & ~n15270;
  assign n15272 = ~n15216 & n15226;
  assign n15273 = ~n15227 & ~n15272;
  assign n15274 = ~n15271 & n15273;
  assign n15275 = ~n15227 & ~n15274;
  assign n15276 = ~n15114 & n15124;
  assign n15277 = ~n15125 & ~n15276;
  assign n15278 = ~n15275 & n15277;
  assign n15279 = n15275 & ~n15277;
  assign n15280 = ~n15278 & ~n15279;
  assign n15281 = n5982 & n12199;
  assign n15282 = n5901 & n12202;
  assign n15283 = n5312 & n12205;
  assign n15284 = n5306 & n12683;
  assign n15285 = ~n15282 & ~n15283;
  assign n15286 = ~n15281 & n15285;
  assign n15287 = ~n15284 & n15286;
  assign n15288 = pi20  & n15287;
  assign n15289 = ~pi20  & ~n15287;
  assign n15290 = ~n15288 & ~n15289;
  assign n15291 = n15280 & ~n15290;
  assign n15292 = ~n15278 & ~n15291;
  assign n15293 = ~n15131 & n15141;
  assign n15294 = ~n15142 & ~n15293;
  assign n15295 = ~n15292 & n15294;
  assign n15296 = n15292 & ~n15294;
  assign n15297 = ~n15295 & ~n15296;
  assign n15298 = n6608 & n12187;
  assign n15299 = n6356 & n12190;
  assign n15300 = n6140 & n12193;
  assign n15301 = n6134 & n12921;
  assign n15302 = ~n15299 & ~n15300;
  assign n15303 = ~n15298 & n15302;
  assign n15304 = ~n15301 & n15303;
  assign n15305 = pi17  & n15304;
  assign n15306 = ~pi17  & ~n15304;
  assign n15307 = ~n15305 & ~n15306;
  assign n15308 = n15297 & ~n15307;
  assign n15309 = ~n15295 & ~n15308;
  assign n15310 = ~n15203 & n15213;
  assign n15311 = ~n15214 & ~n15310;
  assign n15312 = ~n15309 & n15311;
  assign n15313 = ~n15214 & ~n15312;
  assign n15314 = ~n15152 & n15162;
  assign n15315 = ~n15163 & ~n15314;
  assign n15316 = ~n15313 & n15315;
  assign n15317 = n15313 & ~n15315;
  assign n15318 = ~n15316 & ~n15317;
  assign n15319 = n7380 & n12168;
  assign n15320 = n7243 & n12175;
  assign n15321 = n6653 & n12178;
  assign n15322 = n6647 & n12862;
  assign n15323 = ~n15320 & ~n15321;
  assign n15324 = ~n15319 & n15323;
  assign n15325 = ~n15322 & n15324;
  assign n15326 = pi14  & n15325;
  assign n15327 = ~pi14  & ~n15325;
  assign n15328 = ~n15326 & ~n15327;
  assign n15329 = n15318 & ~n15328;
  assign n15330 = ~n15316 & ~n15329;
  assign n15331 = n7548 & ~n12424;
  assign n15332 = n7553 & ~n12165;
  assign n15333 = n13357 & ~n15332;
  assign n15334 = ~n12163 & ~n15333;
  assign n15335 = ~n15331 & ~n15334;
  assign n15336 = pi11  & n15335;
  assign n15337 = ~pi11  & ~n15335;
  assign n15338 = ~n15336 & ~n15337;
  assign n15339 = ~n15330 & ~n15338;
  assign n15340 = n15330 & n15338;
  assign n15341 = ~n15339 & ~n15340;
  assign n15342 = ~n15169 & n15179;
  assign n15343 = ~n15180 & ~n15342;
  assign n15344 = n15341 & n15343;
  assign n15345 = ~n15339 & ~n15344;
  assign n15346 = ~n15194 & ~n15196;
  assign n15347 = ~n15197 & ~n15346;
  assign n15348 = ~n15345 & n15347;
  assign n15349 = n15309 & ~n15311;
  assign n15350 = ~n15312 & ~n15349;
  assign n15351 = n7380 & n12175;
  assign n15352 = n7243 & n12178;
  assign n15353 = n6653 & n12181;
  assign n15354 = n6647 & n12961;
  assign n15355 = ~n15352 & ~n15353;
  assign n15356 = ~n15351 & n15355;
  assign n15357 = ~n15354 & n15356;
  assign n15358 = pi14  & n15357;
  assign n15359 = ~pi14  & ~n15357;
  assign n15360 = ~n15358 & ~n15359;
  assign n15361 = n15350 & ~n15360;
  assign n15362 = n15271 & ~n15273;
  assign n15363 = ~n15274 & ~n15362;
  assign n15364 = n5982 & n12202;
  assign n15365 = n5901 & n12205;
  assign n15366 = n5312 & n12208;
  assign n15367 = n5306 & n12701;
  assign n15368 = ~n15365 & ~n15366;
  assign n15369 = ~n15364 & n15368;
  assign n15370 = ~n15367 & n15369;
  assign n15371 = pi20  & n15370;
  assign n15372 = ~pi20  & ~n15370;
  assign n15373 = ~n15371 & ~n15372;
  assign n15374 = n15363 & ~n15373;
  assign n15375 = n15250 & ~n15252;
  assign n15376 = ~n15253 & ~n15375;
  assign n15377 = n4472 & n12241;
  assign n15378 = n4070 & n12244;
  assign n15379 = n3943 & n12247;
  assign n15380 = n3944 & n14515;
  assign n15381 = ~n15378 & ~n15379;
  assign n15382 = ~n15377 & n15381;
  assign n15383 = ~n15380 & n15382;
  assign n15384 = pi29  & n15383;
  assign n15385 = ~pi29  & ~n15383;
  assign n15386 = ~n15384 & ~n15385;
  assign n15387 = n14910 & ~n14912;
  assign n15388 = ~n14913 & ~n15387;
  assign n15389 = ~n15386 & n15388;
  assign n15390 = n4472 & n12244;
  assign n15391 = n4070 & n12247;
  assign n15392 = n3943 & n12250;
  assign n15393 = n3944 & n14527;
  assign n15394 = ~n15391 & ~n15392;
  assign n15395 = ~n15390 & n15394;
  assign n15396 = ~n15393 & n15395;
  assign n15397 = pi29  & n15396;
  assign n15398 = ~pi29  & ~n15396;
  assign n15399 = ~n15397 & ~n15398;
  assign n15400 = n14906 & ~n14908;
  assign n15401 = ~n14909 & ~n15400;
  assign n15402 = ~n15399 & n15401;
  assign n15403 = n4472 & n12247;
  assign n15404 = n4070 & n12250;
  assign n15405 = n3943 & n12253;
  assign n15406 = n3944 & n14207;
  assign n15407 = ~n15404 & ~n15405;
  assign n15408 = ~n15403 & n15407;
  assign n15409 = ~n15406 & n15408;
  assign n15410 = pi29  & n15409;
  assign n15411 = ~pi29  & ~n15409;
  assign n15412 = ~n15410 & ~n15411;
  assign n15413 = n14902 & ~n14904;
  assign n15414 = ~n14905 & ~n15413;
  assign n15415 = ~n15412 & n15414;
  assign n15416 = n4472 & n12250;
  assign n15417 = n4070 & n12253;
  assign n15418 = n3943 & n12256;
  assign n15419 = n3944 & n14559;
  assign n15420 = ~n15417 & ~n15418;
  assign n15421 = ~n15416 & n15420;
  assign n15422 = ~n15419 & n15421;
  assign n15423 = pi29  & n15422;
  assign n15424 = ~pi29  & ~n15422;
  assign n15425 = ~n15423 & ~n15424;
  assign n15426 = n14898 & ~n14900;
  assign n15427 = ~n14901 & ~n15426;
  assign n15428 = ~n15425 & n15427;
  assign n15429 = n4472 & n12253;
  assign n15430 = n4070 & n12256;
  assign n15431 = n3943 & n12259;
  assign n15432 = n3944 & n14584;
  assign n15433 = ~n15430 & ~n15431;
  assign n15434 = ~n15429 & n15433;
  assign n15435 = ~n15432 & n15434;
  assign n15436 = pi29  & n15435;
  assign n15437 = ~pi29  & ~n15435;
  assign n15438 = ~n15436 & ~n15437;
  assign n15439 = n14894 & ~n14896;
  assign n15440 = ~n14897 & ~n15439;
  assign n15441 = ~n15438 & n15440;
  assign n15442 = n4472 & n12256;
  assign n15443 = n4070 & n12259;
  assign n15444 = n3943 & n12262;
  assign n15445 = n3944 & n14608;
  assign n15446 = ~n15443 & ~n15444;
  assign n15447 = ~n15442 & n15446;
  assign n15448 = ~n15445 & n15447;
  assign n15449 = ~pi29  & ~n15448;
  assign n15450 = pi29  & n15448;
  assign n15451 = ~n15449 & ~n15450;
  assign n15452 = n14890 & ~n14892;
  assign n15453 = ~n14893 & ~n15452;
  assign n15454 = ~n15451 & n15453;
  assign n15455 = n4472 & n12259;
  assign n15456 = n4070 & n12262;
  assign n15457 = n3943 & n12265;
  assign n15458 = n3944 & n14637;
  assign n15459 = ~n15456 & ~n15457;
  assign n15460 = ~n15455 & n15459;
  assign n15461 = ~n15458 & n15460;
  assign n15462 = ~pi29  & ~n15461;
  assign n15463 = pi29  & n15461;
  assign n15464 = ~n15462 & ~n15463;
  assign n15465 = n14886 & ~n14888;
  assign n15466 = ~n14889 & ~n15465;
  assign n15467 = ~n15464 & n15466;
  assign n15468 = n4472 & n12262;
  assign n15469 = n4070 & n12265;
  assign n15470 = n3943 & n12268;
  assign n15471 = n3944 & n14691;
  assign n15472 = ~n15469 & ~n15470;
  assign n15473 = ~n15468 & n15472;
  assign n15474 = ~n15471 & n15473;
  assign n15475 = ~pi29  & ~n15474;
  assign n15476 = pi29  & n15474;
  assign n15477 = ~n15475 & ~n15476;
  assign n15478 = n14882 & ~n14884;
  assign n15479 = ~n14885 & ~n15478;
  assign n15480 = ~n15477 & n15479;
  assign n15481 = n4472 & n12265;
  assign n15482 = n4070 & n12268;
  assign n15483 = n3943 & n12271;
  assign n15484 = n3944 & n14728;
  assign n15485 = ~n15482 & ~n15483;
  assign n15486 = ~n15481 & n15485;
  assign n15487 = ~n15484 & n15486;
  assign n15488 = ~pi29  & ~n15487;
  assign n15489 = pi29  & n15487;
  assign n15490 = ~n15488 & ~n15489;
  assign n15491 = ~n14871 & n14880;
  assign n15492 = ~n14881 & ~n15491;
  assign n15493 = ~n15490 & n15492;
  assign n15494 = n4472 & n12268;
  assign n15495 = n4070 & n12271;
  assign n15496 = n3943 & n12274;
  assign n15497 = n3944 & n14771;
  assign n15498 = ~n15495 & ~n15496;
  assign n15499 = ~n15494 & n15498;
  assign n15500 = ~n15497 & n15499;
  assign n15501 = ~pi29  & ~n15500;
  assign n15502 = pi29  & n15500;
  assign n15503 = ~n15501 & ~n15502;
  assign n15504 = n14829 & n14836;
  assign n15505 = ~n14837 & ~n15504;
  assign n15506 = ~n15503 & n15505;
  assign n15507 = ~n565 & n12281;
  assign n15508 = n3941 & n12281;
  assign n15509 = pi29  & n15508;
  assign n15510 = n4472 & n12279;
  assign n15511 = n4070 & n12281;
  assign n15512 = n3944 & ~n14833;
  assign n15513 = ~n15510 & ~n15511;
  assign n15514 = ~n15512 & n15513;
  assign n15515 = ~n15509 & n15514;
  assign n15516 = n4472 & n12274;
  assign n15517 = n4070 & n12279;
  assign n15518 = n3943 & n12281;
  assign n15519 = n3944 & ~n14876;
  assign n15520 = ~n15517 & ~n15518;
  assign n15521 = ~n15516 & n15520;
  assign n15522 = ~n15519 & n15521;
  assign n15523 = pi29  & n15515;
  assign n15524 = n15522 & n15523;
  assign n15525 = n15507 & n15524;
  assign n15526 = n4472 & n12271;
  assign n15527 = n4070 & n12274;
  assign n15528 = n3943 & n12279;
  assign n15529 = n3944 & n14795;
  assign n15530 = ~n15527 & ~n15528;
  assign n15531 = ~n15526 & n15530;
  assign n15532 = ~n15529 & n15531;
  assign n15533 = ~pi29  & ~n15532;
  assign n15534 = pi29  & n15532;
  assign n15535 = ~n15533 & ~n15534;
  assign n15536 = ~n15507 & ~n15524;
  assign n15537 = ~n15525 & ~n15536;
  assign n15538 = ~n15535 & n15537;
  assign n15539 = ~n15525 & ~n15538;
  assign n15540 = n15503 & ~n15505;
  assign n15541 = ~n15506 & ~n15540;
  assign n15542 = ~n15539 & n15541;
  assign n15543 = ~n15506 & ~n15542;
  assign n15544 = n15490 & ~n15492;
  assign n15545 = ~n15493 & ~n15544;
  assign n15546 = ~n15543 & n15545;
  assign n15547 = ~n15493 & ~n15546;
  assign n15548 = n15477 & ~n15479;
  assign n15549 = ~n15480 & ~n15548;
  assign n15550 = ~n15547 & n15549;
  assign n15551 = ~n15480 & ~n15550;
  assign n15552 = n15464 & ~n15466;
  assign n15553 = ~n15467 & ~n15552;
  assign n15554 = ~n15551 & n15553;
  assign n15555 = ~n15467 & ~n15554;
  assign n15556 = n15451 & ~n15453;
  assign n15557 = ~n15454 & ~n15556;
  assign n15558 = ~n15555 & n15557;
  assign n15559 = ~n15454 & ~n15558;
  assign n15560 = n15438 & ~n15440;
  assign n15561 = ~n15441 & ~n15560;
  assign n15562 = ~n15559 & n15561;
  assign n15563 = ~n15441 & ~n15562;
  assign n15564 = n15425 & ~n15427;
  assign n15565 = ~n15428 & ~n15564;
  assign n15566 = ~n15563 & n15565;
  assign n15567 = ~n15428 & ~n15566;
  assign n15568 = n15412 & ~n15414;
  assign n15569 = ~n15415 & ~n15568;
  assign n15570 = ~n15567 & n15569;
  assign n15571 = ~n15415 & ~n15570;
  assign n15572 = n15399 & ~n15401;
  assign n15573 = ~n15402 & ~n15572;
  assign n15574 = ~n15571 & n15573;
  assign n15575 = ~n15402 & ~n15574;
  assign n15576 = n15386 & ~n15388;
  assign n15577 = ~n15389 & ~n15576;
  assign n15578 = ~n15575 & n15577;
  assign n15579 = ~n15389 & ~n15578;
  assign n15580 = ~n14917 & n14927;
  assign n15581 = ~n14928 & ~n15580;
  assign n15582 = n15579 & ~n15581;
  assign n15583 = ~n15579 & n15581;
  assign n15584 = ~n15582 & ~n15583;
  assign n15585 = n4721 & n12229;
  assign n15586 = n4691 & n12232;
  assign n15587 = n4515 & n12235;
  assign n15588 = n4516 & n13979;
  assign n15589 = ~n15586 & ~n15587;
  assign n15590 = ~n15585 & n15589;
  assign n15591 = ~n15588 & n15590;
  assign n15592 = pi26  & n15591;
  assign n15593 = ~pi26  & ~n15591;
  assign n15594 = ~n15592 & ~n15593;
  assign n15595 = n15584 & n15594;
  assign n15596 = ~n15582 & ~n15595;
  assign n15597 = n15376 & n15596;
  assign n15598 = ~n15376 & ~n15596;
  assign n15599 = ~n15597 & ~n15598;
  assign n15600 = n5267 & n12217;
  assign n15601 = n5185 & n12220;
  assign n15602 = n5121 & n12223;
  assign n15603 = n78 & n13374;
  assign n15604 = ~n15601 & ~n15602;
  assign n15605 = ~n15600 & n15604;
  assign n15606 = ~n15603 & n15605;
  assign n15607 = pi23  & n15606;
  assign n15608 = ~pi23  & ~n15606;
  assign n15609 = ~n15607 & ~n15608;
  assign n15610 = n15599 & ~n15609;
  assign n15611 = ~n15597 & ~n15610;
  assign n15612 = ~n15259 & n15269;
  assign n15613 = ~n15270 & ~n15612;
  assign n15614 = ~n15611 & n15613;
  assign n15615 = n15611 & ~n15613;
  assign n15616 = ~n15614 & ~n15615;
  assign n15617 = n5982 & n12205;
  assign n15618 = n5901 & n12208;
  assign n15619 = n5312 & n12211;
  assign n15620 = n5306 & n13031;
  assign n15621 = ~n15618 & ~n15619;
  assign n15622 = ~n15617 & n15621;
  assign n15623 = ~n15620 & n15622;
  assign n15624 = pi20  & n15623;
  assign n15625 = ~pi20  & ~n15623;
  assign n15626 = ~n15624 & ~n15625;
  assign n15627 = n15616 & ~n15626;
  assign n15628 = ~n15614 & ~n15627;
  assign n15629 = ~n15363 & n15373;
  assign n15630 = ~n15374 & ~n15629;
  assign n15631 = ~n15628 & n15630;
  assign n15632 = ~n15374 & ~n15631;
  assign n15633 = ~n15280 & n15290;
  assign n15634 = ~n15291 & ~n15633;
  assign n15635 = ~n15632 & n15634;
  assign n15636 = n15632 & ~n15634;
  assign n15637 = ~n15635 & ~n15636;
  assign n15638 = n6608 & n12190;
  assign n15639 = n6356 & n12193;
  assign n15640 = n6140 & n12196;
  assign n15641 = n6134 & n12530;
  assign n15642 = ~n15639 & ~n15640;
  assign n15643 = ~n15638 & n15642;
  assign n15644 = ~n15641 & n15643;
  assign n15645 = pi17  & n15644;
  assign n15646 = ~pi17  & ~n15644;
  assign n15647 = ~n15645 & ~n15646;
  assign n15648 = n15637 & ~n15647;
  assign n15649 = ~n15635 & ~n15648;
  assign n15650 = ~n15297 & n15307;
  assign n15651 = ~n15308 & ~n15650;
  assign n15652 = ~n15649 & n15651;
  assign n15653 = n15649 & ~n15651;
  assign n15654 = ~n15652 & ~n15653;
  assign n15655 = n7380 & n12178;
  assign n15656 = n7243 & n12181;
  assign n15657 = n6653 & n12184;
  assign n15658 = n6647 & n12880;
  assign n15659 = ~n15656 & ~n15657;
  assign n15660 = ~n15655 & n15659;
  assign n15661 = ~n15658 & n15660;
  assign n15662 = pi14  & n15661;
  assign n15663 = ~pi14  & ~n15661;
  assign n15664 = ~n15662 & ~n15663;
  assign n15665 = n15654 & ~n15664;
  assign n15666 = ~n15652 & ~n15665;
  assign n15667 = ~n15350 & n15360;
  assign n15668 = ~n15361 & ~n15667;
  assign n15669 = ~n15666 & n15668;
  assign n15670 = ~n15361 & ~n15669;
  assign n15671 = ~n15318 & n15328;
  assign n15672 = ~n15329 & ~n15671;
  assign n15673 = ~n15670 & n15672;
  assign n15674 = n15670 & ~n15672;
  assign n15675 = ~n15673 & ~n15674;
  assign n15676 = n7548 & n13007;
  assign n15677 = n7554 & n12172;
  assign n15678 = ~n8161 & n12165;
  assign n15679 = ~n12163 & ~n13357;
  assign n15680 = ~n15678 & n15679;
  assign n15681 = ~n15677 & ~n15680;
  assign n15682 = ~n15676 & n15681;
  assign n15683 = pi11  & n15682;
  assign n15684 = ~pi11  & ~n15682;
  assign n15685 = ~n15683 & ~n15684;
  assign n15686 = n15675 & ~n15685;
  assign n15687 = ~n15673 & ~n15686;
  assign n15688 = ~n15341 & ~n15343;
  assign n15689 = ~n15344 & ~n15688;
  assign n15690 = ~n15687 & n15689;
  assign n15691 = n15687 & ~n15689;
  assign n15692 = ~n15690 & ~n15691;
  assign n15693 = n15628 & ~n15630;
  assign n15694 = ~n15631 & ~n15693;
  assign n15695 = n6608 & n12193;
  assign n15696 = n6356 & n12196;
  assign n15697 = n6140 & n12199;
  assign n15698 = n6134 & n12594;
  assign n15699 = ~n15696 & ~n15697;
  assign n15700 = ~n15695 & n15699;
  assign n15701 = ~n15698 & n15700;
  assign n15702 = pi17  & n15701;
  assign n15703 = ~pi17  & ~n15701;
  assign n15704 = ~n15702 & ~n15703;
  assign n15705 = n15694 & ~n15704;
  assign n15706 = ~n15584 & ~n15594;
  assign n15707 = ~n15595 & ~n15706;
  assign n15708 = n15575 & ~n15577;
  assign n15709 = ~n15578 & ~n15708;
  assign n15710 = n4721 & n12232;
  assign n15711 = n4691 & n12235;
  assign n15712 = n4515 & n12238;
  assign n15713 = n4516 & n14116;
  assign n15714 = ~n15711 & ~n15712;
  assign n15715 = ~n15710 & n15714;
  assign n15716 = ~n15713 & n15715;
  assign n15717 = pi26  & n15716;
  assign n15718 = ~pi26  & ~n15716;
  assign n15719 = ~n15717 & ~n15718;
  assign n15720 = n15709 & ~n15719;
  assign n15721 = n15571 & ~n15573;
  assign n15722 = ~n15574 & ~n15721;
  assign n15723 = n4721 & n12235;
  assign n15724 = n4691 & n12238;
  assign n15725 = n4515 & n12241;
  assign n15726 = n4516 & n13959;
  assign n15727 = ~n15724 & ~n15725;
  assign n15728 = ~n15723 & n15727;
  assign n15729 = ~n15726 & n15728;
  assign n15730 = pi26  & n15729;
  assign n15731 = ~pi26  & ~n15729;
  assign n15732 = ~n15730 & ~n15731;
  assign n15733 = n15722 & ~n15732;
  assign n15734 = n15567 & ~n15569;
  assign n15735 = ~n15570 & ~n15734;
  assign n15736 = n4721 & n12238;
  assign n15737 = n4691 & n12241;
  assign n15738 = n4515 & n12244;
  assign n15739 = n4516 & n14229;
  assign n15740 = ~n15737 & ~n15738;
  assign n15741 = ~n15736 & n15740;
  assign n15742 = ~n15739 & n15741;
  assign n15743 = pi26  & n15742;
  assign n15744 = ~pi26  & ~n15742;
  assign n15745 = ~n15743 & ~n15744;
  assign n15746 = n15735 & ~n15745;
  assign n15747 = n15563 & ~n15565;
  assign n15748 = ~n15566 & ~n15747;
  assign n15749 = n4721 & n12241;
  assign n15750 = n4691 & n12244;
  assign n15751 = n4515 & n12247;
  assign n15752 = n4516 & n14515;
  assign n15753 = ~n15750 & ~n15751;
  assign n15754 = ~n15749 & n15753;
  assign n15755 = ~n15752 & n15754;
  assign n15756 = pi26  & n15755;
  assign n15757 = ~pi26  & ~n15755;
  assign n15758 = ~n15756 & ~n15757;
  assign n15759 = n15748 & ~n15758;
  assign n15760 = n15559 & ~n15561;
  assign n15761 = ~n15562 & ~n15760;
  assign n15762 = n4721 & n12244;
  assign n15763 = n4691 & n12247;
  assign n15764 = n4515 & n12250;
  assign n15765 = n4516 & n14527;
  assign n15766 = ~n15763 & ~n15764;
  assign n15767 = ~n15762 & n15766;
  assign n15768 = ~n15765 & n15767;
  assign n15769 = pi26  & n15768;
  assign n15770 = ~pi26  & ~n15768;
  assign n15771 = ~n15769 & ~n15770;
  assign n15772 = n15761 & ~n15771;
  assign n15773 = n15555 & ~n15557;
  assign n15774 = ~n15558 & ~n15773;
  assign n15775 = n4721 & n12247;
  assign n15776 = n4691 & n12250;
  assign n15777 = n4515 & n12253;
  assign n15778 = n4516 & n14207;
  assign n15779 = ~n15776 & ~n15777;
  assign n15780 = ~n15775 & n15779;
  assign n15781 = ~n15778 & n15780;
  assign n15782 = pi26  & n15781;
  assign n15783 = ~pi26  & ~n15781;
  assign n15784 = ~n15782 & ~n15783;
  assign n15785 = n15774 & ~n15784;
  assign n15786 = n15551 & ~n15553;
  assign n15787 = ~n15554 & ~n15786;
  assign n15788 = n4721 & n12250;
  assign n15789 = n4691 & n12253;
  assign n15790 = n4515 & n12256;
  assign n15791 = n4516 & n14559;
  assign n15792 = ~n15789 & ~n15790;
  assign n15793 = ~n15788 & n15792;
  assign n15794 = ~n15791 & n15793;
  assign n15795 = pi26  & n15794;
  assign n15796 = ~pi26  & ~n15794;
  assign n15797 = ~n15795 & ~n15796;
  assign n15798 = n15787 & ~n15797;
  assign n15799 = n15547 & ~n15549;
  assign n15800 = ~n15550 & ~n15799;
  assign n15801 = n4721 & n12253;
  assign n15802 = n4691 & n12256;
  assign n15803 = n4515 & n12259;
  assign n15804 = n4516 & n14584;
  assign n15805 = ~n15802 & ~n15803;
  assign n15806 = ~n15801 & n15805;
  assign n15807 = ~n15804 & n15806;
  assign n15808 = pi26  & n15807;
  assign n15809 = ~pi26  & ~n15807;
  assign n15810 = ~n15808 & ~n15809;
  assign n15811 = n15800 & ~n15810;
  assign n15812 = n15543 & ~n15545;
  assign n15813 = ~n15546 & ~n15812;
  assign n15814 = n4721 & n12256;
  assign n15815 = n4515 & n12262;
  assign n15816 = n4691 & n12259;
  assign n15817 = n4516 & n14608;
  assign n15818 = ~n15815 & ~n15816;
  assign n15819 = ~n15814 & n15818;
  assign n15820 = ~n15817 & n15819;
  assign n15821 = pi26  & n15820;
  assign n15822 = ~pi26  & ~n15820;
  assign n15823 = ~n15821 & ~n15822;
  assign n15824 = n15813 & ~n15823;
  assign n15825 = n4721 & n12259;
  assign n15826 = n4691 & n12262;
  assign n15827 = n4515 & n12265;
  assign n15828 = n4516 & n14637;
  assign n15829 = ~n15826 & ~n15827;
  assign n15830 = ~n15825 & n15829;
  assign n15831 = ~n15828 & n15830;
  assign n15832 = pi26  & n15831;
  assign n15833 = ~pi26  & ~n15831;
  assign n15834 = ~n15832 & ~n15833;
  assign n15835 = n15539 & ~n15541;
  assign n15836 = ~n15542 & ~n15835;
  assign n15837 = ~n15834 & n15836;
  assign n15838 = n4721 & n12262;
  assign n15839 = n4515 & n12268;
  assign n15840 = n4691 & n12265;
  assign n15841 = n4516 & n14691;
  assign n15842 = ~n15839 & ~n15840;
  assign n15843 = ~n15838 & n15842;
  assign n15844 = ~n15841 & n15843;
  assign n15845 = ~pi26  & ~n15844;
  assign n15846 = pi26  & n15844;
  assign n15847 = ~n15845 & ~n15846;
  assign n15848 = n15535 & ~n15537;
  assign n15849 = ~n15538 & ~n15848;
  assign n15850 = ~n15847 & n15849;
  assign n15851 = n4721 & n12265;
  assign n15852 = n4691 & n12268;
  assign n15853 = n4515 & n12271;
  assign n15854 = n4516 & n14728;
  assign n15855 = ~n15852 & ~n15853;
  assign n15856 = ~n15851 & n15855;
  assign n15857 = ~n15854 & n15856;
  assign n15858 = ~pi26  & ~n15857;
  assign n15859 = pi26  & n15857;
  assign n15860 = ~n15858 & ~n15859;
  assign n15861 = pi29  & ~n15515;
  assign n15862 = n15522 & ~n15861;
  assign n15863 = ~n15522 & n15861;
  assign n15864 = ~n15862 & ~n15863;
  assign n15865 = ~n15860 & n15864;
  assign n15866 = n4721 & n12268;
  assign n15867 = n4691 & n12271;
  assign n15868 = n4515 & n12274;
  assign n15869 = n4516 & n14771;
  assign n15870 = ~n15867 & ~n15868;
  assign n15871 = ~n15866 & n15870;
  assign n15872 = ~n15869 & n15871;
  assign n15873 = pi26  & n15872;
  assign n15874 = ~pi26  & ~n15872;
  assign n15875 = ~n15873 & ~n15874;
  assign n15876 = n15509 & ~n15514;
  assign n15877 = ~n15515 & ~n15876;
  assign n15878 = ~n15875 & n15877;
  assign n15879 = ~n4512 & n12281;
  assign n15880 = pi26  & n15879;
  assign n15881 = n4721 & n12279;
  assign n15882 = n4691 & n12281;
  assign n15883 = n4516 & ~n14833;
  assign n15884 = ~n15881 & ~n15882;
  assign n15885 = ~n15883 & n15884;
  assign n15886 = ~n15880 & n15885;
  assign n15887 = n4721 & n12274;
  assign n15888 = n4691 & n12279;
  assign n15889 = n4515 & n12281;
  assign n15890 = n4516 & ~n14876;
  assign n15891 = ~n15888 & ~n15889;
  assign n15892 = ~n15887 & n15891;
  assign n15893 = ~n15890 & n15892;
  assign n15894 = pi26  & n15886;
  assign n15895 = n15893 & n15894;
  assign n15896 = n15508 & n15895;
  assign n15897 = n4721 & n12271;
  assign n15898 = n4691 & n12274;
  assign n15899 = n4515 & n12279;
  assign n15900 = n4516 & n14795;
  assign n15901 = ~n15898 & ~n15899;
  assign n15902 = ~n15897 & n15901;
  assign n15903 = ~n15900 & n15902;
  assign n15904 = pi26  & n15903;
  assign n15905 = ~pi26  & ~n15903;
  assign n15906 = ~n15904 & ~n15905;
  assign n15907 = ~n15508 & ~n15895;
  assign n15908 = ~n15896 & ~n15907;
  assign n15909 = ~n15906 & n15908;
  assign n15910 = ~n15896 & ~n15909;
  assign n15911 = n15875 & ~n15877;
  assign n15912 = ~n15878 & ~n15911;
  assign n15913 = ~n15910 & n15912;
  assign n15914 = ~n15878 & ~n15913;
  assign n15915 = n15860 & ~n15864;
  assign n15916 = ~n15865 & ~n15915;
  assign n15917 = ~n15914 & n15916;
  assign n15918 = ~n15865 & ~n15917;
  assign n15919 = n15847 & ~n15849;
  assign n15920 = ~n15850 & ~n15919;
  assign n15921 = ~n15918 & n15920;
  assign n15922 = ~n15850 & ~n15921;
  assign n15923 = n15834 & ~n15836;
  assign n15924 = ~n15837 & ~n15923;
  assign n15925 = ~n15922 & n15924;
  assign n15926 = ~n15837 & ~n15925;
  assign n15927 = ~n15813 & n15823;
  assign n15928 = ~n15824 & ~n15927;
  assign n15929 = ~n15926 & n15928;
  assign n15930 = ~n15824 & ~n15929;
  assign n15931 = ~n15800 & n15810;
  assign n15932 = ~n15811 & ~n15931;
  assign n15933 = ~n15930 & n15932;
  assign n15934 = ~n15811 & ~n15933;
  assign n15935 = ~n15787 & n15797;
  assign n15936 = ~n15798 & ~n15935;
  assign n15937 = ~n15934 & n15936;
  assign n15938 = ~n15798 & ~n15937;
  assign n15939 = ~n15774 & n15784;
  assign n15940 = ~n15785 & ~n15939;
  assign n15941 = ~n15938 & n15940;
  assign n15942 = ~n15785 & ~n15941;
  assign n15943 = ~n15761 & n15771;
  assign n15944 = ~n15772 & ~n15943;
  assign n15945 = ~n15942 & n15944;
  assign n15946 = ~n15772 & ~n15945;
  assign n15947 = ~n15748 & n15758;
  assign n15948 = ~n15759 & ~n15947;
  assign n15949 = ~n15946 & n15948;
  assign n15950 = ~n15759 & ~n15949;
  assign n15951 = ~n15735 & n15745;
  assign n15952 = ~n15746 & ~n15951;
  assign n15953 = ~n15950 & n15952;
  assign n15954 = ~n15746 & ~n15953;
  assign n15955 = ~n15722 & n15732;
  assign n15956 = ~n15733 & ~n15955;
  assign n15957 = ~n15954 & n15956;
  assign n15958 = ~n15733 & ~n15957;
  assign n15959 = ~n15709 & n15719;
  assign n15960 = ~n15720 & ~n15959;
  assign n15961 = ~n15958 & n15960;
  assign n15962 = ~n15720 & ~n15961;
  assign n15963 = ~n15707 & ~n15962;
  assign n15964 = n15707 & n15962;
  assign n15965 = ~n15963 & ~n15964;
  assign n15966 = n5267 & n12220;
  assign n15967 = n5185 & n12223;
  assign n15968 = n5121 & n12226;
  assign n15969 = n78 & n13392;
  assign n15970 = ~n15967 & ~n15968;
  assign n15971 = ~n15966 & n15970;
  assign n15972 = ~n15969 & n15971;
  assign n15973 = pi23  & n15972;
  assign n15974 = ~pi23  & ~n15972;
  assign n15975 = ~n15973 & ~n15974;
  assign n15976 = n15965 & ~n15975;
  assign n15977 = ~n15963 & ~n15976;
  assign n15978 = ~n15599 & n15609;
  assign n15979 = ~n15610 & ~n15978;
  assign n15980 = ~n15977 & n15979;
  assign n15981 = n15977 & ~n15979;
  assign n15982 = ~n15980 & ~n15981;
  assign n15983 = n5982 & n12208;
  assign n15984 = n5901 & n12211;
  assign n15985 = n5312 & n12214;
  assign n15986 = n5306 & n12804;
  assign n15987 = ~n15984 & ~n15985;
  assign n15988 = ~n15983 & n15987;
  assign n15989 = ~n15986 & n15988;
  assign n15990 = pi20  & n15989;
  assign n15991 = ~pi20  & ~n15989;
  assign n15992 = ~n15990 & ~n15991;
  assign n15993 = n15982 & ~n15992;
  assign n15994 = ~n15980 & ~n15993;
  assign n15995 = ~n15616 & n15626;
  assign n15996 = ~n15627 & ~n15995;
  assign n15997 = ~n15994 & n15996;
  assign n15998 = n15994 & ~n15996;
  assign n15999 = ~n15997 & ~n15998;
  assign n16000 = n6608 & n12196;
  assign n16001 = n6356 & n12199;
  assign n16002 = n6140 & n12202;
  assign n16003 = n6134 & n12578;
  assign n16004 = ~n16001 & ~n16002;
  assign n16005 = ~n16000 & n16004;
  assign n16006 = ~n16003 & n16005;
  assign n16007 = pi17  & n16006;
  assign n16008 = ~pi17  & ~n16006;
  assign n16009 = ~n16007 & ~n16008;
  assign n16010 = n15999 & ~n16009;
  assign n16011 = ~n15997 & ~n16010;
  assign n16012 = ~n15694 & n15704;
  assign n16013 = ~n15705 & ~n16012;
  assign n16014 = ~n16011 & n16013;
  assign n16015 = ~n15705 & ~n16014;
  assign n16016 = ~n15637 & n15647;
  assign n16017 = ~n15648 & ~n16016;
  assign n16018 = ~n16015 & n16017;
  assign n16019 = n16015 & ~n16017;
  assign n16020 = ~n16018 & ~n16019;
  assign n16021 = n7380 & n12181;
  assign n16022 = n7243 & n12184;
  assign n16023 = n6653 & n12187;
  assign n16024 = n6647 & n12608;
  assign n16025 = ~n16022 & ~n16023;
  assign n16026 = ~n16021 & n16025;
  assign n16027 = ~n16024 & n16026;
  assign n16028 = pi14  & n16027;
  assign n16029 = ~pi14  & ~n16027;
  assign n16030 = ~n16028 & ~n16029;
  assign n16031 = n16020 & ~n16030;
  assign n16032 = ~n16018 & ~n16031;
  assign n16033 = ~n15654 & n15664;
  assign n16034 = ~n15665 & ~n16033;
  assign n16035 = ~n16032 & n16034;
  assign n16036 = n16032 & ~n16034;
  assign n16037 = ~n16035 & ~n16036;
  assign n16038 = n8161 & n12172;
  assign n16039 = n7847 & n12168;
  assign n16040 = n7554 & n12175;
  assign n16041 = n7548 & n12939;
  assign n16042 = ~n16039 & ~n16040;
  assign n16043 = ~n16038 & n16042;
  assign n16044 = ~n16041 & n16043;
  assign n16045 = pi11  & n16044;
  assign n16046 = ~pi11  & ~n16044;
  assign n16047 = ~n16045 & ~n16046;
  assign n16048 = n16037 & ~n16047;
  assign n16049 = ~n16035 & ~n16048;
  assign n16050 = n8161 & n12166;
  assign n16051 = n7847 & n12172;
  assign n16052 = n7554 & n12168;
  assign n16053 = n7548 & n13106;
  assign n16054 = ~n16050 & ~n16052;
  assign n16055 = ~n16051 & n16054;
  assign n16056 = ~n16053 & n16055;
  assign n16057 = pi11  & n16056;
  assign n16058 = ~pi11  & ~n16056;
  assign n16059 = ~n16057 & ~n16058;
  assign n16060 = ~n16049 & ~n16059;
  assign n16061 = n15666 & ~n15668;
  assign n16062 = ~n15669 & ~n16061;
  assign n16063 = n16049 & n16059;
  assign n16064 = ~n16060 & ~n16063;
  assign n16065 = n16062 & n16064;
  assign n16066 = ~n16060 & ~n16065;
  assign n16067 = ~n15675 & n15685;
  assign n16068 = ~n15686 & ~n16067;
  assign n16069 = ~n16066 & n16068;
  assign n16070 = n16011 & ~n16013;
  assign n16071 = ~n16014 & ~n16070;
  assign n16072 = n7380 & n12184;
  assign n16073 = n7243 & n12187;
  assign n16074 = n6653 & n12190;
  assign n16075 = n6647 & n12845;
  assign n16076 = ~n16073 & ~n16074;
  assign n16077 = ~n16072 & n16076;
  assign n16078 = ~n16075 & n16077;
  assign n16079 = pi14  & n16078;
  assign n16080 = ~pi14  & ~n16078;
  assign n16081 = ~n16079 & ~n16080;
  assign n16082 = n16071 & ~n16081;
  assign n16083 = n5267 & n12223;
  assign n16084 = n5185 & n12226;
  assign n16085 = n5121 & n12229;
  assign n16086 = n78 & n13745;
  assign n16087 = ~n16084 & ~n16085;
  assign n16088 = ~n16083 & n16087;
  assign n16089 = ~n16086 & n16088;
  assign n16090 = ~pi23  & ~n16089;
  assign n16091 = pi23  & n16089;
  assign n16092 = ~n16090 & ~n16091;
  assign n16093 = n15958 & ~n15960;
  assign n16094 = ~n15961 & ~n16093;
  assign n16095 = ~n16092 & n16094;
  assign n16096 = n5267 & n12226;
  assign n16097 = n5185 & n12229;
  assign n16098 = n5121 & n12232;
  assign n16099 = n78 & n13530;
  assign n16100 = ~n16097 & ~n16098;
  assign n16101 = ~n16096 & n16100;
  assign n16102 = ~n16099 & n16101;
  assign n16103 = ~pi23  & ~n16102;
  assign n16104 = pi23  & n16102;
  assign n16105 = ~n16103 & ~n16104;
  assign n16106 = n15954 & ~n15956;
  assign n16107 = ~n15957 & ~n16106;
  assign n16108 = ~n16105 & n16107;
  assign n16109 = n5267 & n12229;
  assign n16110 = n5185 & n12232;
  assign n16111 = n5121 & n12235;
  assign n16112 = n78 & n13979;
  assign n16113 = ~n16110 & ~n16111;
  assign n16114 = ~n16109 & n16113;
  assign n16115 = ~n16112 & n16114;
  assign n16116 = ~pi23  & ~n16115;
  assign n16117 = pi23  & n16115;
  assign n16118 = ~n16116 & ~n16117;
  assign n16119 = n15950 & ~n15952;
  assign n16120 = ~n15953 & ~n16119;
  assign n16121 = ~n16118 & n16120;
  assign n16122 = n5267 & n12232;
  assign n16123 = n5185 & n12235;
  assign n16124 = n5121 & n12238;
  assign n16125 = n78 & n14116;
  assign n16126 = ~n16123 & ~n16124;
  assign n16127 = ~n16122 & n16126;
  assign n16128 = ~n16125 & n16127;
  assign n16129 = ~pi23  & ~n16128;
  assign n16130 = pi23  & n16128;
  assign n16131 = ~n16129 & ~n16130;
  assign n16132 = n15946 & ~n15948;
  assign n16133 = ~n15949 & ~n16132;
  assign n16134 = ~n16131 & n16133;
  assign n16135 = n5267 & n12235;
  assign n16136 = n5185 & n12238;
  assign n16137 = n5121 & n12241;
  assign n16138 = n78 & n13959;
  assign n16139 = ~n16136 & ~n16137;
  assign n16140 = ~n16135 & n16139;
  assign n16141 = ~n16138 & n16140;
  assign n16142 = ~pi23  & ~n16141;
  assign n16143 = pi23  & n16141;
  assign n16144 = ~n16142 & ~n16143;
  assign n16145 = n15942 & ~n15944;
  assign n16146 = ~n15945 & ~n16145;
  assign n16147 = ~n16144 & n16146;
  assign n16148 = n5267 & n12238;
  assign n16149 = n5185 & n12241;
  assign n16150 = n5121 & n12244;
  assign n16151 = n78 & n14229;
  assign n16152 = ~n16149 & ~n16150;
  assign n16153 = ~n16148 & n16152;
  assign n16154 = ~n16151 & n16153;
  assign n16155 = ~pi23  & ~n16154;
  assign n16156 = pi23  & n16154;
  assign n16157 = ~n16155 & ~n16156;
  assign n16158 = n15938 & ~n15940;
  assign n16159 = ~n15941 & ~n16158;
  assign n16160 = ~n16157 & n16159;
  assign n16161 = n5267 & n12241;
  assign n16162 = n5185 & n12244;
  assign n16163 = n5121 & n12247;
  assign n16164 = n78 & n14515;
  assign n16165 = ~n16162 & ~n16163;
  assign n16166 = ~n16161 & n16165;
  assign n16167 = ~n16164 & n16166;
  assign n16168 = ~pi23  & ~n16167;
  assign n16169 = pi23  & n16167;
  assign n16170 = ~n16168 & ~n16169;
  assign n16171 = n15934 & ~n15936;
  assign n16172 = ~n15937 & ~n16171;
  assign n16173 = ~n16170 & n16172;
  assign n16174 = n5267 & n12244;
  assign n16175 = n5185 & n12247;
  assign n16176 = n5121 & n12250;
  assign n16177 = n78 & n14527;
  assign n16178 = ~n16175 & ~n16176;
  assign n16179 = ~n16174 & n16178;
  assign n16180 = ~n16177 & n16179;
  assign n16181 = ~pi23  & ~n16180;
  assign n16182 = pi23  & n16180;
  assign n16183 = ~n16181 & ~n16182;
  assign n16184 = n15930 & ~n15932;
  assign n16185 = ~n15933 & ~n16184;
  assign n16186 = ~n16183 & n16185;
  assign n16187 = n5267 & n12247;
  assign n16188 = n5185 & n12250;
  assign n16189 = n5121 & n12253;
  assign n16190 = n78 & n14207;
  assign n16191 = ~n16188 & ~n16189;
  assign n16192 = ~n16187 & n16191;
  assign n16193 = ~n16190 & n16192;
  assign n16194 = ~pi23  & ~n16193;
  assign n16195 = pi23  & n16193;
  assign n16196 = ~n16194 & ~n16195;
  assign n16197 = n15926 & ~n15928;
  assign n16198 = ~n15929 & ~n16197;
  assign n16199 = ~n16196 & n16198;
  assign n16200 = n5267 & n12250;
  assign n16201 = n5185 & n12253;
  assign n16202 = n5121 & n12256;
  assign n16203 = n78 & n14559;
  assign n16204 = ~n16201 & ~n16202;
  assign n16205 = ~n16200 & n16204;
  assign n16206 = ~n16203 & n16205;
  assign n16207 = ~pi23  & ~n16206;
  assign n16208 = pi23  & n16206;
  assign n16209 = ~n16207 & ~n16208;
  assign n16210 = n15922 & ~n15924;
  assign n16211 = ~n15925 & ~n16210;
  assign n16212 = ~n16209 & n16211;
  assign n16213 = n15918 & ~n15920;
  assign n16214 = ~n15921 & ~n16213;
  assign n16215 = n5267 & n12253;
  assign n16216 = n5185 & n12256;
  assign n16217 = n5121 & n12259;
  assign n16218 = n78 & n14584;
  assign n16219 = ~n16216 & ~n16217;
  assign n16220 = ~n16215 & n16219;
  assign n16221 = ~n16218 & n16220;
  assign n16222 = pi23  & n16221;
  assign n16223 = ~pi23  & ~n16221;
  assign n16224 = ~n16222 & ~n16223;
  assign n16225 = n16214 & ~n16224;
  assign n16226 = n15914 & ~n15916;
  assign n16227 = ~n15917 & ~n16226;
  assign n16228 = n5267 & n12256;
  assign n16229 = n5185 & n12259;
  assign n16230 = n5121 & n12262;
  assign n16231 = n78 & n14608;
  assign n16232 = ~n16229 & ~n16230;
  assign n16233 = ~n16228 & n16232;
  assign n16234 = ~n16231 & n16233;
  assign n16235 = pi23  & n16234;
  assign n16236 = ~pi23  & ~n16234;
  assign n16237 = ~n16235 & ~n16236;
  assign n16238 = n16227 & ~n16237;
  assign n16239 = n5267 & n12259;
  assign n16240 = n5185 & n12262;
  assign n16241 = n5121 & n12265;
  assign n16242 = n78 & n14637;
  assign n16243 = ~n16240 & ~n16241;
  assign n16244 = ~n16239 & n16243;
  assign n16245 = ~n16242 & n16244;
  assign n16246 = ~pi23  & ~n16245;
  assign n16247 = pi23  & n16245;
  assign n16248 = ~n16246 & ~n16247;
  assign n16249 = n15910 & ~n15912;
  assign n16250 = ~n15913 & ~n16249;
  assign n16251 = ~n16248 & n16250;
  assign n16252 = n5267 & n12262;
  assign n16253 = n5185 & n12265;
  assign n16254 = n5121 & n12268;
  assign n16255 = n78 & n14691;
  assign n16256 = ~n16253 & ~n16254;
  assign n16257 = ~n16252 & n16256;
  assign n16258 = ~n16255 & n16257;
  assign n16259 = pi23  & n16258;
  assign n16260 = ~pi23  & ~n16258;
  assign n16261 = ~n16259 & ~n16260;
  assign n16262 = n15906 & ~n15908;
  assign n16263 = ~n15909 & ~n16262;
  assign n16264 = ~n16261 & n16263;
  assign n16265 = n5267 & n12265;
  assign n16266 = n5185 & n12268;
  assign n16267 = n5121 & n12271;
  assign n16268 = n78 & n14728;
  assign n16269 = ~n16266 & ~n16267;
  assign n16270 = ~n16265 & n16269;
  assign n16271 = ~n16268 & n16270;
  assign n16272 = ~pi23  & ~n16271;
  assign n16273 = pi23  & n16271;
  assign n16274 = ~n16272 & ~n16273;
  assign n16275 = pi26  & ~n15886;
  assign n16276 = n15893 & ~n16275;
  assign n16277 = ~n15893 & n16275;
  assign n16278 = ~n16276 & ~n16277;
  assign n16279 = ~n16274 & n16278;
  assign n16280 = n5267 & n12268;
  assign n16281 = n5185 & n12271;
  assign n16282 = n5121 & n12274;
  assign n16283 = n78 & n14771;
  assign n16284 = ~n16281 & ~n16282;
  assign n16285 = ~n16280 & n16284;
  assign n16286 = ~n16283 & n16285;
  assign n16287 = pi23  & n16286;
  assign n16288 = ~pi23  & ~n16286;
  assign n16289 = ~n16287 & ~n16288;
  assign n16290 = n15880 & ~n15885;
  assign n16291 = ~n15886 & ~n16290;
  assign n16292 = ~n16289 & n16291;
  assign n16293 = n74 & n12281;
  assign n16294 = pi23  & n16293;
  assign n16295 = n5267 & n12279;
  assign n16296 = n5185 & n12281;
  assign n16297 = n78 & ~n14833;
  assign n16298 = ~n16295 & ~n16296;
  assign n16299 = ~n16297 & n16298;
  assign n16300 = ~n16294 & n16299;
  assign n16301 = n5267 & n12274;
  assign n16302 = n5185 & n12279;
  assign n16303 = n5121 & n12281;
  assign n16304 = n78 & ~n14876;
  assign n16305 = ~n16302 & ~n16303;
  assign n16306 = ~n16301 & n16305;
  assign n16307 = ~n16304 & n16306;
  assign n16308 = pi23  & n16300;
  assign n16309 = n16307 & n16308;
  assign n16310 = n15879 & n16309;
  assign n16311 = n5267 & n12271;
  assign n16312 = n5185 & n12274;
  assign n16313 = n5121 & n12279;
  assign n16314 = n78 & n14795;
  assign n16315 = ~n16312 & ~n16313;
  assign n16316 = ~n16311 & n16315;
  assign n16317 = ~n16314 & n16316;
  assign n16318 = pi23  & n16317;
  assign n16319 = ~pi23  & ~n16317;
  assign n16320 = ~n16318 & ~n16319;
  assign n16321 = ~n15879 & ~n16309;
  assign n16322 = ~n16310 & ~n16321;
  assign n16323 = ~n16320 & n16322;
  assign n16324 = ~n16310 & ~n16323;
  assign n16325 = n16289 & ~n16291;
  assign n16326 = ~n16292 & ~n16325;
  assign n16327 = ~n16324 & n16326;
  assign n16328 = ~n16292 & ~n16327;
  assign n16329 = n16274 & ~n16278;
  assign n16330 = ~n16279 & ~n16329;
  assign n16331 = ~n16328 & n16330;
  assign n16332 = ~n16279 & ~n16331;
  assign n16333 = n16261 & ~n16263;
  assign n16334 = ~n16264 & ~n16333;
  assign n16335 = ~n16332 & n16334;
  assign n16336 = ~n16264 & ~n16335;
  assign n16337 = n16248 & ~n16250;
  assign n16338 = ~n16251 & ~n16337;
  assign n16339 = ~n16336 & n16338;
  assign n16340 = ~n16251 & ~n16339;
  assign n16341 = ~n16227 & n16237;
  assign n16342 = ~n16238 & ~n16341;
  assign n16343 = ~n16340 & n16342;
  assign n16344 = ~n16238 & ~n16343;
  assign n16345 = ~n16214 & n16224;
  assign n16346 = ~n16225 & ~n16345;
  assign n16347 = ~n16344 & n16346;
  assign n16348 = ~n16225 & ~n16347;
  assign n16349 = n16209 & ~n16211;
  assign n16350 = ~n16212 & ~n16349;
  assign n16351 = ~n16348 & n16350;
  assign n16352 = ~n16212 & ~n16351;
  assign n16353 = n16196 & ~n16198;
  assign n16354 = ~n16199 & ~n16353;
  assign n16355 = ~n16352 & n16354;
  assign n16356 = ~n16199 & ~n16355;
  assign n16357 = n16183 & ~n16185;
  assign n16358 = ~n16186 & ~n16357;
  assign n16359 = ~n16356 & n16358;
  assign n16360 = ~n16186 & ~n16359;
  assign n16361 = n16170 & ~n16172;
  assign n16362 = ~n16173 & ~n16361;
  assign n16363 = ~n16360 & n16362;
  assign n16364 = ~n16173 & ~n16363;
  assign n16365 = n16157 & ~n16159;
  assign n16366 = ~n16160 & ~n16365;
  assign n16367 = ~n16364 & n16366;
  assign n16368 = ~n16160 & ~n16367;
  assign n16369 = n16144 & ~n16146;
  assign n16370 = ~n16147 & ~n16369;
  assign n16371 = ~n16368 & n16370;
  assign n16372 = ~n16147 & ~n16371;
  assign n16373 = n16131 & ~n16133;
  assign n16374 = ~n16134 & ~n16373;
  assign n16375 = ~n16372 & n16374;
  assign n16376 = ~n16134 & ~n16375;
  assign n16377 = n16118 & ~n16120;
  assign n16378 = ~n16121 & ~n16377;
  assign n16379 = ~n16376 & n16378;
  assign n16380 = ~n16121 & ~n16379;
  assign n16381 = n16105 & ~n16107;
  assign n16382 = ~n16108 & ~n16381;
  assign n16383 = ~n16380 & n16382;
  assign n16384 = ~n16108 & ~n16383;
  assign n16385 = n16092 & ~n16094;
  assign n16386 = ~n16095 & ~n16385;
  assign n16387 = ~n16384 & n16386;
  assign n16388 = ~n16095 & ~n16387;
  assign n16389 = ~n15965 & n15975;
  assign n16390 = ~n15976 & ~n16389;
  assign n16391 = ~n16388 & n16390;
  assign n16392 = n16388 & ~n16390;
  assign n16393 = ~n16391 & ~n16392;
  assign n16394 = n5982 & n12211;
  assign n16395 = n5901 & n12214;
  assign n16396 = n5312 & n12217;
  assign n16397 = n5306 & n13203;
  assign n16398 = ~n16395 & ~n16396;
  assign n16399 = ~n16394 & n16398;
  assign n16400 = ~n16397 & n16399;
  assign n16401 = pi20  & n16400;
  assign n16402 = ~pi20  & ~n16400;
  assign n16403 = ~n16401 & ~n16402;
  assign n16404 = n16393 & ~n16403;
  assign n16405 = ~n16391 & ~n16404;
  assign n16406 = ~n15982 & n15992;
  assign n16407 = ~n15993 & ~n16406;
  assign n16408 = ~n16405 & n16407;
  assign n16409 = n16405 & ~n16407;
  assign n16410 = ~n16408 & ~n16409;
  assign n16411 = n6608 & n12199;
  assign n16412 = n6356 & n12202;
  assign n16413 = n6140 & n12205;
  assign n16414 = n6134 & n12683;
  assign n16415 = ~n16412 & ~n16413;
  assign n16416 = ~n16411 & n16415;
  assign n16417 = ~n16414 & n16416;
  assign n16418 = pi17  & n16417;
  assign n16419 = ~pi17  & ~n16417;
  assign n16420 = ~n16418 & ~n16419;
  assign n16421 = n16410 & ~n16420;
  assign n16422 = ~n16408 & ~n16421;
  assign n16423 = ~n15999 & n16009;
  assign n16424 = ~n16010 & ~n16423;
  assign n16425 = ~n16422 & n16424;
  assign n16426 = n16422 & ~n16424;
  assign n16427 = ~n16425 & ~n16426;
  assign n16428 = n7380 & n12187;
  assign n16429 = n7243 & n12190;
  assign n16430 = n6653 & n12193;
  assign n16431 = n6647 & n12921;
  assign n16432 = ~n16429 & ~n16430;
  assign n16433 = ~n16428 & n16432;
  assign n16434 = ~n16431 & n16433;
  assign n16435 = pi14  & n16434;
  assign n16436 = ~pi14  & ~n16434;
  assign n16437 = ~n16435 & ~n16436;
  assign n16438 = n16427 & ~n16437;
  assign n16439 = ~n16425 & ~n16438;
  assign n16440 = ~n16071 & n16081;
  assign n16441 = ~n16082 & ~n16440;
  assign n16442 = ~n16439 & n16441;
  assign n16443 = ~n16082 & ~n16442;
  assign n16444 = ~n16020 & n16030;
  assign n16445 = ~n16031 & ~n16444;
  assign n16446 = ~n16443 & n16445;
  assign n16447 = n16443 & ~n16445;
  assign n16448 = ~n16446 & ~n16447;
  assign n16449 = n8161 & n12168;
  assign n16450 = n7847 & n12175;
  assign n16451 = n7554 & n12178;
  assign n16452 = n7548 & n12862;
  assign n16453 = ~n16450 & ~n16451;
  assign n16454 = ~n16449 & n16453;
  assign n16455 = ~n16452 & n16454;
  assign n16456 = pi11  & n16455;
  assign n16457 = ~pi11  & ~n16455;
  assign n16458 = ~n16456 & ~n16457;
  assign n16459 = n16448 & ~n16458;
  assign n16460 = ~n16446 & ~n16459;
  assign n16461 = n8200 & ~n12424;
  assign n16462 = n8205 & ~n12165;
  assign n16463 = n13513 & ~n16462;
  assign n16464 = ~n12163 & ~n16463;
  assign n16465 = ~n16461 & ~n16464;
  assign n16466 = pi8  & n16465;
  assign n16467 = ~pi8  & ~n16465;
  assign n16468 = ~n16466 & ~n16467;
  assign n16469 = ~n16460 & ~n16468;
  assign n16470 = n16460 & n16468;
  assign n16471 = ~n16469 & ~n16470;
  assign n16472 = ~n16037 & n16047;
  assign n16473 = ~n16048 & ~n16472;
  assign n16474 = n16471 & n16473;
  assign n16475 = ~n16469 & ~n16474;
  assign n16476 = ~n16062 & ~n16064;
  assign n16477 = ~n16065 & ~n16476;
  assign n16478 = ~n16475 & n16477;
  assign n16479 = n16439 & ~n16441;
  assign n16480 = ~n16442 & ~n16479;
  assign n16481 = n8161 & n12175;
  assign n16482 = n7847 & n12178;
  assign n16483 = n7554 & n12181;
  assign n16484 = n7548 & n12961;
  assign n16485 = ~n16482 & ~n16483;
  assign n16486 = ~n16481 & n16485;
  assign n16487 = ~n16484 & n16486;
  assign n16488 = pi11  & n16487;
  assign n16489 = ~pi11  & ~n16487;
  assign n16490 = ~n16488 & ~n16489;
  assign n16491 = n16480 & ~n16490;
  assign n16492 = n16384 & ~n16386;
  assign n16493 = ~n16387 & ~n16492;
  assign n16494 = n5982 & n12214;
  assign n16495 = n5901 & n12217;
  assign n16496 = n5312 & n12220;
  assign n16497 = n5306 & n13187;
  assign n16498 = ~n16495 & ~n16496;
  assign n16499 = ~n16494 & n16498;
  assign n16500 = ~n16497 & n16499;
  assign n16501 = pi20  & n16500;
  assign n16502 = ~pi20  & ~n16500;
  assign n16503 = ~n16501 & ~n16502;
  assign n16504 = n16493 & ~n16503;
  assign n16505 = n16380 & ~n16382;
  assign n16506 = ~n16383 & ~n16505;
  assign n16507 = n5982 & n12217;
  assign n16508 = n5901 & n12220;
  assign n16509 = n5312 & n12223;
  assign n16510 = n5306 & n13374;
  assign n16511 = ~n16508 & ~n16509;
  assign n16512 = ~n16507 & n16511;
  assign n16513 = ~n16510 & n16512;
  assign n16514 = pi20  & n16513;
  assign n16515 = ~pi20  & ~n16513;
  assign n16516 = ~n16514 & ~n16515;
  assign n16517 = n16506 & ~n16516;
  assign n16518 = n16376 & ~n16378;
  assign n16519 = ~n16379 & ~n16518;
  assign n16520 = n5982 & n12220;
  assign n16521 = n5901 & n12223;
  assign n16522 = n5312 & n12226;
  assign n16523 = n5306 & n13392;
  assign n16524 = ~n16521 & ~n16522;
  assign n16525 = ~n16520 & n16524;
  assign n16526 = ~n16523 & n16525;
  assign n16527 = pi20  & n16526;
  assign n16528 = ~pi20  & ~n16526;
  assign n16529 = ~n16527 & ~n16528;
  assign n16530 = n16519 & ~n16529;
  assign n16531 = n16372 & ~n16374;
  assign n16532 = ~n16375 & ~n16531;
  assign n16533 = n5982 & n12223;
  assign n16534 = n5901 & n12226;
  assign n16535 = n5312 & n12229;
  assign n16536 = n5306 & n13745;
  assign n16537 = ~n16534 & ~n16535;
  assign n16538 = ~n16533 & n16537;
  assign n16539 = ~n16536 & n16538;
  assign n16540 = pi20  & n16539;
  assign n16541 = ~pi20  & ~n16539;
  assign n16542 = ~n16540 & ~n16541;
  assign n16543 = n16532 & ~n16542;
  assign n16544 = n16368 & ~n16370;
  assign n16545 = ~n16371 & ~n16544;
  assign n16546 = n5982 & n12226;
  assign n16547 = n5901 & n12229;
  assign n16548 = n5312 & n12232;
  assign n16549 = n5306 & n13530;
  assign n16550 = ~n16547 & ~n16548;
  assign n16551 = ~n16546 & n16550;
  assign n16552 = ~n16549 & n16551;
  assign n16553 = pi20  & n16552;
  assign n16554 = ~pi20  & ~n16552;
  assign n16555 = ~n16553 & ~n16554;
  assign n16556 = n16545 & ~n16555;
  assign n16557 = n16364 & ~n16366;
  assign n16558 = ~n16367 & ~n16557;
  assign n16559 = n5982 & n12229;
  assign n16560 = n5901 & n12232;
  assign n16561 = n5312 & n12235;
  assign n16562 = n5306 & n13979;
  assign n16563 = ~n16560 & ~n16561;
  assign n16564 = ~n16559 & n16563;
  assign n16565 = ~n16562 & n16564;
  assign n16566 = pi20  & n16565;
  assign n16567 = ~pi20  & ~n16565;
  assign n16568 = ~n16566 & ~n16567;
  assign n16569 = n16558 & ~n16568;
  assign n16570 = n16360 & ~n16362;
  assign n16571 = ~n16363 & ~n16570;
  assign n16572 = n5982 & n12232;
  assign n16573 = n5901 & n12235;
  assign n16574 = n5312 & n12238;
  assign n16575 = n5306 & n14116;
  assign n16576 = ~n16573 & ~n16574;
  assign n16577 = ~n16572 & n16576;
  assign n16578 = ~n16575 & n16577;
  assign n16579 = pi20  & n16578;
  assign n16580 = ~pi20  & ~n16578;
  assign n16581 = ~n16579 & ~n16580;
  assign n16582 = n16571 & ~n16581;
  assign n16583 = n16356 & ~n16358;
  assign n16584 = ~n16359 & ~n16583;
  assign n16585 = n5982 & n12235;
  assign n16586 = n5901 & n12238;
  assign n16587 = n5312 & n12241;
  assign n16588 = n5306 & n13959;
  assign n16589 = ~n16586 & ~n16587;
  assign n16590 = ~n16585 & n16589;
  assign n16591 = ~n16588 & n16590;
  assign n16592 = pi20  & n16591;
  assign n16593 = ~pi20  & ~n16591;
  assign n16594 = ~n16592 & ~n16593;
  assign n16595 = n16584 & ~n16594;
  assign n16596 = n16352 & ~n16354;
  assign n16597 = ~n16355 & ~n16596;
  assign n16598 = n5982 & n12238;
  assign n16599 = n5901 & n12241;
  assign n16600 = n5312 & n12244;
  assign n16601 = n5306 & n14229;
  assign n16602 = ~n16599 & ~n16600;
  assign n16603 = ~n16598 & n16602;
  assign n16604 = ~n16601 & n16603;
  assign n16605 = pi20  & n16604;
  assign n16606 = ~pi20  & ~n16604;
  assign n16607 = ~n16605 & ~n16606;
  assign n16608 = n16597 & ~n16607;
  assign n16609 = n16348 & ~n16350;
  assign n16610 = ~n16351 & ~n16609;
  assign n16611 = n5982 & n12241;
  assign n16612 = n5901 & n12244;
  assign n16613 = n5312 & n12247;
  assign n16614 = n5306 & n14515;
  assign n16615 = ~n16612 & ~n16613;
  assign n16616 = ~n16611 & n16615;
  assign n16617 = ~n16614 & n16616;
  assign n16618 = pi20  & n16617;
  assign n16619 = ~pi20  & ~n16617;
  assign n16620 = ~n16618 & ~n16619;
  assign n16621 = n16610 & ~n16620;
  assign n16622 = n5982 & n12244;
  assign n16623 = n5901 & n12247;
  assign n16624 = n5312 & n12250;
  assign n16625 = n5306 & n14527;
  assign n16626 = ~n16623 & ~n16624;
  assign n16627 = ~n16622 & n16626;
  assign n16628 = ~n16625 & n16627;
  assign n16629 = ~pi20  & ~n16628;
  assign n16630 = pi20  & n16628;
  assign n16631 = ~n16629 & ~n16630;
  assign n16632 = n16344 & ~n16346;
  assign n16633 = ~n16347 & ~n16632;
  assign n16634 = ~n16631 & n16633;
  assign n16635 = n5982 & n12247;
  assign n16636 = n5901 & n12250;
  assign n16637 = n5312 & n12253;
  assign n16638 = n5306 & n14207;
  assign n16639 = ~n16636 & ~n16637;
  assign n16640 = ~n16635 & n16639;
  assign n16641 = ~n16638 & n16640;
  assign n16642 = ~pi20  & ~n16641;
  assign n16643 = pi20  & n16641;
  assign n16644 = ~n16642 & ~n16643;
  assign n16645 = n16340 & ~n16342;
  assign n16646 = ~n16343 & ~n16645;
  assign n16647 = ~n16644 & n16646;
  assign n16648 = n16336 & ~n16338;
  assign n16649 = ~n16339 & ~n16648;
  assign n16650 = n5982 & n12250;
  assign n16651 = n5901 & n12253;
  assign n16652 = n5312 & n12256;
  assign n16653 = n5306 & n14559;
  assign n16654 = ~n16651 & ~n16652;
  assign n16655 = ~n16650 & n16654;
  assign n16656 = ~n16653 & n16655;
  assign n16657 = pi20  & n16656;
  assign n16658 = ~pi20  & ~n16656;
  assign n16659 = ~n16657 & ~n16658;
  assign n16660 = n16649 & ~n16659;
  assign n16661 = n16332 & ~n16334;
  assign n16662 = ~n16335 & ~n16661;
  assign n16663 = n5982 & n12253;
  assign n16664 = n5901 & n12256;
  assign n16665 = n5312 & n12259;
  assign n16666 = n5306 & n14584;
  assign n16667 = ~n16664 & ~n16665;
  assign n16668 = ~n16663 & n16667;
  assign n16669 = ~n16666 & n16668;
  assign n16670 = pi20  & n16669;
  assign n16671 = ~pi20  & ~n16669;
  assign n16672 = ~n16670 & ~n16671;
  assign n16673 = n16662 & ~n16672;
  assign n16674 = n16328 & ~n16330;
  assign n16675 = ~n16331 & ~n16674;
  assign n16676 = n5982 & n12256;
  assign n16677 = n5901 & n12259;
  assign n16678 = n5312 & n12262;
  assign n16679 = n5306 & n14608;
  assign n16680 = ~n16677 & ~n16678;
  assign n16681 = ~n16676 & n16680;
  assign n16682 = ~n16679 & n16681;
  assign n16683 = pi20  & n16682;
  assign n16684 = ~pi20  & ~n16682;
  assign n16685 = ~n16683 & ~n16684;
  assign n16686 = n16675 & ~n16685;
  assign n16687 = n5982 & n12259;
  assign n16688 = n5901 & n12262;
  assign n16689 = n5312 & n12265;
  assign n16690 = n5306 & n14637;
  assign n16691 = ~n16688 & ~n16689;
  assign n16692 = ~n16687 & n16691;
  assign n16693 = ~n16690 & n16692;
  assign n16694 = ~pi20  & ~n16693;
  assign n16695 = pi20  & n16693;
  assign n16696 = ~n16694 & ~n16695;
  assign n16697 = n16324 & ~n16326;
  assign n16698 = ~n16327 & ~n16697;
  assign n16699 = ~n16696 & n16698;
  assign n16700 = n5982 & n12262;
  assign n16701 = n5901 & n12265;
  assign n16702 = n5312 & n12268;
  assign n16703 = n5306 & n14691;
  assign n16704 = ~n16701 & ~n16702;
  assign n16705 = ~n16700 & n16704;
  assign n16706 = ~n16703 & n16705;
  assign n16707 = pi20  & n16706;
  assign n16708 = ~pi20  & ~n16706;
  assign n16709 = ~n16707 & ~n16708;
  assign n16710 = n16320 & ~n16322;
  assign n16711 = ~n16323 & ~n16710;
  assign n16712 = ~n16709 & n16711;
  assign n16713 = n5982 & n12265;
  assign n16714 = n5901 & n12268;
  assign n16715 = n5312 & n12271;
  assign n16716 = n5306 & n14728;
  assign n16717 = ~n16714 & ~n16715;
  assign n16718 = ~n16713 & n16717;
  assign n16719 = ~n16716 & n16718;
  assign n16720 = ~pi20  & ~n16719;
  assign n16721 = pi20  & n16719;
  assign n16722 = ~n16720 & ~n16721;
  assign n16723 = pi23  & ~n16300;
  assign n16724 = n16307 & ~n16723;
  assign n16725 = ~n16307 & n16723;
  assign n16726 = ~n16724 & ~n16725;
  assign n16727 = ~n16722 & n16726;
  assign n16728 = n5982 & n12268;
  assign n16729 = n5901 & n12271;
  assign n16730 = n5312 & n12274;
  assign n16731 = n5306 & n14771;
  assign n16732 = ~n16729 & ~n16730;
  assign n16733 = ~n16728 & n16732;
  assign n16734 = ~n16731 & n16733;
  assign n16735 = pi20  & n16734;
  assign n16736 = ~pi20  & ~n16734;
  assign n16737 = ~n16735 & ~n16736;
  assign n16738 = n16294 & ~n16299;
  assign n16739 = ~n16300 & ~n16738;
  assign n16740 = ~n16737 & n16739;
  assign n16741 = n5305 & n12281;
  assign n16742 = pi20  & n16741;
  assign n16743 = n5982 & n12279;
  assign n16744 = n5901 & n12281;
  assign n16745 = n5306 & ~n14833;
  assign n16746 = ~n16743 & ~n16744;
  assign n16747 = ~n16745 & n16746;
  assign n16748 = ~n16742 & n16747;
  assign n16749 = n5982 & n12274;
  assign n16750 = n5901 & n12279;
  assign n16751 = n5312 & n12281;
  assign n16752 = n5306 & ~n14876;
  assign n16753 = ~n16750 & ~n16751;
  assign n16754 = ~n16749 & n16753;
  assign n16755 = ~n16752 & n16754;
  assign n16756 = pi20  & n16748;
  assign n16757 = n16755 & n16756;
  assign n16758 = n16293 & n16757;
  assign n16759 = n5982 & n12271;
  assign n16760 = n5901 & n12274;
  assign n16761 = n5312 & n12279;
  assign n16762 = n5306 & n14795;
  assign n16763 = ~n16760 & ~n16761;
  assign n16764 = ~n16759 & n16763;
  assign n16765 = ~n16762 & n16764;
  assign n16766 = pi20  & n16765;
  assign n16767 = ~pi20  & ~n16765;
  assign n16768 = ~n16766 & ~n16767;
  assign n16769 = ~n16293 & ~n16757;
  assign n16770 = ~n16758 & ~n16769;
  assign n16771 = ~n16768 & n16770;
  assign n16772 = ~n16758 & ~n16771;
  assign n16773 = n16737 & ~n16739;
  assign n16774 = ~n16740 & ~n16773;
  assign n16775 = ~n16772 & n16774;
  assign n16776 = ~n16740 & ~n16775;
  assign n16777 = n16722 & ~n16726;
  assign n16778 = ~n16727 & ~n16777;
  assign n16779 = ~n16776 & n16778;
  assign n16780 = ~n16727 & ~n16779;
  assign n16781 = n16709 & ~n16711;
  assign n16782 = ~n16712 & ~n16781;
  assign n16783 = ~n16780 & n16782;
  assign n16784 = ~n16712 & ~n16783;
  assign n16785 = n16696 & ~n16698;
  assign n16786 = ~n16699 & ~n16785;
  assign n16787 = ~n16784 & n16786;
  assign n16788 = ~n16699 & ~n16787;
  assign n16789 = ~n16675 & n16685;
  assign n16790 = ~n16686 & ~n16789;
  assign n16791 = ~n16788 & n16790;
  assign n16792 = ~n16686 & ~n16791;
  assign n16793 = ~n16662 & n16672;
  assign n16794 = ~n16673 & ~n16793;
  assign n16795 = ~n16792 & n16794;
  assign n16796 = ~n16673 & ~n16795;
  assign n16797 = ~n16649 & n16659;
  assign n16798 = ~n16660 & ~n16797;
  assign n16799 = ~n16796 & n16798;
  assign n16800 = ~n16660 & ~n16799;
  assign n16801 = n16644 & ~n16646;
  assign n16802 = ~n16647 & ~n16801;
  assign n16803 = ~n16800 & n16802;
  assign n16804 = ~n16647 & ~n16803;
  assign n16805 = n16631 & ~n16633;
  assign n16806 = ~n16634 & ~n16805;
  assign n16807 = ~n16804 & n16806;
  assign n16808 = ~n16634 & ~n16807;
  assign n16809 = ~n16610 & n16620;
  assign n16810 = ~n16621 & ~n16809;
  assign n16811 = ~n16808 & n16810;
  assign n16812 = ~n16621 & ~n16811;
  assign n16813 = ~n16597 & n16607;
  assign n16814 = ~n16608 & ~n16813;
  assign n16815 = ~n16812 & n16814;
  assign n16816 = ~n16608 & ~n16815;
  assign n16817 = ~n16584 & n16594;
  assign n16818 = ~n16595 & ~n16817;
  assign n16819 = ~n16816 & n16818;
  assign n16820 = ~n16595 & ~n16819;
  assign n16821 = ~n16571 & n16581;
  assign n16822 = ~n16582 & ~n16821;
  assign n16823 = ~n16820 & n16822;
  assign n16824 = ~n16582 & ~n16823;
  assign n16825 = ~n16558 & n16568;
  assign n16826 = ~n16569 & ~n16825;
  assign n16827 = ~n16824 & n16826;
  assign n16828 = ~n16569 & ~n16827;
  assign n16829 = ~n16545 & n16555;
  assign n16830 = ~n16556 & ~n16829;
  assign n16831 = ~n16828 & n16830;
  assign n16832 = ~n16556 & ~n16831;
  assign n16833 = ~n16532 & n16542;
  assign n16834 = ~n16543 & ~n16833;
  assign n16835 = ~n16832 & n16834;
  assign n16836 = ~n16543 & ~n16835;
  assign n16837 = ~n16519 & n16529;
  assign n16838 = ~n16530 & ~n16837;
  assign n16839 = ~n16836 & n16838;
  assign n16840 = ~n16530 & ~n16839;
  assign n16841 = ~n16506 & n16516;
  assign n16842 = ~n16517 & ~n16841;
  assign n16843 = ~n16840 & n16842;
  assign n16844 = ~n16517 & ~n16843;
  assign n16845 = ~n16493 & n16503;
  assign n16846 = ~n16504 & ~n16845;
  assign n16847 = ~n16844 & n16846;
  assign n16848 = ~n16504 & ~n16847;
  assign n16849 = ~n16393 & n16403;
  assign n16850 = ~n16404 & ~n16849;
  assign n16851 = ~n16848 & n16850;
  assign n16852 = n16848 & ~n16850;
  assign n16853 = ~n16851 & ~n16852;
  assign n16854 = n6608 & n12202;
  assign n16855 = n6356 & n12205;
  assign n16856 = n6140 & n12208;
  assign n16857 = n6134 & n12701;
  assign n16858 = ~n16855 & ~n16856;
  assign n16859 = ~n16854 & n16858;
  assign n16860 = ~n16857 & n16859;
  assign n16861 = pi17  & n16860;
  assign n16862 = ~pi17  & ~n16860;
  assign n16863 = ~n16861 & ~n16862;
  assign n16864 = n16853 & ~n16863;
  assign n16865 = ~n16851 & ~n16864;
  assign n16866 = ~n16410 & n16420;
  assign n16867 = ~n16421 & ~n16866;
  assign n16868 = ~n16865 & n16867;
  assign n16869 = n16865 & ~n16867;
  assign n16870 = ~n16868 & ~n16869;
  assign n16871 = n7380 & n12190;
  assign n16872 = n7243 & n12193;
  assign n16873 = n6653 & n12196;
  assign n16874 = n6647 & n12530;
  assign n16875 = ~n16872 & ~n16873;
  assign n16876 = ~n16871 & n16875;
  assign n16877 = ~n16874 & n16876;
  assign n16878 = pi14  & n16877;
  assign n16879 = ~pi14  & ~n16877;
  assign n16880 = ~n16878 & ~n16879;
  assign n16881 = n16870 & ~n16880;
  assign n16882 = ~n16868 & ~n16881;
  assign n16883 = ~n16427 & n16437;
  assign n16884 = ~n16438 & ~n16883;
  assign n16885 = ~n16882 & n16884;
  assign n16886 = n16882 & ~n16884;
  assign n16887 = ~n16885 & ~n16886;
  assign n16888 = n8161 & n12178;
  assign n16889 = n7847 & n12181;
  assign n16890 = n7554 & n12184;
  assign n16891 = n7548 & n12880;
  assign n16892 = ~n16889 & ~n16890;
  assign n16893 = ~n16888 & n16892;
  assign n16894 = ~n16891 & n16893;
  assign n16895 = pi11  & n16894;
  assign n16896 = ~pi11  & ~n16894;
  assign n16897 = ~n16895 & ~n16896;
  assign n16898 = n16887 & ~n16897;
  assign n16899 = ~n16885 & ~n16898;
  assign n16900 = ~n16480 & n16490;
  assign n16901 = ~n16491 & ~n16900;
  assign n16902 = ~n16899 & n16901;
  assign n16903 = ~n16491 & ~n16902;
  assign n16904 = ~n16448 & n16458;
  assign n16905 = ~n16459 & ~n16904;
  assign n16906 = ~n16903 & n16905;
  assign n16907 = n16903 & ~n16905;
  assign n16908 = ~n16906 & ~n16907;
  assign n16909 = n8200 & n13007;
  assign n16910 = n8206 & n12172;
  assign n16911 = ~n9355 & n12165;
  assign n16912 = ~n12163 & ~n13513;
  assign n16913 = ~n16911 & n16912;
  assign n16914 = ~n16910 & ~n16913;
  assign n16915 = ~n16909 & n16914;
  assign n16916 = pi8  & n16915;
  assign n16917 = ~pi8  & ~n16915;
  assign n16918 = ~n16916 & ~n16917;
  assign n16919 = n16908 & ~n16918;
  assign n16920 = ~n16906 & ~n16919;
  assign n16921 = ~n16471 & ~n16473;
  assign n16922 = ~n16474 & ~n16921;
  assign n16923 = ~n16920 & n16922;
  assign n16924 = n16920 & ~n16922;
  assign n16925 = ~n16923 & ~n16924;
  assign n16926 = n6608 & n12205;
  assign n16927 = n6356 & n12208;
  assign n16928 = n6140 & n12211;
  assign n16929 = n6134 & n13031;
  assign n16930 = ~n16927 & ~n16928;
  assign n16931 = ~n16926 & n16930;
  assign n16932 = ~n16929 & n16931;
  assign n16933 = ~pi17  & ~n16932;
  assign n16934 = pi17  & n16932;
  assign n16935 = ~n16933 & ~n16934;
  assign n16936 = n16844 & ~n16846;
  assign n16937 = ~n16847 & ~n16936;
  assign n16938 = ~n16935 & n16937;
  assign n16939 = n6608 & n12208;
  assign n16940 = n6356 & n12211;
  assign n16941 = n6140 & n12214;
  assign n16942 = n6134 & n12804;
  assign n16943 = ~n16940 & ~n16941;
  assign n16944 = ~n16939 & n16943;
  assign n16945 = ~n16942 & n16944;
  assign n16946 = ~pi17  & ~n16945;
  assign n16947 = pi17  & n16945;
  assign n16948 = ~n16946 & ~n16947;
  assign n16949 = n16840 & ~n16842;
  assign n16950 = ~n16843 & ~n16949;
  assign n16951 = ~n16948 & n16950;
  assign n16952 = n6608 & n12211;
  assign n16953 = n6356 & n12214;
  assign n16954 = n6140 & n12217;
  assign n16955 = n6134 & n13203;
  assign n16956 = ~n16953 & ~n16954;
  assign n16957 = ~n16952 & n16956;
  assign n16958 = ~n16955 & n16957;
  assign n16959 = ~pi17  & ~n16958;
  assign n16960 = pi17  & n16958;
  assign n16961 = ~n16959 & ~n16960;
  assign n16962 = n16836 & ~n16838;
  assign n16963 = ~n16839 & ~n16962;
  assign n16964 = ~n16961 & n16963;
  assign n16965 = n6608 & n12214;
  assign n16966 = n6356 & n12217;
  assign n16967 = n6140 & n12220;
  assign n16968 = n6134 & n13187;
  assign n16969 = ~n16966 & ~n16967;
  assign n16970 = ~n16965 & n16969;
  assign n16971 = ~n16968 & n16970;
  assign n16972 = ~pi17  & ~n16971;
  assign n16973 = pi17  & n16971;
  assign n16974 = ~n16972 & ~n16973;
  assign n16975 = n16832 & ~n16834;
  assign n16976 = ~n16835 & ~n16975;
  assign n16977 = ~n16974 & n16976;
  assign n16978 = n6608 & n12217;
  assign n16979 = n6356 & n12220;
  assign n16980 = n6140 & n12223;
  assign n16981 = n6134 & n13374;
  assign n16982 = ~n16979 & ~n16980;
  assign n16983 = ~n16978 & n16982;
  assign n16984 = ~n16981 & n16983;
  assign n16985 = ~pi17  & ~n16984;
  assign n16986 = pi17  & n16984;
  assign n16987 = ~n16985 & ~n16986;
  assign n16988 = n16828 & ~n16830;
  assign n16989 = ~n16831 & ~n16988;
  assign n16990 = ~n16987 & n16989;
  assign n16991 = n6608 & n12220;
  assign n16992 = n6356 & n12223;
  assign n16993 = n6140 & n12226;
  assign n16994 = n6134 & n13392;
  assign n16995 = ~n16992 & ~n16993;
  assign n16996 = ~n16991 & n16995;
  assign n16997 = ~n16994 & n16996;
  assign n16998 = ~pi17  & ~n16997;
  assign n16999 = pi17  & n16997;
  assign n17000 = ~n16998 & ~n16999;
  assign n17001 = n16824 & ~n16826;
  assign n17002 = ~n16827 & ~n17001;
  assign n17003 = ~n17000 & n17002;
  assign n17004 = n6608 & n12223;
  assign n17005 = n6356 & n12226;
  assign n17006 = n6140 & n12229;
  assign n17007 = n6134 & n13745;
  assign n17008 = ~n17005 & ~n17006;
  assign n17009 = ~n17004 & n17008;
  assign n17010 = ~n17007 & n17009;
  assign n17011 = ~pi17  & ~n17010;
  assign n17012 = pi17  & n17010;
  assign n17013 = ~n17011 & ~n17012;
  assign n17014 = n16820 & ~n16822;
  assign n17015 = ~n16823 & ~n17014;
  assign n17016 = ~n17013 & n17015;
  assign n17017 = n6608 & n12226;
  assign n17018 = n6356 & n12229;
  assign n17019 = n6140 & n12232;
  assign n17020 = n6134 & n13530;
  assign n17021 = ~n17018 & ~n17019;
  assign n17022 = ~n17017 & n17021;
  assign n17023 = ~n17020 & n17022;
  assign n17024 = ~pi17  & ~n17023;
  assign n17025 = pi17  & n17023;
  assign n17026 = ~n17024 & ~n17025;
  assign n17027 = n16816 & ~n16818;
  assign n17028 = ~n16819 & ~n17027;
  assign n17029 = ~n17026 & n17028;
  assign n17030 = n6608 & n12229;
  assign n17031 = n6356 & n12232;
  assign n17032 = n6140 & n12235;
  assign n17033 = n6134 & n13979;
  assign n17034 = ~n17031 & ~n17032;
  assign n17035 = ~n17030 & n17034;
  assign n17036 = ~n17033 & n17035;
  assign n17037 = ~pi17  & ~n17036;
  assign n17038 = pi17  & n17036;
  assign n17039 = ~n17037 & ~n17038;
  assign n17040 = n16812 & ~n16814;
  assign n17041 = ~n16815 & ~n17040;
  assign n17042 = ~n17039 & n17041;
  assign n17043 = n6608 & n12232;
  assign n17044 = n6356 & n12235;
  assign n17045 = n6140 & n12238;
  assign n17046 = n6134 & n14116;
  assign n17047 = ~n17044 & ~n17045;
  assign n17048 = ~n17043 & n17047;
  assign n17049 = ~n17046 & n17048;
  assign n17050 = ~pi17  & ~n17049;
  assign n17051 = pi17  & n17049;
  assign n17052 = ~n17050 & ~n17051;
  assign n17053 = n16808 & ~n16810;
  assign n17054 = ~n16811 & ~n17053;
  assign n17055 = ~n17052 & n17054;
  assign n17056 = n16804 & ~n16806;
  assign n17057 = ~n16807 & ~n17056;
  assign n17058 = n6608 & n12235;
  assign n17059 = n6356 & n12238;
  assign n17060 = n6140 & n12241;
  assign n17061 = n6134 & n13959;
  assign n17062 = ~n17059 & ~n17060;
  assign n17063 = ~n17058 & n17062;
  assign n17064 = ~n17061 & n17063;
  assign n17065 = pi17  & n17064;
  assign n17066 = ~pi17  & ~n17064;
  assign n17067 = ~n17065 & ~n17066;
  assign n17068 = n17057 & ~n17067;
  assign n17069 = n16800 & ~n16802;
  assign n17070 = ~n16803 & ~n17069;
  assign n17071 = n6608 & n12238;
  assign n17072 = n6356 & n12241;
  assign n17073 = n6140 & n12244;
  assign n17074 = n6134 & n14229;
  assign n17075 = ~n17072 & ~n17073;
  assign n17076 = ~n17071 & n17075;
  assign n17077 = ~n17074 & n17076;
  assign n17078 = pi17  & n17077;
  assign n17079 = ~pi17  & ~n17077;
  assign n17080 = ~n17078 & ~n17079;
  assign n17081 = n17070 & ~n17080;
  assign n17082 = n6608 & n12241;
  assign n17083 = n6356 & n12244;
  assign n17084 = n6140 & n12247;
  assign n17085 = n6134 & n14515;
  assign n17086 = ~n17083 & ~n17084;
  assign n17087 = ~n17082 & n17086;
  assign n17088 = ~n17085 & n17087;
  assign n17089 = ~pi17  & ~n17088;
  assign n17090 = pi17  & n17088;
  assign n17091 = ~n17089 & ~n17090;
  assign n17092 = n16796 & ~n16798;
  assign n17093 = ~n16799 & ~n17092;
  assign n17094 = ~n17091 & n17093;
  assign n17095 = n6608 & n12244;
  assign n17096 = n6356 & n12247;
  assign n17097 = n6140 & n12250;
  assign n17098 = n6134 & n14527;
  assign n17099 = ~n17096 & ~n17097;
  assign n17100 = ~n17095 & n17099;
  assign n17101 = ~n17098 & n17100;
  assign n17102 = ~pi17  & ~n17101;
  assign n17103 = pi17  & n17101;
  assign n17104 = ~n17102 & ~n17103;
  assign n17105 = n16792 & ~n16794;
  assign n17106 = ~n16795 & ~n17105;
  assign n17107 = ~n17104 & n17106;
  assign n17108 = n6608 & n12247;
  assign n17109 = n6356 & n12250;
  assign n17110 = n6140 & n12253;
  assign n17111 = n6134 & n14207;
  assign n17112 = ~n17109 & ~n17110;
  assign n17113 = ~n17108 & n17112;
  assign n17114 = ~n17111 & n17113;
  assign n17115 = ~pi17  & ~n17114;
  assign n17116 = pi17  & n17114;
  assign n17117 = ~n17115 & ~n17116;
  assign n17118 = n16788 & ~n16790;
  assign n17119 = ~n16791 & ~n17118;
  assign n17120 = ~n17117 & n17119;
  assign n17121 = n16784 & ~n16786;
  assign n17122 = ~n16787 & ~n17121;
  assign n17123 = n6608 & n12250;
  assign n17124 = n6356 & n12253;
  assign n17125 = n6140 & n12256;
  assign n17126 = n6134 & n14559;
  assign n17127 = ~n17124 & ~n17125;
  assign n17128 = ~n17123 & n17127;
  assign n17129 = ~n17126 & n17128;
  assign n17130 = pi17  & n17129;
  assign n17131 = ~pi17  & ~n17129;
  assign n17132 = ~n17130 & ~n17131;
  assign n17133 = n17122 & ~n17132;
  assign n17134 = n16780 & ~n16782;
  assign n17135 = ~n16783 & ~n17134;
  assign n17136 = n6608 & n12253;
  assign n17137 = n6356 & n12256;
  assign n17138 = n6140 & n12259;
  assign n17139 = n6134 & n14584;
  assign n17140 = ~n17137 & ~n17138;
  assign n17141 = ~n17136 & n17140;
  assign n17142 = ~n17139 & n17141;
  assign n17143 = pi17  & n17142;
  assign n17144 = ~pi17  & ~n17142;
  assign n17145 = ~n17143 & ~n17144;
  assign n17146 = n17135 & ~n17145;
  assign n17147 = n16776 & ~n16778;
  assign n17148 = ~n16779 & ~n17147;
  assign n17149 = n6608 & n12256;
  assign n17150 = n6356 & n12259;
  assign n17151 = n6140 & n12262;
  assign n17152 = n6134 & n14608;
  assign n17153 = ~n17150 & ~n17151;
  assign n17154 = ~n17149 & n17153;
  assign n17155 = ~n17152 & n17154;
  assign n17156 = pi17  & n17155;
  assign n17157 = ~pi17  & ~n17155;
  assign n17158 = ~n17156 & ~n17157;
  assign n17159 = n17148 & ~n17158;
  assign n17160 = n6608 & n12259;
  assign n17161 = n6356 & n12262;
  assign n17162 = n6140 & n12265;
  assign n17163 = n6134 & n14637;
  assign n17164 = ~n17161 & ~n17162;
  assign n17165 = ~n17160 & n17164;
  assign n17166 = ~n17163 & n17165;
  assign n17167 = ~pi17  & ~n17166;
  assign n17168 = pi17  & n17166;
  assign n17169 = ~n17167 & ~n17168;
  assign n17170 = n16772 & ~n16774;
  assign n17171 = ~n16775 & ~n17170;
  assign n17172 = ~n17169 & n17171;
  assign n17173 = n6608 & n12262;
  assign n17174 = n6356 & n12265;
  assign n17175 = n6140 & n12268;
  assign n17176 = n6134 & n14691;
  assign n17177 = ~n17174 & ~n17175;
  assign n17178 = ~n17173 & n17177;
  assign n17179 = ~n17176 & n17178;
  assign n17180 = pi17  & n17179;
  assign n17181 = ~pi17  & ~n17179;
  assign n17182 = ~n17180 & ~n17181;
  assign n17183 = n16768 & ~n16770;
  assign n17184 = ~n16771 & ~n17183;
  assign n17185 = ~n17182 & n17184;
  assign n17186 = n6608 & n12265;
  assign n17187 = n6356 & n12268;
  assign n17188 = n6140 & n12271;
  assign n17189 = n6134 & n14728;
  assign n17190 = ~n17187 & ~n17188;
  assign n17191 = ~n17186 & n17190;
  assign n17192 = ~n17189 & n17191;
  assign n17193 = ~pi17  & ~n17192;
  assign n17194 = pi17  & n17192;
  assign n17195 = ~n17193 & ~n17194;
  assign n17196 = pi20  & ~n16748;
  assign n17197 = n16755 & ~n17196;
  assign n17198 = ~n16755 & n17196;
  assign n17199 = ~n17197 & ~n17198;
  assign n17200 = ~n17195 & n17199;
  assign n17201 = n6608 & n12268;
  assign n17202 = n6356 & n12271;
  assign n17203 = n6140 & n12274;
  assign n17204 = n6134 & n14771;
  assign n17205 = ~n17202 & ~n17203;
  assign n17206 = ~n17201 & n17205;
  assign n17207 = ~n17204 & n17206;
  assign n17208 = pi17  & n17207;
  assign n17209 = ~pi17  & ~n17207;
  assign n17210 = ~n17208 & ~n17209;
  assign n17211 = n16742 & ~n16747;
  assign n17212 = ~n16748 & ~n17211;
  assign n17213 = ~n17210 & n17212;
  assign n17214 = n6130 & n12281;
  assign n17215 = pi17  & n17214;
  assign n17216 = n6608 & n12279;
  assign n17217 = n6356 & n12281;
  assign n17218 = n6134 & ~n14833;
  assign n17219 = ~n17216 & ~n17217;
  assign n17220 = ~n17218 & n17219;
  assign n17221 = ~n17215 & n17220;
  assign n17222 = n6608 & n12274;
  assign n17223 = n6356 & n12279;
  assign n17224 = n6140 & n12281;
  assign n17225 = n6134 & ~n14876;
  assign n17226 = ~n17223 & ~n17224;
  assign n17227 = ~n17222 & n17226;
  assign n17228 = ~n17225 & n17227;
  assign n17229 = pi17  & n17221;
  assign n17230 = n17228 & n17229;
  assign n17231 = n16741 & n17230;
  assign n17232 = n6608 & n12271;
  assign n17233 = n6356 & n12274;
  assign n17234 = n6140 & n12279;
  assign n17235 = n6134 & n14795;
  assign n17236 = ~n17233 & ~n17234;
  assign n17237 = ~n17232 & n17236;
  assign n17238 = ~n17235 & n17237;
  assign n17239 = pi17  & n17238;
  assign n17240 = ~pi17  & ~n17238;
  assign n17241 = ~n17239 & ~n17240;
  assign n17242 = ~n16741 & ~n17230;
  assign n17243 = ~n17231 & ~n17242;
  assign n17244 = ~n17241 & n17243;
  assign n17245 = ~n17231 & ~n17244;
  assign n17246 = n17210 & ~n17212;
  assign n17247 = ~n17213 & ~n17246;
  assign n17248 = ~n17245 & n17247;
  assign n17249 = ~n17213 & ~n17248;
  assign n17250 = n17195 & ~n17199;
  assign n17251 = ~n17200 & ~n17250;
  assign n17252 = ~n17249 & n17251;
  assign n17253 = ~n17200 & ~n17252;
  assign n17254 = n17182 & ~n17184;
  assign n17255 = ~n17185 & ~n17254;
  assign n17256 = ~n17253 & n17255;
  assign n17257 = ~n17185 & ~n17256;
  assign n17258 = n17169 & ~n17171;
  assign n17259 = ~n17172 & ~n17258;
  assign n17260 = ~n17257 & n17259;
  assign n17261 = ~n17172 & ~n17260;
  assign n17262 = ~n17148 & n17158;
  assign n17263 = ~n17159 & ~n17262;
  assign n17264 = ~n17261 & n17263;
  assign n17265 = ~n17159 & ~n17264;
  assign n17266 = ~n17135 & n17145;
  assign n17267 = ~n17146 & ~n17266;
  assign n17268 = ~n17265 & n17267;
  assign n17269 = ~n17146 & ~n17268;
  assign n17270 = ~n17122 & n17132;
  assign n17271 = ~n17133 & ~n17270;
  assign n17272 = ~n17269 & n17271;
  assign n17273 = ~n17133 & ~n17272;
  assign n17274 = n17117 & ~n17119;
  assign n17275 = ~n17120 & ~n17274;
  assign n17276 = ~n17273 & n17275;
  assign n17277 = ~n17120 & ~n17276;
  assign n17278 = n17104 & ~n17106;
  assign n17279 = ~n17107 & ~n17278;
  assign n17280 = ~n17277 & n17279;
  assign n17281 = ~n17107 & ~n17280;
  assign n17282 = n17091 & ~n17093;
  assign n17283 = ~n17094 & ~n17282;
  assign n17284 = ~n17281 & n17283;
  assign n17285 = ~n17094 & ~n17284;
  assign n17286 = ~n17070 & n17080;
  assign n17287 = ~n17081 & ~n17286;
  assign n17288 = ~n17285 & n17287;
  assign n17289 = ~n17081 & ~n17288;
  assign n17290 = ~n17057 & n17067;
  assign n17291 = ~n17068 & ~n17290;
  assign n17292 = ~n17289 & n17291;
  assign n17293 = ~n17068 & ~n17292;
  assign n17294 = n17052 & ~n17054;
  assign n17295 = ~n17055 & ~n17294;
  assign n17296 = ~n17293 & n17295;
  assign n17297 = ~n17055 & ~n17296;
  assign n17298 = n17039 & ~n17041;
  assign n17299 = ~n17042 & ~n17298;
  assign n17300 = ~n17297 & n17299;
  assign n17301 = ~n17042 & ~n17300;
  assign n17302 = n17026 & ~n17028;
  assign n17303 = ~n17029 & ~n17302;
  assign n17304 = ~n17301 & n17303;
  assign n17305 = ~n17029 & ~n17304;
  assign n17306 = n17013 & ~n17015;
  assign n17307 = ~n17016 & ~n17306;
  assign n17308 = ~n17305 & n17307;
  assign n17309 = ~n17016 & ~n17308;
  assign n17310 = n17000 & ~n17002;
  assign n17311 = ~n17003 & ~n17310;
  assign n17312 = ~n17309 & n17311;
  assign n17313 = ~n17003 & ~n17312;
  assign n17314 = n16987 & ~n16989;
  assign n17315 = ~n16990 & ~n17314;
  assign n17316 = ~n17313 & n17315;
  assign n17317 = ~n16990 & ~n17316;
  assign n17318 = n16974 & ~n16976;
  assign n17319 = ~n16977 & ~n17318;
  assign n17320 = ~n17317 & n17319;
  assign n17321 = ~n16977 & ~n17320;
  assign n17322 = n16961 & ~n16963;
  assign n17323 = ~n16964 & ~n17322;
  assign n17324 = ~n17321 & n17323;
  assign n17325 = ~n16964 & ~n17324;
  assign n17326 = n16948 & ~n16950;
  assign n17327 = ~n16951 & ~n17326;
  assign n17328 = ~n17325 & n17327;
  assign n17329 = ~n16951 & ~n17328;
  assign n17330 = n16935 & ~n16937;
  assign n17331 = ~n16938 & ~n17330;
  assign n17332 = ~n17329 & n17331;
  assign n17333 = ~n16938 & ~n17332;
  assign n17334 = ~n16853 & n16863;
  assign n17335 = ~n16864 & ~n17334;
  assign n17336 = ~n17333 & n17335;
  assign n17337 = n17333 & ~n17335;
  assign n17338 = ~n17336 & ~n17337;
  assign n17339 = n7380 & n12193;
  assign n17340 = n7243 & n12196;
  assign n17341 = n6653 & n12199;
  assign n17342 = n6647 & n12594;
  assign n17343 = ~n17340 & ~n17341;
  assign n17344 = ~n17339 & n17343;
  assign n17345 = ~n17342 & n17344;
  assign n17346 = pi14  & n17345;
  assign n17347 = ~pi14  & ~n17345;
  assign n17348 = ~n17346 & ~n17347;
  assign n17349 = n17338 & ~n17348;
  assign n17350 = ~n17336 & ~n17349;
  assign n17351 = ~n16870 & n16880;
  assign n17352 = ~n16881 & ~n17351;
  assign n17353 = ~n17350 & n17352;
  assign n17354 = n17350 & ~n17352;
  assign n17355 = ~n17353 & ~n17354;
  assign n17356 = n8161 & n12181;
  assign n17357 = n7847 & n12184;
  assign n17358 = n7554 & n12187;
  assign n17359 = n7548 & n12608;
  assign n17360 = ~n17357 & ~n17358;
  assign n17361 = ~n17356 & n17360;
  assign n17362 = ~n17359 & n17361;
  assign n17363 = pi11  & n17362;
  assign n17364 = ~pi11  & ~n17362;
  assign n17365 = ~n17363 & ~n17364;
  assign n17366 = n17355 & ~n17365;
  assign n17367 = ~n17353 & ~n17366;
  assign n17368 = ~n16887 & n16897;
  assign n17369 = ~n16898 & ~n17368;
  assign n17370 = ~n17367 & n17369;
  assign n17371 = n17367 & ~n17369;
  assign n17372 = ~n17370 & ~n17371;
  assign n17373 = n9355 & n12172;
  assign n17374 = n8939 & n12168;
  assign n17375 = n8206 & n12175;
  assign n17376 = n8200 & n12939;
  assign n17377 = ~n17374 & ~n17375;
  assign n17378 = ~n17373 & n17377;
  assign n17379 = ~n17376 & n17378;
  assign n17380 = pi8  & n17379;
  assign n17381 = ~pi8  & ~n17379;
  assign n17382 = ~n17380 & ~n17381;
  assign n17383 = n17372 & ~n17382;
  assign n17384 = ~n17370 & ~n17383;
  assign n17385 = n9355 & n12166;
  assign n17386 = n8939 & n12172;
  assign n17387 = n8206 & n12168;
  assign n17388 = n8200 & n13106;
  assign n17389 = ~n17385 & ~n17387;
  assign n17390 = ~n17386 & n17389;
  assign n17391 = ~n17388 & n17390;
  assign n17392 = pi8  & n17391;
  assign n17393 = ~pi8  & ~n17391;
  assign n17394 = ~n17392 & ~n17393;
  assign n17395 = ~n17384 & ~n17394;
  assign n17396 = n16899 & ~n16901;
  assign n17397 = ~n16902 & ~n17396;
  assign n17398 = n17384 & n17394;
  assign n17399 = ~n17395 & ~n17398;
  assign n17400 = n17397 & n17399;
  assign n17401 = ~n17395 & ~n17400;
  assign n17402 = ~n16908 & n16918;
  assign n17403 = ~n16919 & ~n17402;
  assign n17404 = ~n17401 & n17403;
  assign n17405 = n17329 & ~n17331;
  assign n17406 = ~n17332 & ~n17405;
  assign n17407 = n7380 & n12196;
  assign n17408 = n7243 & n12199;
  assign n17409 = n6653 & n12202;
  assign n17410 = n6647 & n12578;
  assign n17411 = ~n17408 & ~n17409;
  assign n17412 = ~n17407 & n17411;
  assign n17413 = ~n17410 & n17412;
  assign n17414 = pi14  & n17413;
  assign n17415 = ~pi14  & ~n17413;
  assign n17416 = ~n17414 & ~n17415;
  assign n17417 = n17406 & ~n17416;
  assign n17418 = n17325 & ~n17327;
  assign n17419 = ~n17328 & ~n17418;
  assign n17420 = n7380 & n12199;
  assign n17421 = n7243 & n12202;
  assign n17422 = n6653 & n12205;
  assign n17423 = n6647 & n12683;
  assign n17424 = ~n17421 & ~n17422;
  assign n17425 = ~n17420 & n17424;
  assign n17426 = ~n17423 & n17425;
  assign n17427 = pi14  & n17426;
  assign n17428 = ~pi14  & ~n17426;
  assign n17429 = ~n17427 & ~n17428;
  assign n17430 = n17419 & ~n17429;
  assign n17431 = n17321 & ~n17323;
  assign n17432 = ~n17324 & ~n17431;
  assign n17433 = n7380 & n12202;
  assign n17434 = n7243 & n12205;
  assign n17435 = n6653 & n12208;
  assign n17436 = n6647 & n12701;
  assign n17437 = ~n17434 & ~n17435;
  assign n17438 = ~n17433 & n17437;
  assign n17439 = ~n17436 & n17438;
  assign n17440 = pi14  & n17439;
  assign n17441 = ~pi14  & ~n17439;
  assign n17442 = ~n17440 & ~n17441;
  assign n17443 = n17432 & ~n17442;
  assign n17444 = n17317 & ~n17319;
  assign n17445 = ~n17320 & ~n17444;
  assign n17446 = n7380 & n12205;
  assign n17447 = n7243 & n12208;
  assign n17448 = n6653 & n12211;
  assign n17449 = n6647 & n13031;
  assign n17450 = ~n17447 & ~n17448;
  assign n17451 = ~n17446 & n17450;
  assign n17452 = ~n17449 & n17451;
  assign n17453 = pi14  & n17452;
  assign n17454 = ~pi14  & ~n17452;
  assign n17455 = ~n17453 & ~n17454;
  assign n17456 = n17445 & ~n17455;
  assign n17457 = n17313 & ~n17315;
  assign n17458 = ~n17316 & ~n17457;
  assign n17459 = n7380 & n12208;
  assign n17460 = n7243 & n12211;
  assign n17461 = n6653 & n12214;
  assign n17462 = n6647 & n12804;
  assign n17463 = ~n17460 & ~n17461;
  assign n17464 = ~n17459 & n17463;
  assign n17465 = ~n17462 & n17464;
  assign n17466 = pi14  & n17465;
  assign n17467 = ~pi14  & ~n17465;
  assign n17468 = ~n17466 & ~n17467;
  assign n17469 = n17458 & ~n17468;
  assign n17470 = n17309 & ~n17311;
  assign n17471 = ~n17312 & ~n17470;
  assign n17472 = n7380 & n12211;
  assign n17473 = n7243 & n12214;
  assign n17474 = n6653 & n12217;
  assign n17475 = n6647 & n13203;
  assign n17476 = ~n17473 & ~n17474;
  assign n17477 = ~n17472 & n17476;
  assign n17478 = ~n17475 & n17477;
  assign n17479 = pi14  & n17478;
  assign n17480 = ~pi14  & ~n17478;
  assign n17481 = ~n17479 & ~n17480;
  assign n17482 = n17471 & ~n17481;
  assign n17483 = n17305 & ~n17307;
  assign n17484 = ~n17308 & ~n17483;
  assign n17485 = n7380 & n12214;
  assign n17486 = n7243 & n12217;
  assign n17487 = n6653 & n12220;
  assign n17488 = n6647 & n13187;
  assign n17489 = ~n17486 & ~n17487;
  assign n17490 = ~n17485 & n17489;
  assign n17491 = ~n17488 & n17490;
  assign n17492 = pi14  & n17491;
  assign n17493 = ~pi14  & ~n17491;
  assign n17494 = ~n17492 & ~n17493;
  assign n17495 = n17484 & ~n17494;
  assign n17496 = n17301 & ~n17303;
  assign n17497 = ~n17304 & ~n17496;
  assign n17498 = n7380 & n12217;
  assign n17499 = n7243 & n12220;
  assign n17500 = n6653 & n12223;
  assign n17501 = n6647 & n13374;
  assign n17502 = ~n17499 & ~n17500;
  assign n17503 = ~n17498 & n17502;
  assign n17504 = ~n17501 & n17503;
  assign n17505 = pi14  & n17504;
  assign n17506 = ~pi14  & ~n17504;
  assign n17507 = ~n17505 & ~n17506;
  assign n17508 = n17497 & ~n17507;
  assign n17509 = n17297 & ~n17299;
  assign n17510 = ~n17300 & ~n17509;
  assign n17511 = n7380 & n12220;
  assign n17512 = n7243 & n12223;
  assign n17513 = n6653 & n12226;
  assign n17514 = n6647 & n13392;
  assign n17515 = ~n17512 & ~n17513;
  assign n17516 = ~n17511 & n17515;
  assign n17517 = ~n17514 & n17516;
  assign n17518 = pi14  & n17517;
  assign n17519 = ~pi14  & ~n17517;
  assign n17520 = ~n17518 & ~n17519;
  assign n17521 = n17510 & ~n17520;
  assign n17522 = n17293 & ~n17295;
  assign n17523 = ~n17296 & ~n17522;
  assign n17524 = n7380 & n12223;
  assign n17525 = n7243 & n12226;
  assign n17526 = n6653 & n12229;
  assign n17527 = n6647 & n13745;
  assign n17528 = ~n17525 & ~n17526;
  assign n17529 = ~n17524 & n17528;
  assign n17530 = ~n17527 & n17529;
  assign n17531 = pi14  & n17530;
  assign n17532 = ~pi14  & ~n17530;
  assign n17533 = ~n17531 & ~n17532;
  assign n17534 = n17523 & ~n17533;
  assign n17535 = n7380 & n12226;
  assign n17536 = n7243 & n12229;
  assign n17537 = n6653 & n12232;
  assign n17538 = n6647 & n13530;
  assign n17539 = ~n17536 & ~n17537;
  assign n17540 = ~n17535 & n17539;
  assign n17541 = ~n17538 & n17540;
  assign n17542 = ~pi14  & ~n17541;
  assign n17543 = pi14  & n17541;
  assign n17544 = ~n17542 & ~n17543;
  assign n17545 = n17289 & ~n17291;
  assign n17546 = ~n17292 & ~n17545;
  assign n17547 = ~n17544 & n17546;
  assign n17548 = n7380 & n12229;
  assign n17549 = n7243 & n12232;
  assign n17550 = n6653 & n12235;
  assign n17551 = n6647 & n13979;
  assign n17552 = ~n17549 & ~n17550;
  assign n17553 = ~n17548 & n17552;
  assign n17554 = ~n17551 & n17553;
  assign n17555 = ~pi14  & ~n17554;
  assign n17556 = pi14  & n17554;
  assign n17557 = ~n17555 & ~n17556;
  assign n17558 = n17285 & ~n17287;
  assign n17559 = ~n17288 & ~n17558;
  assign n17560 = ~n17557 & n17559;
  assign n17561 = n17281 & ~n17283;
  assign n17562 = ~n17284 & ~n17561;
  assign n17563 = n7380 & n12232;
  assign n17564 = n7243 & n12235;
  assign n17565 = n6653 & n12238;
  assign n17566 = n6647 & n14116;
  assign n17567 = ~n17564 & ~n17565;
  assign n17568 = ~n17563 & n17567;
  assign n17569 = ~n17566 & n17568;
  assign n17570 = pi14  & n17569;
  assign n17571 = ~pi14  & ~n17569;
  assign n17572 = ~n17570 & ~n17571;
  assign n17573 = n17562 & ~n17572;
  assign n17574 = n17277 & ~n17279;
  assign n17575 = ~n17280 & ~n17574;
  assign n17576 = n7380 & n12235;
  assign n17577 = n7243 & n12238;
  assign n17578 = n6653 & n12241;
  assign n17579 = n6647 & n13959;
  assign n17580 = ~n17577 & ~n17578;
  assign n17581 = ~n17576 & n17580;
  assign n17582 = ~n17579 & n17581;
  assign n17583 = pi14  & n17582;
  assign n17584 = ~pi14  & ~n17582;
  assign n17585 = ~n17583 & ~n17584;
  assign n17586 = n17575 & ~n17585;
  assign n17587 = n17273 & ~n17275;
  assign n17588 = ~n17276 & ~n17587;
  assign n17589 = n7380 & n12238;
  assign n17590 = n7243 & n12241;
  assign n17591 = n6653 & n12244;
  assign n17592 = n6647 & n14229;
  assign n17593 = ~n17590 & ~n17591;
  assign n17594 = ~n17589 & n17593;
  assign n17595 = ~n17592 & n17594;
  assign n17596 = pi14  & n17595;
  assign n17597 = ~pi14  & ~n17595;
  assign n17598 = ~n17596 & ~n17597;
  assign n17599 = n17588 & ~n17598;
  assign n17600 = n7380 & n12241;
  assign n17601 = n7243 & n12244;
  assign n17602 = n6653 & n12247;
  assign n17603 = n6647 & n14515;
  assign n17604 = ~n17601 & ~n17602;
  assign n17605 = ~n17600 & n17604;
  assign n17606 = ~n17603 & n17605;
  assign n17607 = ~pi14  & ~n17606;
  assign n17608 = pi14  & n17606;
  assign n17609 = ~n17607 & ~n17608;
  assign n17610 = n17269 & ~n17271;
  assign n17611 = ~n17272 & ~n17610;
  assign n17612 = ~n17609 & n17611;
  assign n17613 = n7380 & n12244;
  assign n17614 = n7243 & n12247;
  assign n17615 = n6653 & n12250;
  assign n17616 = n6647 & n14527;
  assign n17617 = ~n17614 & ~n17615;
  assign n17618 = ~n17613 & n17617;
  assign n17619 = ~n17616 & n17618;
  assign n17620 = ~pi14  & ~n17619;
  assign n17621 = pi14  & n17619;
  assign n17622 = ~n17620 & ~n17621;
  assign n17623 = n17265 & ~n17267;
  assign n17624 = ~n17268 & ~n17623;
  assign n17625 = ~n17622 & n17624;
  assign n17626 = n7380 & n12247;
  assign n17627 = n7243 & n12250;
  assign n17628 = n6653 & n12253;
  assign n17629 = n6647 & n14207;
  assign n17630 = ~n17627 & ~n17628;
  assign n17631 = ~n17626 & n17630;
  assign n17632 = ~n17629 & n17631;
  assign n17633 = ~pi14  & ~n17632;
  assign n17634 = pi14  & n17632;
  assign n17635 = ~n17633 & ~n17634;
  assign n17636 = n17261 & ~n17263;
  assign n17637 = ~n17264 & ~n17636;
  assign n17638 = ~n17635 & n17637;
  assign n17639 = n17257 & ~n17259;
  assign n17640 = ~n17260 & ~n17639;
  assign n17641 = n7380 & n12250;
  assign n17642 = n7243 & n12253;
  assign n17643 = n6653 & n12256;
  assign n17644 = n6647 & n14559;
  assign n17645 = ~n17642 & ~n17643;
  assign n17646 = ~n17641 & n17645;
  assign n17647 = ~n17644 & n17646;
  assign n17648 = pi14  & n17647;
  assign n17649 = ~pi14  & ~n17647;
  assign n17650 = ~n17648 & ~n17649;
  assign n17651 = n17640 & ~n17650;
  assign n17652 = n17253 & ~n17255;
  assign n17653 = ~n17256 & ~n17652;
  assign n17654 = n7380 & n12253;
  assign n17655 = n7243 & n12256;
  assign n17656 = n6653 & n12259;
  assign n17657 = n6647 & n14584;
  assign n17658 = ~n17655 & ~n17656;
  assign n17659 = ~n17654 & n17658;
  assign n17660 = ~n17657 & n17659;
  assign n17661 = pi14  & n17660;
  assign n17662 = ~pi14  & ~n17660;
  assign n17663 = ~n17661 & ~n17662;
  assign n17664 = n17653 & ~n17663;
  assign n17665 = n17249 & ~n17251;
  assign n17666 = ~n17252 & ~n17665;
  assign n17667 = n7380 & n12256;
  assign n17668 = n7243 & n12259;
  assign n17669 = n6653 & n12262;
  assign n17670 = n6647 & n14608;
  assign n17671 = ~n17668 & ~n17669;
  assign n17672 = ~n17667 & n17671;
  assign n17673 = ~n17670 & n17672;
  assign n17674 = pi14  & n17673;
  assign n17675 = ~pi14  & ~n17673;
  assign n17676 = ~n17674 & ~n17675;
  assign n17677 = n17666 & ~n17676;
  assign n17678 = n7380 & n12259;
  assign n17679 = n7243 & n12262;
  assign n17680 = n6653 & n12265;
  assign n17681 = n6647 & n14637;
  assign n17682 = ~n17679 & ~n17680;
  assign n17683 = ~n17678 & n17682;
  assign n17684 = ~n17681 & n17683;
  assign n17685 = ~pi14  & ~n17684;
  assign n17686 = pi14  & n17684;
  assign n17687 = ~n17685 & ~n17686;
  assign n17688 = n17245 & ~n17247;
  assign n17689 = ~n17248 & ~n17688;
  assign n17690 = ~n17687 & n17689;
  assign n17691 = n7380 & n12262;
  assign n17692 = n7243 & n12265;
  assign n17693 = n6653 & n12268;
  assign n17694 = n6647 & n14691;
  assign n17695 = ~n17692 & ~n17693;
  assign n17696 = ~n17691 & n17695;
  assign n17697 = ~n17694 & n17696;
  assign n17698 = pi14  & n17697;
  assign n17699 = ~pi14  & ~n17697;
  assign n17700 = ~n17698 & ~n17699;
  assign n17701 = n17241 & ~n17243;
  assign n17702 = ~n17244 & ~n17701;
  assign n17703 = ~n17700 & n17702;
  assign n17704 = n7380 & n12265;
  assign n17705 = n7243 & n12268;
  assign n17706 = n6653 & n12271;
  assign n17707 = n6647 & n14728;
  assign n17708 = ~n17705 & ~n17706;
  assign n17709 = ~n17704 & n17708;
  assign n17710 = ~n17707 & n17709;
  assign n17711 = ~pi14  & ~n17710;
  assign n17712 = pi14  & n17710;
  assign n17713 = ~n17711 & ~n17712;
  assign n17714 = pi17  & ~n17221;
  assign n17715 = n17228 & ~n17714;
  assign n17716 = ~n17228 & n17714;
  assign n17717 = ~n17715 & ~n17716;
  assign n17718 = ~n17713 & n17717;
  assign n17719 = n7380 & n12268;
  assign n17720 = n7243 & n12271;
  assign n17721 = n6653 & n12274;
  assign n17722 = n6647 & n14771;
  assign n17723 = ~n17720 & ~n17721;
  assign n17724 = ~n17719 & n17723;
  assign n17725 = ~n17722 & n17724;
  assign n17726 = pi14  & n17725;
  assign n17727 = ~pi14  & ~n17725;
  assign n17728 = ~n17726 & ~n17727;
  assign n17729 = n17215 & ~n17220;
  assign n17730 = ~n17221 & ~n17729;
  assign n17731 = ~n17728 & n17730;
  assign n17732 = n6643 & n12281;
  assign n17733 = pi14  & n17732;
  assign n17734 = n7380 & n12279;
  assign n17735 = n7243 & n12281;
  assign n17736 = n6647 & ~n14833;
  assign n17737 = ~n17734 & ~n17735;
  assign n17738 = ~n17736 & n17737;
  assign n17739 = ~n17733 & n17738;
  assign n17740 = n7380 & n12274;
  assign n17741 = n7243 & n12279;
  assign n17742 = n6653 & n12281;
  assign n17743 = n6647 & ~n14876;
  assign n17744 = ~n17741 & ~n17742;
  assign n17745 = ~n17740 & n17744;
  assign n17746 = ~n17743 & n17745;
  assign n17747 = pi14  & n17739;
  assign n17748 = n17746 & n17747;
  assign n17749 = n17214 & n17748;
  assign n17750 = n7380 & n12271;
  assign n17751 = n7243 & n12274;
  assign n17752 = n6653 & n12279;
  assign n17753 = n6647 & n14795;
  assign n17754 = ~n17751 & ~n17752;
  assign n17755 = ~n17750 & n17754;
  assign n17756 = ~n17753 & n17755;
  assign n17757 = pi14  & n17756;
  assign n17758 = ~pi14  & ~n17756;
  assign n17759 = ~n17757 & ~n17758;
  assign n17760 = ~n17214 & ~n17748;
  assign n17761 = ~n17749 & ~n17760;
  assign n17762 = ~n17759 & n17761;
  assign n17763 = ~n17749 & ~n17762;
  assign n17764 = n17728 & ~n17730;
  assign n17765 = ~n17731 & ~n17764;
  assign n17766 = ~n17763 & n17765;
  assign n17767 = ~n17731 & ~n17766;
  assign n17768 = n17713 & ~n17717;
  assign n17769 = ~n17718 & ~n17768;
  assign n17770 = ~n17767 & n17769;
  assign n17771 = ~n17718 & ~n17770;
  assign n17772 = n17700 & ~n17702;
  assign n17773 = ~n17703 & ~n17772;
  assign n17774 = ~n17771 & n17773;
  assign n17775 = ~n17703 & ~n17774;
  assign n17776 = n17687 & ~n17689;
  assign n17777 = ~n17690 & ~n17776;
  assign n17778 = ~n17775 & n17777;
  assign n17779 = ~n17690 & ~n17778;
  assign n17780 = ~n17666 & n17676;
  assign n17781 = ~n17677 & ~n17780;
  assign n17782 = ~n17779 & n17781;
  assign n17783 = ~n17677 & ~n17782;
  assign n17784 = ~n17653 & n17663;
  assign n17785 = ~n17664 & ~n17784;
  assign n17786 = ~n17783 & n17785;
  assign n17787 = ~n17664 & ~n17786;
  assign n17788 = ~n17640 & n17650;
  assign n17789 = ~n17651 & ~n17788;
  assign n17790 = ~n17787 & n17789;
  assign n17791 = ~n17651 & ~n17790;
  assign n17792 = n17635 & ~n17637;
  assign n17793 = ~n17638 & ~n17792;
  assign n17794 = ~n17791 & n17793;
  assign n17795 = ~n17638 & ~n17794;
  assign n17796 = n17622 & ~n17624;
  assign n17797 = ~n17625 & ~n17796;
  assign n17798 = ~n17795 & n17797;
  assign n17799 = ~n17625 & ~n17798;
  assign n17800 = n17609 & ~n17611;
  assign n17801 = ~n17612 & ~n17800;
  assign n17802 = ~n17799 & n17801;
  assign n17803 = ~n17612 & ~n17802;
  assign n17804 = ~n17588 & n17598;
  assign n17805 = ~n17599 & ~n17804;
  assign n17806 = ~n17803 & n17805;
  assign n17807 = ~n17599 & ~n17806;
  assign n17808 = ~n17575 & n17585;
  assign n17809 = ~n17586 & ~n17808;
  assign n17810 = ~n17807 & n17809;
  assign n17811 = ~n17586 & ~n17810;
  assign n17812 = ~n17562 & n17572;
  assign n17813 = ~n17573 & ~n17812;
  assign n17814 = ~n17811 & n17813;
  assign n17815 = ~n17573 & ~n17814;
  assign n17816 = n17557 & ~n17559;
  assign n17817 = ~n17560 & ~n17816;
  assign n17818 = ~n17815 & n17817;
  assign n17819 = ~n17560 & ~n17818;
  assign n17820 = n17544 & ~n17546;
  assign n17821 = ~n17547 & ~n17820;
  assign n17822 = ~n17819 & n17821;
  assign n17823 = ~n17547 & ~n17822;
  assign n17824 = ~n17523 & n17533;
  assign n17825 = ~n17534 & ~n17824;
  assign n17826 = ~n17823 & n17825;
  assign n17827 = ~n17534 & ~n17826;
  assign n17828 = ~n17510 & n17520;
  assign n17829 = ~n17521 & ~n17828;
  assign n17830 = ~n17827 & n17829;
  assign n17831 = ~n17521 & ~n17830;
  assign n17832 = ~n17497 & n17507;
  assign n17833 = ~n17508 & ~n17832;
  assign n17834 = ~n17831 & n17833;
  assign n17835 = ~n17508 & ~n17834;
  assign n17836 = ~n17484 & n17494;
  assign n17837 = ~n17495 & ~n17836;
  assign n17838 = ~n17835 & n17837;
  assign n17839 = ~n17495 & ~n17838;
  assign n17840 = ~n17471 & n17481;
  assign n17841 = ~n17482 & ~n17840;
  assign n17842 = ~n17839 & n17841;
  assign n17843 = ~n17482 & ~n17842;
  assign n17844 = ~n17458 & n17468;
  assign n17845 = ~n17469 & ~n17844;
  assign n17846 = ~n17843 & n17845;
  assign n17847 = ~n17469 & ~n17846;
  assign n17848 = ~n17445 & n17455;
  assign n17849 = ~n17456 & ~n17848;
  assign n17850 = ~n17847 & n17849;
  assign n17851 = ~n17456 & ~n17850;
  assign n17852 = ~n17432 & n17442;
  assign n17853 = ~n17443 & ~n17852;
  assign n17854 = ~n17851 & n17853;
  assign n17855 = ~n17443 & ~n17854;
  assign n17856 = ~n17419 & n17429;
  assign n17857 = ~n17430 & ~n17856;
  assign n17858 = ~n17855 & n17857;
  assign n17859 = ~n17430 & ~n17858;
  assign n17860 = ~n17406 & n17416;
  assign n17861 = ~n17417 & ~n17860;
  assign n17862 = ~n17859 & n17861;
  assign n17863 = ~n17417 & ~n17862;
  assign n17864 = ~n17338 & n17348;
  assign n17865 = ~n17349 & ~n17864;
  assign n17866 = ~n17863 & n17865;
  assign n17867 = n17863 & ~n17865;
  assign n17868 = ~n17866 & ~n17867;
  assign n17869 = n8161 & n12184;
  assign n17870 = n7847 & n12187;
  assign n17871 = n7554 & n12190;
  assign n17872 = n7548 & n12845;
  assign n17873 = ~n17870 & ~n17871;
  assign n17874 = ~n17869 & n17873;
  assign n17875 = ~n17872 & n17874;
  assign n17876 = pi11  & n17875;
  assign n17877 = ~pi11  & ~n17875;
  assign n17878 = ~n17876 & ~n17877;
  assign n17879 = n17868 & ~n17878;
  assign n17880 = ~n17866 & ~n17879;
  assign n17881 = ~n17355 & n17365;
  assign n17882 = ~n17366 & ~n17881;
  assign n17883 = ~n17880 & n17882;
  assign n17884 = n17880 & ~n17882;
  assign n17885 = ~n17883 & ~n17884;
  assign n17886 = n9355 & n12168;
  assign n17887 = n8939 & n12175;
  assign n17888 = n8206 & n12178;
  assign n17889 = n8200 & n12862;
  assign n17890 = ~n17887 & ~n17888;
  assign n17891 = ~n17886 & n17890;
  assign n17892 = ~n17889 & n17891;
  assign n17893 = pi8  & n17892;
  assign n17894 = ~pi8  & ~n17892;
  assign n17895 = ~n17893 & ~n17894;
  assign n17896 = n17885 & ~n17895;
  assign n17897 = ~n17883 & ~n17896;
  assign n17898 = n9830 & ~n12424;
  assign n17899 = n9835 & ~n12165;
  assign n17900 = n13942 & ~n17899;
  assign n17901 = ~n12163 & ~n17900;
  assign n17902 = ~n17898 & ~n17901;
  assign n17903 = pi5  & n17902;
  assign n17904 = ~pi5  & ~n17902;
  assign n17905 = ~n17903 & ~n17904;
  assign n17906 = ~n17897 & ~n17905;
  assign n17907 = n17897 & n17905;
  assign n17908 = ~n17906 & ~n17907;
  assign n17909 = ~n17372 & n17382;
  assign n17910 = ~n17383 & ~n17909;
  assign n17911 = n17908 & n17910;
  assign n17912 = ~n17906 & ~n17911;
  assign n17913 = ~n17397 & ~n17399;
  assign n17914 = ~n17400 & ~n17913;
  assign n17915 = ~n17912 & n17914;
  assign n17916 = n8161 & n12187;
  assign n17917 = n7847 & n12190;
  assign n17918 = n7554 & n12193;
  assign n17919 = n7548 & n12921;
  assign n17920 = ~n17917 & ~n17918;
  assign n17921 = ~n17916 & n17920;
  assign n17922 = ~n17919 & n17921;
  assign n17923 = ~pi11  & ~n17922;
  assign n17924 = pi11  & n17922;
  assign n17925 = ~n17923 & ~n17924;
  assign n17926 = n17859 & ~n17861;
  assign n17927 = ~n17862 & ~n17926;
  assign n17928 = ~n17925 & n17927;
  assign n17929 = n8161 & n12190;
  assign n17930 = n7847 & n12193;
  assign n17931 = n7554 & n12196;
  assign n17932 = n7548 & n12530;
  assign n17933 = ~n17930 & ~n17931;
  assign n17934 = ~n17929 & n17933;
  assign n17935 = ~n17932 & n17934;
  assign n17936 = ~pi11  & ~n17935;
  assign n17937 = pi11  & n17935;
  assign n17938 = ~n17936 & ~n17937;
  assign n17939 = n17855 & ~n17857;
  assign n17940 = ~n17858 & ~n17939;
  assign n17941 = ~n17938 & n17940;
  assign n17942 = n8161 & n12193;
  assign n17943 = n7847 & n12196;
  assign n17944 = n7554 & n12199;
  assign n17945 = n7548 & n12594;
  assign n17946 = ~n17943 & ~n17944;
  assign n17947 = ~n17942 & n17946;
  assign n17948 = ~n17945 & n17947;
  assign n17949 = ~pi11  & ~n17948;
  assign n17950 = pi11  & n17948;
  assign n17951 = ~n17949 & ~n17950;
  assign n17952 = n17851 & ~n17853;
  assign n17953 = ~n17854 & ~n17952;
  assign n17954 = ~n17951 & n17953;
  assign n17955 = n8161 & n12196;
  assign n17956 = n7847 & n12199;
  assign n17957 = n7554 & n12202;
  assign n17958 = n7548 & n12578;
  assign n17959 = ~n17956 & ~n17957;
  assign n17960 = ~n17955 & n17959;
  assign n17961 = ~n17958 & n17960;
  assign n17962 = ~pi11  & ~n17961;
  assign n17963 = pi11  & n17961;
  assign n17964 = ~n17962 & ~n17963;
  assign n17965 = n17847 & ~n17849;
  assign n17966 = ~n17850 & ~n17965;
  assign n17967 = ~n17964 & n17966;
  assign n17968 = n8161 & n12199;
  assign n17969 = n7847 & n12202;
  assign n17970 = n7554 & n12205;
  assign n17971 = n7548 & n12683;
  assign n17972 = ~n17969 & ~n17970;
  assign n17973 = ~n17968 & n17972;
  assign n17974 = ~n17971 & n17973;
  assign n17975 = ~pi11  & ~n17974;
  assign n17976 = pi11  & n17974;
  assign n17977 = ~n17975 & ~n17976;
  assign n17978 = n17843 & ~n17845;
  assign n17979 = ~n17846 & ~n17978;
  assign n17980 = ~n17977 & n17979;
  assign n17981 = n8161 & n12202;
  assign n17982 = n7847 & n12205;
  assign n17983 = n7554 & n12208;
  assign n17984 = n7548 & n12701;
  assign n17985 = ~n17982 & ~n17983;
  assign n17986 = ~n17981 & n17985;
  assign n17987 = ~n17984 & n17986;
  assign n17988 = ~pi11  & ~n17987;
  assign n17989 = pi11  & n17987;
  assign n17990 = ~n17988 & ~n17989;
  assign n17991 = n17839 & ~n17841;
  assign n17992 = ~n17842 & ~n17991;
  assign n17993 = ~n17990 & n17992;
  assign n17994 = n8161 & n12205;
  assign n17995 = n7847 & n12208;
  assign n17996 = n7554 & n12211;
  assign n17997 = n7548 & n13031;
  assign n17998 = ~n17995 & ~n17996;
  assign n17999 = ~n17994 & n17998;
  assign n18000 = ~n17997 & n17999;
  assign n18001 = ~pi11  & ~n18000;
  assign n18002 = pi11  & n18000;
  assign n18003 = ~n18001 & ~n18002;
  assign n18004 = n17835 & ~n17837;
  assign n18005 = ~n17838 & ~n18004;
  assign n18006 = ~n18003 & n18005;
  assign n18007 = n8161 & n12208;
  assign n18008 = n7847 & n12211;
  assign n18009 = n7554 & n12214;
  assign n18010 = n7548 & n12804;
  assign n18011 = ~n18008 & ~n18009;
  assign n18012 = ~n18007 & n18011;
  assign n18013 = ~n18010 & n18012;
  assign n18014 = ~pi11  & ~n18013;
  assign n18015 = pi11  & n18013;
  assign n18016 = ~n18014 & ~n18015;
  assign n18017 = n17831 & ~n17833;
  assign n18018 = ~n17834 & ~n18017;
  assign n18019 = ~n18016 & n18018;
  assign n18020 = n8161 & n12211;
  assign n18021 = n7847 & n12214;
  assign n18022 = n7554 & n12217;
  assign n18023 = n7548 & n13203;
  assign n18024 = ~n18021 & ~n18022;
  assign n18025 = ~n18020 & n18024;
  assign n18026 = ~n18023 & n18025;
  assign n18027 = ~pi11  & ~n18026;
  assign n18028 = pi11  & n18026;
  assign n18029 = ~n18027 & ~n18028;
  assign n18030 = n17827 & ~n17829;
  assign n18031 = ~n17830 & ~n18030;
  assign n18032 = ~n18029 & n18031;
  assign n18033 = n8161 & n12214;
  assign n18034 = n7847 & n12217;
  assign n18035 = n7554 & n12220;
  assign n18036 = n7548 & n13187;
  assign n18037 = ~n18034 & ~n18035;
  assign n18038 = ~n18033 & n18037;
  assign n18039 = ~n18036 & n18038;
  assign n18040 = ~pi11  & ~n18039;
  assign n18041 = pi11  & n18039;
  assign n18042 = ~n18040 & ~n18041;
  assign n18043 = n17823 & ~n17825;
  assign n18044 = ~n17826 & ~n18043;
  assign n18045 = ~n18042 & n18044;
  assign n18046 = n17819 & ~n17821;
  assign n18047 = ~n17822 & ~n18046;
  assign n18048 = n8161 & n12217;
  assign n18049 = n7847 & n12220;
  assign n18050 = n7554 & n12223;
  assign n18051 = n7548 & n13374;
  assign n18052 = ~n18049 & ~n18050;
  assign n18053 = ~n18048 & n18052;
  assign n18054 = ~n18051 & n18053;
  assign n18055 = pi11  & n18054;
  assign n18056 = ~pi11  & ~n18054;
  assign n18057 = ~n18055 & ~n18056;
  assign n18058 = n18047 & ~n18057;
  assign n18059 = n17815 & ~n17817;
  assign n18060 = ~n17818 & ~n18059;
  assign n18061 = n8161 & n12220;
  assign n18062 = n7847 & n12223;
  assign n18063 = n7554 & n12226;
  assign n18064 = n7548 & n13392;
  assign n18065 = ~n18062 & ~n18063;
  assign n18066 = ~n18061 & n18065;
  assign n18067 = ~n18064 & n18066;
  assign n18068 = pi11  & n18067;
  assign n18069 = ~pi11  & ~n18067;
  assign n18070 = ~n18068 & ~n18069;
  assign n18071 = n18060 & ~n18070;
  assign n18072 = n8161 & n12223;
  assign n18073 = n7847 & n12226;
  assign n18074 = n7554 & n12229;
  assign n18075 = n7548 & n13745;
  assign n18076 = ~n18073 & ~n18074;
  assign n18077 = ~n18072 & n18076;
  assign n18078 = ~n18075 & n18077;
  assign n18079 = ~pi11  & ~n18078;
  assign n18080 = pi11  & n18078;
  assign n18081 = ~n18079 & ~n18080;
  assign n18082 = n17811 & ~n17813;
  assign n18083 = ~n17814 & ~n18082;
  assign n18084 = ~n18081 & n18083;
  assign n18085 = n8161 & n12226;
  assign n18086 = n7847 & n12229;
  assign n18087 = n7554 & n12232;
  assign n18088 = n7548 & n13530;
  assign n18089 = ~n18086 & ~n18087;
  assign n18090 = ~n18085 & n18089;
  assign n18091 = ~n18088 & n18090;
  assign n18092 = ~pi11  & ~n18091;
  assign n18093 = pi11  & n18091;
  assign n18094 = ~n18092 & ~n18093;
  assign n18095 = n17807 & ~n17809;
  assign n18096 = ~n17810 & ~n18095;
  assign n18097 = ~n18094 & n18096;
  assign n18098 = n8161 & n12229;
  assign n18099 = n7847 & n12232;
  assign n18100 = n7554 & n12235;
  assign n18101 = n7548 & n13979;
  assign n18102 = ~n18099 & ~n18100;
  assign n18103 = ~n18098 & n18102;
  assign n18104 = ~n18101 & n18103;
  assign n18105 = ~pi11  & ~n18104;
  assign n18106 = pi11  & n18104;
  assign n18107 = ~n18105 & ~n18106;
  assign n18108 = n17803 & ~n17805;
  assign n18109 = ~n17806 & ~n18108;
  assign n18110 = ~n18107 & n18109;
  assign n18111 = n17799 & ~n17801;
  assign n18112 = ~n17802 & ~n18111;
  assign n18113 = n8161 & n12232;
  assign n18114 = n7847 & n12235;
  assign n18115 = n7554 & n12238;
  assign n18116 = n7548 & n14116;
  assign n18117 = ~n18114 & ~n18115;
  assign n18118 = ~n18113 & n18117;
  assign n18119 = ~n18116 & n18118;
  assign n18120 = pi11  & n18119;
  assign n18121 = ~pi11  & ~n18119;
  assign n18122 = ~n18120 & ~n18121;
  assign n18123 = n18112 & ~n18122;
  assign n18124 = n17795 & ~n17797;
  assign n18125 = ~n17798 & ~n18124;
  assign n18126 = n8161 & n12235;
  assign n18127 = n7847 & n12238;
  assign n18128 = n7554 & n12241;
  assign n18129 = n7548 & n13959;
  assign n18130 = ~n18127 & ~n18128;
  assign n18131 = ~n18126 & n18130;
  assign n18132 = ~n18129 & n18131;
  assign n18133 = pi11  & n18132;
  assign n18134 = ~pi11  & ~n18132;
  assign n18135 = ~n18133 & ~n18134;
  assign n18136 = n18125 & ~n18135;
  assign n18137 = n17791 & ~n17793;
  assign n18138 = ~n17794 & ~n18137;
  assign n18139 = n8161 & n12238;
  assign n18140 = n7847 & n12241;
  assign n18141 = n7554 & n12244;
  assign n18142 = n7548 & n14229;
  assign n18143 = ~n18140 & ~n18141;
  assign n18144 = ~n18139 & n18143;
  assign n18145 = ~n18142 & n18144;
  assign n18146 = pi11  & n18145;
  assign n18147 = ~pi11  & ~n18145;
  assign n18148 = ~n18146 & ~n18147;
  assign n18149 = n18138 & ~n18148;
  assign n18150 = n8161 & n12241;
  assign n18151 = n7847 & n12244;
  assign n18152 = n7554 & n12247;
  assign n18153 = n7548 & n14515;
  assign n18154 = ~n18151 & ~n18152;
  assign n18155 = ~n18150 & n18154;
  assign n18156 = ~n18153 & n18155;
  assign n18157 = ~pi11  & ~n18156;
  assign n18158 = pi11  & n18156;
  assign n18159 = ~n18157 & ~n18158;
  assign n18160 = n17787 & ~n17789;
  assign n18161 = ~n17790 & ~n18160;
  assign n18162 = ~n18159 & n18161;
  assign n18163 = n8161 & n12244;
  assign n18164 = n7847 & n12247;
  assign n18165 = n7554 & n12250;
  assign n18166 = n7548 & n14527;
  assign n18167 = ~n18164 & ~n18165;
  assign n18168 = ~n18163 & n18167;
  assign n18169 = ~n18166 & n18168;
  assign n18170 = ~pi11  & ~n18169;
  assign n18171 = pi11  & n18169;
  assign n18172 = ~n18170 & ~n18171;
  assign n18173 = n17783 & ~n17785;
  assign n18174 = ~n17786 & ~n18173;
  assign n18175 = ~n18172 & n18174;
  assign n18176 = n8161 & n12247;
  assign n18177 = n7847 & n12250;
  assign n18178 = n7554 & n12253;
  assign n18179 = n7548 & n14207;
  assign n18180 = ~n18177 & ~n18178;
  assign n18181 = ~n18176 & n18180;
  assign n18182 = ~n18179 & n18181;
  assign n18183 = ~pi11  & ~n18182;
  assign n18184 = pi11  & n18182;
  assign n18185 = ~n18183 & ~n18184;
  assign n18186 = n17779 & ~n17781;
  assign n18187 = ~n17782 & ~n18186;
  assign n18188 = ~n18185 & n18187;
  assign n18189 = n17775 & ~n17777;
  assign n18190 = ~n17778 & ~n18189;
  assign n18191 = n8161 & n12250;
  assign n18192 = n7847 & n12253;
  assign n18193 = n7554 & n12256;
  assign n18194 = n7548 & n14559;
  assign n18195 = ~n18192 & ~n18193;
  assign n18196 = ~n18191 & n18195;
  assign n18197 = ~n18194 & n18196;
  assign n18198 = pi11  & n18197;
  assign n18199 = ~pi11  & ~n18197;
  assign n18200 = ~n18198 & ~n18199;
  assign n18201 = n18190 & ~n18200;
  assign n18202 = n17771 & ~n17773;
  assign n18203 = ~n17774 & ~n18202;
  assign n18204 = n8161 & n12253;
  assign n18205 = n7847 & n12256;
  assign n18206 = n7554 & n12259;
  assign n18207 = n7548 & n14584;
  assign n18208 = ~n18205 & ~n18206;
  assign n18209 = ~n18204 & n18208;
  assign n18210 = ~n18207 & n18209;
  assign n18211 = pi11  & n18210;
  assign n18212 = ~pi11  & ~n18210;
  assign n18213 = ~n18211 & ~n18212;
  assign n18214 = n18203 & ~n18213;
  assign n18215 = n17767 & ~n17769;
  assign n18216 = ~n17770 & ~n18215;
  assign n18217 = n8161 & n12256;
  assign n18218 = n7847 & n12259;
  assign n18219 = n7554 & n12262;
  assign n18220 = n7548 & n14608;
  assign n18221 = ~n18218 & ~n18219;
  assign n18222 = ~n18217 & n18221;
  assign n18223 = ~n18220 & n18222;
  assign n18224 = pi11  & n18223;
  assign n18225 = ~pi11  & ~n18223;
  assign n18226 = ~n18224 & ~n18225;
  assign n18227 = n18216 & ~n18226;
  assign n18228 = n8161 & n12259;
  assign n18229 = n7847 & n12262;
  assign n18230 = n7554 & n12265;
  assign n18231 = n7548 & n14637;
  assign n18232 = ~n18229 & ~n18230;
  assign n18233 = ~n18228 & n18232;
  assign n18234 = ~n18231 & n18233;
  assign n18235 = ~pi11  & ~n18234;
  assign n18236 = pi11  & n18234;
  assign n18237 = ~n18235 & ~n18236;
  assign n18238 = n17763 & ~n17765;
  assign n18239 = ~n17766 & ~n18238;
  assign n18240 = ~n18237 & n18239;
  assign n18241 = n8161 & n12262;
  assign n18242 = n7847 & n12265;
  assign n18243 = n7554 & n12268;
  assign n18244 = n7548 & n14691;
  assign n18245 = ~n18242 & ~n18243;
  assign n18246 = ~n18241 & n18245;
  assign n18247 = ~n18244 & n18246;
  assign n18248 = pi11  & n18247;
  assign n18249 = ~pi11  & ~n18247;
  assign n18250 = ~n18248 & ~n18249;
  assign n18251 = n17759 & ~n17761;
  assign n18252 = ~n17762 & ~n18251;
  assign n18253 = ~n18250 & n18252;
  assign n18254 = n8161 & n12265;
  assign n18255 = n7847 & n12268;
  assign n18256 = n7554 & n12271;
  assign n18257 = n7548 & n14728;
  assign n18258 = ~n18255 & ~n18256;
  assign n18259 = ~n18254 & n18258;
  assign n18260 = ~n18257 & n18259;
  assign n18261 = ~pi11  & ~n18260;
  assign n18262 = pi11  & n18260;
  assign n18263 = ~n18261 & ~n18262;
  assign n18264 = pi14  & ~n17739;
  assign n18265 = n17746 & ~n18264;
  assign n18266 = ~n17746 & n18264;
  assign n18267 = ~n18265 & ~n18266;
  assign n18268 = ~n18263 & n18267;
  assign n18269 = n8161 & n12268;
  assign n18270 = n7847 & n12271;
  assign n18271 = n7554 & n12274;
  assign n18272 = n7548 & n14771;
  assign n18273 = ~n18270 & ~n18271;
  assign n18274 = ~n18269 & n18273;
  assign n18275 = ~n18272 & n18274;
  assign n18276 = pi11  & n18275;
  assign n18277 = ~pi11  & ~n18275;
  assign n18278 = ~n18276 & ~n18277;
  assign n18279 = n17733 & ~n17738;
  assign n18280 = ~n17739 & ~n18279;
  assign n18281 = ~n18278 & n18280;
  assign n18282 = n7547 & n12281;
  assign n18283 = pi11  & n18282;
  assign n18284 = n8161 & n12279;
  assign n18285 = n7847 & n12281;
  assign n18286 = n7548 & ~n14833;
  assign n18287 = ~n18284 & ~n18285;
  assign n18288 = ~n18286 & n18287;
  assign n18289 = ~n18283 & n18288;
  assign n18290 = n8161 & n12274;
  assign n18291 = n7847 & n12279;
  assign n18292 = n7554 & n12281;
  assign n18293 = n7548 & ~n14876;
  assign n18294 = ~n18291 & ~n18292;
  assign n18295 = ~n18290 & n18294;
  assign n18296 = ~n18293 & n18295;
  assign n18297 = pi11  & n18289;
  assign n18298 = n18296 & n18297;
  assign n18299 = n17732 & n18298;
  assign n18300 = n8161 & n12271;
  assign n18301 = n7847 & n12274;
  assign n18302 = n7554 & n12279;
  assign n18303 = n7548 & n14795;
  assign n18304 = ~n18301 & ~n18302;
  assign n18305 = ~n18300 & n18304;
  assign n18306 = ~n18303 & n18305;
  assign n18307 = pi11  & n18306;
  assign n18308 = ~pi11  & ~n18306;
  assign n18309 = ~n18307 & ~n18308;
  assign n18310 = ~n17732 & ~n18298;
  assign n18311 = ~n18299 & ~n18310;
  assign n18312 = ~n18309 & n18311;
  assign n18313 = ~n18299 & ~n18312;
  assign n18314 = n18278 & ~n18280;
  assign n18315 = ~n18281 & ~n18314;
  assign n18316 = ~n18313 & n18315;
  assign n18317 = ~n18281 & ~n18316;
  assign n18318 = n18263 & ~n18267;
  assign n18319 = ~n18268 & ~n18318;
  assign n18320 = ~n18317 & n18319;
  assign n18321 = ~n18268 & ~n18320;
  assign n18322 = n18250 & ~n18252;
  assign n18323 = ~n18253 & ~n18322;
  assign n18324 = ~n18321 & n18323;
  assign n18325 = ~n18253 & ~n18324;
  assign n18326 = n18237 & ~n18239;
  assign n18327 = ~n18240 & ~n18326;
  assign n18328 = ~n18325 & n18327;
  assign n18329 = ~n18240 & ~n18328;
  assign n18330 = ~n18216 & n18226;
  assign n18331 = ~n18227 & ~n18330;
  assign n18332 = ~n18329 & n18331;
  assign n18333 = ~n18227 & ~n18332;
  assign n18334 = ~n18203 & n18213;
  assign n18335 = ~n18214 & ~n18334;
  assign n18336 = ~n18333 & n18335;
  assign n18337 = ~n18214 & ~n18336;
  assign n18338 = ~n18190 & n18200;
  assign n18339 = ~n18201 & ~n18338;
  assign n18340 = ~n18337 & n18339;
  assign n18341 = ~n18201 & ~n18340;
  assign n18342 = n18185 & ~n18187;
  assign n18343 = ~n18188 & ~n18342;
  assign n18344 = ~n18341 & n18343;
  assign n18345 = ~n18188 & ~n18344;
  assign n18346 = n18172 & ~n18174;
  assign n18347 = ~n18175 & ~n18346;
  assign n18348 = ~n18345 & n18347;
  assign n18349 = ~n18175 & ~n18348;
  assign n18350 = n18159 & ~n18161;
  assign n18351 = ~n18162 & ~n18350;
  assign n18352 = ~n18349 & n18351;
  assign n18353 = ~n18162 & ~n18352;
  assign n18354 = ~n18138 & n18148;
  assign n18355 = ~n18149 & ~n18354;
  assign n18356 = ~n18353 & n18355;
  assign n18357 = ~n18149 & ~n18356;
  assign n18358 = ~n18125 & n18135;
  assign n18359 = ~n18136 & ~n18358;
  assign n18360 = ~n18357 & n18359;
  assign n18361 = ~n18136 & ~n18360;
  assign n18362 = ~n18112 & n18122;
  assign n18363 = ~n18123 & ~n18362;
  assign n18364 = ~n18361 & n18363;
  assign n18365 = ~n18123 & ~n18364;
  assign n18366 = n18107 & ~n18109;
  assign n18367 = ~n18110 & ~n18366;
  assign n18368 = ~n18365 & n18367;
  assign n18369 = ~n18110 & ~n18368;
  assign n18370 = n18094 & ~n18096;
  assign n18371 = ~n18097 & ~n18370;
  assign n18372 = ~n18369 & n18371;
  assign n18373 = ~n18097 & ~n18372;
  assign n18374 = n18081 & ~n18083;
  assign n18375 = ~n18084 & ~n18374;
  assign n18376 = ~n18373 & n18375;
  assign n18377 = ~n18084 & ~n18376;
  assign n18378 = ~n18060 & n18070;
  assign n18379 = ~n18071 & ~n18378;
  assign n18380 = ~n18377 & n18379;
  assign n18381 = ~n18071 & ~n18380;
  assign n18382 = ~n18047 & n18057;
  assign n18383 = ~n18058 & ~n18382;
  assign n18384 = ~n18381 & n18383;
  assign n18385 = ~n18058 & ~n18384;
  assign n18386 = n18042 & ~n18044;
  assign n18387 = ~n18045 & ~n18386;
  assign n18388 = ~n18385 & n18387;
  assign n18389 = ~n18045 & ~n18388;
  assign n18390 = n18029 & ~n18031;
  assign n18391 = ~n18032 & ~n18390;
  assign n18392 = ~n18389 & n18391;
  assign n18393 = ~n18032 & ~n18392;
  assign n18394 = n18016 & ~n18018;
  assign n18395 = ~n18019 & ~n18394;
  assign n18396 = ~n18393 & n18395;
  assign n18397 = ~n18019 & ~n18396;
  assign n18398 = n18003 & ~n18005;
  assign n18399 = ~n18006 & ~n18398;
  assign n18400 = ~n18397 & n18399;
  assign n18401 = ~n18006 & ~n18400;
  assign n18402 = n17990 & ~n17992;
  assign n18403 = ~n17993 & ~n18402;
  assign n18404 = ~n18401 & n18403;
  assign n18405 = ~n17993 & ~n18404;
  assign n18406 = n17977 & ~n17979;
  assign n18407 = ~n17980 & ~n18406;
  assign n18408 = ~n18405 & n18407;
  assign n18409 = ~n17980 & ~n18408;
  assign n18410 = n17964 & ~n17966;
  assign n18411 = ~n17967 & ~n18410;
  assign n18412 = ~n18409 & n18411;
  assign n18413 = ~n17967 & ~n18412;
  assign n18414 = n17951 & ~n17953;
  assign n18415 = ~n17954 & ~n18414;
  assign n18416 = ~n18413 & n18415;
  assign n18417 = ~n17954 & ~n18416;
  assign n18418 = n17938 & ~n17940;
  assign n18419 = ~n17941 & ~n18418;
  assign n18420 = ~n18417 & n18419;
  assign n18421 = ~n17941 & ~n18420;
  assign n18422 = n17925 & ~n17927;
  assign n18423 = ~n17928 & ~n18422;
  assign n18424 = ~n18421 & n18423;
  assign n18425 = ~n17928 & ~n18424;
  assign n18426 = ~n17868 & n17878;
  assign n18427 = ~n17879 & ~n18426;
  assign n18428 = ~n18425 & n18427;
  assign n18429 = n18425 & ~n18427;
  assign n18430 = ~n18428 & ~n18429;
  assign n18431 = n9355 & n12175;
  assign n18432 = n8939 & n12178;
  assign n18433 = n8206 & n12181;
  assign n18434 = n8200 & n12961;
  assign n18435 = ~n18432 & ~n18433;
  assign n18436 = ~n18431 & n18435;
  assign n18437 = ~n18434 & n18436;
  assign n18438 = pi8  & n18437;
  assign n18439 = ~pi8  & ~n18437;
  assign n18440 = ~n18438 & ~n18439;
  assign n18441 = n18430 & ~n18440;
  assign n18442 = ~n18428 & ~n18441;
  assign n18443 = ~n17885 & n17895;
  assign n18444 = ~n17896 & ~n18443;
  assign n18445 = ~n18442 & n18444;
  assign n18446 = n18442 & ~n18444;
  assign n18447 = ~n18445 & ~n18446;
  assign n18448 = n9830 & n13007;
  assign n18449 = n9836 & n12172;
  assign n18450 = ~n71 & n12165;
  assign n18451 = ~n12163 & ~n13942;
  assign n18452 = ~n18450 & n18451;
  assign n18453 = ~n18449 & ~n18452;
  assign n18454 = ~n18448 & n18453;
  assign n18455 = pi5  & n18454;
  assign n18456 = ~pi5  & ~n18454;
  assign n18457 = ~n18455 & ~n18456;
  assign n18458 = n18447 & ~n18457;
  assign n18459 = ~n18445 & ~n18458;
  assign n18460 = ~n17908 & ~n17910;
  assign n18461 = ~n17911 & ~n18460;
  assign n18462 = ~n18459 & n18461;
  assign n18463 = n18459 & ~n18461;
  assign n18464 = ~n18462 & ~n18463;
  assign n18465 = n18421 & ~n18423;
  assign n18466 = ~n18424 & ~n18465;
  assign n18467 = n9355 & n12178;
  assign n18468 = n8939 & n12181;
  assign n18469 = n8206 & n12184;
  assign n18470 = n8200 & n12880;
  assign n18471 = ~n18468 & ~n18469;
  assign n18472 = ~n18467 & n18471;
  assign n18473 = ~n18470 & n18472;
  assign n18474 = pi8  & n18473;
  assign n18475 = ~pi8  & ~n18473;
  assign n18476 = ~n18474 & ~n18475;
  assign n18477 = n18466 & ~n18476;
  assign n18478 = n18417 & ~n18419;
  assign n18479 = ~n18420 & ~n18478;
  assign n18480 = n9355 & n12181;
  assign n18481 = n8939 & n12184;
  assign n18482 = n8206 & n12187;
  assign n18483 = n8200 & n12608;
  assign n18484 = ~n18481 & ~n18482;
  assign n18485 = ~n18480 & n18484;
  assign n18486 = ~n18483 & n18485;
  assign n18487 = pi8  & n18486;
  assign n18488 = ~pi8  & ~n18486;
  assign n18489 = ~n18487 & ~n18488;
  assign n18490 = n18479 & ~n18489;
  assign n18491 = n18413 & ~n18415;
  assign n18492 = ~n18416 & ~n18491;
  assign n18493 = n9355 & n12184;
  assign n18494 = n8939 & n12187;
  assign n18495 = n8206 & n12190;
  assign n18496 = n8200 & n12845;
  assign n18497 = ~n18494 & ~n18495;
  assign n18498 = ~n18493 & n18497;
  assign n18499 = ~n18496 & n18498;
  assign n18500 = pi8  & n18499;
  assign n18501 = ~pi8  & ~n18499;
  assign n18502 = ~n18500 & ~n18501;
  assign n18503 = n18492 & ~n18502;
  assign n18504 = n18409 & ~n18411;
  assign n18505 = ~n18412 & ~n18504;
  assign n18506 = n9355 & n12187;
  assign n18507 = n8939 & n12190;
  assign n18508 = n8206 & n12193;
  assign n18509 = n8200 & n12921;
  assign n18510 = ~n18507 & ~n18508;
  assign n18511 = ~n18506 & n18510;
  assign n18512 = ~n18509 & n18511;
  assign n18513 = pi8  & n18512;
  assign n18514 = ~pi8  & ~n18512;
  assign n18515 = ~n18513 & ~n18514;
  assign n18516 = n18505 & ~n18515;
  assign n18517 = n18405 & ~n18407;
  assign n18518 = ~n18408 & ~n18517;
  assign n18519 = n9355 & n12190;
  assign n18520 = n8939 & n12193;
  assign n18521 = n8206 & n12196;
  assign n18522 = n8200 & n12530;
  assign n18523 = ~n18520 & ~n18521;
  assign n18524 = ~n18519 & n18523;
  assign n18525 = ~n18522 & n18524;
  assign n18526 = pi8  & n18525;
  assign n18527 = ~pi8  & ~n18525;
  assign n18528 = ~n18526 & ~n18527;
  assign n18529 = n18518 & ~n18528;
  assign n18530 = n18401 & ~n18403;
  assign n18531 = ~n18404 & ~n18530;
  assign n18532 = n9355 & n12193;
  assign n18533 = n8939 & n12196;
  assign n18534 = n8206 & n12199;
  assign n18535 = n8200 & n12594;
  assign n18536 = ~n18533 & ~n18534;
  assign n18537 = ~n18532 & n18536;
  assign n18538 = ~n18535 & n18537;
  assign n18539 = pi8  & n18538;
  assign n18540 = ~pi8  & ~n18538;
  assign n18541 = ~n18539 & ~n18540;
  assign n18542 = n18531 & ~n18541;
  assign n18543 = n18397 & ~n18399;
  assign n18544 = ~n18400 & ~n18543;
  assign n18545 = n9355 & n12196;
  assign n18546 = n8939 & n12199;
  assign n18547 = n8206 & n12202;
  assign n18548 = n8200 & n12578;
  assign n18549 = ~n18546 & ~n18547;
  assign n18550 = ~n18545 & n18549;
  assign n18551 = ~n18548 & n18550;
  assign n18552 = pi8  & n18551;
  assign n18553 = ~pi8  & ~n18551;
  assign n18554 = ~n18552 & ~n18553;
  assign n18555 = n18544 & ~n18554;
  assign n18556 = n18393 & ~n18395;
  assign n18557 = ~n18396 & ~n18556;
  assign n18558 = n9355 & n12199;
  assign n18559 = n8939 & n12202;
  assign n18560 = n8206 & n12205;
  assign n18561 = n8200 & n12683;
  assign n18562 = ~n18559 & ~n18560;
  assign n18563 = ~n18558 & n18562;
  assign n18564 = ~n18561 & n18563;
  assign n18565 = pi8  & n18564;
  assign n18566 = ~pi8  & ~n18564;
  assign n18567 = ~n18565 & ~n18566;
  assign n18568 = n18557 & ~n18567;
  assign n18569 = n18389 & ~n18391;
  assign n18570 = ~n18392 & ~n18569;
  assign n18571 = n9355 & n12202;
  assign n18572 = n8939 & n12205;
  assign n18573 = n8206 & n12208;
  assign n18574 = n8200 & n12701;
  assign n18575 = ~n18572 & ~n18573;
  assign n18576 = ~n18571 & n18575;
  assign n18577 = ~n18574 & n18576;
  assign n18578 = pi8  & n18577;
  assign n18579 = ~pi8  & ~n18577;
  assign n18580 = ~n18578 & ~n18579;
  assign n18581 = n18570 & ~n18580;
  assign n18582 = n18385 & ~n18387;
  assign n18583 = ~n18388 & ~n18582;
  assign n18584 = n9355 & n12205;
  assign n18585 = n8939 & n12208;
  assign n18586 = n8206 & n12211;
  assign n18587 = n8200 & n13031;
  assign n18588 = ~n18585 & ~n18586;
  assign n18589 = ~n18584 & n18588;
  assign n18590 = ~n18587 & n18589;
  assign n18591 = pi8  & n18590;
  assign n18592 = ~pi8  & ~n18590;
  assign n18593 = ~n18591 & ~n18592;
  assign n18594 = n18583 & ~n18593;
  assign n18595 = n9355 & n12208;
  assign n18596 = n8939 & n12211;
  assign n18597 = n8206 & n12214;
  assign n18598 = n8200 & n12804;
  assign n18599 = ~n18596 & ~n18597;
  assign n18600 = ~n18595 & n18599;
  assign n18601 = ~n18598 & n18600;
  assign n18602 = ~pi8  & ~n18601;
  assign n18603 = pi8  & n18601;
  assign n18604 = ~n18602 & ~n18603;
  assign n18605 = n18381 & ~n18383;
  assign n18606 = ~n18384 & ~n18605;
  assign n18607 = ~n18604 & n18606;
  assign n18608 = n9355 & n12211;
  assign n18609 = n8939 & n12214;
  assign n18610 = n8206 & n12217;
  assign n18611 = n8200 & n13203;
  assign n18612 = ~n18609 & ~n18610;
  assign n18613 = ~n18608 & n18612;
  assign n18614 = ~n18611 & n18613;
  assign n18615 = ~pi8  & ~n18614;
  assign n18616 = pi8  & n18614;
  assign n18617 = ~n18615 & ~n18616;
  assign n18618 = n18377 & ~n18379;
  assign n18619 = ~n18380 & ~n18618;
  assign n18620 = ~n18617 & n18619;
  assign n18621 = n18373 & ~n18375;
  assign n18622 = ~n18376 & ~n18621;
  assign n18623 = n9355 & n12214;
  assign n18624 = n8939 & n12217;
  assign n18625 = n8206 & n12220;
  assign n18626 = n8200 & n13187;
  assign n18627 = ~n18624 & ~n18625;
  assign n18628 = ~n18623 & n18627;
  assign n18629 = ~n18626 & n18628;
  assign n18630 = pi8  & n18629;
  assign n18631 = ~pi8  & ~n18629;
  assign n18632 = ~n18630 & ~n18631;
  assign n18633 = n18622 & ~n18632;
  assign n18634 = n18369 & ~n18371;
  assign n18635 = ~n18372 & ~n18634;
  assign n18636 = n9355 & n12217;
  assign n18637 = n8939 & n12220;
  assign n18638 = n8206 & n12223;
  assign n18639 = n8200 & n13374;
  assign n18640 = ~n18637 & ~n18638;
  assign n18641 = ~n18636 & n18640;
  assign n18642 = ~n18639 & n18641;
  assign n18643 = pi8  & n18642;
  assign n18644 = ~pi8  & ~n18642;
  assign n18645 = ~n18643 & ~n18644;
  assign n18646 = n18635 & ~n18645;
  assign n18647 = n18365 & ~n18367;
  assign n18648 = ~n18368 & ~n18647;
  assign n18649 = n9355 & n12220;
  assign n18650 = n8939 & n12223;
  assign n18651 = n8206 & n12226;
  assign n18652 = n8200 & n13392;
  assign n18653 = ~n18650 & ~n18651;
  assign n18654 = ~n18649 & n18653;
  assign n18655 = ~n18652 & n18654;
  assign n18656 = pi8  & n18655;
  assign n18657 = ~pi8  & ~n18655;
  assign n18658 = ~n18656 & ~n18657;
  assign n18659 = n18648 & ~n18658;
  assign n18660 = n9355 & n12223;
  assign n18661 = n8939 & n12226;
  assign n18662 = n8206 & n12229;
  assign n18663 = n8200 & n13745;
  assign n18664 = ~n18661 & ~n18662;
  assign n18665 = ~n18660 & n18664;
  assign n18666 = ~n18663 & n18665;
  assign n18667 = ~pi8  & ~n18666;
  assign n18668 = pi8  & n18666;
  assign n18669 = ~n18667 & ~n18668;
  assign n18670 = n18361 & ~n18363;
  assign n18671 = ~n18364 & ~n18670;
  assign n18672 = ~n18669 & n18671;
  assign n18673 = n9355 & n12226;
  assign n18674 = n8939 & n12229;
  assign n18675 = n8206 & n12232;
  assign n18676 = n8200 & n13530;
  assign n18677 = ~n18674 & ~n18675;
  assign n18678 = ~n18673 & n18677;
  assign n18679 = ~n18676 & n18678;
  assign n18680 = ~pi8  & ~n18679;
  assign n18681 = pi8  & n18679;
  assign n18682 = ~n18680 & ~n18681;
  assign n18683 = n18357 & ~n18359;
  assign n18684 = ~n18360 & ~n18683;
  assign n18685 = ~n18682 & n18684;
  assign n18686 = n9355 & n12229;
  assign n18687 = n8939 & n12232;
  assign n18688 = n8206 & n12235;
  assign n18689 = n8200 & n13979;
  assign n18690 = ~n18687 & ~n18688;
  assign n18691 = ~n18686 & n18690;
  assign n18692 = ~n18689 & n18691;
  assign n18693 = ~pi8  & ~n18692;
  assign n18694 = pi8  & n18692;
  assign n18695 = ~n18693 & ~n18694;
  assign n18696 = n18353 & ~n18355;
  assign n18697 = ~n18356 & ~n18696;
  assign n18698 = ~n18695 & n18697;
  assign n18699 = n18349 & ~n18351;
  assign n18700 = ~n18352 & ~n18699;
  assign n18701 = n9355 & n12232;
  assign n18702 = n8939 & n12235;
  assign n18703 = n8206 & n12238;
  assign n18704 = n8200 & n14116;
  assign n18705 = ~n18702 & ~n18703;
  assign n18706 = ~n18701 & n18705;
  assign n18707 = ~n18704 & n18706;
  assign n18708 = pi8  & n18707;
  assign n18709 = ~pi8  & ~n18707;
  assign n18710 = ~n18708 & ~n18709;
  assign n18711 = n18700 & ~n18710;
  assign n18712 = n18345 & ~n18347;
  assign n18713 = ~n18348 & ~n18712;
  assign n18714 = n9355 & n12235;
  assign n18715 = n8939 & n12238;
  assign n18716 = n8206 & n12241;
  assign n18717 = n8200 & n13959;
  assign n18718 = ~n18715 & ~n18716;
  assign n18719 = ~n18714 & n18718;
  assign n18720 = ~n18717 & n18719;
  assign n18721 = pi8  & n18720;
  assign n18722 = ~pi8  & ~n18720;
  assign n18723 = ~n18721 & ~n18722;
  assign n18724 = n18713 & ~n18723;
  assign n18725 = n18341 & ~n18343;
  assign n18726 = ~n18344 & ~n18725;
  assign n18727 = n9355 & n12238;
  assign n18728 = n8939 & n12241;
  assign n18729 = n8206 & n12244;
  assign n18730 = n8200 & n14229;
  assign n18731 = ~n18728 & ~n18729;
  assign n18732 = ~n18727 & n18731;
  assign n18733 = ~n18730 & n18732;
  assign n18734 = pi8  & n18733;
  assign n18735 = ~pi8  & ~n18733;
  assign n18736 = ~n18734 & ~n18735;
  assign n18737 = n18726 & ~n18736;
  assign n18738 = n9355 & n12241;
  assign n18739 = n8939 & n12244;
  assign n18740 = n8206 & n12247;
  assign n18741 = n8200 & n14515;
  assign n18742 = ~n18739 & ~n18740;
  assign n18743 = ~n18738 & n18742;
  assign n18744 = ~n18741 & n18743;
  assign n18745 = ~pi8  & ~n18744;
  assign n18746 = pi8  & n18744;
  assign n18747 = ~n18745 & ~n18746;
  assign n18748 = n18337 & ~n18339;
  assign n18749 = ~n18340 & ~n18748;
  assign n18750 = ~n18747 & n18749;
  assign n18751 = n9355 & n12244;
  assign n18752 = n8939 & n12247;
  assign n18753 = n8206 & n12250;
  assign n18754 = n8200 & n14527;
  assign n18755 = ~n18752 & ~n18753;
  assign n18756 = ~n18751 & n18755;
  assign n18757 = ~n18754 & n18756;
  assign n18758 = ~pi8  & ~n18757;
  assign n18759 = pi8  & n18757;
  assign n18760 = ~n18758 & ~n18759;
  assign n18761 = n18333 & ~n18335;
  assign n18762 = ~n18336 & ~n18761;
  assign n18763 = ~n18760 & n18762;
  assign n18764 = n9355 & n12247;
  assign n18765 = n8939 & n12250;
  assign n18766 = n8206 & n12253;
  assign n18767 = n8200 & n14207;
  assign n18768 = ~n18765 & ~n18766;
  assign n18769 = ~n18764 & n18768;
  assign n18770 = ~n18767 & n18769;
  assign n18771 = ~pi8  & ~n18770;
  assign n18772 = pi8  & n18770;
  assign n18773 = ~n18771 & ~n18772;
  assign n18774 = n18329 & ~n18331;
  assign n18775 = ~n18332 & ~n18774;
  assign n18776 = ~n18773 & n18775;
  assign n18777 = n18325 & ~n18327;
  assign n18778 = ~n18328 & ~n18777;
  assign n18779 = n9355 & n12250;
  assign n18780 = n8939 & n12253;
  assign n18781 = n8206 & n12256;
  assign n18782 = n8200 & n14559;
  assign n18783 = ~n18780 & ~n18781;
  assign n18784 = ~n18779 & n18783;
  assign n18785 = ~n18782 & n18784;
  assign n18786 = pi8  & n18785;
  assign n18787 = ~pi8  & ~n18785;
  assign n18788 = ~n18786 & ~n18787;
  assign n18789 = n18778 & ~n18788;
  assign n18790 = n18321 & ~n18323;
  assign n18791 = ~n18324 & ~n18790;
  assign n18792 = n9355 & n12253;
  assign n18793 = n8939 & n12256;
  assign n18794 = n8206 & n12259;
  assign n18795 = n8200 & n14584;
  assign n18796 = ~n18793 & ~n18794;
  assign n18797 = ~n18792 & n18796;
  assign n18798 = ~n18795 & n18797;
  assign n18799 = pi8  & n18798;
  assign n18800 = ~pi8  & ~n18798;
  assign n18801 = ~n18799 & ~n18800;
  assign n18802 = n18791 & ~n18801;
  assign n18803 = n18317 & ~n18319;
  assign n18804 = ~n18320 & ~n18803;
  assign n18805 = n9355 & n12256;
  assign n18806 = n8939 & n12259;
  assign n18807 = n8206 & n12262;
  assign n18808 = n8200 & n14608;
  assign n18809 = ~n18806 & ~n18807;
  assign n18810 = ~n18805 & n18809;
  assign n18811 = ~n18808 & n18810;
  assign n18812 = pi8  & n18811;
  assign n18813 = ~pi8  & ~n18811;
  assign n18814 = ~n18812 & ~n18813;
  assign n18815 = n18804 & ~n18814;
  assign n18816 = n9355 & n12259;
  assign n18817 = n8939 & n12262;
  assign n18818 = n8206 & n12265;
  assign n18819 = n8200 & n14637;
  assign n18820 = ~n18817 & ~n18818;
  assign n18821 = ~n18816 & n18820;
  assign n18822 = ~n18819 & n18821;
  assign n18823 = ~pi8  & ~n18822;
  assign n18824 = pi8  & n18822;
  assign n18825 = ~n18823 & ~n18824;
  assign n18826 = n18313 & ~n18315;
  assign n18827 = ~n18316 & ~n18826;
  assign n18828 = ~n18825 & n18827;
  assign n18829 = n9355 & n12262;
  assign n18830 = n8939 & n12265;
  assign n18831 = n8206 & n12268;
  assign n18832 = n8200 & n14691;
  assign n18833 = ~n18830 & ~n18831;
  assign n18834 = ~n18829 & n18833;
  assign n18835 = ~n18832 & n18834;
  assign n18836 = pi8  & n18835;
  assign n18837 = ~pi8  & ~n18835;
  assign n18838 = ~n18836 & ~n18837;
  assign n18839 = n18309 & ~n18311;
  assign n18840 = ~n18312 & ~n18839;
  assign n18841 = ~n18838 & n18840;
  assign n18842 = n9355 & n12265;
  assign n18843 = n8939 & n12268;
  assign n18844 = n8206 & n12271;
  assign n18845 = n8200 & n14728;
  assign n18846 = ~n18843 & ~n18844;
  assign n18847 = ~n18842 & n18846;
  assign n18848 = ~n18845 & n18847;
  assign n18849 = ~pi8  & ~n18848;
  assign n18850 = pi8  & n18848;
  assign n18851 = ~n18849 & ~n18850;
  assign n18852 = pi11  & ~n18289;
  assign n18853 = n18296 & ~n18852;
  assign n18854 = ~n18296 & n18852;
  assign n18855 = ~n18853 & ~n18854;
  assign n18856 = ~n18851 & n18855;
  assign n18857 = n9355 & n12268;
  assign n18858 = n8939 & n12271;
  assign n18859 = n8206 & n12274;
  assign n18860 = n8200 & n14771;
  assign n18861 = ~n18858 & ~n18859;
  assign n18862 = ~n18857 & n18861;
  assign n18863 = ~n18860 & n18862;
  assign n18864 = pi8  & n18863;
  assign n18865 = ~pi8  & ~n18863;
  assign n18866 = ~n18864 & ~n18865;
  assign n18867 = n18283 & ~n18288;
  assign n18868 = ~n18289 & ~n18867;
  assign n18869 = ~n18866 & n18868;
  assign n18870 = n8199 & n12281;
  assign n18871 = pi8  & n18870;
  assign n18872 = n9355 & n12279;
  assign n18873 = n8939 & n12281;
  assign n18874 = n8200 & ~n14833;
  assign n18875 = ~n18872 & ~n18873;
  assign n18876 = ~n18874 & n18875;
  assign n18877 = ~n18871 & n18876;
  assign n18878 = n9355 & n12274;
  assign n18879 = n8939 & n12279;
  assign n18880 = n8206 & n12281;
  assign n18881 = n8200 & ~n14876;
  assign n18882 = ~n18879 & ~n18880;
  assign n18883 = ~n18878 & n18882;
  assign n18884 = ~n18881 & n18883;
  assign n18885 = pi8  & n18877;
  assign n18886 = n18884 & n18885;
  assign n18887 = n18282 & n18886;
  assign n18888 = n9355 & n12271;
  assign n18889 = n8939 & n12274;
  assign n18890 = n8206 & n12279;
  assign n18891 = n8200 & n14795;
  assign n18892 = ~n18889 & ~n18890;
  assign n18893 = ~n18888 & n18892;
  assign n18894 = ~n18891 & n18893;
  assign n18895 = pi8  & n18894;
  assign n18896 = ~pi8  & ~n18894;
  assign n18897 = ~n18895 & ~n18896;
  assign n18898 = ~n18282 & ~n18886;
  assign n18899 = ~n18887 & ~n18898;
  assign n18900 = ~n18897 & n18899;
  assign n18901 = ~n18887 & ~n18900;
  assign n18902 = n18866 & ~n18868;
  assign n18903 = ~n18869 & ~n18902;
  assign n18904 = ~n18901 & n18903;
  assign n18905 = ~n18869 & ~n18904;
  assign n18906 = n18851 & ~n18855;
  assign n18907 = ~n18856 & ~n18906;
  assign n18908 = ~n18905 & n18907;
  assign n18909 = ~n18856 & ~n18908;
  assign n18910 = n18838 & ~n18840;
  assign n18911 = ~n18841 & ~n18910;
  assign n18912 = ~n18909 & n18911;
  assign n18913 = ~n18841 & ~n18912;
  assign n18914 = n18825 & ~n18827;
  assign n18915 = ~n18828 & ~n18914;
  assign n18916 = ~n18913 & n18915;
  assign n18917 = ~n18828 & ~n18916;
  assign n18918 = ~n18804 & n18814;
  assign n18919 = ~n18815 & ~n18918;
  assign n18920 = ~n18917 & n18919;
  assign n18921 = ~n18815 & ~n18920;
  assign n18922 = ~n18791 & n18801;
  assign n18923 = ~n18802 & ~n18922;
  assign n18924 = ~n18921 & n18923;
  assign n18925 = ~n18802 & ~n18924;
  assign n18926 = ~n18778 & n18788;
  assign n18927 = ~n18789 & ~n18926;
  assign n18928 = ~n18925 & n18927;
  assign n18929 = ~n18789 & ~n18928;
  assign n18930 = n18773 & ~n18775;
  assign n18931 = ~n18776 & ~n18930;
  assign n18932 = ~n18929 & n18931;
  assign n18933 = ~n18776 & ~n18932;
  assign n18934 = n18760 & ~n18762;
  assign n18935 = ~n18763 & ~n18934;
  assign n18936 = ~n18933 & n18935;
  assign n18937 = ~n18763 & ~n18936;
  assign n18938 = n18747 & ~n18749;
  assign n18939 = ~n18750 & ~n18938;
  assign n18940 = ~n18937 & n18939;
  assign n18941 = ~n18750 & ~n18940;
  assign n18942 = ~n18726 & n18736;
  assign n18943 = ~n18737 & ~n18942;
  assign n18944 = ~n18941 & n18943;
  assign n18945 = ~n18737 & ~n18944;
  assign n18946 = ~n18713 & n18723;
  assign n18947 = ~n18724 & ~n18946;
  assign n18948 = ~n18945 & n18947;
  assign n18949 = ~n18724 & ~n18948;
  assign n18950 = ~n18700 & n18710;
  assign n18951 = ~n18711 & ~n18950;
  assign n18952 = ~n18949 & n18951;
  assign n18953 = ~n18711 & ~n18952;
  assign n18954 = n18695 & ~n18697;
  assign n18955 = ~n18698 & ~n18954;
  assign n18956 = ~n18953 & n18955;
  assign n18957 = ~n18698 & ~n18956;
  assign n18958 = n18682 & ~n18684;
  assign n18959 = ~n18685 & ~n18958;
  assign n18960 = ~n18957 & n18959;
  assign n18961 = ~n18685 & ~n18960;
  assign n18962 = n18669 & ~n18671;
  assign n18963 = ~n18672 & ~n18962;
  assign n18964 = ~n18961 & n18963;
  assign n18965 = ~n18672 & ~n18964;
  assign n18966 = ~n18648 & n18658;
  assign n18967 = ~n18659 & ~n18966;
  assign n18968 = ~n18965 & n18967;
  assign n18969 = ~n18659 & ~n18968;
  assign n18970 = ~n18635 & n18645;
  assign n18971 = ~n18646 & ~n18970;
  assign n18972 = ~n18969 & n18971;
  assign n18973 = ~n18646 & ~n18972;
  assign n18974 = ~n18622 & n18632;
  assign n18975 = ~n18633 & ~n18974;
  assign n18976 = ~n18973 & n18975;
  assign n18977 = ~n18633 & ~n18976;
  assign n18978 = n18617 & ~n18619;
  assign n18979 = ~n18620 & ~n18978;
  assign n18980 = ~n18977 & n18979;
  assign n18981 = ~n18620 & ~n18980;
  assign n18982 = n18604 & ~n18606;
  assign n18983 = ~n18607 & ~n18982;
  assign n18984 = ~n18981 & n18983;
  assign n18985 = ~n18607 & ~n18984;
  assign n18986 = ~n18583 & n18593;
  assign n18987 = ~n18594 & ~n18986;
  assign n18988 = ~n18985 & n18987;
  assign n18989 = ~n18594 & ~n18988;
  assign n18990 = ~n18570 & n18580;
  assign n18991 = ~n18581 & ~n18990;
  assign n18992 = ~n18989 & n18991;
  assign n18993 = ~n18581 & ~n18992;
  assign n18994 = ~n18557 & n18567;
  assign n18995 = ~n18568 & ~n18994;
  assign n18996 = ~n18993 & n18995;
  assign n18997 = ~n18568 & ~n18996;
  assign n18998 = ~n18544 & n18554;
  assign n18999 = ~n18555 & ~n18998;
  assign n19000 = ~n18997 & n18999;
  assign n19001 = ~n18555 & ~n19000;
  assign n19002 = ~n18531 & n18541;
  assign n19003 = ~n18542 & ~n19002;
  assign n19004 = ~n19001 & n19003;
  assign n19005 = ~n18542 & ~n19004;
  assign n19006 = ~n18518 & n18528;
  assign n19007 = ~n18529 & ~n19006;
  assign n19008 = ~n19005 & n19007;
  assign n19009 = ~n18529 & ~n19008;
  assign n19010 = ~n18505 & n18515;
  assign n19011 = ~n18516 & ~n19010;
  assign n19012 = ~n19009 & n19011;
  assign n19013 = ~n18516 & ~n19012;
  assign n19014 = ~n18492 & n18502;
  assign n19015 = ~n18503 & ~n19014;
  assign n19016 = ~n19013 & n19015;
  assign n19017 = ~n18503 & ~n19016;
  assign n19018 = ~n18479 & n18489;
  assign n19019 = ~n18490 & ~n19018;
  assign n19020 = ~n19017 & n19019;
  assign n19021 = ~n18490 & ~n19020;
  assign n19022 = ~n18466 & n18476;
  assign n19023 = ~n18477 & ~n19022;
  assign n19024 = ~n19021 & n19023;
  assign n19025 = ~n18477 & ~n19024;
  assign n19026 = ~n18430 & n18440;
  assign n19027 = ~n18441 & ~n19026;
  assign n19028 = ~n19025 & n19027;
  assign n19029 = n19025 & ~n19027;
  assign n19030 = ~n19028 & ~n19029;
  assign n19031 = n71 & n12166;
  assign n19032 = n10329 & n12172;
  assign n19033 = n9836 & n12168;
  assign n19034 = n9830 & n13106;
  assign n19035 = ~n19031 & ~n19033;
  assign n19036 = ~n19032 & n19035;
  assign n19037 = ~n19034 & n19036;
  assign n19038 = pi5  & n19037;
  assign n19039 = ~pi5  & ~n19037;
  assign n19040 = ~n19038 & ~n19039;
  assign n19041 = n19030 & ~n19040;
  assign n19042 = ~n19028 & ~n19041;
  assign n19043 = ~n18447 & n18457;
  assign n19044 = ~n18458 & ~n19043;
  assign n19045 = ~n19042 & n19044;
  assign n19046 = n19042 & ~n19044;
  assign n19047 = ~n19045 & ~n19046;
  assign n19048 = n71 & n12172;
  assign n19049 = n10329 & n12168;
  assign n19050 = n9836 & n12175;
  assign n19051 = n9830 & n12939;
  assign n19052 = ~n19049 & ~n19050;
  assign n19053 = ~n19048 & n19052;
  assign n19054 = ~n19051 & n19053;
  assign n19055 = ~pi5  & ~n19054;
  assign n19056 = pi5  & n19054;
  assign n19057 = ~n19055 & ~n19056;
  assign n19058 = n19021 & ~n19023;
  assign n19059 = ~n19024 & ~n19058;
  assign n19060 = ~n19057 & n19059;
  assign n19061 = n10884 & ~n12424;
  assign n19062 = n10883 & ~n12165;
  assign n19063 = ~n11463 & ~n11476;
  assign n19064 = ~n19062 & n19063;
  assign n19065 = ~n12163 & ~n19064;
  assign n19066 = ~n19061 & ~n19065;
  assign n19067 = pi2  & n19066;
  assign n19068 = ~pi2  & ~n19066;
  assign n19069 = ~n19067 & ~n19068;
  assign n19070 = n19057 & ~n19059;
  assign n19071 = ~n19060 & ~n19070;
  assign n19072 = ~n19069 & n19071;
  assign n19073 = ~n19060 & ~n19072;
  assign n19074 = ~n19030 & n19040;
  assign n19075 = ~n19041 & ~n19074;
  assign n19076 = ~n19073 & n19075;
  assign n19077 = n19073 & ~n19075;
  assign n19078 = ~n19076 & ~n19077;
  assign n19079 = n71 & n12168;
  assign n19080 = n10329 & n12175;
  assign n19081 = n9836 & n12178;
  assign n19082 = n9830 & n12862;
  assign n19083 = ~n19080 & ~n19081;
  assign n19084 = ~n19079 & n19083;
  assign n19085 = ~n19082 & n19084;
  assign n19086 = ~pi5  & ~n19085;
  assign n19087 = pi5  & n19085;
  assign n19088 = ~n19086 & ~n19087;
  assign n19089 = n19017 & ~n19019;
  assign n19090 = ~n19020 & ~n19089;
  assign n19091 = ~n19088 & n19090;
  assign n19092 = n71 & n12175;
  assign n19093 = n10329 & n12178;
  assign n19094 = n9836 & n12181;
  assign n19095 = n9830 & n12961;
  assign n19096 = ~n19093 & ~n19094;
  assign n19097 = ~n19092 & n19096;
  assign n19098 = ~n19095 & n19097;
  assign n19099 = ~pi5  & ~n19098;
  assign n19100 = pi5  & n19098;
  assign n19101 = ~n19099 & ~n19100;
  assign n19102 = n19013 & ~n19015;
  assign n19103 = ~n19016 & ~n19102;
  assign n19104 = ~n19101 & n19103;
  assign n19105 = n71 & n12178;
  assign n19106 = n10329 & n12181;
  assign n19107 = n9836 & n12184;
  assign n19108 = n9830 & n12880;
  assign n19109 = ~n19106 & ~n19107;
  assign n19110 = ~n19105 & n19109;
  assign n19111 = ~n19108 & n19110;
  assign n19112 = ~pi5  & ~n19111;
  assign n19113 = pi5  & n19111;
  assign n19114 = ~n19112 & ~n19113;
  assign n19115 = n19009 & ~n19011;
  assign n19116 = ~n19012 & ~n19115;
  assign n19117 = ~n19114 & n19116;
  assign n19118 = n71 & n12181;
  assign n19119 = n10329 & n12184;
  assign n19120 = n9836 & n12187;
  assign n19121 = n9830 & n12608;
  assign n19122 = ~n19119 & ~n19120;
  assign n19123 = ~n19118 & n19122;
  assign n19124 = ~n19121 & n19123;
  assign n19125 = ~pi5  & ~n19124;
  assign n19126 = pi5  & n19124;
  assign n19127 = ~n19125 & ~n19126;
  assign n19128 = n19005 & ~n19007;
  assign n19129 = ~n19008 & ~n19128;
  assign n19130 = ~n19127 & n19129;
  assign n19131 = n71 & n12184;
  assign n19132 = n10329 & n12187;
  assign n19133 = n9836 & n12190;
  assign n19134 = n9830 & n12845;
  assign n19135 = ~n19132 & ~n19133;
  assign n19136 = ~n19131 & n19135;
  assign n19137 = ~n19134 & n19136;
  assign n19138 = ~pi5  & ~n19137;
  assign n19139 = pi5  & n19137;
  assign n19140 = ~n19138 & ~n19139;
  assign n19141 = n19001 & ~n19003;
  assign n19142 = ~n19004 & ~n19141;
  assign n19143 = ~n19140 & n19142;
  assign n19144 = n71 & n12187;
  assign n19145 = n10329 & n12190;
  assign n19146 = n9836 & n12193;
  assign n19147 = n9830 & n12921;
  assign n19148 = ~n19145 & ~n19146;
  assign n19149 = ~n19144 & n19148;
  assign n19150 = ~n19147 & n19149;
  assign n19151 = ~pi5  & ~n19150;
  assign n19152 = pi5  & n19150;
  assign n19153 = ~n19151 & ~n19152;
  assign n19154 = n18997 & ~n18999;
  assign n19155 = ~n19000 & ~n19154;
  assign n19156 = ~n19153 & n19155;
  assign n19157 = n71 & n12190;
  assign n19158 = n10329 & n12193;
  assign n19159 = n9836 & n12196;
  assign n19160 = n9830 & n12530;
  assign n19161 = ~n19158 & ~n19159;
  assign n19162 = ~n19157 & n19161;
  assign n19163 = ~n19160 & n19162;
  assign n19164 = ~pi5  & ~n19163;
  assign n19165 = pi5  & n19163;
  assign n19166 = ~n19164 & ~n19165;
  assign n19167 = n18993 & ~n18995;
  assign n19168 = ~n18996 & ~n19167;
  assign n19169 = ~n19166 & n19168;
  assign n19170 = n71 & n12193;
  assign n19171 = n10329 & n12196;
  assign n19172 = n9836 & n12199;
  assign n19173 = n9830 & n12594;
  assign n19174 = ~n19171 & ~n19172;
  assign n19175 = ~n19170 & n19174;
  assign n19176 = ~n19173 & n19175;
  assign n19177 = ~pi5  & ~n19176;
  assign n19178 = pi5  & n19176;
  assign n19179 = ~n19177 & ~n19178;
  assign n19180 = n18989 & ~n18991;
  assign n19181 = ~n18992 & ~n19180;
  assign n19182 = ~n19179 & n19181;
  assign n19183 = n71 & n12196;
  assign n19184 = n10329 & n12199;
  assign n19185 = n9836 & n12202;
  assign n19186 = n9830 & n12578;
  assign n19187 = ~n19184 & ~n19185;
  assign n19188 = ~n19183 & n19187;
  assign n19189 = ~n19186 & n19188;
  assign n19190 = ~pi5  & ~n19189;
  assign n19191 = pi5  & n19189;
  assign n19192 = ~n19190 & ~n19191;
  assign n19193 = n18985 & ~n18987;
  assign n19194 = ~n18988 & ~n19193;
  assign n19195 = ~n19192 & n19194;
  assign n19196 = n18981 & ~n18983;
  assign n19197 = ~n18984 & ~n19196;
  assign n19198 = n71 & n12199;
  assign n19199 = n10329 & n12202;
  assign n19200 = n9836 & n12205;
  assign n19201 = n9830 & n12683;
  assign n19202 = ~n19199 & ~n19200;
  assign n19203 = ~n19198 & n19202;
  assign n19204 = ~n19201 & n19203;
  assign n19205 = pi5  & n19204;
  assign n19206 = ~pi5  & ~n19204;
  assign n19207 = ~n19205 & ~n19206;
  assign n19208 = n19197 & ~n19207;
  assign n19209 = n18977 & ~n18979;
  assign n19210 = ~n18980 & ~n19209;
  assign n19211 = n71 & n12202;
  assign n19212 = n10329 & n12205;
  assign n19213 = n9836 & n12208;
  assign n19214 = n9830 & n12701;
  assign n19215 = ~n19212 & ~n19213;
  assign n19216 = ~n19211 & n19215;
  assign n19217 = ~n19214 & n19216;
  assign n19218 = pi5  & n19217;
  assign n19219 = ~pi5  & ~n19217;
  assign n19220 = ~n19218 & ~n19219;
  assign n19221 = n19210 & ~n19220;
  assign n19222 = n71 & n12205;
  assign n19223 = n10329 & n12208;
  assign n19224 = n9836 & n12211;
  assign n19225 = n9830 & n13031;
  assign n19226 = ~n19223 & ~n19224;
  assign n19227 = ~n19222 & n19226;
  assign n19228 = ~n19225 & n19227;
  assign n19229 = ~pi5  & ~n19228;
  assign n19230 = pi5  & n19228;
  assign n19231 = ~n19229 & ~n19230;
  assign n19232 = n18973 & ~n18975;
  assign n19233 = ~n18976 & ~n19232;
  assign n19234 = ~n19231 & n19233;
  assign n19235 = n71 & n12208;
  assign n19236 = n10329 & n12211;
  assign n19237 = n9836 & n12214;
  assign n19238 = n9830 & n12804;
  assign n19239 = ~n19236 & ~n19237;
  assign n19240 = ~n19235 & n19239;
  assign n19241 = ~n19238 & n19240;
  assign n19242 = ~pi5  & ~n19241;
  assign n19243 = pi5  & n19241;
  assign n19244 = ~n19242 & ~n19243;
  assign n19245 = n18969 & ~n18971;
  assign n19246 = ~n18972 & ~n19245;
  assign n19247 = ~n19244 & n19246;
  assign n19248 = n71 & n12211;
  assign n19249 = n10329 & n12214;
  assign n19250 = n9836 & n12217;
  assign n19251 = n9830 & n13203;
  assign n19252 = ~n19249 & ~n19250;
  assign n19253 = ~n19248 & n19252;
  assign n19254 = ~n19251 & n19253;
  assign n19255 = ~pi5  & ~n19254;
  assign n19256 = pi5  & n19254;
  assign n19257 = ~n19255 & ~n19256;
  assign n19258 = n18965 & ~n18967;
  assign n19259 = ~n18968 & ~n19258;
  assign n19260 = ~n19257 & n19259;
  assign n19261 = n18961 & ~n18963;
  assign n19262 = ~n18964 & ~n19261;
  assign n19263 = n71 & n12214;
  assign n19264 = n10329 & n12217;
  assign n19265 = n9836 & n12220;
  assign n19266 = n9830 & n13187;
  assign n19267 = ~n19264 & ~n19265;
  assign n19268 = ~n19263 & n19267;
  assign n19269 = ~n19266 & n19268;
  assign n19270 = pi5  & n19269;
  assign n19271 = ~pi5  & ~n19269;
  assign n19272 = ~n19270 & ~n19271;
  assign n19273 = n19262 & ~n19272;
  assign n19274 = n18957 & ~n18959;
  assign n19275 = ~n18960 & ~n19274;
  assign n19276 = n71 & n12217;
  assign n19277 = n10329 & n12220;
  assign n19278 = n9836 & n12223;
  assign n19279 = n9830 & n13374;
  assign n19280 = ~n19277 & ~n19278;
  assign n19281 = ~n19276 & n19280;
  assign n19282 = ~n19279 & n19281;
  assign n19283 = pi5  & n19282;
  assign n19284 = ~pi5  & ~n19282;
  assign n19285 = ~n19283 & ~n19284;
  assign n19286 = n19275 & ~n19285;
  assign n19287 = n18953 & ~n18955;
  assign n19288 = ~n18956 & ~n19287;
  assign n19289 = n71 & n12220;
  assign n19290 = n10329 & n12223;
  assign n19291 = n9836 & n12226;
  assign n19292 = n9830 & n13392;
  assign n19293 = ~n19290 & ~n19291;
  assign n19294 = ~n19289 & n19293;
  assign n19295 = ~n19292 & n19294;
  assign n19296 = pi5  & n19295;
  assign n19297 = ~pi5  & ~n19295;
  assign n19298 = ~n19296 & ~n19297;
  assign n19299 = n19288 & ~n19298;
  assign n19300 = n71 & n12223;
  assign n19301 = n10329 & n12226;
  assign n19302 = n9836 & n12229;
  assign n19303 = n9830 & n13745;
  assign n19304 = ~n19301 & ~n19302;
  assign n19305 = ~n19300 & n19304;
  assign n19306 = ~n19303 & n19305;
  assign n19307 = ~pi5  & ~n19306;
  assign n19308 = pi5  & n19306;
  assign n19309 = ~n19307 & ~n19308;
  assign n19310 = n18949 & ~n18951;
  assign n19311 = ~n18952 & ~n19310;
  assign n19312 = ~n19309 & n19311;
  assign n19313 = n71 & n12226;
  assign n19314 = n10329 & n12229;
  assign n19315 = n9836 & n12232;
  assign n19316 = n9830 & n13530;
  assign n19317 = ~n19314 & ~n19315;
  assign n19318 = ~n19313 & n19317;
  assign n19319 = ~n19316 & n19318;
  assign n19320 = ~pi5  & ~n19319;
  assign n19321 = pi5  & n19319;
  assign n19322 = ~n19320 & ~n19321;
  assign n19323 = n18945 & ~n18947;
  assign n19324 = ~n18948 & ~n19323;
  assign n19325 = ~n19322 & n19324;
  assign n19326 = n71 & n12229;
  assign n19327 = n10329 & n12232;
  assign n19328 = n9836 & n12235;
  assign n19329 = n9830 & n13979;
  assign n19330 = ~n19327 & ~n19328;
  assign n19331 = ~n19326 & n19330;
  assign n19332 = ~n19329 & n19331;
  assign n19333 = ~pi5  & ~n19332;
  assign n19334 = pi5  & n19332;
  assign n19335 = ~n19333 & ~n19334;
  assign n19336 = n18941 & ~n18943;
  assign n19337 = ~n18944 & ~n19336;
  assign n19338 = ~n19335 & n19337;
  assign n19339 = n18937 & ~n18939;
  assign n19340 = ~n18940 & ~n19339;
  assign n19341 = n71 & n12232;
  assign n19342 = n10329 & n12235;
  assign n19343 = n9836 & n12238;
  assign n19344 = n9830 & n14116;
  assign n19345 = ~n19342 & ~n19343;
  assign n19346 = ~n19341 & n19345;
  assign n19347 = ~n19344 & n19346;
  assign n19348 = pi5  & n19347;
  assign n19349 = ~pi5  & ~n19347;
  assign n19350 = ~n19348 & ~n19349;
  assign n19351 = n19340 & ~n19350;
  assign n19352 = n18933 & ~n18935;
  assign n19353 = ~n18936 & ~n19352;
  assign n19354 = n71 & n12235;
  assign n19355 = n10329 & n12238;
  assign n19356 = n9836 & n12241;
  assign n19357 = n9830 & n13959;
  assign n19358 = ~n19355 & ~n19356;
  assign n19359 = ~n19354 & n19358;
  assign n19360 = ~n19357 & n19359;
  assign n19361 = pi5  & n19360;
  assign n19362 = ~pi5  & ~n19360;
  assign n19363 = ~n19361 & ~n19362;
  assign n19364 = n19353 & ~n19363;
  assign n19365 = n18929 & ~n18931;
  assign n19366 = ~n18932 & ~n19365;
  assign n19367 = n71 & n12238;
  assign n19368 = n10329 & n12241;
  assign n19369 = n9836 & n12244;
  assign n19370 = n9830 & n14229;
  assign n19371 = ~n19368 & ~n19369;
  assign n19372 = ~n19367 & n19371;
  assign n19373 = ~n19370 & n19372;
  assign n19374 = pi5  & n19373;
  assign n19375 = ~pi5  & ~n19373;
  assign n19376 = ~n19374 & ~n19375;
  assign n19377 = n19366 & ~n19376;
  assign n19378 = n71 & n12241;
  assign n19379 = n10329 & n12244;
  assign n19380 = n9836 & n12247;
  assign n19381 = n9830 & n14515;
  assign n19382 = ~n19379 & ~n19380;
  assign n19383 = ~n19378 & n19382;
  assign n19384 = ~n19381 & n19383;
  assign n19385 = ~pi5  & ~n19384;
  assign n19386 = pi5  & n19384;
  assign n19387 = ~n19385 & ~n19386;
  assign n19388 = n18925 & ~n18927;
  assign n19389 = ~n18928 & ~n19388;
  assign n19390 = ~n19387 & n19389;
  assign n19391 = n71 & n12244;
  assign n19392 = n10329 & n12247;
  assign n19393 = n9836 & n12250;
  assign n19394 = n9830 & n14527;
  assign n19395 = ~n19392 & ~n19393;
  assign n19396 = ~n19391 & n19395;
  assign n19397 = ~n19394 & n19396;
  assign n19398 = ~pi5  & ~n19397;
  assign n19399 = pi5  & n19397;
  assign n19400 = ~n19398 & ~n19399;
  assign n19401 = n18921 & ~n18923;
  assign n19402 = ~n18924 & ~n19401;
  assign n19403 = ~n19400 & n19402;
  assign n19404 = n71 & n12247;
  assign n19405 = n10329 & n12250;
  assign n19406 = n9836 & n12253;
  assign n19407 = n9830 & n14207;
  assign n19408 = ~n19405 & ~n19406;
  assign n19409 = ~n19404 & n19408;
  assign n19410 = ~n19407 & n19409;
  assign n19411 = ~pi5  & ~n19410;
  assign n19412 = pi5  & n19410;
  assign n19413 = ~n19411 & ~n19412;
  assign n19414 = n18917 & ~n18919;
  assign n19415 = ~n18920 & ~n19414;
  assign n19416 = ~n19413 & n19415;
  assign n19417 = n18913 & ~n18915;
  assign n19418 = ~n18916 & ~n19417;
  assign n19419 = n71 & n12250;
  assign n19420 = n10329 & n12253;
  assign n19421 = n9836 & n12256;
  assign n19422 = n9830 & n14559;
  assign n19423 = ~n19420 & ~n19421;
  assign n19424 = ~n19419 & n19423;
  assign n19425 = ~n19422 & n19424;
  assign n19426 = pi5  & n19425;
  assign n19427 = ~pi5  & ~n19425;
  assign n19428 = ~n19426 & ~n19427;
  assign n19429 = n19418 & ~n19428;
  assign n19430 = n18909 & ~n18911;
  assign n19431 = ~n18912 & ~n19430;
  assign n19432 = n71 & n12253;
  assign n19433 = n10329 & n12256;
  assign n19434 = n9836 & n12259;
  assign n19435 = n9830 & n14584;
  assign n19436 = ~n19433 & ~n19434;
  assign n19437 = ~n19432 & n19436;
  assign n19438 = ~n19435 & n19437;
  assign n19439 = pi5  & n19438;
  assign n19440 = ~pi5  & ~n19438;
  assign n19441 = ~n19439 & ~n19440;
  assign n19442 = n19431 & ~n19441;
  assign n19443 = n18905 & ~n18907;
  assign n19444 = ~n18908 & ~n19443;
  assign n19445 = n71 & n12256;
  assign n19446 = n10329 & n12259;
  assign n19447 = n9836 & n12262;
  assign n19448 = n9830 & n14608;
  assign n19449 = ~n19446 & ~n19447;
  assign n19450 = ~n19445 & n19449;
  assign n19451 = ~n19448 & n19450;
  assign n19452 = pi5  & n19451;
  assign n19453 = ~pi5  & ~n19451;
  assign n19454 = ~n19452 & ~n19453;
  assign n19455 = n19444 & ~n19454;
  assign n19456 = n71 & n12259;
  assign n19457 = n10329 & n12262;
  assign n19458 = n9836 & n12265;
  assign n19459 = n9830 & n14637;
  assign n19460 = ~n19457 & ~n19458;
  assign n19461 = ~n19456 & n19460;
  assign n19462 = ~n19459 & n19461;
  assign n19463 = ~pi5  & ~n19462;
  assign n19464 = pi5  & n19462;
  assign n19465 = ~n19463 & ~n19464;
  assign n19466 = n18901 & ~n18903;
  assign n19467 = ~n18904 & ~n19466;
  assign n19468 = ~n19465 & n19467;
  assign n19469 = n71 & n12262;
  assign n19470 = n10329 & n12265;
  assign n19471 = n9836 & n12268;
  assign n19472 = n9830 & n14691;
  assign n19473 = ~n19470 & ~n19471;
  assign n19474 = ~n19469 & n19473;
  assign n19475 = ~n19472 & n19474;
  assign n19476 = pi5  & n19475;
  assign n19477 = ~pi5  & ~n19475;
  assign n19478 = ~n19476 & ~n19477;
  assign n19479 = n18897 & ~n18899;
  assign n19480 = ~n18900 & ~n19479;
  assign n19481 = ~n19478 & n19480;
  assign n19482 = n71 & n12265;
  assign n19483 = n10329 & n12268;
  assign n19484 = n9836 & n12271;
  assign n19485 = n9830 & n14728;
  assign n19486 = ~n19483 & ~n19484;
  assign n19487 = ~n19482 & n19486;
  assign n19488 = ~n19485 & n19487;
  assign n19489 = ~pi5  & ~n19488;
  assign n19490 = pi5  & n19488;
  assign n19491 = ~n19489 & ~n19490;
  assign n19492 = pi8  & ~n18877;
  assign n19493 = n18884 & ~n19492;
  assign n19494 = ~n18884 & n19492;
  assign n19495 = ~n19493 & ~n19494;
  assign n19496 = ~n19491 & n19495;
  assign n19497 = n71 & n12268;
  assign n19498 = n10329 & n12271;
  assign n19499 = n9836 & n12274;
  assign n19500 = n9830 & n14771;
  assign n19501 = ~n19498 & ~n19499;
  assign n19502 = ~n19497 & n19501;
  assign n19503 = ~n19500 & n19502;
  assign n19504 = pi5  & n19503;
  assign n19505 = ~pi5  & ~n19503;
  assign n19506 = ~n19504 & ~n19505;
  assign n19507 = n18871 & ~n18876;
  assign n19508 = ~n18877 & ~n19507;
  assign n19509 = ~n19506 & n19508;
  assign n19510 = n67 & n12281;
  assign n19511 = pi5  & n19510;
  assign n19512 = n71 & n12279;
  assign n19513 = n10329 & n12281;
  assign n19514 = n9830 & ~n14833;
  assign n19515 = ~n19512 & ~n19513;
  assign n19516 = ~n19514 & n19515;
  assign n19517 = ~n19511 & n19516;
  assign n19518 = n71 & n12274;
  assign n19519 = n10329 & n12279;
  assign n19520 = n9836 & n12281;
  assign n19521 = n9830 & ~n14876;
  assign n19522 = ~n19519 & ~n19520;
  assign n19523 = ~n19518 & n19522;
  assign n19524 = ~n19521 & n19523;
  assign n19525 = pi5  & n19517;
  assign n19526 = n19524 & n19525;
  assign n19527 = n18870 & n19526;
  assign n19528 = n71 & n12271;
  assign n19529 = n10329 & n12274;
  assign n19530 = n9836 & n12279;
  assign n19531 = n9830 & n14795;
  assign n19532 = ~n19529 & ~n19530;
  assign n19533 = ~n19528 & n19532;
  assign n19534 = ~n19531 & n19533;
  assign n19535 = pi5  & n19534;
  assign n19536 = ~pi5  & ~n19534;
  assign n19537 = ~n19535 & ~n19536;
  assign n19538 = ~n18870 & ~n19526;
  assign n19539 = ~n19527 & ~n19538;
  assign n19540 = ~n19537 & n19539;
  assign n19541 = ~n19527 & ~n19540;
  assign n19542 = n19506 & ~n19508;
  assign n19543 = ~n19509 & ~n19542;
  assign n19544 = ~n19541 & n19543;
  assign n19545 = ~n19509 & ~n19544;
  assign n19546 = n19491 & ~n19495;
  assign n19547 = ~n19496 & ~n19546;
  assign n19548 = ~n19545 & n19547;
  assign n19549 = ~n19496 & ~n19548;
  assign n19550 = n19478 & ~n19480;
  assign n19551 = ~n19481 & ~n19550;
  assign n19552 = ~n19549 & n19551;
  assign n19553 = ~n19481 & ~n19552;
  assign n19554 = n19465 & ~n19467;
  assign n19555 = ~n19468 & ~n19554;
  assign n19556 = ~n19553 & n19555;
  assign n19557 = ~n19468 & ~n19556;
  assign n19558 = ~n19444 & n19454;
  assign n19559 = ~n19455 & ~n19558;
  assign n19560 = ~n19557 & n19559;
  assign n19561 = ~n19455 & ~n19560;
  assign n19562 = ~n19431 & n19441;
  assign n19563 = ~n19442 & ~n19562;
  assign n19564 = ~n19561 & n19563;
  assign n19565 = ~n19442 & ~n19564;
  assign n19566 = ~n19418 & n19428;
  assign n19567 = ~n19429 & ~n19566;
  assign n19568 = ~n19565 & n19567;
  assign n19569 = ~n19429 & ~n19568;
  assign n19570 = n19413 & ~n19415;
  assign n19571 = ~n19416 & ~n19570;
  assign n19572 = ~n19569 & n19571;
  assign n19573 = ~n19416 & ~n19572;
  assign n19574 = n19400 & ~n19402;
  assign n19575 = ~n19403 & ~n19574;
  assign n19576 = ~n19573 & n19575;
  assign n19577 = ~n19403 & ~n19576;
  assign n19578 = n19387 & ~n19389;
  assign n19579 = ~n19390 & ~n19578;
  assign n19580 = ~n19577 & n19579;
  assign n19581 = ~n19390 & ~n19580;
  assign n19582 = ~n19366 & n19376;
  assign n19583 = ~n19377 & ~n19582;
  assign n19584 = ~n19581 & n19583;
  assign n19585 = ~n19377 & ~n19584;
  assign n19586 = ~n19353 & n19363;
  assign n19587 = ~n19364 & ~n19586;
  assign n19588 = ~n19585 & n19587;
  assign n19589 = ~n19364 & ~n19588;
  assign n19590 = ~n19340 & n19350;
  assign n19591 = ~n19351 & ~n19590;
  assign n19592 = ~n19589 & n19591;
  assign n19593 = ~n19351 & ~n19592;
  assign n19594 = n19335 & ~n19337;
  assign n19595 = ~n19338 & ~n19594;
  assign n19596 = ~n19593 & n19595;
  assign n19597 = ~n19338 & ~n19596;
  assign n19598 = n19322 & ~n19324;
  assign n19599 = ~n19325 & ~n19598;
  assign n19600 = ~n19597 & n19599;
  assign n19601 = ~n19325 & ~n19600;
  assign n19602 = n19309 & ~n19311;
  assign n19603 = ~n19312 & ~n19602;
  assign n19604 = ~n19601 & n19603;
  assign n19605 = ~n19312 & ~n19604;
  assign n19606 = ~n19288 & n19298;
  assign n19607 = ~n19299 & ~n19606;
  assign n19608 = ~n19605 & n19607;
  assign n19609 = ~n19299 & ~n19608;
  assign n19610 = ~n19275 & n19285;
  assign n19611 = ~n19286 & ~n19610;
  assign n19612 = ~n19609 & n19611;
  assign n19613 = ~n19286 & ~n19612;
  assign n19614 = ~n19262 & n19272;
  assign n19615 = ~n19273 & ~n19614;
  assign n19616 = ~n19613 & n19615;
  assign n19617 = ~n19273 & ~n19616;
  assign n19618 = n19257 & ~n19259;
  assign n19619 = ~n19260 & ~n19618;
  assign n19620 = ~n19617 & n19619;
  assign n19621 = ~n19260 & ~n19620;
  assign n19622 = n19244 & ~n19246;
  assign n19623 = ~n19247 & ~n19622;
  assign n19624 = ~n19621 & n19623;
  assign n19625 = ~n19247 & ~n19624;
  assign n19626 = n19231 & ~n19233;
  assign n19627 = ~n19234 & ~n19626;
  assign n19628 = ~n19625 & n19627;
  assign n19629 = ~n19234 & ~n19628;
  assign n19630 = ~n19210 & n19220;
  assign n19631 = ~n19221 & ~n19630;
  assign n19632 = ~n19629 & n19631;
  assign n19633 = ~n19221 & ~n19632;
  assign n19634 = ~n19197 & n19207;
  assign n19635 = ~n19208 & ~n19634;
  assign n19636 = ~n19633 & n19635;
  assign n19637 = ~n19208 & ~n19636;
  assign n19638 = n19192 & ~n19194;
  assign n19639 = ~n19195 & ~n19638;
  assign n19640 = ~n19637 & n19639;
  assign n19641 = ~n19195 & ~n19640;
  assign n19642 = n19179 & ~n19181;
  assign n19643 = ~n19182 & ~n19642;
  assign n19644 = ~n19641 & n19643;
  assign n19645 = ~n19182 & ~n19644;
  assign n19646 = n19166 & ~n19168;
  assign n19647 = ~n19169 & ~n19646;
  assign n19648 = ~n19645 & n19647;
  assign n19649 = ~n19169 & ~n19648;
  assign n19650 = n19153 & ~n19155;
  assign n19651 = ~n19156 & ~n19650;
  assign n19652 = ~n19649 & n19651;
  assign n19653 = ~n19156 & ~n19652;
  assign n19654 = n19140 & ~n19142;
  assign n19655 = ~n19143 & ~n19654;
  assign n19656 = ~n19653 & n19655;
  assign n19657 = ~n19143 & ~n19656;
  assign n19658 = n19127 & ~n19129;
  assign n19659 = ~n19130 & ~n19658;
  assign n19660 = ~n19657 & n19659;
  assign n19661 = ~n19130 & ~n19660;
  assign n19662 = n19114 & ~n19116;
  assign n19663 = ~n19117 & ~n19662;
  assign n19664 = ~n19661 & n19663;
  assign n19665 = ~n19117 & ~n19664;
  assign n19666 = n19101 & ~n19103;
  assign n19667 = ~n19104 & ~n19666;
  assign n19668 = ~n19665 & n19667;
  assign n19669 = ~n19104 & ~n19668;
  assign n19670 = n19088 & ~n19090;
  assign n19671 = ~n19091 & ~n19670;
  assign n19672 = ~n19669 & n19671;
  assign n19673 = ~n19091 & ~n19672;
  assign n19674 = n19069 & ~n19071;
  assign n19675 = ~n19072 & ~n19674;
  assign n19676 = ~n19673 & n19675;
  assign n19677 = n19673 & ~n19675;
  assign n19678 = ~n19676 & ~n19677;
  assign n19679 = n19669 & ~n19671;
  assign n19680 = ~n19672 & ~n19679;
  assign n19681 = n10884 & n13007;
  assign n19682 = n10883 & n12172;
  assign n19683 = ~n11476 & n12165;
  assign n19684 = ~n12163 & ~n19063;
  assign n19685 = ~n19683 & n19684;
  assign n19686 = ~n19682 & ~n19685;
  assign n19687 = ~n19681 & n19686;
  assign n19688 = pi2  & n19687;
  assign n19689 = ~pi2  & ~n19687;
  assign n19690 = ~n19688 & ~n19689;
  assign n19691 = n19680 & ~n19690;
  assign n19692 = n19665 & ~n19667;
  assign n19693 = ~n19668 & ~n19692;
  assign n19694 = n11476 & n12166;
  assign n19695 = n11463 & n12172;
  assign n19696 = n10883 & n12168;
  assign n19697 = n10884 & n13106;
  assign n19698 = ~n19694 & ~n19696;
  assign n19699 = ~n19695 & n19698;
  assign n19700 = ~n19697 & n19699;
  assign n19701 = pi2  & n19700;
  assign n19702 = ~pi2  & ~n19700;
  assign n19703 = ~n19701 & ~n19702;
  assign n19704 = n19693 & ~n19703;
  assign n19705 = n19661 & ~n19663;
  assign n19706 = ~n19664 & ~n19705;
  assign n19707 = n11476 & n12172;
  assign n19708 = n11463 & n12168;
  assign n19709 = n10883 & n12175;
  assign n19710 = n10884 & n12939;
  assign n19711 = ~n19708 & ~n19709;
  assign n19712 = ~n19707 & n19711;
  assign n19713 = ~n19710 & n19712;
  assign n19714 = pi2  & n19713;
  assign n19715 = ~pi2  & ~n19713;
  assign n19716 = ~n19714 & ~n19715;
  assign n19717 = n19706 & ~n19716;
  assign n19718 = n19657 & ~n19659;
  assign n19719 = ~n19660 & ~n19718;
  assign n19720 = n11476 & n12168;
  assign n19721 = n11463 & n12175;
  assign n19722 = n10883 & n12178;
  assign n19723 = n10884 & n12862;
  assign n19724 = ~n19721 & ~n19722;
  assign n19725 = ~n19720 & n19724;
  assign n19726 = ~n19723 & n19725;
  assign n19727 = pi2  & n19726;
  assign n19728 = ~pi2  & ~n19726;
  assign n19729 = ~n19727 & ~n19728;
  assign n19730 = n19719 & ~n19729;
  assign n19731 = n19653 & ~n19655;
  assign n19732 = ~n19656 & ~n19731;
  assign n19733 = n11476 & n12175;
  assign n19734 = n11463 & n12178;
  assign n19735 = n10883 & n12181;
  assign n19736 = n10884 & n12961;
  assign n19737 = ~n19734 & ~n19735;
  assign n19738 = ~n19733 & n19737;
  assign n19739 = ~n19736 & n19738;
  assign n19740 = pi2  & n19739;
  assign n19741 = ~pi2  & ~n19739;
  assign n19742 = ~n19740 & ~n19741;
  assign n19743 = n19732 & ~n19742;
  assign n19744 = n19649 & ~n19651;
  assign n19745 = ~n19652 & ~n19744;
  assign n19746 = n11476 & n12178;
  assign n19747 = n11463 & n12181;
  assign n19748 = n10883 & n12184;
  assign n19749 = n10884 & n12880;
  assign n19750 = ~n19747 & ~n19748;
  assign n19751 = ~n19746 & n19750;
  assign n19752 = ~n19749 & n19751;
  assign n19753 = pi2  & n19752;
  assign n19754 = ~pi2  & ~n19752;
  assign n19755 = ~n19753 & ~n19754;
  assign n19756 = n19745 & ~n19755;
  assign n19757 = n19645 & ~n19647;
  assign n19758 = ~n19648 & ~n19757;
  assign n19759 = n11476 & n12181;
  assign n19760 = n11463 & n12184;
  assign n19761 = n10883 & n12187;
  assign n19762 = n10884 & n12608;
  assign n19763 = ~n19760 & ~n19761;
  assign n19764 = ~n19759 & n19763;
  assign n19765 = ~n19762 & n19764;
  assign n19766 = pi2  & n19765;
  assign n19767 = ~pi2  & ~n19765;
  assign n19768 = ~n19766 & ~n19767;
  assign n19769 = n19758 & ~n19768;
  assign n19770 = n19641 & ~n19643;
  assign n19771 = ~n19644 & ~n19770;
  assign n19772 = n11476 & n12184;
  assign n19773 = n11463 & n12187;
  assign n19774 = n10883 & n12190;
  assign n19775 = n10884 & n12845;
  assign n19776 = ~n19773 & ~n19774;
  assign n19777 = ~n19772 & n19776;
  assign n19778 = ~n19775 & n19777;
  assign n19779 = pi2  & n19778;
  assign n19780 = ~pi2  & ~n19778;
  assign n19781 = ~n19779 & ~n19780;
  assign n19782 = n19771 & ~n19781;
  assign n19783 = n19637 & ~n19639;
  assign n19784 = ~n19640 & ~n19783;
  assign n19785 = n11476 & n12187;
  assign n19786 = n11463 & n12190;
  assign n19787 = n10883 & n12193;
  assign n19788 = n10884 & n12921;
  assign n19789 = ~n19786 & ~n19787;
  assign n19790 = ~n19785 & n19789;
  assign n19791 = ~n19788 & n19790;
  assign n19792 = pi2  & n19791;
  assign n19793 = ~pi2  & ~n19791;
  assign n19794 = ~n19792 & ~n19793;
  assign n19795 = n19784 & ~n19794;
  assign n19796 = ~n19784 & n19794;
  assign n19797 = ~n19795 & ~n19796;
  assign n19798 = n19633 & ~n19635;
  assign n19799 = ~n19636 & ~n19798;
  assign n19800 = n19629 & ~n19631;
  assign n19801 = ~n19632 & ~n19800;
  assign n19802 = n11476 & n12196;
  assign n19803 = n11463 & n12199;
  assign n19804 = n10883 & n12202;
  assign n19805 = n10884 & n12578;
  assign n19806 = ~n19803 & ~n19804;
  assign n19807 = ~n19802 & n19806;
  assign n19808 = ~n19805 & n19807;
  assign n19809 = pi2  & n19808;
  assign n19810 = ~pi2  & ~n19808;
  assign n19811 = ~n19809 & ~n19810;
  assign n19812 = n11476 & n12199;
  assign n19813 = n11463 & n12202;
  assign n19814 = n10883 & n12205;
  assign n19815 = n10884 & n12683;
  assign n19816 = ~n19813 & ~n19814;
  assign n19817 = ~n19812 & n19816;
  assign n19818 = ~n19815 & n19817;
  assign n19819 = pi2  & n19818;
  assign n19820 = ~pi2  & ~n19818;
  assign n19821 = ~n19819 & ~n19820;
  assign n19822 = n11476 & n12202;
  assign n19823 = n11463 & n12205;
  assign n19824 = n10883 & n12208;
  assign n19825 = n10884 & n12701;
  assign n19826 = ~n19823 & ~n19824;
  assign n19827 = ~n19822 & n19826;
  assign n19828 = ~n19825 & n19827;
  assign n19829 = pi2  & n19828;
  assign n19830 = ~pi2  & ~n19828;
  assign n19831 = ~n19829 & ~n19830;
  assign n19832 = n19613 & ~n19615;
  assign n19833 = ~n19616 & ~n19832;
  assign n19834 = n19609 & ~n19611;
  assign n19835 = ~n19612 & ~n19834;
  assign n19836 = n19605 & ~n19607;
  assign n19837 = ~n19608 & ~n19836;
  assign n19838 = n11476 & n12214;
  assign n19839 = n11463 & n12217;
  assign n19840 = n10883 & n12220;
  assign n19841 = n10884 & n13187;
  assign n19842 = ~n19839 & ~n19840;
  assign n19843 = ~n19838 & n19842;
  assign n19844 = ~n19841 & n19843;
  assign n19845 = pi2  & n19844;
  assign n19846 = ~pi2  & ~n19844;
  assign n19847 = ~n19845 & ~n19846;
  assign n19848 = n11476 & n12217;
  assign n19849 = n11463 & n12220;
  assign n19850 = n10883 & n12223;
  assign n19851 = n10884 & n13374;
  assign n19852 = ~n19849 & ~n19850;
  assign n19853 = ~n19848 & n19852;
  assign n19854 = ~n19851 & n19853;
  assign n19855 = pi2  & n19854;
  assign n19856 = ~pi2  & ~n19854;
  assign n19857 = ~n19855 & ~n19856;
  assign n19858 = n11476 & n12220;
  assign n19859 = n11463 & n12223;
  assign n19860 = n10883 & n12226;
  assign n19861 = n10884 & n13392;
  assign n19862 = ~n19859 & ~n19860;
  assign n19863 = ~n19858 & n19862;
  assign n19864 = ~n19861 & n19863;
  assign n19865 = pi2  & n19864;
  assign n19866 = ~pi2  & ~n19864;
  assign n19867 = ~n19865 & ~n19866;
  assign n19868 = n19589 & ~n19591;
  assign n19869 = ~n19592 & ~n19868;
  assign n19870 = n19585 & ~n19587;
  assign n19871 = ~n19588 & ~n19870;
  assign n19872 = n19581 & ~n19583;
  assign n19873 = ~n19584 & ~n19872;
  assign n19874 = n11476 & n12232;
  assign n19875 = n11463 & n12235;
  assign n19876 = n10883 & n12238;
  assign n19877 = n10884 & n14116;
  assign n19878 = ~n19875 & ~n19876;
  assign n19879 = ~n19874 & n19878;
  assign n19880 = ~n19877 & n19879;
  assign n19881 = pi2  & n19880;
  assign n19882 = ~pi2  & ~n19880;
  assign n19883 = ~n19881 & ~n19882;
  assign n19884 = n11476 & n12235;
  assign n19885 = n11463 & n12238;
  assign n19886 = n10883 & n12241;
  assign n19887 = n10884 & n13959;
  assign n19888 = ~n19885 & ~n19886;
  assign n19889 = ~n19884 & n19888;
  assign n19890 = ~n19887 & n19889;
  assign n19891 = pi2  & n19890;
  assign n19892 = ~pi2  & ~n19890;
  assign n19893 = ~n19891 & ~n19892;
  assign n19894 = n11476 & n12238;
  assign n19895 = n11463 & n12241;
  assign n19896 = n10883 & n12244;
  assign n19897 = n10884 & n14229;
  assign n19898 = ~n19895 & ~n19896;
  assign n19899 = ~n19894 & n19898;
  assign n19900 = ~n19897 & n19899;
  assign n19901 = pi2  & n19900;
  assign n19902 = ~pi2  & ~n19900;
  assign n19903 = ~n19901 & ~n19902;
  assign n19904 = n19565 & ~n19567;
  assign n19905 = ~n19568 & ~n19904;
  assign n19906 = n19561 & ~n19563;
  assign n19907 = ~n19564 & ~n19906;
  assign n19908 = n19557 & ~n19559;
  assign n19909 = ~n19560 & ~n19908;
  assign n19910 = n11476 & n12250;
  assign n19911 = n11463 & n12253;
  assign n19912 = n10883 & n12256;
  assign n19913 = n10884 & n14559;
  assign n19914 = ~n19911 & ~n19912;
  assign n19915 = ~n19910 & n19914;
  assign n19916 = ~n19913 & n19915;
  assign n19917 = pi2  & n19916;
  assign n19918 = ~pi2  & ~n19916;
  assign n19919 = ~n19917 & ~n19918;
  assign n19920 = n11476 & n12253;
  assign n19921 = n11463 & n12256;
  assign n19922 = n10883 & n12259;
  assign n19923 = n10884 & n14584;
  assign n19924 = ~n19921 & ~n19922;
  assign n19925 = ~n19920 & n19924;
  assign n19926 = ~n19923 & n19925;
  assign n19927 = pi2  & n19926;
  assign n19928 = ~pi2  & ~n19926;
  assign n19929 = ~n19927 & ~n19928;
  assign n19930 = n11476 & n12256;
  assign n19931 = n11463 & n12259;
  assign n19932 = n10883 & n12262;
  assign n19933 = n10884 & n14608;
  assign n19934 = ~n19931 & ~n19932;
  assign n19935 = ~n19930 & n19934;
  assign n19936 = ~n19933 & n19935;
  assign n19937 = pi2  & n19936;
  assign n19938 = ~pi2  & ~n19936;
  assign n19939 = ~n19937 & ~n19938;
  assign n19940 = n19541 & ~n19543;
  assign n19941 = ~n19544 & ~n19940;
  assign n19942 = n11476 & n12262;
  assign n19943 = n11463 & n12265;
  assign n19944 = n10883 & n12268;
  assign n19945 = n10884 & n14691;
  assign n19946 = ~n19943 & ~n19944;
  assign n19947 = ~n19942 & n19946;
  assign n19948 = ~n19945 & n19947;
  assign n19949 = pi2  & n19948;
  assign n19950 = ~pi2  & ~n19948;
  assign n19951 = ~n19949 & ~n19950;
  assign n19952 = pi5  & ~n19517;
  assign n19953 = n19524 & ~n19952;
  assign n19954 = ~n19524 & n19952;
  assign n19955 = ~n19953 & ~n19954;
  assign n19956 = n11476 & n12274;
  assign n19957 = ~n12274 & n14833;
  assign n19958 = n10884 & ~n19957;
  assign n19959 = pi1  & ~n10884;
  assign n19960 = n12279 & n19959;
  assign n19961 = pi2  & ~n12281;
  assign n19962 = ~n19960 & n19961;
  assign n19963 = ~n19956 & n19962;
  assign n19964 = ~n19958 & n19963;
  assign n19965 = ~n19510 & ~n19964;
  assign n19966 = n11476 & n12271;
  assign n19967 = n11463 & n12274;
  assign n19968 = n10883 & n12279;
  assign n19969 = n10884 & n14795;
  assign n19970 = ~n19967 & ~n19968;
  assign n19971 = ~n19966 & n19970;
  assign n19972 = ~n19969 & n19971;
  assign n19973 = ~pi2  & ~n19972;
  assign n19974 = pi2  & n19972;
  assign n19975 = ~n19973 & ~n19974;
  assign n19976 = ~n19965 & ~n19975;
  assign n19977 = n11476 & n12268;
  assign n19978 = n11463 & n12271;
  assign n19979 = n10883 & n12274;
  assign n19980 = n10884 & n14771;
  assign n19981 = ~n19978 & ~n19979;
  assign n19982 = ~n19977 & n19981;
  assign n19983 = ~n19980 & n19982;
  assign n19984 = pi2  & n19983;
  assign n19985 = ~pi2  & ~n19983;
  assign n19986 = ~n19984 & ~n19985;
  assign n19987 = n19976 & ~n19986;
  assign n19988 = ~n19976 & n19986;
  assign n19989 = n19511 & ~n19516;
  assign n19990 = ~n19517 & ~n19989;
  assign n19991 = ~n19988 & n19990;
  assign n19992 = ~n19987 & ~n19991;
  assign n19993 = n19955 & ~n19992;
  assign n19994 = ~n19955 & n19992;
  assign n19995 = n11476 & n12265;
  assign n19996 = n11463 & n12268;
  assign n19997 = n10883 & n12271;
  assign n19998 = n10884 & n14728;
  assign n19999 = ~n19996 & ~n19997;
  assign n20000 = ~n19995 & n19999;
  assign n20001 = ~n19998 & n20000;
  assign n20002 = pi2  & ~n20001;
  assign n20003 = ~pi2  & n20001;
  assign n20004 = ~n20002 & ~n20003;
  assign n20005 = ~n19994 & n20004;
  assign n20006 = ~n19993 & ~n20005;
  assign n20007 = ~n19951 & ~n20006;
  assign n20008 = n19951 & n20006;
  assign n20009 = n19537 & ~n19539;
  assign n20010 = ~n19540 & ~n20009;
  assign n20011 = ~n20008 & n20010;
  assign n20012 = ~n20007 & ~n20011;
  assign n20013 = n19941 & ~n20012;
  assign n20014 = ~n19941 & n20012;
  assign n20015 = n11476 & n12259;
  assign n20016 = n11463 & n12262;
  assign n20017 = n10883 & n12265;
  assign n20018 = n10884 & n14637;
  assign n20019 = ~n20016 & ~n20017;
  assign n20020 = ~n20015 & n20019;
  assign n20021 = ~n20018 & n20020;
  assign n20022 = pi2  & ~n20021;
  assign n20023 = ~pi2  & n20021;
  assign n20024 = ~n20022 & ~n20023;
  assign n20025 = ~n20014 & n20024;
  assign n20026 = ~n20013 & ~n20025;
  assign n20027 = ~n19939 & ~n20026;
  assign n20028 = n19939 & n20026;
  assign n20029 = n19545 & ~n19547;
  assign n20030 = ~n19548 & ~n20029;
  assign n20031 = ~n20028 & n20030;
  assign n20032 = ~n20027 & ~n20031;
  assign n20033 = ~n19929 & ~n20032;
  assign n20034 = n19929 & n20032;
  assign n20035 = n19549 & ~n19551;
  assign n20036 = ~n19552 & ~n20035;
  assign n20037 = ~n20034 & n20036;
  assign n20038 = ~n20033 & ~n20037;
  assign n20039 = ~n19919 & ~n20038;
  assign n20040 = n19919 & n20038;
  assign n20041 = n19553 & ~n19555;
  assign n20042 = ~n19556 & ~n20041;
  assign n20043 = ~n20040 & n20042;
  assign n20044 = ~n20039 & ~n20043;
  assign n20045 = n19909 & ~n20044;
  assign n20046 = ~n19909 & n20044;
  assign n20047 = n11476 & n12247;
  assign n20048 = n11463 & n12250;
  assign n20049 = n10883 & n12253;
  assign n20050 = n10884 & n14207;
  assign n20051 = ~n20048 & ~n20049;
  assign n20052 = ~n20047 & n20051;
  assign n20053 = ~n20050 & n20052;
  assign n20054 = pi2  & ~n20053;
  assign n20055 = ~pi2  & n20053;
  assign n20056 = ~n20054 & ~n20055;
  assign n20057 = ~n20046 & n20056;
  assign n20058 = ~n20045 & ~n20057;
  assign n20059 = n19907 & ~n20058;
  assign n20060 = ~n19907 & n20058;
  assign n20061 = n11476 & n12244;
  assign n20062 = n11463 & n12247;
  assign n20063 = n10883 & n12250;
  assign n20064 = n10884 & n14527;
  assign n20065 = ~n20062 & ~n20063;
  assign n20066 = ~n20061 & n20065;
  assign n20067 = ~n20064 & n20066;
  assign n20068 = pi2  & ~n20067;
  assign n20069 = ~pi2  & n20067;
  assign n20070 = ~n20068 & ~n20069;
  assign n20071 = ~n20060 & n20070;
  assign n20072 = ~n20059 & ~n20071;
  assign n20073 = n19905 & ~n20072;
  assign n20074 = ~n19905 & n20072;
  assign n20075 = n11476 & n12241;
  assign n20076 = n11463 & n12244;
  assign n20077 = n10883 & n12247;
  assign n20078 = n10884 & n14515;
  assign n20079 = ~n20076 & ~n20077;
  assign n20080 = ~n20075 & n20079;
  assign n20081 = ~n20078 & n20080;
  assign n20082 = pi2  & ~n20081;
  assign n20083 = ~pi2  & n20081;
  assign n20084 = ~n20082 & ~n20083;
  assign n20085 = ~n20074 & n20084;
  assign n20086 = ~n20073 & ~n20085;
  assign n20087 = ~n19903 & ~n20086;
  assign n20088 = n19903 & n20086;
  assign n20089 = n19569 & ~n19571;
  assign n20090 = ~n19572 & ~n20089;
  assign n20091 = ~n20088 & n20090;
  assign n20092 = ~n20087 & ~n20091;
  assign n20093 = ~n19893 & ~n20092;
  assign n20094 = n19893 & n20092;
  assign n20095 = n19573 & ~n19575;
  assign n20096 = ~n19576 & ~n20095;
  assign n20097 = ~n20094 & n20096;
  assign n20098 = ~n20093 & ~n20097;
  assign n20099 = ~n19883 & ~n20098;
  assign n20100 = n19883 & n20098;
  assign n20101 = n19577 & ~n19579;
  assign n20102 = ~n19580 & ~n20101;
  assign n20103 = ~n20100 & n20102;
  assign n20104 = ~n20099 & ~n20103;
  assign n20105 = n19873 & ~n20104;
  assign n20106 = ~n19873 & n20104;
  assign n20107 = n11476 & n12229;
  assign n20108 = n11463 & n12232;
  assign n20109 = n10883 & n12235;
  assign n20110 = n10884 & n13979;
  assign n20111 = ~n20108 & ~n20109;
  assign n20112 = ~n20107 & n20111;
  assign n20113 = ~n20110 & n20112;
  assign n20114 = pi2  & ~n20113;
  assign n20115 = ~pi2  & n20113;
  assign n20116 = ~n20114 & ~n20115;
  assign n20117 = ~n20106 & n20116;
  assign n20118 = ~n20105 & ~n20117;
  assign n20119 = n19871 & ~n20118;
  assign n20120 = ~n19871 & n20118;
  assign n20121 = n11476 & n12226;
  assign n20122 = n11463 & n12229;
  assign n20123 = n10883 & n12232;
  assign n20124 = n10884 & n13530;
  assign n20125 = ~n20122 & ~n20123;
  assign n20126 = ~n20121 & n20125;
  assign n20127 = ~n20124 & n20126;
  assign n20128 = pi2  & ~n20127;
  assign n20129 = ~pi2  & n20127;
  assign n20130 = ~n20128 & ~n20129;
  assign n20131 = ~n20120 & n20130;
  assign n20132 = ~n20119 & ~n20131;
  assign n20133 = n19869 & ~n20132;
  assign n20134 = ~n19869 & n20132;
  assign n20135 = n11476 & n12223;
  assign n20136 = n11463 & n12226;
  assign n20137 = n10883 & n12229;
  assign n20138 = n10884 & n13745;
  assign n20139 = ~n20136 & ~n20137;
  assign n20140 = ~n20135 & n20139;
  assign n20141 = ~n20138 & n20140;
  assign n20142 = pi2  & ~n20141;
  assign n20143 = ~pi2  & n20141;
  assign n20144 = ~n20142 & ~n20143;
  assign n20145 = ~n20134 & n20144;
  assign n20146 = ~n20133 & ~n20145;
  assign n20147 = ~n19867 & ~n20146;
  assign n20148 = n19867 & n20146;
  assign n20149 = n19593 & ~n19595;
  assign n20150 = ~n19596 & ~n20149;
  assign n20151 = ~n20148 & n20150;
  assign n20152 = ~n20147 & ~n20151;
  assign n20153 = ~n19857 & ~n20152;
  assign n20154 = n19857 & n20152;
  assign n20155 = n19597 & ~n19599;
  assign n20156 = ~n19600 & ~n20155;
  assign n20157 = ~n20154 & n20156;
  assign n20158 = ~n20153 & ~n20157;
  assign n20159 = ~n19847 & ~n20158;
  assign n20160 = n19847 & n20158;
  assign n20161 = n19601 & ~n19603;
  assign n20162 = ~n19604 & ~n20161;
  assign n20163 = ~n20160 & n20162;
  assign n20164 = ~n20159 & ~n20163;
  assign n20165 = n19837 & ~n20164;
  assign n20166 = ~n19837 & n20164;
  assign n20167 = n11476 & n12211;
  assign n20168 = n11463 & n12214;
  assign n20169 = n10883 & n12217;
  assign n20170 = n10884 & n13203;
  assign n20171 = ~n20168 & ~n20169;
  assign n20172 = ~n20167 & n20171;
  assign n20173 = ~n20170 & n20172;
  assign n20174 = pi2  & ~n20173;
  assign n20175 = ~pi2  & n20173;
  assign n20176 = ~n20174 & ~n20175;
  assign n20177 = ~n20166 & n20176;
  assign n20178 = ~n20165 & ~n20177;
  assign n20179 = n19835 & ~n20178;
  assign n20180 = ~n19835 & n20178;
  assign n20181 = n11476 & n12208;
  assign n20182 = n11463 & n12211;
  assign n20183 = n10883 & n12214;
  assign n20184 = n10884 & n12804;
  assign n20185 = ~n20182 & ~n20183;
  assign n20186 = ~n20181 & n20185;
  assign n20187 = ~n20184 & n20186;
  assign n20188 = pi2  & ~n20187;
  assign n20189 = ~pi2  & n20187;
  assign n20190 = ~n20188 & ~n20189;
  assign n20191 = ~n20180 & n20190;
  assign n20192 = ~n20179 & ~n20191;
  assign n20193 = n19833 & ~n20192;
  assign n20194 = ~n19833 & n20192;
  assign n20195 = n11476 & n12205;
  assign n20196 = n11463 & n12208;
  assign n20197 = n10883 & n12211;
  assign n20198 = n10884 & n13031;
  assign n20199 = ~n20196 & ~n20197;
  assign n20200 = ~n20195 & n20199;
  assign n20201 = ~n20198 & n20200;
  assign n20202 = pi2  & ~n20201;
  assign n20203 = ~pi2  & n20201;
  assign n20204 = ~n20202 & ~n20203;
  assign n20205 = ~n20194 & n20204;
  assign n20206 = ~n20193 & ~n20205;
  assign n20207 = ~n19831 & ~n20206;
  assign n20208 = n19831 & n20206;
  assign n20209 = n19617 & ~n19619;
  assign n20210 = ~n19620 & ~n20209;
  assign n20211 = ~n20208 & n20210;
  assign n20212 = ~n20207 & ~n20211;
  assign n20213 = ~n19821 & ~n20212;
  assign n20214 = n19821 & n20212;
  assign n20215 = n19621 & ~n19623;
  assign n20216 = ~n19624 & ~n20215;
  assign n20217 = ~n20214 & n20216;
  assign n20218 = ~n20213 & ~n20217;
  assign n20219 = ~n19811 & ~n20218;
  assign n20220 = n19811 & n20218;
  assign n20221 = n19625 & ~n19627;
  assign n20222 = ~n19628 & ~n20221;
  assign n20223 = ~n20220 & n20222;
  assign n20224 = ~n20219 & ~n20223;
  assign n20225 = n19801 & ~n20224;
  assign n20226 = ~n19801 & n20224;
  assign n20227 = n11476 & n12193;
  assign n20228 = n11463 & n12196;
  assign n20229 = n10883 & n12199;
  assign n20230 = n10884 & n12594;
  assign n20231 = ~n20228 & ~n20229;
  assign n20232 = ~n20227 & n20231;
  assign n20233 = ~n20230 & n20232;
  assign n20234 = pi2  & ~n20233;
  assign n20235 = ~pi2  & n20233;
  assign n20236 = ~n20234 & ~n20235;
  assign n20237 = ~n20226 & n20236;
  assign n20238 = ~n20225 & ~n20237;
  assign n20239 = n19799 & ~n20238;
  assign n20240 = ~n19799 & n20238;
  assign n20241 = n11476 & n12190;
  assign n20242 = n11463 & n12193;
  assign n20243 = n10883 & n12196;
  assign n20244 = n10884 & n12530;
  assign n20245 = ~n20242 & ~n20243;
  assign n20246 = ~n20241 & n20245;
  assign n20247 = ~n20244 & n20246;
  assign n20248 = pi2  & ~n20247;
  assign n20249 = ~pi2  & n20247;
  assign n20250 = ~n20248 & ~n20249;
  assign n20251 = ~n20240 & n20250;
  assign n20252 = ~n20239 & ~n20251;
  assign n20253 = n19797 & ~n20252;
  assign n20254 = ~n19795 & ~n20253;
  assign n20255 = ~n19771 & n19781;
  assign n20256 = ~n19782 & ~n20255;
  assign n20257 = ~n20254 & n20256;
  assign n20258 = ~n19782 & ~n20257;
  assign n20259 = ~n19758 & n19768;
  assign n20260 = ~n19769 & ~n20259;
  assign n20261 = ~n20258 & n20260;
  assign n20262 = ~n19769 & ~n20261;
  assign n20263 = ~n19745 & n19755;
  assign n20264 = ~n19756 & ~n20263;
  assign n20265 = ~n20262 & n20264;
  assign n20266 = ~n19756 & ~n20265;
  assign n20267 = ~n19732 & n19742;
  assign n20268 = ~n19743 & ~n20267;
  assign n20269 = ~n20266 & n20268;
  assign n20270 = ~n19743 & ~n20269;
  assign n20271 = ~n19719 & n19729;
  assign n20272 = ~n19730 & ~n20271;
  assign n20273 = ~n20270 & n20272;
  assign n20274 = ~n19730 & ~n20273;
  assign n20275 = ~n19706 & n19716;
  assign n20276 = ~n19717 & ~n20275;
  assign n20277 = ~n20274 & n20276;
  assign n20278 = ~n19717 & ~n20277;
  assign n20279 = ~n19693 & n19703;
  assign n20280 = ~n19704 & ~n20279;
  assign n20281 = ~n20278 & n20280;
  assign n20282 = ~n19704 & ~n20281;
  assign n20283 = ~n19680 & n19690;
  assign n20284 = ~n19691 & ~n20283;
  assign n20285 = ~n20282 & n20284;
  assign n20286 = ~n19691 & ~n20285;
  assign n20287 = n19678 & ~n20286;
  assign n20288 = ~n19676 & ~n20287;
  assign n20289 = n19078 & ~n20288;
  assign n20290 = ~n19076 & ~n20289;
  assign n20291 = n19047 & ~n20290;
  assign n20292 = ~n19045 & ~n20291;
  assign n20293 = n18464 & ~n20292;
  assign n20294 = ~n18462 & ~n20293;
  assign n20295 = n17912 & ~n17914;
  assign n20296 = ~n17915 & ~n20295;
  assign n20297 = ~n20294 & n20296;
  assign n20298 = ~n17915 & ~n20297;
  assign n20299 = n17401 & ~n17403;
  assign n20300 = ~n17404 & ~n20299;
  assign n20301 = ~n20298 & n20300;
  assign n20302 = ~n17404 & ~n20301;
  assign n20303 = n16925 & ~n20302;
  assign n20304 = ~n16923 & ~n20303;
  assign n20305 = n16475 & ~n16477;
  assign n20306 = ~n16478 & ~n20305;
  assign n20307 = ~n20304 & n20306;
  assign n20308 = ~n16478 & ~n20307;
  assign n20309 = n16066 & ~n16068;
  assign n20310 = ~n16069 & ~n20309;
  assign n20311 = ~n20308 & n20310;
  assign n20312 = ~n16069 & ~n20311;
  assign n20313 = n15692 & ~n20312;
  assign n20314 = ~n15690 & ~n20313;
  assign n20315 = n15345 & ~n15347;
  assign n20316 = ~n15348 & ~n20315;
  assign n20317 = ~n20314 & n20316;
  assign n20318 = ~n15348 & ~n20317;
  assign n20319 = n15198 & ~n15200;
  assign n20320 = ~n15201 & ~n20319;
  assign n20321 = ~n20318 & n20320;
  assign n20322 = ~n15201 & ~n20321;
  assign n20323 = n15052 & ~n20322;
  assign n20324 = ~n15050 & ~n20323;
  assign n20325 = n14479 & ~n14481;
  assign n20326 = ~n14482 & ~n20325;
  assign n20327 = ~n20324 & n20326;
  assign n20328 = ~n14482 & ~n20327;
  assign n20329 = n14349 & ~n14351;
  assign n20330 = ~n14352 & ~n20329;
  assign n20331 = ~n20328 & n20330;
  assign n20332 = ~n14352 & ~n20331;
  assign n20333 = n14083 & ~n20332;
  assign n20334 = ~n14081 & ~n20333;
  assign n20335 = n13851 & ~n13853;
  assign n20336 = ~n13854 & ~n20335;
  assign n20337 = ~n20334 & n20336;
  assign n20338 = ~n13854 & ~n20337;
  assign n20339 = n13722 & ~n13724;
  assign n20340 = ~n13725 & ~n20339;
  assign n20341 = ~n20338 & n20340;
  assign n20342 = ~n13725 & ~n20341;
  assign n20343 = n13627 & ~n20342;
  assign n20344 = ~n13625 & ~n20343;
  assign n20345 = n13277 & ~n13279;
  assign n20346 = ~n13280 & ~n20345;
  assign n20347 = ~n20344 & n20346;
  assign n20348 = ~n13280 & ~n20347;
  assign n20349 = n13024 & n13120;
  assign n20350 = ~n13121 & ~n20349;
  assign n20351 = ~n20348 & n20350;
  assign n20352 = ~n13121 & ~n20351;
  assign n20353 = n13022 & ~n20352;
  assign n20354 = ~n13022 & n20352;
  assign n20355 = ~n20353 & ~n20354;
  assign n20356 = n71 & n20355;
  assign n20357 = n20348 & ~n20350;
  assign n20358 = ~n20351 & ~n20357;
  assign n20359 = n10329 & n20358;
  assign n20360 = n20344 & ~n20346;
  assign n20361 = ~n20347 & ~n20360;
  assign n20362 = n9836 & n20361;
  assign n20363 = n20358 & n20361;
  assign n20364 = ~n13627 & n20342;
  assign n20365 = ~n20343 & ~n20364;
  assign n20366 = n20361 & n20365;
  assign n20367 = n20338 & ~n20340;
  assign n20368 = ~n20341 & ~n20367;
  assign n20369 = n20365 & n20368;
  assign n20370 = n20334 & ~n20336;
  assign n20371 = ~n20337 & ~n20370;
  assign n20372 = n20368 & n20371;
  assign n20373 = ~n14083 & n20332;
  assign n20374 = ~n20333 & ~n20373;
  assign n20375 = n20371 & n20374;
  assign n20376 = n20328 & ~n20330;
  assign n20377 = ~n20331 & ~n20376;
  assign n20378 = n20374 & n20377;
  assign n20379 = n20324 & ~n20326;
  assign n20380 = ~n20327 & ~n20379;
  assign n20381 = n20377 & n20380;
  assign n20382 = ~n15052 & n20322;
  assign n20383 = ~n20323 & ~n20382;
  assign n20384 = n20380 & n20383;
  assign n20385 = n20318 & ~n20320;
  assign n20386 = ~n20321 & ~n20385;
  assign n20387 = n20383 & n20386;
  assign n20388 = n20314 & ~n20316;
  assign n20389 = ~n20317 & ~n20388;
  assign n20390 = n20386 & n20389;
  assign n20391 = ~n15692 & n20312;
  assign n20392 = ~n20313 & ~n20391;
  assign n20393 = n20389 & n20392;
  assign n20394 = n20308 & ~n20310;
  assign n20395 = ~n20311 & ~n20394;
  assign n20396 = n20392 & n20395;
  assign n20397 = n20304 & ~n20306;
  assign n20398 = ~n20307 & ~n20397;
  assign n20399 = n20395 & n20398;
  assign n20400 = ~n16925 & n20302;
  assign n20401 = ~n20303 & ~n20400;
  assign n20402 = n20398 & n20401;
  assign n20403 = n20298 & ~n20300;
  assign n20404 = ~n20301 & ~n20403;
  assign n20405 = n20401 & n20404;
  assign n20406 = n20294 & ~n20296;
  assign n20407 = ~n20297 & ~n20406;
  assign n20408 = n20404 & n20407;
  assign n20409 = ~n18464 & n20292;
  assign n20410 = ~n20293 & ~n20409;
  assign n20411 = n20407 & n20410;
  assign n20412 = ~n19047 & n20290;
  assign n20413 = ~n20291 & ~n20412;
  assign n20414 = n20410 & n20413;
  assign n20415 = ~n19078 & n20288;
  assign n20416 = ~n20289 & ~n20415;
  assign n20417 = n20413 & n20416;
  assign n20418 = ~n19678 & n20286;
  assign n20419 = ~n20287 & ~n20418;
  assign n20420 = n20416 & n20419;
  assign n20421 = n20282 & ~n20284;
  assign n20422 = ~n20285 & ~n20421;
  assign n20423 = n20419 & n20422;
  assign n20424 = n20278 & ~n20280;
  assign n20425 = ~n20281 & ~n20424;
  assign n20426 = n20422 & n20425;
  assign n20427 = n20274 & ~n20276;
  assign n20428 = ~n20277 & ~n20427;
  assign n20429 = n20425 & n20428;
  assign n20430 = n20270 & ~n20272;
  assign n20431 = ~n20273 & ~n20430;
  assign n20432 = n20428 & n20431;
  assign n20433 = n20266 & ~n20268;
  assign n20434 = ~n20269 & ~n20433;
  assign n20435 = n20431 & n20434;
  assign n20436 = n20262 & ~n20264;
  assign n20437 = ~n20265 & ~n20436;
  assign n20438 = n20434 & n20437;
  assign n20439 = n20258 & ~n20260;
  assign n20440 = ~n20261 & ~n20439;
  assign n20441 = n20437 & n20440;
  assign n20442 = ~n20437 & ~n20440;
  assign n20443 = ~n20441 & ~n20442;
  assign n20444 = n20254 & ~n20256;
  assign n20445 = ~n20257 & ~n20444;
  assign n20446 = ~n19797 & n20252;
  assign n20447 = ~n20253 & ~n20446;
  assign n20448 = n20445 & ~n20447;
  assign n20449 = ~n20440 & n20448;
  assign n20450 = n20445 & ~n20449;
  assign n20451 = n20443 & n20450;
  assign n20452 = ~n20441 & ~n20451;
  assign n20453 = ~n20434 & ~n20437;
  assign n20454 = ~n20438 & ~n20453;
  assign n20455 = ~n20452 & n20454;
  assign n20456 = ~n20438 & ~n20455;
  assign n20457 = ~n20431 & ~n20434;
  assign n20458 = ~n20435 & ~n20457;
  assign n20459 = ~n20456 & n20458;
  assign n20460 = ~n20435 & ~n20459;
  assign n20461 = ~n20428 & ~n20431;
  assign n20462 = ~n20432 & ~n20461;
  assign n20463 = ~n20460 & n20462;
  assign n20464 = ~n20432 & ~n20463;
  assign n20465 = ~n20425 & ~n20428;
  assign n20466 = ~n20429 & ~n20465;
  assign n20467 = ~n20464 & n20466;
  assign n20468 = ~n20429 & ~n20467;
  assign n20469 = ~n20422 & ~n20425;
  assign n20470 = ~n20426 & ~n20469;
  assign n20471 = ~n20468 & n20470;
  assign n20472 = ~n20426 & ~n20471;
  assign n20473 = ~n20419 & ~n20422;
  assign n20474 = ~n20423 & ~n20473;
  assign n20475 = ~n20472 & n20474;
  assign n20476 = ~n20423 & ~n20475;
  assign n20477 = ~n20416 & ~n20419;
  assign n20478 = ~n20420 & ~n20477;
  assign n20479 = ~n20476 & n20478;
  assign n20480 = ~n20420 & ~n20479;
  assign n20481 = ~n20413 & ~n20416;
  assign n20482 = ~n20417 & ~n20481;
  assign n20483 = ~n20480 & n20482;
  assign n20484 = ~n20417 & ~n20483;
  assign n20485 = ~n20410 & ~n20413;
  assign n20486 = ~n20414 & ~n20485;
  assign n20487 = ~n20484 & n20486;
  assign n20488 = ~n20414 & ~n20487;
  assign n20489 = ~n20407 & ~n20410;
  assign n20490 = ~n20411 & ~n20489;
  assign n20491 = ~n20488 & n20490;
  assign n20492 = ~n20411 & ~n20491;
  assign n20493 = ~n20404 & ~n20407;
  assign n20494 = ~n20408 & ~n20493;
  assign n20495 = ~n20492 & n20494;
  assign n20496 = ~n20408 & ~n20495;
  assign n20497 = ~n20401 & ~n20404;
  assign n20498 = ~n20405 & ~n20497;
  assign n20499 = ~n20496 & n20498;
  assign n20500 = ~n20405 & ~n20499;
  assign n20501 = ~n20398 & ~n20401;
  assign n20502 = ~n20402 & ~n20501;
  assign n20503 = ~n20500 & n20502;
  assign n20504 = ~n20402 & ~n20503;
  assign n20505 = ~n20395 & ~n20398;
  assign n20506 = ~n20399 & ~n20505;
  assign n20507 = ~n20504 & n20506;
  assign n20508 = ~n20399 & ~n20507;
  assign n20509 = ~n20392 & ~n20395;
  assign n20510 = ~n20396 & ~n20509;
  assign n20511 = ~n20508 & n20510;
  assign n20512 = ~n20396 & ~n20511;
  assign n20513 = ~n20389 & ~n20392;
  assign n20514 = ~n20393 & ~n20513;
  assign n20515 = ~n20512 & n20514;
  assign n20516 = ~n20393 & ~n20515;
  assign n20517 = ~n20386 & ~n20389;
  assign n20518 = ~n20390 & ~n20517;
  assign n20519 = ~n20516 & n20518;
  assign n20520 = ~n20390 & ~n20519;
  assign n20521 = ~n20383 & ~n20386;
  assign n20522 = ~n20387 & ~n20521;
  assign n20523 = ~n20520 & n20522;
  assign n20524 = ~n20387 & ~n20523;
  assign n20525 = ~n20380 & ~n20383;
  assign n20526 = ~n20384 & ~n20525;
  assign n20527 = ~n20524 & n20526;
  assign n20528 = ~n20384 & ~n20527;
  assign n20529 = ~n20377 & ~n20380;
  assign n20530 = ~n20381 & ~n20529;
  assign n20531 = ~n20528 & n20530;
  assign n20532 = ~n20381 & ~n20531;
  assign n20533 = ~n20374 & ~n20377;
  assign n20534 = ~n20378 & ~n20533;
  assign n20535 = ~n20532 & n20534;
  assign n20536 = ~n20378 & ~n20535;
  assign n20537 = ~n20371 & ~n20374;
  assign n20538 = ~n20375 & ~n20537;
  assign n20539 = ~n20536 & n20538;
  assign n20540 = ~n20375 & ~n20539;
  assign n20541 = ~n20368 & ~n20371;
  assign n20542 = ~n20372 & ~n20541;
  assign n20543 = ~n20540 & n20542;
  assign n20544 = ~n20372 & ~n20543;
  assign n20545 = ~n20365 & ~n20368;
  assign n20546 = ~n20369 & ~n20545;
  assign n20547 = ~n20544 & n20546;
  assign n20548 = ~n20369 & ~n20547;
  assign n20549 = ~n20361 & ~n20365;
  assign n20550 = ~n20366 & ~n20549;
  assign n20551 = ~n20548 & n20550;
  assign n20552 = ~n20366 & ~n20551;
  assign n20553 = ~n20358 & ~n20361;
  assign n20554 = ~n20363 & ~n20553;
  assign n20555 = ~n20552 & n20554;
  assign n20556 = ~n20363 & ~n20555;
  assign n20557 = n20355 & n20358;
  assign n20558 = ~n20355 & ~n20358;
  assign n20559 = ~n20557 & ~n20558;
  assign n20560 = ~n20556 & n20559;
  assign n20561 = n20556 & ~n20559;
  assign n20562 = ~n20560 & ~n20561;
  assign n20563 = n9830 & n20562;
  assign n20564 = ~n20359 & ~n20362;
  assign n20565 = ~n20356 & n20564;
  assign n20566 = ~n20563 & n20565;
  assign n20567 = ~pi5  & ~n20566;
  assign n20568 = pi5  & n20566;
  assign n20569 = ~n20567 & ~n20568;
  assign n20570 = n8161 & n20380;
  assign n20571 = n7847 & n20383;
  assign n20572 = n7554 & n20386;
  assign n20573 = n20524 & ~n20526;
  assign n20574 = ~n20527 & ~n20573;
  assign n20575 = n7548 & n20574;
  assign n20576 = ~n20571 & ~n20572;
  assign n20577 = ~n20570 & n20576;
  assign n20578 = ~n20575 & n20577;
  assign n20579 = ~pi11  & ~n20578;
  assign n20580 = pi11  & n20578;
  assign n20581 = ~n20579 & ~n20580;
  assign n20582 = n7380 & n20392;
  assign n20583 = n7243 & n20395;
  assign n20584 = n6653 & n20398;
  assign n20585 = n20508 & ~n20510;
  assign n20586 = ~n20511 & ~n20585;
  assign n20587 = n6647 & n20586;
  assign n20588 = ~n20583 & ~n20584;
  assign n20589 = ~n20582 & n20588;
  assign n20590 = ~n20587 & n20589;
  assign n20591 = ~pi14  & ~n20590;
  assign n20592 = pi14  & n20590;
  assign n20593 = ~n20591 & ~n20592;
  assign n20594 = n5267 & n20428;
  assign n20595 = n5185 & n20431;
  assign n20596 = n5121 & n20434;
  assign n20597 = n20460 & ~n20462;
  assign n20598 = ~n20463 & ~n20597;
  assign n20599 = n78 & n20598;
  assign n20600 = ~n20595 & ~n20596;
  assign n20601 = ~n20594 & n20600;
  assign n20602 = ~n20599 & n20601;
  assign n20603 = pi23  & n20602;
  assign n20604 = ~pi23  & ~n20602;
  assign n20605 = ~n20603 & ~n20604;
  assign n20606 = n4721 & n20437;
  assign n20607 = n4691 & n20440;
  assign n20608 = n4515 & n20445;
  assign n20609 = ~n20443 & ~n20450;
  assign n20610 = ~n20451 & ~n20609;
  assign n20611 = n4516 & n20610;
  assign n20612 = ~n20607 & ~n20608;
  assign n20613 = ~n20606 & n20612;
  assign n20614 = ~n20611 & n20613;
  assign n20615 = pi26  & n20614;
  assign n20616 = ~pi26  & ~n20614;
  assign n20617 = ~n20615 & ~n20616;
  assign n20618 = n3941 & n20447;
  assign n20619 = ~n4512 & n20447;
  assign n20620 = pi26  & n20619;
  assign n20621 = n4721 & n20445;
  assign n20622 = n4691 & n20447;
  assign n20623 = ~n20445 & n20447;
  assign n20624 = ~n20448 & ~n20623;
  assign n20625 = n4516 & ~n20624;
  assign n20626 = ~n20621 & ~n20622;
  assign n20627 = ~n20625 & n20626;
  assign n20628 = ~n20620 & n20627;
  assign n20629 = n4721 & n20440;
  assign n20630 = n4691 & n20445;
  assign n20631 = n4515 & n20447;
  assign n20632 = n20440 & ~n20448;
  assign n20633 = ~n20449 & ~n20632;
  assign n20634 = n4516 & ~n20633;
  assign n20635 = ~n20630 & ~n20631;
  assign n20636 = ~n20629 & n20635;
  assign n20637 = ~n20634 & n20636;
  assign n20638 = pi26  & n20628;
  assign n20639 = n20637 & n20638;
  assign n20640 = n20618 & n20639;
  assign n20641 = ~n20618 & ~n20639;
  assign n20642 = ~n20640 & ~n20641;
  assign n20643 = ~n20617 & n20642;
  assign n20644 = n20617 & ~n20642;
  assign n20645 = ~n20643 & ~n20644;
  assign n20646 = ~n20605 & n20645;
  assign n20647 = n5267 & n20431;
  assign n20648 = n5185 & n20434;
  assign n20649 = n5121 & n20437;
  assign n20650 = n20456 & ~n20458;
  assign n20651 = ~n20459 & ~n20650;
  assign n20652 = n78 & n20651;
  assign n20653 = ~n20648 & ~n20649;
  assign n20654 = ~n20647 & n20653;
  assign n20655 = ~n20652 & n20654;
  assign n20656 = ~pi23  & ~n20655;
  assign n20657 = pi23  & n20655;
  assign n20658 = ~n20656 & ~n20657;
  assign n20659 = pi26  & ~n20628;
  assign n20660 = n20637 & ~n20659;
  assign n20661 = ~n20637 & n20659;
  assign n20662 = ~n20660 & ~n20661;
  assign n20663 = ~n20658 & n20662;
  assign n20664 = n5267 & n20434;
  assign n20665 = n5185 & n20437;
  assign n20666 = n5121 & n20440;
  assign n20667 = n20452 & ~n20454;
  assign n20668 = ~n20455 & ~n20667;
  assign n20669 = n78 & n20668;
  assign n20670 = ~n20665 & ~n20666;
  assign n20671 = ~n20664 & n20670;
  assign n20672 = ~n20669 & n20671;
  assign n20673 = pi23  & n20672;
  assign n20674 = ~pi23  & ~n20672;
  assign n20675 = ~n20673 & ~n20674;
  assign n20676 = n20620 & ~n20627;
  assign n20677 = ~n20628 & ~n20676;
  assign n20678 = ~n20675 & n20677;
  assign n20679 = n74 & n20447;
  assign n20680 = pi23  & n20679;
  assign n20681 = n5267 & n20445;
  assign n20682 = n5185 & n20447;
  assign n20683 = n78 & ~n20624;
  assign n20684 = ~n20681 & ~n20682;
  assign n20685 = ~n20683 & n20684;
  assign n20686 = ~n20680 & n20685;
  assign n20687 = n5267 & n20440;
  assign n20688 = n5185 & n20445;
  assign n20689 = n5121 & n20447;
  assign n20690 = n78 & ~n20633;
  assign n20691 = ~n20688 & ~n20689;
  assign n20692 = ~n20687 & n20691;
  assign n20693 = ~n20690 & n20692;
  assign n20694 = pi23  & n20686;
  assign n20695 = n20693 & n20694;
  assign n20696 = n20619 & n20695;
  assign n20697 = n5267 & n20437;
  assign n20698 = n5185 & n20440;
  assign n20699 = n5121 & n20445;
  assign n20700 = n78 & n20610;
  assign n20701 = ~n20698 & ~n20699;
  assign n20702 = ~n20697 & n20701;
  assign n20703 = ~n20700 & n20702;
  assign n20704 = pi23  & n20703;
  assign n20705 = ~pi23  & ~n20703;
  assign n20706 = ~n20704 & ~n20705;
  assign n20707 = ~n20619 & ~n20695;
  assign n20708 = ~n20696 & ~n20707;
  assign n20709 = ~n20706 & n20708;
  assign n20710 = ~n20696 & ~n20709;
  assign n20711 = n20675 & ~n20677;
  assign n20712 = ~n20678 & ~n20711;
  assign n20713 = ~n20710 & n20712;
  assign n20714 = ~n20678 & ~n20713;
  assign n20715 = n20658 & ~n20662;
  assign n20716 = ~n20663 & ~n20715;
  assign n20717 = ~n20714 & n20716;
  assign n20718 = ~n20663 & ~n20717;
  assign n20719 = n20605 & ~n20645;
  assign n20720 = ~n20646 & ~n20719;
  assign n20721 = ~n20718 & n20720;
  assign n20722 = ~n20646 & ~n20721;
  assign n20723 = n5267 & n20425;
  assign n20724 = n5185 & n20428;
  assign n20725 = n5121 & n20431;
  assign n20726 = n20464 & ~n20466;
  assign n20727 = ~n20467 & ~n20726;
  assign n20728 = n78 & n20727;
  assign n20729 = ~n20724 & ~n20725;
  assign n20730 = ~n20723 & n20729;
  assign n20731 = ~n20728 & n20730;
  assign n20732 = ~pi23  & ~n20731;
  assign n20733 = pi23  & n20731;
  assign n20734 = ~n20732 & ~n20733;
  assign n20735 = ~n20640 & ~n20643;
  assign n20736 = n4721 & n20434;
  assign n20737 = n4691 & n20437;
  assign n20738 = n4515 & n20440;
  assign n20739 = n4516 & n20668;
  assign n20740 = ~n20737 & ~n20738;
  assign n20741 = ~n20736 & n20740;
  assign n20742 = ~n20739 & n20741;
  assign n20743 = pi26  & n20742;
  assign n20744 = ~pi26  & ~n20742;
  assign n20745 = ~n20743 & ~n20744;
  assign n20746 = pi29  & n20618;
  assign n20747 = n4472 & n20445;
  assign n20748 = n4070 & n20447;
  assign n20749 = n3944 & ~n20624;
  assign n20750 = ~n20747 & ~n20748;
  assign n20751 = ~n20749 & n20750;
  assign n20752 = n20746 & ~n20751;
  assign n20753 = ~n20746 & n20751;
  assign n20754 = ~n20752 & ~n20753;
  assign n20755 = ~n20745 & n20754;
  assign n20756 = n20745 & ~n20754;
  assign n20757 = ~n20755 & ~n20756;
  assign n20758 = ~n20735 & n20757;
  assign n20759 = n20735 & ~n20757;
  assign n20760 = ~n20758 & ~n20759;
  assign n20761 = ~n20734 & n20760;
  assign n20762 = n20734 & ~n20760;
  assign n20763 = ~n20761 & ~n20762;
  assign n20764 = ~n20722 & n20763;
  assign n20765 = n20722 & ~n20763;
  assign n20766 = ~n20764 & ~n20765;
  assign n20767 = n5982 & n20416;
  assign n20768 = n5901 & n20419;
  assign n20769 = n5312 & n20422;
  assign n20770 = n20476 & ~n20478;
  assign n20771 = ~n20479 & ~n20770;
  assign n20772 = n5306 & n20771;
  assign n20773 = ~n20768 & ~n20769;
  assign n20774 = ~n20767 & n20773;
  assign n20775 = ~n20772 & n20774;
  assign n20776 = pi20  & n20775;
  assign n20777 = ~pi20  & ~n20775;
  assign n20778 = ~n20776 & ~n20777;
  assign n20779 = n20766 & ~n20778;
  assign n20780 = n20718 & ~n20720;
  assign n20781 = ~n20721 & ~n20780;
  assign n20782 = n5982 & n20419;
  assign n20783 = n5901 & n20422;
  assign n20784 = n5312 & n20425;
  assign n20785 = n20472 & ~n20474;
  assign n20786 = ~n20475 & ~n20785;
  assign n20787 = n5306 & n20786;
  assign n20788 = ~n20783 & ~n20784;
  assign n20789 = ~n20782 & n20788;
  assign n20790 = ~n20787 & n20789;
  assign n20791 = pi20  & n20790;
  assign n20792 = ~pi20  & ~n20790;
  assign n20793 = ~n20791 & ~n20792;
  assign n20794 = n20781 & ~n20793;
  assign n20795 = n20714 & ~n20716;
  assign n20796 = ~n20717 & ~n20795;
  assign n20797 = n5982 & n20422;
  assign n20798 = n5901 & n20425;
  assign n20799 = n5312 & n20428;
  assign n20800 = n20468 & ~n20470;
  assign n20801 = ~n20471 & ~n20800;
  assign n20802 = n5306 & n20801;
  assign n20803 = ~n20798 & ~n20799;
  assign n20804 = ~n20797 & n20803;
  assign n20805 = ~n20802 & n20804;
  assign n20806 = pi20  & n20805;
  assign n20807 = ~pi20  & ~n20805;
  assign n20808 = ~n20806 & ~n20807;
  assign n20809 = n20796 & ~n20808;
  assign n20810 = n5982 & n20425;
  assign n20811 = n5901 & n20428;
  assign n20812 = n5312 & n20431;
  assign n20813 = n5306 & n20727;
  assign n20814 = ~n20811 & ~n20812;
  assign n20815 = ~n20810 & n20814;
  assign n20816 = ~n20813 & n20815;
  assign n20817 = ~pi20  & ~n20816;
  assign n20818 = pi20  & n20816;
  assign n20819 = ~n20817 & ~n20818;
  assign n20820 = n20710 & ~n20712;
  assign n20821 = ~n20713 & ~n20820;
  assign n20822 = ~n20819 & n20821;
  assign n20823 = n5982 & n20428;
  assign n20824 = n5901 & n20431;
  assign n20825 = n5312 & n20434;
  assign n20826 = n5306 & n20598;
  assign n20827 = ~n20824 & ~n20825;
  assign n20828 = ~n20823 & n20827;
  assign n20829 = ~n20826 & n20828;
  assign n20830 = pi20  & n20829;
  assign n20831 = ~pi20  & ~n20829;
  assign n20832 = ~n20830 & ~n20831;
  assign n20833 = n20706 & ~n20708;
  assign n20834 = ~n20709 & ~n20833;
  assign n20835 = ~n20832 & n20834;
  assign n20836 = n5982 & n20431;
  assign n20837 = n5901 & n20434;
  assign n20838 = n5312 & n20437;
  assign n20839 = n5306 & n20651;
  assign n20840 = ~n20837 & ~n20838;
  assign n20841 = ~n20836 & n20840;
  assign n20842 = ~n20839 & n20841;
  assign n20843 = ~pi20  & ~n20842;
  assign n20844 = pi20  & n20842;
  assign n20845 = ~n20843 & ~n20844;
  assign n20846 = pi23  & ~n20686;
  assign n20847 = n20693 & ~n20846;
  assign n20848 = ~n20693 & n20846;
  assign n20849 = ~n20847 & ~n20848;
  assign n20850 = ~n20845 & n20849;
  assign n20851 = n5982 & n20434;
  assign n20852 = n5901 & n20437;
  assign n20853 = n5312 & n20440;
  assign n20854 = n5306 & n20668;
  assign n20855 = ~n20852 & ~n20853;
  assign n20856 = ~n20851 & n20855;
  assign n20857 = ~n20854 & n20856;
  assign n20858 = pi20  & n20857;
  assign n20859 = ~pi20  & ~n20857;
  assign n20860 = ~n20858 & ~n20859;
  assign n20861 = n20680 & ~n20685;
  assign n20862 = ~n20686 & ~n20861;
  assign n20863 = ~n20860 & n20862;
  assign n20864 = n5305 & n20447;
  assign n20865 = pi20  & n20864;
  assign n20866 = n5982 & n20445;
  assign n20867 = n5901 & n20447;
  assign n20868 = n5306 & ~n20624;
  assign n20869 = ~n20866 & ~n20867;
  assign n20870 = ~n20868 & n20869;
  assign n20871 = ~n20865 & n20870;
  assign n20872 = n5982 & n20440;
  assign n20873 = n5901 & n20445;
  assign n20874 = n5312 & n20447;
  assign n20875 = n5306 & ~n20633;
  assign n20876 = ~n20873 & ~n20874;
  assign n20877 = ~n20872 & n20876;
  assign n20878 = ~n20875 & n20877;
  assign n20879 = pi20  & n20871;
  assign n20880 = n20878 & n20879;
  assign n20881 = n20679 & n20880;
  assign n20882 = n5982 & n20437;
  assign n20883 = n5901 & n20440;
  assign n20884 = n5312 & n20445;
  assign n20885 = n5306 & n20610;
  assign n20886 = ~n20883 & ~n20884;
  assign n20887 = ~n20882 & n20886;
  assign n20888 = ~n20885 & n20887;
  assign n20889 = pi20  & n20888;
  assign n20890 = ~pi20  & ~n20888;
  assign n20891 = ~n20889 & ~n20890;
  assign n20892 = ~n20679 & ~n20880;
  assign n20893 = ~n20881 & ~n20892;
  assign n20894 = ~n20891 & n20893;
  assign n20895 = ~n20881 & ~n20894;
  assign n20896 = n20860 & ~n20862;
  assign n20897 = ~n20863 & ~n20896;
  assign n20898 = ~n20895 & n20897;
  assign n20899 = ~n20863 & ~n20898;
  assign n20900 = n20845 & ~n20849;
  assign n20901 = ~n20850 & ~n20900;
  assign n20902 = ~n20899 & n20901;
  assign n20903 = ~n20850 & ~n20902;
  assign n20904 = n20832 & ~n20834;
  assign n20905 = ~n20835 & ~n20904;
  assign n20906 = ~n20903 & n20905;
  assign n20907 = ~n20835 & ~n20906;
  assign n20908 = n20819 & ~n20821;
  assign n20909 = ~n20822 & ~n20908;
  assign n20910 = ~n20907 & n20909;
  assign n20911 = ~n20822 & ~n20910;
  assign n20912 = ~n20796 & n20808;
  assign n20913 = ~n20809 & ~n20912;
  assign n20914 = ~n20911 & n20913;
  assign n20915 = ~n20809 & ~n20914;
  assign n20916 = ~n20781 & n20793;
  assign n20917 = ~n20794 & ~n20916;
  assign n20918 = ~n20915 & n20917;
  assign n20919 = ~n20794 & ~n20918;
  assign n20920 = ~n20766 & n20778;
  assign n20921 = ~n20779 & ~n20920;
  assign n20922 = ~n20919 & n20921;
  assign n20923 = ~n20779 & ~n20922;
  assign n20924 = n5982 & n20413;
  assign n20925 = n5901 & n20416;
  assign n20926 = n5312 & n20419;
  assign n20927 = n20480 & ~n20482;
  assign n20928 = ~n20483 & ~n20927;
  assign n20929 = n5306 & n20928;
  assign n20930 = ~n20925 & ~n20926;
  assign n20931 = ~n20924 & n20930;
  assign n20932 = ~n20929 & n20931;
  assign n20933 = ~pi20  & ~n20932;
  assign n20934 = pi20  & n20932;
  assign n20935 = ~n20933 & ~n20934;
  assign n20936 = ~n20761 & ~n20764;
  assign n20937 = ~n20755 & ~n20758;
  assign n20938 = n4721 & n20431;
  assign n20939 = n4691 & n20434;
  assign n20940 = n4515 & n20437;
  assign n20941 = n4516 & n20651;
  assign n20942 = ~n20939 & ~n20940;
  assign n20943 = ~n20938 & n20942;
  assign n20944 = ~n20941 & n20943;
  assign n20945 = ~pi26  & ~n20944;
  assign n20946 = pi26  & n20944;
  assign n20947 = ~n20945 & ~n20946;
  assign n20948 = pi29  & ~n20753;
  assign n20949 = n4472 & n20440;
  assign n20950 = n4070 & n20445;
  assign n20951 = n3943 & n20447;
  assign n20952 = n3944 & ~n20633;
  assign n20953 = ~n20950 & ~n20951;
  assign n20954 = ~n20949 & n20953;
  assign n20955 = ~n20952 & n20954;
  assign n20956 = ~n20948 & n20955;
  assign n20957 = n20948 & ~n20955;
  assign n20958 = ~n20956 & ~n20957;
  assign n20959 = ~n20947 & n20958;
  assign n20960 = n20947 & ~n20958;
  assign n20961 = ~n20959 & ~n20960;
  assign n20962 = ~n20937 & n20961;
  assign n20963 = n20937 & ~n20961;
  assign n20964 = ~n20962 & ~n20963;
  assign n20965 = n5267 & n20422;
  assign n20966 = n5185 & n20425;
  assign n20967 = n5121 & n20428;
  assign n20968 = n78 & n20801;
  assign n20969 = ~n20966 & ~n20967;
  assign n20970 = ~n20965 & n20969;
  assign n20971 = ~n20968 & n20970;
  assign n20972 = pi23  & n20971;
  assign n20973 = ~pi23  & ~n20971;
  assign n20974 = ~n20972 & ~n20973;
  assign n20975 = n20964 & ~n20974;
  assign n20976 = ~n20964 & n20974;
  assign n20977 = ~n20975 & ~n20976;
  assign n20978 = ~n20936 & n20977;
  assign n20979 = n20936 & ~n20977;
  assign n20980 = ~n20978 & ~n20979;
  assign n20981 = ~n20935 & n20980;
  assign n20982 = n20935 & ~n20980;
  assign n20983 = ~n20981 & ~n20982;
  assign n20984 = ~n20923 & n20983;
  assign n20985 = n20923 & ~n20983;
  assign n20986 = ~n20984 & ~n20985;
  assign n20987 = n6608 & n20404;
  assign n20988 = n6356 & n20407;
  assign n20989 = n6140 & n20410;
  assign n20990 = n20492 & ~n20494;
  assign n20991 = ~n20495 & ~n20990;
  assign n20992 = n6134 & n20991;
  assign n20993 = ~n20988 & ~n20989;
  assign n20994 = ~n20987 & n20993;
  assign n20995 = ~n20992 & n20994;
  assign n20996 = pi17  & n20995;
  assign n20997 = ~pi17  & ~n20995;
  assign n20998 = ~n20996 & ~n20997;
  assign n20999 = n20986 & ~n20998;
  assign n21000 = n6608 & n20407;
  assign n21001 = n6356 & n20410;
  assign n21002 = n6140 & n20413;
  assign n21003 = n20488 & ~n20490;
  assign n21004 = ~n20491 & ~n21003;
  assign n21005 = n6134 & n21004;
  assign n21006 = ~n21001 & ~n21002;
  assign n21007 = ~n21000 & n21006;
  assign n21008 = ~n21005 & n21007;
  assign n21009 = ~pi17  & ~n21008;
  assign n21010 = pi17  & n21008;
  assign n21011 = ~n21009 & ~n21010;
  assign n21012 = n20919 & ~n20921;
  assign n21013 = ~n20922 & ~n21012;
  assign n21014 = ~n21011 & n21013;
  assign n21015 = n6608 & n20410;
  assign n21016 = n6356 & n20413;
  assign n21017 = n6140 & n20416;
  assign n21018 = n20484 & ~n20486;
  assign n21019 = ~n20487 & ~n21018;
  assign n21020 = n6134 & n21019;
  assign n21021 = ~n21016 & ~n21017;
  assign n21022 = ~n21015 & n21021;
  assign n21023 = ~n21020 & n21022;
  assign n21024 = ~pi17  & ~n21023;
  assign n21025 = pi17  & n21023;
  assign n21026 = ~n21024 & ~n21025;
  assign n21027 = n20915 & ~n20917;
  assign n21028 = ~n20918 & ~n21027;
  assign n21029 = ~n21026 & n21028;
  assign n21030 = n6608 & n20413;
  assign n21031 = n6356 & n20416;
  assign n21032 = n6140 & n20419;
  assign n21033 = n6134 & n20928;
  assign n21034 = ~n21031 & ~n21032;
  assign n21035 = ~n21030 & n21034;
  assign n21036 = ~n21033 & n21035;
  assign n21037 = ~pi17  & ~n21036;
  assign n21038 = pi17  & n21036;
  assign n21039 = ~n21037 & ~n21038;
  assign n21040 = n20911 & ~n20913;
  assign n21041 = ~n20914 & ~n21040;
  assign n21042 = ~n21039 & n21041;
  assign n21043 = n20907 & ~n20909;
  assign n21044 = ~n20910 & ~n21043;
  assign n21045 = n6608 & n20416;
  assign n21046 = n6356 & n20419;
  assign n21047 = n6140 & n20422;
  assign n21048 = n6134 & n20771;
  assign n21049 = ~n21046 & ~n21047;
  assign n21050 = ~n21045 & n21049;
  assign n21051 = ~n21048 & n21050;
  assign n21052 = pi17  & n21051;
  assign n21053 = ~pi17  & ~n21051;
  assign n21054 = ~n21052 & ~n21053;
  assign n21055 = n21044 & ~n21054;
  assign n21056 = n20903 & ~n20905;
  assign n21057 = ~n20906 & ~n21056;
  assign n21058 = n6608 & n20419;
  assign n21059 = n6356 & n20422;
  assign n21060 = n6140 & n20425;
  assign n21061 = n6134 & n20786;
  assign n21062 = ~n21059 & ~n21060;
  assign n21063 = ~n21058 & n21062;
  assign n21064 = ~n21061 & n21063;
  assign n21065 = pi17  & n21064;
  assign n21066 = ~pi17  & ~n21064;
  assign n21067 = ~n21065 & ~n21066;
  assign n21068 = n21057 & ~n21067;
  assign n21069 = n20899 & ~n20901;
  assign n21070 = ~n20902 & ~n21069;
  assign n21071 = n6608 & n20422;
  assign n21072 = n6356 & n20425;
  assign n21073 = n6140 & n20428;
  assign n21074 = n6134 & n20801;
  assign n21075 = ~n21072 & ~n21073;
  assign n21076 = ~n21071 & n21075;
  assign n21077 = ~n21074 & n21076;
  assign n21078 = pi17  & n21077;
  assign n21079 = ~pi17  & ~n21077;
  assign n21080 = ~n21078 & ~n21079;
  assign n21081 = n21070 & ~n21080;
  assign n21082 = n6608 & n20425;
  assign n21083 = n6356 & n20428;
  assign n21084 = n6140 & n20431;
  assign n21085 = n6134 & n20727;
  assign n21086 = ~n21083 & ~n21084;
  assign n21087 = ~n21082 & n21086;
  assign n21088 = ~n21085 & n21087;
  assign n21089 = ~pi17  & ~n21088;
  assign n21090 = pi17  & n21088;
  assign n21091 = ~n21089 & ~n21090;
  assign n21092 = n20895 & ~n20897;
  assign n21093 = ~n20898 & ~n21092;
  assign n21094 = ~n21091 & n21093;
  assign n21095 = n6608 & n20428;
  assign n21096 = n6356 & n20431;
  assign n21097 = n6140 & n20434;
  assign n21098 = n6134 & n20598;
  assign n21099 = ~n21096 & ~n21097;
  assign n21100 = ~n21095 & n21099;
  assign n21101 = ~n21098 & n21100;
  assign n21102 = pi17  & n21101;
  assign n21103 = ~pi17  & ~n21101;
  assign n21104 = ~n21102 & ~n21103;
  assign n21105 = n20891 & ~n20893;
  assign n21106 = ~n20894 & ~n21105;
  assign n21107 = ~n21104 & n21106;
  assign n21108 = n6608 & n20431;
  assign n21109 = n6356 & n20434;
  assign n21110 = n6140 & n20437;
  assign n21111 = n6134 & n20651;
  assign n21112 = ~n21109 & ~n21110;
  assign n21113 = ~n21108 & n21112;
  assign n21114 = ~n21111 & n21113;
  assign n21115 = ~pi17  & ~n21114;
  assign n21116 = pi17  & n21114;
  assign n21117 = ~n21115 & ~n21116;
  assign n21118 = pi20  & ~n20871;
  assign n21119 = n20878 & ~n21118;
  assign n21120 = ~n20878 & n21118;
  assign n21121 = ~n21119 & ~n21120;
  assign n21122 = ~n21117 & n21121;
  assign n21123 = n6608 & n20434;
  assign n21124 = n6356 & n20437;
  assign n21125 = n6140 & n20440;
  assign n21126 = n6134 & n20668;
  assign n21127 = ~n21124 & ~n21125;
  assign n21128 = ~n21123 & n21127;
  assign n21129 = ~n21126 & n21128;
  assign n21130 = pi17  & n21129;
  assign n21131 = ~pi17  & ~n21129;
  assign n21132 = ~n21130 & ~n21131;
  assign n21133 = n20865 & ~n20870;
  assign n21134 = ~n20871 & ~n21133;
  assign n21135 = ~n21132 & n21134;
  assign n21136 = n6130 & n20447;
  assign n21137 = pi17  & n21136;
  assign n21138 = n6608 & n20445;
  assign n21139 = n6356 & n20447;
  assign n21140 = n6134 & ~n20624;
  assign n21141 = ~n21138 & ~n21139;
  assign n21142 = ~n21140 & n21141;
  assign n21143 = ~n21137 & n21142;
  assign n21144 = n6608 & n20440;
  assign n21145 = n6356 & n20445;
  assign n21146 = n6140 & n20447;
  assign n21147 = n6134 & ~n20633;
  assign n21148 = ~n21145 & ~n21146;
  assign n21149 = ~n21144 & n21148;
  assign n21150 = ~n21147 & n21149;
  assign n21151 = pi17  & n21143;
  assign n21152 = n21150 & n21151;
  assign n21153 = n20864 & n21152;
  assign n21154 = n6608 & n20437;
  assign n21155 = n6356 & n20440;
  assign n21156 = n6140 & n20445;
  assign n21157 = n6134 & n20610;
  assign n21158 = ~n21155 & ~n21156;
  assign n21159 = ~n21154 & n21158;
  assign n21160 = ~n21157 & n21159;
  assign n21161 = pi17  & n21160;
  assign n21162 = ~pi17  & ~n21160;
  assign n21163 = ~n21161 & ~n21162;
  assign n21164 = ~n20864 & ~n21152;
  assign n21165 = ~n21153 & ~n21164;
  assign n21166 = ~n21163 & n21165;
  assign n21167 = ~n21153 & ~n21166;
  assign n21168 = n21132 & ~n21134;
  assign n21169 = ~n21135 & ~n21168;
  assign n21170 = ~n21167 & n21169;
  assign n21171 = ~n21135 & ~n21170;
  assign n21172 = n21117 & ~n21121;
  assign n21173 = ~n21122 & ~n21172;
  assign n21174 = ~n21171 & n21173;
  assign n21175 = ~n21122 & ~n21174;
  assign n21176 = n21104 & ~n21106;
  assign n21177 = ~n21107 & ~n21176;
  assign n21178 = ~n21175 & n21177;
  assign n21179 = ~n21107 & ~n21178;
  assign n21180 = n21091 & ~n21093;
  assign n21181 = ~n21094 & ~n21180;
  assign n21182 = ~n21179 & n21181;
  assign n21183 = ~n21094 & ~n21182;
  assign n21184 = ~n21070 & n21080;
  assign n21185 = ~n21081 & ~n21184;
  assign n21186 = ~n21183 & n21185;
  assign n21187 = ~n21081 & ~n21186;
  assign n21188 = ~n21057 & n21067;
  assign n21189 = ~n21068 & ~n21188;
  assign n21190 = ~n21187 & n21189;
  assign n21191 = ~n21068 & ~n21190;
  assign n21192 = ~n21044 & n21054;
  assign n21193 = ~n21055 & ~n21192;
  assign n21194 = ~n21191 & n21193;
  assign n21195 = ~n21055 & ~n21194;
  assign n21196 = n21039 & ~n21041;
  assign n21197 = ~n21042 & ~n21196;
  assign n21198 = ~n21195 & n21197;
  assign n21199 = ~n21042 & ~n21198;
  assign n21200 = n21026 & ~n21028;
  assign n21201 = ~n21029 & ~n21200;
  assign n21202 = ~n21199 & n21201;
  assign n21203 = ~n21029 & ~n21202;
  assign n21204 = n21011 & ~n21013;
  assign n21205 = ~n21014 & ~n21204;
  assign n21206 = ~n21203 & n21205;
  assign n21207 = ~n21014 & ~n21206;
  assign n21208 = ~n20986 & n20998;
  assign n21209 = ~n20999 & ~n21208;
  assign n21210 = ~n21207 & n21209;
  assign n21211 = ~n20999 & ~n21210;
  assign n21212 = ~n20981 & ~n20984;
  assign n21213 = n5982 & n20410;
  assign n21214 = n5901 & n20413;
  assign n21215 = n5312 & n20416;
  assign n21216 = n5306 & n21019;
  assign n21217 = ~n21214 & ~n21215;
  assign n21218 = ~n21213 & n21217;
  assign n21219 = ~n21216 & n21218;
  assign n21220 = ~pi20  & ~n21219;
  assign n21221 = pi20  & n21219;
  assign n21222 = ~n21220 & ~n21221;
  assign n21223 = ~n20975 & ~n20978;
  assign n21224 = ~n20959 & ~n20962;
  assign n21225 = n4721 & n20428;
  assign n21226 = n4691 & n20431;
  assign n21227 = n4515 & n20434;
  assign n21228 = n4516 & n20598;
  assign n21229 = ~n21226 & ~n21227;
  assign n21230 = ~n21225 & n21229;
  assign n21231 = ~n21228 & n21230;
  assign n21232 = ~pi26  & ~n21231;
  assign n21233 = pi26  & n21231;
  assign n21234 = ~n21232 & ~n21233;
  assign n21235 = n4472 & n20437;
  assign n21236 = n4070 & n20440;
  assign n21237 = n3943 & n20445;
  assign n21238 = n3944 & n20610;
  assign n21239 = ~n21236 & ~n21237;
  assign n21240 = ~n21235 & n21239;
  assign n21241 = ~n21238 & n21240;
  assign n21242 = ~pi29  & ~n21241;
  assign n21243 = pi29  & n21241;
  assign n21244 = ~n21242 & ~n21243;
  assign n21245 = ~n565 & n20447;
  assign n21246 = pi29  & n20753;
  assign n21247 = n20955 & n21246;
  assign n21248 = n21245 & n21247;
  assign n21249 = ~n21245 & ~n21247;
  assign n21250 = ~n21248 & ~n21249;
  assign n21251 = ~n21244 & n21250;
  assign n21252 = n21244 & ~n21250;
  assign n21253 = ~n21251 & ~n21252;
  assign n21254 = ~n21234 & n21253;
  assign n21255 = n21234 & ~n21253;
  assign n21256 = ~n21254 & ~n21255;
  assign n21257 = ~n21224 & n21256;
  assign n21258 = n21224 & ~n21256;
  assign n21259 = ~n21257 & ~n21258;
  assign n21260 = n5267 & n20419;
  assign n21261 = n5185 & n20422;
  assign n21262 = n5121 & n20425;
  assign n21263 = n78 & n20786;
  assign n21264 = ~n21261 & ~n21262;
  assign n21265 = ~n21260 & n21264;
  assign n21266 = ~n21263 & n21265;
  assign n21267 = pi23  & n21266;
  assign n21268 = ~pi23  & ~n21266;
  assign n21269 = ~n21267 & ~n21268;
  assign n21270 = n21259 & ~n21269;
  assign n21271 = ~n21259 & n21269;
  assign n21272 = ~n21270 & ~n21271;
  assign n21273 = ~n21223 & n21272;
  assign n21274 = n21223 & ~n21272;
  assign n21275 = ~n21273 & ~n21274;
  assign n21276 = ~n21222 & n21275;
  assign n21277 = n21222 & ~n21275;
  assign n21278 = ~n21276 & ~n21277;
  assign n21279 = ~n21212 & n21278;
  assign n21280 = n21212 & ~n21278;
  assign n21281 = ~n21279 & ~n21280;
  assign n21282 = n6608 & n20401;
  assign n21283 = n6356 & n20404;
  assign n21284 = n6140 & n20407;
  assign n21285 = n20496 & ~n20498;
  assign n21286 = ~n20499 & ~n21285;
  assign n21287 = n6134 & n21286;
  assign n21288 = ~n21283 & ~n21284;
  assign n21289 = ~n21282 & n21288;
  assign n21290 = ~n21287 & n21289;
  assign n21291 = pi17  & n21290;
  assign n21292 = ~pi17  & ~n21290;
  assign n21293 = ~n21291 & ~n21292;
  assign n21294 = n21281 & ~n21293;
  assign n21295 = ~n21281 & n21293;
  assign n21296 = ~n21294 & ~n21295;
  assign n21297 = ~n21211 & n21296;
  assign n21298 = n21211 & ~n21296;
  assign n21299 = ~n21297 & ~n21298;
  assign n21300 = ~n20593 & n21299;
  assign n21301 = n7380 & n20395;
  assign n21302 = n7243 & n20398;
  assign n21303 = n6653 & n20401;
  assign n21304 = n20504 & ~n20506;
  assign n21305 = ~n20507 & ~n21304;
  assign n21306 = n6647 & n21305;
  assign n21307 = ~n21302 & ~n21303;
  assign n21308 = ~n21301 & n21307;
  assign n21309 = ~n21306 & n21308;
  assign n21310 = ~pi14  & ~n21309;
  assign n21311 = pi14  & n21309;
  assign n21312 = ~n21310 & ~n21311;
  assign n21313 = n21207 & ~n21209;
  assign n21314 = ~n21210 & ~n21313;
  assign n21315 = ~n21312 & n21314;
  assign n21316 = n21203 & ~n21205;
  assign n21317 = ~n21206 & ~n21316;
  assign n21318 = n7380 & n20398;
  assign n21319 = n7243 & n20401;
  assign n21320 = n6653 & n20404;
  assign n21321 = n20500 & ~n20502;
  assign n21322 = ~n20503 & ~n21321;
  assign n21323 = n6647 & n21322;
  assign n21324 = ~n21319 & ~n21320;
  assign n21325 = ~n21318 & n21324;
  assign n21326 = ~n21323 & n21325;
  assign n21327 = pi14  & n21326;
  assign n21328 = ~pi14  & ~n21326;
  assign n21329 = ~n21327 & ~n21328;
  assign n21330 = n21317 & ~n21329;
  assign n21331 = n21199 & ~n21201;
  assign n21332 = ~n21202 & ~n21331;
  assign n21333 = n7380 & n20401;
  assign n21334 = n7243 & n20404;
  assign n21335 = n6653 & n20407;
  assign n21336 = n6647 & n21286;
  assign n21337 = ~n21334 & ~n21335;
  assign n21338 = ~n21333 & n21337;
  assign n21339 = ~n21336 & n21338;
  assign n21340 = pi14  & n21339;
  assign n21341 = ~pi14  & ~n21339;
  assign n21342 = ~n21340 & ~n21341;
  assign n21343 = n21332 & ~n21342;
  assign n21344 = n21195 & ~n21197;
  assign n21345 = ~n21198 & ~n21344;
  assign n21346 = n7380 & n20404;
  assign n21347 = n7243 & n20407;
  assign n21348 = n6653 & n20410;
  assign n21349 = n6647 & n20991;
  assign n21350 = ~n21347 & ~n21348;
  assign n21351 = ~n21346 & n21350;
  assign n21352 = ~n21349 & n21351;
  assign n21353 = pi14  & n21352;
  assign n21354 = ~pi14  & ~n21352;
  assign n21355 = ~n21353 & ~n21354;
  assign n21356 = n21345 & ~n21355;
  assign n21357 = n7380 & n20407;
  assign n21358 = n7243 & n20410;
  assign n21359 = n6653 & n20413;
  assign n21360 = n6647 & n21004;
  assign n21361 = ~n21358 & ~n21359;
  assign n21362 = ~n21357 & n21361;
  assign n21363 = ~n21360 & n21362;
  assign n21364 = ~pi14  & ~n21363;
  assign n21365 = pi14  & n21363;
  assign n21366 = ~n21364 & ~n21365;
  assign n21367 = n21191 & ~n21193;
  assign n21368 = ~n21194 & ~n21367;
  assign n21369 = ~n21366 & n21368;
  assign n21370 = n7380 & n20410;
  assign n21371 = n7243 & n20413;
  assign n21372 = n6653 & n20416;
  assign n21373 = n6647 & n21019;
  assign n21374 = ~n21371 & ~n21372;
  assign n21375 = ~n21370 & n21374;
  assign n21376 = ~n21373 & n21375;
  assign n21377 = ~pi14  & ~n21376;
  assign n21378 = pi14  & n21376;
  assign n21379 = ~n21377 & ~n21378;
  assign n21380 = n21187 & ~n21189;
  assign n21381 = ~n21190 & ~n21380;
  assign n21382 = ~n21379 & n21381;
  assign n21383 = n7380 & n20413;
  assign n21384 = n7243 & n20416;
  assign n21385 = n6653 & n20419;
  assign n21386 = n6647 & n20928;
  assign n21387 = ~n21384 & ~n21385;
  assign n21388 = ~n21383 & n21387;
  assign n21389 = ~n21386 & n21388;
  assign n21390 = ~pi14  & ~n21389;
  assign n21391 = pi14  & n21389;
  assign n21392 = ~n21390 & ~n21391;
  assign n21393 = n21183 & ~n21185;
  assign n21394 = ~n21186 & ~n21393;
  assign n21395 = ~n21392 & n21394;
  assign n21396 = n21179 & ~n21181;
  assign n21397 = ~n21182 & ~n21396;
  assign n21398 = n7380 & n20416;
  assign n21399 = n7243 & n20419;
  assign n21400 = n6653 & n20422;
  assign n21401 = n6647 & n20771;
  assign n21402 = ~n21399 & ~n21400;
  assign n21403 = ~n21398 & n21402;
  assign n21404 = ~n21401 & n21403;
  assign n21405 = pi14  & n21404;
  assign n21406 = ~pi14  & ~n21404;
  assign n21407 = ~n21405 & ~n21406;
  assign n21408 = n21397 & ~n21407;
  assign n21409 = n21175 & ~n21177;
  assign n21410 = ~n21178 & ~n21409;
  assign n21411 = n7380 & n20419;
  assign n21412 = n7243 & n20422;
  assign n21413 = n6653 & n20425;
  assign n21414 = n6647 & n20786;
  assign n21415 = ~n21412 & ~n21413;
  assign n21416 = ~n21411 & n21415;
  assign n21417 = ~n21414 & n21416;
  assign n21418 = pi14  & n21417;
  assign n21419 = ~pi14  & ~n21417;
  assign n21420 = ~n21418 & ~n21419;
  assign n21421 = n21410 & ~n21420;
  assign n21422 = n21171 & ~n21173;
  assign n21423 = ~n21174 & ~n21422;
  assign n21424 = n7380 & n20422;
  assign n21425 = n7243 & n20425;
  assign n21426 = n6653 & n20428;
  assign n21427 = n6647 & n20801;
  assign n21428 = ~n21425 & ~n21426;
  assign n21429 = ~n21424 & n21428;
  assign n21430 = ~n21427 & n21429;
  assign n21431 = pi14  & n21430;
  assign n21432 = ~pi14  & ~n21430;
  assign n21433 = ~n21431 & ~n21432;
  assign n21434 = n21423 & ~n21433;
  assign n21435 = n7380 & n20425;
  assign n21436 = n7243 & n20428;
  assign n21437 = n6653 & n20431;
  assign n21438 = n6647 & n20727;
  assign n21439 = ~n21436 & ~n21437;
  assign n21440 = ~n21435 & n21439;
  assign n21441 = ~n21438 & n21440;
  assign n21442 = ~pi14  & ~n21441;
  assign n21443 = pi14  & n21441;
  assign n21444 = ~n21442 & ~n21443;
  assign n21445 = n21167 & ~n21169;
  assign n21446 = ~n21170 & ~n21445;
  assign n21447 = ~n21444 & n21446;
  assign n21448 = n7380 & n20428;
  assign n21449 = n7243 & n20431;
  assign n21450 = n6653 & n20434;
  assign n21451 = n6647 & n20598;
  assign n21452 = ~n21449 & ~n21450;
  assign n21453 = ~n21448 & n21452;
  assign n21454 = ~n21451 & n21453;
  assign n21455 = pi14  & n21454;
  assign n21456 = ~pi14  & ~n21454;
  assign n21457 = ~n21455 & ~n21456;
  assign n21458 = n21163 & ~n21165;
  assign n21459 = ~n21166 & ~n21458;
  assign n21460 = ~n21457 & n21459;
  assign n21461 = n7380 & n20431;
  assign n21462 = n7243 & n20434;
  assign n21463 = n6653 & n20437;
  assign n21464 = n6647 & n20651;
  assign n21465 = ~n21462 & ~n21463;
  assign n21466 = ~n21461 & n21465;
  assign n21467 = ~n21464 & n21466;
  assign n21468 = ~pi14  & ~n21467;
  assign n21469 = pi14  & n21467;
  assign n21470 = ~n21468 & ~n21469;
  assign n21471 = pi17  & ~n21143;
  assign n21472 = n21150 & ~n21471;
  assign n21473 = ~n21150 & n21471;
  assign n21474 = ~n21472 & ~n21473;
  assign n21475 = ~n21470 & n21474;
  assign n21476 = n7380 & n20434;
  assign n21477 = n7243 & n20437;
  assign n21478 = n6653 & n20440;
  assign n21479 = n6647 & n20668;
  assign n21480 = ~n21477 & ~n21478;
  assign n21481 = ~n21476 & n21480;
  assign n21482 = ~n21479 & n21481;
  assign n21483 = pi14  & n21482;
  assign n21484 = ~pi14  & ~n21482;
  assign n21485 = ~n21483 & ~n21484;
  assign n21486 = n21137 & ~n21142;
  assign n21487 = ~n21143 & ~n21486;
  assign n21488 = ~n21485 & n21487;
  assign n21489 = n6643 & n20447;
  assign n21490 = pi14  & n21489;
  assign n21491 = n7380 & n20445;
  assign n21492 = n7243 & n20447;
  assign n21493 = n6647 & ~n20624;
  assign n21494 = ~n21491 & ~n21492;
  assign n21495 = ~n21493 & n21494;
  assign n21496 = ~n21490 & n21495;
  assign n21497 = n7380 & n20440;
  assign n21498 = n7243 & n20445;
  assign n21499 = n6653 & n20447;
  assign n21500 = n6647 & ~n20633;
  assign n21501 = ~n21498 & ~n21499;
  assign n21502 = ~n21497 & n21501;
  assign n21503 = ~n21500 & n21502;
  assign n21504 = pi14  & n21496;
  assign n21505 = n21503 & n21504;
  assign n21506 = n21136 & n21505;
  assign n21507 = n7380 & n20437;
  assign n21508 = n7243 & n20440;
  assign n21509 = n6653 & n20445;
  assign n21510 = n6647 & n20610;
  assign n21511 = ~n21508 & ~n21509;
  assign n21512 = ~n21507 & n21511;
  assign n21513 = ~n21510 & n21512;
  assign n21514 = pi14  & n21513;
  assign n21515 = ~pi14  & ~n21513;
  assign n21516 = ~n21514 & ~n21515;
  assign n21517 = ~n21136 & ~n21505;
  assign n21518 = ~n21506 & ~n21517;
  assign n21519 = ~n21516 & n21518;
  assign n21520 = ~n21506 & ~n21519;
  assign n21521 = n21485 & ~n21487;
  assign n21522 = ~n21488 & ~n21521;
  assign n21523 = ~n21520 & n21522;
  assign n21524 = ~n21488 & ~n21523;
  assign n21525 = n21470 & ~n21474;
  assign n21526 = ~n21475 & ~n21525;
  assign n21527 = ~n21524 & n21526;
  assign n21528 = ~n21475 & ~n21527;
  assign n21529 = n21457 & ~n21459;
  assign n21530 = ~n21460 & ~n21529;
  assign n21531 = ~n21528 & n21530;
  assign n21532 = ~n21460 & ~n21531;
  assign n21533 = n21444 & ~n21446;
  assign n21534 = ~n21447 & ~n21533;
  assign n21535 = ~n21532 & n21534;
  assign n21536 = ~n21447 & ~n21535;
  assign n21537 = ~n21423 & n21433;
  assign n21538 = ~n21434 & ~n21537;
  assign n21539 = ~n21536 & n21538;
  assign n21540 = ~n21434 & ~n21539;
  assign n21541 = ~n21410 & n21420;
  assign n21542 = ~n21421 & ~n21541;
  assign n21543 = ~n21540 & n21542;
  assign n21544 = ~n21421 & ~n21543;
  assign n21545 = ~n21397 & n21407;
  assign n21546 = ~n21408 & ~n21545;
  assign n21547 = ~n21544 & n21546;
  assign n21548 = ~n21408 & ~n21547;
  assign n21549 = n21392 & ~n21394;
  assign n21550 = ~n21395 & ~n21549;
  assign n21551 = ~n21548 & n21550;
  assign n21552 = ~n21395 & ~n21551;
  assign n21553 = n21379 & ~n21381;
  assign n21554 = ~n21382 & ~n21553;
  assign n21555 = ~n21552 & n21554;
  assign n21556 = ~n21382 & ~n21555;
  assign n21557 = n21366 & ~n21368;
  assign n21558 = ~n21369 & ~n21557;
  assign n21559 = ~n21556 & n21558;
  assign n21560 = ~n21369 & ~n21559;
  assign n21561 = ~n21345 & n21355;
  assign n21562 = ~n21356 & ~n21561;
  assign n21563 = ~n21560 & n21562;
  assign n21564 = ~n21356 & ~n21563;
  assign n21565 = ~n21332 & n21342;
  assign n21566 = ~n21343 & ~n21565;
  assign n21567 = ~n21564 & n21566;
  assign n21568 = ~n21343 & ~n21567;
  assign n21569 = ~n21317 & n21329;
  assign n21570 = ~n21330 & ~n21569;
  assign n21571 = ~n21568 & n21570;
  assign n21572 = ~n21330 & ~n21571;
  assign n21573 = n21312 & ~n21314;
  assign n21574 = ~n21315 & ~n21573;
  assign n21575 = ~n21572 & n21574;
  assign n21576 = ~n21315 & ~n21575;
  assign n21577 = n20593 & ~n21299;
  assign n21578 = ~n21300 & ~n21577;
  assign n21579 = ~n21576 & n21578;
  assign n21580 = ~n21300 & ~n21579;
  assign n21581 = ~n21294 & ~n21297;
  assign n21582 = n6608 & n20398;
  assign n21583 = n6356 & n20401;
  assign n21584 = n6140 & n20404;
  assign n21585 = n6134 & n21322;
  assign n21586 = ~n21583 & ~n21584;
  assign n21587 = ~n21582 & n21586;
  assign n21588 = ~n21585 & n21587;
  assign n21589 = ~pi17  & ~n21588;
  assign n21590 = pi17  & n21588;
  assign n21591 = ~n21589 & ~n21590;
  assign n21592 = ~n21276 & ~n21279;
  assign n21593 = ~n21270 & ~n21273;
  assign n21594 = n5267 & n20416;
  assign n21595 = n5185 & n20419;
  assign n21596 = n5121 & n20422;
  assign n21597 = n78 & n20771;
  assign n21598 = ~n21595 & ~n21596;
  assign n21599 = ~n21594 & n21598;
  assign n21600 = ~n21597 & n21599;
  assign n21601 = ~pi23  & ~n21600;
  assign n21602 = pi23  & n21600;
  assign n21603 = ~n21601 & ~n21602;
  assign n21604 = ~n21254 & ~n21257;
  assign n21605 = n4721 & n20425;
  assign n21606 = n4691 & n20428;
  assign n21607 = n4515 & n20431;
  assign n21608 = n4516 & n20727;
  assign n21609 = ~n21606 & ~n21607;
  assign n21610 = ~n21605 & n21609;
  assign n21611 = ~n21608 & n21610;
  assign n21612 = pi26  & n21611;
  assign n21613 = ~pi26  & ~n21611;
  assign n21614 = ~n21612 & ~n21613;
  assign n21615 = ~n21248 & ~n21251;
  assign n21616 = n4472 & n20434;
  assign n21617 = n4070 & n20437;
  assign n21618 = n3943 & n20440;
  assign n21619 = n3944 & n20668;
  assign n21620 = ~n21617 & ~n21618;
  assign n21621 = ~n21616 & n21620;
  assign n21622 = ~n21619 & n21621;
  assign n21623 = ~pi29  & ~n21622;
  assign n21624 = pi29  & n21622;
  assign n21625 = ~n21623 & ~n21624;
  assign n21626 = ~n250 & ~n321;
  assign n21627 = ~n389 & n21626;
  assign n21628 = n386 & n1117;
  assign n21629 = n1125 & n1243;
  assign n21630 = n1346 & n1760;
  assign n21631 = n5369 & n21630;
  assign n21632 = n21628 & n21629;
  assign n21633 = n21627 & n21632;
  assign n21634 = n21631 & n21633;
  assign n21635 = ~n126 & ~n175;
  assign n21636 = ~n221 & ~n234;
  assign n21637 = n21635 & n21636;
  assign n21638 = n309 & n603;
  assign n21639 = n1121 & n1233;
  assign n21640 = n1631 & n2903;
  assign n21641 = n3380 & n4156;
  assign n21642 = n21640 & n21641;
  assign n21643 = n21638 & n21639;
  assign n21644 = n576 & n21637;
  assign n21645 = n4770 & n21644;
  assign n21646 = n21642 & n21643;
  assign n21647 = n13141 & n21646;
  assign n21648 = n21645 & n21647;
  assign n21649 = ~n165 & ~n208;
  assign n21650 = ~n213 & ~n644;
  assign n21651 = ~n682 & n21650;
  assign n21652 = n1157 & n21649;
  assign n21653 = n1380 & n1904;
  assign n21654 = n21652 & n21653;
  assign n21655 = n2228 & n21651;
  assign n21656 = n2825 & n21655;
  assign n21657 = n1872 & n21654;
  assign n21658 = n7019 & n14739;
  assign n21659 = n21657 & n21658;
  assign n21660 = n21656 & n21659;
  assign n21661 = n21634 & n21660;
  assign n21662 = n14659 & n21648;
  assign n21663 = n21661 & n21662;
  assign n21664 = n3896 & n20445;
  assign n21665 = n3683 & n20447;
  assign n21666 = n566 & ~n20624;
  assign n21667 = ~n21664 & ~n21665;
  assign n21668 = ~n21666 & n21667;
  assign n21669 = ~n21663 & ~n21668;
  assign n21670 = n21663 & n21668;
  assign n21671 = ~n21669 & ~n21670;
  assign n21672 = ~n21625 & n21671;
  assign n21673 = n21625 & ~n21671;
  assign n21674 = ~n21672 & ~n21673;
  assign n21675 = ~n21615 & n21674;
  assign n21676 = n21615 & ~n21674;
  assign n21677 = ~n21675 & ~n21676;
  assign n21678 = ~n21614 & n21677;
  assign n21679 = n21614 & ~n21677;
  assign n21680 = ~n21678 & ~n21679;
  assign n21681 = ~n21604 & n21680;
  assign n21682 = n21604 & ~n21680;
  assign n21683 = ~n21681 & ~n21682;
  assign n21684 = ~n21603 & n21683;
  assign n21685 = n21603 & ~n21683;
  assign n21686 = ~n21684 & ~n21685;
  assign n21687 = n21593 & ~n21686;
  assign n21688 = ~n21593 & n21686;
  assign n21689 = ~n21687 & ~n21688;
  assign n21690 = n5982 & n20407;
  assign n21691 = n5901 & n20410;
  assign n21692 = n5312 & n20413;
  assign n21693 = n5306 & n21004;
  assign n21694 = ~n21691 & ~n21692;
  assign n21695 = ~n21690 & n21694;
  assign n21696 = ~n21693 & n21695;
  assign n21697 = pi20  & n21696;
  assign n21698 = ~pi20  & ~n21696;
  assign n21699 = ~n21697 & ~n21698;
  assign n21700 = n21689 & ~n21699;
  assign n21701 = ~n21689 & n21699;
  assign n21702 = ~n21700 & ~n21701;
  assign n21703 = ~n21592 & n21702;
  assign n21704 = n21592 & ~n21702;
  assign n21705 = ~n21703 & ~n21704;
  assign n21706 = ~n21591 & n21705;
  assign n21707 = n21591 & ~n21705;
  assign n21708 = ~n21706 & ~n21707;
  assign n21709 = ~n21581 & n21708;
  assign n21710 = n21581 & ~n21708;
  assign n21711 = ~n21709 & ~n21710;
  assign n21712 = n7380 & n20389;
  assign n21713 = n7243 & n20392;
  assign n21714 = n6653 & n20395;
  assign n21715 = n20512 & ~n20514;
  assign n21716 = ~n20515 & ~n21715;
  assign n21717 = n6647 & n21716;
  assign n21718 = ~n21713 & ~n21714;
  assign n21719 = ~n21712 & n21718;
  assign n21720 = ~n21717 & n21719;
  assign n21721 = pi14  & n21720;
  assign n21722 = ~pi14  & ~n21720;
  assign n21723 = ~n21721 & ~n21722;
  assign n21724 = n21711 & ~n21723;
  assign n21725 = ~n21711 & n21723;
  assign n21726 = ~n21724 & ~n21725;
  assign n21727 = ~n21580 & n21726;
  assign n21728 = n21580 & ~n21726;
  assign n21729 = ~n21727 & ~n21728;
  assign n21730 = ~n20581 & n21729;
  assign n21731 = n21576 & ~n21578;
  assign n21732 = ~n21579 & ~n21731;
  assign n21733 = n8161 & n20383;
  assign n21734 = n7847 & n20386;
  assign n21735 = n7554 & n20389;
  assign n21736 = n20520 & ~n20522;
  assign n21737 = ~n20523 & ~n21736;
  assign n21738 = n7548 & n21737;
  assign n21739 = ~n21734 & ~n21735;
  assign n21740 = ~n21733 & n21739;
  assign n21741 = ~n21738 & n21740;
  assign n21742 = pi11  & n21741;
  assign n21743 = ~pi11  & ~n21741;
  assign n21744 = ~n21742 & ~n21743;
  assign n21745 = n21732 & ~n21744;
  assign n21746 = n21572 & ~n21574;
  assign n21747 = ~n21575 & ~n21746;
  assign n21748 = n8161 & n20386;
  assign n21749 = n7847 & n20389;
  assign n21750 = n7554 & n20392;
  assign n21751 = n20516 & ~n20518;
  assign n21752 = ~n20519 & ~n21751;
  assign n21753 = n7548 & n21752;
  assign n21754 = ~n21749 & ~n21750;
  assign n21755 = ~n21748 & n21754;
  assign n21756 = ~n21753 & n21755;
  assign n21757 = pi11  & n21756;
  assign n21758 = ~pi11  & ~n21756;
  assign n21759 = ~n21757 & ~n21758;
  assign n21760 = n21747 & ~n21759;
  assign n21761 = n8161 & n20389;
  assign n21762 = n7847 & n20392;
  assign n21763 = n7554 & n20395;
  assign n21764 = n7548 & n21716;
  assign n21765 = ~n21762 & ~n21763;
  assign n21766 = ~n21761 & n21765;
  assign n21767 = ~n21764 & n21766;
  assign n21768 = ~pi11  & ~n21767;
  assign n21769 = pi11  & n21767;
  assign n21770 = ~n21768 & ~n21769;
  assign n21771 = n21568 & ~n21570;
  assign n21772 = ~n21571 & ~n21771;
  assign n21773 = ~n21770 & n21772;
  assign n21774 = n8161 & n20392;
  assign n21775 = n7847 & n20395;
  assign n21776 = n7554 & n20398;
  assign n21777 = n7548 & n20586;
  assign n21778 = ~n21775 & ~n21776;
  assign n21779 = ~n21774 & n21778;
  assign n21780 = ~n21777 & n21779;
  assign n21781 = ~pi11  & ~n21780;
  assign n21782 = pi11  & n21780;
  assign n21783 = ~n21781 & ~n21782;
  assign n21784 = n21564 & ~n21566;
  assign n21785 = ~n21567 & ~n21784;
  assign n21786 = ~n21783 & n21785;
  assign n21787 = n8161 & n20395;
  assign n21788 = n7847 & n20398;
  assign n21789 = n7554 & n20401;
  assign n21790 = n7548 & n21305;
  assign n21791 = ~n21788 & ~n21789;
  assign n21792 = ~n21787 & n21791;
  assign n21793 = ~n21790 & n21792;
  assign n21794 = ~pi11  & ~n21793;
  assign n21795 = pi11  & n21793;
  assign n21796 = ~n21794 & ~n21795;
  assign n21797 = n21560 & ~n21562;
  assign n21798 = ~n21563 & ~n21797;
  assign n21799 = ~n21796 & n21798;
  assign n21800 = n21556 & ~n21558;
  assign n21801 = ~n21559 & ~n21800;
  assign n21802 = n8161 & n20398;
  assign n21803 = n7847 & n20401;
  assign n21804 = n7554 & n20404;
  assign n21805 = n7548 & n21322;
  assign n21806 = ~n21803 & ~n21804;
  assign n21807 = ~n21802 & n21806;
  assign n21808 = ~n21805 & n21807;
  assign n21809 = pi11  & n21808;
  assign n21810 = ~pi11  & ~n21808;
  assign n21811 = ~n21809 & ~n21810;
  assign n21812 = n21801 & ~n21811;
  assign n21813 = n21552 & ~n21554;
  assign n21814 = ~n21555 & ~n21813;
  assign n21815 = n8161 & n20401;
  assign n21816 = n7847 & n20404;
  assign n21817 = n7554 & n20407;
  assign n21818 = n7548 & n21286;
  assign n21819 = ~n21816 & ~n21817;
  assign n21820 = ~n21815 & n21819;
  assign n21821 = ~n21818 & n21820;
  assign n21822 = pi11  & n21821;
  assign n21823 = ~pi11  & ~n21821;
  assign n21824 = ~n21822 & ~n21823;
  assign n21825 = n21814 & ~n21824;
  assign n21826 = n21548 & ~n21550;
  assign n21827 = ~n21551 & ~n21826;
  assign n21828 = n8161 & n20404;
  assign n21829 = n7847 & n20407;
  assign n21830 = n7554 & n20410;
  assign n21831 = n7548 & n20991;
  assign n21832 = ~n21829 & ~n21830;
  assign n21833 = ~n21828 & n21832;
  assign n21834 = ~n21831 & n21833;
  assign n21835 = pi11  & n21834;
  assign n21836 = ~pi11  & ~n21834;
  assign n21837 = ~n21835 & ~n21836;
  assign n21838 = n21827 & ~n21837;
  assign n21839 = n8161 & n20407;
  assign n21840 = n7847 & n20410;
  assign n21841 = n7554 & n20413;
  assign n21842 = n7548 & n21004;
  assign n21843 = ~n21840 & ~n21841;
  assign n21844 = ~n21839 & n21843;
  assign n21845 = ~n21842 & n21844;
  assign n21846 = ~pi11  & ~n21845;
  assign n21847 = pi11  & n21845;
  assign n21848 = ~n21846 & ~n21847;
  assign n21849 = n21544 & ~n21546;
  assign n21850 = ~n21547 & ~n21849;
  assign n21851 = ~n21848 & n21850;
  assign n21852 = n8161 & n20410;
  assign n21853 = n7847 & n20413;
  assign n21854 = n7554 & n20416;
  assign n21855 = n7548 & n21019;
  assign n21856 = ~n21853 & ~n21854;
  assign n21857 = ~n21852 & n21856;
  assign n21858 = ~n21855 & n21857;
  assign n21859 = ~pi11  & ~n21858;
  assign n21860 = pi11  & n21858;
  assign n21861 = ~n21859 & ~n21860;
  assign n21862 = n21540 & ~n21542;
  assign n21863 = ~n21543 & ~n21862;
  assign n21864 = ~n21861 & n21863;
  assign n21865 = n8161 & n20413;
  assign n21866 = n7847 & n20416;
  assign n21867 = n7554 & n20419;
  assign n21868 = n7548 & n20928;
  assign n21869 = ~n21866 & ~n21867;
  assign n21870 = ~n21865 & n21869;
  assign n21871 = ~n21868 & n21870;
  assign n21872 = ~pi11  & ~n21871;
  assign n21873 = pi11  & n21871;
  assign n21874 = ~n21872 & ~n21873;
  assign n21875 = n21536 & ~n21538;
  assign n21876 = ~n21539 & ~n21875;
  assign n21877 = ~n21874 & n21876;
  assign n21878 = n21532 & ~n21534;
  assign n21879 = ~n21535 & ~n21878;
  assign n21880 = n8161 & n20416;
  assign n21881 = n7847 & n20419;
  assign n21882 = n7554 & n20422;
  assign n21883 = n7548 & n20771;
  assign n21884 = ~n21881 & ~n21882;
  assign n21885 = ~n21880 & n21884;
  assign n21886 = ~n21883 & n21885;
  assign n21887 = pi11  & n21886;
  assign n21888 = ~pi11  & ~n21886;
  assign n21889 = ~n21887 & ~n21888;
  assign n21890 = n21879 & ~n21889;
  assign n21891 = n21528 & ~n21530;
  assign n21892 = ~n21531 & ~n21891;
  assign n21893 = n8161 & n20419;
  assign n21894 = n7847 & n20422;
  assign n21895 = n7554 & n20425;
  assign n21896 = n7548 & n20786;
  assign n21897 = ~n21894 & ~n21895;
  assign n21898 = ~n21893 & n21897;
  assign n21899 = ~n21896 & n21898;
  assign n21900 = pi11  & n21899;
  assign n21901 = ~pi11  & ~n21899;
  assign n21902 = ~n21900 & ~n21901;
  assign n21903 = n21892 & ~n21902;
  assign n21904 = n21524 & ~n21526;
  assign n21905 = ~n21527 & ~n21904;
  assign n21906 = n8161 & n20422;
  assign n21907 = n7847 & n20425;
  assign n21908 = n7554 & n20428;
  assign n21909 = n7548 & n20801;
  assign n21910 = ~n21907 & ~n21908;
  assign n21911 = ~n21906 & n21910;
  assign n21912 = ~n21909 & n21911;
  assign n21913 = pi11  & n21912;
  assign n21914 = ~pi11  & ~n21912;
  assign n21915 = ~n21913 & ~n21914;
  assign n21916 = n21905 & ~n21915;
  assign n21917 = n8161 & n20425;
  assign n21918 = n7847 & n20428;
  assign n21919 = n7554 & n20431;
  assign n21920 = n7548 & n20727;
  assign n21921 = ~n21918 & ~n21919;
  assign n21922 = ~n21917 & n21921;
  assign n21923 = ~n21920 & n21922;
  assign n21924 = ~pi11  & ~n21923;
  assign n21925 = pi11  & n21923;
  assign n21926 = ~n21924 & ~n21925;
  assign n21927 = n21520 & ~n21522;
  assign n21928 = ~n21523 & ~n21927;
  assign n21929 = ~n21926 & n21928;
  assign n21930 = n8161 & n20428;
  assign n21931 = n7847 & n20431;
  assign n21932 = n7554 & n20434;
  assign n21933 = n7548 & n20598;
  assign n21934 = ~n21931 & ~n21932;
  assign n21935 = ~n21930 & n21934;
  assign n21936 = ~n21933 & n21935;
  assign n21937 = pi11  & n21936;
  assign n21938 = ~pi11  & ~n21936;
  assign n21939 = ~n21937 & ~n21938;
  assign n21940 = n21516 & ~n21518;
  assign n21941 = ~n21519 & ~n21940;
  assign n21942 = ~n21939 & n21941;
  assign n21943 = n8161 & n20431;
  assign n21944 = n7847 & n20434;
  assign n21945 = n7554 & n20437;
  assign n21946 = n7548 & n20651;
  assign n21947 = ~n21944 & ~n21945;
  assign n21948 = ~n21943 & n21947;
  assign n21949 = ~n21946 & n21948;
  assign n21950 = ~pi11  & ~n21949;
  assign n21951 = pi11  & n21949;
  assign n21952 = ~n21950 & ~n21951;
  assign n21953 = pi14  & ~n21496;
  assign n21954 = n21503 & ~n21953;
  assign n21955 = ~n21503 & n21953;
  assign n21956 = ~n21954 & ~n21955;
  assign n21957 = ~n21952 & n21956;
  assign n21958 = n8161 & n20434;
  assign n21959 = n7847 & n20437;
  assign n21960 = n7554 & n20440;
  assign n21961 = n7548 & n20668;
  assign n21962 = ~n21959 & ~n21960;
  assign n21963 = ~n21958 & n21962;
  assign n21964 = ~n21961 & n21963;
  assign n21965 = pi11  & n21964;
  assign n21966 = ~pi11  & ~n21964;
  assign n21967 = ~n21965 & ~n21966;
  assign n21968 = n21490 & ~n21495;
  assign n21969 = ~n21496 & ~n21968;
  assign n21970 = ~n21967 & n21969;
  assign n21971 = n7547 & n20447;
  assign n21972 = pi11  & n21971;
  assign n21973 = n8161 & n20445;
  assign n21974 = n7847 & n20447;
  assign n21975 = n7548 & ~n20624;
  assign n21976 = ~n21973 & ~n21974;
  assign n21977 = ~n21975 & n21976;
  assign n21978 = ~n21972 & n21977;
  assign n21979 = n8161 & n20440;
  assign n21980 = n7847 & n20445;
  assign n21981 = n7554 & n20447;
  assign n21982 = n7548 & ~n20633;
  assign n21983 = ~n21980 & ~n21981;
  assign n21984 = ~n21979 & n21983;
  assign n21985 = ~n21982 & n21984;
  assign n21986 = pi11  & n21978;
  assign n21987 = n21985 & n21986;
  assign n21988 = n21489 & n21987;
  assign n21989 = n8161 & n20437;
  assign n21990 = n7847 & n20440;
  assign n21991 = n7554 & n20445;
  assign n21992 = n7548 & n20610;
  assign n21993 = ~n21990 & ~n21991;
  assign n21994 = ~n21989 & n21993;
  assign n21995 = ~n21992 & n21994;
  assign n21996 = pi11  & n21995;
  assign n21997 = ~pi11  & ~n21995;
  assign n21998 = ~n21996 & ~n21997;
  assign n21999 = ~n21489 & ~n21987;
  assign n22000 = ~n21988 & ~n21999;
  assign n22001 = ~n21998 & n22000;
  assign n22002 = ~n21988 & ~n22001;
  assign n22003 = n21967 & ~n21969;
  assign n22004 = ~n21970 & ~n22003;
  assign n22005 = ~n22002 & n22004;
  assign n22006 = ~n21970 & ~n22005;
  assign n22007 = n21952 & ~n21956;
  assign n22008 = ~n21957 & ~n22007;
  assign n22009 = ~n22006 & n22008;
  assign n22010 = ~n21957 & ~n22009;
  assign n22011 = n21939 & ~n21941;
  assign n22012 = ~n21942 & ~n22011;
  assign n22013 = ~n22010 & n22012;
  assign n22014 = ~n21942 & ~n22013;
  assign n22015 = n21926 & ~n21928;
  assign n22016 = ~n21929 & ~n22015;
  assign n22017 = ~n22014 & n22016;
  assign n22018 = ~n21929 & ~n22017;
  assign n22019 = ~n21905 & n21915;
  assign n22020 = ~n21916 & ~n22019;
  assign n22021 = ~n22018 & n22020;
  assign n22022 = ~n21916 & ~n22021;
  assign n22023 = ~n21892 & n21902;
  assign n22024 = ~n21903 & ~n22023;
  assign n22025 = ~n22022 & n22024;
  assign n22026 = ~n21903 & ~n22025;
  assign n22027 = ~n21879 & n21889;
  assign n22028 = ~n21890 & ~n22027;
  assign n22029 = ~n22026 & n22028;
  assign n22030 = ~n21890 & ~n22029;
  assign n22031 = n21874 & ~n21876;
  assign n22032 = ~n21877 & ~n22031;
  assign n22033 = ~n22030 & n22032;
  assign n22034 = ~n21877 & ~n22033;
  assign n22035 = n21861 & ~n21863;
  assign n22036 = ~n21864 & ~n22035;
  assign n22037 = ~n22034 & n22036;
  assign n22038 = ~n21864 & ~n22037;
  assign n22039 = n21848 & ~n21850;
  assign n22040 = ~n21851 & ~n22039;
  assign n22041 = ~n22038 & n22040;
  assign n22042 = ~n21851 & ~n22041;
  assign n22043 = ~n21827 & n21837;
  assign n22044 = ~n21838 & ~n22043;
  assign n22045 = ~n22042 & n22044;
  assign n22046 = ~n21838 & ~n22045;
  assign n22047 = ~n21814 & n21824;
  assign n22048 = ~n21825 & ~n22047;
  assign n22049 = ~n22046 & n22048;
  assign n22050 = ~n21825 & ~n22049;
  assign n22051 = ~n21801 & n21811;
  assign n22052 = ~n21812 & ~n22051;
  assign n22053 = ~n22050 & n22052;
  assign n22054 = ~n21812 & ~n22053;
  assign n22055 = n21796 & ~n21798;
  assign n22056 = ~n21799 & ~n22055;
  assign n22057 = ~n22054 & n22056;
  assign n22058 = ~n21799 & ~n22057;
  assign n22059 = n21783 & ~n21785;
  assign n22060 = ~n21786 & ~n22059;
  assign n22061 = ~n22058 & n22060;
  assign n22062 = ~n21786 & ~n22061;
  assign n22063 = n21770 & ~n21772;
  assign n22064 = ~n21773 & ~n22063;
  assign n22065 = ~n22062 & n22064;
  assign n22066 = ~n21773 & ~n22065;
  assign n22067 = ~n21747 & n21759;
  assign n22068 = ~n21760 & ~n22067;
  assign n22069 = ~n22066 & n22068;
  assign n22070 = ~n21760 & ~n22069;
  assign n22071 = ~n21732 & n21744;
  assign n22072 = ~n21745 & ~n22071;
  assign n22073 = ~n22070 & n22072;
  assign n22074 = ~n21745 & ~n22073;
  assign n22075 = n20581 & ~n21729;
  assign n22076 = ~n21730 & ~n22075;
  assign n22077 = ~n22074 & n22076;
  assign n22078 = ~n21730 & ~n22077;
  assign n22079 = n8161 & n20377;
  assign n22080 = n7847 & n20380;
  assign n22081 = n7554 & n20383;
  assign n22082 = n20528 & ~n20530;
  assign n22083 = ~n20531 & ~n22082;
  assign n22084 = n7548 & n22083;
  assign n22085 = ~n22080 & ~n22081;
  assign n22086 = ~n22079 & n22085;
  assign n22087 = ~n22084 & n22086;
  assign n22088 = ~pi11  & ~n22087;
  assign n22089 = pi11  & n22087;
  assign n22090 = ~n22088 & ~n22089;
  assign n22091 = ~n21724 & ~n21727;
  assign n22092 = ~n21706 & ~n21709;
  assign n22093 = n6608 & n20395;
  assign n22094 = n6356 & n20398;
  assign n22095 = n6140 & n20401;
  assign n22096 = n6134 & n21305;
  assign n22097 = ~n22094 & ~n22095;
  assign n22098 = ~n22093 & n22097;
  assign n22099 = ~n22096 & n22098;
  assign n22100 = ~pi17  & ~n22099;
  assign n22101 = pi17  & n22099;
  assign n22102 = ~n22100 & ~n22101;
  assign n22103 = ~n21700 & ~n21703;
  assign n22104 = ~n21684 & ~n21688;
  assign n22105 = n5267 & n20413;
  assign n22106 = n5185 & n20416;
  assign n22107 = n5121 & n20419;
  assign n22108 = n78 & n20928;
  assign n22109 = ~n22106 & ~n22107;
  assign n22110 = ~n22105 & n22109;
  assign n22111 = ~n22108 & n22110;
  assign n22112 = ~pi23  & ~n22111;
  assign n22113 = pi23  & n22111;
  assign n22114 = ~n22112 & ~n22113;
  assign n22115 = ~n21678 & ~n21681;
  assign n22116 = ~n21672 & ~n21675;
  assign n22117 = n4472 & n20431;
  assign n22118 = n4070 & n20434;
  assign n22119 = n3943 & n20437;
  assign n22120 = n3944 & n20651;
  assign n22121 = ~n22118 & ~n22119;
  assign n22122 = ~n22117 & n22121;
  assign n22123 = ~n22120 & n22122;
  assign n22124 = ~pi29  & ~n22123;
  assign n22125 = pi29  & n22123;
  assign n22126 = ~n22124 & ~n22125;
  assign n22127 = ~n162 & ~n290;
  assign n22128 = ~n446 & n22127;
  assign n22129 = ~n250 & ~n382;
  assign n22130 = ~n492 & ~n683;
  assign n22131 = n22129 & n22130;
  assign n22132 = n150 & n742;
  assign n22133 = n1356 & n1689;
  assign n22134 = n1969 & n5002;
  assign n22135 = n12716 & n22134;
  assign n22136 = n22132 & n22133;
  assign n22137 = n22128 & n22131;
  assign n22138 = n22136 & n22137;
  assign n22139 = n1867 & n22135;
  assign n22140 = n4146 & n4582;
  assign n22141 = n22139 & n22140;
  assign n22142 = n5696 & n22138;
  assign n22143 = n22141 & n22142;
  assign n22144 = n6950 & n22143;
  assign n22145 = n14659 & n22144;
  assign n22146 = n21669 & ~n22145;
  assign n22147 = ~n21669 & n22145;
  assign n22148 = ~n22146 & ~n22147;
  assign n22149 = n3896 & n20440;
  assign n22150 = n3683 & n20445;
  assign n22151 = n564 & n20447;
  assign n22152 = n566 & ~n20633;
  assign n22153 = ~n22150 & ~n22151;
  assign n22154 = ~n22149 & n22153;
  assign n22155 = ~n22152 & n22154;
  assign n22156 = n22148 & ~n22155;
  assign n22157 = ~n22148 & n22155;
  assign n22158 = ~n22156 & ~n22157;
  assign n22159 = ~n22126 & n22158;
  assign n22160 = n22126 & ~n22158;
  assign n22161 = ~n22159 & ~n22160;
  assign n22162 = n22116 & ~n22161;
  assign n22163 = ~n22116 & n22161;
  assign n22164 = ~n22162 & ~n22163;
  assign n22165 = n4721 & n20422;
  assign n22166 = n4691 & n20425;
  assign n22167 = n4515 & n20428;
  assign n22168 = n4516 & n20801;
  assign n22169 = ~n22166 & ~n22167;
  assign n22170 = ~n22165 & n22169;
  assign n22171 = ~n22168 & n22170;
  assign n22172 = pi26  & n22171;
  assign n22173 = ~pi26  & ~n22171;
  assign n22174 = ~n22172 & ~n22173;
  assign n22175 = n22164 & ~n22174;
  assign n22176 = ~n22164 & n22174;
  assign n22177 = ~n22175 & ~n22176;
  assign n22178 = ~n22115 & n22177;
  assign n22179 = n22115 & ~n22177;
  assign n22180 = ~n22178 & ~n22179;
  assign n22181 = ~n22114 & n22180;
  assign n22182 = n22114 & ~n22180;
  assign n22183 = ~n22181 & ~n22182;
  assign n22184 = n22104 & ~n22183;
  assign n22185 = ~n22104 & n22183;
  assign n22186 = ~n22184 & ~n22185;
  assign n22187 = n5982 & n20404;
  assign n22188 = n5901 & n20407;
  assign n22189 = n5312 & n20410;
  assign n22190 = n5306 & n20991;
  assign n22191 = ~n22188 & ~n22189;
  assign n22192 = ~n22187 & n22191;
  assign n22193 = ~n22190 & n22192;
  assign n22194 = pi20  & n22193;
  assign n22195 = ~pi20  & ~n22193;
  assign n22196 = ~n22194 & ~n22195;
  assign n22197 = n22186 & ~n22196;
  assign n22198 = ~n22186 & n22196;
  assign n22199 = ~n22197 & ~n22198;
  assign n22200 = ~n22103 & n22199;
  assign n22201 = n22103 & ~n22199;
  assign n22202 = ~n22200 & ~n22201;
  assign n22203 = ~n22102 & n22202;
  assign n22204 = n22102 & ~n22202;
  assign n22205 = ~n22203 & ~n22204;
  assign n22206 = n22092 & ~n22205;
  assign n22207 = ~n22092 & n22205;
  assign n22208 = ~n22206 & ~n22207;
  assign n22209 = n7380 & n20386;
  assign n22210 = n7243 & n20389;
  assign n22211 = n6653 & n20392;
  assign n22212 = n6647 & n21752;
  assign n22213 = ~n22210 & ~n22211;
  assign n22214 = ~n22209 & n22213;
  assign n22215 = ~n22212 & n22214;
  assign n22216 = pi14  & n22215;
  assign n22217 = ~pi14  & ~n22215;
  assign n22218 = ~n22216 & ~n22217;
  assign n22219 = n22208 & ~n22218;
  assign n22220 = ~n22208 & n22218;
  assign n22221 = ~n22219 & ~n22220;
  assign n22222 = ~n22091 & n22221;
  assign n22223 = n22091 & ~n22221;
  assign n22224 = ~n22222 & ~n22223;
  assign n22225 = ~n22090 & n22224;
  assign n22226 = n22090 & ~n22224;
  assign n22227 = ~n22225 & ~n22226;
  assign n22228 = ~n22078 & n22227;
  assign n22229 = n22078 & ~n22227;
  assign n22230 = ~n22228 & ~n22229;
  assign n22231 = n9355 & n20368;
  assign n22232 = n8939 & n20371;
  assign n22233 = n8206 & n20374;
  assign n22234 = n20540 & ~n20542;
  assign n22235 = ~n20543 & ~n22234;
  assign n22236 = n8200 & n22235;
  assign n22237 = ~n22232 & ~n22233;
  assign n22238 = ~n22231 & n22237;
  assign n22239 = ~n22236 & n22238;
  assign n22240 = pi8  & n22239;
  assign n22241 = ~pi8  & ~n22239;
  assign n22242 = ~n22240 & ~n22241;
  assign n22243 = n22230 & ~n22242;
  assign n22244 = n22074 & ~n22076;
  assign n22245 = ~n22077 & ~n22244;
  assign n22246 = n9355 & n20371;
  assign n22247 = n8939 & n20374;
  assign n22248 = n8206 & n20377;
  assign n22249 = n20536 & ~n20538;
  assign n22250 = ~n20539 & ~n22249;
  assign n22251 = n8200 & n22250;
  assign n22252 = ~n22247 & ~n22248;
  assign n22253 = ~n22246 & n22252;
  assign n22254 = ~n22251 & n22253;
  assign n22255 = pi8  & n22254;
  assign n22256 = ~pi8  & ~n22254;
  assign n22257 = ~n22255 & ~n22256;
  assign n22258 = n22245 & ~n22257;
  assign n22259 = n9355 & n20374;
  assign n22260 = n8939 & n20377;
  assign n22261 = n8206 & n20380;
  assign n22262 = n20532 & ~n20534;
  assign n22263 = ~n20535 & ~n22262;
  assign n22264 = n8200 & n22263;
  assign n22265 = ~n22260 & ~n22261;
  assign n22266 = ~n22259 & n22265;
  assign n22267 = ~n22264 & n22266;
  assign n22268 = ~pi8  & ~n22267;
  assign n22269 = pi8  & n22267;
  assign n22270 = ~n22268 & ~n22269;
  assign n22271 = n22070 & ~n22072;
  assign n22272 = ~n22073 & ~n22271;
  assign n22273 = ~n22270 & n22272;
  assign n22274 = n9355 & n20377;
  assign n22275 = n8939 & n20380;
  assign n22276 = n8206 & n20383;
  assign n22277 = n8200 & n22083;
  assign n22278 = ~n22275 & ~n22276;
  assign n22279 = ~n22274 & n22278;
  assign n22280 = ~n22277 & n22279;
  assign n22281 = ~pi8  & ~n22280;
  assign n22282 = pi8  & n22280;
  assign n22283 = ~n22281 & ~n22282;
  assign n22284 = n22066 & ~n22068;
  assign n22285 = ~n22069 & ~n22284;
  assign n22286 = ~n22283 & n22285;
  assign n22287 = n22062 & ~n22064;
  assign n22288 = ~n22065 & ~n22287;
  assign n22289 = n9355 & n20380;
  assign n22290 = n8939 & n20383;
  assign n22291 = n8206 & n20386;
  assign n22292 = n8200 & n20574;
  assign n22293 = ~n22290 & ~n22291;
  assign n22294 = ~n22289 & n22293;
  assign n22295 = ~n22292 & n22294;
  assign n22296 = pi8  & n22295;
  assign n22297 = ~pi8  & ~n22295;
  assign n22298 = ~n22296 & ~n22297;
  assign n22299 = n22288 & ~n22298;
  assign n22300 = n22058 & ~n22060;
  assign n22301 = ~n22061 & ~n22300;
  assign n22302 = n9355 & n20383;
  assign n22303 = n8939 & n20386;
  assign n22304 = n8206 & n20389;
  assign n22305 = n8200 & n21737;
  assign n22306 = ~n22303 & ~n22304;
  assign n22307 = ~n22302 & n22306;
  assign n22308 = ~n22305 & n22307;
  assign n22309 = pi8  & n22308;
  assign n22310 = ~pi8  & ~n22308;
  assign n22311 = ~n22309 & ~n22310;
  assign n22312 = n22301 & ~n22311;
  assign n22313 = n22054 & ~n22056;
  assign n22314 = ~n22057 & ~n22313;
  assign n22315 = n9355 & n20386;
  assign n22316 = n8939 & n20389;
  assign n22317 = n8206 & n20392;
  assign n22318 = n8200 & n21752;
  assign n22319 = ~n22316 & ~n22317;
  assign n22320 = ~n22315 & n22319;
  assign n22321 = ~n22318 & n22320;
  assign n22322 = pi8  & n22321;
  assign n22323 = ~pi8  & ~n22321;
  assign n22324 = ~n22322 & ~n22323;
  assign n22325 = n22314 & ~n22324;
  assign n22326 = n9355 & n20389;
  assign n22327 = n8939 & n20392;
  assign n22328 = n8206 & n20395;
  assign n22329 = n8200 & n21716;
  assign n22330 = ~n22327 & ~n22328;
  assign n22331 = ~n22326 & n22330;
  assign n22332 = ~n22329 & n22331;
  assign n22333 = ~pi8  & ~n22332;
  assign n22334 = pi8  & n22332;
  assign n22335 = ~n22333 & ~n22334;
  assign n22336 = n22050 & ~n22052;
  assign n22337 = ~n22053 & ~n22336;
  assign n22338 = ~n22335 & n22337;
  assign n22339 = n9355 & n20392;
  assign n22340 = n8939 & n20395;
  assign n22341 = n8206 & n20398;
  assign n22342 = n8200 & n20586;
  assign n22343 = ~n22340 & ~n22341;
  assign n22344 = ~n22339 & n22343;
  assign n22345 = ~n22342 & n22344;
  assign n22346 = ~pi8  & ~n22345;
  assign n22347 = pi8  & n22345;
  assign n22348 = ~n22346 & ~n22347;
  assign n22349 = n22046 & ~n22048;
  assign n22350 = ~n22049 & ~n22349;
  assign n22351 = ~n22348 & n22350;
  assign n22352 = n9355 & n20395;
  assign n22353 = n8939 & n20398;
  assign n22354 = n8206 & n20401;
  assign n22355 = n8200 & n21305;
  assign n22356 = ~n22353 & ~n22354;
  assign n22357 = ~n22352 & n22356;
  assign n22358 = ~n22355 & n22357;
  assign n22359 = ~pi8  & ~n22358;
  assign n22360 = pi8  & n22358;
  assign n22361 = ~n22359 & ~n22360;
  assign n22362 = n22042 & ~n22044;
  assign n22363 = ~n22045 & ~n22362;
  assign n22364 = ~n22361 & n22363;
  assign n22365 = n22038 & ~n22040;
  assign n22366 = ~n22041 & ~n22365;
  assign n22367 = n9355 & n20398;
  assign n22368 = n8939 & n20401;
  assign n22369 = n8206 & n20404;
  assign n22370 = n8200 & n21322;
  assign n22371 = ~n22368 & ~n22369;
  assign n22372 = ~n22367 & n22371;
  assign n22373 = ~n22370 & n22372;
  assign n22374 = pi8  & n22373;
  assign n22375 = ~pi8  & ~n22373;
  assign n22376 = ~n22374 & ~n22375;
  assign n22377 = n22366 & ~n22376;
  assign n22378 = n22034 & ~n22036;
  assign n22379 = ~n22037 & ~n22378;
  assign n22380 = n9355 & n20401;
  assign n22381 = n8939 & n20404;
  assign n22382 = n8206 & n20407;
  assign n22383 = n8200 & n21286;
  assign n22384 = ~n22381 & ~n22382;
  assign n22385 = ~n22380 & n22384;
  assign n22386 = ~n22383 & n22385;
  assign n22387 = pi8  & n22386;
  assign n22388 = ~pi8  & ~n22386;
  assign n22389 = ~n22387 & ~n22388;
  assign n22390 = n22379 & ~n22389;
  assign n22391 = n22030 & ~n22032;
  assign n22392 = ~n22033 & ~n22391;
  assign n22393 = n9355 & n20404;
  assign n22394 = n8939 & n20407;
  assign n22395 = n8206 & n20410;
  assign n22396 = n8200 & n20991;
  assign n22397 = ~n22394 & ~n22395;
  assign n22398 = ~n22393 & n22397;
  assign n22399 = ~n22396 & n22398;
  assign n22400 = pi8  & n22399;
  assign n22401 = ~pi8  & ~n22399;
  assign n22402 = ~n22400 & ~n22401;
  assign n22403 = n22392 & ~n22402;
  assign n22404 = n9355 & n20407;
  assign n22405 = n8939 & n20410;
  assign n22406 = n8206 & n20413;
  assign n22407 = n8200 & n21004;
  assign n22408 = ~n22405 & ~n22406;
  assign n22409 = ~n22404 & n22408;
  assign n22410 = ~n22407 & n22409;
  assign n22411 = ~pi8  & ~n22410;
  assign n22412 = pi8  & n22410;
  assign n22413 = ~n22411 & ~n22412;
  assign n22414 = n22026 & ~n22028;
  assign n22415 = ~n22029 & ~n22414;
  assign n22416 = ~n22413 & n22415;
  assign n22417 = n9355 & n20410;
  assign n22418 = n8939 & n20413;
  assign n22419 = n8206 & n20416;
  assign n22420 = n8200 & n21019;
  assign n22421 = ~n22418 & ~n22419;
  assign n22422 = ~n22417 & n22421;
  assign n22423 = ~n22420 & n22422;
  assign n22424 = ~pi8  & ~n22423;
  assign n22425 = pi8  & n22423;
  assign n22426 = ~n22424 & ~n22425;
  assign n22427 = n22022 & ~n22024;
  assign n22428 = ~n22025 & ~n22427;
  assign n22429 = ~n22426 & n22428;
  assign n22430 = n9355 & n20413;
  assign n22431 = n8939 & n20416;
  assign n22432 = n8206 & n20419;
  assign n22433 = n8200 & n20928;
  assign n22434 = ~n22431 & ~n22432;
  assign n22435 = ~n22430 & n22434;
  assign n22436 = ~n22433 & n22435;
  assign n22437 = ~pi8  & ~n22436;
  assign n22438 = pi8  & n22436;
  assign n22439 = ~n22437 & ~n22438;
  assign n22440 = n22018 & ~n22020;
  assign n22441 = ~n22021 & ~n22440;
  assign n22442 = ~n22439 & n22441;
  assign n22443 = n22014 & ~n22016;
  assign n22444 = ~n22017 & ~n22443;
  assign n22445 = n9355 & n20416;
  assign n22446 = n8939 & n20419;
  assign n22447 = n8206 & n20422;
  assign n22448 = n8200 & n20771;
  assign n22449 = ~n22446 & ~n22447;
  assign n22450 = ~n22445 & n22449;
  assign n22451 = ~n22448 & n22450;
  assign n22452 = pi8  & n22451;
  assign n22453 = ~pi8  & ~n22451;
  assign n22454 = ~n22452 & ~n22453;
  assign n22455 = n22444 & ~n22454;
  assign n22456 = n22010 & ~n22012;
  assign n22457 = ~n22013 & ~n22456;
  assign n22458 = n9355 & n20419;
  assign n22459 = n8939 & n20422;
  assign n22460 = n8206 & n20425;
  assign n22461 = n8200 & n20786;
  assign n22462 = ~n22459 & ~n22460;
  assign n22463 = ~n22458 & n22462;
  assign n22464 = ~n22461 & n22463;
  assign n22465 = pi8  & n22464;
  assign n22466 = ~pi8  & ~n22464;
  assign n22467 = ~n22465 & ~n22466;
  assign n22468 = n22457 & ~n22467;
  assign n22469 = n22006 & ~n22008;
  assign n22470 = ~n22009 & ~n22469;
  assign n22471 = n9355 & n20422;
  assign n22472 = n8939 & n20425;
  assign n22473 = n8206 & n20428;
  assign n22474 = n8200 & n20801;
  assign n22475 = ~n22472 & ~n22473;
  assign n22476 = ~n22471 & n22475;
  assign n22477 = ~n22474 & n22476;
  assign n22478 = pi8  & n22477;
  assign n22479 = ~pi8  & ~n22477;
  assign n22480 = ~n22478 & ~n22479;
  assign n22481 = n22470 & ~n22480;
  assign n22482 = n9355 & n20425;
  assign n22483 = n8939 & n20428;
  assign n22484 = n8206 & n20431;
  assign n22485 = n8200 & n20727;
  assign n22486 = ~n22483 & ~n22484;
  assign n22487 = ~n22482 & n22486;
  assign n22488 = ~n22485 & n22487;
  assign n22489 = ~pi8  & ~n22488;
  assign n22490 = pi8  & n22488;
  assign n22491 = ~n22489 & ~n22490;
  assign n22492 = n22002 & ~n22004;
  assign n22493 = ~n22005 & ~n22492;
  assign n22494 = ~n22491 & n22493;
  assign n22495 = n9355 & n20428;
  assign n22496 = n8939 & n20431;
  assign n22497 = n8206 & n20434;
  assign n22498 = n8200 & n20598;
  assign n22499 = ~n22496 & ~n22497;
  assign n22500 = ~n22495 & n22499;
  assign n22501 = ~n22498 & n22500;
  assign n22502 = pi8  & n22501;
  assign n22503 = ~pi8  & ~n22501;
  assign n22504 = ~n22502 & ~n22503;
  assign n22505 = n21998 & ~n22000;
  assign n22506 = ~n22001 & ~n22505;
  assign n22507 = ~n22504 & n22506;
  assign n22508 = n9355 & n20431;
  assign n22509 = n8939 & n20434;
  assign n22510 = n8206 & n20437;
  assign n22511 = n8200 & n20651;
  assign n22512 = ~n22509 & ~n22510;
  assign n22513 = ~n22508 & n22512;
  assign n22514 = ~n22511 & n22513;
  assign n22515 = ~pi8  & ~n22514;
  assign n22516 = pi8  & n22514;
  assign n22517 = ~n22515 & ~n22516;
  assign n22518 = pi11  & ~n21978;
  assign n22519 = n21985 & ~n22518;
  assign n22520 = ~n21985 & n22518;
  assign n22521 = ~n22519 & ~n22520;
  assign n22522 = ~n22517 & n22521;
  assign n22523 = n9355 & n20434;
  assign n22524 = n8939 & n20437;
  assign n22525 = n8206 & n20440;
  assign n22526 = n8200 & n20668;
  assign n22527 = ~n22524 & ~n22525;
  assign n22528 = ~n22523 & n22527;
  assign n22529 = ~n22526 & n22528;
  assign n22530 = pi8  & n22529;
  assign n22531 = ~pi8  & ~n22529;
  assign n22532 = ~n22530 & ~n22531;
  assign n22533 = n21972 & ~n21977;
  assign n22534 = ~n21978 & ~n22533;
  assign n22535 = ~n22532 & n22534;
  assign n22536 = n8199 & n20447;
  assign n22537 = pi8  & n22536;
  assign n22538 = n9355 & n20445;
  assign n22539 = n8939 & n20447;
  assign n22540 = n8200 & ~n20624;
  assign n22541 = ~n22538 & ~n22539;
  assign n22542 = ~n22540 & n22541;
  assign n22543 = ~n22537 & n22542;
  assign n22544 = n9355 & n20440;
  assign n22545 = n8939 & n20445;
  assign n22546 = n8206 & n20447;
  assign n22547 = n8200 & ~n20633;
  assign n22548 = ~n22545 & ~n22546;
  assign n22549 = ~n22544 & n22548;
  assign n22550 = ~n22547 & n22549;
  assign n22551 = pi8  & n22543;
  assign n22552 = n22550 & n22551;
  assign n22553 = n21971 & n22552;
  assign n22554 = n9355 & n20437;
  assign n22555 = n8939 & n20440;
  assign n22556 = n8206 & n20445;
  assign n22557 = n8200 & n20610;
  assign n22558 = ~n22555 & ~n22556;
  assign n22559 = ~n22554 & n22558;
  assign n22560 = ~n22557 & n22559;
  assign n22561 = pi8  & n22560;
  assign n22562 = ~pi8  & ~n22560;
  assign n22563 = ~n22561 & ~n22562;
  assign n22564 = ~n21971 & ~n22552;
  assign n22565 = ~n22553 & ~n22564;
  assign n22566 = ~n22563 & n22565;
  assign n22567 = ~n22553 & ~n22566;
  assign n22568 = n22532 & ~n22534;
  assign n22569 = ~n22535 & ~n22568;
  assign n22570 = ~n22567 & n22569;
  assign n22571 = ~n22535 & ~n22570;
  assign n22572 = n22517 & ~n22521;
  assign n22573 = ~n22522 & ~n22572;
  assign n22574 = ~n22571 & n22573;
  assign n22575 = ~n22522 & ~n22574;
  assign n22576 = n22504 & ~n22506;
  assign n22577 = ~n22507 & ~n22576;
  assign n22578 = ~n22575 & n22577;
  assign n22579 = ~n22507 & ~n22578;
  assign n22580 = n22491 & ~n22493;
  assign n22581 = ~n22494 & ~n22580;
  assign n22582 = ~n22579 & n22581;
  assign n22583 = ~n22494 & ~n22582;
  assign n22584 = ~n22470 & n22480;
  assign n22585 = ~n22481 & ~n22584;
  assign n22586 = ~n22583 & n22585;
  assign n22587 = ~n22481 & ~n22586;
  assign n22588 = ~n22457 & n22467;
  assign n22589 = ~n22468 & ~n22588;
  assign n22590 = ~n22587 & n22589;
  assign n22591 = ~n22468 & ~n22590;
  assign n22592 = ~n22444 & n22454;
  assign n22593 = ~n22455 & ~n22592;
  assign n22594 = ~n22591 & n22593;
  assign n22595 = ~n22455 & ~n22594;
  assign n22596 = n22439 & ~n22441;
  assign n22597 = ~n22442 & ~n22596;
  assign n22598 = ~n22595 & n22597;
  assign n22599 = ~n22442 & ~n22598;
  assign n22600 = n22426 & ~n22428;
  assign n22601 = ~n22429 & ~n22600;
  assign n22602 = ~n22599 & n22601;
  assign n22603 = ~n22429 & ~n22602;
  assign n22604 = n22413 & ~n22415;
  assign n22605 = ~n22416 & ~n22604;
  assign n22606 = ~n22603 & n22605;
  assign n22607 = ~n22416 & ~n22606;
  assign n22608 = ~n22392 & n22402;
  assign n22609 = ~n22403 & ~n22608;
  assign n22610 = ~n22607 & n22609;
  assign n22611 = ~n22403 & ~n22610;
  assign n22612 = ~n22379 & n22389;
  assign n22613 = ~n22390 & ~n22612;
  assign n22614 = ~n22611 & n22613;
  assign n22615 = ~n22390 & ~n22614;
  assign n22616 = ~n22366 & n22376;
  assign n22617 = ~n22377 & ~n22616;
  assign n22618 = ~n22615 & n22617;
  assign n22619 = ~n22377 & ~n22618;
  assign n22620 = n22361 & ~n22363;
  assign n22621 = ~n22364 & ~n22620;
  assign n22622 = ~n22619 & n22621;
  assign n22623 = ~n22364 & ~n22622;
  assign n22624 = n22348 & ~n22350;
  assign n22625 = ~n22351 & ~n22624;
  assign n22626 = ~n22623 & n22625;
  assign n22627 = ~n22351 & ~n22626;
  assign n22628 = n22335 & ~n22337;
  assign n22629 = ~n22338 & ~n22628;
  assign n22630 = ~n22627 & n22629;
  assign n22631 = ~n22338 & ~n22630;
  assign n22632 = ~n22314 & n22324;
  assign n22633 = ~n22325 & ~n22632;
  assign n22634 = ~n22631 & n22633;
  assign n22635 = ~n22325 & ~n22634;
  assign n22636 = ~n22301 & n22311;
  assign n22637 = ~n22312 & ~n22636;
  assign n22638 = ~n22635 & n22637;
  assign n22639 = ~n22312 & ~n22638;
  assign n22640 = ~n22288 & n22298;
  assign n22641 = ~n22299 & ~n22640;
  assign n22642 = ~n22639 & n22641;
  assign n22643 = ~n22299 & ~n22642;
  assign n22644 = n22283 & ~n22285;
  assign n22645 = ~n22286 & ~n22644;
  assign n22646 = ~n22643 & n22645;
  assign n22647 = ~n22286 & ~n22646;
  assign n22648 = n22270 & ~n22272;
  assign n22649 = ~n22273 & ~n22648;
  assign n22650 = ~n22647 & n22649;
  assign n22651 = ~n22273 & ~n22650;
  assign n22652 = ~n22245 & n22257;
  assign n22653 = ~n22258 & ~n22652;
  assign n22654 = ~n22651 & n22653;
  assign n22655 = ~n22258 & ~n22654;
  assign n22656 = ~n22230 & n22242;
  assign n22657 = ~n22243 & ~n22656;
  assign n22658 = ~n22655 & n22657;
  assign n22659 = ~n22243 & ~n22658;
  assign n22660 = ~n22225 & ~n22228;
  assign n22661 = n8161 & n20374;
  assign n22662 = n7847 & n20377;
  assign n22663 = n7554 & n20380;
  assign n22664 = n7548 & n22263;
  assign n22665 = ~n22662 & ~n22663;
  assign n22666 = ~n22661 & n22665;
  assign n22667 = ~n22664 & n22666;
  assign n22668 = ~pi11  & ~n22667;
  assign n22669 = pi11  & n22667;
  assign n22670 = ~n22668 & ~n22669;
  assign n22671 = ~n22219 & ~n22222;
  assign n22672 = ~n22203 & ~n22207;
  assign n22673 = n6608 & n20392;
  assign n22674 = n6356 & n20395;
  assign n22675 = n6140 & n20398;
  assign n22676 = n6134 & n20586;
  assign n22677 = ~n22674 & ~n22675;
  assign n22678 = ~n22673 & n22677;
  assign n22679 = ~n22676 & n22678;
  assign n22680 = ~pi17  & ~n22679;
  assign n22681 = pi17  & n22679;
  assign n22682 = ~n22680 & ~n22681;
  assign n22683 = ~n22197 & ~n22200;
  assign n22684 = ~n22181 & ~n22185;
  assign n22685 = n5267 & n20410;
  assign n22686 = n5185 & n20413;
  assign n22687 = n5121 & n20416;
  assign n22688 = n78 & n21019;
  assign n22689 = ~n22686 & ~n22687;
  assign n22690 = ~n22685 & n22689;
  assign n22691 = ~n22688 & n22690;
  assign n22692 = ~pi23  & ~n22691;
  assign n22693 = pi23  & n22691;
  assign n22694 = ~n22692 & ~n22693;
  assign n22695 = ~n22175 & ~n22178;
  assign n22696 = ~n22159 & ~n22163;
  assign n22697 = n4472 & n20428;
  assign n22698 = n4070 & n20431;
  assign n22699 = n3943 & n20434;
  assign n22700 = n3944 & n20598;
  assign n22701 = ~n22698 & ~n22699;
  assign n22702 = ~n22697 & n22701;
  assign n22703 = ~n22700 & n22702;
  assign n22704 = ~pi29  & ~n22703;
  assign n22705 = pi29  & n22703;
  assign n22706 = ~n22704 & ~n22705;
  assign n22707 = ~n22146 & ~n22156;
  assign n22708 = ~n287 & ~n690;
  assign n22709 = n969 & n22708;
  assign n22710 = ~n243 & ~n447;
  assign n22711 = n166 & n22710;
  assign n22712 = n464 & n524;
  assign n22713 = n731 & n940;
  assign n22714 = n2660 & n3628;
  assign n22715 = n5550 & n22714;
  assign n22716 = n22712 & n22713;
  assign n22717 = n22709 & n22711;
  assign n22718 = n22716 & n22717;
  assign n22719 = n2379 & n22715;
  assign n22720 = n22718 & n22719;
  assign n22721 = n4568 & n5795;
  assign n22722 = n22720 & n22721;
  assign n22723 = n1779 & n22722;
  assign n22724 = n2696 & n22723;
  assign n22725 = n3896 & n20437;
  assign n22726 = n564 & n20445;
  assign n22727 = n3683 & n20440;
  assign n22728 = n566 & n20610;
  assign n22729 = ~n22726 & ~n22727;
  assign n22730 = ~n22725 & n22729;
  assign n22731 = ~n22728 & n22730;
  assign n22732 = ~n22724 & ~n22731;
  assign n22733 = n22724 & n22731;
  assign n22734 = ~n22732 & ~n22733;
  assign n22735 = ~n22707 & n22734;
  assign n22736 = n22707 & ~n22734;
  assign n22737 = ~n22735 & ~n22736;
  assign n22738 = ~n22706 & n22737;
  assign n22739 = n22706 & ~n22737;
  assign n22740 = ~n22738 & ~n22739;
  assign n22741 = n22696 & ~n22740;
  assign n22742 = ~n22696 & n22740;
  assign n22743 = ~n22741 & ~n22742;
  assign n22744 = n4721 & n20419;
  assign n22745 = n4691 & n20422;
  assign n22746 = n4515 & n20425;
  assign n22747 = n4516 & n20786;
  assign n22748 = ~n22745 & ~n22746;
  assign n22749 = ~n22744 & n22748;
  assign n22750 = ~n22747 & n22749;
  assign n22751 = pi26  & n22750;
  assign n22752 = ~pi26  & ~n22750;
  assign n22753 = ~n22751 & ~n22752;
  assign n22754 = n22743 & ~n22753;
  assign n22755 = ~n22743 & n22753;
  assign n22756 = ~n22754 & ~n22755;
  assign n22757 = ~n22695 & n22756;
  assign n22758 = n22695 & ~n22756;
  assign n22759 = ~n22757 & ~n22758;
  assign n22760 = ~n22694 & n22759;
  assign n22761 = n22694 & ~n22759;
  assign n22762 = ~n22760 & ~n22761;
  assign n22763 = n22684 & ~n22762;
  assign n22764 = ~n22684 & n22762;
  assign n22765 = ~n22763 & ~n22764;
  assign n22766 = n5982 & n20401;
  assign n22767 = n5901 & n20404;
  assign n22768 = n5312 & n20407;
  assign n22769 = n5306 & n21286;
  assign n22770 = ~n22767 & ~n22768;
  assign n22771 = ~n22766 & n22770;
  assign n22772 = ~n22769 & n22771;
  assign n22773 = pi20  & n22772;
  assign n22774 = ~pi20  & ~n22772;
  assign n22775 = ~n22773 & ~n22774;
  assign n22776 = n22765 & ~n22775;
  assign n22777 = ~n22765 & n22775;
  assign n22778 = ~n22776 & ~n22777;
  assign n22779 = ~n22683 & n22778;
  assign n22780 = n22683 & ~n22778;
  assign n22781 = ~n22779 & ~n22780;
  assign n22782 = ~n22682 & n22781;
  assign n22783 = n22682 & ~n22781;
  assign n22784 = ~n22782 & ~n22783;
  assign n22785 = n22672 & ~n22784;
  assign n22786 = ~n22672 & n22784;
  assign n22787 = ~n22785 & ~n22786;
  assign n22788 = n7380 & n20383;
  assign n22789 = n7243 & n20386;
  assign n22790 = n6653 & n20389;
  assign n22791 = n6647 & n21737;
  assign n22792 = ~n22789 & ~n22790;
  assign n22793 = ~n22788 & n22792;
  assign n22794 = ~n22791 & n22793;
  assign n22795 = pi14  & n22794;
  assign n22796 = ~pi14  & ~n22794;
  assign n22797 = ~n22795 & ~n22796;
  assign n22798 = n22787 & ~n22797;
  assign n22799 = ~n22787 & n22797;
  assign n22800 = ~n22798 & ~n22799;
  assign n22801 = ~n22671 & n22800;
  assign n22802 = n22671 & ~n22800;
  assign n22803 = ~n22801 & ~n22802;
  assign n22804 = ~n22670 & n22803;
  assign n22805 = n22670 & ~n22803;
  assign n22806 = ~n22804 & ~n22805;
  assign n22807 = n22660 & ~n22806;
  assign n22808 = ~n22660 & n22806;
  assign n22809 = ~n22807 & ~n22808;
  assign n22810 = n9355 & n20365;
  assign n22811 = n8939 & n20368;
  assign n22812 = n8206 & n20371;
  assign n22813 = n20544 & ~n20546;
  assign n22814 = ~n20547 & ~n22813;
  assign n22815 = n8200 & n22814;
  assign n22816 = ~n22811 & ~n22812;
  assign n22817 = ~n22810 & n22816;
  assign n22818 = ~n22815 & n22817;
  assign n22819 = pi8  & n22818;
  assign n22820 = ~pi8  & ~n22818;
  assign n22821 = ~n22819 & ~n22820;
  assign n22822 = n22809 & ~n22821;
  assign n22823 = ~n22809 & n22821;
  assign n22824 = ~n22822 & ~n22823;
  assign n22825 = ~n22659 & n22824;
  assign n22826 = n22659 & ~n22824;
  assign n22827 = ~n22825 & ~n22826;
  assign n22828 = ~n20569 & n22827;
  assign n22829 = n71 & n20358;
  assign n22830 = n10329 & n20361;
  assign n22831 = n9836 & n20365;
  assign n22832 = n20552 & ~n20554;
  assign n22833 = ~n20555 & ~n22832;
  assign n22834 = n9830 & n22833;
  assign n22835 = ~n22830 & ~n22831;
  assign n22836 = ~n22829 & n22835;
  assign n22837 = ~n22834 & n22836;
  assign n22838 = ~pi5  & ~n22837;
  assign n22839 = pi5  & n22837;
  assign n22840 = ~n22838 & ~n22839;
  assign n22841 = n22655 & ~n22657;
  assign n22842 = ~n22658 & ~n22841;
  assign n22843 = ~n22840 & n22842;
  assign n22844 = n71 & n20361;
  assign n22845 = n10329 & n20365;
  assign n22846 = n9836 & n20368;
  assign n22847 = n20548 & ~n20550;
  assign n22848 = ~n20551 & ~n22847;
  assign n22849 = n9830 & n22848;
  assign n22850 = ~n22845 & ~n22846;
  assign n22851 = ~n22844 & n22850;
  assign n22852 = ~n22849 & n22851;
  assign n22853 = ~pi5  & ~n22852;
  assign n22854 = pi5  & n22852;
  assign n22855 = ~n22853 & ~n22854;
  assign n22856 = n22651 & ~n22653;
  assign n22857 = ~n22654 & ~n22856;
  assign n22858 = ~n22855 & n22857;
  assign n22859 = n22647 & ~n22649;
  assign n22860 = ~n22650 & ~n22859;
  assign n22861 = n71 & n20365;
  assign n22862 = n10329 & n20368;
  assign n22863 = n9836 & n20371;
  assign n22864 = n9830 & n22814;
  assign n22865 = ~n22862 & ~n22863;
  assign n22866 = ~n22861 & n22865;
  assign n22867 = ~n22864 & n22866;
  assign n22868 = pi5  & n22867;
  assign n22869 = ~pi5  & ~n22867;
  assign n22870 = ~n22868 & ~n22869;
  assign n22871 = n22860 & ~n22870;
  assign n22872 = n22643 & ~n22645;
  assign n22873 = ~n22646 & ~n22872;
  assign n22874 = n71 & n20368;
  assign n22875 = n10329 & n20371;
  assign n22876 = n9836 & n20374;
  assign n22877 = n9830 & n22235;
  assign n22878 = ~n22875 & ~n22876;
  assign n22879 = ~n22874 & n22878;
  assign n22880 = ~n22877 & n22879;
  assign n22881 = pi5  & n22880;
  assign n22882 = ~pi5  & ~n22880;
  assign n22883 = ~n22881 & ~n22882;
  assign n22884 = n22873 & ~n22883;
  assign n22885 = n71 & n20371;
  assign n22886 = n10329 & n20374;
  assign n22887 = n9836 & n20377;
  assign n22888 = n9830 & n22250;
  assign n22889 = ~n22886 & ~n22887;
  assign n22890 = ~n22885 & n22889;
  assign n22891 = ~n22888 & n22890;
  assign n22892 = ~pi5  & ~n22891;
  assign n22893 = pi5  & n22891;
  assign n22894 = ~n22892 & ~n22893;
  assign n22895 = n22639 & ~n22641;
  assign n22896 = ~n22642 & ~n22895;
  assign n22897 = ~n22894 & n22896;
  assign n22898 = n71 & n20374;
  assign n22899 = n10329 & n20377;
  assign n22900 = n9836 & n20380;
  assign n22901 = n9830 & n22263;
  assign n22902 = ~n22899 & ~n22900;
  assign n22903 = ~n22898 & n22902;
  assign n22904 = ~n22901 & n22903;
  assign n22905 = ~pi5  & ~n22904;
  assign n22906 = pi5  & n22904;
  assign n22907 = ~n22905 & ~n22906;
  assign n22908 = n22635 & ~n22637;
  assign n22909 = ~n22638 & ~n22908;
  assign n22910 = ~n22907 & n22909;
  assign n22911 = n71 & n20377;
  assign n22912 = n10329 & n20380;
  assign n22913 = n9836 & n20383;
  assign n22914 = n9830 & n22083;
  assign n22915 = ~n22912 & ~n22913;
  assign n22916 = ~n22911 & n22915;
  assign n22917 = ~n22914 & n22916;
  assign n22918 = ~pi5  & ~n22917;
  assign n22919 = pi5  & n22917;
  assign n22920 = ~n22918 & ~n22919;
  assign n22921 = n22631 & ~n22633;
  assign n22922 = ~n22634 & ~n22921;
  assign n22923 = ~n22920 & n22922;
  assign n22924 = n22627 & ~n22629;
  assign n22925 = ~n22630 & ~n22924;
  assign n22926 = n71 & n20380;
  assign n22927 = n10329 & n20383;
  assign n22928 = n9836 & n20386;
  assign n22929 = n9830 & n20574;
  assign n22930 = ~n22927 & ~n22928;
  assign n22931 = ~n22926 & n22930;
  assign n22932 = ~n22929 & n22931;
  assign n22933 = pi5  & n22932;
  assign n22934 = ~pi5  & ~n22932;
  assign n22935 = ~n22933 & ~n22934;
  assign n22936 = n22925 & ~n22935;
  assign n22937 = n22623 & ~n22625;
  assign n22938 = ~n22626 & ~n22937;
  assign n22939 = n71 & n20383;
  assign n22940 = n10329 & n20386;
  assign n22941 = n9836 & n20389;
  assign n22942 = n9830 & n21737;
  assign n22943 = ~n22940 & ~n22941;
  assign n22944 = ~n22939 & n22943;
  assign n22945 = ~n22942 & n22944;
  assign n22946 = pi5  & n22945;
  assign n22947 = ~pi5  & ~n22945;
  assign n22948 = ~n22946 & ~n22947;
  assign n22949 = n22938 & ~n22948;
  assign n22950 = n22619 & ~n22621;
  assign n22951 = ~n22622 & ~n22950;
  assign n22952 = n71 & n20386;
  assign n22953 = n10329 & n20389;
  assign n22954 = n9836 & n20392;
  assign n22955 = n9830 & n21752;
  assign n22956 = ~n22953 & ~n22954;
  assign n22957 = ~n22952 & n22956;
  assign n22958 = ~n22955 & n22957;
  assign n22959 = pi5  & n22958;
  assign n22960 = ~pi5  & ~n22958;
  assign n22961 = ~n22959 & ~n22960;
  assign n22962 = n22951 & ~n22961;
  assign n22963 = n71 & n20389;
  assign n22964 = n10329 & n20392;
  assign n22965 = n9836 & n20395;
  assign n22966 = n9830 & n21716;
  assign n22967 = ~n22964 & ~n22965;
  assign n22968 = ~n22963 & n22967;
  assign n22969 = ~n22966 & n22968;
  assign n22970 = ~pi5  & ~n22969;
  assign n22971 = pi5  & n22969;
  assign n22972 = ~n22970 & ~n22971;
  assign n22973 = n22615 & ~n22617;
  assign n22974 = ~n22618 & ~n22973;
  assign n22975 = ~n22972 & n22974;
  assign n22976 = n71 & n20392;
  assign n22977 = n10329 & n20395;
  assign n22978 = n9836 & n20398;
  assign n22979 = n9830 & n20586;
  assign n22980 = ~n22977 & ~n22978;
  assign n22981 = ~n22976 & n22980;
  assign n22982 = ~n22979 & n22981;
  assign n22983 = ~pi5  & ~n22982;
  assign n22984 = pi5  & n22982;
  assign n22985 = ~n22983 & ~n22984;
  assign n22986 = n22611 & ~n22613;
  assign n22987 = ~n22614 & ~n22986;
  assign n22988 = ~n22985 & n22987;
  assign n22989 = n71 & n20395;
  assign n22990 = n10329 & n20398;
  assign n22991 = n9836 & n20401;
  assign n22992 = n9830 & n21305;
  assign n22993 = ~n22990 & ~n22991;
  assign n22994 = ~n22989 & n22993;
  assign n22995 = ~n22992 & n22994;
  assign n22996 = ~pi5  & ~n22995;
  assign n22997 = pi5  & n22995;
  assign n22998 = ~n22996 & ~n22997;
  assign n22999 = n22607 & ~n22609;
  assign n23000 = ~n22610 & ~n22999;
  assign n23001 = ~n22998 & n23000;
  assign n23002 = n22603 & ~n22605;
  assign n23003 = ~n22606 & ~n23002;
  assign n23004 = n71 & n20398;
  assign n23005 = n10329 & n20401;
  assign n23006 = n9836 & n20404;
  assign n23007 = n9830 & n21322;
  assign n23008 = ~n23005 & ~n23006;
  assign n23009 = ~n23004 & n23008;
  assign n23010 = ~n23007 & n23009;
  assign n23011 = pi5  & n23010;
  assign n23012 = ~pi5  & ~n23010;
  assign n23013 = ~n23011 & ~n23012;
  assign n23014 = n23003 & ~n23013;
  assign n23015 = n22599 & ~n22601;
  assign n23016 = ~n22602 & ~n23015;
  assign n23017 = n71 & n20401;
  assign n23018 = n10329 & n20404;
  assign n23019 = n9836 & n20407;
  assign n23020 = n9830 & n21286;
  assign n23021 = ~n23018 & ~n23019;
  assign n23022 = ~n23017 & n23021;
  assign n23023 = ~n23020 & n23022;
  assign n23024 = pi5  & n23023;
  assign n23025 = ~pi5  & ~n23023;
  assign n23026 = ~n23024 & ~n23025;
  assign n23027 = n23016 & ~n23026;
  assign n23028 = n22595 & ~n22597;
  assign n23029 = ~n22598 & ~n23028;
  assign n23030 = n71 & n20404;
  assign n23031 = n10329 & n20407;
  assign n23032 = n9836 & n20410;
  assign n23033 = n9830 & n20991;
  assign n23034 = ~n23031 & ~n23032;
  assign n23035 = ~n23030 & n23034;
  assign n23036 = ~n23033 & n23035;
  assign n23037 = pi5  & n23036;
  assign n23038 = ~pi5  & ~n23036;
  assign n23039 = ~n23037 & ~n23038;
  assign n23040 = n23029 & ~n23039;
  assign n23041 = n71 & n20407;
  assign n23042 = n10329 & n20410;
  assign n23043 = n9836 & n20413;
  assign n23044 = n9830 & n21004;
  assign n23045 = ~n23042 & ~n23043;
  assign n23046 = ~n23041 & n23045;
  assign n23047 = ~n23044 & n23046;
  assign n23048 = ~pi5  & ~n23047;
  assign n23049 = pi5  & n23047;
  assign n23050 = ~n23048 & ~n23049;
  assign n23051 = n22591 & ~n22593;
  assign n23052 = ~n22594 & ~n23051;
  assign n23053 = ~n23050 & n23052;
  assign n23054 = n71 & n20410;
  assign n23055 = n10329 & n20413;
  assign n23056 = n9836 & n20416;
  assign n23057 = n9830 & n21019;
  assign n23058 = ~n23055 & ~n23056;
  assign n23059 = ~n23054 & n23058;
  assign n23060 = ~n23057 & n23059;
  assign n23061 = ~pi5  & ~n23060;
  assign n23062 = pi5  & n23060;
  assign n23063 = ~n23061 & ~n23062;
  assign n23064 = n22587 & ~n22589;
  assign n23065 = ~n22590 & ~n23064;
  assign n23066 = ~n23063 & n23065;
  assign n23067 = n71 & n20413;
  assign n23068 = n10329 & n20416;
  assign n23069 = n9836 & n20419;
  assign n23070 = n9830 & n20928;
  assign n23071 = ~n23068 & ~n23069;
  assign n23072 = ~n23067 & n23071;
  assign n23073 = ~n23070 & n23072;
  assign n23074 = ~pi5  & ~n23073;
  assign n23075 = pi5  & n23073;
  assign n23076 = ~n23074 & ~n23075;
  assign n23077 = n22583 & ~n22585;
  assign n23078 = ~n22586 & ~n23077;
  assign n23079 = ~n23076 & n23078;
  assign n23080 = n22579 & ~n22581;
  assign n23081 = ~n22582 & ~n23080;
  assign n23082 = n71 & n20416;
  assign n23083 = n10329 & n20419;
  assign n23084 = n9836 & n20422;
  assign n23085 = n9830 & n20771;
  assign n23086 = ~n23083 & ~n23084;
  assign n23087 = ~n23082 & n23086;
  assign n23088 = ~n23085 & n23087;
  assign n23089 = pi5  & n23088;
  assign n23090 = ~pi5  & ~n23088;
  assign n23091 = ~n23089 & ~n23090;
  assign n23092 = n23081 & ~n23091;
  assign n23093 = n22575 & ~n22577;
  assign n23094 = ~n22578 & ~n23093;
  assign n23095 = n71 & n20419;
  assign n23096 = n10329 & n20422;
  assign n23097 = n9836 & n20425;
  assign n23098 = n9830 & n20786;
  assign n23099 = ~n23096 & ~n23097;
  assign n23100 = ~n23095 & n23099;
  assign n23101 = ~n23098 & n23100;
  assign n23102 = pi5  & n23101;
  assign n23103 = ~pi5  & ~n23101;
  assign n23104 = ~n23102 & ~n23103;
  assign n23105 = n23094 & ~n23104;
  assign n23106 = n22571 & ~n22573;
  assign n23107 = ~n22574 & ~n23106;
  assign n23108 = n71 & n20422;
  assign n23109 = n10329 & n20425;
  assign n23110 = n9836 & n20428;
  assign n23111 = n9830 & n20801;
  assign n23112 = ~n23109 & ~n23110;
  assign n23113 = ~n23108 & n23112;
  assign n23114 = ~n23111 & n23113;
  assign n23115 = pi5  & n23114;
  assign n23116 = ~pi5  & ~n23114;
  assign n23117 = ~n23115 & ~n23116;
  assign n23118 = n23107 & ~n23117;
  assign n23119 = n71 & n20425;
  assign n23120 = n10329 & n20428;
  assign n23121 = n9836 & n20431;
  assign n23122 = n9830 & n20727;
  assign n23123 = ~n23120 & ~n23121;
  assign n23124 = ~n23119 & n23123;
  assign n23125 = ~n23122 & n23124;
  assign n23126 = ~pi5  & ~n23125;
  assign n23127 = pi5  & n23125;
  assign n23128 = ~n23126 & ~n23127;
  assign n23129 = n22567 & ~n22569;
  assign n23130 = ~n22570 & ~n23129;
  assign n23131 = ~n23128 & n23130;
  assign n23132 = n71 & n20428;
  assign n23133 = n10329 & n20431;
  assign n23134 = n9836 & n20434;
  assign n23135 = n9830 & n20598;
  assign n23136 = ~n23133 & ~n23134;
  assign n23137 = ~n23132 & n23136;
  assign n23138 = ~n23135 & n23137;
  assign n23139 = pi5  & n23138;
  assign n23140 = ~pi5  & ~n23138;
  assign n23141 = ~n23139 & ~n23140;
  assign n23142 = n22563 & ~n22565;
  assign n23143 = ~n22566 & ~n23142;
  assign n23144 = ~n23141 & n23143;
  assign n23145 = n71 & n20431;
  assign n23146 = n10329 & n20434;
  assign n23147 = n9836 & n20437;
  assign n23148 = n9830 & n20651;
  assign n23149 = ~n23146 & ~n23147;
  assign n23150 = ~n23145 & n23149;
  assign n23151 = ~n23148 & n23150;
  assign n23152 = ~pi5  & ~n23151;
  assign n23153 = pi5  & n23151;
  assign n23154 = ~n23152 & ~n23153;
  assign n23155 = pi8  & ~n22543;
  assign n23156 = n22550 & ~n23155;
  assign n23157 = ~n22550 & n23155;
  assign n23158 = ~n23156 & ~n23157;
  assign n23159 = ~n23154 & n23158;
  assign n23160 = n71 & n20434;
  assign n23161 = n10329 & n20437;
  assign n23162 = n9836 & n20440;
  assign n23163 = n9830 & n20668;
  assign n23164 = ~n23161 & ~n23162;
  assign n23165 = ~n23160 & n23164;
  assign n23166 = ~n23163 & n23165;
  assign n23167 = pi5  & n23166;
  assign n23168 = ~pi5  & ~n23166;
  assign n23169 = ~n23167 & ~n23168;
  assign n23170 = n22537 & ~n22542;
  assign n23171 = ~n22543 & ~n23170;
  assign n23172 = ~n23169 & n23171;
  assign n23173 = n67 & n20447;
  assign n23174 = pi5  & n23173;
  assign n23175 = n71 & n20445;
  assign n23176 = n10329 & n20447;
  assign n23177 = n9830 & ~n20624;
  assign n23178 = ~n23175 & ~n23176;
  assign n23179 = ~n23177 & n23178;
  assign n23180 = ~n23174 & n23179;
  assign n23181 = n71 & n20440;
  assign n23182 = n10329 & n20445;
  assign n23183 = n9836 & n20447;
  assign n23184 = n9830 & ~n20633;
  assign n23185 = ~n23182 & ~n23183;
  assign n23186 = ~n23181 & n23185;
  assign n23187 = ~n23184 & n23186;
  assign n23188 = pi5  & n23180;
  assign n23189 = n23187 & n23188;
  assign n23190 = n22536 & n23189;
  assign n23191 = n71 & n20437;
  assign n23192 = n10329 & n20440;
  assign n23193 = n9836 & n20445;
  assign n23194 = n9830 & n20610;
  assign n23195 = ~n23192 & ~n23193;
  assign n23196 = ~n23191 & n23195;
  assign n23197 = ~n23194 & n23196;
  assign n23198 = pi5  & n23197;
  assign n23199 = ~pi5  & ~n23197;
  assign n23200 = ~n23198 & ~n23199;
  assign n23201 = ~n22536 & ~n23189;
  assign n23202 = ~n23190 & ~n23201;
  assign n23203 = ~n23200 & n23202;
  assign n23204 = ~n23190 & ~n23203;
  assign n23205 = n23169 & ~n23171;
  assign n23206 = ~n23172 & ~n23205;
  assign n23207 = ~n23204 & n23206;
  assign n23208 = ~n23172 & ~n23207;
  assign n23209 = n23154 & ~n23158;
  assign n23210 = ~n23159 & ~n23209;
  assign n23211 = ~n23208 & n23210;
  assign n23212 = ~n23159 & ~n23211;
  assign n23213 = n23141 & ~n23143;
  assign n23214 = ~n23144 & ~n23213;
  assign n23215 = ~n23212 & n23214;
  assign n23216 = ~n23144 & ~n23215;
  assign n23217 = n23128 & ~n23130;
  assign n23218 = ~n23131 & ~n23217;
  assign n23219 = ~n23216 & n23218;
  assign n23220 = ~n23131 & ~n23219;
  assign n23221 = ~n23107 & n23117;
  assign n23222 = ~n23118 & ~n23221;
  assign n23223 = ~n23220 & n23222;
  assign n23224 = ~n23118 & ~n23223;
  assign n23225 = ~n23094 & n23104;
  assign n23226 = ~n23105 & ~n23225;
  assign n23227 = ~n23224 & n23226;
  assign n23228 = ~n23105 & ~n23227;
  assign n23229 = ~n23081 & n23091;
  assign n23230 = ~n23092 & ~n23229;
  assign n23231 = ~n23228 & n23230;
  assign n23232 = ~n23092 & ~n23231;
  assign n23233 = n23076 & ~n23078;
  assign n23234 = ~n23079 & ~n23233;
  assign n23235 = ~n23232 & n23234;
  assign n23236 = ~n23079 & ~n23235;
  assign n23237 = n23063 & ~n23065;
  assign n23238 = ~n23066 & ~n23237;
  assign n23239 = ~n23236 & n23238;
  assign n23240 = ~n23066 & ~n23239;
  assign n23241 = n23050 & ~n23052;
  assign n23242 = ~n23053 & ~n23241;
  assign n23243 = ~n23240 & n23242;
  assign n23244 = ~n23053 & ~n23243;
  assign n23245 = ~n23029 & n23039;
  assign n23246 = ~n23040 & ~n23245;
  assign n23247 = ~n23244 & n23246;
  assign n23248 = ~n23040 & ~n23247;
  assign n23249 = ~n23016 & n23026;
  assign n23250 = ~n23027 & ~n23249;
  assign n23251 = ~n23248 & n23250;
  assign n23252 = ~n23027 & ~n23251;
  assign n23253 = ~n23003 & n23013;
  assign n23254 = ~n23014 & ~n23253;
  assign n23255 = ~n23252 & n23254;
  assign n23256 = ~n23014 & ~n23255;
  assign n23257 = n22998 & ~n23000;
  assign n23258 = ~n23001 & ~n23257;
  assign n23259 = ~n23256 & n23258;
  assign n23260 = ~n23001 & ~n23259;
  assign n23261 = n22985 & ~n22987;
  assign n23262 = ~n22988 & ~n23261;
  assign n23263 = ~n23260 & n23262;
  assign n23264 = ~n22988 & ~n23263;
  assign n23265 = n22972 & ~n22974;
  assign n23266 = ~n22975 & ~n23265;
  assign n23267 = ~n23264 & n23266;
  assign n23268 = ~n22975 & ~n23267;
  assign n23269 = ~n22951 & n22961;
  assign n23270 = ~n22962 & ~n23269;
  assign n23271 = ~n23268 & n23270;
  assign n23272 = ~n22962 & ~n23271;
  assign n23273 = ~n22938 & n22948;
  assign n23274 = ~n22949 & ~n23273;
  assign n23275 = ~n23272 & n23274;
  assign n23276 = ~n22949 & ~n23275;
  assign n23277 = ~n22925 & n22935;
  assign n23278 = ~n22936 & ~n23277;
  assign n23279 = ~n23276 & n23278;
  assign n23280 = ~n22936 & ~n23279;
  assign n23281 = n22920 & ~n22922;
  assign n23282 = ~n22923 & ~n23281;
  assign n23283 = ~n23280 & n23282;
  assign n23284 = ~n22923 & ~n23283;
  assign n23285 = n22907 & ~n22909;
  assign n23286 = ~n22910 & ~n23285;
  assign n23287 = ~n23284 & n23286;
  assign n23288 = ~n22910 & ~n23287;
  assign n23289 = n22894 & ~n22896;
  assign n23290 = ~n22897 & ~n23289;
  assign n23291 = ~n23288 & n23290;
  assign n23292 = ~n22897 & ~n23291;
  assign n23293 = ~n22873 & n22883;
  assign n23294 = ~n22884 & ~n23293;
  assign n23295 = ~n23292 & n23294;
  assign n23296 = ~n22884 & ~n23295;
  assign n23297 = ~n22860 & n22870;
  assign n23298 = ~n22871 & ~n23297;
  assign n23299 = ~n23296 & n23298;
  assign n23300 = ~n22871 & ~n23299;
  assign n23301 = n22855 & ~n22857;
  assign n23302 = ~n22858 & ~n23301;
  assign n23303 = ~n23300 & n23302;
  assign n23304 = ~n22858 & ~n23303;
  assign n23305 = n22840 & ~n22842;
  assign n23306 = ~n22843 & ~n23305;
  assign n23307 = ~n23304 & n23306;
  assign n23308 = ~n22843 & ~n23307;
  assign n23309 = n20569 & ~n22827;
  assign n23310 = ~n22828 & ~n23309;
  assign n23311 = ~n23308 & n23310;
  assign n23312 = ~n22828 & ~n23311;
  assign n23313 = ~n13020 & ~n20353;
  assign n23314 = ~n12872 & ~n12950;
  assign n23315 = ~n12926 & ~n12929;
  assign n23316 = ~n12911 & ~n12914;
  assign n23317 = ~n77 & n12426;
  assign n23318 = ~n12163 & ~n23317;
  assign n23319 = pi23  & ~n23318;
  assign n23320 = ~pi23  & n23318;
  assign n23321 = ~n23319 & ~n23320;
  assign n23322 = ~n315 & ~n335;
  assign n23323 = ~n577 & ~n666;
  assign n23324 = n23322 & n23323;
  assign n23325 = n166 & n1086;
  assign n23326 = n1157 & n1710;
  assign n23327 = n4274 & n6976;
  assign n23328 = n23326 & n23327;
  assign n23329 = n23324 & n23325;
  assign n23330 = n6880 & n23329;
  assign n23331 = n852 & n23328;
  assign n23332 = n23330 & n23331;
  assign n23333 = n5367 & n23332;
  assign n23334 = n13450 & n14850;
  assign n23335 = n23333 & n23334;
  assign n23336 = n12731 & n23335;
  assign n23337 = n12910 & n23336;
  assign n23338 = ~n12910 & ~n23336;
  assign n23339 = ~n23337 & ~n23338;
  assign n23340 = n23321 & n23339;
  assign n23341 = ~n23321 & ~n23339;
  assign n23342 = ~n23340 & ~n23341;
  assign n23343 = ~n23316 & n23342;
  assign n23344 = n23316 & ~n23342;
  assign n23345 = ~n23343 & ~n23344;
  assign n23346 = n3896 & n12184;
  assign n23347 = n3683 & n12187;
  assign n23348 = n564 & n12190;
  assign n23349 = n566 & n12845;
  assign n23350 = ~n23347 & ~n23348;
  assign n23351 = ~n23346 & n23350;
  assign n23352 = ~n23349 & n23351;
  assign n23353 = n23345 & ~n23352;
  assign n23354 = ~n23345 & n23352;
  assign n23355 = ~n23353 & ~n23354;
  assign n23356 = n23315 & ~n23355;
  assign n23357 = ~n23315 & n23355;
  assign n23358 = ~n23356 & ~n23357;
  assign n23359 = n4472 & n12175;
  assign n23360 = n4070 & n12178;
  assign n23361 = n3943 & n12181;
  assign n23362 = n3944 & n12961;
  assign n23363 = ~n23360 & ~n23361;
  assign n23364 = ~n23359 & n23363;
  assign n23365 = ~n23362 & n23364;
  assign n23366 = pi29  & n23365;
  assign n23367 = ~pi29  & ~n23365;
  assign n23368 = ~n23366 & ~n23367;
  assign n23369 = n23358 & ~n23368;
  assign n23370 = ~n23358 & n23368;
  assign n23371 = ~n23369 & ~n23370;
  assign n23372 = ~n12932 & ~n12947;
  assign n23373 = n4721 & n12166;
  assign n23374 = n4691 & n12172;
  assign n23375 = n4515 & n12168;
  assign n23376 = n4516 & n13106;
  assign n23377 = ~n23373 & ~n23375;
  assign n23378 = ~n23374 & n23377;
  assign n23379 = ~n23376 & n23378;
  assign n23380 = pi26  & n23379;
  assign n23381 = ~pi26  & ~n23379;
  assign n23382 = ~n23380 & ~n23381;
  assign n23383 = ~n23372 & ~n23382;
  assign n23384 = n23372 & n23382;
  assign n23385 = ~n23383 & ~n23384;
  assign n23386 = n23371 & n23385;
  assign n23387 = ~n23371 & ~n23385;
  assign n23388 = ~n23386 & ~n23387;
  assign n23389 = ~n23314 & n23388;
  assign n23390 = n23314 & ~n23388;
  assign n23391 = ~n23389 & ~n23390;
  assign n23392 = ~n23313 & n23391;
  assign n23393 = n23313 & ~n23391;
  assign n23394 = ~n23392 & ~n23393;
  assign n23395 = n71 & n23394;
  assign n23396 = n10329 & n20355;
  assign n23397 = n9836 & n20358;
  assign n23398 = ~n20557 & ~n20560;
  assign n23399 = n20355 & n23394;
  assign n23400 = ~n20355 & ~n23394;
  assign n23401 = ~n23399 & ~n23400;
  assign n23402 = ~n23398 & n23401;
  assign n23403 = n23398 & ~n23401;
  assign n23404 = ~n23402 & ~n23403;
  assign n23405 = n9830 & n23404;
  assign n23406 = ~n23396 & ~n23397;
  assign n23407 = ~n23395 & n23406;
  assign n23408 = ~n23405 & n23407;
  assign n23409 = ~pi5  & ~n23408;
  assign n23410 = pi5  & n23408;
  assign n23411 = ~n23409 & ~n23410;
  assign n23412 = ~n22822 & ~n22825;
  assign n23413 = ~n22804 & ~n22808;
  assign n23414 = n8161 & n20371;
  assign n23415 = n7847 & n20374;
  assign n23416 = n7554 & n20377;
  assign n23417 = n7548 & n22250;
  assign n23418 = ~n23415 & ~n23416;
  assign n23419 = ~n23414 & n23418;
  assign n23420 = ~n23417 & n23419;
  assign n23421 = ~pi11  & ~n23420;
  assign n23422 = pi11  & n23420;
  assign n23423 = ~n23421 & ~n23422;
  assign n23424 = ~n22798 & ~n22801;
  assign n23425 = ~n22782 & ~n22786;
  assign n23426 = n6608 & n20389;
  assign n23427 = n6356 & n20392;
  assign n23428 = n6140 & n20395;
  assign n23429 = n6134 & n21716;
  assign n23430 = ~n23427 & ~n23428;
  assign n23431 = ~n23426 & n23430;
  assign n23432 = ~n23429 & n23431;
  assign n23433 = ~pi17  & ~n23432;
  assign n23434 = pi17  & n23432;
  assign n23435 = ~n23433 & ~n23434;
  assign n23436 = ~n22776 & ~n22779;
  assign n23437 = ~n22760 & ~n22764;
  assign n23438 = n5267 & n20407;
  assign n23439 = n5185 & n20410;
  assign n23440 = n5121 & n20413;
  assign n23441 = n78 & n21004;
  assign n23442 = ~n23439 & ~n23440;
  assign n23443 = ~n23438 & n23442;
  assign n23444 = ~n23441 & n23443;
  assign n23445 = ~pi23  & ~n23444;
  assign n23446 = pi23  & n23444;
  assign n23447 = ~n23445 & ~n23446;
  assign n23448 = ~n22754 & ~n22757;
  assign n23449 = ~n22738 & ~n22742;
  assign n23450 = n4472 & n20425;
  assign n23451 = n4070 & n20428;
  assign n23452 = n3943 & n20431;
  assign n23453 = n3944 & n20727;
  assign n23454 = ~n23451 & ~n23452;
  assign n23455 = ~n23450 & n23454;
  assign n23456 = ~n23453 & n23455;
  assign n23457 = ~pi29  & ~n23456;
  assign n23458 = pi29  & n23456;
  assign n23459 = ~n23457 & ~n23458;
  assign n23460 = ~n22732 & ~n22735;
  assign n23461 = ~n213 & ~n447;
  assign n23462 = ~n544 & ~n585;
  assign n23463 = ~n588 & n23462;
  assign n23464 = n765 & n23461;
  assign n23465 = n1595 & n2360;
  assign n23466 = n4911 & n23465;
  assign n23467 = n23463 & n23464;
  assign n23468 = n1053 & n6189;
  assign n23469 = n23467 & n23468;
  assign n23470 = n12456 & n23466;
  assign n23471 = n23469 & n23470;
  assign n23472 = n12443 & n23471;
  assign n23473 = n12897 & n23472;
  assign n23474 = n14710 & n23473;
  assign n23475 = n3896 & n20434;
  assign n23476 = n564 & n20440;
  assign n23477 = n3683 & n20437;
  assign n23478 = n566 & n20668;
  assign n23479 = ~n23476 & ~n23477;
  assign n23480 = ~n23475 & n23479;
  assign n23481 = ~n23478 & n23480;
  assign n23482 = ~n23474 & ~n23481;
  assign n23483 = n23474 & n23481;
  assign n23484 = ~n23482 & ~n23483;
  assign n23485 = ~n23460 & n23484;
  assign n23486 = n23460 & ~n23484;
  assign n23487 = ~n23485 & ~n23486;
  assign n23488 = ~n23459 & n23487;
  assign n23489 = n23459 & ~n23487;
  assign n23490 = ~n23488 & ~n23489;
  assign n23491 = n23449 & ~n23490;
  assign n23492 = ~n23449 & n23490;
  assign n23493 = ~n23491 & ~n23492;
  assign n23494 = n4721 & n20416;
  assign n23495 = n4691 & n20419;
  assign n23496 = n4515 & n20422;
  assign n23497 = n4516 & n20771;
  assign n23498 = ~n23495 & ~n23496;
  assign n23499 = ~n23494 & n23498;
  assign n23500 = ~n23497 & n23499;
  assign n23501 = pi26  & n23500;
  assign n23502 = ~pi26  & ~n23500;
  assign n23503 = ~n23501 & ~n23502;
  assign n23504 = n23493 & ~n23503;
  assign n23505 = ~n23493 & n23503;
  assign n23506 = ~n23504 & ~n23505;
  assign n23507 = ~n23448 & n23506;
  assign n23508 = n23448 & ~n23506;
  assign n23509 = ~n23507 & ~n23508;
  assign n23510 = ~n23447 & n23509;
  assign n23511 = n23447 & ~n23509;
  assign n23512 = ~n23510 & ~n23511;
  assign n23513 = n23437 & ~n23512;
  assign n23514 = ~n23437 & n23512;
  assign n23515 = ~n23513 & ~n23514;
  assign n23516 = n5982 & n20398;
  assign n23517 = n5901 & n20401;
  assign n23518 = n5312 & n20404;
  assign n23519 = n5306 & n21322;
  assign n23520 = ~n23517 & ~n23518;
  assign n23521 = ~n23516 & n23520;
  assign n23522 = ~n23519 & n23521;
  assign n23523 = pi20  & n23522;
  assign n23524 = ~pi20  & ~n23522;
  assign n23525 = ~n23523 & ~n23524;
  assign n23526 = n23515 & ~n23525;
  assign n23527 = ~n23515 & n23525;
  assign n23528 = ~n23526 & ~n23527;
  assign n23529 = ~n23436 & n23528;
  assign n23530 = n23436 & ~n23528;
  assign n23531 = ~n23529 & ~n23530;
  assign n23532 = ~n23435 & n23531;
  assign n23533 = n23435 & ~n23531;
  assign n23534 = ~n23532 & ~n23533;
  assign n23535 = n23425 & ~n23534;
  assign n23536 = ~n23425 & n23534;
  assign n23537 = ~n23535 & ~n23536;
  assign n23538 = n7380 & n20380;
  assign n23539 = n7243 & n20383;
  assign n23540 = n6653 & n20386;
  assign n23541 = n6647 & n20574;
  assign n23542 = ~n23539 & ~n23540;
  assign n23543 = ~n23538 & n23542;
  assign n23544 = ~n23541 & n23543;
  assign n23545 = pi14  & n23544;
  assign n23546 = ~pi14  & ~n23544;
  assign n23547 = ~n23545 & ~n23546;
  assign n23548 = n23537 & ~n23547;
  assign n23549 = ~n23537 & n23547;
  assign n23550 = ~n23548 & ~n23549;
  assign n23551 = ~n23424 & n23550;
  assign n23552 = n23424 & ~n23550;
  assign n23553 = ~n23551 & ~n23552;
  assign n23554 = ~n23423 & n23553;
  assign n23555 = n23423 & ~n23553;
  assign n23556 = ~n23554 & ~n23555;
  assign n23557 = n23413 & ~n23556;
  assign n23558 = ~n23413 & n23556;
  assign n23559 = ~n23557 & ~n23558;
  assign n23560 = n9355 & n20361;
  assign n23561 = n8939 & n20365;
  assign n23562 = n8206 & n20368;
  assign n23563 = n8200 & n22848;
  assign n23564 = ~n23561 & ~n23562;
  assign n23565 = ~n23560 & n23564;
  assign n23566 = ~n23563 & n23565;
  assign n23567 = pi8  & n23566;
  assign n23568 = ~pi8  & ~n23566;
  assign n23569 = ~n23567 & ~n23568;
  assign n23570 = n23559 & ~n23569;
  assign n23571 = ~n23559 & n23569;
  assign n23572 = ~n23570 & ~n23571;
  assign n23573 = ~n23412 & n23572;
  assign n23574 = n23412 & ~n23572;
  assign n23575 = ~n23573 & ~n23574;
  assign n23576 = ~n23411 & n23575;
  assign n23577 = n23411 & ~n23575;
  assign n23578 = ~n23576 & ~n23577;
  assign n23579 = n23312 & ~n23578;
  assign n23580 = ~n23312 & n23578;
  assign n23581 = ~n23579 & ~n23580;
  assign n23582 = ~n23357 & ~n23369;
  assign n23583 = ~n23343 & ~n23353;
  assign n23584 = ~n23338 & ~n23340;
  assign n23585 = ~n222 & ~n536;
  assign n23586 = n719 & n23585;
  assign n23587 = n737 & n743;
  assign n23588 = n1710 & n23587;
  assign n23589 = n7069 & n23586;
  assign n23590 = n23588 & n23589;
  assign n23591 = ~n122 & ~n509;
  assign n23592 = ~n641 & n23591;
  assign n23593 = n386 & n1118;
  assign n23594 = n1124 & n2903;
  assign n23595 = n23593 & n23594;
  assign n23596 = n23592 & n23595;
  assign n23597 = n810 & n23596;
  assign n23598 = n23590 & n23597;
  assign n23599 = n264 & n23598;
  assign n23600 = n986 & n23599;
  assign n23601 = ~n23584 & n23600;
  assign n23602 = n23584 & ~n23600;
  assign n23603 = ~n23601 & ~n23602;
  assign n23604 = n3896 & n12181;
  assign n23605 = n564 & n12187;
  assign n23606 = n3683 & n12184;
  assign n23607 = n566 & n12608;
  assign n23608 = ~n23605 & ~n23606;
  assign n23609 = ~n23604 & n23608;
  assign n23610 = ~n23607 & n23609;
  assign n23611 = n23603 & ~n23610;
  assign n23612 = ~n23603 & n23610;
  assign n23613 = ~n23611 & ~n23612;
  assign n23614 = ~n23583 & n23613;
  assign n23615 = n23583 & ~n23613;
  assign n23616 = ~n23614 & ~n23615;
  assign n23617 = n4472 & n12168;
  assign n23618 = n4070 & n12175;
  assign n23619 = n3943 & n12178;
  assign n23620 = n3944 & n12862;
  assign n23621 = ~n23618 & ~n23619;
  assign n23622 = ~n23617 & n23621;
  assign n23623 = ~n23620 & n23622;
  assign n23624 = pi29  & n23623;
  assign n23625 = ~pi29  & ~n23623;
  assign n23626 = ~n23624 & ~n23625;
  assign n23627 = n23616 & ~n23626;
  assign n23628 = ~n23616 & n23626;
  assign n23629 = ~n23627 & ~n23628;
  assign n23630 = ~n23582 & n23629;
  assign n23631 = n23582 & ~n23629;
  assign n23632 = ~n23630 & ~n23631;
  assign n23633 = n4691 & ~n12165;
  assign n23634 = ~n4721 & ~n23633;
  assign n23635 = ~n12163 & ~n23634;
  assign n23636 = n4516 & n13007;
  assign n23637 = n4515 & n12172;
  assign n23638 = ~n23636 & ~n23637;
  assign n23639 = ~n23635 & n23638;
  assign n23640 = pi26  & n23639;
  assign n23641 = ~pi26  & ~n23639;
  assign n23642 = ~n23640 & ~n23641;
  assign n23643 = n23632 & ~n23642;
  assign n23644 = ~n23630 & ~n23643;
  assign n23645 = ~n23601 & ~n23611;
  assign n23646 = ~n494 & ~n509;
  assign n23647 = n211 & n23646;
  assign n23648 = n782 & n14817;
  assign n23649 = n23647 & n23648;
  assign n23650 = n1471 & n1834;
  assign n23651 = n23649 & n23650;
  assign n23652 = n764 & n23651;
  assign n23653 = n724 & n23652;
  assign n23654 = n264 & n23653;
  assign n23655 = n839 & n23654;
  assign n23656 = n881 & n23655;
  assign n23657 = ~n23600 & n23656;
  assign n23658 = n23600 & ~n23656;
  assign n23659 = ~n23657 & ~n23658;
  assign n23660 = n3896 & n12178;
  assign n23661 = n3683 & n12181;
  assign n23662 = n564 & n12184;
  assign n23663 = n566 & n12880;
  assign n23664 = ~n23661 & ~n23662;
  assign n23665 = ~n23660 & n23664;
  assign n23666 = ~n23663 & n23665;
  assign n23667 = n23659 & ~n23666;
  assign n23668 = ~n23659 & n23666;
  assign n23669 = ~n23667 & ~n23668;
  assign n23670 = n23645 & ~n23669;
  assign n23671 = ~n23645 & n23669;
  assign n23672 = ~n23670 & ~n23671;
  assign n23673 = ~n23614 & ~n23627;
  assign n23674 = ~n23672 & n23673;
  assign n23675 = n23672 & ~n23673;
  assign n23676 = ~n23674 & ~n23675;
  assign n23677 = n4472 & n12172;
  assign n23678 = n4070 & n12168;
  assign n23679 = n3943 & n12175;
  assign n23680 = n3944 & n12939;
  assign n23681 = ~n23678 & ~n23679;
  assign n23682 = ~n23677 & n23681;
  assign n23683 = ~n23680 & n23682;
  assign n23684 = pi29  & n23683;
  assign n23685 = ~pi29  & ~n23683;
  assign n23686 = ~n23684 & ~n23685;
  assign n23687 = n12165 & ~n23638;
  assign n23688 = n4509 & n4514;
  assign n23689 = ~n12163 & ~n23688;
  assign n23690 = pi26  & ~n23689;
  assign n23691 = ~pi26  & n23689;
  assign n23692 = ~n23690 & ~n23691;
  assign n23693 = ~n23687 & ~n23692;
  assign n23694 = pi26  & n23687;
  assign n23695 = ~n23693 & ~n23694;
  assign n23696 = ~n23686 & ~n23695;
  assign n23697 = n23686 & n23695;
  assign n23698 = ~n23696 & ~n23697;
  assign n23699 = ~n23676 & ~n23698;
  assign n23700 = n23676 & n23698;
  assign n23701 = ~n23699 & ~n23700;
  assign n23702 = ~n23644 & n23701;
  assign n23703 = ~n23383 & ~n23386;
  assign n23704 = ~n23632 & n23642;
  assign n23705 = ~n23643 & ~n23704;
  assign n23706 = ~n23703 & n23705;
  assign n23707 = ~n23389 & ~n23392;
  assign n23708 = n23703 & ~n23705;
  assign n23709 = ~n23706 & ~n23708;
  assign n23710 = ~n23707 & n23709;
  assign n23711 = ~n23706 & ~n23710;
  assign n23712 = n23644 & ~n23701;
  assign n23713 = ~n23702 & ~n23712;
  assign n23714 = ~n23711 & n23713;
  assign n23715 = ~n23702 & ~n23714;
  assign n23716 = ~n23671 & ~n23675;
  assign n23717 = ~n23658 & ~n23667;
  assign n23718 = n519 & n617;
  assign n23719 = ~n494 & ~n568;
  assign n23720 = n732 & n23719;
  assign n23721 = n638 & n23720;
  assign n23722 = n373 & n23721;
  assign n23723 = n23718 & n23722;
  assign n23724 = n23600 & n23723;
  assign n23725 = ~n23600 & ~n23723;
  assign n23726 = ~n23724 & ~n23725;
  assign n23727 = n23692 & n23726;
  assign n23728 = ~n23692 & ~n23726;
  assign n23729 = ~n23727 & ~n23728;
  assign n23730 = ~n23717 & n23729;
  assign n23731 = n23717 & ~n23729;
  assign n23732 = ~n23730 & ~n23731;
  assign n23733 = n3896 & n12175;
  assign n23734 = n3683 & n12178;
  assign n23735 = n564 & n12181;
  assign n23736 = n566 & n12961;
  assign n23737 = ~n23734 & ~n23735;
  assign n23738 = ~n23733 & n23737;
  assign n23739 = ~n23736 & n23738;
  assign n23740 = n23732 & ~n23739;
  assign n23741 = ~n23732 & n23739;
  assign n23742 = ~n23740 & ~n23741;
  assign n23743 = n4472 & n12166;
  assign n23744 = n4070 & n12172;
  assign n23745 = n3943 & n12168;
  assign n23746 = n3944 & n13106;
  assign n23747 = ~n23743 & ~n23745;
  assign n23748 = ~n23744 & n23747;
  assign n23749 = ~n23746 & n23748;
  assign n23750 = pi29  & n23749;
  assign n23751 = ~pi29  & ~n23749;
  assign n23752 = ~n23750 & ~n23751;
  assign n23753 = n23742 & ~n23752;
  assign n23754 = ~n23742 & n23752;
  assign n23755 = ~n23753 & ~n23754;
  assign n23756 = n23716 & ~n23755;
  assign n23757 = ~n23716 & n23755;
  assign n23758 = ~n23756 & ~n23757;
  assign n23759 = ~n23696 & ~n23700;
  assign n23760 = n23758 & ~n23759;
  assign n23761 = ~n23758 & n23759;
  assign n23762 = ~n23760 & ~n23761;
  assign n23763 = n23715 & ~n23762;
  assign n23764 = ~n23715 & n23762;
  assign n23765 = ~n23763 & ~n23764;
  assign n23766 = n11476 & n23765;
  assign n23767 = n23711 & ~n23713;
  assign n23768 = ~n23714 & ~n23767;
  assign n23769 = n11463 & n23768;
  assign n23770 = n23707 & ~n23709;
  assign n23771 = ~n23710 & ~n23770;
  assign n23772 = n10883 & n23771;
  assign n23773 = n23768 & n23771;
  assign n23774 = n23394 & n23771;
  assign n23775 = ~n23399 & ~n23402;
  assign n23776 = ~n23394 & ~n23771;
  assign n23777 = ~n23774 & ~n23776;
  assign n23778 = ~n23775 & n23777;
  assign n23779 = ~n23774 & ~n23778;
  assign n23780 = ~n23768 & ~n23771;
  assign n23781 = ~n23773 & ~n23780;
  assign n23782 = ~n23779 & n23781;
  assign n23783 = ~n23773 & ~n23782;
  assign n23784 = n23765 & n23768;
  assign n23785 = ~n23765 & ~n23768;
  assign n23786 = ~n23784 & ~n23785;
  assign n23787 = ~n23783 & n23786;
  assign n23788 = n23783 & ~n23786;
  assign n23789 = ~n23787 & ~n23788;
  assign n23790 = n10884 & n23789;
  assign n23791 = ~n23769 & ~n23772;
  assign n23792 = ~n23766 & n23791;
  assign n23793 = ~n23790 & n23792;
  assign n23794 = pi2  & n23793;
  assign n23795 = ~pi2  & ~n23793;
  assign n23796 = ~n23794 & ~n23795;
  assign n23797 = n23581 & ~n23796;
  assign n23798 = ~n23581 & n23796;
  assign n23799 = ~n23797 & ~n23798;
  assign n23800 = n11476 & n23768;
  assign n23801 = n11463 & n23771;
  assign n23802 = n10883 & n23394;
  assign n23803 = n23779 & ~n23781;
  assign n23804 = ~n23782 & ~n23803;
  assign n23805 = n10884 & n23804;
  assign n23806 = ~n23801 & ~n23802;
  assign n23807 = ~n23800 & n23806;
  assign n23808 = ~n23805 & n23807;
  assign n23809 = pi2  & n23808;
  assign n23810 = ~pi2  & ~n23808;
  assign n23811 = ~n23809 & ~n23810;
  assign n23812 = n11476 & n23771;
  assign n23813 = n11463 & n23394;
  assign n23814 = n10883 & n20355;
  assign n23815 = n23775 & ~n23777;
  assign n23816 = ~n23778 & ~n23815;
  assign n23817 = n10884 & n23816;
  assign n23818 = ~n23813 & ~n23814;
  assign n23819 = ~n23812 & n23818;
  assign n23820 = ~n23817 & n23819;
  assign n23821 = pi2  & n23820;
  assign n23822 = ~pi2  & ~n23820;
  assign n23823 = ~n23821 & ~n23822;
  assign n23824 = n11476 & n23394;
  assign n23825 = n11463 & n20355;
  assign n23826 = n10883 & n20358;
  assign n23827 = n10884 & n23404;
  assign n23828 = ~n23825 & ~n23826;
  assign n23829 = ~n23824 & n23828;
  assign n23830 = ~n23827 & n23829;
  assign n23831 = pi2  & n23830;
  assign n23832 = ~pi2  & ~n23830;
  assign n23833 = ~n23831 & ~n23832;
  assign n23834 = n23296 & ~n23298;
  assign n23835 = ~n23299 & ~n23834;
  assign n23836 = n23292 & ~n23294;
  assign n23837 = ~n23295 & ~n23836;
  assign n23838 = n11476 & n20361;
  assign n23839 = n11463 & n20365;
  assign n23840 = n10883 & n20368;
  assign n23841 = n10884 & n22848;
  assign n23842 = ~n23839 & ~n23840;
  assign n23843 = ~n23838 & n23842;
  assign n23844 = ~n23841 & n23843;
  assign n23845 = pi2  & n23844;
  assign n23846 = ~pi2  & ~n23844;
  assign n23847 = ~n23845 & ~n23846;
  assign n23848 = n11476 & n20365;
  assign n23849 = n11463 & n20368;
  assign n23850 = n10883 & n20371;
  assign n23851 = n10884 & n22814;
  assign n23852 = ~n23849 & ~n23850;
  assign n23853 = ~n23848 & n23852;
  assign n23854 = ~n23851 & n23853;
  assign n23855 = pi2  & n23854;
  assign n23856 = ~pi2  & ~n23854;
  assign n23857 = ~n23855 & ~n23856;
  assign n23858 = n11476 & n20368;
  assign n23859 = n11463 & n20371;
  assign n23860 = n10883 & n20374;
  assign n23861 = n10884 & n22235;
  assign n23862 = ~n23859 & ~n23860;
  assign n23863 = ~n23858 & n23862;
  assign n23864 = ~n23861 & n23863;
  assign n23865 = pi2  & n23864;
  assign n23866 = ~pi2  & ~n23864;
  assign n23867 = ~n23865 & ~n23866;
  assign n23868 = n23276 & ~n23278;
  assign n23869 = ~n23279 & ~n23868;
  assign n23870 = n23272 & ~n23274;
  assign n23871 = ~n23275 & ~n23870;
  assign n23872 = n23268 & ~n23270;
  assign n23873 = ~n23271 & ~n23872;
  assign n23874 = n11476 & n20380;
  assign n23875 = n11463 & n20383;
  assign n23876 = n10883 & n20386;
  assign n23877 = n10884 & n20574;
  assign n23878 = ~n23875 & ~n23876;
  assign n23879 = ~n23874 & n23878;
  assign n23880 = ~n23877 & n23879;
  assign n23881 = pi2  & n23880;
  assign n23882 = ~pi2  & ~n23880;
  assign n23883 = ~n23881 & ~n23882;
  assign n23884 = n11476 & n20383;
  assign n23885 = n11463 & n20386;
  assign n23886 = n10883 & n20389;
  assign n23887 = n10884 & n21737;
  assign n23888 = ~n23885 & ~n23886;
  assign n23889 = ~n23884 & n23888;
  assign n23890 = ~n23887 & n23889;
  assign n23891 = pi2  & n23890;
  assign n23892 = ~pi2  & ~n23890;
  assign n23893 = ~n23891 & ~n23892;
  assign n23894 = n11476 & n20386;
  assign n23895 = n11463 & n20389;
  assign n23896 = n10883 & n20392;
  assign n23897 = n10884 & n21752;
  assign n23898 = ~n23895 & ~n23896;
  assign n23899 = ~n23894 & n23898;
  assign n23900 = ~n23897 & n23899;
  assign n23901 = pi2  & n23900;
  assign n23902 = ~pi2  & ~n23900;
  assign n23903 = ~n23901 & ~n23902;
  assign n23904 = n23252 & ~n23254;
  assign n23905 = ~n23255 & ~n23904;
  assign n23906 = n23248 & ~n23250;
  assign n23907 = ~n23251 & ~n23906;
  assign n23908 = n23244 & ~n23246;
  assign n23909 = ~n23247 & ~n23908;
  assign n23910 = n11476 & n20398;
  assign n23911 = n11463 & n20401;
  assign n23912 = n10883 & n20404;
  assign n23913 = n10884 & n21322;
  assign n23914 = ~n23911 & ~n23912;
  assign n23915 = ~n23910 & n23914;
  assign n23916 = ~n23913 & n23915;
  assign n23917 = pi2  & n23916;
  assign n23918 = ~pi2  & ~n23916;
  assign n23919 = ~n23917 & ~n23918;
  assign n23920 = n11476 & n20401;
  assign n23921 = n11463 & n20404;
  assign n23922 = n10883 & n20407;
  assign n23923 = n10884 & n21286;
  assign n23924 = ~n23921 & ~n23922;
  assign n23925 = ~n23920 & n23924;
  assign n23926 = ~n23923 & n23925;
  assign n23927 = pi2  & n23926;
  assign n23928 = ~pi2  & ~n23926;
  assign n23929 = ~n23927 & ~n23928;
  assign n23930 = n11476 & n20404;
  assign n23931 = n11463 & n20407;
  assign n23932 = n10883 & n20410;
  assign n23933 = n10884 & n20991;
  assign n23934 = ~n23931 & ~n23932;
  assign n23935 = ~n23930 & n23934;
  assign n23936 = ~n23933 & n23935;
  assign n23937 = pi2  & n23936;
  assign n23938 = ~pi2  & ~n23936;
  assign n23939 = ~n23937 & ~n23938;
  assign n23940 = n23228 & ~n23230;
  assign n23941 = ~n23231 & ~n23940;
  assign n23942 = n23224 & ~n23226;
  assign n23943 = ~n23227 & ~n23942;
  assign n23944 = n23220 & ~n23222;
  assign n23945 = ~n23223 & ~n23944;
  assign n23946 = n11476 & n20416;
  assign n23947 = n11463 & n20419;
  assign n23948 = n10883 & n20422;
  assign n23949 = n10884 & n20771;
  assign n23950 = ~n23947 & ~n23948;
  assign n23951 = ~n23946 & n23950;
  assign n23952 = ~n23949 & n23951;
  assign n23953 = pi2  & n23952;
  assign n23954 = ~pi2  & ~n23952;
  assign n23955 = ~n23953 & ~n23954;
  assign n23956 = n11476 & n20419;
  assign n23957 = n11463 & n20422;
  assign n23958 = n10883 & n20425;
  assign n23959 = n10884 & n20786;
  assign n23960 = ~n23957 & ~n23958;
  assign n23961 = ~n23956 & n23960;
  assign n23962 = ~n23959 & n23961;
  assign n23963 = pi2  & n23962;
  assign n23964 = ~pi2  & ~n23962;
  assign n23965 = ~n23963 & ~n23964;
  assign n23966 = n11476 & n20422;
  assign n23967 = n11463 & n20425;
  assign n23968 = n10883 & n20428;
  assign n23969 = n10884 & n20801;
  assign n23970 = ~n23967 & ~n23968;
  assign n23971 = ~n23966 & n23970;
  assign n23972 = ~n23969 & n23971;
  assign n23973 = pi2  & n23972;
  assign n23974 = ~pi2  & ~n23972;
  assign n23975 = ~n23973 & ~n23974;
  assign n23976 = n23204 & ~n23206;
  assign n23977 = ~n23207 & ~n23976;
  assign n23978 = n11476 & n20428;
  assign n23979 = n11463 & n20431;
  assign n23980 = n10883 & n20434;
  assign n23981 = n10884 & n20598;
  assign n23982 = ~n23979 & ~n23980;
  assign n23983 = ~n23978 & n23982;
  assign n23984 = ~n23981 & n23983;
  assign n23985 = pi2  & n23984;
  assign n23986 = ~pi2  & ~n23984;
  assign n23987 = ~n23985 & ~n23986;
  assign n23988 = pi5  & ~n23180;
  assign n23989 = n23187 & ~n23988;
  assign n23990 = ~n23187 & n23988;
  assign n23991 = ~n23989 & ~n23990;
  assign n23992 = n11476 & n20440;
  assign n23993 = ~n20440 & n20624;
  assign n23994 = n10884 & ~n23993;
  assign n23995 = n19959 & n20445;
  assign n23996 = pi2  & ~n20447;
  assign n23997 = ~n23995 & n23996;
  assign n23998 = ~n23992 & n23997;
  assign n23999 = ~n23994 & n23998;
  assign n24000 = ~n23173 & ~n23999;
  assign n24001 = n11476 & n20437;
  assign n24002 = n11463 & n20440;
  assign n24003 = n10883 & n20445;
  assign n24004 = n10884 & n20610;
  assign n24005 = ~n24002 & ~n24003;
  assign n24006 = ~n24001 & n24005;
  assign n24007 = ~n24004 & n24006;
  assign n24008 = ~pi2  & ~n24007;
  assign n24009 = pi2  & n24007;
  assign n24010 = ~n24008 & ~n24009;
  assign n24011 = ~n24000 & ~n24010;
  assign n24012 = n11476 & n20434;
  assign n24013 = n11463 & n20437;
  assign n24014 = n10883 & n20440;
  assign n24015 = n10884 & n20668;
  assign n24016 = ~n24013 & ~n24014;
  assign n24017 = ~n24012 & n24016;
  assign n24018 = ~n24015 & n24017;
  assign n24019 = pi2  & n24018;
  assign n24020 = ~pi2  & ~n24018;
  assign n24021 = ~n24019 & ~n24020;
  assign n24022 = n24011 & ~n24021;
  assign n24023 = ~n24011 & n24021;
  assign n24024 = n23174 & ~n23179;
  assign n24025 = ~n23180 & ~n24024;
  assign n24026 = ~n24023 & n24025;
  assign n24027 = ~n24022 & ~n24026;
  assign n24028 = n23991 & ~n24027;
  assign n24029 = ~n23991 & n24027;
  assign n24030 = n11476 & n20431;
  assign n24031 = n11463 & n20434;
  assign n24032 = n10883 & n20437;
  assign n24033 = n10884 & n20651;
  assign n24034 = ~n24031 & ~n24032;
  assign n24035 = ~n24030 & n24034;
  assign n24036 = ~n24033 & n24035;
  assign n24037 = pi2  & ~n24036;
  assign n24038 = ~pi2  & n24036;
  assign n24039 = ~n24037 & ~n24038;
  assign n24040 = ~n24029 & n24039;
  assign n24041 = ~n24028 & ~n24040;
  assign n24042 = ~n23987 & ~n24041;
  assign n24043 = n23987 & n24041;
  assign n24044 = n23200 & ~n23202;
  assign n24045 = ~n23203 & ~n24044;
  assign n24046 = ~n24043 & n24045;
  assign n24047 = ~n24042 & ~n24046;
  assign n24048 = n23977 & ~n24047;
  assign n24049 = ~n23977 & n24047;
  assign n24050 = n11476 & n20425;
  assign n24051 = n11463 & n20428;
  assign n24052 = n10883 & n20431;
  assign n24053 = n10884 & n20727;
  assign n24054 = ~n24051 & ~n24052;
  assign n24055 = ~n24050 & n24054;
  assign n24056 = ~n24053 & n24055;
  assign n24057 = pi2  & ~n24056;
  assign n24058 = ~pi2  & n24056;
  assign n24059 = ~n24057 & ~n24058;
  assign n24060 = ~n24049 & n24059;
  assign n24061 = ~n24048 & ~n24060;
  assign n24062 = ~n23975 & ~n24061;
  assign n24063 = n23975 & n24061;
  assign n24064 = n23208 & ~n23210;
  assign n24065 = ~n23211 & ~n24064;
  assign n24066 = ~n24063 & n24065;
  assign n24067 = ~n24062 & ~n24066;
  assign n24068 = ~n23965 & ~n24067;
  assign n24069 = n23965 & n24067;
  assign n24070 = n23212 & ~n23214;
  assign n24071 = ~n23215 & ~n24070;
  assign n24072 = ~n24069 & n24071;
  assign n24073 = ~n24068 & ~n24072;
  assign n24074 = ~n23955 & ~n24073;
  assign n24075 = n23955 & n24073;
  assign n24076 = n23216 & ~n23218;
  assign n24077 = ~n23219 & ~n24076;
  assign n24078 = ~n24075 & n24077;
  assign n24079 = ~n24074 & ~n24078;
  assign n24080 = n23945 & ~n24079;
  assign n24081 = ~n23945 & n24079;
  assign n24082 = n11476 & n20413;
  assign n24083 = n11463 & n20416;
  assign n24084 = n10883 & n20419;
  assign n24085 = n10884 & n20928;
  assign n24086 = ~n24083 & ~n24084;
  assign n24087 = ~n24082 & n24086;
  assign n24088 = ~n24085 & n24087;
  assign n24089 = pi2  & ~n24088;
  assign n24090 = ~pi2  & n24088;
  assign n24091 = ~n24089 & ~n24090;
  assign n24092 = ~n24081 & n24091;
  assign n24093 = ~n24080 & ~n24092;
  assign n24094 = n23943 & ~n24093;
  assign n24095 = ~n23943 & n24093;
  assign n24096 = n11476 & n20410;
  assign n24097 = n11463 & n20413;
  assign n24098 = n10883 & n20416;
  assign n24099 = n10884 & n21019;
  assign n24100 = ~n24097 & ~n24098;
  assign n24101 = ~n24096 & n24100;
  assign n24102 = ~n24099 & n24101;
  assign n24103 = pi2  & ~n24102;
  assign n24104 = ~pi2  & n24102;
  assign n24105 = ~n24103 & ~n24104;
  assign n24106 = ~n24095 & n24105;
  assign n24107 = ~n24094 & ~n24106;
  assign n24108 = n23941 & ~n24107;
  assign n24109 = ~n23941 & n24107;
  assign n24110 = n11476 & n20407;
  assign n24111 = n11463 & n20410;
  assign n24112 = n10883 & n20413;
  assign n24113 = n10884 & n21004;
  assign n24114 = ~n24111 & ~n24112;
  assign n24115 = ~n24110 & n24114;
  assign n24116 = ~n24113 & n24115;
  assign n24117 = pi2  & ~n24116;
  assign n24118 = ~pi2  & n24116;
  assign n24119 = ~n24117 & ~n24118;
  assign n24120 = ~n24109 & n24119;
  assign n24121 = ~n24108 & ~n24120;
  assign n24122 = ~n23939 & ~n24121;
  assign n24123 = n23939 & n24121;
  assign n24124 = n23232 & ~n23234;
  assign n24125 = ~n23235 & ~n24124;
  assign n24126 = ~n24123 & n24125;
  assign n24127 = ~n24122 & ~n24126;
  assign n24128 = ~n23929 & ~n24127;
  assign n24129 = n23929 & n24127;
  assign n24130 = n23236 & ~n23238;
  assign n24131 = ~n23239 & ~n24130;
  assign n24132 = ~n24129 & n24131;
  assign n24133 = ~n24128 & ~n24132;
  assign n24134 = ~n23919 & ~n24133;
  assign n24135 = n23919 & n24133;
  assign n24136 = n23240 & ~n23242;
  assign n24137 = ~n23243 & ~n24136;
  assign n24138 = ~n24135 & n24137;
  assign n24139 = ~n24134 & ~n24138;
  assign n24140 = n23909 & ~n24139;
  assign n24141 = ~n23909 & n24139;
  assign n24142 = n11476 & n20395;
  assign n24143 = n11463 & n20398;
  assign n24144 = n10883 & n20401;
  assign n24145 = n10884 & n21305;
  assign n24146 = ~n24143 & ~n24144;
  assign n24147 = ~n24142 & n24146;
  assign n24148 = ~n24145 & n24147;
  assign n24149 = pi2  & ~n24148;
  assign n24150 = ~pi2  & n24148;
  assign n24151 = ~n24149 & ~n24150;
  assign n24152 = ~n24141 & n24151;
  assign n24153 = ~n24140 & ~n24152;
  assign n24154 = n23907 & ~n24153;
  assign n24155 = ~n23907 & n24153;
  assign n24156 = n11476 & n20392;
  assign n24157 = n11463 & n20395;
  assign n24158 = n10883 & n20398;
  assign n24159 = n10884 & n20586;
  assign n24160 = ~n24157 & ~n24158;
  assign n24161 = ~n24156 & n24160;
  assign n24162 = ~n24159 & n24161;
  assign n24163 = pi2  & ~n24162;
  assign n24164 = ~pi2  & n24162;
  assign n24165 = ~n24163 & ~n24164;
  assign n24166 = ~n24155 & n24165;
  assign n24167 = ~n24154 & ~n24166;
  assign n24168 = n23905 & ~n24167;
  assign n24169 = ~n23905 & n24167;
  assign n24170 = n11476 & n20389;
  assign n24171 = n11463 & n20392;
  assign n24172 = n10883 & n20395;
  assign n24173 = n10884 & n21716;
  assign n24174 = ~n24171 & ~n24172;
  assign n24175 = ~n24170 & n24174;
  assign n24176 = ~n24173 & n24175;
  assign n24177 = pi2  & ~n24176;
  assign n24178 = ~pi2  & n24176;
  assign n24179 = ~n24177 & ~n24178;
  assign n24180 = ~n24169 & n24179;
  assign n24181 = ~n24168 & ~n24180;
  assign n24182 = ~n23903 & ~n24181;
  assign n24183 = n23903 & n24181;
  assign n24184 = n23256 & ~n23258;
  assign n24185 = ~n23259 & ~n24184;
  assign n24186 = ~n24183 & n24185;
  assign n24187 = ~n24182 & ~n24186;
  assign n24188 = ~n23893 & ~n24187;
  assign n24189 = n23893 & n24187;
  assign n24190 = n23260 & ~n23262;
  assign n24191 = ~n23263 & ~n24190;
  assign n24192 = ~n24189 & n24191;
  assign n24193 = ~n24188 & ~n24192;
  assign n24194 = ~n23883 & ~n24193;
  assign n24195 = n23883 & n24193;
  assign n24196 = n23264 & ~n23266;
  assign n24197 = ~n23267 & ~n24196;
  assign n24198 = ~n24195 & n24197;
  assign n24199 = ~n24194 & ~n24198;
  assign n24200 = n23873 & ~n24199;
  assign n24201 = ~n23873 & n24199;
  assign n24202 = n11476 & n20377;
  assign n24203 = n11463 & n20380;
  assign n24204 = n10883 & n20383;
  assign n24205 = n10884 & n22083;
  assign n24206 = ~n24203 & ~n24204;
  assign n24207 = ~n24202 & n24206;
  assign n24208 = ~n24205 & n24207;
  assign n24209 = pi2  & ~n24208;
  assign n24210 = ~pi2  & n24208;
  assign n24211 = ~n24209 & ~n24210;
  assign n24212 = ~n24201 & n24211;
  assign n24213 = ~n24200 & ~n24212;
  assign n24214 = n23871 & ~n24213;
  assign n24215 = ~n23871 & n24213;
  assign n24216 = n11476 & n20374;
  assign n24217 = n11463 & n20377;
  assign n24218 = n10883 & n20380;
  assign n24219 = n10884 & n22263;
  assign n24220 = ~n24217 & ~n24218;
  assign n24221 = ~n24216 & n24220;
  assign n24222 = ~n24219 & n24221;
  assign n24223 = pi2  & ~n24222;
  assign n24224 = ~pi2  & n24222;
  assign n24225 = ~n24223 & ~n24224;
  assign n24226 = ~n24215 & n24225;
  assign n24227 = ~n24214 & ~n24226;
  assign n24228 = n23869 & ~n24227;
  assign n24229 = ~n23869 & n24227;
  assign n24230 = n11476 & n20371;
  assign n24231 = n11463 & n20374;
  assign n24232 = n10883 & n20377;
  assign n24233 = n10884 & n22250;
  assign n24234 = ~n24231 & ~n24232;
  assign n24235 = ~n24230 & n24234;
  assign n24236 = ~n24233 & n24235;
  assign n24237 = pi2  & ~n24236;
  assign n24238 = ~pi2  & n24236;
  assign n24239 = ~n24237 & ~n24238;
  assign n24240 = ~n24229 & n24239;
  assign n24241 = ~n24228 & ~n24240;
  assign n24242 = ~n23867 & ~n24241;
  assign n24243 = n23867 & n24241;
  assign n24244 = n23280 & ~n23282;
  assign n24245 = ~n23283 & ~n24244;
  assign n24246 = ~n24243 & n24245;
  assign n24247 = ~n24242 & ~n24246;
  assign n24248 = ~n23857 & ~n24247;
  assign n24249 = n23857 & n24247;
  assign n24250 = n23284 & ~n23286;
  assign n24251 = ~n23287 & ~n24250;
  assign n24252 = ~n24249 & n24251;
  assign n24253 = ~n24248 & ~n24252;
  assign n24254 = ~n23847 & ~n24253;
  assign n24255 = n23847 & n24253;
  assign n24256 = n23288 & ~n23290;
  assign n24257 = ~n23291 & ~n24256;
  assign n24258 = ~n24255 & n24257;
  assign n24259 = ~n24254 & ~n24258;
  assign n24260 = n23837 & ~n24259;
  assign n24261 = ~n23837 & n24259;
  assign n24262 = n11476 & n20358;
  assign n24263 = n11463 & n20361;
  assign n24264 = n10883 & n20365;
  assign n24265 = n10884 & n22833;
  assign n24266 = ~n24263 & ~n24264;
  assign n24267 = ~n24262 & n24266;
  assign n24268 = ~n24265 & n24267;
  assign n24269 = pi2  & ~n24268;
  assign n24270 = ~pi2  & n24268;
  assign n24271 = ~n24269 & ~n24270;
  assign n24272 = ~n24261 & n24271;
  assign n24273 = ~n24260 & ~n24272;
  assign n24274 = n23835 & ~n24273;
  assign n24275 = ~n23835 & n24273;
  assign n24276 = n11476 & n20355;
  assign n24277 = n11463 & n20358;
  assign n24278 = n10883 & n20361;
  assign n24279 = n10884 & n20562;
  assign n24280 = ~n24277 & ~n24278;
  assign n24281 = ~n24276 & n24280;
  assign n24282 = ~n24279 & n24281;
  assign n24283 = pi2  & ~n24282;
  assign n24284 = ~pi2  & n24282;
  assign n24285 = ~n24283 & ~n24284;
  assign n24286 = ~n24275 & n24285;
  assign n24287 = ~n24274 & ~n24286;
  assign n24288 = ~n23833 & ~n24287;
  assign n24289 = n23833 & n24287;
  assign n24290 = n23300 & ~n23302;
  assign n24291 = ~n23303 & ~n24290;
  assign n24292 = ~n24289 & n24291;
  assign n24293 = ~n24288 & ~n24292;
  assign n24294 = ~n23823 & ~n24293;
  assign n24295 = n23823 & n24293;
  assign n24296 = n23304 & ~n23306;
  assign n24297 = ~n23307 & ~n24296;
  assign n24298 = ~n24295 & n24297;
  assign n24299 = ~n24294 & ~n24298;
  assign n24300 = ~n23811 & ~n24299;
  assign n24301 = n23811 & n24299;
  assign n24302 = n23308 & ~n23310;
  assign n24303 = ~n23311 & ~n24302;
  assign n24304 = ~n24301 & n24303;
  assign n24305 = ~n24300 & ~n24304;
  assign n24306 = n23799 & ~n24305;
  assign n24307 = ~n23797 & ~n24306;
  assign n24308 = ~n23576 & ~n23580;
  assign n24309 = n71 & n23771;
  assign n24310 = n10329 & n23394;
  assign n24311 = n9836 & n20355;
  assign n24312 = n9830 & n23816;
  assign n24313 = ~n24310 & ~n24311;
  assign n24314 = ~n24309 & n24313;
  assign n24315 = ~n24312 & n24314;
  assign n24316 = ~pi5  & ~n24315;
  assign n24317 = pi5  & n24315;
  assign n24318 = ~n24316 & ~n24317;
  assign n24319 = ~n23570 & ~n23573;
  assign n24320 = ~n23554 & ~n23558;
  assign n24321 = n8161 & n20368;
  assign n24322 = n7847 & n20371;
  assign n24323 = n7554 & n20374;
  assign n24324 = n7548 & n22235;
  assign n24325 = ~n24322 & ~n24323;
  assign n24326 = ~n24321 & n24325;
  assign n24327 = ~n24324 & n24326;
  assign n24328 = ~pi11  & ~n24327;
  assign n24329 = pi11  & n24327;
  assign n24330 = ~n24328 & ~n24329;
  assign n24331 = ~n23548 & ~n23551;
  assign n24332 = ~n23532 & ~n23536;
  assign n24333 = n6608 & n20386;
  assign n24334 = n6356 & n20389;
  assign n24335 = n6140 & n20392;
  assign n24336 = n6134 & n21752;
  assign n24337 = ~n24334 & ~n24335;
  assign n24338 = ~n24333 & n24337;
  assign n24339 = ~n24336 & n24338;
  assign n24340 = ~pi17  & ~n24339;
  assign n24341 = pi17  & n24339;
  assign n24342 = ~n24340 & ~n24341;
  assign n24343 = ~n23526 & ~n23529;
  assign n24344 = ~n23510 & ~n23514;
  assign n24345 = n5267 & n20404;
  assign n24346 = n5185 & n20407;
  assign n24347 = n5121 & n20410;
  assign n24348 = n78 & n20991;
  assign n24349 = ~n24346 & ~n24347;
  assign n24350 = ~n24345 & n24349;
  assign n24351 = ~n24348 & n24350;
  assign n24352 = ~pi23  & ~n24351;
  assign n24353 = pi23  & n24351;
  assign n24354 = ~n24352 & ~n24353;
  assign n24355 = ~n23504 & ~n23507;
  assign n24356 = ~n23488 & ~n23492;
  assign n24357 = n4472 & n20422;
  assign n24358 = n4070 & n20425;
  assign n24359 = n3943 & n20428;
  assign n24360 = n3944 & n20801;
  assign n24361 = ~n24358 & ~n24359;
  assign n24362 = ~n24357 & n24361;
  assign n24363 = ~n24360 & n24362;
  assign n24364 = ~pi29  & ~n24363;
  assign n24365 = pi29  & n24363;
  assign n24366 = ~n24364 & ~n24365;
  assign n24367 = ~n23482 & ~n23485;
  assign n24368 = n969 & n1085;
  assign n24369 = n1300 & n1756;
  assign n24370 = n2150 & n2478;
  assign n24371 = n3627 & n12450;
  assign n24372 = n24370 & n24371;
  assign n24373 = n24368 & n24369;
  assign n24374 = n2626 & n24373;
  assign n24375 = n5342 & n24372;
  assign n24376 = n12625 & n24375;
  assign n24377 = n4426 & n24374;
  assign n24378 = n24376 & n24377;
  assign n24379 = n4949 & n24378;
  assign n24380 = n12733 & n24379;
  assign n24381 = n3896 & n20431;
  assign n24382 = n564 & n20437;
  assign n24383 = n3683 & n20434;
  assign n24384 = n566 & n20651;
  assign n24385 = ~n24382 & ~n24383;
  assign n24386 = ~n24381 & n24385;
  assign n24387 = ~n24384 & n24386;
  assign n24388 = ~n24380 & ~n24387;
  assign n24389 = n24380 & n24387;
  assign n24390 = ~n24388 & ~n24389;
  assign n24391 = ~n24367 & n24390;
  assign n24392 = n24367 & ~n24390;
  assign n24393 = ~n24391 & ~n24392;
  assign n24394 = ~n24366 & n24393;
  assign n24395 = n24366 & ~n24393;
  assign n24396 = ~n24394 & ~n24395;
  assign n24397 = n24356 & ~n24396;
  assign n24398 = ~n24356 & n24396;
  assign n24399 = ~n24397 & ~n24398;
  assign n24400 = n4721 & n20413;
  assign n24401 = n4691 & n20416;
  assign n24402 = n4515 & n20419;
  assign n24403 = n4516 & n20928;
  assign n24404 = ~n24401 & ~n24402;
  assign n24405 = ~n24400 & n24404;
  assign n24406 = ~n24403 & n24405;
  assign n24407 = pi26  & n24406;
  assign n24408 = ~pi26  & ~n24406;
  assign n24409 = ~n24407 & ~n24408;
  assign n24410 = n24399 & ~n24409;
  assign n24411 = ~n24399 & n24409;
  assign n24412 = ~n24410 & ~n24411;
  assign n24413 = ~n24355 & n24412;
  assign n24414 = n24355 & ~n24412;
  assign n24415 = ~n24413 & ~n24414;
  assign n24416 = ~n24354 & n24415;
  assign n24417 = n24354 & ~n24415;
  assign n24418 = ~n24416 & ~n24417;
  assign n24419 = n24344 & ~n24418;
  assign n24420 = ~n24344 & n24418;
  assign n24421 = ~n24419 & ~n24420;
  assign n24422 = n5982 & n20395;
  assign n24423 = n5901 & n20398;
  assign n24424 = n5312 & n20401;
  assign n24425 = n5306 & n21305;
  assign n24426 = ~n24423 & ~n24424;
  assign n24427 = ~n24422 & n24426;
  assign n24428 = ~n24425 & n24427;
  assign n24429 = pi20  & n24428;
  assign n24430 = ~pi20  & ~n24428;
  assign n24431 = ~n24429 & ~n24430;
  assign n24432 = n24421 & ~n24431;
  assign n24433 = ~n24421 & n24431;
  assign n24434 = ~n24432 & ~n24433;
  assign n24435 = ~n24343 & n24434;
  assign n24436 = n24343 & ~n24434;
  assign n24437 = ~n24435 & ~n24436;
  assign n24438 = ~n24342 & n24437;
  assign n24439 = n24342 & ~n24437;
  assign n24440 = ~n24438 & ~n24439;
  assign n24441 = n24332 & ~n24440;
  assign n24442 = ~n24332 & n24440;
  assign n24443 = ~n24441 & ~n24442;
  assign n24444 = n7380 & n20377;
  assign n24445 = n7243 & n20380;
  assign n24446 = n6653 & n20383;
  assign n24447 = n6647 & n22083;
  assign n24448 = ~n24445 & ~n24446;
  assign n24449 = ~n24444 & n24448;
  assign n24450 = ~n24447 & n24449;
  assign n24451 = pi14  & n24450;
  assign n24452 = ~pi14  & ~n24450;
  assign n24453 = ~n24451 & ~n24452;
  assign n24454 = n24443 & ~n24453;
  assign n24455 = ~n24443 & n24453;
  assign n24456 = ~n24454 & ~n24455;
  assign n24457 = ~n24331 & n24456;
  assign n24458 = n24331 & ~n24456;
  assign n24459 = ~n24457 & ~n24458;
  assign n24460 = ~n24330 & n24459;
  assign n24461 = n24330 & ~n24459;
  assign n24462 = ~n24460 & ~n24461;
  assign n24463 = n24320 & ~n24462;
  assign n24464 = ~n24320 & n24462;
  assign n24465 = ~n24463 & ~n24464;
  assign n24466 = n9355 & n20358;
  assign n24467 = n8939 & n20361;
  assign n24468 = n8206 & n20365;
  assign n24469 = n8200 & n22833;
  assign n24470 = ~n24467 & ~n24468;
  assign n24471 = ~n24466 & n24470;
  assign n24472 = ~n24469 & n24471;
  assign n24473 = pi8  & n24472;
  assign n24474 = ~pi8  & ~n24472;
  assign n24475 = ~n24473 & ~n24474;
  assign n24476 = n24465 & ~n24475;
  assign n24477 = ~n24465 & n24475;
  assign n24478 = ~n24476 & ~n24477;
  assign n24479 = ~n24319 & n24478;
  assign n24480 = n24319 & ~n24478;
  assign n24481 = ~n24479 & ~n24480;
  assign n24482 = ~n24318 & n24481;
  assign n24483 = n24318 & ~n24481;
  assign n24484 = ~n24482 & ~n24483;
  assign n24485 = n24308 & ~n24484;
  assign n24486 = ~n24308 & n24484;
  assign n24487 = ~n24485 & ~n24486;
  assign n24488 = ~n23760 & ~n23764;
  assign n24489 = ~n23753 & ~n23757;
  assign n24490 = ~n23730 & ~n23740;
  assign n24491 = ~n23725 & ~n23727;
  assign n24492 = n533 & ~n568;
  assign n24493 = n712 & n24492;
  assign n24494 = n23718 & n24493;
  assign n24495 = ~n24491 & n24494;
  assign n24496 = n24491 & ~n24494;
  assign n24497 = ~n24495 & ~n24496;
  assign n24498 = n3896 & n12168;
  assign n24499 = n3683 & n12175;
  assign n24500 = n564 & n12178;
  assign n24501 = n566 & n12862;
  assign n24502 = ~n24499 & ~n24500;
  assign n24503 = ~n24498 & n24502;
  assign n24504 = ~n24501 & n24503;
  assign n24505 = n24497 & ~n24504;
  assign n24506 = ~n24497 & n24504;
  assign n24507 = ~n24505 & ~n24506;
  assign n24508 = n24490 & ~n24507;
  assign n24509 = ~n24490 & n24507;
  assign n24510 = ~n24508 & ~n24509;
  assign n24511 = n4472 & ~n12163;
  assign n24512 = n3944 & n13007;
  assign n24513 = n4070 & n12166;
  assign n24514 = n3943 & n12172;
  assign n24515 = ~n24511 & ~n24513;
  assign n24516 = ~n24514 & n24515;
  assign n24517 = ~n24512 & n24516;
  assign n24518 = pi29  & n24517;
  assign n24519 = ~pi29  & ~n24517;
  assign n24520 = ~n24518 & ~n24519;
  assign n24521 = n24510 & ~n24520;
  assign n24522 = ~n24510 & n24520;
  assign n24523 = ~n24521 & ~n24522;
  assign n24524 = ~n24489 & n24523;
  assign n24525 = n24489 & ~n24523;
  assign n24526 = ~n24524 & ~n24525;
  assign n24527 = ~n24488 & n24526;
  assign n24528 = n24488 & ~n24526;
  assign n24529 = ~n24527 & ~n24528;
  assign n24530 = n11476 & n24529;
  assign n24531 = n11463 & n23765;
  assign n24532 = n10883 & n23768;
  assign n24533 = ~n23784 & ~n23787;
  assign n24534 = n23765 & n24529;
  assign n24535 = ~n23765 & ~n24529;
  assign n24536 = ~n24534 & ~n24535;
  assign n24537 = ~n24533 & n24536;
  assign n24538 = n24533 & ~n24536;
  assign n24539 = ~n24537 & ~n24538;
  assign n24540 = n10884 & n24539;
  assign n24541 = ~n24531 & ~n24532;
  assign n24542 = ~n24530 & n24541;
  assign n24543 = ~n24540 & n24542;
  assign n24544 = pi2  & n24543;
  assign n24545 = ~pi2  & ~n24543;
  assign n24546 = ~n24544 & ~n24545;
  assign n24547 = n24487 & ~n24546;
  assign n24548 = ~n24487 & n24546;
  assign n24549 = ~n24547 & ~n24548;
  assign n24550 = ~n24307 & n24549;
  assign n24551 = n24307 & ~n24549;
  assign n24552 = ~n24550 & ~n24551;
  assign n24553 = ~n23799 & n24305;
  assign n24554 = ~n24306 & ~n24553;
  assign n24555 = n24552 & n24554;
  assign n24556 = ~n24552 & ~n24554;
  assign po0  = ~n24555 & ~n24556;
  assign n24558 = ~n24547 & ~n24550;
  assign n24559 = ~n24482 & ~n24486;
  assign n24560 = n71 & n23768;
  assign n24561 = n10329 & n23771;
  assign n24562 = n9836 & n23394;
  assign n24563 = n9830 & n23804;
  assign n24564 = ~n24561 & ~n24562;
  assign n24565 = ~n24560 & n24564;
  assign n24566 = ~n24563 & n24565;
  assign n24567 = ~pi5  & ~n24566;
  assign n24568 = pi5  & n24566;
  assign n24569 = ~n24567 & ~n24568;
  assign n24570 = ~n24476 & ~n24479;
  assign n24571 = ~n24460 & ~n24464;
  assign n24572 = n8161 & n20365;
  assign n24573 = n7847 & n20368;
  assign n24574 = n7554 & n20371;
  assign n24575 = n7548 & n22814;
  assign n24576 = ~n24573 & ~n24574;
  assign n24577 = ~n24572 & n24576;
  assign n24578 = ~n24575 & n24577;
  assign n24579 = ~pi11  & ~n24578;
  assign n24580 = pi11  & n24578;
  assign n24581 = ~n24579 & ~n24580;
  assign n24582 = ~n24454 & ~n24457;
  assign n24583 = ~n24438 & ~n24442;
  assign n24584 = n6608 & n20383;
  assign n24585 = n6356 & n20386;
  assign n24586 = n6140 & n20389;
  assign n24587 = n6134 & n21737;
  assign n24588 = ~n24585 & ~n24586;
  assign n24589 = ~n24584 & n24588;
  assign n24590 = ~n24587 & n24589;
  assign n24591 = ~pi17  & ~n24590;
  assign n24592 = pi17  & n24590;
  assign n24593 = ~n24591 & ~n24592;
  assign n24594 = ~n24432 & ~n24435;
  assign n24595 = ~n24416 & ~n24420;
  assign n24596 = n5267 & n20401;
  assign n24597 = n5185 & n20404;
  assign n24598 = n5121 & n20407;
  assign n24599 = n78 & n21286;
  assign n24600 = ~n24597 & ~n24598;
  assign n24601 = ~n24596 & n24600;
  assign n24602 = ~n24599 & n24601;
  assign n24603 = ~pi23  & ~n24602;
  assign n24604 = pi23  & n24602;
  assign n24605 = ~n24603 & ~n24604;
  assign n24606 = ~n24410 & ~n24413;
  assign n24607 = ~n24394 & ~n24398;
  assign n24608 = n4472 & n20419;
  assign n24609 = n4070 & n20422;
  assign n24610 = n3943 & n20425;
  assign n24611 = n3944 & n20786;
  assign n24612 = ~n24609 & ~n24610;
  assign n24613 = ~n24608 & n24612;
  assign n24614 = ~n24611 & n24613;
  assign n24615 = pi29  & n24614;
  assign n24616 = ~pi29  & ~n24614;
  assign n24617 = ~n24615 & ~n24616;
  assign n24618 = ~n24388 & ~n24391;
  assign n24619 = ~n177 & ~n509;
  assign n24620 = n403 & n24619;
  assign n24621 = n1014 & n2109;
  assign n24622 = n2150 & n2231;
  assign n24623 = n2271 & n2366;
  assign n24624 = n2390 & n24623;
  assign n24625 = n24621 & n24622;
  assign n24626 = n1153 & n24620;
  assign n24627 = n2740 & n24626;
  assign n24628 = n24624 & n24625;
  assign n24629 = n6952 & n24628;
  assign n24630 = n7027 & n24627;
  assign n24631 = n24629 & n24630;
  assign n24632 = n3119 & n13467;
  assign n24633 = n24631 & n24632;
  assign n24634 = n1262 & n24633;
  assign n24635 = n3896 & n20428;
  assign n24636 = n564 & n20434;
  assign n24637 = n3683 & n20431;
  assign n24638 = n566 & n20598;
  assign n24639 = ~n24636 & ~n24637;
  assign n24640 = ~n24635 & n24639;
  assign n24641 = ~n24638 & n24640;
  assign n24642 = ~n24634 & ~n24641;
  assign n24643 = n24634 & n24641;
  assign n24644 = ~n24642 & ~n24643;
  assign n24645 = ~n24618 & n24644;
  assign n24646 = n24618 & ~n24644;
  assign n24647 = ~n24645 & ~n24646;
  assign n24648 = ~n24617 & n24647;
  assign n24649 = n24617 & ~n24647;
  assign n24650 = ~n24648 & ~n24649;
  assign n24651 = ~n24607 & n24650;
  assign n24652 = n24607 & ~n24650;
  assign n24653 = ~n24651 & ~n24652;
  assign n24654 = n4721 & n20410;
  assign n24655 = n4691 & n20413;
  assign n24656 = n4515 & n20416;
  assign n24657 = n4516 & n21019;
  assign n24658 = ~n24655 & ~n24656;
  assign n24659 = ~n24654 & n24658;
  assign n24660 = ~n24657 & n24659;
  assign n24661 = pi26  & n24660;
  assign n24662 = ~pi26  & ~n24660;
  assign n24663 = ~n24661 & ~n24662;
  assign n24664 = n24653 & ~n24663;
  assign n24665 = ~n24653 & n24663;
  assign n24666 = ~n24664 & ~n24665;
  assign n24667 = ~n24606 & n24666;
  assign n24668 = n24606 & ~n24666;
  assign n24669 = ~n24667 & ~n24668;
  assign n24670 = ~n24605 & n24669;
  assign n24671 = n24605 & ~n24669;
  assign n24672 = ~n24670 & ~n24671;
  assign n24673 = n24595 & ~n24672;
  assign n24674 = ~n24595 & n24672;
  assign n24675 = ~n24673 & ~n24674;
  assign n24676 = n5982 & n20392;
  assign n24677 = n5901 & n20395;
  assign n24678 = n5312 & n20398;
  assign n24679 = n5306 & n20586;
  assign n24680 = ~n24677 & ~n24678;
  assign n24681 = ~n24676 & n24680;
  assign n24682 = ~n24679 & n24681;
  assign n24683 = pi20  & n24682;
  assign n24684 = ~pi20  & ~n24682;
  assign n24685 = ~n24683 & ~n24684;
  assign n24686 = n24675 & ~n24685;
  assign n24687 = ~n24675 & n24685;
  assign n24688 = ~n24686 & ~n24687;
  assign n24689 = ~n24594 & n24688;
  assign n24690 = n24594 & ~n24688;
  assign n24691 = ~n24689 & ~n24690;
  assign n24692 = ~n24593 & n24691;
  assign n24693 = n24593 & ~n24691;
  assign n24694 = ~n24692 & ~n24693;
  assign n24695 = n24583 & ~n24694;
  assign n24696 = ~n24583 & n24694;
  assign n24697 = ~n24695 & ~n24696;
  assign n24698 = n7380 & n20374;
  assign n24699 = n7243 & n20377;
  assign n24700 = n6653 & n20380;
  assign n24701 = n6647 & n22263;
  assign n24702 = ~n24699 & ~n24700;
  assign n24703 = ~n24698 & n24702;
  assign n24704 = ~n24701 & n24703;
  assign n24705 = pi14  & n24704;
  assign n24706 = ~pi14  & ~n24704;
  assign n24707 = ~n24705 & ~n24706;
  assign n24708 = n24697 & ~n24707;
  assign n24709 = ~n24697 & n24707;
  assign n24710 = ~n24708 & ~n24709;
  assign n24711 = ~n24582 & n24710;
  assign n24712 = n24582 & ~n24710;
  assign n24713 = ~n24711 & ~n24712;
  assign n24714 = ~n24581 & n24713;
  assign n24715 = n24581 & ~n24713;
  assign n24716 = ~n24714 & ~n24715;
  assign n24717 = n24571 & ~n24716;
  assign n24718 = ~n24571 & n24716;
  assign n24719 = ~n24717 & ~n24718;
  assign n24720 = n9355 & n20355;
  assign n24721 = n8939 & n20358;
  assign n24722 = n8206 & n20361;
  assign n24723 = n8200 & n20562;
  assign n24724 = ~n24721 & ~n24722;
  assign n24725 = ~n24720 & n24724;
  assign n24726 = ~n24723 & n24725;
  assign n24727 = pi8  & n24726;
  assign n24728 = ~pi8  & ~n24726;
  assign n24729 = ~n24727 & ~n24728;
  assign n24730 = n24719 & ~n24729;
  assign n24731 = ~n24719 & n24729;
  assign n24732 = ~n24730 & ~n24731;
  assign n24733 = ~n24570 & n24732;
  assign n24734 = n24570 & ~n24732;
  assign n24735 = ~n24733 & ~n24734;
  assign n24736 = ~n24569 & n24735;
  assign n24737 = n24569 & ~n24735;
  assign n24738 = ~n24736 & ~n24737;
  assign n24739 = n24559 & ~n24738;
  assign n24740 = ~n24559 & n24738;
  assign n24741 = ~n24739 & ~n24740;
  assign n24742 = ~n24524 & ~n24527;
  assign n24743 = ~n24509 & ~n24521;
  assign n24744 = ~n24495 & ~n24505;
  assign n24745 = n491 & n535;
  assign n24746 = n24494 & ~n24745;
  assign n24747 = ~n24494 & n24745;
  assign n24748 = ~n24746 & ~n24747;
  assign n24749 = ~n24744 & n24748;
  assign n24750 = n24744 & ~n24748;
  assign n24751 = ~n24749 & ~n24750;
  assign n24752 = n3944 & ~n12424;
  assign n24753 = n3943 & ~n12165;
  assign n24754 = ~n4070 & ~n4472;
  assign n24755 = ~n24753 & n24754;
  assign n24756 = ~n12163 & ~n24755;
  assign n24757 = ~n24752 & ~n24756;
  assign n24758 = ~pi29  & ~n24757;
  assign n24759 = pi29  & n24757;
  assign n24760 = ~n24758 & ~n24759;
  assign n24761 = n3896 & n12172;
  assign n24762 = n3683 & n12168;
  assign n24763 = n564 & n12175;
  assign n24764 = n566 & n12939;
  assign n24765 = ~n24762 & ~n24763;
  assign n24766 = ~n24761 & n24765;
  assign n24767 = ~n24764 & n24766;
  assign n24768 = ~n24760 & ~n24767;
  assign n24769 = n24760 & n24767;
  assign n24770 = ~n24768 & ~n24769;
  assign n24771 = n24751 & n24770;
  assign n24772 = ~n24751 & ~n24770;
  assign n24773 = ~n24771 & ~n24772;
  assign n24774 = ~n24743 & n24773;
  assign n24775 = n24743 & ~n24773;
  assign n24776 = ~n24774 & ~n24775;
  assign n24777 = ~n24742 & n24776;
  assign n24778 = n24742 & ~n24776;
  assign n24779 = ~n24777 & ~n24778;
  assign n24780 = n11476 & n24779;
  assign n24781 = n11463 & n24529;
  assign n24782 = n10883 & n23765;
  assign n24783 = ~n24534 & ~n24537;
  assign n24784 = ~n24529 & ~n24779;
  assign n24785 = n24529 & n24779;
  assign n24786 = ~n24784 & ~n24785;
  assign n24787 = ~n24783 & n24786;
  assign n24788 = n24783 & ~n24786;
  assign n24789 = ~n24787 & ~n24788;
  assign n24790 = n10884 & n24789;
  assign n24791 = ~n24781 & ~n24782;
  assign n24792 = ~n24780 & n24791;
  assign n24793 = ~n24790 & n24792;
  assign n24794 = pi2  & n24793;
  assign n24795 = ~pi2  & ~n24793;
  assign n24796 = ~n24794 & ~n24795;
  assign n24797 = n24741 & ~n24796;
  assign n24798 = ~n24741 & n24796;
  assign n24799 = ~n24797 & ~n24798;
  assign n24800 = ~n24558 & n24799;
  assign n24801 = n24558 & ~n24799;
  assign n24802 = ~n24800 & ~n24801;
  assign n24803 = n24555 & n24802;
  assign n24804 = ~n24555 & ~n24802;
  assign po1  = ~n24803 & ~n24804;
  assign n24806 = ~n24797 & ~n24800;
  assign n24807 = ~n24736 & ~n24740;
  assign n24808 = n71 & n23765;
  assign n24809 = n10329 & n23768;
  assign n24810 = n9836 & n23771;
  assign n24811 = n9830 & n23789;
  assign n24812 = ~n24809 & ~n24810;
  assign n24813 = ~n24808 & n24812;
  assign n24814 = ~n24811 & n24813;
  assign n24815 = ~pi5  & ~n24814;
  assign n24816 = pi5  & n24814;
  assign n24817 = ~n24815 & ~n24816;
  assign n24818 = ~n24730 & ~n24733;
  assign n24819 = ~n24714 & ~n24718;
  assign n24820 = n8161 & n20361;
  assign n24821 = n7847 & n20365;
  assign n24822 = n7554 & n20368;
  assign n24823 = n7548 & n22848;
  assign n24824 = ~n24821 & ~n24822;
  assign n24825 = ~n24820 & n24824;
  assign n24826 = ~n24823 & n24825;
  assign n24827 = ~pi11  & ~n24826;
  assign n24828 = pi11  & n24826;
  assign n24829 = ~n24827 & ~n24828;
  assign n24830 = ~n24708 & ~n24711;
  assign n24831 = ~n24692 & ~n24696;
  assign n24832 = n6608 & n20380;
  assign n24833 = n6356 & n20383;
  assign n24834 = n6140 & n20386;
  assign n24835 = n6134 & n20574;
  assign n24836 = ~n24833 & ~n24834;
  assign n24837 = ~n24832 & n24836;
  assign n24838 = ~n24835 & n24837;
  assign n24839 = ~pi17  & ~n24838;
  assign n24840 = pi17  & n24838;
  assign n24841 = ~n24839 & ~n24840;
  assign n24842 = ~n24686 & ~n24689;
  assign n24843 = ~n24670 & ~n24674;
  assign n24844 = n5267 & n20398;
  assign n24845 = n5185 & n20401;
  assign n24846 = n5121 & n20404;
  assign n24847 = n78 & n21322;
  assign n24848 = ~n24845 & ~n24846;
  assign n24849 = ~n24844 & n24848;
  assign n24850 = ~n24847 & n24849;
  assign n24851 = ~pi23  & ~n24850;
  assign n24852 = pi23  & n24850;
  assign n24853 = ~n24851 & ~n24852;
  assign n24854 = ~n24664 & ~n24667;
  assign n24855 = ~n24648 & ~n24651;
  assign n24856 = n4472 & n20416;
  assign n24857 = n4070 & n20419;
  assign n24858 = n3943 & n20422;
  assign n24859 = n3944 & n20771;
  assign n24860 = ~n24857 & ~n24858;
  assign n24861 = ~n24856 & n24860;
  assign n24862 = ~n24859 & n24861;
  assign n24863 = pi29  & n24862;
  assign n24864 = ~pi29  & ~n24862;
  assign n24865 = ~n24863 & ~n24864;
  assign n24866 = ~n24642 & ~n24645;
  assign n24867 = ~n126 & ~n539;
  assign n24868 = ~n541 & n24867;
  assign n24869 = n252 & n738;
  assign n24870 = n765 & n1157;
  assign n24871 = n1161 & n3085;
  assign n24872 = n24870 & n24871;
  assign n24873 = n24868 & n24869;
  assign n24874 = n1583 & n12765;
  assign n24875 = n13493 & n24874;
  assign n24876 = n24872 & n24873;
  assign n24877 = n2581 & n7060;
  assign n24878 = n24876 & n24877;
  assign n24879 = n4371 & n24875;
  assign n24880 = n24878 & n24879;
  assign n24881 = n2418 & n24880;
  assign n24882 = n4404 & n24881;
  assign n24883 = n3896 & n20425;
  assign n24884 = n564 & n20431;
  assign n24885 = n3683 & n20428;
  assign n24886 = n566 & n20727;
  assign n24887 = ~n24884 & ~n24885;
  assign n24888 = ~n24883 & n24887;
  assign n24889 = ~n24886 & n24888;
  assign n24890 = ~n24882 & ~n24889;
  assign n24891 = n24882 & n24889;
  assign n24892 = ~n24890 & ~n24891;
  assign n24893 = ~n24866 & n24892;
  assign n24894 = n24866 & ~n24892;
  assign n24895 = ~n24893 & ~n24894;
  assign n24896 = ~n24865 & n24895;
  assign n24897 = n24865 & ~n24895;
  assign n24898 = ~n24896 & ~n24897;
  assign n24899 = ~n24855 & n24898;
  assign n24900 = n24855 & ~n24898;
  assign n24901 = ~n24899 & ~n24900;
  assign n24902 = n4721 & n20407;
  assign n24903 = n4691 & n20410;
  assign n24904 = n4515 & n20413;
  assign n24905 = n4516 & n21004;
  assign n24906 = ~n24903 & ~n24904;
  assign n24907 = ~n24902 & n24906;
  assign n24908 = ~n24905 & n24907;
  assign n24909 = pi26  & n24908;
  assign n24910 = ~pi26  & ~n24908;
  assign n24911 = ~n24909 & ~n24910;
  assign n24912 = n24901 & ~n24911;
  assign n24913 = ~n24901 & n24911;
  assign n24914 = ~n24912 & ~n24913;
  assign n24915 = ~n24854 & n24914;
  assign n24916 = n24854 & ~n24914;
  assign n24917 = ~n24915 & ~n24916;
  assign n24918 = ~n24853 & n24917;
  assign n24919 = n24853 & ~n24917;
  assign n24920 = ~n24918 & ~n24919;
  assign n24921 = n24843 & ~n24920;
  assign n24922 = ~n24843 & n24920;
  assign n24923 = ~n24921 & ~n24922;
  assign n24924 = n5982 & n20389;
  assign n24925 = n5901 & n20392;
  assign n24926 = n5312 & n20395;
  assign n24927 = n5306 & n21716;
  assign n24928 = ~n24925 & ~n24926;
  assign n24929 = ~n24924 & n24928;
  assign n24930 = ~n24927 & n24929;
  assign n24931 = pi20  & n24930;
  assign n24932 = ~pi20  & ~n24930;
  assign n24933 = ~n24931 & ~n24932;
  assign n24934 = n24923 & ~n24933;
  assign n24935 = ~n24923 & n24933;
  assign n24936 = ~n24934 & ~n24935;
  assign n24937 = ~n24842 & n24936;
  assign n24938 = n24842 & ~n24936;
  assign n24939 = ~n24937 & ~n24938;
  assign n24940 = ~n24841 & n24939;
  assign n24941 = n24841 & ~n24939;
  assign n24942 = ~n24940 & ~n24941;
  assign n24943 = n24831 & ~n24942;
  assign n24944 = ~n24831 & n24942;
  assign n24945 = ~n24943 & ~n24944;
  assign n24946 = n7380 & n20371;
  assign n24947 = n7243 & n20374;
  assign n24948 = n6653 & n20377;
  assign n24949 = n6647 & n22250;
  assign n24950 = ~n24947 & ~n24948;
  assign n24951 = ~n24946 & n24950;
  assign n24952 = ~n24949 & n24951;
  assign n24953 = pi14  & n24952;
  assign n24954 = ~pi14  & ~n24952;
  assign n24955 = ~n24953 & ~n24954;
  assign n24956 = n24945 & ~n24955;
  assign n24957 = ~n24945 & n24955;
  assign n24958 = ~n24956 & ~n24957;
  assign n24959 = ~n24830 & n24958;
  assign n24960 = n24830 & ~n24958;
  assign n24961 = ~n24959 & ~n24960;
  assign n24962 = ~n24829 & n24961;
  assign n24963 = n24829 & ~n24961;
  assign n24964 = ~n24962 & ~n24963;
  assign n24965 = n24819 & ~n24964;
  assign n24966 = ~n24819 & n24964;
  assign n24967 = ~n24965 & ~n24966;
  assign n24968 = n9355 & n23394;
  assign n24969 = n8939 & n20355;
  assign n24970 = n8206 & n20358;
  assign n24971 = n8200 & n23404;
  assign n24972 = ~n24969 & ~n24970;
  assign n24973 = ~n24968 & n24972;
  assign n24974 = ~n24971 & n24973;
  assign n24975 = pi8  & n24974;
  assign n24976 = ~pi8  & ~n24974;
  assign n24977 = ~n24975 & ~n24976;
  assign n24978 = n24967 & ~n24977;
  assign n24979 = ~n24967 & n24977;
  assign n24980 = ~n24978 & ~n24979;
  assign n24981 = ~n24818 & n24980;
  assign n24982 = n24818 & ~n24980;
  assign n24983 = ~n24981 & ~n24982;
  assign n24984 = ~n24817 & n24983;
  assign n24985 = n24817 & ~n24983;
  assign n24986 = ~n24984 & ~n24985;
  assign n24987 = n24807 & ~n24986;
  assign n24988 = ~n24807 & n24986;
  assign n24989 = ~n24987 & ~n24988;
  assign n24990 = ~n24774 & ~n24777;
  assign n24991 = ~n24768 & ~n24771;
  assign n24992 = ~n24747 & ~n24749;
  assign n24993 = ~n3937 & n3942;
  assign n24994 = ~n12163 & ~n24993;
  assign n24995 = pi29  & ~n24994;
  assign n24996 = ~pi29  & n24994;
  assign n24997 = ~n24995 & ~n24996;
  assign n24998 = n12158 & n24745;
  assign n24999 = ~n12158 & ~n24745;
  assign n25000 = ~n24998 & ~n24999;
  assign n25001 = n24997 & n25000;
  assign n25002 = ~n24997 & ~n25000;
  assign n25003 = ~n25001 & ~n25002;
  assign n25004 = n3896 & n12166;
  assign n25005 = n3683 & n12172;
  assign n25006 = n564 & n12168;
  assign n25007 = n566 & n13106;
  assign n25008 = ~n25004 & ~n25006;
  assign n25009 = ~n25005 & n25008;
  assign n25010 = ~n25007 & n25009;
  assign n25011 = n25003 & ~n25010;
  assign n25012 = ~n25003 & n25010;
  assign n25013 = ~n25011 & ~n25012;
  assign n25014 = ~n24992 & n25013;
  assign n25015 = n24992 & ~n25013;
  assign n25016 = ~n25014 & ~n25015;
  assign n25017 = ~n24991 & n25016;
  assign n25018 = n24991 & ~n25016;
  assign n25019 = ~n25017 & ~n25018;
  assign n25020 = ~n24990 & n25019;
  assign n25021 = n24990 & ~n25019;
  assign n25022 = ~n25020 & ~n25021;
  assign n25023 = n11476 & n25022;
  assign n25024 = n11463 & n24779;
  assign n25025 = n10883 & n24529;
  assign n25026 = ~n24785 & ~n24787;
  assign n25027 = ~n24779 & ~n25022;
  assign n25028 = n24779 & n25022;
  assign n25029 = ~n25027 & ~n25028;
  assign n25030 = ~n25026 & n25029;
  assign n25031 = n25026 & ~n25029;
  assign n25032 = ~n25030 & ~n25031;
  assign n25033 = n10884 & n25032;
  assign n25034 = ~n25024 & ~n25025;
  assign n25035 = ~n25023 & n25034;
  assign n25036 = ~n25033 & n25035;
  assign n25037 = pi2  & n25036;
  assign n25038 = ~pi2  & ~n25036;
  assign n25039 = ~n25037 & ~n25038;
  assign n25040 = n24989 & ~n25039;
  assign n25041 = ~n24989 & n25039;
  assign n25042 = ~n25040 & ~n25041;
  assign n25043 = ~n24806 & n25042;
  assign n25044 = n24806 & ~n25042;
  assign n25045 = ~n25043 & ~n25044;
  assign n25046 = n24803 & n25045;
  assign n25047 = ~n24803 & ~n25045;
  assign po2  = ~n25046 & ~n25047;
  assign n25049 = ~n25040 & ~n25043;
  assign n25050 = ~n24984 & ~n24988;
  assign n25051 = n71 & n24529;
  assign n25052 = n10329 & n23765;
  assign n25053 = n9836 & n23768;
  assign n25054 = n9830 & n24539;
  assign n25055 = ~n25052 & ~n25053;
  assign n25056 = ~n25051 & n25055;
  assign n25057 = ~n25054 & n25056;
  assign n25058 = ~pi5  & ~n25057;
  assign n25059 = pi5  & n25057;
  assign n25060 = ~n25058 & ~n25059;
  assign n25061 = ~n24978 & ~n24981;
  assign n25062 = ~n24962 & ~n24966;
  assign n25063 = n8161 & n20358;
  assign n25064 = n7847 & n20361;
  assign n25065 = n7554 & n20365;
  assign n25066 = n7548 & n22833;
  assign n25067 = ~n25064 & ~n25065;
  assign n25068 = ~n25063 & n25067;
  assign n25069 = ~n25066 & n25068;
  assign n25070 = ~pi11  & ~n25069;
  assign n25071 = pi11  & n25069;
  assign n25072 = ~n25070 & ~n25071;
  assign n25073 = ~n24956 & ~n24959;
  assign n25074 = ~n24940 & ~n24944;
  assign n25075 = n6608 & n20377;
  assign n25076 = n6356 & n20380;
  assign n25077 = n6140 & n20383;
  assign n25078 = n6134 & n22083;
  assign n25079 = ~n25076 & ~n25077;
  assign n25080 = ~n25075 & n25079;
  assign n25081 = ~n25078 & n25080;
  assign n25082 = ~pi17  & ~n25081;
  assign n25083 = pi17  & n25081;
  assign n25084 = ~n25082 & ~n25083;
  assign n25085 = ~n24934 & ~n24937;
  assign n25086 = ~n24918 & ~n24922;
  assign n25087 = n5267 & n20395;
  assign n25088 = n5185 & n20398;
  assign n25089 = n5121 & n20401;
  assign n25090 = n78 & n21305;
  assign n25091 = ~n25088 & ~n25089;
  assign n25092 = ~n25087 & n25091;
  assign n25093 = ~n25090 & n25092;
  assign n25094 = ~pi23  & ~n25093;
  assign n25095 = pi23  & n25093;
  assign n25096 = ~n25094 & ~n25095;
  assign n25097 = ~n24912 & ~n24915;
  assign n25098 = ~n24896 & ~n24899;
  assign n25099 = n4472 & n20413;
  assign n25100 = n4070 & n20416;
  assign n25101 = n3943 & n20419;
  assign n25102 = n3944 & n20928;
  assign n25103 = ~n25100 & ~n25101;
  assign n25104 = ~n25099 & n25103;
  assign n25105 = ~n25102 & n25104;
  assign n25106 = pi29  & n25105;
  assign n25107 = ~pi29  & ~n25105;
  assign n25108 = ~n25106 & ~n25107;
  assign n25109 = ~n24890 & ~n24893;
  assign n25110 = n366 & n1041;
  assign n25111 = n1247 & n25110;
  assign n25112 = ~n91 & ~n553;
  assign n25113 = n927 & n25112;
  assign n25114 = n1077 & n1432;
  assign n25115 = n3085 & n25114;
  assign n25116 = n2445 & n25113;
  assign n25117 = n2454 & n5340;
  assign n25118 = n25116 & n25117;
  assign n25119 = n25111 & n25115;
  assign n25120 = n25118 & n25119;
  assign n25121 = n14539 & n25120;
  assign n25122 = n2922 & n25121;
  assign n25123 = n4178 & n7084;
  assign n25124 = n25122 & n25123;
  assign n25125 = n3896 & n20422;
  assign n25126 = n564 & n20428;
  assign n25127 = n3683 & n20425;
  assign n25128 = n566 & n20801;
  assign n25129 = ~n25126 & ~n25127;
  assign n25130 = ~n25125 & n25129;
  assign n25131 = ~n25128 & n25130;
  assign n25132 = ~n25124 & ~n25131;
  assign n25133 = n25124 & n25131;
  assign n25134 = ~n25132 & ~n25133;
  assign n25135 = ~n25109 & n25134;
  assign n25136 = n25109 & ~n25134;
  assign n25137 = ~n25135 & ~n25136;
  assign n25138 = ~n25108 & n25137;
  assign n25139 = n25108 & ~n25137;
  assign n25140 = ~n25138 & ~n25139;
  assign n25141 = ~n25098 & n25140;
  assign n25142 = n25098 & ~n25140;
  assign n25143 = ~n25141 & ~n25142;
  assign n25144 = n4721 & n20404;
  assign n25145 = n4691 & n20407;
  assign n25146 = n4515 & n20410;
  assign n25147 = n4516 & n20991;
  assign n25148 = ~n25145 & ~n25146;
  assign n25149 = ~n25144 & n25148;
  assign n25150 = ~n25147 & n25149;
  assign n25151 = pi26  & n25150;
  assign n25152 = ~pi26  & ~n25150;
  assign n25153 = ~n25151 & ~n25152;
  assign n25154 = n25143 & ~n25153;
  assign n25155 = ~n25143 & n25153;
  assign n25156 = ~n25154 & ~n25155;
  assign n25157 = ~n25097 & n25156;
  assign n25158 = n25097 & ~n25156;
  assign n25159 = ~n25157 & ~n25158;
  assign n25160 = ~n25096 & n25159;
  assign n25161 = n25096 & ~n25159;
  assign n25162 = ~n25160 & ~n25161;
  assign n25163 = n25086 & ~n25162;
  assign n25164 = ~n25086 & n25162;
  assign n25165 = ~n25163 & ~n25164;
  assign n25166 = n5982 & n20386;
  assign n25167 = n5901 & n20389;
  assign n25168 = n5312 & n20392;
  assign n25169 = n5306 & n21752;
  assign n25170 = ~n25167 & ~n25168;
  assign n25171 = ~n25166 & n25170;
  assign n25172 = ~n25169 & n25171;
  assign n25173 = pi20  & n25172;
  assign n25174 = ~pi20  & ~n25172;
  assign n25175 = ~n25173 & ~n25174;
  assign n25176 = n25165 & ~n25175;
  assign n25177 = ~n25165 & n25175;
  assign n25178 = ~n25176 & ~n25177;
  assign n25179 = ~n25085 & n25178;
  assign n25180 = n25085 & ~n25178;
  assign n25181 = ~n25179 & ~n25180;
  assign n25182 = ~n25084 & n25181;
  assign n25183 = n25084 & ~n25181;
  assign n25184 = ~n25182 & ~n25183;
  assign n25185 = n25074 & ~n25184;
  assign n25186 = ~n25074 & n25184;
  assign n25187 = ~n25185 & ~n25186;
  assign n25188 = n7380 & n20368;
  assign n25189 = n7243 & n20371;
  assign n25190 = n6653 & n20374;
  assign n25191 = n6647 & n22235;
  assign n25192 = ~n25189 & ~n25190;
  assign n25193 = ~n25188 & n25192;
  assign n25194 = ~n25191 & n25193;
  assign n25195 = pi14  & n25194;
  assign n25196 = ~pi14  & ~n25194;
  assign n25197 = ~n25195 & ~n25196;
  assign n25198 = n25187 & ~n25197;
  assign n25199 = ~n25187 & n25197;
  assign n25200 = ~n25198 & ~n25199;
  assign n25201 = ~n25073 & n25200;
  assign n25202 = n25073 & ~n25200;
  assign n25203 = ~n25201 & ~n25202;
  assign n25204 = ~n25072 & n25203;
  assign n25205 = n25072 & ~n25203;
  assign n25206 = ~n25204 & ~n25205;
  assign n25207 = n25062 & ~n25206;
  assign n25208 = ~n25062 & n25206;
  assign n25209 = ~n25207 & ~n25208;
  assign n25210 = n9355 & n23771;
  assign n25211 = n8939 & n23394;
  assign n25212 = n8206 & n20355;
  assign n25213 = n8200 & n23816;
  assign n25214 = ~n25211 & ~n25212;
  assign n25215 = ~n25210 & n25214;
  assign n25216 = ~n25213 & n25215;
  assign n25217 = pi8  & n25216;
  assign n25218 = ~pi8  & ~n25216;
  assign n25219 = ~n25217 & ~n25218;
  assign n25220 = n25209 & ~n25219;
  assign n25221 = ~n25209 & n25219;
  assign n25222 = ~n25220 & ~n25221;
  assign n25223 = ~n25061 & n25222;
  assign n25224 = n25061 & ~n25222;
  assign n25225 = ~n25223 & ~n25224;
  assign n25226 = ~n25060 & n25225;
  assign n25227 = n25060 & ~n25225;
  assign n25228 = ~n25226 & ~n25227;
  assign n25229 = n25050 & ~n25228;
  assign n25230 = ~n25050 & n25228;
  assign n25231 = ~n25229 & ~n25230;
  assign n25232 = ~n25011 & ~n25014;
  assign n25233 = ~n24999 & ~n25001;
  assign n25234 = n562 & ~n25233;
  assign n25235 = ~n562 & n25233;
  assign n25236 = ~n25234 & ~n25235;
  assign n25237 = n3896 & ~n12163;
  assign n25238 = n566 & n13007;
  assign n25239 = n3683 & n12166;
  assign n25240 = n564 & n12172;
  assign n25241 = ~n25237 & ~n25239;
  assign n25242 = ~n25240 & n25241;
  assign n25243 = ~n25238 & n25242;
  assign n25244 = n25236 & ~n25243;
  assign n25245 = ~n25236 & n25243;
  assign n25246 = ~n25244 & ~n25245;
  assign n25247 = n25232 & ~n25246;
  assign n25248 = ~n25232 & n25246;
  assign n25249 = ~n25247 & ~n25248;
  assign n25250 = ~n25017 & ~n25020;
  assign n25251 = ~n25249 & n25250;
  assign n25252 = n25249 & ~n25250;
  assign n25253 = ~n25251 & ~n25252;
  assign n25254 = n11476 & n25253;
  assign n25255 = n11463 & n25022;
  assign n25256 = n10883 & n24779;
  assign n25257 = ~n25028 & ~n25030;
  assign n25258 = n25022 & n25253;
  assign n25259 = ~n25022 & ~n25253;
  assign n25260 = ~n25258 & ~n25259;
  assign n25261 = ~n25257 & n25260;
  assign n25262 = n25257 & ~n25260;
  assign n25263 = ~n25261 & ~n25262;
  assign n25264 = n10884 & n25263;
  assign n25265 = ~n25255 & ~n25256;
  assign n25266 = ~n25254 & n25265;
  assign n25267 = ~n25264 & n25266;
  assign n25268 = pi2  & n25267;
  assign n25269 = ~pi2  & ~n25267;
  assign n25270 = ~n25268 & ~n25269;
  assign n25271 = n25231 & ~n25270;
  assign n25272 = ~n25231 & n25270;
  assign n25273 = ~n25271 & ~n25272;
  assign n25274 = ~n25049 & n25273;
  assign n25275 = n25049 & ~n25273;
  assign n25276 = ~n25274 & ~n25275;
  assign n25277 = n25046 & n25276;
  assign n25278 = ~n25046 & ~n25276;
  assign po3  = ~n25277 & ~n25278;
  assign n25280 = ~n25271 & ~n25274;
  assign n25281 = ~n25226 & ~n25230;
  assign n25282 = n71 & n24779;
  assign n25283 = n10329 & n24529;
  assign n25284 = n9836 & n23765;
  assign n25285 = n9830 & n24789;
  assign n25286 = ~n25283 & ~n25284;
  assign n25287 = ~n25282 & n25286;
  assign n25288 = ~n25285 & n25287;
  assign n25289 = ~pi5  & ~n25288;
  assign n25290 = pi5  & n25288;
  assign n25291 = ~n25289 & ~n25290;
  assign n25292 = ~n25220 & ~n25223;
  assign n25293 = ~n25204 & ~n25208;
  assign n25294 = n8161 & n20355;
  assign n25295 = n7847 & n20358;
  assign n25296 = n7554 & n20361;
  assign n25297 = n7548 & n20562;
  assign n25298 = ~n25295 & ~n25296;
  assign n25299 = ~n25294 & n25298;
  assign n25300 = ~n25297 & n25299;
  assign n25301 = ~pi11  & ~n25300;
  assign n25302 = pi11  & n25300;
  assign n25303 = ~n25301 & ~n25302;
  assign n25304 = ~n25198 & ~n25201;
  assign n25305 = ~n25182 & ~n25186;
  assign n25306 = n6608 & n20374;
  assign n25307 = n6356 & n20377;
  assign n25308 = n6140 & n20380;
  assign n25309 = n6134 & n22263;
  assign n25310 = ~n25307 & ~n25308;
  assign n25311 = ~n25306 & n25310;
  assign n25312 = ~n25309 & n25311;
  assign n25313 = ~pi17  & ~n25312;
  assign n25314 = pi17  & n25312;
  assign n25315 = ~n25313 & ~n25314;
  assign n25316 = ~n25176 & ~n25179;
  assign n25317 = ~n25160 & ~n25164;
  assign n25318 = n5267 & n20392;
  assign n25319 = n5185 & n20395;
  assign n25320 = n5121 & n20398;
  assign n25321 = n78 & n20586;
  assign n25322 = ~n25319 & ~n25320;
  assign n25323 = ~n25318 & n25322;
  assign n25324 = ~n25321 & n25323;
  assign n25325 = ~pi23  & ~n25324;
  assign n25326 = pi23  & n25324;
  assign n25327 = ~n25325 & ~n25326;
  assign n25328 = ~n25154 & ~n25157;
  assign n25329 = ~n25138 & ~n25141;
  assign n25330 = n4472 & n20410;
  assign n25331 = n4070 & n20413;
  assign n25332 = n3943 & n20416;
  assign n25333 = n3944 & n21019;
  assign n25334 = ~n25331 & ~n25332;
  assign n25335 = ~n25330 & n25334;
  assign n25336 = ~n25333 & n25335;
  assign n25337 = pi29  & n25336;
  assign n25338 = ~pi29  & ~n25336;
  assign n25339 = ~n25337 & ~n25338;
  assign n25340 = ~n25132 & ~n25135;
  assign n25341 = ~n126 & ~n315;
  assign n25342 = ~n421 & ~n701;
  assign n25343 = n25341 & n25342;
  assign n25344 = n1014 & n1238;
  assign n25345 = n2390 & n2785;
  assign n25346 = n6440 & n13337;
  assign n25347 = n25345 & n25346;
  assign n25348 = n25343 & n25344;
  assign n25349 = n25347 & n25348;
  assign n25350 = ~n300 & ~n388;
  assign n25351 = ~n541 & n25350;
  assign n25352 = n146 & n201;
  assign n25353 = n885 & n1112;
  assign n25354 = n1344 & n2472;
  assign n25355 = n2787 & n5681;
  assign n25356 = n25354 & n25355;
  assign n25357 = n25352 & n25353;
  assign n25358 = n1084 & n25351;
  assign n25359 = n1966 & n2144;
  assign n25360 = n25358 & n25359;
  assign n25361 = n25356 & n25357;
  assign n25362 = n2732 & n25361;
  assign n25363 = n25349 & n25360;
  assign n25364 = n25362 & n25363;
  assign n25365 = n4342 & n25364;
  assign n25366 = n5022 & n25365;
  assign n25367 = n3896 & n20419;
  assign n25368 = n564 & n20425;
  assign n25369 = n3683 & n20422;
  assign n25370 = n566 & n20786;
  assign n25371 = ~n25368 & ~n25369;
  assign n25372 = ~n25367 & n25371;
  assign n25373 = ~n25370 & n25372;
  assign n25374 = ~n25366 & ~n25373;
  assign n25375 = n25366 & n25373;
  assign n25376 = ~n25374 & ~n25375;
  assign n25377 = ~n25340 & n25376;
  assign n25378 = n25340 & ~n25376;
  assign n25379 = ~n25377 & ~n25378;
  assign n25380 = ~n25339 & n25379;
  assign n25381 = n25339 & ~n25379;
  assign n25382 = ~n25380 & ~n25381;
  assign n25383 = ~n25329 & n25382;
  assign n25384 = n25329 & ~n25382;
  assign n25385 = ~n25383 & ~n25384;
  assign n25386 = n4721 & n20401;
  assign n25387 = n4691 & n20404;
  assign n25388 = n4515 & n20407;
  assign n25389 = n4516 & n21286;
  assign n25390 = ~n25387 & ~n25388;
  assign n25391 = ~n25386 & n25390;
  assign n25392 = ~n25389 & n25391;
  assign n25393 = pi26  & n25392;
  assign n25394 = ~pi26  & ~n25392;
  assign n25395 = ~n25393 & ~n25394;
  assign n25396 = n25385 & ~n25395;
  assign n25397 = ~n25385 & n25395;
  assign n25398 = ~n25396 & ~n25397;
  assign n25399 = ~n25328 & n25398;
  assign n25400 = n25328 & ~n25398;
  assign n25401 = ~n25399 & ~n25400;
  assign n25402 = ~n25327 & n25401;
  assign n25403 = n25327 & ~n25401;
  assign n25404 = ~n25402 & ~n25403;
  assign n25405 = n25317 & ~n25404;
  assign n25406 = ~n25317 & n25404;
  assign n25407 = ~n25405 & ~n25406;
  assign n25408 = n5982 & n20383;
  assign n25409 = n5901 & n20386;
  assign n25410 = n5312 & n20389;
  assign n25411 = n5306 & n21737;
  assign n25412 = ~n25409 & ~n25410;
  assign n25413 = ~n25408 & n25412;
  assign n25414 = ~n25411 & n25413;
  assign n25415 = pi20  & n25414;
  assign n25416 = ~pi20  & ~n25414;
  assign n25417 = ~n25415 & ~n25416;
  assign n25418 = n25407 & ~n25417;
  assign n25419 = ~n25407 & n25417;
  assign n25420 = ~n25418 & ~n25419;
  assign n25421 = ~n25316 & n25420;
  assign n25422 = n25316 & ~n25420;
  assign n25423 = ~n25421 & ~n25422;
  assign n25424 = ~n25315 & n25423;
  assign n25425 = n25315 & ~n25423;
  assign n25426 = ~n25424 & ~n25425;
  assign n25427 = n25305 & ~n25426;
  assign n25428 = ~n25305 & n25426;
  assign n25429 = ~n25427 & ~n25428;
  assign n25430 = n7380 & n20365;
  assign n25431 = n7243 & n20368;
  assign n25432 = n6653 & n20371;
  assign n25433 = n6647 & n22814;
  assign n25434 = ~n25431 & ~n25432;
  assign n25435 = ~n25430 & n25434;
  assign n25436 = ~n25433 & n25435;
  assign n25437 = pi14  & n25436;
  assign n25438 = ~pi14  & ~n25436;
  assign n25439 = ~n25437 & ~n25438;
  assign n25440 = n25429 & ~n25439;
  assign n25441 = ~n25429 & n25439;
  assign n25442 = ~n25440 & ~n25441;
  assign n25443 = ~n25304 & n25442;
  assign n25444 = n25304 & ~n25442;
  assign n25445 = ~n25443 & ~n25444;
  assign n25446 = ~n25303 & n25445;
  assign n25447 = n25303 & ~n25445;
  assign n25448 = ~n25446 & ~n25447;
  assign n25449 = n25293 & ~n25448;
  assign n25450 = ~n25293 & n25448;
  assign n25451 = ~n25449 & ~n25450;
  assign n25452 = n9355 & n23768;
  assign n25453 = n8939 & n23771;
  assign n25454 = n8206 & n23394;
  assign n25455 = n8200 & n23804;
  assign n25456 = ~n25453 & ~n25454;
  assign n25457 = ~n25452 & n25456;
  assign n25458 = ~n25455 & n25457;
  assign n25459 = pi8  & n25458;
  assign n25460 = ~pi8  & ~n25458;
  assign n25461 = ~n25459 & ~n25460;
  assign n25462 = n25451 & ~n25461;
  assign n25463 = ~n25451 & n25461;
  assign n25464 = ~n25462 & ~n25463;
  assign n25465 = ~n25292 & n25464;
  assign n25466 = n25292 & ~n25464;
  assign n25467 = ~n25465 & ~n25466;
  assign n25468 = ~n25291 & n25467;
  assign n25469 = n25291 & ~n25467;
  assign n25470 = ~n25468 & ~n25469;
  assign n25471 = n25281 & ~n25470;
  assign n25472 = ~n25281 & n25470;
  assign n25473 = ~n25471 & ~n25472;
  assign n25474 = n566 & ~n12424;
  assign n25475 = n564 & ~n12165;
  assign n25476 = ~n3683 & ~n3896;
  assign n25477 = ~n25475 & n25476;
  assign n25478 = ~n12163 & ~n25477;
  assign n25479 = ~n25474 & ~n25478;
  assign n25480 = n562 & n25479;
  assign n25481 = ~n562 & ~n25479;
  assign n25482 = ~n25480 & ~n25481;
  assign n25483 = ~n25234 & ~n25244;
  assign n25484 = n25482 & n25483;
  assign n25485 = ~n25482 & ~n25483;
  assign n25486 = ~n25484 & ~n25485;
  assign n25487 = ~n25248 & ~n25252;
  assign n25488 = ~n25486 & n25487;
  assign n25489 = n25486 & ~n25487;
  assign n25490 = ~n25488 & ~n25489;
  assign n25491 = n11476 & n25490;
  assign n25492 = n11463 & n25253;
  assign n25493 = n10883 & n25022;
  assign n25494 = ~n25258 & ~n25261;
  assign n25495 = ~n25253 & ~n25490;
  assign n25496 = n25253 & n25490;
  assign n25497 = ~n25495 & ~n25496;
  assign n25498 = ~n25494 & n25497;
  assign n25499 = n25494 & ~n25497;
  assign n25500 = ~n25498 & ~n25499;
  assign n25501 = n10884 & n25500;
  assign n25502 = ~n25492 & ~n25493;
  assign n25503 = ~n25491 & n25502;
  assign n25504 = ~n25501 & n25503;
  assign n25505 = pi2  & n25504;
  assign n25506 = ~pi2  & ~n25504;
  assign n25507 = ~n25505 & ~n25506;
  assign n25508 = n25473 & ~n25507;
  assign n25509 = ~n25473 & n25507;
  assign n25510 = ~n25508 & ~n25509;
  assign n25511 = ~n25280 & n25510;
  assign n25512 = n25280 & ~n25510;
  assign n25513 = ~n25511 & ~n25512;
  assign n25514 = n25277 & n25513;
  assign n25515 = ~n25277 & ~n25513;
  assign po4  = ~n25514 & ~n25515;
  assign n25517 = ~n25508 & ~n25511;
  assign n25518 = ~n25468 & ~n25472;
  assign n25519 = n71 & n25022;
  assign n25520 = n10329 & n24779;
  assign n25521 = n9836 & n24529;
  assign n25522 = n9830 & n25032;
  assign n25523 = ~n25520 & ~n25521;
  assign n25524 = ~n25519 & n25523;
  assign n25525 = ~n25522 & n25524;
  assign n25526 = ~pi5  & ~n25525;
  assign n25527 = pi5  & n25525;
  assign n25528 = ~n25526 & ~n25527;
  assign n25529 = ~n25462 & ~n25465;
  assign n25530 = ~n25446 & ~n25450;
  assign n25531 = n8161 & n23394;
  assign n25532 = n7847 & n20355;
  assign n25533 = n7554 & n20358;
  assign n25534 = n7548 & n23404;
  assign n25535 = ~n25532 & ~n25533;
  assign n25536 = ~n25531 & n25535;
  assign n25537 = ~n25534 & n25536;
  assign n25538 = ~pi11  & ~n25537;
  assign n25539 = pi11  & n25537;
  assign n25540 = ~n25538 & ~n25539;
  assign n25541 = ~n25440 & ~n25443;
  assign n25542 = ~n25424 & ~n25428;
  assign n25543 = n6608 & n20371;
  assign n25544 = n6356 & n20374;
  assign n25545 = n6140 & n20377;
  assign n25546 = n6134 & n22250;
  assign n25547 = ~n25544 & ~n25545;
  assign n25548 = ~n25543 & n25547;
  assign n25549 = ~n25546 & n25548;
  assign n25550 = ~pi17  & ~n25549;
  assign n25551 = pi17  & n25549;
  assign n25552 = ~n25550 & ~n25551;
  assign n25553 = ~n25418 & ~n25421;
  assign n25554 = ~n25402 & ~n25406;
  assign n25555 = n5267 & n20389;
  assign n25556 = n5185 & n20392;
  assign n25557 = n5121 & n20395;
  assign n25558 = n78 & n21716;
  assign n25559 = ~n25556 & ~n25557;
  assign n25560 = ~n25555 & n25559;
  assign n25561 = ~n25558 & n25560;
  assign n25562 = ~pi23  & ~n25561;
  assign n25563 = pi23  & n25561;
  assign n25564 = ~n25562 & ~n25563;
  assign n25565 = ~n25396 & ~n25399;
  assign n25566 = ~n25380 & ~n25383;
  assign n25567 = n4472 & n20407;
  assign n25568 = n4070 & n20410;
  assign n25569 = n3943 & n20413;
  assign n25570 = n3944 & n21004;
  assign n25571 = ~n25568 & ~n25569;
  assign n25572 = ~n25567 & n25571;
  assign n25573 = ~n25570 & n25572;
  assign n25574 = pi29  & n25573;
  assign n25575 = ~pi29  & ~n25573;
  assign n25576 = ~n25574 & ~n25575;
  assign n25577 = ~n25374 & ~n25377;
  assign n25578 = ~n195 & ~n216;
  assign n25579 = ~n405 & ~n470;
  assign n25580 = ~n572 & ~n648;
  assign n25581 = ~n667 & n25580;
  assign n25582 = n25578 & n25579;
  assign n25583 = n523 & n1054;
  assign n25584 = n1594 & n2374;
  assign n25585 = n5574 & n25584;
  assign n25586 = n25582 & n25583;
  assign n25587 = n25581 & n25586;
  assign n25588 = n1081 & n25585;
  assign n25589 = n4160 & n25588;
  assign n25590 = n4110 & n25587;
  assign n25591 = n25589 & n25590;
  assign n25592 = n5786 & n25591;
  assign n25593 = n14752 & n25592;
  assign n25594 = n3896 & n20416;
  assign n25595 = n564 & n20422;
  assign n25596 = n3683 & n20419;
  assign n25597 = n566 & n20771;
  assign n25598 = ~n25595 & ~n25596;
  assign n25599 = ~n25594 & n25598;
  assign n25600 = ~n25597 & n25599;
  assign n25601 = ~n25593 & ~n25600;
  assign n25602 = n25593 & n25600;
  assign n25603 = ~n25601 & ~n25602;
  assign n25604 = ~n25577 & n25603;
  assign n25605 = n25577 & ~n25603;
  assign n25606 = ~n25604 & ~n25605;
  assign n25607 = ~n25576 & n25606;
  assign n25608 = n25576 & ~n25606;
  assign n25609 = ~n25607 & ~n25608;
  assign n25610 = ~n25566 & n25609;
  assign n25611 = n25566 & ~n25609;
  assign n25612 = ~n25610 & ~n25611;
  assign n25613 = n4721 & n20398;
  assign n25614 = n4691 & n20401;
  assign n25615 = n4515 & n20404;
  assign n25616 = n4516 & n21322;
  assign n25617 = ~n25614 & ~n25615;
  assign n25618 = ~n25613 & n25617;
  assign n25619 = ~n25616 & n25618;
  assign n25620 = pi26  & n25619;
  assign n25621 = ~pi26  & ~n25619;
  assign n25622 = ~n25620 & ~n25621;
  assign n25623 = n25612 & ~n25622;
  assign n25624 = ~n25612 & n25622;
  assign n25625 = ~n25623 & ~n25624;
  assign n25626 = ~n25565 & n25625;
  assign n25627 = n25565 & ~n25625;
  assign n25628 = ~n25626 & ~n25627;
  assign n25629 = ~n25564 & n25628;
  assign n25630 = n25564 & ~n25628;
  assign n25631 = ~n25629 & ~n25630;
  assign n25632 = n25554 & ~n25631;
  assign n25633 = ~n25554 & n25631;
  assign n25634 = ~n25632 & ~n25633;
  assign n25635 = n5982 & n20380;
  assign n25636 = n5901 & n20383;
  assign n25637 = n5312 & n20386;
  assign n25638 = n5306 & n20574;
  assign n25639 = ~n25636 & ~n25637;
  assign n25640 = ~n25635 & n25639;
  assign n25641 = ~n25638 & n25640;
  assign n25642 = pi20  & n25641;
  assign n25643 = ~pi20  & ~n25641;
  assign n25644 = ~n25642 & ~n25643;
  assign n25645 = n25634 & ~n25644;
  assign n25646 = ~n25634 & n25644;
  assign n25647 = ~n25645 & ~n25646;
  assign n25648 = ~n25553 & n25647;
  assign n25649 = n25553 & ~n25647;
  assign n25650 = ~n25648 & ~n25649;
  assign n25651 = ~n25552 & n25650;
  assign n25652 = n25552 & ~n25650;
  assign n25653 = ~n25651 & ~n25652;
  assign n25654 = n25542 & ~n25653;
  assign n25655 = ~n25542 & n25653;
  assign n25656 = ~n25654 & ~n25655;
  assign n25657 = n7380 & n20361;
  assign n25658 = n7243 & n20365;
  assign n25659 = n6653 & n20368;
  assign n25660 = n6647 & n22848;
  assign n25661 = ~n25658 & ~n25659;
  assign n25662 = ~n25657 & n25661;
  assign n25663 = ~n25660 & n25662;
  assign n25664 = pi14  & n25663;
  assign n25665 = ~pi14  & ~n25663;
  assign n25666 = ~n25664 & ~n25665;
  assign n25667 = n25656 & ~n25666;
  assign n25668 = ~n25656 & n25666;
  assign n25669 = ~n25667 & ~n25668;
  assign n25670 = ~n25541 & n25669;
  assign n25671 = n25541 & ~n25669;
  assign n25672 = ~n25670 & ~n25671;
  assign n25673 = ~n25540 & n25672;
  assign n25674 = n25540 & ~n25672;
  assign n25675 = ~n25673 & ~n25674;
  assign n25676 = n25530 & ~n25675;
  assign n25677 = ~n25530 & n25675;
  assign n25678 = ~n25676 & ~n25677;
  assign n25679 = n9355 & n23765;
  assign n25680 = n8939 & n23768;
  assign n25681 = n8206 & n23771;
  assign n25682 = n8200 & n23789;
  assign n25683 = ~n25680 & ~n25681;
  assign n25684 = ~n25679 & n25683;
  assign n25685 = ~n25682 & n25684;
  assign n25686 = pi8  & n25685;
  assign n25687 = ~pi8  & ~n25685;
  assign n25688 = ~n25686 & ~n25687;
  assign n25689 = n25678 & ~n25688;
  assign n25690 = ~n25678 & n25688;
  assign n25691 = ~n25689 & ~n25690;
  assign n25692 = ~n25529 & n25691;
  assign n25693 = n25529 & ~n25691;
  assign n25694 = ~n25692 & ~n25693;
  assign n25695 = ~n25528 & n25694;
  assign n25696 = n25528 & ~n25694;
  assign n25697 = ~n25695 & ~n25696;
  assign n25698 = n25518 & ~n25697;
  assign n25699 = ~n25518 & n25697;
  assign n25700 = ~n25698 & ~n25699;
  assign n25701 = ~n25485 & ~n25489;
  assign n25702 = ~pi31  & n105;
  assign n25703 = ~n12163 & ~n25702;
  assign n25704 = n25480 & ~n25703;
  assign n25705 = ~n25480 & n25703;
  assign n25706 = ~n25704 & ~n25705;
  assign n25707 = n25701 & n25706;
  assign n25708 = ~n25701 & ~n25706;
  assign n25709 = ~n25707 & ~n25708;
  assign n25710 = n11476 & n25709;
  assign n25711 = n11463 & n25490;
  assign n25712 = n10883 & n25253;
  assign n25713 = ~n25496 & ~n25498;
  assign n25714 = n25490 & n25709;
  assign n25715 = ~n25490 & ~n25709;
  assign n25716 = ~n25714 & ~n25715;
  assign n25717 = ~n25713 & n25716;
  assign n25718 = n25713 & ~n25716;
  assign n25719 = ~n25717 & ~n25718;
  assign n25720 = n10884 & n25719;
  assign n25721 = ~n25711 & ~n25712;
  assign n25722 = ~n25710 & n25721;
  assign n25723 = ~n25720 & n25722;
  assign n25724 = pi2  & n25723;
  assign n25725 = ~pi2  & ~n25723;
  assign n25726 = ~n25724 & ~n25725;
  assign n25727 = n25700 & ~n25726;
  assign n25728 = ~n25700 & n25726;
  assign n25729 = ~n25727 & ~n25728;
  assign n25730 = ~n25517 & n25729;
  assign n25731 = n25517 & ~n25729;
  assign n25732 = ~n25730 & ~n25731;
  assign n25733 = n25514 & n25732;
  assign n25734 = ~n25514 & ~n25732;
  assign po5  = ~n25733 & ~n25734;
  assign n25736 = ~n25695 & ~n25699;
  assign n25737 = n71 & n25253;
  assign n25738 = n10329 & n25022;
  assign n25739 = n9836 & n24779;
  assign n25740 = n9830 & n25263;
  assign n25741 = ~n25738 & ~n25739;
  assign n25742 = ~n25737 & n25741;
  assign n25743 = ~n25740 & n25742;
  assign n25744 = ~pi5  & ~n25743;
  assign n25745 = pi5  & n25743;
  assign n25746 = ~n25744 & ~n25745;
  assign n25747 = ~n25689 & ~n25692;
  assign n25748 = ~n25673 & ~n25677;
  assign n25749 = n8161 & n23771;
  assign n25750 = n7847 & n23394;
  assign n25751 = n7554 & n20355;
  assign n25752 = n7548 & n23816;
  assign n25753 = ~n25750 & ~n25751;
  assign n25754 = ~n25749 & n25753;
  assign n25755 = ~n25752 & n25754;
  assign n25756 = ~pi11  & ~n25755;
  assign n25757 = pi11  & n25755;
  assign n25758 = ~n25756 & ~n25757;
  assign n25759 = ~n25667 & ~n25670;
  assign n25760 = ~n25651 & ~n25655;
  assign n25761 = n6608 & n20368;
  assign n25762 = n6356 & n20371;
  assign n25763 = n6140 & n20374;
  assign n25764 = n6134 & n22235;
  assign n25765 = ~n25762 & ~n25763;
  assign n25766 = ~n25761 & n25765;
  assign n25767 = ~n25764 & n25766;
  assign n25768 = ~pi17  & ~n25767;
  assign n25769 = pi17  & n25767;
  assign n25770 = ~n25768 & ~n25769;
  assign n25771 = ~n25645 & ~n25648;
  assign n25772 = ~n25629 & ~n25633;
  assign n25773 = n5267 & n20386;
  assign n25774 = n5185 & n20389;
  assign n25775 = n5121 & n20392;
  assign n25776 = n78 & n21752;
  assign n25777 = ~n25774 & ~n25775;
  assign n25778 = ~n25773 & n25777;
  assign n25779 = ~n25776 & n25778;
  assign n25780 = ~pi23  & ~n25779;
  assign n25781 = pi23  & n25779;
  assign n25782 = ~n25780 & ~n25781;
  assign n25783 = ~n25623 & ~n25626;
  assign n25784 = ~n25607 & ~n25610;
  assign n25785 = n4472 & n20404;
  assign n25786 = n4070 & n20407;
  assign n25787 = n3943 & n20410;
  assign n25788 = n3944 & n20991;
  assign n25789 = ~n25786 & ~n25787;
  assign n25790 = ~n25785 & n25789;
  assign n25791 = ~n25788 & n25790;
  assign n25792 = pi29  & n25791;
  assign n25793 = ~pi29  & ~n25791;
  assign n25794 = ~n25792 & ~n25793;
  assign n25795 = ~n25601 & ~n25604;
  assign n25796 = ~n250 & ~n553;
  assign n25797 = n850 & n25796;
  assign n25798 = n2300 & n2493;
  assign n25799 = n5529 & n25798;
  assign n25800 = n25797 & n25799;
  assign n25801 = ~n279 & ~n311;
  assign n25802 = ~n389 & ~n465;
  assign n25803 = ~n467 & ~n522;
  assign n25804 = n25802 & n25803;
  assign n25805 = n201 & n25801;
  assign n25806 = n885 & n969;
  assign n25807 = n1117 & n1357;
  assign n25808 = n1394 & n1431;
  assign n25809 = n2050 & n25808;
  assign n25810 = n25806 & n25807;
  assign n25811 = n25804 & n25805;
  assign n25812 = n25810 & n25811;
  assign n25813 = n25111 & n25809;
  assign n25814 = n25812 & n25813;
  assign n25815 = n13495 & n25800;
  assign n25816 = n25814 & n25815;
  assign n25817 = n3119 & n5561;
  assign n25818 = n13915 & n25817;
  assign n25819 = n25816 & n25818;
  assign n25820 = n3896 & n20413;
  assign n25821 = n564 & n20419;
  assign n25822 = n3683 & n20416;
  assign n25823 = n566 & n20928;
  assign n25824 = ~n25821 & ~n25822;
  assign n25825 = ~n25820 & n25824;
  assign n25826 = ~n25823 & n25825;
  assign n25827 = ~n25819 & ~n25826;
  assign n25828 = n25819 & n25826;
  assign n25829 = ~n25827 & ~n25828;
  assign n25830 = ~n25795 & n25829;
  assign n25831 = n25795 & ~n25829;
  assign n25832 = ~n25830 & ~n25831;
  assign n25833 = ~n25794 & n25832;
  assign n25834 = n25794 & ~n25832;
  assign n25835 = ~n25833 & ~n25834;
  assign n25836 = ~n25784 & n25835;
  assign n25837 = n25784 & ~n25835;
  assign n25838 = ~n25836 & ~n25837;
  assign n25839 = n4721 & n20395;
  assign n25840 = n4691 & n20398;
  assign n25841 = n4515 & n20401;
  assign n25842 = n4516 & n21305;
  assign n25843 = ~n25840 & ~n25841;
  assign n25844 = ~n25839 & n25843;
  assign n25845 = ~n25842 & n25844;
  assign n25846 = pi26  & n25845;
  assign n25847 = ~pi26  & ~n25845;
  assign n25848 = ~n25846 & ~n25847;
  assign n25849 = n25838 & ~n25848;
  assign n25850 = ~n25838 & n25848;
  assign n25851 = ~n25849 & ~n25850;
  assign n25852 = ~n25783 & n25851;
  assign n25853 = n25783 & ~n25851;
  assign n25854 = ~n25852 & ~n25853;
  assign n25855 = ~n25782 & n25854;
  assign n25856 = n25782 & ~n25854;
  assign n25857 = ~n25855 & ~n25856;
  assign n25858 = n25772 & ~n25857;
  assign n25859 = ~n25772 & n25857;
  assign n25860 = ~n25858 & ~n25859;
  assign n25861 = n5982 & n20377;
  assign n25862 = n5901 & n20380;
  assign n25863 = n5312 & n20383;
  assign n25864 = n5306 & n22083;
  assign n25865 = ~n25862 & ~n25863;
  assign n25866 = ~n25861 & n25865;
  assign n25867 = ~n25864 & n25866;
  assign n25868 = pi20  & n25867;
  assign n25869 = ~pi20  & ~n25867;
  assign n25870 = ~n25868 & ~n25869;
  assign n25871 = n25860 & ~n25870;
  assign n25872 = ~n25860 & n25870;
  assign n25873 = ~n25871 & ~n25872;
  assign n25874 = ~n25771 & n25873;
  assign n25875 = n25771 & ~n25873;
  assign n25876 = ~n25874 & ~n25875;
  assign n25877 = ~n25770 & n25876;
  assign n25878 = n25770 & ~n25876;
  assign n25879 = ~n25877 & ~n25878;
  assign n25880 = n25760 & ~n25879;
  assign n25881 = ~n25760 & n25879;
  assign n25882 = ~n25880 & ~n25881;
  assign n25883 = n7380 & n20358;
  assign n25884 = n7243 & n20361;
  assign n25885 = n6653 & n20365;
  assign n25886 = n6647 & n22833;
  assign n25887 = ~n25884 & ~n25885;
  assign n25888 = ~n25883 & n25887;
  assign n25889 = ~n25886 & n25888;
  assign n25890 = pi14  & n25889;
  assign n25891 = ~pi14  & ~n25889;
  assign n25892 = ~n25890 & ~n25891;
  assign n25893 = n25882 & ~n25892;
  assign n25894 = ~n25882 & n25892;
  assign n25895 = ~n25893 & ~n25894;
  assign n25896 = ~n25759 & n25895;
  assign n25897 = n25759 & ~n25895;
  assign n25898 = ~n25896 & ~n25897;
  assign n25899 = ~n25758 & n25898;
  assign n25900 = n25758 & ~n25898;
  assign n25901 = ~n25899 & ~n25900;
  assign n25902 = n25748 & ~n25901;
  assign n25903 = ~n25748 & n25901;
  assign n25904 = ~n25902 & ~n25903;
  assign n25905 = n9355 & n24529;
  assign n25906 = n8939 & n23765;
  assign n25907 = n8206 & n23768;
  assign n25908 = n8200 & n24539;
  assign n25909 = ~n25906 & ~n25907;
  assign n25910 = ~n25905 & n25909;
  assign n25911 = ~n25908 & n25910;
  assign n25912 = pi8  & n25911;
  assign n25913 = ~pi8  & ~n25911;
  assign n25914 = ~n25912 & ~n25913;
  assign n25915 = n25904 & ~n25914;
  assign n25916 = ~n25904 & n25914;
  assign n25917 = ~n25915 & ~n25916;
  assign n25918 = ~n25747 & n25917;
  assign n25919 = n25747 & ~n25917;
  assign n25920 = ~n25918 & ~n25919;
  assign n25921 = ~n25746 & n25920;
  assign n25922 = n25746 & ~n25920;
  assign n25923 = ~n25921 & ~n25922;
  assign n25924 = ~n19063 & n25709;
  assign n25925 = ~n25714 & ~n25717;
  assign n25926 = n10884 & ~n25925;
  assign n25927 = n10883 & n25490;
  assign n25928 = ~n25924 & ~n25927;
  assign n25929 = ~n25926 & n25928;
  assign n25930 = pi2  & n25929;
  assign n25931 = ~pi2  & ~n25929;
  assign n25932 = ~n25930 & ~n25931;
  assign n25933 = n25923 & ~n25932;
  assign n25934 = ~n25923 & n25932;
  assign n25935 = ~n25933 & ~n25934;
  assign n25936 = n25736 & ~n25935;
  assign n25937 = ~n25736 & n25935;
  assign n25938 = ~n25936 & ~n25937;
  assign n25939 = ~n25727 & ~n25730;
  assign n25940 = ~n25938 & n25939;
  assign n25941 = n25938 & ~n25939;
  assign n25942 = ~n25940 & ~n25941;
  assign n25943 = n25733 & n25942;
  assign n25944 = ~n25733 & ~n25942;
  assign po6  = ~n25943 & ~n25944;
  assign n25946 = ~n25921 & ~n25933;
  assign n25947 = ~n25915 & ~n25918;
  assign n25948 = ~n25899 & ~n25903;
  assign n25949 = ~n25893 & ~n25896;
  assign n25950 = ~n25877 & ~n25881;
  assign n25951 = ~n25871 & ~n25874;
  assign n25952 = ~n25855 & ~n25859;
  assign n25953 = ~n25833 & ~n25836;
  assign n25954 = ~n25827 & ~n25830;
  assign n25955 = ~n307 & ~n379;
  assign n25956 = ~n494 & ~n666;
  assign n25957 = n25955 & n25956;
  assign n25958 = n624 & n1015;
  assign n25959 = n3079 & n13338;
  assign n25960 = n25958 & n25959;
  assign n25961 = n2806 & n25957;
  assign n25962 = n12649 & n13311;
  assign n25963 = n25961 & n25962;
  assign n25964 = n7055 & n25960;
  assign n25965 = n25963 & n25964;
  assign n25966 = n260 & n2638;
  assign n25967 = n12470 & n25966;
  assign n25968 = n25965 & n25967;
  assign n25969 = n3168 & n25968;
  assign n25970 = n881 & n25969;
  assign n25971 = pi2  & ~n25709;
  assign n25972 = n13900 & n25709;
  assign n25973 = ~n25971 & ~n25972;
  assign n25974 = ~n25970 & ~n25973;
  assign n25975 = n25970 & n25973;
  assign n25976 = ~n25974 & ~n25975;
  assign n25977 = n3896 & n20410;
  assign n25978 = n3683 & n20413;
  assign n25979 = n564 & n20416;
  assign n25980 = n566 & n21019;
  assign n25981 = ~n25978 & ~n25979;
  assign n25982 = ~n25977 & n25981;
  assign n25983 = ~n25980 & n25982;
  assign n25984 = ~n25976 & n25983;
  assign n25985 = n25976 & ~n25983;
  assign n25986 = ~n25984 & ~n25985;
  assign n25987 = n25954 & ~n25986;
  assign n25988 = ~n25954 & n25986;
  assign n25989 = ~n25987 & ~n25988;
  assign n25990 = n4472 & n20401;
  assign n25991 = n4070 & n20404;
  assign n25992 = n3943 & n20407;
  assign n25993 = n3944 & n21286;
  assign n25994 = ~n25991 & ~n25992;
  assign n25995 = ~n25990 & n25994;
  assign n25996 = ~n25993 & n25995;
  assign n25997 = pi29  & n25996;
  assign n25998 = ~pi29  & ~n25996;
  assign n25999 = ~n25997 & ~n25998;
  assign n26000 = n25989 & ~n25999;
  assign n26001 = ~n25989 & n25999;
  assign n26002 = ~n26000 & ~n26001;
  assign n26003 = ~n25953 & n26002;
  assign n26004 = n25953 & ~n26002;
  assign n26005 = ~n26003 & ~n26004;
  assign n26006 = n4721 & n20392;
  assign n26007 = n4691 & n20395;
  assign n26008 = n4515 & n20398;
  assign n26009 = n4516 & n20586;
  assign n26010 = ~n26007 & ~n26008;
  assign n26011 = ~n26006 & n26010;
  assign n26012 = ~n26009 & n26011;
  assign n26013 = pi26  & n26012;
  assign n26014 = ~pi26  & ~n26012;
  assign n26015 = ~n26013 & ~n26014;
  assign n26016 = n26005 & n26015;
  assign n26017 = ~n26005 & ~n26015;
  assign n26018 = ~n26016 & ~n26017;
  assign n26019 = ~n25849 & ~n25852;
  assign n26020 = n26018 & n26019;
  assign n26021 = ~n26018 & ~n26019;
  assign n26022 = ~n26020 & ~n26021;
  assign n26023 = n5267 & n20383;
  assign n26024 = n5185 & n20386;
  assign n26025 = n5121 & n20389;
  assign n26026 = n78 & n21737;
  assign n26027 = ~n26024 & ~n26025;
  assign n26028 = ~n26023 & n26027;
  assign n26029 = ~n26026 & n26028;
  assign n26030 = pi23  & n26029;
  assign n26031 = ~pi23  & ~n26029;
  assign n26032 = ~n26030 & ~n26031;
  assign n26033 = n26022 & ~n26032;
  assign n26034 = ~n26022 & n26032;
  assign n26035 = ~n26033 & ~n26034;
  assign n26036 = n25952 & ~n26035;
  assign n26037 = ~n25952 & n26035;
  assign n26038 = ~n26036 & ~n26037;
  assign n26039 = n5982 & n20374;
  assign n26040 = n5901 & n20377;
  assign n26041 = n5312 & n20380;
  assign n26042 = n5306 & n22263;
  assign n26043 = ~n26040 & ~n26041;
  assign n26044 = ~n26039 & n26043;
  assign n26045 = ~n26042 & n26044;
  assign n26046 = pi20  & n26045;
  assign n26047 = ~pi20  & ~n26045;
  assign n26048 = ~n26046 & ~n26047;
  assign n26049 = n26038 & ~n26048;
  assign n26050 = ~n26038 & n26048;
  assign n26051 = ~n26049 & ~n26050;
  assign n26052 = n25951 & ~n26051;
  assign n26053 = ~n25951 & n26051;
  assign n26054 = ~n26052 & ~n26053;
  assign n26055 = n6608 & n20365;
  assign n26056 = n6356 & n20368;
  assign n26057 = n6140 & n20371;
  assign n26058 = n6134 & n22814;
  assign n26059 = ~n26056 & ~n26057;
  assign n26060 = ~n26055 & n26059;
  assign n26061 = ~n26058 & n26060;
  assign n26062 = pi17  & n26061;
  assign n26063 = ~pi17  & ~n26061;
  assign n26064 = ~n26062 & ~n26063;
  assign n26065 = n26054 & ~n26064;
  assign n26066 = ~n26054 & n26064;
  assign n26067 = ~n26065 & ~n26066;
  assign n26068 = n25950 & ~n26067;
  assign n26069 = ~n25950 & n26067;
  assign n26070 = ~n26068 & ~n26069;
  assign n26071 = n7380 & n20355;
  assign n26072 = n7243 & n20358;
  assign n26073 = n6653 & n20361;
  assign n26074 = n6647 & n20562;
  assign n26075 = ~n26072 & ~n26073;
  assign n26076 = ~n26071 & n26075;
  assign n26077 = ~n26074 & n26076;
  assign n26078 = pi14  & n26077;
  assign n26079 = ~pi14  & ~n26077;
  assign n26080 = ~n26078 & ~n26079;
  assign n26081 = n26070 & ~n26080;
  assign n26082 = ~n26070 & n26080;
  assign n26083 = ~n26081 & ~n26082;
  assign n26084 = n25949 & ~n26083;
  assign n26085 = ~n25949 & n26083;
  assign n26086 = ~n26084 & ~n26085;
  assign n26087 = n8161 & n23768;
  assign n26088 = n7847 & n23771;
  assign n26089 = n7554 & n23394;
  assign n26090 = n7548 & n23804;
  assign n26091 = ~n26088 & ~n26089;
  assign n26092 = ~n26087 & n26091;
  assign n26093 = ~n26090 & n26092;
  assign n26094 = pi11  & n26093;
  assign n26095 = ~pi11  & ~n26093;
  assign n26096 = ~n26094 & ~n26095;
  assign n26097 = n26086 & ~n26096;
  assign n26098 = ~n26086 & n26096;
  assign n26099 = ~n26097 & ~n26098;
  assign n26100 = n25948 & ~n26099;
  assign n26101 = ~n25948 & n26099;
  assign n26102 = ~n26100 & ~n26101;
  assign n26103 = n9355 & n24779;
  assign n26104 = n8939 & n24529;
  assign n26105 = n8206 & n23765;
  assign n26106 = n8200 & n24789;
  assign n26107 = ~n26104 & ~n26105;
  assign n26108 = ~n26103 & n26107;
  assign n26109 = ~n26106 & n26108;
  assign n26110 = pi8  & n26109;
  assign n26111 = ~pi8  & ~n26109;
  assign n26112 = ~n26110 & ~n26111;
  assign n26113 = n26102 & ~n26112;
  assign n26114 = ~n26102 & n26112;
  assign n26115 = ~n26113 & ~n26114;
  assign n26116 = n25947 & ~n26115;
  assign n26117 = ~n25947 & n26115;
  assign n26118 = ~n26116 & ~n26117;
  assign n26119 = n71 & n25490;
  assign n26120 = n10329 & n25253;
  assign n26121 = n9836 & n25022;
  assign n26122 = n9830 & n25500;
  assign n26123 = ~n26120 & ~n26121;
  assign n26124 = ~n26119 & n26123;
  assign n26125 = ~n26122 & n26124;
  assign n26126 = pi5  & n26125;
  assign n26127 = ~pi5  & ~n26125;
  assign n26128 = ~n26126 & ~n26127;
  assign n26129 = n26118 & ~n26128;
  assign n26130 = ~n26118 & n26128;
  assign n26131 = ~n26129 & ~n26130;
  assign n26132 = n25946 & ~n26131;
  assign n26133 = ~n25946 & n26131;
  assign n26134 = ~n26132 & ~n26133;
  assign n26135 = ~n25937 & ~n25941;
  assign n26136 = ~n26134 & n26135;
  assign n26137 = n26134 & ~n26135;
  assign n26138 = ~n26136 & ~n26137;
  assign n26139 = n25943 & n26138;
  assign n26140 = ~n25943 & ~n26138;
  assign po7  = ~n26139 & ~n26140;
  assign n26142 = ~n26117 & ~n26129;
  assign n26143 = ~n26101 & ~n26113;
  assign n26144 = ~n26085 & ~n26097;
  assign n26145 = ~n26069 & ~n26081;
  assign n26146 = ~n26053 & ~n26065;
  assign n26147 = ~n26037 & ~n26049;
  assign n26148 = ~n26021 & ~n26033;
  assign n26149 = n4721 & n20389;
  assign n26150 = n4691 & n20392;
  assign n26151 = n4515 & n20395;
  assign n26152 = n4516 & n21716;
  assign n26153 = ~n26150 & ~n26151;
  assign n26154 = ~n26149 & n26153;
  assign n26155 = ~n26152 & n26154;
  assign n26156 = pi26  & n26155;
  assign n26157 = ~pi26  & ~n26155;
  assign n26158 = ~n26156 & ~n26157;
  assign n26159 = ~n25988 & ~n26000;
  assign n26160 = ~n285 & ~n467;
  assign n26161 = ~n646 & n26160;
  assign n26162 = n471 & n26161;
  assign n26163 = n14839 & n26162;
  assign n26164 = ~n134 & ~n310;
  assign n26165 = ~n364 & ~n463;
  assign n26166 = n26164 & n26165;
  assign n26167 = n337 & n403;
  assign n26168 = n600 & n1355;
  assign n26169 = n1508 & n1754;
  assign n26170 = n2193 & n2599;
  assign n26171 = n3085 & n4156;
  assign n26172 = n26170 & n26171;
  assign n26173 = n26168 & n26169;
  assign n26174 = n26166 & n26167;
  assign n26175 = n22128 & n26174;
  assign n26176 = n26172 & n26173;
  assign n26177 = n26175 & n26176;
  assign n26178 = n2059 & n26163;
  assign n26179 = n26177 & n26178;
  assign n26180 = n2851 & n26179;
  assign n26181 = n14816 & n26180;
  assign n26182 = ~n25973 & ~n26181;
  assign n26183 = n25973 & n26181;
  assign n26184 = ~n26182 & ~n26183;
  assign n26185 = ~n25975 & ~n25983;
  assign n26186 = ~n25974 & ~n26185;
  assign n26187 = n26184 & ~n26186;
  assign n26188 = ~n26184 & n26186;
  assign n26189 = ~n26187 & ~n26188;
  assign n26190 = n3896 & n20407;
  assign n26191 = n3683 & n20410;
  assign n26192 = n564 & n20413;
  assign n26193 = n566 & n21004;
  assign n26194 = ~n26191 & ~n26192;
  assign n26195 = ~n26190 & n26194;
  assign n26196 = ~n26193 & n26195;
  assign n26197 = n26189 & ~n26196;
  assign n26198 = ~n26189 & n26196;
  assign n26199 = ~n26197 & ~n26198;
  assign n26200 = n26159 & ~n26199;
  assign n26201 = ~n26159 & n26199;
  assign n26202 = ~n26200 & ~n26201;
  assign n26203 = n4472 & n20398;
  assign n26204 = n4070 & n20401;
  assign n26205 = n3943 & n20404;
  assign n26206 = n3944 & n21322;
  assign n26207 = ~n26204 & ~n26205;
  assign n26208 = ~n26203 & n26207;
  assign n26209 = ~n26206 & n26208;
  assign n26210 = pi29  & n26209;
  assign n26211 = ~pi29  & ~n26209;
  assign n26212 = ~n26210 & ~n26211;
  assign n26213 = n26202 & ~n26212;
  assign n26214 = ~n26202 & n26212;
  assign n26215 = ~n26213 & ~n26214;
  assign n26216 = ~n26158 & n26215;
  assign n26217 = n26158 & ~n26215;
  assign n26218 = ~n26216 & ~n26217;
  assign n26219 = ~n26004 & ~n26016;
  assign n26220 = ~n26218 & ~n26219;
  assign n26221 = n26218 & n26219;
  assign n26222 = ~n26220 & ~n26221;
  assign n26223 = n5267 & n20380;
  assign n26224 = n5185 & n20383;
  assign n26225 = n5121 & n20386;
  assign n26226 = n78 & n20574;
  assign n26227 = ~n26224 & ~n26225;
  assign n26228 = ~n26223 & n26227;
  assign n26229 = ~n26226 & n26228;
  assign n26230 = pi23  & n26229;
  assign n26231 = ~pi23  & ~n26229;
  assign n26232 = ~n26230 & ~n26231;
  assign n26233 = n26222 & ~n26232;
  assign n26234 = ~n26222 & n26232;
  assign n26235 = ~n26233 & ~n26234;
  assign n26236 = n26148 & ~n26235;
  assign n26237 = ~n26148 & n26235;
  assign n26238 = ~n26236 & ~n26237;
  assign n26239 = n5982 & n20371;
  assign n26240 = n5901 & n20374;
  assign n26241 = n5312 & n20377;
  assign n26242 = n5306 & n22250;
  assign n26243 = ~n26240 & ~n26241;
  assign n26244 = ~n26239 & n26243;
  assign n26245 = ~n26242 & n26244;
  assign n26246 = pi20  & n26245;
  assign n26247 = ~pi20  & ~n26245;
  assign n26248 = ~n26246 & ~n26247;
  assign n26249 = n26238 & ~n26248;
  assign n26250 = ~n26238 & n26248;
  assign n26251 = ~n26249 & ~n26250;
  assign n26252 = n26147 & ~n26251;
  assign n26253 = ~n26147 & n26251;
  assign n26254 = ~n26252 & ~n26253;
  assign n26255 = n6608 & n20361;
  assign n26256 = n6356 & n20365;
  assign n26257 = n6140 & n20368;
  assign n26258 = n6134 & n22848;
  assign n26259 = ~n26256 & ~n26257;
  assign n26260 = ~n26255 & n26259;
  assign n26261 = ~n26258 & n26260;
  assign n26262 = pi17  & n26261;
  assign n26263 = ~pi17  & ~n26261;
  assign n26264 = ~n26262 & ~n26263;
  assign n26265 = n26254 & ~n26264;
  assign n26266 = ~n26254 & n26264;
  assign n26267 = ~n26265 & ~n26266;
  assign n26268 = n26146 & ~n26267;
  assign n26269 = ~n26146 & n26267;
  assign n26270 = ~n26268 & ~n26269;
  assign n26271 = n7380 & n23394;
  assign n26272 = n7243 & n20355;
  assign n26273 = n6653 & n20358;
  assign n26274 = n6647 & n23404;
  assign n26275 = ~n26272 & ~n26273;
  assign n26276 = ~n26271 & n26275;
  assign n26277 = ~n26274 & n26276;
  assign n26278 = pi14  & n26277;
  assign n26279 = ~pi14  & ~n26277;
  assign n26280 = ~n26278 & ~n26279;
  assign n26281 = n26270 & ~n26280;
  assign n26282 = ~n26270 & n26280;
  assign n26283 = ~n26281 & ~n26282;
  assign n26284 = n26145 & ~n26283;
  assign n26285 = ~n26145 & n26283;
  assign n26286 = ~n26284 & ~n26285;
  assign n26287 = n8161 & n23765;
  assign n26288 = n7847 & n23768;
  assign n26289 = n7554 & n23771;
  assign n26290 = n7548 & n23789;
  assign n26291 = ~n26288 & ~n26289;
  assign n26292 = ~n26287 & n26291;
  assign n26293 = ~n26290 & n26292;
  assign n26294 = pi11  & n26293;
  assign n26295 = ~pi11  & ~n26293;
  assign n26296 = ~n26294 & ~n26295;
  assign n26297 = n26286 & ~n26296;
  assign n26298 = ~n26286 & n26296;
  assign n26299 = ~n26297 & ~n26298;
  assign n26300 = n26144 & ~n26299;
  assign n26301 = ~n26144 & n26299;
  assign n26302 = ~n26300 & ~n26301;
  assign n26303 = n9355 & n25022;
  assign n26304 = n8939 & n24779;
  assign n26305 = n8206 & n24529;
  assign n26306 = n8200 & n25032;
  assign n26307 = ~n26304 & ~n26305;
  assign n26308 = ~n26303 & n26307;
  assign n26309 = ~n26306 & n26308;
  assign n26310 = pi8  & n26309;
  assign n26311 = ~pi8  & ~n26309;
  assign n26312 = ~n26310 & ~n26311;
  assign n26313 = n26302 & ~n26312;
  assign n26314 = ~n26302 & n26312;
  assign n26315 = ~n26313 & ~n26314;
  assign n26316 = n26143 & ~n26315;
  assign n26317 = ~n26143 & n26315;
  assign n26318 = ~n26316 & ~n26317;
  assign n26319 = n71 & n25709;
  assign n26320 = n10329 & n25490;
  assign n26321 = n9836 & n25253;
  assign n26322 = n9830 & n25719;
  assign n26323 = ~n26320 & ~n26321;
  assign n26324 = ~n26319 & n26323;
  assign n26325 = ~n26322 & n26324;
  assign n26326 = pi5  & n26325;
  assign n26327 = ~pi5  & ~n26325;
  assign n26328 = ~n26326 & ~n26327;
  assign n26329 = n26318 & ~n26328;
  assign n26330 = ~n26318 & n26328;
  assign n26331 = ~n26329 & ~n26330;
  assign n26332 = n26142 & ~n26331;
  assign n26333 = ~n26142 & n26331;
  assign n26334 = ~n26332 & ~n26333;
  assign n26335 = ~n26133 & ~n26137;
  assign n26336 = ~n26334 & n26335;
  assign n26337 = n26334 & ~n26335;
  assign n26338 = ~n26336 & ~n26337;
  assign n26339 = n26139 & n26338;
  assign n26340 = ~n26139 & ~n26338;
  assign po8  = ~n26339 & ~n26340;
  assign n26342 = ~n26317 & ~n26329;
  assign n26343 = ~n26301 & ~n26313;
  assign n26344 = ~n13942 & n25709;
  assign n26345 = n9836 & n25490;
  assign n26346 = n9830 & ~n25925;
  assign n26347 = ~n26344 & ~n26345;
  assign n26348 = ~n26346 & n26347;
  assign n26349 = pi5  & n26348;
  assign n26350 = ~pi5  & ~n26348;
  assign n26351 = ~n26349 & ~n26350;
  assign n26352 = ~n26343 & ~n26351;
  assign n26353 = n26343 & n26351;
  assign n26354 = ~n26352 & ~n26353;
  assign n26355 = ~n26285 & ~n26297;
  assign n26356 = ~n26269 & ~n26281;
  assign n26357 = ~n26253 & ~n26265;
  assign n26358 = ~n26237 & ~n26249;
  assign n26359 = ~n26221 & ~n26233;
  assign n26360 = ~n26213 & ~n26216;
  assign n26361 = n4721 & n20386;
  assign n26362 = n4691 & n20389;
  assign n26363 = n4515 & n20392;
  assign n26364 = n4516 & n21752;
  assign n26365 = ~n26362 & ~n26363;
  assign n26366 = ~n26361 & n26365;
  assign n26367 = ~n26364 & n26366;
  assign n26368 = pi26  & n26367;
  assign n26369 = ~pi26  & ~n26367;
  assign n26370 = ~n26368 & ~n26369;
  assign n26371 = ~n26197 & ~n26201;
  assign n26372 = ~n26182 & ~n26187;
  assign n26373 = ~n92 & ~n580;
  assign n26374 = ~n676 & n26373;
  assign n26375 = n882 & n927;
  assign n26376 = n1944 & n3078;
  assign n26377 = n3351 & n5372;
  assign n26378 = n26376 & n26377;
  assign n26379 = n26374 & n26375;
  assign n26380 = n3074 & n26379;
  assign n26381 = n4086 & n26378;
  assign n26382 = n14138 & n26381;
  assign n26383 = n1519 & n26380;
  assign n26384 = n5702 & n26383;
  assign n26385 = n26382 & n26384;
  assign n26386 = n2880 & n26385;
  assign n26387 = n1707 & n26386;
  assign n26388 = ~n25973 & ~n26387;
  assign n26389 = n25973 & n26387;
  assign n26390 = ~n26388 & ~n26389;
  assign n26391 = ~n26372 & n26390;
  assign n26392 = n26372 & ~n26390;
  assign n26393 = ~n26391 & ~n26392;
  assign n26394 = n3896 & n20404;
  assign n26395 = n3683 & n20407;
  assign n26396 = n564 & n20410;
  assign n26397 = n566 & n20991;
  assign n26398 = ~n26395 & ~n26396;
  assign n26399 = ~n26394 & n26398;
  assign n26400 = ~n26397 & n26399;
  assign n26401 = n26393 & ~n26400;
  assign n26402 = ~n26393 & n26400;
  assign n26403 = ~n26401 & ~n26402;
  assign n26404 = n26371 & ~n26403;
  assign n26405 = ~n26371 & n26403;
  assign n26406 = ~n26404 & ~n26405;
  assign n26407 = n4472 & n20395;
  assign n26408 = n4070 & n20398;
  assign n26409 = n3943 & n20401;
  assign n26410 = n3944 & n21305;
  assign n26411 = ~n26408 & ~n26409;
  assign n26412 = ~n26407 & n26411;
  assign n26413 = ~n26410 & n26412;
  assign n26414 = pi29  & n26413;
  assign n26415 = ~pi29  & ~n26413;
  assign n26416 = ~n26414 & ~n26415;
  assign n26417 = n26406 & ~n26416;
  assign n26418 = ~n26406 & n26416;
  assign n26419 = ~n26417 & ~n26418;
  assign n26420 = ~n26370 & n26419;
  assign n26421 = n26370 & ~n26419;
  assign n26422 = ~n26420 & ~n26421;
  assign n26423 = n26360 & ~n26422;
  assign n26424 = ~n26360 & n26422;
  assign n26425 = ~n26423 & ~n26424;
  assign n26426 = n5267 & n20377;
  assign n26427 = n5185 & n20380;
  assign n26428 = n5121 & n20383;
  assign n26429 = n78 & n22083;
  assign n26430 = ~n26427 & ~n26428;
  assign n26431 = ~n26426 & n26430;
  assign n26432 = ~n26429 & n26431;
  assign n26433 = pi23  & n26432;
  assign n26434 = ~pi23  & ~n26432;
  assign n26435 = ~n26433 & ~n26434;
  assign n26436 = n26425 & ~n26435;
  assign n26437 = ~n26425 & n26435;
  assign n26438 = ~n26436 & ~n26437;
  assign n26439 = n26359 & ~n26438;
  assign n26440 = ~n26359 & n26438;
  assign n26441 = ~n26439 & ~n26440;
  assign n26442 = n5982 & n20368;
  assign n26443 = n5901 & n20371;
  assign n26444 = n5312 & n20374;
  assign n26445 = n5306 & n22235;
  assign n26446 = ~n26443 & ~n26444;
  assign n26447 = ~n26442 & n26446;
  assign n26448 = ~n26445 & n26447;
  assign n26449 = pi20  & n26448;
  assign n26450 = ~pi20  & ~n26448;
  assign n26451 = ~n26449 & ~n26450;
  assign n26452 = n26441 & ~n26451;
  assign n26453 = ~n26441 & n26451;
  assign n26454 = ~n26452 & ~n26453;
  assign n26455 = n26358 & ~n26454;
  assign n26456 = ~n26358 & n26454;
  assign n26457 = ~n26455 & ~n26456;
  assign n26458 = n6608 & n20358;
  assign n26459 = n6356 & n20361;
  assign n26460 = n6140 & n20365;
  assign n26461 = n6134 & n22833;
  assign n26462 = ~n26459 & ~n26460;
  assign n26463 = ~n26458 & n26462;
  assign n26464 = ~n26461 & n26463;
  assign n26465 = pi17  & n26464;
  assign n26466 = ~pi17  & ~n26464;
  assign n26467 = ~n26465 & ~n26466;
  assign n26468 = n26457 & ~n26467;
  assign n26469 = ~n26457 & n26467;
  assign n26470 = ~n26468 & ~n26469;
  assign n26471 = n26357 & ~n26470;
  assign n26472 = ~n26357 & n26470;
  assign n26473 = ~n26471 & ~n26472;
  assign n26474 = n7380 & n23771;
  assign n26475 = n7243 & n23394;
  assign n26476 = n6653 & n20355;
  assign n26477 = n6647 & n23816;
  assign n26478 = ~n26475 & ~n26476;
  assign n26479 = ~n26474 & n26478;
  assign n26480 = ~n26477 & n26479;
  assign n26481 = pi14  & n26480;
  assign n26482 = ~pi14  & ~n26480;
  assign n26483 = ~n26481 & ~n26482;
  assign n26484 = n26473 & ~n26483;
  assign n26485 = ~n26473 & n26483;
  assign n26486 = ~n26484 & ~n26485;
  assign n26487 = n26356 & ~n26486;
  assign n26488 = ~n26356 & n26486;
  assign n26489 = ~n26487 & ~n26488;
  assign n26490 = n8161 & n24529;
  assign n26491 = n7847 & n23765;
  assign n26492 = n7554 & n23768;
  assign n26493 = n7548 & n24539;
  assign n26494 = ~n26491 & ~n26492;
  assign n26495 = ~n26490 & n26494;
  assign n26496 = ~n26493 & n26495;
  assign n26497 = pi11  & n26496;
  assign n26498 = ~pi11  & ~n26496;
  assign n26499 = ~n26497 & ~n26498;
  assign n26500 = n26489 & ~n26499;
  assign n26501 = ~n26489 & n26499;
  assign n26502 = ~n26500 & ~n26501;
  assign n26503 = n26355 & ~n26502;
  assign n26504 = ~n26355 & n26502;
  assign n26505 = ~n26503 & ~n26504;
  assign n26506 = n9355 & n25253;
  assign n26507 = n8939 & n25022;
  assign n26508 = n8206 & n24779;
  assign n26509 = n8200 & n25263;
  assign n26510 = ~n26507 & ~n26508;
  assign n26511 = ~n26506 & n26510;
  assign n26512 = ~n26509 & n26511;
  assign n26513 = pi8  & n26512;
  assign n26514 = ~pi8  & ~n26512;
  assign n26515 = ~n26513 & ~n26514;
  assign n26516 = n26505 & ~n26515;
  assign n26517 = ~n26505 & n26515;
  assign n26518 = ~n26516 & ~n26517;
  assign n26519 = n26354 & n26518;
  assign n26520 = ~n26354 & ~n26518;
  assign n26521 = ~n26519 & ~n26520;
  assign n26522 = n26342 & ~n26521;
  assign n26523 = ~n26342 & n26521;
  assign n26524 = ~n26522 & ~n26523;
  assign n26525 = ~n26333 & ~n26337;
  assign n26526 = ~n26524 & n26525;
  assign n26527 = n26524 & ~n26525;
  assign n26528 = ~n26526 & ~n26527;
  assign n26529 = n26339 & n26528;
  assign n26530 = ~n26339 & ~n26528;
  assign po9  = ~n26529 & ~n26530;
  assign n26532 = ~n26523 & ~n26527;
  assign n26533 = ~n26352 & ~n26519;
  assign n26534 = ~n26488 & ~n26500;
  assign n26535 = ~n26456 & ~n26468;
  assign n26536 = ~n26440 & ~n26452;
  assign n26537 = ~n26424 & ~n26436;
  assign n26538 = ~n26417 & ~n26420;
  assign n26539 = n4721 & n20383;
  assign n26540 = n4691 & n20386;
  assign n26541 = n4515 & n20389;
  assign n26542 = n4516 & n21737;
  assign n26543 = ~n26540 & ~n26541;
  assign n26544 = ~n26539 & n26543;
  assign n26545 = ~n26542 & n26544;
  assign n26546 = pi26  & n26545;
  assign n26547 = ~pi26  & ~n26545;
  assign n26548 = ~n26546 & ~n26547;
  assign n26549 = ~n26401 & ~n26405;
  assign n26550 = ~n26388 & ~n26391;
  assign n26551 = ~n13943 & n25709;
  assign n26552 = ~pi5  & n26551;
  assign n26553 = pi5  & ~n26551;
  assign n26554 = ~n26552 & ~n26553;
  assign n26555 = ~n466 & ~n483;
  assign n26556 = ~n662 & ~n683;
  assign n26557 = n26555 & n26556;
  assign n26558 = n146 & n497;
  assign n26559 = n1862 & n1911;
  assign n26560 = n3154 & n4932;
  assign n26561 = n26559 & n26560;
  assign n26562 = n26557 & n26558;
  assign n26563 = n5551 & n26562;
  assign n26564 = n12771 & n26561;
  assign n26565 = n26563 & n26564;
  assign n26566 = n21634 & n26565;
  assign n26567 = n4285 & n26566;
  assign n26568 = n2596 & n26567;
  assign n26569 = n25973 & ~n26568;
  assign n26570 = ~n25973 & n26568;
  assign n26571 = ~n26569 & ~n26570;
  assign n26572 = n26554 & n26571;
  assign n26573 = ~n26554 & ~n26571;
  assign n26574 = ~n26572 & ~n26573;
  assign n26575 = ~n26550 & n26574;
  assign n26576 = n26550 & ~n26574;
  assign n26577 = ~n26575 & ~n26576;
  assign n26578 = n3896 & n20401;
  assign n26579 = n3683 & n20404;
  assign n26580 = n564 & n20407;
  assign n26581 = n566 & n21286;
  assign n26582 = ~n26579 & ~n26580;
  assign n26583 = ~n26578 & n26582;
  assign n26584 = ~n26581 & n26583;
  assign n26585 = n26577 & ~n26584;
  assign n26586 = ~n26577 & n26584;
  assign n26587 = ~n26585 & ~n26586;
  assign n26588 = n26549 & ~n26587;
  assign n26589 = ~n26549 & n26587;
  assign n26590 = ~n26588 & ~n26589;
  assign n26591 = n4472 & n20392;
  assign n26592 = n4070 & n20395;
  assign n26593 = n3943 & n20398;
  assign n26594 = n3944 & n20586;
  assign n26595 = ~n26592 & ~n26593;
  assign n26596 = ~n26591 & n26595;
  assign n26597 = ~n26594 & n26596;
  assign n26598 = pi29  & n26597;
  assign n26599 = ~pi29  & ~n26597;
  assign n26600 = ~n26598 & ~n26599;
  assign n26601 = n26590 & ~n26600;
  assign n26602 = ~n26590 & n26600;
  assign n26603 = ~n26601 & ~n26602;
  assign n26604 = ~n26548 & n26603;
  assign n26605 = n26548 & ~n26603;
  assign n26606 = ~n26604 & ~n26605;
  assign n26607 = n26538 & ~n26606;
  assign n26608 = ~n26538 & n26606;
  assign n26609 = ~n26607 & ~n26608;
  assign n26610 = n5267 & n20374;
  assign n26611 = n5185 & n20377;
  assign n26612 = n5121 & n20380;
  assign n26613 = n78 & n22263;
  assign n26614 = ~n26611 & ~n26612;
  assign n26615 = ~n26610 & n26614;
  assign n26616 = ~n26613 & n26615;
  assign n26617 = pi23  & n26616;
  assign n26618 = ~pi23  & ~n26616;
  assign n26619 = ~n26617 & ~n26618;
  assign n26620 = n26609 & ~n26619;
  assign n26621 = ~n26609 & n26619;
  assign n26622 = ~n26620 & ~n26621;
  assign n26623 = n26537 & ~n26622;
  assign n26624 = ~n26537 & n26622;
  assign n26625 = ~n26623 & ~n26624;
  assign n26626 = n5982 & n20365;
  assign n26627 = n5901 & n20368;
  assign n26628 = n5312 & n20371;
  assign n26629 = n5306 & n22814;
  assign n26630 = ~n26627 & ~n26628;
  assign n26631 = ~n26626 & n26630;
  assign n26632 = ~n26629 & n26631;
  assign n26633 = pi20  & n26632;
  assign n26634 = ~pi20  & ~n26632;
  assign n26635 = ~n26633 & ~n26634;
  assign n26636 = n26625 & ~n26635;
  assign n26637 = ~n26625 & n26635;
  assign n26638 = ~n26636 & ~n26637;
  assign n26639 = n26536 & ~n26638;
  assign n26640 = ~n26536 & n26638;
  assign n26641 = ~n26639 & ~n26640;
  assign n26642 = n6608 & n20355;
  assign n26643 = n6356 & n20358;
  assign n26644 = n6140 & n20361;
  assign n26645 = n6134 & n20562;
  assign n26646 = ~n26643 & ~n26644;
  assign n26647 = ~n26642 & n26646;
  assign n26648 = ~n26645 & n26647;
  assign n26649 = pi17  & n26648;
  assign n26650 = ~pi17  & ~n26648;
  assign n26651 = ~n26649 & ~n26650;
  assign n26652 = n26641 & ~n26651;
  assign n26653 = ~n26641 & n26651;
  assign n26654 = ~n26652 & ~n26653;
  assign n26655 = n26535 & ~n26654;
  assign n26656 = ~n26535 & n26654;
  assign n26657 = ~n26655 & ~n26656;
  assign n26658 = ~n26472 & ~n26484;
  assign n26659 = n7380 & n23768;
  assign n26660 = n7243 & n23771;
  assign n26661 = n6653 & n23394;
  assign n26662 = n6647 & n23804;
  assign n26663 = ~n26660 & ~n26661;
  assign n26664 = ~n26659 & n26663;
  assign n26665 = ~n26662 & n26664;
  assign n26666 = pi14  & n26665;
  assign n26667 = ~pi14  & ~n26665;
  assign n26668 = ~n26666 & ~n26667;
  assign n26669 = ~n26658 & ~n26668;
  assign n26670 = n26658 & n26668;
  assign n26671 = ~n26669 & ~n26670;
  assign n26672 = ~n26657 & ~n26671;
  assign n26673 = n26657 & n26671;
  assign n26674 = ~n26672 & ~n26673;
  assign n26675 = n8161 & n24779;
  assign n26676 = n7847 & n24529;
  assign n26677 = n7554 & n23765;
  assign n26678 = n7548 & n24789;
  assign n26679 = ~n26676 & ~n26677;
  assign n26680 = ~n26675 & n26679;
  assign n26681 = ~n26678 & n26680;
  assign n26682 = pi11  & n26681;
  assign n26683 = ~pi11  & ~n26681;
  assign n26684 = ~n26682 & ~n26683;
  assign n26685 = n26674 & ~n26684;
  assign n26686 = ~n26674 & n26684;
  assign n26687 = ~n26685 & ~n26686;
  assign n26688 = n26534 & ~n26687;
  assign n26689 = ~n26534 & n26687;
  assign n26690 = ~n26688 & ~n26689;
  assign n26691 = ~n26504 & ~n26516;
  assign n26692 = n9355 & n25490;
  assign n26693 = n8939 & n25253;
  assign n26694 = n8206 & n25022;
  assign n26695 = n8200 & n25500;
  assign n26696 = ~n26693 & ~n26694;
  assign n26697 = ~n26692 & n26696;
  assign n26698 = ~n26695 & n26697;
  assign n26699 = pi8  & n26698;
  assign n26700 = ~pi8  & ~n26698;
  assign n26701 = ~n26699 & ~n26700;
  assign n26702 = ~n26691 & ~n26701;
  assign n26703 = n26691 & n26701;
  assign n26704 = ~n26702 & ~n26703;
  assign n26705 = ~n26690 & ~n26704;
  assign n26706 = n26690 & n26704;
  assign n26707 = ~n26705 & ~n26706;
  assign n26708 = ~n26533 & n26707;
  assign n26709 = n26533 & ~n26707;
  assign n26710 = ~n26708 & ~n26709;
  assign n26711 = ~n26532 & n26710;
  assign n26712 = n26532 & ~n26710;
  assign n26713 = ~n26711 & ~n26712;
  assign n26714 = ~n26529 & ~n26713;
  assign n26715 = n26529 & n26713;
  assign po10  = ~n26714 & ~n26715;
  assign n26717 = ~n26708 & ~n26711;
  assign n26718 = ~n26702 & ~n26706;
  assign n26719 = ~n26685 & ~n26689;
  assign n26720 = ~n26669 & ~n26673;
  assign n26721 = ~n26652 & ~n26656;
  assign n26722 = ~n26636 & ~n26640;
  assign n26723 = ~n26620 & ~n26624;
  assign n26724 = ~n26604 & ~n26608;
  assign n26725 = ~n26589 & ~n26601;
  assign n26726 = ~n26575 & ~n26585;
  assign n26727 = ~n26569 & ~n26572;
  assign n26728 = n840 & n926;
  assign n26729 = n1347 & n1754;
  assign n26730 = n2049 & n2086;
  assign n26731 = n13406 & n26730;
  assign n26732 = n26728 & n26729;
  assign n26733 = n2000 & n26732;
  assign n26734 = n6439 & n26731;
  assign n26735 = n7059 & n26734;
  assign n26736 = n1131 & n26733;
  assign n26737 = n26735 & n26736;
  assign n26738 = ~n92 & ~n216;
  assign n26739 = ~n235 & ~n406;
  assign n26740 = ~n421 & n26739;
  assign n26741 = n1232 & n26738;
  assign n26742 = n1237 & n1242;
  assign n26743 = n2271 & n2455;
  assign n26744 = n4267 & n4384;
  assign n26745 = n26743 & n26744;
  assign n26746 = n26741 & n26742;
  assign n26747 = n3345 & n26740;
  assign n26748 = n26746 & n26747;
  assign n26749 = n1592 & n26745;
  assign n26750 = n7021 & n26749;
  assign n26751 = n2177 & n26748;
  assign n26752 = n26750 & n26751;
  assign n26753 = n26737 & n26752;
  assign n26754 = n1500 & n26753;
  assign n26755 = ~n26727 & n26754;
  assign n26756 = n26727 & ~n26754;
  assign n26757 = ~n26755 & ~n26756;
  assign n26758 = n3896 & n20398;
  assign n26759 = n3683 & n20401;
  assign n26760 = n564 & n20404;
  assign n26761 = n566 & n21322;
  assign n26762 = ~n26759 & ~n26760;
  assign n26763 = ~n26758 & n26762;
  assign n26764 = ~n26761 & n26763;
  assign n26765 = n26757 & ~n26764;
  assign n26766 = ~n26757 & n26764;
  assign n26767 = ~n26765 & ~n26766;
  assign n26768 = n26726 & ~n26767;
  assign n26769 = ~n26726 & n26767;
  assign n26770 = ~n26768 & ~n26769;
  assign n26771 = n4472 & n20389;
  assign n26772 = n4070 & n20392;
  assign n26773 = n3943 & n20395;
  assign n26774 = n3944 & n21716;
  assign n26775 = ~n26772 & ~n26773;
  assign n26776 = ~n26771 & n26775;
  assign n26777 = ~n26774 & n26776;
  assign n26778 = pi29  & n26777;
  assign n26779 = ~pi29  & ~n26777;
  assign n26780 = ~n26778 & ~n26779;
  assign n26781 = n26770 & ~n26780;
  assign n26782 = ~n26770 & n26780;
  assign n26783 = ~n26781 & ~n26782;
  assign n26784 = ~n26725 & n26783;
  assign n26785 = n26725 & ~n26783;
  assign n26786 = ~n26784 & ~n26785;
  assign n26787 = n4721 & n20380;
  assign n26788 = n4691 & n20383;
  assign n26789 = n4515 & n20386;
  assign n26790 = n4516 & n20574;
  assign n26791 = ~n26788 & ~n26789;
  assign n26792 = ~n26787 & n26791;
  assign n26793 = ~n26790 & n26792;
  assign n26794 = pi26  & n26793;
  assign n26795 = ~pi26  & ~n26793;
  assign n26796 = ~n26794 & ~n26795;
  assign n26797 = n26786 & ~n26796;
  assign n26798 = ~n26786 & n26796;
  assign n26799 = ~n26797 & ~n26798;
  assign n26800 = n26724 & ~n26799;
  assign n26801 = ~n26724 & n26799;
  assign n26802 = ~n26800 & ~n26801;
  assign n26803 = n5267 & n20371;
  assign n26804 = n5185 & n20374;
  assign n26805 = n5121 & n20377;
  assign n26806 = n78 & n22250;
  assign n26807 = ~n26804 & ~n26805;
  assign n26808 = ~n26803 & n26807;
  assign n26809 = ~n26806 & n26808;
  assign n26810 = pi23  & n26809;
  assign n26811 = ~pi23  & ~n26809;
  assign n26812 = ~n26810 & ~n26811;
  assign n26813 = n26802 & ~n26812;
  assign n26814 = ~n26802 & n26812;
  assign n26815 = ~n26813 & ~n26814;
  assign n26816 = n26723 & ~n26815;
  assign n26817 = ~n26723 & n26815;
  assign n26818 = ~n26816 & ~n26817;
  assign n26819 = n5982 & n20361;
  assign n26820 = n5901 & n20365;
  assign n26821 = n5312 & n20368;
  assign n26822 = n5306 & n22848;
  assign n26823 = ~n26820 & ~n26821;
  assign n26824 = ~n26819 & n26823;
  assign n26825 = ~n26822 & n26824;
  assign n26826 = pi20  & n26825;
  assign n26827 = ~pi20  & ~n26825;
  assign n26828 = ~n26826 & ~n26827;
  assign n26829 = n26818 & ~n26828;
  assign n26830 = ~n26818 & n26828;
  assign n26831 = ~n26829 & ~n26830;
  assign n26832 = n26722 & ~n26831;
  assign n26833 = ~n26722 & n26831;
  assign n26834 = ~n26832 & ~n26833;
  assign n26835 = n6608 & n23394;
  assign n26836 = n6356 & n20355;
  assign n26837 = n6140 & n20358;
  assign n26838 = n6134 & n23404;
  assign n26839 = ~n26836 & ~n26837;
  assign n26840 = ~n26835 & n26839;
  assign n26841 = ~n26838 & n26840;
  assign n26842 = pi17  & n26841;
  assign n26843 = ~pi17  & ~n26841;
  assign n26844 = ~n26842 & ~n26843;
  assign n26845 = n26834 & ~n26844;
  assign n26846 = ~n26834 & n26844;
  assign n26847 = ~n26845 & ~n26846;
  assign n26848 = n26721 & ~n26847;
  assign n26849 = ~n26721 & n26847;
  assign n26850 = ~n26848 & ~n26849;
  assign n26851 = n7380 & n23765;
  assign n26852 = n7243 & n23768;
  assign n26853 = n6653 & n23771;
  assign n26854 = n6647 & n23789;
  assign n26855 = ~n26852 & ~n26853;
  assign n26856 = ~n26851 & n26855;
  assign n26857 = ~n26854 & n26856;
  assign n26858 = pi14  & n26857;
  assign n26859 = ~pi14  & ~n26857;
  assign n26860 = ~n26858 & ~n26859;
  assign n26861 = n26850 & ~n26860;
  assign n26862 = ~n26850 & n26860;
  assign n26863 = ~n26861 & ~n26862;
  assign n26864 = ~n26720 & n26863;
  assign n26865 = n26720 & ~n26863;
  assign n26866 = ~n26864 & ~n26865;
  assign n26867 = n8161 & n25022;
  assign n26868 = n7847 & n24779;
  assign n26869 = n7554 & n24529;
  assign n26870 = n7548 & n25032;
  assign n26871 = ~n26868 & ~n26869;
  assign n26872 = ~n26867 & n26871;
  assign n26873 = ~n26870 & n26872;
  assign n26874 = pi11  & n26873;
  assign n26875 = ~pi11  & ~n26873;
  assign n26876 = ~n26874 & ~n26875;
  assign n26877 = n26866 & ~n26876;
  assign n26878 = ~n26866 & n26876;
  assign n26879 = ~n26877 & ~n26878;
  assign n26880 = n26719 & ~n26879;
  assign n26881 = ~n26719 & n26879;
  assign n26882 = ~n26880 & ~n26881;
  assign n26883 = n9355 & n25709;
  assign n26884 = n8939 & n25490;
  assign n26885 = n8206 & n25253;
  assign n26886 = n8200 & n25719;
  assign n26887 = ~n26884 & ~n26885;
  assign n26888 = ~n26883 & n26887;
  assign n26889 = ~n26886 & n26888;
  assign n26890 = pi8  & n26889;
  assign n26891 = ~pi8  & ~n26889;
  assign n26892 = ~n26890 & ~n26891;
  assign n26893 = n26882 & ~n26892;
  assign n26894 = ~n26882 & n26892;
  assign n26895 = ~n26893 & ~n26894;
  assign n26896 = ~n26718 & n26895;
  assign n26897 = n26718 & ~n26895;
  assign n26898 = ~n26896 & ~n26897;
  assign n26899 = n26717 & ~n26898;
  assign n26900 = ~n26717 & n26898;
  assign n26901 = ~n26899 & ~n26900;
  assign n26902 = n26715 & n26901;
  assign n26903 = ~n26715 & ~n26901;
  assign po11  = ~n26902 & ~n26903;
  assign n26905 = ~n26881 & ~n26893;
  assign n26906 = ~n26864 & ~n26877;
  assign n26907 = ~n13513 & n25709;
  assign n26908 = n8206 & n25490;
  assign n26909 = n8200 & ~n25925;
  assign n26910 = ~n26907 & ~n26908;
  assign n26911 = ~n26909 & n26910;
  assign n26912 = pi8  & n26911;
  assign n26913 = ~pi8  & ~n26911;
  assign n26914 = ~n26912 & ~n26913;
  assign n26915 = ~n26906 & ~n26914;
  assign n26916 = n26906 & n26914;
  assign n26917 = ~n26915 & ~n26916;
  assign n26918 = ~n26849 & ~n26861;
  assign n26919 = ~n26833 & ~n26845;
  assign n26920 = ~n26817 & ~n26829;
  assign n26921 = ~n26801 & ~n26813;
  assign n26922 = ~n26784 & ~n26797;
  assign n26923 = n4721 & n20377;
  assign n26924 = n4691 & n20380;
  assign n26925 = n4515 & n20383;
  assign n26926 = n4516 & n22083;
  assign n26927 = ~n26924 & ~n26925;
  assign n26928 = ~n26923 & n26927;
  assign n26929 = ~n26926 & n26928;
  assign n26930 = pi26  & n26929;
  assign n26931 = ~pi26  & ~n26929;
  assign n26932 = ~n26930 & ~n26931;
  assign n26933 = ~n26769 & ~n26781;
  assign n26934 = ~n26755 & ~n26765;
  assign n26935 = ~n334 & ~n469;
  assign n26936 = ~n553 & n26935;
  assign n26937 = n523 & n1760;
  assign n26938 = n2473 & n3071;
  assign n26939 = n3073 & n26938;
  assign n26940 = n26936 & n26937;
  assign n26941 = n3808 & n4934;
  assign n26942 = n26940 & n26941;
  assign n26943 = n1782 & n26939;
  assign n26944 = n26942 & n26943;
  assign n26945 = n3091 & n26944;
  assign n26946 = ~n163 & ~n251;
  assign n26947 = ~n316 & ~n421;
  assign n26948 = ~n577 & n26947;
  assign n26949 = n744 & n26946;
  assign n26950 = n5682 & n26949;
  assign n26951 = n26948 & n26950;
  assign n26952 = ~n162 & ~n307;
  assign n26953 = ~n459 & ~n671;
  assign n26954 = n26952 & n26953;
  assign n26955 = n428 & n2870;
  assign n26956 = n26954 & n26955;
  assign n26957 = n6882 & n12457;
  assign n26958 = n26956 & n26957;
  assign n26959 = n4263 & n26958;
  assign n26960 = n26951 & n26959;
  assign n26961 = n4155 & n26960;
  assign n26962 = n26945 & n26961;
  assign n26963 = n12751 & n26962;
  assign n26964 = ~n26754 & n26963;
  assign n26965 = n26754 & ~n26963;
  assign n26966 = ~n26964 & ~n26965;
  assign n26967 = ~n26934 & n26966;
  assign n26968 = n26934 & ~n26966;
  assign n26969 = ~n26967 & ~n26968;
  assign n26970 = n3896 & n20395;
  assign n26971 = n3683 & n20398;
  assign n26972 = n564 & n20401;
  assign n26973 = n566 & n21305;
  assign n26974 = ~n26971 & ~n26972;
  assign n26975 = ~n26970 & n26974;
  assign n26976 = ~n26973 & n26975;
  assign n26977 = n26969 & ~n26976;
  assign n26978 = ~n26969 & n26976;
  assign n26979 = ~n26977 & ~n26978;
  assign n26980 = n26933 & ~n26979;
  assign n26981 = ~n26933 & n26979;
  assign n26982 = ~n26980 & ~n26981;
  assign n26983 = n4472 & n20386;
  assign n26984 = n4070 & n20389;
  assign n26985 = n3943 & n20392;
  assign n26986 = n3944 & n21752;
  assign n26987 = ~n26984 & ~n26985;
  assign n26988 = ~n26983 & n26987;
  assign n26989 = ~n26986 & n26988;
  assign n26990 = pi29  & n26989;
  assign n26991 = ~pi29  & ~n26989;
  assign n26992 = ~n26990 & ~n26991;
  assign n26993 = n26982 & ~n26992;
  assign n26994 = ~n26982 & n26992;
  assign n26995 = ~n26993 & ~n26994;
  assign n26996 = ~n26932 & n26995;
  assign n26997 = n26932 & ~n26995;
  assign n26998 = ~n26996 & ~n26997;
  assign n26999 = n26922 & ~n26998;
  assign n27000 = ~n26922 & n26998;
  assign n27001 = ~n26999 & ~n27000;
  assign n27002 = n5267 & n20368;
  assign n27003 = n5185 & n20371;
  assign n27004 = n5121 & n20374;
  assign n27005 = n78 & n22235;
  assign n27006 = ~n27003 & ~n27004;
  assign n27007 = ~n27002 & n27006;
  assign n27008 = ~n27005 & n27007;
  assign n27009 = pi23  & n27008;
  assign n27010 = ~pi23  & ~n27008;
  assign n27011 = ~n27009 & ~n27010;
  assign n27012 = n27001 & ~n27011;
  assign n27013 = ~n27001 & n27011;
  assign n27014 = ~n27012 & ~n27013;
  assign n27015 = n26921 & ~n27014;
  assign n27016 = ~n26921 & n27014;
  assign n27017 = ~n27015 & ~n27016;
  assign n27018 = n5982 & n20358;
  assign n27019 = n5901 & n20361;
  assign n27020 = n5312 & n20365;
  assign n27021 = n5306 & n22833;
  assign n27022 = ~n27019 & ~n27020;
  assign n27023 = ~n27018 & n27022;
  assign n27024 = ~n27021 & n27023;
  assign n27025 = pi20  & n27024;
  assign n27026 = ~pi20  & ~n27024;
  assign n27027 = ~n27025 & ~n27026;
  assign n27028 = n27017 & ~n27027;
  assign n27029 = ~n27017 & n27027;
  assign n27030 = ~n27028 & ~n27029;
  assign n27031 = n26920 & ~n27030;
  assign n27032 = ~n26920 & n27030;
  assign n27033 = ~n27031 & ~n27032;
  assign n27034 = n6608 & n23771;
  assign n27035 = n6356 & n23394;
  assign n27036 = n6140 & n20355;
  assign n27037 = n6134 & n23816;
  assign n27038 = ~n27035 & ~n27036;
  assign n27039 = ~n27034 & n27038;
  assign n27040 = ~n27037 & n27039;
  assign n27041 = pi17  & n27040;
  assign n27042 = ~pi17  & ~n27040;
  assign n27043 = ~n27041 & ~n27042;
  assign n27044 = n27033 & ~n27043;
  assign n27045 = ~n27033 & n27043;
  assign n27046 = ~n27044 & ~n27045;
  assign n27047 = n26919 & ~n27046;
  assign n27048 = ~n26919 & n27046;
  assign n27049 = ~n27047 & ~n27048;
  assign n27050 = n7380 & n24529;
  assign n27051 = n7243 & n23765;
  assign n27052 = n6653 & n23768;
  assign n27053 = n6647 & n24539;
  assign n27054 = ~n27051 & ~n27052;
  assign n27055 = ~n27050 & n27054;
  assign n27056 = ~n27053 & n27055;
  assign n27057 = pi14  & n27056;
  assign n27058 = ~pi14  & ~n27056;
  assign n27059 = ~n27057 & ~n27058;
  assign n27060 = n27049 & ~n27059;
  assign n27061 = ~n27049 & n27059;
  assign n27062 = ~n27060 & ~n27061;
  assign n27063 = n26918 & ~n27062;
  assign n27064 = ~n26918 & n27062;
  assign n27065 = ~n27063 & ~n27064;
  assign n27066 = n8161 & n25253;
  assign n27067 = n7847 & n25022;
  assign n27068 = n7554 & n24779;
  assign n27069 = n7548 & n25263;
  assign n27070 = ~n27067 & ~n27068;
  assign n27071 = ~n27066 & n27070;
  assign n27072 = ~n27069 & n27071;
  assign n27073 = pi11  & n27072;
  assign n27074 = ~pi11  & ~n27072;
  assign n27075 = ~n27073 & ~n27074;
  assign n27076 = n27065 & ~n27075;
  assign n27077 = ~n27065 & n27075;
  assign n27078 = ~n27076 & ~n27077;
  assign n27079 = n26917 & n27078;
  assign n27080 = ~n26917 & ~n27078;
  assign n27081 = ~n27079 & ~n27080;
  assign n27082 = n26905 & ~n27081;
  assign n27083 = ~n26905 & n27081;
  assign n27084 = ~n27082 & ~n27083;
  assign n27085 = ~n26896 & ~n26900;
  assign n27086 = ~n27084 & n27085;
  assign n27087 = n27084 & ~n27085;
  assign n27088 = ~n27086 & ~n27087;
  assign n27089 = n26902 & n27088;
  assign n27090 = ~n26902 & ~n27088;
  assign po12  = ~n27089 & ~n27090;
  assign n27092 = ~n27083 & ~n27087;
  assign n27093 = ~n26915 & ~n27079;
  assign n27094 = ~n27048 & ~n27060;
  assign n27095 = ~n27016 & ~n27028;
  assign n27096 = ~n27000 & ~n27012;
  assign n27097 = ~n26993 & ~n26996;
  assign n27098 = ~n26977 & ~n26981;
  assign n27099 = n4472 & n20383;
  assign n27100 = n4070 & n20386;
  assign n27101 = n3943 & n20389;
  assign n27102 = n3944 & n21737;
  assign n27103 = ~n27100 & ~n27101;
  assign n27104 = ~n27099 & n27103;
  assign n27105 = ~n27102 & n27104;
  assign n27106 = pi29  & n27105;
  assign n27107 = ~pi29  & ~n27105;
  assign n27108 = ~n27106 & ~n27107;
  assign n27109 = ~n26965 & ~n26967;
  assign n27110 = ~n13514 & n25709;
  assign n27111 = pi8  & ~n27110;
  assign n27112 = ~pi8  & n27110;
  assign n27113 = ~n27111 & ~n27112;
  assign n27114 = ~n308 & ~n591;
  assign n27115 = n211 & n27114;
  assign n27116 = n930 & n1041;
  assign n27117 = n1862 & n27116;
  assign n27118 = n1123 & n27115;
  assign n27119 = n1396 & n2225;
  assign n27120 = n12734 & n27119;
  assign n27121 = n27117 & n27118;
  assign n27122 = n12720 & n27121;
  assign n27123 = n27120 & n27122;
  assign n27124 = n2765 & n27123;
  assign n27125 = n1299 & n3340;
  assign n27126 = n27124 & n27125;
  assign n27127 = n26754 & n27126;
  assign n27128 = ~n26754 & ~n27126;
  assign n27129 = ~n27127 & ~n27128;
  assign n27130 = n27113 & n27129;
  assign n27131 = ~n27113 & ~n27129;
  assign n27132 = ~n27130 & ~n27131;
  assign n27133 = ~n27109 & n27132;
  assign n27134 = n27109 & ~n27132;
  assign n27135 = ~n27133 & ~n27134;
  assign n27136 = n3896 & n20392;
  assign n27137 = n3683 & n20395;
  assign n27138 = n564 & n20398;
  assign n27139 = n566 & n20586;
  assign n27140 = ~n27137 & ~n27138;
  assign n27141 = ~n27136 & n27140;
  assign n27142 = ~n27139 & n27141;
  assign n27143 = n27135 & ~n27142;
  assign n27144 = ~n27135 & n27142;
  assign n27145 = ~n27143 & ~n27144;
  assign n27146 = ~n27108 & n27145;
  assign n27147 = n27108 & ~n27145;
  assign n27148 = ~n27146 & ~n27147;
  assign n27149 = n27098 & ~n27148;
  assign n27150 = ~n27098 & n27148;
  assign n27151 = ~n27149 & ~n27150;
  assign n27152 = n4721 & n20374;
  assign n27153 = n4691 & n20377;
  assign n27154 = n4515 & n20380;
  assign n27155 = n4516 & n22263;
  assign n27156 = ~n27153 & ~n27154;
  assign n27157 = ~n27152 & n27156;
  assign n27158 = ~n27155 & n27157;
  assign n27159 = pi26  & n27158;
  assign n27160 = ~pi26  & ~n27158;
  assign n27161 = ~n27159 & ~n27160;
  assign n27162 = n27151 & ~n27161;
  assign n27163 = ~n27151 & n27161;
  assign n27164 = ~n27162 & ~n27163;
  assign n27165 = n27097 & ~n27164;
  assign n27166 = ~n27097 & n27164;
  assign n27167 = ~n27165 & ~n27166;
  assign n27168 = n5267 & n20365;
  assign n27169 = n5185 & n20368;
  assign n27170 = n5121 & n20371;
  assign n27171 = n78 & n22814;
  assign n27172 = ~n27169 & ~n27170;
  assign n27173 = ~n27168 & n27172;
  assign n27174 = ~n27171 & n27173;
  assign n27175 = pi23  & n27174;
  assign n27176 = ~pi23  & ~n27174;
  assign n27177 = ~n27175 & ~n27176;
  assign n27178 = n27167 & ~n27177;
  assign n27179 = ~n27167 & n27177;
  assign n27180 = ~n27178 & ~n27179;
  assign n27181 = n27096 & ~n27180;
  assign n27182 = ~n27096 & n27180;
  assign n27183 = ~n27181 & ~n27182;
  assign n27184 = n5982 & n20355;
  assign n27185 = n5901 & n20358;
  assign n27186 = n5312 & n20361;
  assign n27187 = n5306 & n20562;
  assign n27188 = ~n27185 & ~n27186;
  assign n27189 = ~n27184 & n27188;
  assign n27190 = ~n27187 & n27189;
  assign n27191 = pi20  & n27190;
  assign n27192 = ~pi20  & ~n27190;
  assign n27193 = ~n27191 & ~n27192;
  assign n27194 = n27183 & ~n27193;
  assign n27195 = ~n27183 & n27193;
  assign n27196 = ~n27194 & ~n27195;
  assign n27197 = n27095 & ~n27196;
  assign n27198 = ~n27095 & n27196;
  assign n27199 = ~n27197 & ~n27198;
  assign n27200 = ~n27032 & ~n27044;
  assign n27201 = n6608 & n23768;
  assign n27202 = n6356 & n23771;
  assign n27203 = n6140 & n23394;
  assign n27204 = n6134 & n23804;
  assign n27205 = ~n27202 & ~n27203;
  assign n27206 = ~n27201 & n27205;
  assign n27207 = ~n27204 & n27206;
  assign n27208 = pi17  & n27207;
  assign n27209 = ~pi17  & ~n27207;
  assign n27210 = ~n27208 & ~n27209;
  assign n27211 = ~n27200 & ~n27210;
  assign n27212 = n27200 & n27210;
  assign n27213 = ~n27211 & ~n27212;
  assign n27214 = ~n27199 & ~n27213;
  assign n27215 = n27199 & n27213;
  assign n27216 = ~n27214 & ~n27215;
  assign n27217 = n7380 & n24779;
  assign n27218 = n7243 & n24529;
  assign n27219 = n6653 & n23765;
  assign n27220 = n6647 & n24789;
  assign n27221 = ~n27218 & ~n27219;
  assign n27222 = ~n27217 & n27221;
  assign n27223 = ~n27220 & n27222;
  assign n27224 = pi14  & n27223;
  assign n27225 = ~pi14  & ~n27223;
  assign n27226 = ~n27224 & ~n27225;
  assign n27227 = n27216 & ~n27226;
  assign n27228 = ~n27216 & n27226;
  assign n27229 = ~n27227 & ~n27228;
  assign n27230 = n27094 & ~n27229;
  assign n27231 = ~n27094 & n27229;
  assign n27232 = ~n27230 & ~n27231;
  assign n27233 = ~n27064 & ~n27076;
  assign n27234 = n8161 & n25490;
  assign n27235 = n7847 & n25253;
  assign n27236 = n7554 & n25022;
  assign n27237 = n7548 & n25500;
  assign n27238 = ~n27235 & ~n27236;
  assign n27239 = ~n27234 & n27238;
  assign n27240 = ~n27237 & n27239;
  assign n27241 = pi11  & n27240;
  assign n27242 = ~pi11  & ~n27240;
  assign n27243 = ~n27241 & ~n27242;
  assign n27244 = ~n27233 & ~n27243;
  assign n27245 = n27233 & n27243;
  assign n27246 = ~n27244 & ~n27245;
  assign n27247 = ~n27232 & ~n27246;
  assign n27248 = n27232 & n27246;
  assign n27249 = ~n27247 & ~n27248;
  assign n27250 = ~n27093 & n27249;
  assign n27251 = n27093 & ~n27249;
  assign n27252 = ~n27250 & ~n27251;
  assign n27253 = ~n27092 & n27252;
  assign n27254 = n27092 & ~n27252;
  assign n27255 = ~n27253 & ~n27254;
  assign n27256 = ~n27089 & ~n27255;
  assign n27257 = n27089 & n27255;
  assign po13  = ~n27256 & ~n27257;
  assign n27259 = ~n27250 & ~n27253;
  assign n27260 = ~n27244 & ~n27248;
  assign n27261 = ~n27227 & ~n27231;
  assign n27262 = n7380 & n25022;
  assign n27263 = n7243 & n24779;
  assign n27264 = n6653 & n24529;
  assign n27265 = n6647 & n25032;
  assign n27266 = ~n27263 & ~n27264;
  assign n27267 = ~n27262 & n27266;
  assign n27268 = ~n27265 & n27267;
  assign n27269 = pi14  & n27268;
  assign n27270 = ~pi14  & ~n27268;
  assign n27271 = ~n27269 & ~n27270;
  assign n27272 = ~n27211 & ~n27215;
  assign n27273 = ~n27194 & ~n27198;
  assign n27274 = ~n27178 & ~n27182;
  assign n27275 = ~n27162 & ~n27166;
  assign n27276 = ~n27146 & ~n27150;
  assign n27277 = ~n27128 & ~n27130;
  assign n27278 = ~n210 & ~n391;
  assign n27279 = ~n577 & n27278;
  assign n27280 = n931 & n3248;
  assign n27281 = n3763 & n14185;
  assign n27282 = n27280 & n27281;
  assign n27283 = n2307 & n27279;
  assign n27284 = n3230 & n14646;
  assign n27285 = n27283 & n27284;
  assign n27286 = n5337 & n27282;
  assign n27287 = n27285 & n27286;
  assign n27288 = n13341 & n27287;
  assign n27289 = n1036 & n27288;
  assign n27290 = n2515 & n27289;
  assign n27291 = ~n27277 & n27290;
  assign n27292 = n27277 & ~n27290;
  assign n27293 = ~n27291 & ~n27292;
  assign n27294 = n3896 & n20389;
  assign n27295 = n3683 & n20392;
  assign n27296 = n564 & n20395;
  assign n27297 = n566 & n21716;
  assign n27298 = ~n27295 & ~n27296;
  assign n27299 = ~n27294 & n27298;
  assign n27300 = ~n27297 & n27299;
  assign n27301 = ~n27293 & ~n27300;
  assign n27302 = n27293 & n27300;
  assign n27303 = ~n27301 & ~n27302;
  assign n27304 = ~n27133 & ~n27143;
  assign n27305 = n27303 & n27304;
  assign n27306 = ~n27303 & ~n27304;
  assign n27307 = ~n27305 & ~n27306;
  assign n27308 = n4472 & n20380;
  assign n27309 = n4070 & n20383;
  assign n27310 = n3943 & n20386;
  assign n27311 = n3944 & n20574;
  assign n27312 = ~n27309 & ~n27310;
  assign n27313 = ~n27308 & n27312;
  assign n27314 = ~n27311 & n27313;
  assign n27315 = pi29  & n27314;
  assign n27316 = ~pi29  & ~n27314;
  assign n27317 = ~n27315 & ~n27316;
  assign n27318 = n27307 & ~n27317;
  assign n27319 = ~n27307 & n27317;
  assign n27320 = ~n27318 & ~n27319;
  assign n27321 = ~n27276 & n27320;
  assign n27322 = n27276 & ~n27320;
  assign n27323 = ~n27321 & ~n27322;
  assign n27324 = n4721 & n20371;
  assign n27325 = n4691 & n20374;
  assign n27326 = n4515 & n20377;
  assign n27327 = n4516 & n22250;
  assign n27328 = ~n27325 & ~n27326;
  assign n27329 = ~n27324 & n27328;
  assign n27330 = ~n27327 & n27329;
  assign n27331 = pi26  & n27330;
  assign n27332 = ~pi26  & ~n27330;
  assign n27333 = ~n27331 & ~n27332;
  assign n27334 = n27323 & ~n27333;
  assign n27335 = ~n27323 & n27333;
  assign n27336 = ~n27334 & ~n27335;
  assign n27337 = n27275 & ~n27336;
  assign n27338 = ~n27275 & n27336;
  assign n27339 = ~n27337 & ~n27338;
  assign n27340 = n5267 & n20361;
  assign n27341 = n5185 & n20365;
  assign n27342 = n5121 & n20368;
  assign n27343 = n78 & n22848;
  assign n27344 = ~n27341 & ~n27342;
  assign n27345 = ~n27340 & n27344;
  assign n27346 = ~n27343 & n27345;
  assign n27347 = pi23  & n27346;
  assign n27348 = ~pi23  & ~n27346;
  assign n27349 = ~n27347 & ~n27348;
  assign n27350 = n27339 & ~n27349;
  assign n27351 = ~n27339 & n27349;
  assign n27352 = ~n27350 & ~n27351;
  assign n27353 = n27274 & ~n27352;
  assign n27354 = ~n27274 & n27352;
  assign n27355 = ~n27353 & ~n27354;
  assign n27356 = n5982 & n23394;
  assign n27357 = n5901 & n20355;
  assign n27358 = n5312 & n20358;
  assign n27359 = n5306 & n23404;
  assign n27360 = ~n27357 & ~n27358;
  assign n27361 = ~n27356 & n27360;
  assign n27362 = ~n27359 & n27361;
  assign n27363 = pi20  & n27362;
  assign n27364 = ~pi20  & ~n27362;
  assign n27365 = ~n27363 & ~n27364;
  assign n27366 = n27355 & ~n27365;
  assign n27367 = ~n27355 & n27365;
  assign n27368 = ~n27366 & ~n27367;
  assign n27369 = n27273 & ~n27368;
  assign n27370 = ~n27273 & n27368;
  assign n27371 = ~n27369 & ~n27370;
  assign n27372 = n6608 & n23765;
  assign n27373 = n6356 & n23768;
  assign n27374 = n6140 & n23771;
  assign n27375 = n6134 & n23789;
  assign n27376 = ~n27373 & ~n27374;
  assign n27377 = ~n27372 & n27376;
  assign n27378 = ~n27375 & n27377;
  assign n27379 = pi17  & n27378;
  assign n27380 = ~pi17  & ~n27378;
  assign n27381 = ~n27379 & ~n27380;
  assign n27382 = n27371 & ~n27381;
  assign n27383 = ~n27371 & n27381;
  assign n27384 = ~n27382 & ~n27383;
  assign n27385 = ~n27272 & n27384;
  assign n27386 = n27272 & ~n27384;
  assign n27387 = ~n27385 & ~n27386;
  assign n27388 = ~n27271 & n27387;
  assign n27389 = n27271 & ~n27387;
  assign n27390 = ~n27388 & ~n27389;
  assign n27391 = n27261 & ~n27390;
  assign n27392 = ~n27261 & n27390;
  assign n27393 = ~n27391 & ~n27392;
  assign n27394 = n8161 & n25709;
  assign n27395 = n7847 & n25490;
  assign n27396 = n7554 & n25253;
  assign n27397 = n7548 & n25719;
  assign n27398 = ~n27395 & ~n27396;
  assign n27399 = ~n27394 & n27398;
  assign n27400 = ~n27397 & n27399;
  assign n27401 = pi11  & n27400;
  assign n27402 = ~pi11  & ~n27400;
  assign n27403 = ~n27401 & ~n27402;
  assign n27404 = n27393 & ~n27403;
  assign n27405 = ~n27393 & n27403;
  assign n27406 = ~n27404 & ~n27405;
  assign n27407 = ~n27260 & n27406;
  assign n27408 = n27260 & ~n27406;
  assign n27409 = ~n27407 & ~n27408;
  assign n27410 = n27259 & ~n27409;
  assign n27411 = ~n27259 & n27409;
  assign n27412 = ~n27410 & ~n27411;
  assign n27413 = n27257 & n27412;
  assign n27414 = ~n27257 & ~n27412;
  assign po14  = ~n27413 & ~n27414;
  assign n27416 = ~n27392 & ~n27404;
  assign n27417 = ~n27385 & ~n27388;
  assign n27418 = ~n13357 & n25709;
  assign n27419 = n7554 & n25490;
  assign n27420 = n7548 & ~n25925;
  assign n27421 = ~n27418 & ~n27419;
  assign n27422 = ~n27420 & n27421;
  assign n27423 = pi11  & n27422;
  assign n27424 = ~pi11  & ~n27422;
  assign n27425 = ~n27423 & ~n27424;
  assign n27426 = ~n27417 & ~n27425;
  assign n27427 = n27417 & n27425;
  assign n27428 = ~n27426 & ~n27427;
  assign n27429 = ~n27370 & ~n27382;
  assign n27430 = ~n27354 & ~n27366;
  assign n27431 = ~n27338 & ~n27350;
  assign n27432 = ~n27321 & ~n27334;
  assign n27433 = ~n27306 & ~n27318;
  assign n27434 = n4472 & n20377;
  assign n27435 = n4070 & n20380;
  assign n27436 = n3943 & n20383;
  assign n27437 = n3944 & n22083;
  assign n27438 = ~n27435 & ~n27436;
  assign n27439 = ~n27434 & n27438;
  assign n27440 = ~n27437 & n27439;
  assign n27441 = pi29  & n27440;
  assign n27442 = ~pi29  & ~n27440;
  assign n27443 = ~n27441 & ~n27442;
  assign n27444 = ~n243 & ~n379;
  assign n27445 = ~n542 & n27444;
  assign n27446 = n1203 & n1561;
  assign n27447 = n1808 & n2063;
  assign n27448 = n2092 & n3352;
  assign n27449 = n27447 & n27448;
  assign n27450 = n14844 & n27446;
  assign n27451 = n1158 & n27445;
  assign n27452 = n3378 & n27451;
  assign n27453 = n27449 & n27450;
  assign n27454 = n27452 & n27453;
  assign n27455 = n12715 & n14167;
  assign n27456 = n27454 & n27455;
  assign n27457 = n5786 & n27456;
  assign n27458 = n26737 & n27457;
  assign n27459 = ~n27290 & n27458;
  assign n27460 = n27290 & ~n27458;
  assign n27461 = ~n27459 & ~n27460;
  assign n27462 = ~n27292 & ~n27302;
  assign n27463 = n27461 & n27462;
  assign n27464 = ~n27461 & ~n27462;
  assign n27465 = ~n27463 & ~n27464;
  assign n27466 = n3896 & n20386;
  assign n27467 = n3683 & n20389;
  assign n27468 = n564 & n20392;
  assign n27469 = n566 & n21752;
  assign n27470 = ~n27467 & ~n27468;
  assign n27471 = ~n27466 & n27470;
  assign n27472 = ~n27469 & n27471;
  assign n27473 = n27465 & ~n27472;
  assign n27474 = ~n27465 & n27472;
  assign n27475 = ~n27473 & ~n27474;
  assign n27476 = ~n27443 & n27475;
  assign n27477 = n27443 & ~n27475;
  assign n27478 = ~n27476 & ~n27477;
  assign n27479 = ~n27433 & n27478;
  assign n27480 = n27433 & ~n27478;
  assign n27481 = ~n27479 & ~n27480;
  assign n27482 = n4721 & n20368;
  assign n27483 = n4691 & n20371;
  assign n27484 = n4515 & n20374;
  assign n27485 = n4516 & n22235;
  assign n27486 = ~n27483 & ~n27484;
  assign n27487 = ~n27482 & n27486;
  assign n27488 = ~n27485 & n27487;
  assign n27489 = pi26  & n27488;
  assign n27490 = ~pi26  & ~n27488;
  assign n27491 = ~n27489 & ~n27490;
  assign n27492 = n27481 & ~n27491;
  assign n27493 = ~n27481 & n27491;
  assign n27494 = ~n27492 & ~n27493;
  assign n27495 = n27432 & ~n27494;
  assign n27496 = ~n27432 & n27494;
  assign n27497 = ~n27495 & ~n27496;
  assign n27498 = n5267 & n20358;
  assign n27499 = n5185 & n20361;
  assign n27500 = n5121 & n20365;
  assign n27501 = n78 & n22833;
  assign n27502 = ~n27499 & ~n27500;
  assign n27503 = ~n27498 & n27502;
  assign n27504 = ~n27501 & n27503;
  assign n27505 = pi23  & n27504;
  assign n27506 = ~pi23  & ~n27504;
  assign n27507 = ~n27505 & ~n27506;
  assign n27508 = n27497 & ~n27507;
  assign n27509 = ~n27497 & n27507;
  assign n27510 = ~n27508 & ~n27509;
  assign n27511 = n27431 & ~n27510;
  assign n27512 = ~n27431 & n27510;
  assign n27513 = ~n27511 & ~n27512;
  assign n27514 = n5982 & n23771;
  assign n27515 = n5901 & n23394;
  assign n27516 = n5312 & n20355;
  assign n27517 = n5306 & n23816;
  assign n27518 = ~n27515 & ~n27516;
  assign n27519 = ~n27514 & n27518;
  assign n27520 = ~n27517 & n27519;
  assign n27521 = pi20  & n27520;
  assign n27522 = ~pi20  & ~n27520;
  assign n27523 = ~n27521 & ~n27522;
  assign n27524 = n27513 & ~n27523;
  assign n27525 = ~n27513 & n27523;
  assign n27526 = ~n27524 & ~n27525;
  assign n27527 = n27430 & ~n27526;
  assign n27528 = ~n27430 & n27526;
  assign n27529 = ~n27527 & ~n27528;
  assign n27530 = n6608 & n24529;
  assign n27531 = n6356 & n23765;
  assign n27532 = n6140 & n23768;
  assign n27533 = n6134 & n24539;
  assign n27534 = ~n27531 & ~n27532;
  assign n27535 = ~n27530 & n27534;
  assign n27536 = ~n27533 & n27535;
  assign n27537 = pi17  & n27536;
  assign n27538 = ~pi17  & ~n27536;
  assign n27539 = ~n27537 & ~n27538;
  assign n27540 = n27529 & ~n27539;
  assign n27541 = ~n27529 & n27539;
  assign n27542 = ~n27540 & ~n27541;
  assign n27543 = n27429 & ~n27542;
  assign n27544 = ~n27429 & n27542;
  assign n27545 = ~n27543 & ~n27544;
  assign n27546 = n7380 & n25253;
  assign n27547 = n7243 & n25022;
  assign n27548 = n6653 & n24779;
  assign n27549 = n6647 & n25263;
  assign n27550 = ~n27547 & ~n27548;
  assign n27551 = ~n27546 & n27550;
  assign n27552 = ~n27549 & n27551;
  assign n27553 = pi14  & n27552;
  assign n27554 = ~pi14  & ~n27552;
  assign n27555 = ~n27553 & ~n27554;
  assign n27556 = n27545 & ~n27555;
  assign n27557 = ~n27545 & n27555;
  assign n27558 = ~n27556 & ~n27557;
  assign n27559 = n27428 & n27558;
  assign n27560 = ~n27428 & ~n27558;
  assign n27561 = ~n27559 & ~n27560;
  assign n27562 = n27416 & ~n27561;
  assign n27563 = ~n27416 & n27561;
  assign n27564 = ~n27562 & ~n27563;
  assign n27565 = ~n27407 & ~n27411;
  assign n27566 = ~n27564 & n27565;
  assign n27567 = n27564 & ~n27565;
  assign n27568 = ~n27566 & ~n27567;
  assign n27569 = n27413 & n27568;
  assign n27570 = ~n27413 & ~n27568;
  assign po15  = ~n27569 & ~n27570;
  assign n27572 = ~n27563 & ~n27567;
  assign n27573 = ~n27426 & ~n27559;
  assign n27574 = ~n27528 & ~n27540;
  assign n27575 = ~n27496 & ~n27508;
  assign n27576 = ~n27479 & ~n27492;
  assign n27577 = n4721 & n20365;
  assign n27578 = n4691 & n20368;
  assign n27579 = n4515 & n20371;
  assign n27580 = n4516 & n22814;
  assign n27581 = ~n27578 & ~n27579;
  assign n27582 = ~n27577 & n27581;
  assign n27583 = ~n27580 & n27582;
  assign n27584 = pi26  & n27583;
  assign n27585 = ~pi26  & ~n27583;
  assign n27586 = ~n27584 & ~n27585;
  assign n27587 = n4472 & n20374;
  assign n27588 = n4070 & n20377;
  assign n27589 = n3943 & n20380;
  assign n27590 = n3944 & n22263;
  assign n27591 = ~n27588 & ~n27589;
  assign n27592 = ~n27587 & n27591;
  assign n27593 = ~n27590 & n27592;
  assign n27594 = pi29  & n27593;
  assign n27595 = ~pi29  & ~n27593;
  assign n27596 = ~n27594 & ~n27595;
  assign n27597 = ~n27473 & ~n27476;
  assign n27598 = ~n27460 & ~n27463;
  assign n27599 = ~n13358 & n25709;
  assign n27600 = pi11  & ~n27599;
  assign n27601 = ~pi11  & n27599;
  assign n27602 = ~n27600 & ~n27601;
  assign n27603 = ~n134 & ~n405;
  assign n27604 = n573 & n27603;
  assign n27605 = n737 & n1113;
  assign n27606 = n1560 & n3271;
  assign n27607 = n3379 & n27606;
  assign n27608 = n27604 & n27605;
  assign n27609 = n5547 & n12486;
  assign n27610 = n27608 & n27609;
  assign n27611 = n2886 & n27607;
  assign n27612 = n5532 & n27611;
  assign n27613 = n27610 & n27612;
  assign n27614 = n2203 & n27613;
  assign n27615 = n1193 & n2251;
  assign n27616 = n27614 & n27615;
  assign n27617 = n27290 & n27616;
  assign n27618 = ~n27290 & ~n27616;
  assign n27619 = ~n27617 & ~n27618;
  assign n27620 = n27602 & n27619;
  assign n27621 = ~n27602 & ~n27619;
  assign n27622 = ~n27620 & ~n27621;
  assign n27623 = n3896 & n20383;
  assign n27624 = n3683 & n20386;
  assign n27625 = n564 & n20389;
  assign n27626 = n566 & n21737;
  assign n27627 = ~n27624 & ~n27625;
  assign n27628 = ~n27623 & n27627;
  assign n27629 = ~n27626 & n27628;
  assign n27630 = n27622 & ~n27629;
  assign n27631 = ~n27622 & n27629;
  assign n27632 = ~n27630 & ~n27631;
  assign n27633 = ~n27598 & n27632;
  assign n27634 = n27598 & ~n27632;
  assign n27635 = ~n27633 & ~n27634;
  assign n27636 = ~n27597 & n27635;
  assign n27637 = n27597 & ~n27635;
  assign n27638 = ~n27636 & ~n27637;
  assign n27639 = ~n27596 & n27638;
  assign n27640 = n27596 & ~n27638;
  assign n27641 = ~n27639 & ~n27640;
  assign n27642 = ~n27586 & n27641;
  assign n27643 = n27586 & ~n27641;
  assign n27644 = ~n27642 & ~n27643;
  assign n27645 = n27576 & ~n27644;
  assign n27646 = ~n27576 & n27644;
  assign n27647 = ~n27645 & ~n27646;
  assign n27648 = n5267 & n20355;
  assign n27649 = n5185 & n20358;
  assign n27650 = n5121 & n20361;
  assign n27651 = n78 & n20562;
  assign n27652 = ~n27649 & ~n27650;
  assign n27653 = ~n27648 & n27652;
  assign n27654 = ~n27651 & n27653;
  assign n27655 = pi23  & n27654;
  assign n27656 = ~pi23  & ~n27654;
  assign n27657 = ~n27655 & ~n27656;
  assign n27658 = n27647 & ~n27657;
  assign n27659 = ~n27647 & n27657;
  assign n27660 = ~n27658 & ~n27659;
  assign n27661 = n27575 & ~n27660;
  assign n27662 = ~n27575 & n27660;
  assign n27663 = ~n27661 & ~n27662;
  assign n27664 = ~n27512 & ~n27524;
  assign n27665 = n5982 & n23768;
  assign n27666 = n5901 & n23771;
  assign n27667 = n5312 & n23394;
  assign n27668 = n5306 & n23804;
  assign n27669 = ~n27666 & ~n27667;
  assign n27670 = ~n27665 & n27669;
  assign n27671 = ~n27668 & n27670;
  assign n27672 = pi20  & n27671;
  assign n27673 = ~pi20  & ~n27671;
  assign n27674 = ~n27672 & ~n27673;
  assign n27675 = ~n27664 & ~n27674;
  assign n27676 = n27664 & n27674;
  assign n27677 = ~n27675 & ~n27676;
  assign n27678 = ~n27663 & ~n27677;
  assign n27679 = n27663 & n27677;
  assign n27680 = ~n27678 & ~n27679;
  assign n27681 = n6608 & n24779;
  assign n27682 = n6356 & n24529;
  assign n27683 = n6140 & n23765;
  assign n27684 = n6134 & n24789;
  assign n27685 = ~n27682 & ~n27683;
  assign n27686 = ~n27681 & n27685;
  assign n27687 = ~n27684 & n27686;
  assign n27688 = pi17  & n27687;
  assign n27689 = ~pi17  & ~n27687;
  assign n27690 = ~n27688 & ~n27689;
  assign n27691 = n27680 & ~n27690;
  assign n27692 = ~n27680 & n27690;
  assign n27693 = ~n27691 & ~n27692;
  assign n27694 = n27574 & ~n27693;
  assign n27695 = ~n27574 & n27693;
  assign n27696 = ~n27694 & ~n27695;
  assign n27697 = ~n27544 & ~n27556;
  assign n27698 = n7380 & n25490;
  assign n27699 = n7243 & n25253;
  assign n27700 = n6653 & n25022;
  assign n27701 = n6647 & n25500;
  assign n27702 = ~n27699 & ~n27700;
  assign n27703 = ~n27698 & n27702;
  assign n27704 = ~n27701 & n27703;
  assign n27705 = pi14  & n27704;
  assign n27706 = ~pi14  & ~n27704;
  assign n27707 = ~n27705 & ~n27706;
  assign n27708 = ~n27697 & ~n27707;
  assign n27709 = n27697 & n27707;
  assign n27710 = ~n27708 & ~n27709;
  assign n27711 = ~n27696 & ~n27710;
  assign n27712 = n27696 & n27710;
  assign n27713 = ~n27711 & ~n27712;
  assign n27714 = ~n27573 & n27713;
  assign n27715 = n27573 & ~n27713;
  assign n27716 = ~n27714 & ~n27715;
  assign n27717 = ~n27572 & n27716;
  assign n27718 = n27572 & ~n27716;
  assign n27719 = ~n27717 & ~n27718;
  assign n27720 = ~n27569 & ~n27719;
  assign n27721 = n27569 & n27719;
  assign po16  = ~n27720 & ~n27721;
  assign n27723 = ~n27714 & ~n27717;
  assign n27724 = ~n27708 & ~n27712;
  assign n27725 = ~n27691 & ~n27695;
  assign n27726 = ~n27675 & ~n27679;
  assign n27727 = ~n27658 & ~n27662;
  assign n27728 = ~n27642 & ~n27646;
  assign n27729 = ~n27636 & ~n27639;
  assign n27730 = ~n27618 & ~n27620;
  assign n27731 = ~n662 & n919;
  assign n27732 = n1713 & n2234;
  assign n27733 = n2830 & n2925;
  assign n27734 = n3080 & n27733;
  assign n27735 = n27731 & n27732;
  assign n27736 = n669 & n2313;
  assign n27737 = n27735 & n27736;
  assign n27738 = n12539 & n27734;
  assign n27739 = n27737 & n27738;
  assign n27740 = n25349 & n25800;
  assign n27741 = n27739 & n27740;
  assign n27742 = n12496 & n27741;
  assign n27743 = n14179 & n27742;
  assign n27744 = ~n27730 & n27743;
  assign n27745 = n27730 & ~n27743;
  assign n27746 = ~n27744 & ~n27745;
  assign n27747 = n3896 & n20380;
  assign n27748 = n3683 & n20383;
  assign n27749 = n564 & n20386;
  assign n27750 = n566 & n20574;
  assign n27751 = ~n27748 & ~n27749;
  assign n27752 = ~n27747 & n27751;
  assign n27753 = ~n27750 & n27752;
  assign n27754 = ~n27746 & ~n27753;
  assign n27755 = n27746 & n27753;
  assign n27756 = ~n27754 & ~n27755;
  assign n27757 = ~n27630 & ~n27633;
  assign n27758 = n27756 & n27757;
  assign n27759 = ~n27756 & ~n27757;
  assign n27760 = ~n27758 & ~n27759;
  assign n27761 = n4472 & n20371;
  assign n27762 = n4070 & n20374;
  assign n27763 = n3943 & n20377;
  assign n27764 = n3944 & n22250;
  assign n27765 = ~n27762 & ~n27763;
  assign n27766 = ~n27761 & n27765;
  assign n27767 = ~n27764 & n27766;
  assign n27768 = pi29  & n27767;
  assign n27769 = ~pi29  & ~n27767;
  assign n27770 = ~n27768 & ~n27769;
  assign n27771 = n27760 & ~n27770;
  assign n27772 = ~n27760 & n27770;
  assign n27773 = ~n27771 & ~n27772;
  assign n27774 = ~n27729 & n27773;
  assign n27775 = n27729 & ~n27773;
  assign n27776 = ~n27774 & ~n27775;
  assign n27777 = n4721 & n20361;
  assign n27778 = n4691 & n20365;
  assign n27779 = n4515 & n20368;
  assign n27780 = n4516 & n22848;
  assign n27781 = ~n27778 & ~n27779;
  assign n27782 = ~n27777 & n27781;
  assign n27783 = ~n27780 & n27782;
  assign n27784 = pi26  & n27783;
  assign n27785 = ~pi26  & ~n27783;
  assign n27786 = ~n27784 & ~n27785;
  assign n27787 = n27776 & ~n27786;
  assign n27788 = ~n27776 & n27786;
  assign n27789 = ~n27787 & ~n27788;
  assign n27790 = n27728 & ~n27789;
  assign n27791 = ~n27728 & n27789;
  assign n27792 = ~n27790 & ~n27791;
  assign n27793 = n5267 & n23394;
  assign n27794 = n5185 & n20355;
  assign n27795 = n5121 & n20358;
  assign n27796 = n78 & n23404;
  assign n27797 = ~n27794 & ~n27795;
  assign n27798 = ~n27793 & n27797;
  assign n27799 = ~n27796 & n27798;
  assign n27800 = pi23  & n27799;
  assign n27801 = ~pi23  & ~n27799;
  assign n27802 = ~n27800 & ~n27801;
  assign n27803 = n27792 & ~n27802;
  assign n27804 = ~n27792 & n27802;
  assign n27805 = ~n27803 & ~n27804;
  assign n27806 = n27727 & ~n27805;
  assign n27807 = ~n27727 & n27805;
  assign n27808 = ~n27806 & ~n27807;
  assign n27809 = n5982 & n23765;
  assign n27810 = n5901 & n23768;
  assign n27811 = n5312 & n23771;
  assign n27812 = n5306 & n23789;
  assign n27813 = ~n27810 & ~n27811;
  assign n27814 = ~n27809 & n27813;
  assign n27815 = ~n27812 & n27814;
  assign n27816 = pi20  & n27815;
  assign n27817 = ~pi20  & ~n27815;
  assign n27818 = ~n27816 & ~n27817;
  assign n27819 = n27808 & ~n27818;
  assign n27820 = ~n27808 & n27818;
  assign n27821 = ~n27819 & ~n27820;
  assign n27822 = ~n27726 & n27821;
  assign n27823 = n27726 & ~n27821;
  assign n27824 = ~n27822 & ~n27823;
  assign n27825 = n6608 & n25022;
  assign n27826 = n6356 & n24779;
  assign n27827 = n6140 & n24529;
  assign n27828 = n6134 & n25032;
  assign n27829 = ~n27826 & ~n27827;
  assign n27830 = ~n27825 & n27829;
  assign n27831 = ~n27828 & n27830;
  assign n27832 = pi17  & n27831;
  assign n27833 = ~pi17  & ~n27831;
  assign n27834 = ~n27832 & ~n27833;
  assign n27835 = n27824 & ~n27834;
  assign n27836 = ~n27824 & n27834;
  assign n27837 = ~n27835 & ~n27836;
  assign n27838 = n27725 & ~n27837;
  assign n27839 = ~n27725 & n27837;
  assign n27840 = ~n27838 & ~n27839;
  assign n27841 = n7380 & n25709;
  assign n27842 = n7243 & n25490;
  assign n27843 = n6653 & n25253;
  assign n27844 = n6647 & n25719;
  assign n27845 = ~n27842 & ~n27843;
  assign n27846 = ~n27841 & n27845;
  assign n27847 = ~n27844 & n27846;
  assign n27848 = pi14  & n27847;
  assign n27849 = ~pi14  & ~n27847;
  assign n27850 = ~n27848 & ~n27849;
  assign n27851 = n27840 & ~n27850;
  assign n27852 = ~n27840 & n27850;
  assign n27853 = ~n27851 & ~n27852;
  assign n27854 = ~n27724 & n27853;
  assign n27855 = n27724 & ~n27853;
  assign n27856 = ~n27854 & ~n27855;
  assign n27857 = n27723 & ~n27856;
  assign n27858 = ~n27723 & n27856;
  assign n27859 = ~n27857 & ~n27858;
  assign n27860 = n27721 & n27859;
  assign n27861 = ~n27721 & ~n27859;
  assign po17  = ~n27860 & ~n27861;
  assign n27863 = ~n27839 & ~n27851;
  assign n27864 = ~n27822 & ~n27835;
  assign n27865 = ~n12787 & n25709;
  assign n27866 = n6653 & n25490;
  assign n27867 = n6647 & ~n25925;
  assign n27868 = ~n27865 & ~n27866;
  assign n27869 = ~n27867 & n27868;
  assign n27870 = pi14  & n27869;
  assign n27871 = ~pi14  & ~n27869;
  assign n27872 = ~n27870 & ~n27871;
  assign n27873 = ~n27864 & ~n27872;
  assign n27874 = n27864 & n27872;
  assign n27875 = ~n27873 & ~n27874;
  assign n27876 = ~n27807 & ~n27819;
  assign n27877 = ~n27791 & ~n27803;
  assign n27878 = ~n27774 & ~n27787;
  assign n27879 = n4721 & n20358;
  assign n27880 = n4691 & n20361;
  assign n27881 = n4515 & n20365;
  assign n27882 = n4516 & n22833;
  assign n27883 = ~n27880 & ~n27881;
  assign n27884 = ~n27879 & n27883;
  assign n27885 = ~n27882 & n27884;
  assign n27886 = pi26  & n27885;
  assign n27887 = ~pi26  & ~n27885;
  assign n27888 = ~n27886 & ~n27887;
  assign n27889 = ~n125 & ~n288;
  assign n27890 = ~n334 & ~n381;
  assign n27891 = ~n387 & ~n425;
  assign n27892 = ~n673 & ~n687;
  assign n27893 = n27891 & n27892;
  assign n27894 = n27889 & n27890;
  assign n27895 = n281 & n1593;
  assign n27896 = n3855 & n27895;
  assign n27897 = n27893 & n27894;
  assign n27898 = n27896 & n27897;
  assign n27899 = n2888 & n3769;
  assign n27900 = n27898 & n27899;
  assign n27901 = n952 & n3636;
  assign n27902 = n5696 & n27901;
  assign n27903 = n3153 & n27900;
  assign n27904 = n27902 & n27903;
  assign n27905 = n4324 & n27904;
  assign n27906 = ~n27743 & n27905;
  assign n27907 = n27743 & ~n27905;
  assign n27908 = ~n27906 & ~n27907;
  assign n27909 = n3896 & n20377;
  assign n27910 = n3683 & n20380;
  assign n27911 = n564 & n20383;
  assign n27912 = n566 & n22083;
  assign n27913 = ~n27910 & ~n27911;
  assign n27914 = ~n27909 & n27913;
  assign n27915 = ~n27912 & n27914;
  assign n27916 = n27908 & ~n27915;
  assign n27917 = ~n27908 & n27915;
  assign n27918 = ~n27916 & ~n27917;
  assign n27919 = ~n27745 & ~n27755;
  assign n27920 = ~n27918 & ~n27919;
  assign n27921 = n27918 & n27919;
  assign n27922 = ~n27920 & ~n27921;
  assign n27923 = ~n27759 & ~n27771;
  assign n27924 = ~n27922 & n27923;
  assign n27925 = n27922 & ~n27923;
  assign n27926 = ~n27924 & ~n27925;
  assign n27927 = n4472 & n20368;
  assign n27928 = n4070 & n20371;
  assign n27929 = n3943 & n20374;
  assign n27930 = n3944 & n22235;
  assign n27931 = ~n27928 & ~n27929;
  assign n27932 = ~n27927 & n27931;
  assign n27933 = ~n27930 & n27932;
  assign n27934 = pi29  & n27933;
  assign n27935 = ~pi29  & ~n27933;
  assign n27936 = ~n27934 & ~n27935;
  assign n27937 = n27926 & ~n27936;
  assign n27938 = ~n27926 & n27936;
  assign n27939 = ~n27937 & ~n27938;
  assign n27940 = ~n27888 & n27939;
  assign n27941 = n27888 & ~n27939;
  assign n27942 = ~n27940 & ~n27941;
  assign n27943 = n27878 & ~n27942;
  assign n27944 = ~n27878 & n27942;
  assign n27945 = ~n27943 & ~n27944;
  assign n27946 = n5267 & n23771;
  assign n27947 = n5185 & n23394;
  assign n27948 = n5121 & n20355;
  assign n27949 = n78 & n23816;
  assign n27950 = ~n27947 & ~n27948;
  assign n27951 = ~n27946 & n27950;
  assign n27952 = ~n27949 & n27951;
  assign n27953 = pi23  & n27952;
  assign n27954 = ~pi23  & ~n27952;
  assign n27955 = ~n27953 & ~n27954;
  assign n27956 = n27945 & ~n27955;
  assign n27957 = ~n27945 & n27955;
  assign n27958 = ~n27956 & ~n27957;
  assign n27959 = n27877 & ~n27958;
  assign n27960 = ~n27877 & n27958;
  assign n27961 = ~n27959 & ~n27960;
  assign n27962 = n5982 & n24529;
  assign n27963 = n5901 & n23765;
  assign n27964 = n5312 & n23768;
  assign n27965 = n5306 & n24539;
  assign n27966 = ~n27963 & ~n27964;
  assign n27967 = ~n27962 & n27966;
  assign n27968 = ~n27965 & n27967;
  assign n27969 = pi20  & n27968;
  assign n27970 = ~pi20  & ~n27968;
  assign n27971 = ~n27969 & ~n27970;
  assign n27972 = n27961 & ~n27971;
  assign n27973 = ~n27961 & n27971;
  assign n27974 = ~n27972 & ~n27973;
  assign n27975 = n27876 & ~n27974;
  assign n27976 = ~n27876 & n27974;
  assign n27977 = ~n27975 & ~n27976;
  assign n27978 = n6608 & n25253;
  assign n27979 = n6356 & n25022;
  assign n27980 = n6140 & n24779;
  assign n27981 = n6134 & n25263;
  assign n27982 = ~n27979 & ~n27980;
  assign n27983 = ~n27978 & n27982;
  assign n27984 = ~n27981 & n27983;
  assign n27985 = pi17  & n27984;
  assign n27986 = ~pi17  & ~n27984;
  assign n27987 = ~n27985 & ~n27986;
  assign n27988 = n27977 & ~n27987;
  assign n27989 = ~n27977 & n27987;
  assign n27990 = ~n27988 & ~n27989;
  assign n27991 = n27875 & n27990;
  assign n27992 = ~n27875 & ~n27990;
  assign n27993 = ~n27991 & ~n27992;
  assign n27994 = n27863 & ~n27993;
  assign n27995 = ~n27863 & n27993;
  assign n27996 = ~n27994 & ~n27995;
  assign n27997 = ~n27854 & ~n27858;
  assign n27998 = ~n27996 & n27997;
  assign n27999 = n27996 & ~n27997;
  assign n28000 = ~n27998 & ~n27999;
  assign n28001 = n27860 & n28000;
  assign n28002 = ~n27860 & ~n28000;
  assign po18  = ~n28001 & ~n28002;
  assign n28004 = ~n27995 & ~n27999;
  assign n28005 = ~n27873 & ~n27991;
  assign n28006 = ~n27960 & ~n27972;
  assign n28007 = ~n27937 & ~n27940;
  assign n28008 = ~n27921 & ~n27925;
  assign n28009 = ~n27907 & ~n27916;
  assign n28010 = ~n12788 & n25709;
  assign n28011 = pi14  & ~n28010;
  assign n28012 = ~pi14  & n28010;
  assign n28013 = ~n28011 & ~n28012;
  assign n28014 = ~n536 & ~n683;
  assign n28015 = n1306 & n28014;
  assign n28016 = n1265 & n28015;
  assign n28017 = n3197 & n4273;
  assign n28018 = n13881 & n28017;
  assign n28019 = n13409 & n28016;
  assign n28020 = n28018 & n28019;
  assign n28021 = n1880 & n7067;
  assign n28022 = n28020 & n28021;
  assign n28023 = n13153 & n28022;
  assign n28024 = n2128 & n28023;
  assign n28025 = n27743 & n28024;
  assign n28026 = ~n27743 & ~n28024;
  assign n28027 = ~n28025 & ~n28026;
  assign n28028 = n28013 & n28027;
  assign n28029 = ~n28013 & ~n28027;
  assign n28030 = ~n28028 & ~n28029;
  assign n28031 = ~n28009 & n28030;
  assign n28032 = n28009 & ~n28030;
  assign n28033 = ~n28031 & ~n28032;
  assign n28034 = n3896 & n20374;
  assign n28035 = n3683 & n20377;
  assign n28036 = n564 & n20380;
  assign n28037 = n566 & n22263;
  assign n28038 = ~n28035 & ~n28036;
  assign n28039 = ~n28034 & n28038;
  assign n28040 = ~n28037 & n28039;
  assign n28041 = n28033 & n28040;
  assign n28042 = ~n28033 & ~n28040;
  assign n28043 = ~n28041 & ~n28042;
  assign n28044 = n4472 & n20365;
  assign n28045 = n4070 & n20368;
  assign n28046 = n3943 & n20371;
  assign n28047 = n3944 & n22814;
  assign n28048 = ~n28045 & ~n28046;
  assign n28049 = ~n28044 & n28048;
  assign n28050 = ~n28047 & n28049;
  assign n28051 = pi29  & n28050;
  assign n28052 = ~pi29  & ~n28050;
  assign n28053 = ~n28051 & ~n28052;
  assign n28054 = ~n28043 & ~n28053;
  assign n28055 = n28043 & n28053;
  assign n28056 = ~n28054 & ~n28055;
  assign n28057 = n28008 & ~n28056;
  assign n28058 = ~n28008 & n28056;
  assign n28059 = ~n28057 & ~n28058;
  assign n28060 = n4721 & n20355;
  assign n28061 = n4691 & n20358;
  assign n28062 = n4515 & n20361;
  assign n28063 = n4516 & n20562;
  assign n28064 = ~n28061 & ~n28062;
  assign n28065 = ~n28060 & n28064;
  assign n28066 = ~n28063 & n28065;
  assign n28067 = pi26  & n28066;
  assign n28068 = ~pi26  & ~n28066;
  assign n28069 = ~n28067 & ~n28068;
  assign n28070 = n28059 & ~n28069;
  assign n28071 = ~n28059 & n28069;
  assign n28072 = ~n28070 & ~n28071;
  assign n28073 = n28007 & ~n28072;
  assign n28074 = ~n28007 & n28072;
  assign n28075 = ~n28073 & ~n28074;
  assign n28076 = ~n27944 & ~n27956;
  assign n28077 = n5267 & n23768;
  assign n28078 = n5185 & n23771;
  assign n28079 = n5121 & n23394;
  assign n28080 = n78 & n23804;
  assign n28081 = ~n28078 & ~n28079;
  assign n28082 = ~n28077 & n28081;
  assign n28083 = ~n28080 & n28082;
  assign n28084 = pi23  & n28083;
  assign n28085 = ~pi23  & ~n28083;
  assign n28086 = ~n28084 & ~n28085;
  assign n28087 = ~n28076 & ~n28086;
  assign n28088 = n28076 & n28086;
  assign n28089 = ~n28087 & ~n28088;
  assign n28090 = ~n28075 & ~n28089;
  assign n28091 = n28075 & n28089;
  assign n28092 = ~n28090 & ~n28091;
  assign n28093 = n5982 & n24779;
  assign n28094 = n5901 & n24529;
  assign n28095 = n5312 & n23765;
  assign n28096 = n5306 & n24789;
  assign n28097 = ~n28094 & ~n28095;
  assign n28098 = ~n28093 & n28097;
  assign n28099 = ~n28096 & n28098;
  assign n28100 = pi20  & n28099;
  assign n28101 = ~pi20  & ~n28099;
  assign n28102 = ~n28100 & ~n28101;
  assign n28103 = n28092 & ~n28102;
  assign n28104 = ~n28092 & n28102;
  assign n28105 = ~n28103 & ~n28104;
  assign n28106 = n28006 & ~n28105;
  assign n28107 = ~n28006 & n28105;
  assign n28108 = ~n28106 & ~n28107;
  assign n28109 = ~n27976 & ~n27988;
  assign n28110 = n6608 & n25490;
  assign n28111 = n6356 & n25253;
  assign n28112 = n6140 & n25022;
  assign n28113 = n6134 & n25500;
  assign n28114 = ~n28111 & ~n28112;
  assign n28115 = ~n28110 & n28114;
  assign n28116 = ~n28113 & n28115;
  assign n28117 = pi17  & n28116;
  assign n28118 = ~pi17  & ~n28116;
  assign n28119 = ~n28117 & ~n28118;
  assign n28120 = ~n28109 & ~n28119;
  assign n28121 = n28109 & n28119;
  assign n28122 = ~n28120 & ~n28121;
  assign n28123 = ~n28108 & ~n28122;
  assign n28124 = n28108 & n28122;
  assign n28125 = ~n28123 & ~n28124;
  assign n28126 = ~n28005 & n28125;
  assign n28127 = n28005 & ~n28125;
  assign n28128 = ~n28126 & ~n28127;
  assign n28129 = ~n28004 & n28128;
  assign n28130 = n28004 & ~n28128;
  assign n28131 = ~n28129 & ~n28130;
  assign n28132 = ~n28001 & ~n28131;
  assign n28133 = n28001 & n28131;
  assign po19  = ~n28132 & ~n28133;
  assign n28135 = ~n28126 & ~n28129;
  assign n28136 = ~n28120 & ~n28124;
  assign n28137 = ~n28103 & ~n28107;
  assign n28138 = n5982 & n25022;
  assign n28139 = n5901 & n24779;
  assign n28140 = n5312 & n24529;
  assign n28141 = n5306 & n25032;
  assign n28142 = ~n28139 & ~n28140;
  assign n28143 = ~n28138 & n28142;
  assign n28144 = ~n28141 & n28143;
  assign n28145 = pi20  & n28144;
  assign n28146 = ~pi20  & ~n28144;
  assign n28147 = ~n28145 & ~n28146;
  assign n28148 = ~n28087 & ~n28091;
  assign n28149 = ~n28070 & ~n28074;
  assign n28150 = ~n28054 & ~n28058;
  assign n28151 = ~n28026 & ~n28028;
  assign n28152 = ~n466 & ~n601;
  assign n28153 = n166 & n28152;
  assign n28154 = n524 & n904;
  assign n28155 = n923 & n1868;
  assign n28156 = n2008 & n2599;
  assign n28157 = n14801 & n28156;
  assign n28158 = n28154 & n28155;
  assign n28159 = n2169 & n28153;
  assign n28160 = n28158 & n28159;
  assign n28161 = n945 & n28157;
  assign n28162 = n28160 & n28161;
  assign n28163 = n6225 & n13458;
  assign n28164 = n28162 & n28163;
  assign n28165 = n5543 & n28164;
  assign n28166 = n3340 & n28165;
  assign n28167 = ~n28151 & n28166;
  assign n28168 = n28151 & ~n28166;
  assign n28169 = ~n28167 & ~n28168;
  assign n28170 = n3896 & n20371;
  assign n28171 = n3683 & n20374;
  assign n28172 = n564 & n20377;
  assign n28173 = n566 & n22250;
  assign n28174 = ~n28171 & ~n28172;
  assign n28175 = ~n28170 & n28174;
  assign n28176 = ~n28173 & n28175;
  assign n28177 = ~n28169 & ~n28176;
  assign n28178 = n28169 & n28176;
  assign n28179 = ~n28177 & ~n28178;
  assign n28180 = ~n28032 & ~n28041;
  assign n28181 = n28179 & ~n28180;
  assign n28182 = ~n28179 & n28180;
  assign n28183 = ~n28181 & ~n28182;
  assign n28184 = n4472 & n20361;
  assign n28185 = n4070 & n20365;
  assign n28186 = n3943 & n20368;
  assign n28187 = n3944 & n22848;
  assign n28188 = ~n28185 & ~n28186;
  assign n28189 = ~n28184 & n28188;
  assign n28190 = ~n28187 & n28189;
  assign n28191 = pi29  & n28190;
  assign n28192 = ~pi29  & ~n28190;
  assign n28193 = ~n28191 & ~n28192;
  assign n28194 = n28183 & ~n28193;
  assign n28195 = ~n28183 & n28193;
  assign n28196 = ~n28194 & ~n28195;
  assign n28197 = ~n28150 & n28196;
  assign n28198 = n28150 & ~n28196;
  assign n28199 = ~n28197 & ~n28198;
  assign n28200 = n4721 & n23394;
  assign n28201 = n4691 & n20355;
  assign n28202 = n4515 & n20358;
  assign n28203 = n4516 & n23404;
  assign n28204 = ~n28201 & ~n28202;
  assign n28205 = ~n28200 & n28204;
  assign n28206 = ~n28203 & n28205;
  assign n28207 = pi26  & n28206;
  assign n28208 = ~pi26  & ~n28206;
  assign n28209 = ~n28207 & ~n28208;
  assign n28210 = n28199 & ~n28209;
  assign n28211 = ~n28199 & n28209;
  assign n28212 = ~n28210 & ~n28211;
  assign n28213 = n28149 & ~n28212;
  assign n28214 = ~n28149 & n28212;
  assign n28215 = ~n28213 & ~n28214;
  assign n28216 = n5267 & n23765;
  assign n28217 = n5185 & n23768;
  assign n28218 = n5121 & n23771;
  assign n28219 = n78 & n23789;
  assign n28220 = ~n28217 & ~n28218;
  assign n28221 = ~n28216 & n28220;
  assign n28222 = ~n28219 & n28221;
  assign n28223 = pi23  & n28222;
  assign n28224 = ~pi23  & ~n28222;
  assign n28225 = ~n28223 & ~n28224;
  assign n28226 = n28215 & ~n28225;
  assign n28227 = ~n28215 & n28225;
  assign n28228 = ~n28226 & ~n28227;
  assign n28229 = ~n28148 & n28228;
  assign n28230 = n28148 & ~n28228;
  assign n28231 = ~n28229 & ~n28230;
  assign n28232 = ~n28147 & n28231;
  assign n28233 = n28147 & ~n28231;
  assign n28234 = ~n28232 & ~n28233;
  assign n28235 = n28137 & ~n28234;
  assign n28236 = ~n28137 & n28234;
  assign n28237 = ~n28235 & ~n28236;
  assign n28238 = n6608 & n25709;
  assign n28239 = n6356 & n25490;
  assign n28240 = n6140 & n25253;
  assign n28241 = n6134 & n25719;
  assign n28242 = ~n28239 & ~n28240;
  assign n28243 = ~n28238 & n28242;
  assign n28244 = ~n28241 & n28243;
  assign n28245 = pi17  & n28244;
  assign n28246 = ~pi17  & ~n28244;
  assign n28247 = ~n28245 & ~n28246;
  assign n28248 = n28237 & ~n28247;
  assign n28249 = ~n28237 & n28247;
  assign n28250 = ~n28248 & ~n28249;
  assign n28251 = ~n28136 & n28250;
  assign n28252 = n28136 & ~n28250;
  assign n28253 = ~n28251 & ~n28252;
  assign n28254 = n28135 & ~n28253;
  assign n28255 = ~n28135 & n28253;
  assign n28256 = ~n28254 & ~n28255;
  assign n28257 = n28133 & n28256;
  assign n28258 = ~n28133 & ~n28256;
  assign po20  = ~n28257 & ~n28258;
  assign n28260 = ~n28236 & ~n28248;
  assign n28261 = ~n28229 & ~n28232;
  assign n28262 = ~n12666 & n25709;
  assign n28263 = n6140 & n25490;
  assign n28264 = n6134 & ~n25925;
  assign n28265 = ~n28262 & ~n28263;
  assign n28266 = ~n28264 & n28265;
  assign n28267 = pi17  & n28266;
  assign n28268 = ~pi17  & ~n28266;
  assign n28269 = ~n28267 & ~n28268;
  assign n28270 = ~n28261 & ~n28269;
  assign n28271 = n28261 & n28269;
  assign n28272 = ~n28270 & ~n28271;
  assign n28273 = ~n28214 & ~n28226;
  assign n28274 = ~n28197 & ~n28210;
  assign n28275 = ~n28182 & ~n28194;
  assign n28276 = n4472 & n20358;
  assign n28277 = n4070 & n20361;
  assign n28278 = n3943 & n20365;
  assign n28279 = n3944 & n22833;
  assign n28280 = ~n28277 & ~n28278;
  assign n28281 = ~n28276 & n28280;
  assign n28282 = ~n28279 & n28281;
  assign n28283 = pi29  & n28282;
  assign n28284 = ~pi29  & ~n28282;
  assign n28285 = ~n28283 & ~n28284;
  assign n28286 = ~n405 & n14753;
  assign n28287 = ~n144 & ~n422;
  assign n28288 = ~n482 & ~n650;
  assign n28289 = n28287 & n28288;
  assign n28290 = n237 & n1242;
  assign n28291 = n1374 & n1465;
  assign n28292 = n2234 & n2737;
  assign n28293 = n28291 & n28292;
  assign n28294 = n28289 & n28290;
  assign n28295 = n28293 & n28294;
  assign n28296 = n847 & n3176;
  assign n28297 = n28286 & n28296;
  assign n28298 = n28295 & n28297;
  assign n28299 = n3838 & n28298;
  assign n28300 = n1941 & n5737;
  assign n28301 = n28299 & n28300;
  assign n28302 = n28166 & ~n28301;
  assign n28303 = ~n28166 & n28301;
  assign n28304 = ~n28302 & ~n28303;
  assign n28305 = ~n28168 & ~n28178;
  assign n28306 = n28304 & n28305;
  assign n28307 = ~n28304 & ~n28305;
  assign n28308 = ~n28306 & ~n28307;
  assign n28309 = n3896 & n20368;
  assign n28310 = n3683 & n20371;
  assign n28311 = n564 & n20374;
  assign n28312 = n566 & n22235;
  assign n28313 = ~n28310 & ~n28311;
  assign n28314 = ~n28309 & n28313;
  assign n28315 = ~n28312 & n28314;
  assign n28316 = n28308 & ~n28315;
  assign n28317 = ~n28308 & n28315;
  assign n28318 = ~n28316 & ~n28317;
  assign n28319 = ~n28285 & n28318;
  assign n28320 = n28285 & ~n28318;
  assign n28321 = ~n28319 & ~n28320;
  assign n28322 = ~n28275 & n28321;
  assign n28323 = n28275 & ~n28321;
  assign n28324 = ~n28322 & ~n28323;
  assign n28325 = n4721 & n23771;
  assign n28326 = n4691 & n23394;
  assign n28327 = n4515 & n20355;
  assign n28328 = n4516 & n23816;
  assign n28329 = ~n28326 & ~n28327;
  assign n28330 = ~n28325 & n28329;
  assign n28331 = ~n28328 & n28330;
  assign n28332 = pi26  & n28331;
  assign n28333 = ~pi26  & ~n28331;
  assign n28334 = ~n28332 & ~n28333;
  assign n28335 = n28324 & ~n28334;
  assign n28336 = ~n28324 & n28334;
  assign n28337 = ~n28335 & ~n28336;
  assign n28338 = n28274 & ~n28337;
  assign n28339 = ~n28274 & n28337;
  assign n28340 = ~n28338 & ~n28339;
  assign n28341 = n5267 & n24529;
  assign n28342 = n5185 & n23765;
  assign n28343 = n5121 & n23768;
  assign n28344 = n78 & n24539;
  assign n28345 = ~n28342 & ~n28343;
  assign n28346 = ~n28341 & n28345;
  assign n28347 = ~n28344 & n28346;
  assign n28348 = pi23  & n28347;
  assign n28349 = ~pi23  & ~n28347;
  assign n28350 = ~n28348 & ~n28349;
  assign n28351 = n28340 & ~n28350;
  assign n28352 = ~n28340 & n28350;
  assign n28353 = ~n28351 & ~n28352;
  assign n28354 = n28273 & ~n28353;
  assign n28355 = ~n28273 & n28353;
  assign n28356 = ~n28354 & ~n28355;
  assign n28357 = n5982 & n25253;
  assign n28358 = n5901 & n25022;
  assign n28359 = n5312 & n24779;
  assign n28360 = n5306 & n25263;
  assign n28361 = ~n28358 & ~n28359;
  assign n28362 = ~n28357 & n28361;
  assign n28363 = ~n28360 & n28362;
  assign n28364 = pi20  & n28363;
  assign n28365 = ~pi20  & ~n28363;
  assign n28366 = ~n28364 & ~n28365;
  assign n28367 = n28356 & ~n28366;
  assign n28368 = ~n28356 & n28366;
  assign n28369 = ~n28367 & ~n28368;
  assign n28370 = n28272 & n28369;
  assign n28371 = ~n28272 & ~n28369;
  assign n28372 = ~n28370 & ~n28371;
  assign n28373 = n28260 & ~n28372;
  assign n28374 = ~n28260 & n28372;
  assign n28375 = ~n28373 & ~n28374;
  assign n28376 = ~n28251 & ~n28255;
  assign n28377 = ~n28375 & n28376;
  assign n28378 = n28375 & ~n28376;
  assign n28379 = ~n28377 & ~n28378;
  assign n28380 = n28257 & n28379;
  assign n28381 = ~n28257 & ~n28379;
  assign po21  = ~n28380 & ~n28381;
  assign n28383 = ~n28374 & ~n28378;
  assign n28384 = ~n28270 & ~n28370;
  assign n28385 = ~n28339 & ~n28351;
  assign n28386 = n5267 & n24779;
  assign n28387 = n5185 & n24529;
  assign n28388 = n5121 & n23765;
  assign n28389 = n78 & n24789;
  assign n28390 = ~n28387 & ~n28388;
  assign n28391 = ~n28386 & n28390;
  assign n28392 = ~n28389 & n28391;
  assign n28393 = pi23  & n28392;
  assign n28394 = ~pi23  & ~n28392;
  assign n28395 = ~n28393 & ~n28394;
  assign n28396 = n4472 & n20355;
  assign n28397 = n4070 & n20358;
  assign n28398 = n3943 & n20361;
  assign n28399 = n3944 & n20562;
  assign n28400 = ~n28397 & ~n28398;
  assign n28401 = ~n28396 & n28400;
  assign n28402 = ~n28399 & n28401;
  assign n28403 = pi29  & n28402;
  assign n28404 = ~pi29  & ~n28402;
  assign n28405 = ~n28403 & ~n28404;
  assign n28406 = ~n28316 & ~n28319;
  assign n28407 = ~n28303 & ~n28306;
  assign n28408 = ~n12667 & n25709;
  assign n28409 = pi17  & ~n28408;
  assign n28410 = ~pi17  & n28408;
  assign n28411 = ~n28409 & ~n28410;
  assign n28412 = ~n144 & ~n356;
  assign n28413 = ~n407 & n28412;
  assign n28414 = n1355 & n1739;
  assign n28415 = n28413 & n28414;
  assign n28416 = n1972 & n22709;
  assign n28417 = n28415 & n28416;
  assign n28418 = n1789 & n3349;
  assign n28419 = n12437 & n28418;
  assign n28420 = n28417 & n28419;
  assign n28421 = n1484 & n28420;
  assign n28422 = n4604 & n5356;
  assign n28423 = n28421 & n28422;
  assign n28424 = n28301 & n28423;
  assign n28425 = ~n28301 & ~n28423;
  assign n28426 = ~n28424 & ~n28425;
  assign n28427 = n28411 & n28426;
  assign n28428 = ~n28411 & ~n28426;
  assign n28429 = ~n28427 & ~n28428;
  assign n28430 = n3896 & n20365;
  assign n28431 = n3683 & n20368;
  assign n28432 = n564 & n20371;
  assign n28433 = n566 & n22814;
  assign n28434 = ~n28431 & ~n28432;
  assign n28435 = ~n28430 & n28434;
  assign n28436 = ~n28433 & n28435;
  assign n28437 = n28429 & ~n28436;
  assign n28438 = ~n28429 & n28436;
  assign n28439 = ~n28437 & ~n28438;
  assign n28440 = ~n28407 & n28439;
  assign n28441 = n28407 & ~n28439;
  assign n28442 = ~n28440 & ~n28441;
  assign n28443 = ~n28406 & n28442;
  assign n28444 = n28406 & ~n28442;
  assign n28445 = ~n28443 & ~n28444;
  assign n28446 = ~n28405 & n28445;
  assign n28447 = n28405 & ~n28445;
  assign n28448 = ~n28446 & ~n28447;
  assign n28449 = ~n28322 & ~n28335;
  assign n28450 = n4721 & n23768;
  assign n28451 = n4691 & n23771;
  assign n28452 = n4515 & n23394;
  assign n28453 = n4516 & n23804;
  assign n28454 = ~n28451 & ~n28452;
  assign n28455 = ~n28450 & n28454;
  assign n28456 = ~n28453 & n28455;
  assign n28457 = pi26  & n28456;
  assign n28458 = ~pi26  & ~n28456;
  assign n28459 = ~n28457 & ~n28458;
  assign n28460 = ~n28449 & ~n28459;
  assign n28461 = n28449 & n28459;
  assign n28462 = ~n28460 & ~n28461;
  assign n28463 = n28448 & n28462;
  assign n28464 = ~n28448 & ~n28462;
  assign n28465 = ~n28463 & ~n28464;
  assign n28466 = ~n28395 & n28465;
  assign n28467 = n28395 & ~n28465;
  assign n28468 = ~n28466 & ~n28467;
  assign n28469 = n28385 & ~n28468;
  assign n28470 = ~n28385 & n28468;
  assign n28471 = ~n28469 & ~n28470;
  assign n28472 = ~n28355 & ~n28367;
  assign n28473 = n5982 & n25490;
  assign n28474 = n5901 & n25253;
  assign n28475 = n5312 & n25022;
  assign n28476 = n5306 & n25500;
  assign n28477 = ~n28474 & ~n28475;
  assign n28478 = ~n28473 & n28477;
  assign n28479 = ~n28476 & n28478;
  assign n28480 = pi20  & n28479;
  assign n28481 = ~pi20  & ~n28479;
  assign n28482 = ~n28480 & ~n28481;
  assign n28483 = ~n28472 & ~n28482;
  assign n28484 = n28472 & n28482;
  assign n28485 = ~n28483 & ~n28484;
  assign n28486 = ~n28471 & ~n28485;
  assign n28487 = n28471 & n28485;
  assign n28488 = ~n28486 & ~n28487;
  assign n28489 = ~n28384 & n28488;
  assign n28490 = n28384 & ~n28488;
  assign n28491 = ~n28489 & ~n28490;
  assign n28492 = ~n28383 & n28491;
  assign n28493 = n28383 & ~n28491;
  assign n28494 = ~n28492 & ~n28493;
  assign n28495 = ~n28380 & ~n28494;
  assign n28496 = n28380 & n28494;
  assign po22  = ~n28495 & ~n28496;
  assign n28498 = ~n28489 & ~n28492;
  assign n28499 = ~n28483 & ~n28487;
  assign n28500 = ~n28466 & ~n28470;
  assign n28501 = ~n28460 & ~n28463;
  assign n28502 = ~n28443 & ~n28446;
  assign n28503 = ~n28425 & ~n28427;
  assign n28504 = ~n118 & ~n139;
  assign n28505 = ~n277 & ~n388;
  assign n28506 = ~n602 & ~n683;
  assign n28507 = n28505 & n28506;
  assign n28508 = n1121 & n28504;
  assign n28509 = n1469 & n1534;
  assign n28510 = n4767 & n28509;
  assign n28511 = n28507 & n28508;
  assign n28512 = n3256 & n12126;
  assign n28513 = n28511 & n28512;
  assign n28514 = n28510 & n28513;
  assign n28515 = n1182 & n3202;
  assign n28516 = n28514 & n28515;
  assign n28517 = n6854 & n28516;
  assign n28518 = n26945 & n28517;
  assign n28519 = ~n28503 & n28518;
  assign n28520 = n28503 & ~n28518;
  assign n28521 = ~n28519 & ~n28520;
  assign n28522 = n3896 & n20361;
  assign n28523 = n3683 & n20365;
  assign n28524 = n564 & n20368;
  assign n28525 = n566 & n22848;
  assign n28526 = ~n28523 & ~n28524;
  assign n28527 = ~n28522 & n28526;
  assign n28528 = ~n28525 & n28527;
  assign n28529 = ~n28521 & ~n28528;
  assign n28530 = n28521 & n28528;
  assign n28531 = ~n28529 & ~n28530;
  assign n28532 = ~n28437 & ~n28440;
  assign n28533 = n28531 & n28532;
  assign n28534 = ~n28531 & ~n28532;
  assign n28535 = ~n28533 & ~n28534;
  assign n28536 = n4472 & n23394;
  assign n28537 = n4070 & n20355;
  assign n28538 = n3943 & n20358;
  assign n28539 = n3944 & n23404;
  assign n28540 = ~n28537 & ~n28538;
  assign n28541 = ~n28536 & n28540;
  assign n28542 = ~n28539 & n28541;
  assign n28543 = pi29  & n28542;
  assign n28544 = ~pi29  & ~n28542;
  assign n28545 = ~n28543 & ~n28544;
  assign n28546 = n28535 & ~n28545;
  assign n28547 = ~n28535 & n28545;
  assign n28548 = ~n28546 & ~n28547;
  assign n28549 = ~n28502 & n28548;
  assign n28550 = n28502 & ~n28548;
  assign n28551 = ~n28549 & ~n28550;
  assign n28552 = n4721 & n23765;
  assign n28553 = n4691 & n23768;
  assign n28554 = n4515 & n23771;
  assign n28555 = n4516 & n23789;
  assign n28556 = ~n28553 & ~n28554;
  assign n28557 = ~n28552 & n28556;
  assign n28558 = ~n28555 & n28557;
  assign n28559 = pi26  & n28558;
  assign n28560 = ~pi26  & ~n28558;
  assign n28561 = ~n28559 & ~n28560;
  assign n28562 = n28551 & ~n28561;
  assign n28563 = ~n28551 & n28561;
  assign n28564 = ~n28562 & ~n28563;
  assign n28565 = ~n28501 & n28564;
  assign n28566 = n28501 & ~n28564;
  assign n28567 = ~n28565 & ~n28566;
  assign n28568 = n5267 & n25022;
  assign n28569 = n5185 & n24779;
  assign n28570 = n5121 & n24529;
  assign n28571 = n78 & n25032;
  assign n28572 = ~n28569 & ~n28570;
  assign n28573 = ~n28568 & n28572;
  assign n28574 = ~n28571 & n28573;
  assign n28575 = pi23  & n28574;
  assign n28576 = ~pi23  & ~n28574;
  assign n28577 = ~n28575 & ~n28576;
  assign n28578 = n28567 & ~n28577;
  assign n28579 = ~n28567 & n28577;
  assign n28580 = ~n28578 & ~n28579;
  assign n28581 = n28500 & ~n28580;
  assign n28582 = ~n28500 & n28580;
  assign n28583 = ~n28581 & ~n28582;
  assign n28584 = n5982 & n25709;
  assign n28585 = n5901 & n25490;
  assign n28586 = n5312 & n25253;
  assign n28587 = n5306 & n25719;
  assign n28588 = ~n28585 & ~n28586;
  assign n28589 = ~n28584 & n28588;
  assign n28590 = ~n28587 & n28589;
  assign n28591 = pi20  & n28590;
  assign n28592 = ~pi20  & ~n28590;
  assign n28593 = ~n28591 & ~n28592;
  assign n28594 = n28583 & ~n28593;
  assign n28595 = ~n28583 & n28593;
  assign n28596 = ~n28594 & ~n28595;
  assign n28597 = ~n28499 & n28596;
  assign n28598 = n28499 & ~n28596;
  assign n28599 = ~n28597 & ~n28598;
  assign n28600 = n28498 & ~n28599;
  assign n28601 = ~n28498 & n28599;
  assign n28602 = ~n28600 & ~n28601;
  assign n28603 = n28496 & n28602;
  assign n28604 = ~n28496 & ~n28602;
  assign po23  = ~n28603 & ~n28604;
  assign n28606 = ~n28582 & ~n28594;
  assign n28607 = ~n28565 & ~n28578;
  assign n28608 = ~n12513 & n25709;
  assign n28609 = n5312 & n25490;
  assign n28610 = n5306 & ~n25925;
  assign n28611 = ~n28608 & ~n28609;
  assign n28612 = ~n28610 & n28611;
  assign n28613 = pi20  & n28612;
  assign n28614 = ~pi20  & ~n28612;
  assign n28615 = ~n28613 & ~n28614;
  assign n28616 = ~n28607 & ~n28615;
  assign n28617 = n28607 & n28615;
  assign n28618 = ~n28616 & ~n28617;
  assign n28619 = ~n28549 & ~n28562;
  assign n28620 = n4721 & n24529;
  assign n28621 = n4691 & n23765;
  assign n28622 = n4515 & n23768;
  assign n28623 = n4516 & n24539;
  assign n28624 = ~n28621 & ~n28622;
  assign n28625 = ~n28620 & n28624;
  assign n28626 = ~n28623 & n28625;
  assign n28627 = pi26  & n28626;
  assign n28628 = ~pi26  & ~n28626;
  assign n28629 = ~n28627 & ~n28628;
  assign n28630 = ~n296 & ~n546;
  assign n28631 = n1203 & n28630;
  assign n28632 = n1398 & n3323;
  assign n28633 = n12753 & n28632;
  assign n28634 = n12467 & n28631;
  assign n28635 = n28633 & n28634;
  assign n28636 = n28286 & n28635;
  assign n28637 = n4591 & n26163;
  assign n28638 = n28636 & n28637;
  assign n28639 = n5030 & n6894;
  assign n28640 = n28638 & n28639;
  assign n28641 = n1500 & n28640;
  assign n28642 = ~n28518 & n28641;
  assign n28643 = n28518 & ~n28641;
  assign n28644 = ~n28642 & ~n28643;
  assign n28645 = n3896 & n20358;
  assign n28646 = n3683 & n20361;
  assign n28647 = n564 & n20365;
  assign n28648 = n566 & n22833;
  assign n28649 = ~n28646 & ~n28647;
  assign n28650 = ~n28645 & n28649;
  assign n28651 = ~n28648 & n28650;
  assign n28652 = n28644 & ~n28651;
  assign n28653 = ~n28644 & n28651;
  assign n28654 = ~n28652 & ~n28653;
  assign n28655 = ~n28520 & ~n28530;
  assign n28656 = ~n28654 & ~n28655;
  assign n28657 = n28654 & n28655;
  assign n28658 = ~n28656 & ~n28657;
  assign n28659 = ~n28534 & ~n28546;
  assign n28660 = ~n28658 & n28659;
  assign n28661 = n28658 & ~n28659;
  assign n28662 = ~n28660 & ~n28661;
  assign n28663 = n4472 & n23771;
  assign n28664 = n4070 & n23394;
  assign n28665 = n3943 & n20355;
  assign n28666 = n3944 & n23816;
  assign n28667 = ~n28664 & ~n28665;
  assign n28668 = ~n28663 & n28667;
  assign n28669 = ~n28666 & n28668;
  assign n28670 = pi29  & n28669;
  assign n28671 = ~pi29  & ~n28669;
  assign n28672 = ~n28670 & ~n28671;
  assign n28673 = n28662 & ~n28672;
  assign n28674 = ~n28662 & n28672;
  assign n28675 = ~n28673 & ~n28674;
  assign n28676 = ~n28629 & n28675;
  assign n28677 = n28629 & ~n28675;
  assign n28678 = ~n28676 & ~n28677;
  assign n28679 = n28619 & ~n28678;
  assign n28680 = ~n28619 & n28678;
  assign n28681 = ~n28679 & ~n28680;
  assign n28682 = n5267 & n25253;
  assign n28683 = n5185 & n25022;
  assign n28684 = n5121 & n24779;
  assign n28685 = n78 & n25263;
  assign n28686 = ~n28683 & ~n28684;
  assign n28687 = ~n28682 & n28686;
  assign n28688 = ~n28685 & n28687;
  assign n28689 = pi23  & n28688;
  assign n28690 = ~pi23  & ~n28688;
  assign n28691 = ~n28689 & ~n28690;
  assign n28692 = n28681 & ~n28691;
  assign n28693 = ~n28681 & n28691;
  assign n28694 = ~n28692 & ~n28693;
  assign n28695 = n28618 & n28694;
  assign n28696 = ~n28618 & ~n28694;
  assign n28697 = ~n28695 & ~n28696;
  assign n28698 = n28606 & ~n28697;
  assign n28699 = ~n28606 & n28697;
  assign n28700 = ~n28698 & ~n28699;
  assign n28701 = ~n28597 & ~n28601;
  assign n28702 = ~n28700 & n28701;
  assign n28703 = n28700 & ~n28701;
  assign n28704 = ~n28702 & ~n28703;
  assign n28705 = n28603 & n28704;
  assign n28706 = ~n28603 & ~n28704;
  assign po24  = ~n28705 & ~n28706;
  assign n28708 = ~n28699 & ~n28703;
  assign n28709 = ~n28616 & ~n28695;
  assign n28710 = ~n28673 & ~n28676;
  assign n28711 = ~n28643 & ~n28652;
  assign n28712 = ~n12514 & n25709;
  assign n28713 = pi20  & ~n28712;
  assign n28714 = ~pi20  & n28712;
  assign n28715 = ~n28713 & ~n28714;
  assign n28716 = ~n360 & ~n536;
  assign n28717 = ~n545 & ~n687;
  assign n28718 = n28716 & n28717;
  assign n28719 = n1015 & n1115;
  assign n28720 = n1201 & n1630;
  assign n28721 = n12626 & n28720;
  assign n28722 = n28718 & n28719;
  assign n28723 = n437 & n901;
  assign n28724 = n3400 & n28723;
  assign n28725 = n28721 & n28722;
  assign n28726 = n3176 & n13918;
  assign n28727 = n28725 & n28726;
  assign n28728 = n14737 & n28724;
  assign n28729 = n28727 & n28728;
  assign n28730 = n1861 & n28729;
  assign n28731 = n4928 & n28730;
  assign n28732 = n28518 & n28731;
  assign n28733 = ~n28518 & ~n28731;
  assign n28734 = ~n28732 & ~n28733;
  assign n28735 = n28715 & n28734;
  assign n28736 = ~n28715 & ~n28734;
  assign n28737 = ~n28735 & ~n28736;
  assign n28738 = ~n28711 & n28737;
  assign n28739 = n28711 & ~n28737;
  assign n28740 = ~n28738 & ~n28739;
  assign n28741 = n3896 & n20355;
  assign n28742 = n3683 & n20358;
  assign n28743 = n564 & n20361;
  assign n28744 = n566 & n20562;
  assign n28745 = ~n28742 & ~n28743;
  assign n28746 = ~n28741 & n28745;
  assign n28747 = ~n28744 & n28746;
  assign n28748 = n28740 & n28747;
  assign n28749 = ~n28740 & ~n28747;
  assign n28750 = ~n28748 & ~n28749;
  assign n28751 = ~n28657 & ~n28661;
  assign n28752 = n28750 & n28751;
  assign n28753 = ~n28750 & ~n28751;
  assign n28754 = ~n28752 & ~n28753;
  assign n28755 = n4472 & n23768;
  assign n28756 = n4070 & n23771;
  assign n28757 = n3943 & n23394;
  assign n28758 = n3944 & n23804;
  assign n28759 = ~n28756 & ~n28757;
  assign n28760 = ~n28755 & n28759;
  assign n28761 = ~n28758 & n28760;
  assign n28762 = pi29  & n28761;
  assign n28763 = ~pi29  & ~n28761;
  assign n28764 = ~n28762 & ~n28763;
  assign n28765 = n28754 & ~n28764;
  assign n28766 = ~n28754 & n28764;
  assign n28767 = ~n28765 & ~n28766;
  assign n28768 = n4721 & n24779;
  assign n28769 = n4691 & n24529;
  assign n28770 = n4515 & n23765;
  assign n28771 = n4516 & n24789;
  assign n28772 = ~n28769 & ~n28770;
  assign n28773 = ~n28768 & n28772;
  assign n28774 = ~n28771 & n28773;
  assign n28775 = pi26  & n28774;
  assign n28776 = ~pi26  & ~n28774;
  assign n28777 = ~n28775 & ~n28776;
  assign n28778 = n28767 & ~n28777;
  assign n28779 = ~n28767 & n28777;
  assign n28780 = ~n28778 & ~n28779;
  assign n28781 = n28710 & ~n28780;
  assign n28782 = ~n28710 & n28780;
  assign n28783 = ~n28781 & ~n28782;
  assign n28784 = ~n28680 & ~n28692;
  assign n28785 = n5267 & n25490;
  assign n28786 = n5185 & n25253;
  assign n28787 = n5121 & n25022;
  assign n28788 = n78 & n25500;
  assign n28789 = ~n28786 & ~n28787;
  assign n28790 = ~n28785 & n28789;
  assign n28791 = ~n28788 & n28790;
  assign n28792 = pi23  & n28791;
  assign n28793 = ~pi23  & ~n28791;
  assign n28794 = ~n28792 & ~n28793;
  assign n28795 = ~n28784 & ~n28794;
  assign n28796 = n28784 & n28794;
  assign n28797 = ~n28795 & ~n28796;
  assign n28798 = ~n28783 & ~n28797;
  assign n28799 = n28783 & n28797;
  assign n28800 = ~n28798 & ~n28799;
  assign n28801 = ~n28709 & n28800;
  assign n28802 = n28709 & ~n28800;
  assign n28803 = ~n28801 & ~n28802;
  assign n28804 = ~n28708 & n28803;
  assign n28805 = n28708 & ~n28803;
  assign n28806 = ~n28804 & ~n28805;
  assign n28807 = ~n28705 & ~n28806;
  assign n28808 = n28705 & n28806;
  assign po25  = ~n28807 & ~n28808;
  assign n28810 = ~n28801 & ~n28804;
  assign n28811 = ~n28795 & ~n28799;
  assign n28812 = ~n28753 & ~n28765;
  assign n28813 = ~n28733 & ~n28735;
  assign n28814 = ~n375 & ~n420;
  assign n28815 = ~n572 & n28814;
  assign n28816 = n2097 & n2365;
  assign n28817 = n2452 & n5368;
  assign n28818 = n14711 & n28817;
  assign n28819 = n28815 & n28816;
  assign n28820 = n1207 & n28819;
  assign n28821 = n2423 & n28818;
  assign n28822 = n28820 & n28821;
  assign n28823 = n4271 & n14806;
  assign n28824 = n28822 & n28823;
  assign n28825 = n2490 & n13450;
  assign n28826 = n28824 & n28825;
  assign n28827 = n4604 & n28826;
  assign n28828 = ~n28813 & n28827;
  assign n28829 = n28813 & ~n28827;
  assign n28830 = ~n28828 & ~n28829;
  assign n28831 = n3896 & n23394;
  assign n28832 = n3683 & n20355;
  assign n28833 = n564 & n20358;
  assign n28834 = n566 & n23404;
  assign n28835 = ~n28832 & ~n28833;
  assign n28836 = ~n28831 & n28835;
  assign n28837 = ~n28834 & n28836;
  assign n28838 = ~n28830 & ~n28837;
  assign n28839 = n28830 & n28837;
  assign n28840 = ~n28838 & ~n28839;
  assign n28841 = ~n28739 & ~n28748;
  assign n28842 = n28840 & ~n28841;
  assign n28843 = ~n28840 & n28841;
  assign n28844 = ~n28842 & ~n28843;
  assign n28845 = n4472 & n23765;
  assign n28846 = n4070 & n23768;
  assign n28847 = n3943 & n23771;
  assign n28848 = n3944 & n23789;
  assign n28849 = ~n28846 & ~n28847;
  assign n28850 = ~n28845 & n28849;
  assign n28851 = ~n28848 & n28850;
  assign n28852 = pi29  & n28851;
  assign n28853 = ~pi29  & ~n28851;
  assign n28854 = ~n28852 & ~n28853;
  assign n28855 = n28844 & ~n28854;
  assign n28856 = ~n28844 & n28854;
  assign n28857 = ~n28855 & ~n28856;
  assign n28858 = ~n28812 & n28857;
  assign n28859 = n28812 & ~n28857;
  assign n28860 = ~n28858 & ~n28859;
  assign n28861 = n4721 & n25022;
  assign n28862 = n4691 & n24779;
  assign n28863 = n4515 & n24529;
  assign n28864 = n4516 & n25032;
  assign n28865 = ~n28862 & ~n28863;
  assign n28866 = ~n28861 & n28865;
  assign n28867 = ~n28864 & n28866;
  assign n28868 = pi26  & n28867;
  assign n28869 = ~pi26  & ~n28867;
  assign n28870 = ~n28868 & ~n28869;
  assign n28871 = n28860 & n28870;
  assign n28872 = ~n28860 & ~n28870;
  assign n28873 = ~n28871 & ~n28872;
  assign n28874 = ~n28778 & ~n28782;
  assign n28875 = n28873 & n28874;
  assign n28876 = ~n28873 & ~n28874;
  assign n28877 = ~n28875 & ~n28876;
  assign n28878 = n5267 & n25709;
  assign n28879 = n5185 & n25490;
  assign n28880 = n5121 & n25253;
  assign n28881 = n78 & n25719;
  assign n28882 = ~n28879 & ~n28880;
  assign n28883 = ~n28878 & n28882;
  assign n28884 = ~n28881 & n28883;
  assign n28885 = pi23  & n28884;
  assign n28886 = ~pi23  & ~n28884;
  assign n28887 = ~n28885 & ~n28886;
  assign n28888 = n28877 & ~n28887;
  assign n28889 = ~n28877 & n28887;
  assign n28890 = ~n28888 & ~n28889;
  assign n28891 = ~n28811 & n28890;
  assign n28892 = n28811 & ~n28890;
  assign n28893 = ~n28891 & ~n28892;
  assign n28894 = n28810 & ~n28893;
  assign n28895 = ~n28810 & n28893;
  assign n28896 = ~n28894 & ~n28895;
  assign n28897 = n28808 & n28896;
  assign n28898 = ~n28808 & ~n28896;
  assign po26  = ~n28897 & ~n28898;
  assign n28900 = ~n28876 & ~n28888;
  assign n28901 = ~n12426 & n25709;
  assign n28902 = n5121 & n25490;
  assign n28903 = n78 & ~n25925;
  assign n28904 = ~n28901 & ~n28902;
  assign n28905 = ~n28903 & n28904;
  assign n28906 = pi23  & n28905;
  assign n28907 = ~pi23  & ~n28905;
  assign n28908 = ~n28906 & ~n28907;
  assign n28909 = ~n28859 & ~n28871;
  assign n28910 = ~n28908 & n28909;
  assign n28911 = n28908 & ~n28909;
  assign n28912 = ~n28910 & ~n28911;
  assign n28913 = n4721 & n25253;
  assign n28914 = n4691 & n25022;
  assign n28915 = n4515 & n24779;
  assign n28916 = n4516 & n25263;
  assign n28917 = ~n28914 & ~n28915;
  assign n28918 = ~n28913 & n28917;
  assign n28919 = ~n28916 & n28918;
  assign n28920 = pi26  & n28919;
  assign n28921 = ~pi26  & ~n28919;
  assign n28922 = ~n28920 & ~n28921;
  assign n28923 = ~n28843 & ~n28855;
  assign n28924 = ~n202 & ~n280;
  assign n28925 = ~n290 & ~n424;
  assign n28926 = n28924 & n28925;
  assign n28927 = n471 & n1203;
  assign n28928 = n1208 & n1354;
  assign n28929 = n1909 & n2097;
  assign n28930 = n28928 & n28929;
  assign n28931 = n28926 & n28927;
  assign n28932 = n12128 & n14644;
  assign n28933 = n28931 & n28932;
  assign n28934 = n28930 & n28933;
  assign n28935 = n23590 & n26951;
  assign n28936 = n28934 & n28935;
  assign n28937 = n21648 & n28936;
  assign n28938 = n3728 & n28937;
  assign n28939 = n28827 & ~n28938;
  assign n28940 = ~n28827 & n28938;
  assign n28941 = ~n28939 & ~n28940;
  assign n28942 = ~n28829 & ~n28839;
  assign n28943 = n28941 & n28942;
  assign n28944 = ~n28941 & ~n28942;
  assign n28945 = ~n28943 & ~n28944;
  assign n28946 = n3896 & n23771;
  assign n28947 = n3683 & n23394;
  assign n28948 = n564 & n20355;
  assign n28949 = n566 & n23816;
  assign n28950 = ~n28947 & ~n28948;
  assign n28951 = ~n28946 & n28950;
  assign n28952 = ~n28949 & n28951;
  assign n28953 = n28945 & ~n28952;
  assign n28954 = ~n28945 & n28952;
  assign n28955 = ~n28953 & ~n28954;
  assign n28956 = n28923 & ~n28955;
  assign n28957 = ~n28923 & n28955;
  assign n28958 = ~n28956 & ~n28957;
  assign n28959 = n4472 & n24529;
  assign n28960 = n4070 & n23765;
  assign n28961 = n3943 & n23768;
  assign n28962 = n3944 & n24539;
  assign n28963 = ~n28960 & ~n28961;
  assign n28964 = ~n28959 & n28963;
  assign n28965 = ~n28962 & n28964;
  assign n28966 = pi29  & n28965;
  assign n28967 = ~pi29  & ~n28965;
  assign n28968 = ~n28966 & ~n28967;
  assign n28969 = n28958 & ~n28968;
  assign n28970 = ~n28958 & n28968;
  assign n28971 = ~n28969 & ~n28970;
  assign n28972 = ~n28922 & n28971;
  assign n28973 = n28922 & ~n28971;
  assign n28974 = ~n28972 & ~n28973;
  assign n28975 = n28912 & n28974;
  assign n28976 = ~n28912 & ~n28974;
  assign n28977 = ~n28975 & ~n28976;
  assign n28978 = n28900 & ~n28977;
  assign n28979 = ~n28900 & n28977;
  assign n28980 = ~n28978 & ~n28979;
  assign n28981 = ~n28891 & ~n28895;
  assign n28982 = ~n28980 & n28981;
  assign n28983 = n28980 & ~n28981;
  assign n28984 = ~n28982 & ~n28983;
  assign n28985 = n28897 & n28984;
  assign n28986 = ~n28897 & ~n28984;
  assign po27  = ~n28985 & ~n28986;
  assign n28988 = ~n28979 & ~n28983;
  assign n28989 = ~n28910 & ~n28975;
  assign n28990 = ~n28953 & ~n28957;
  assign n28991 = ~n28940 & ~n28943;
  assign n28992 = ~n23317 & n25709;
  assign n28993 = pi23  & ~n28992;
  assign n28994 = ~pi23  & n28992;
  assign n28995 = ~n28993 & ~n28994;
  assign n28996 = ~n250 & ~n544;
  assign n28997 = n392 & n28996;
  assign n28998 = n664 & n1246;
  assign n28999 = n5527 & n28998;
  assign n29000 = n14662 & n28997;
  assign n29001 = n249 & n29000;
  assign n29002 = n5371 & n28999;
  assign n29003 = n29001 & n29002;
  assign n29004 = n353 & n29003;
  assign n29005 = n611 & n29004;
  assign n29006 = n3660 & n29005;
  assign n29007 = n28938 & n29006;
  assign n29008 = ~n28938 & ~n29006;
  assign n29009 = ~n29007 & ~n29008;
  assign n29010 = n28995 & n29009;
  assign n29011 = ~n28995 & ~n29009;
  assign n29012 = ~n29010 & ~n29011;
  assign n29013 = ~n28991 & n29012;
  assign n29014 = n28991 & ~n29012;
  assign n29015 = ~n29013 & ~n29014;
  assign n29016 = n3896 & n23768;
  assign n29017 = n3683 & n23771;
  assign n29018 = n564 & n23394;
  assign n29019 = n566 & n23804;
  assign n29020 = ~n29017 & ~n29018;
  assign n29021 = ~n29016 & n29020;
  assign n29022 = ~n29019 & n29021;
  assign n29023 = n29015 & ~n29022;
  assign n29024 = ~n29015 & n29022;
  assign n29025 = ~n29023 & ~n29024;
  assign n29026 = n28990 & ~n29025;
  assign n29027 = ~n28990 & n29025;
  assign n29028 = ~n29026 & ~n29027;
  assign n29029 = n4472 & n24779;
  assign n29030 = n4070 & n24529;
  assign n29031 = n3943 & n23765;
  assign n29032 = n3944 & n24789;
  assign n29033 = ~n29030 & ~n29031;
  assign n29034 = ~n29029 & n29033;
  assign n29035 = ~n29032 & n29034;
  assign n29036 = pi29  & n29035;
  assign n29037 = ~pi29  & ~n29035;
  assign n29038 = ~n29036 & ~n29037;
  assign n29039 = n29028 & ~n29038;
  assign n29040 = ~n29028 & n29038;
  assign n29041 = ~n29039 & ~n29040;
  assign n29042 = ~n28969 & ~n28972;
  assign n29043 = n4721 & n25490;
  assign n29044 = n4691 & n25253;
  assign n29045 = n4515 & n25022;
  assign n29046 = n4516 & n25500;
  assign n29047 = ~n29044 & ~n29045;
  assign n29048 = ~n29043 & n29047;
  assign n29049 = ~n29046 & n29048;
  assign n29050 = pi26  & n29049;
  assign n29051 = ~pi26  & ~n29049;
  assign n29052 = ~n29050 & ~n29051;
  assign n29053 = ~n29042 & ~n29052;
  assign n29054 = n29042 & n29052;
  assign n29055 = ~n29053 & ~n29054;
  assign n29056 = n29041 & n29055;
  assign n29057 = ~n29041 & ~n29055;
  assign n29058 = ~n29056 & ~n29057;
  assign n29059 = ~n28989 & n29058;
  assign n29060 = n28989 & ~n29058;
  assign n29061 = ~n29059 & ~n29060;
  assign n29062 = ~n28988 & n29061;
  assign n29063 = n28988 & ~n29061;
  assign n29064 = ~n29062 & ~n29063;
  assign n29065 = ~n28985 & ~n29064;
  assign n29066 = n28985 & n29064;
  assign po28  = ~n29065 & ~n29066;
  assign n29068 = ~n29059 & ~n29062;
  assign n29069 = ~n29053 & ~n29056;
  assign n29070 = ~n29027 & ~n29039;
  assign n29071 = ~n29008 & ~n29010;
  assign n29072 = ~n360 & ~n375;
  assign n29073 = n357 & n29072;
  assign n29074 = n464 & n921;
  assign n29075 = n1342 & n2008;
  assign n29076 = n2220 & n2450;
  assign n29077 = n4418 & n29076;
  assign n29078 = n29074 & n29075;
  assign n29079 = n29073 & n29078;
  assign n29080 = n6938 & n29077;
  assign n29081 = n13882 & n29080;
  assign n29082 = n333 & n29079;
  assign n29083 = n29081 & n29082;
  assign n29084 = n788 & n29083;
  assign n29085 = n14671 & n29084;
  assign n29086 = n23718 & n29085;
  assign n29087 = ~n29071 & n29086;
  assign n29088 = n29071 & ~n29086;
  assign n29089 = ~n29087 & ~n29088;
  assign n29090 = n3896 & n23765;
  assign n29091 = n3683 & n23768;
  assign n29092 = n564 & n23771;
  assign n29093 = n566 & n23789;
  assign n29094 = ~n29091 & ~n29092;
  assign n29095 = ~n29090 & n29094;
  assign n29096 = ~n29093 & n29095;
  assign n29097 = ~n29089 & ~n29096;
  assign n29098 = n29089 & n29096;
  assign n29099 = ~n29097 & ~n29098;
  assign n29100 = ~n29013 & ~n29023;
  assign n29101 = n29099 & n29100;
  assign n29102 = ~n29099 & ~n29100;
  assign n29103 = ~n29101 & ~n29102;
  assign n29104 = n4472 & n25022;
  assign n29105 = n4070 & n24779;
  assign n29106 = n3943 & n24529;
  assign n29107 = n3944 & n25032;
  assign n29108 = ~n29105 & ~n29106;
  assign n29109 = ~n29104 & n29108;
  assign n29110 = ~n29107 & n29109;
  assign n29111 = pi29  & n29110;
  assign n29112 = ~pi29  & ~n29110;
  assign n29113 = ~n29111 & ~n29112;
  assign n29114 = n29103 & ~n29113;
  assign n29115 = ~n29103 & n29113;
  assign n29116 = ~n29114 & ~n29115;
  assign n29117 = ~n29070 & n29116;
  assign n29118 = n29070 & ~n29116;
  assign n29119 = ~n29117 & ~n29118;
  assign n29120 = n4721 & n25709;
  assign n29121 = n4691 & n25490;
  assign n29122 = n4515 & n25253;
  assign n29123 = n4516 & n25719;
  assign n29124 = ~n29121 & ~n29122;
  assign n29125 = ~n29120 & n29124;
  assign n29126 = ~n29123 & n29125;
  assign n29127 = pi26  & n29126;
  assign n29128 = ~pi26  & ~n29126;
  assign n29129 = ~n29127 & ~n29128;
  assign n29130 = n29119 & ~n29129;
  assign n29131 = ~n29119 & n29129;
  assign n29132 = ~n29130 & ~n29131;
  assign n29133 = ~n29069 & n29132;
  assign n29134 = n29069 & ~n29132;
  assign n29135 = ~n29133 & ~n29134;
  assign n29136 = n29068 & ~n29135;
  assign n29137 = ~n29068 & n29135;
  assign n29138 = ~n29136 & ~n29137;
  assign n29139 = n29066 & n29138;
  assign n29140 = ~n29066 & ~n29138;
  assign po29  = ~n29139 & ~n29140;
  assign n29142 = ~n29133 & ~n29137;
  assign n29143 = ~n29117 & ~n29130;
  assign n29144 = ~n29102 & ~n29114;
  assign n29145 = n191 & n3599;
  assign n29146 = n306 & n29145;
  assign n29147 = n456 & n562;
  assign n29148 = n713 & n29147;
  assign n29149 = n29146 & n29148;
  assign n29150 = n23718 & n29149;
  assign n29151 = ~n29086 & n29150;
  assign n29152 = n29086 & ~n29150;
  assign n29153 = ~n29151 & ~n29152;
  assign n29154 = ~n29088 & ~n29098;
  assign n29155 = n29153 & n29154;
  assign n29156 = ~n29153 & ~n29154;
  assign n29157 = ~n29155 & ~n29156;
  assign n29158 = n3896 & n24529;
  assign n29159 = n3683 & n23765;
  assign n29160 = n564 & n23768;
  assign n29161 = n566 & n24539;
  assign n29162 = ~n29159 & ~n29160;
  assign n29163 = ~n29158 & n29162;
  assign n29164 = ~n29161 & n29163;
  assign n29165 = n29157 & ~n29164;
  assign n29166 = ~n29157 & n29164;
  assign n29167 = ~n29165 & ~n29166;
  assign n29168 = n29144 & ~n29167;
  assign n29169 = ~n29144 & n29167;
  assign n29170 = ~n29168 & ~n29169;
  assign n29171 = n4515 & n25490;
  assign n29172 = n4516 & ~n25925;
  assign n29173 = ~n4514 & ~n4516;
  assign n29174 = n25709 & n29173;
  assign n29175 = ~n29171 & ~n29174;
  assign n29176 = ~n29172 & n29175;
  assign n29177 = ~pi26  & ~n29176;
  assign n29178 = pi26  & n29176;
  assign n29179 = ~n29177 & ~n29178;
  assign n29180 = n4472 & n25253;
  assign n29181 = n4070 & n25022;
  assign n29182 = n3943 & n24779;
  assign n29183 = n3944 & n25263;
  assign n29184 = ~n29181 & ~n29182;
  assign n29185 = ~n29180 & n29184;
  assign n29186 = ~n29183 & n29185;
  assign n29187 = pi29  & n29186;
  assign n29188 = ~pi29  & ~n29186;
  assign n29189 = ~n29187 & ~n29188;
  assign n29190 = ~n29179 & ~n29189;
  assign n29191 = n29179 & n29189;
  assign n29192 = ~n29190 & ~n29191;
  assign n29193 = ~n29170 & ~n29192;
  assign n29194 = n29170 & n29192;
  assign n29195 = ~n29193 & ~n29194;
  assign n29196 = ~n29143 & n29195;
  assign n29197 = n29143 & ~n29195;
  assign n29198 = ~n29196 & ~n29197;
  assign n29199 = ~n29142 & n29198;
  assign n29200 = n29142 & ~n29198;
  assign n29201 = ~n29199 & ~n29200;
  assign n29202 = ~n29139 & ~n29201;
  assign n29203 = n29139 & n29201;
  assign po30  = ~n29202 & ~n29203;
  assign n29205 = ~n23688 & n25709;
  assign n29206 = n29203 & ~n29205;
  assign n29207 = ~n29203 & n29205;
  assign n29208 = ~n29206 & ~n29207;
  assign n29209 = ~n29196 & ~n29199;
  assign n29210 = ~n29190 & ~n29194;
  assign n29211 = n29209 & ~n29210;
  assign n29212 = ~n29209 & n29210;
  assign n29213 = ~n29211 & ~n29212;
  assign n29214 = n29086 & n29213;
  assign n29215 = ~n29086 & ~n29213;
  assign n29216 = ~n29214 & ~n29215;
  assign n29217 = n534 & n618;
  assign n29218 = pi26  & ~n29217;
  assign n29219 = ~pi26  & n29217;
  assign n29220 = ~n29218 & ~n29219;
  assign n29221 = ~n29165 & ~n29169;
  assign n29222 = ~n29152 & ~n29155;
  assign n29223 = n29221 & ~n29222;
  assign n29224 = ~n29221 & n29222;
  assign n29225 = ~n29223 & ~n29224;
  assign n29226 = n4472 & n25490;
  assign n29227 = n4070 & n25253;
  assign n29228 = n3943 & n25022;
  assign n29229 = n3944 & n25500;
  assign n29230 = ~n29227 & ~n29228;
  assign n29231 = ~n29226 & n29230;
  assign n29232 = ~n29229 & n29231;
  assign n29233 = pi29  & ~n29232;
  assign n29234 = ~pi29  & n29232;
  assign n29235 = ~n29233 & ~n29234;
  assign n29236 = n3896 & n24779;
  assign n29237 = n3683 & n24529;
  assign n29238 = n564 & n23765;
  assign n29239 = n566 & n24789;
  assign n29240 = ~n29237 & ~n29238;
  assign n29241 = ~n29236 & n29240;
  assign n29242 = ~n29239 & n29241;
  assign n29243 = n29235 & ~n29242;
  assign n29244 = ~n29235 & n29242;
  assign n29245 = ~n29243 & ~n29244;
  assign n29246 = n29225 & n29245;
  assign n29247 = ~n29225 & ~n29245;
  assign n29248 = ~n29246 & ~n29247;
  assign n29249 = n29220 & ~n29248;
  assign n29250 = ~n29220 & n29248;
  assign n29251 = ~n29249 & ~n29250;
  assign n29252 = n29216 & ~n29251;
  assign n29253 = ~n29216 & n29251;
  assign n29254 = ~n29252 & ~n29253;
  assign n29255 = n29208 & n29254;
  assign n29256 = ~n29208 & ~n29254;
  assign po31  = n29255 | n29256;
endmodule
