module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 ,
    pi131 , pi132 , pi133 , pi134 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 ,
    pi130 , pi131 , pi132 , pi133 , pi134 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ;
  wire n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396,
    n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426,
    n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894,
    n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924,
    n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170,
    n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182,
    n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200,
    n3201, n3202, n3203, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212,
    n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242,
    n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272,
    n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302,
    n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332,
    n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362,
    n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3390, n3391, n3392,
    n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416,
    n3417, n3418, n3419, n3420, n3421, n3422,
    n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3439, n3440,
    n3441, n3442, n3443, n3444, n3445, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476,
    n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722,
    n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782,
    n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052,
    n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292,
    n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334,
    n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346,
    n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382,
    n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412,
    n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430,
    n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442,
    n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466,
    n4467, n4468, n4469, n4470, n4471, n4472,
    n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496,
    n4497, n4498, n4499, n4500, n4501, n4502,
    n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526,
    n4527, n4528, n4529, n4530, n4531, n4532,
    n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562,
    n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586,
    n4587, n4588, n4589, n4590, n4591, n4592,
    n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622,
    n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700,
    n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708, n4709, n4710, n4711, n4712,
    n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924;
  assign n264 = ~pi130  & ~pi131 ;
  assign n265 = pi77  & pi128 ;
  assign n266 = pi78  & ~pi128 ;
  assign n267 = ~pi78  & ~pi128 ;
  assign n268 = ~pi77  & pi128 ;
  assign n269 = ~n267 & ~n268;
  assign n270 = ~n265 & ~n266;
  assign n271 = pi129  & n265;
  assign n272 = pi129  & n266;
  assign n273 = ~n271 & ~n272;
  assign n274 = pi129  & n4545;
  assign n275 = pi80  & ~pi128 ;
  assign n276 = pi79  & pi128 ;
  assign n277 = ~pi79  & pi128 ;
  assign n278 = ~pi80  & ~pi128 ;
  assign n279 = ~n277 & ~n278;
  assign n280 = ~n275 & ~n276;
  assign n281 = ~pi129  & n275;
  assign n282 = ~pi129  & n276;
  assign n283 = ~n281 & ~n282;
  assign n284 = ~pi129  & n4547;
  assign n285 = pi129  & ~n4545;
  assign n286 = ~pi129  & ~n4547;
  assign n287 = ~n285 & ~n286;
  assign n288 = n4546 & n4548;
  assign n289 = n264 & n4549;
  assign n290 = pi130  & ~pi131 ;
  assign n291 = pi73  & pi128 ;
  assign n292 = pi74  & ~pi128 ;
  assign n293 = ~pi74  & ~pi128 ;
  assign n294 = ~pi73  & pi128 ;
  assign n295 = ~n293 & ~n294;
  assign n296 = ~n291 & ~n292;
  assign n297 = pi129  & n291;
  assign n298 = pi129  & n292;
  assign n299 = ~n297 & ~n298;
  assign n300 = pi129  & n4550;
  assign n301 = pi76  & ~pi128 ;
  assign n302 = pi75  & pi128 ;
  assign n303 = ~pi75  & pi128 ;
  assign n304 = ~pi76  & ~pi128 ;
  assign n305 = ~n303 & ~n304;
  assign n306 = ~n301 & ~n302;
  assign n307 = ~pi129  & n301;
  assign n308 = ~pi129  & n302;
  assign n309 = ~n307 & ~n308;
  assign n310 = ~pi129  & n4552;
  assign n311 = pi129  & ~n4550;
  assign n312 = ~pi129  & ~n4552;
  assign n313 = ~n311 & ~n312;
  assign n314 = n4551 & n4553;
  assign n315 = n290 & n4554;
  assign n316 = ~n289 & ~n315;
  assign n317 = pi130  & pi131 ;
  assign n318 = pi65  & pi128 ;
  assign n319 = pi66  & ~pi128 ;
  assign n320 = ~pi66  & ~pi128 ;
  assign n321 = ~pi65  & pi128 ;
  assign n322 = ~n320 & ~n321;
  assign n323 = ~n318 & ~n319;
  assign n324 = pi129  & n318;
  assign n325 = pi129  & n319;
  assign n326 = ~n324 & ~n325;
  assign n327 = pi129  & n4555;
  assign n328 = pi68  & ~pi128 ;
  assign n329 = pi67  & pi128 ;
  assign n330 = ~pi67  & pi128 ;
  assign n331 = ~pi68  & ~pi128 ;
  assign n332 = ~n330 & ~n331;
  assign n333 = ~n328 & ~n329;
  assign n334 = ~pi129  & n328;
  assign n335 = ~pi129  & n329;
  assign n336 = ~n334 & ~n335;
  assign n337 = ~pi129  & n4557;
  assign n338 = pi129  & ~n4555;
  assign n339 = ~pi129  & ~n4557;
  assign n340 = ~n338 & ~n339;
  assign n341 = n4556 & n4558;
  assign n342 = n317 & n4559;
  assign n343 = ~pi130  & pi131 ;
  assign n344 = pi69  & pi128 ;
  assign n345 = pi70  & ~pi128 ;
  assign n346 = ~pi70  & ~pi128 ;
  assign n347 = ~pi69  & pi128 ;
  assign n348 = ~n346 & ~n347;
  assign n349 = ~n344 & ~n345;
  assign n350 = pi129  & n344;
  assign n351 = pi129  & n345;
  assign n352 = ~n350 & ~n351;
  assign n353 = pi129  & n4560;
  assign n354 = pi72  & ~pi128 ;
  assign n355 = pi71  & pi128 ;
  assign n356 = ~pi71  & pi128 ;
  assign n357 = ~pi72  & ~pi128 ;
  assign n358 = ~n356 & ~n357;
  assign n359 = ~n354 & ~n355;
  assign n360 = ~pi129  & n354;
  assign n361 = ~pi129  & n355;
  assign n362 = ~n360 & ~n361;
  assign n363 = ~pi129  & n4562;
  assign n364 = pi129  & ~n4560;
  assign n365 = ~pi129  & ~n4562;
  assign n366 = ~n364 & ~n365;
  assign n367 = n4561 & n4563;
  assign n368 = n343 & n4564;
  assign n369 = ~n342 & ~n368;
  assign n370 = n316 & n369;
  assign n371 = pi132  & pi133 ;
  assign n372 = ~n370 & n371;
  assign n373 = pi93  & pi128 ;
  assign n374 = pi94  & ~pi128 ;
  assign n375 = ~pi94  & ~pi128 ;
  assign n376 = ~pi93  & pi128 ;
  assign n377 = ~n375 & ~n376;
  assign n378 = ~n373 & ~n374;
  assign n379 = pi129  & n373;
  assign n380 = pi129  & n374;
  assign n381 = ~n379 & ~n380;
  assign n382 = pi129  & n4565;
  assign n383 = pi96  & ~pi128 ;
  assign n384 = pi95  & pi128 ;
  assign n385 = ~pi95  & pi128 ;
  assign n386 = ~pi96  & ~pi128 ;
  assign n387 = ~n385 & ~n386;
  assign n388 = ~n383 & ~n384;
  assign n389 = ~pi129  & n383;
  assign n390 = ~pi129  & n384;
  assign n391 = ~n389 & ~n390;
  assign n392 = ~pi129  & n4567;
  assign n393 = pi129  & ~n4565;
  assign n394 = ~pi129  & ~n4567;
  assign n395 = ~n393 & ~n394;
  assign n396 = n4566 & n4568;
  assign n397 = n264 & n4569;
  assign n398 = pi89  & pi128 ;
  assign n399 = pi90  & ~pi128 ;
  assign n400 = ~pi90  & ~pi128 ;
  assign n401 = ~pi89  & pi128 ;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~n398 & ~n399;
  assign n404 = pi129  & n398;
  assign n405 = pi129  & n399;
  assign n406 = ~n404 & ~n405;
  assign n407 = pi129  & n4570;
  assign n408 = pi92  & ~pi128 ;
  assign n409 = pi91  & pi128 ;
  assign n410 = ~pi91  & pi128 ;
  assign n411 = ~pi92  & ~pi128 ;
  assign n412 = ~n410 & ~n411;
  assign n413 = ~n408 & ~n409;
  assign n414 = ~pi129  & n408;
  assign n415 = ~pi129  & n409;
  assign n416 = ~n414 & ~n415;
  assign n417 = ~pi129  & n4572;
  assign n418 = pi129  & ~n4570;
  assign n419 = ~pi129  & ~n4572;
  assign n420 = ~n418 & ~n419;
  assign n421 = n4571 & n4573;
  assign n422 = n290 & n4574;
  assign n423 = ~n397 & ~n422;
  assign n424 = pi81  & pi128 ;
  assign n425 = pi82  & ~pi128 ;
  assign n426 = ~pi82  & ~pi128 ;
  assign n427 = ~pi81  & pi128 ;
  assign n428 = ~n426 & ~n427;
  assign n429 = ~n424 & ~n425;
  assign n430 = pi129  & n424;
  assign n431 = pi129  & n425;
  assign n432 = ~n430 & ~n431;
  assign n433 = pi129  & n4575;
  assign n434 = pi84  & ~pi128 ;
  assign n435 = pi83  & pi128 ;
  assign n436 = ~pi83  & pi128 ;
  assign n437 = ~pi84  & ~pi128 ;
  assign n438 = ~n436 & ~n437;
  assign n439 = ~n434 & ~n435;
  assign n440 = ~pi129  & n434;
  assign n441 = ~pi129  & n435;
  assign n442 = ~n440 & ~n441;
  assign n443 = ~pi129  & n4577;
  assign n444 = pi129  & ~n4575;
  assign n445 = ~pi129  & ~n4577;
  assign n446 = ~n444 & ~n445;
  assign n447 = n4576 & n4578;
  assign n448 = n317 & n4579;
  assign n449 = pi85  & pi128 ;
  assign n450 = pi86  & ~pi128 ;
  assign n451 = ~pi86  & ~pi128 ;
  assign n452 = ~pi85  & pi128 ;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~n449 & ~n450;
  assign n455 = pi129  & n449;
  assign n456 = pi129  & n450;
  assign n457 = ~n455 & ~n456;
  assign n458 = pi129  & n4580;
  assign n459 = pi88  & ~pi128 ;
  assign n460 = pi87  & pi128 ;
  assign n461 = ~pi87  & pi128 ;
  assign n462 = ~pi88  & ~pi128 ;
  assign n463 = ~n461 & ~n462;
  assign n464 = ~n459 & ~n460;
  assign n465 = ~pi129  & n459;
  assign n466 = ~pi129  & n460;
  assign n467 = ~n465 & ~n466;
  assign n468 = ~pi129  & n4582;
  assign n469 = pi129  & ~n4580;
  assign n470 = ~pi129  & ~n4582;
  assign n471 = ~n469 & ~n470;
  assign n472 = n4581 & n4583;
  assign n473 = n343 & n4584;
  assign n474 = ~n448 & ~n473;
  assign n475 = n423 & n474;
  assign n476 = ~pi132  & pi133 ;
  assign n477 = ~n475 & n476;
  assign n478 = ~n372 & ~n477;
  assign n479 = pi125  & pi128 ;
  assign n480 = pi126  & ~pi128 ;
  assign n481 = ~pi126  & ~pi128 ;
  assign n482 = ~pi125  & pi128 ;
  assign n483 = ~n481 & ~n482;
  assign n484 = ~n479 & ~n480;
  assign n485 = pi129  & n479;
  assign n486 = pi129  & n480;
  assign n487 = ~n485 & ~n486;
  assign n488 = pi129  & n4585;
  assign n489 = pi0  & ~pi128 ;
  assign n490 = pi127  & pi128 ;
  assign n491 = ~pi127  & pi128 ;
  assign n492 = ~pi0  & ~pi128 ;
  assign n493 = ~n491 & ~n492;
  assign n494 = ~n489 & ~n490;
  assign n495 = ~pi129  & n489;
  assign n496 = ~pi129  & n490;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~pi129  & n4587;
  assign n499 = pi129  & ~n4585;
  assign n500 = ~pi129  & ~n4587;
  assign n501 = ~n499 & ~n500;
  assign n502 = n4586 & n4588;
  assign n503 = n264 & n4589;
  assign n504 = pi121  & pi128 ;
  assign n505 = pi122  & ~pi128 ;
  assign n506 = ~pi122  & ~pi128 ;
  assign n507 = ~pi121  & pi128 ;
  assign n508 = ~n506 & ~n507;
  assign n509 = ~n504 & ~n505;
  assign n510 = pi129  & n504;
  assign n511 = pi129  & n505;
  assign n512 = ~n510 & ~n511;
  assign n513 = pi129  & n4590;
  assign n514 = pi124  & ~pi128 ;
  assign n515 = pi123  & pi128 ;
  assign n516 = ~pi123  & pi128 ;
  assign n517 = ~pi124  & ~pi128 ;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n514 & ~n515;
  assign n520 = ~pi129  & n514;
  assign n521 = ~pi129  & n515;
  assign n522 = ~n520 & ~n521;
  assign n523 = ~pi129  & n4592;
  assign n524 = pi129  & ~n4590;
  assign n525 = ~pi129  & ~n4592;
  assign n526 = ~n524 & ~n525;
  assign n527 = n4591 & n4593;
  assign n528 = n290 & n4594;
  assign n529 = ~n503 & ~n528;
  assign n530 = pi113  & pi128 ;
  assign n531 = pi114  & ~pi128 ;
  assign n532 = ~pi114  & ~pi128 ;
  assign n533 = ~pi113  & pi128 ;
  assign n534 = ~n532 & ~n533;
  assign n535 = ~n530 & ~n531;
  assign n536 = pi129  & n530;
  assign n537 = pi129  & n531;
  assign n538 = ~n536 & ~n537;
  assign n539 = pi129  & n4595;
  assign n540 = pi116  & ~pi128 ;
  assign n541 = pi115  & pi128 ;
  assign n542 = ~pi115  & pi128 ;
  assign n543 = ~pi116  & ~pi128 ;
  assign n544 = ~n542 & ~n543;
  assign n545 = ~n540 & ~n541;
  assign n546 = ~pi129  & n540;
  assign n547 = ~pi129  & n541;
  assign n548 = ~n546 & ~n547;
  assign n549 = ~pi129  & n4597;
  assign n550 = pi129  & ~n4595;
  assign n551 = ~pi129  & ~n4597;
  assign n552 = ~n550 & ~n551;
  assign n553 = n4596 & n4598;
  assign n554 = n317 & n4599;
  assign n555 = pi117  & pi128 ;
  assign n556 = pi118  & ~pi128 ;
  assign n557 = ~pi118  & ~pi128 ;
  assign n558 = ~pi117  & pi128 ;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~n555 & ~n556;
  assign n561 = pi129  & n555;
  assign n562 = pi129  & n556;
  assign n563 = ~n561 & ~n562;
  assign n564 = pi129  & n4600;
  assign n565 = pi120  & ~pi128 ;
  assign n566 = pi119  & pi128 ;
  assign n567 = ~pi119  & pi128 ;
  assign n568 = ~pi120  & ~pi128 ;
  assign n569 = ~n567 & ~n568;
  assign n570 = ~n565 & ~n566;
  assign n571 = ~pi129  & n565;
  assign n572 = ~pi129  & n566;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~pi129  & n4602;
  assign n575 = pi129  & ~n4600;
  assign n576 = ~pi129  & ~n4602;
  assign n577 = ~n575 & ~n576;
  assign n578 = n4601 & n4603;
  assign n579 = n343 & n4604;
  assign n580 = ~n554 & ~n579;
  assign n581 = n529 & n580;
  assign n582 = ~pi132  & ~pi133 ;
  assign n583 = ~n581 & n582;
  assign n584 = pi109  & pi128 ;
  assign n585 = pi110  & ~pi128 ;
  assign n586 = ~pi110  & ~pi128 ;
  assign n587 = ~pi109  & pi128 ;
  assign n588 = ~n586 & ~n587;
  assign n589 = ~n584 & ~n585;
  assign n590 = pi129  & n584;
  assign n591 = pi129  & n585;
  assign n592 = ~n590 & ~n591;
  assign n593 = pi129  & n4605;
  assign n594 = pi112  & ~pi128 ;
  assign n595 = pi111  & pi128 ;
  assign n596 = ~pi111  & pi128 ;
  assign n597 = ~pi112  & ~pi128 ;
  assign n598 = ~n596 & ~n597;
  assign n599 = ~n594 & ~n595;
  assign n600 = ~pi129  & n594;
  assign n601 = ~pi129  & n595;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~pi129  & n4607;
  assign n604 = pi129  & ~n4605;
  assign n605 = ~pi129  & ~n4607;
  assign n606 = ~n604 & ~n605;
  assign n607 = n4606 & n4608;
  assign n608 = n264 & n4609;
  assign n609 = pi105  & pi128 ;
  assign n610 = pi106  & ~pi128 ;
  assign n611 = ~pi106  & ~pi128 ;
  assign n612 = ~pi105  & pi128 ;
  assign n613 = ~n611 & ~n612;
  assign n614 = ~n609 & ~n610;
  assign n615 = pi129  & n609;
  assign n616 = pi129  & n610;
  assign n617 = ~n615 & ~n616;
  assign n618 = pi129  & n4610;
  assign n619 = pi108  & ~pi128 ;
  assign n620 = pi107  & pi128 ;
  assign n621 = ~pi107  & pi128 ;
  assign n622 = ~pi108  & ~pi128 ;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~n619 & ~n620;
  assign n625 = ~pi129  & n619;
  assign n626 = ~pi129  & n620;
  assign n627 = ~n625 & ~n626;
  assign n628 = ~pi129  & n4612;
  assign n629 = pi129  & ~n4610;
  assign n630 = ~pi129  & ~n4612;
  assign n631 = ~n629 & ~n630;
  assign n632 = n4611 & n4613;
  assign n633 = n290 & n4614;
  assign n634 = ~n608 & ~n633;
  assign n635 = pi97  & pi128 ;
  assign n636 = pi98  & ~pi128 ;
  assign n637 = ~pi98  & ~pi128 ;
  assign n638 = ~pi97  & pi128 ;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~n635 & ~n636;
  assign n641 = pi129  & n635;
  assign n642 = pi129  & n636;
  assign n643 = ~n641 & ~n642;
  assign n644 = pi129  & n4615;
  assign n645 = pi100  & ~pi128 ;
  assign n646 = pi99  & pi128 ;
  assign n647 = ~pi99  & pi128 ;
  assign n648 = ~pi100  & ~pi128 ;
  assign n649 = ~n647 & ~n648;
  assign n650 = ~n645 & ~n646;
  assign n651 = ~pi129  & n645;
  assign n652 = ~pi129  & n646;
  assign n653 = ~n651 & ~n652;
  assign n654 = ~pi129  & n4617;
  assign n655 = pi129  & ~n4615;
  assign n656 = ~pi129  & ~n4617;
  assign n657 = ~n655 & ~n656;
  assign n658 = n4616 & n4618;
  assign n659 = n317 & n4619;
  assign n660 = pi101  & pi128 ;
  assign n661 = pi102  & ~pi128 ;
  assign n662 = ~pi102  & ~pi128 ;
  assign n663 = ~pi101  & pi128 ;
  assign n664 = ~n662 & ~n663;
  assign n665 = ~n660 & ~n661;
  assign n666 = pi129  & n660;
  assign n667 = pi129  & n661;
  assign n668 = ~n666 & ~n667;
  assign n669 = pi129  & n4620;
  assign n670 = pi104  & ~pi128 ;
  assign n671 = pi103  & pi128 ;
  assign n672 = ~pi103  & pi128 ;
  assign n673 = ~pi104  & ~pi128 ;
  assign n674 = ~n672 & ~n673;
  assign n675 = ~n670 & ~n671;
  assign n676 = ~pi129  & n670;
  assign n677 = ~pi129  & n671;
  assign n678 = ~n676 & ~n677;
  assign n679 = ~pi129  & n4622;
  assign n680 = pi129  & ~n4620;
  assign n681 = ~pi129  & ~n4622;
  assign n682 = ~n680 & ~n681;
  assign n683 = n4621 & n4623;
  assign n684 = n343 & n4624;
  assign n685 = ~n659 & ~n684;
  assign n686 = n634 & n685;
  assign n687 = pi132  & ~pi133 ;
  assign n688 = ~n686 & n687;
  assign n689 = ~n583 & ~n688;
  assign n690 = n478 & n689;
  assign n691 = ~pi134  & ~n690;
  assign n692 = pi13  & pi128 ;
  assign n693 = pi14  & ~pi128 ;
  assign n694 = ~pi14  & ~pi128 ;
  assign n695 = ~pi13  & pi128 ;
  assign n696 = ~n694 & ~n695;
  assign n697 = ~n692 & ~n693;
  assign n698 = pi129  & n692;
  assign n699 = pi129  & n693;
  assign n700 = ~n698 & ~n699;
  assign n701 = pi129  & n4625;
  assign n702 = pi16  & ~pi128 ;
  assign n703 = pi15  & pi128 ;
  assign n704 = ~pi15  & pi128 ;
  assign n705 = ~pi16  & ~pi128 ;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n702 & ~n703;
  assign n708 = ~pi129  & n702;
  assign n709 = ~pi129  & n703;
  assign n710 = ~n708 & ~n709;
  assign n711 = ~pi129  & n4627;
  assign n712 = pi129  & ~n4625;
  assign n713 = ~pi129  & ~n4627;
  assign n714 = ~n712 & ~n713;
  assign n715 = n4626 & n4628;
  assign n716 = n264 & n4629;
  assign n717 = pi9  & pi128 ;
  assign n718 = pi10  & ~pi128 ;
  assign n719 = ~pi10  & ~pi128 ;
  assign n720 = ~pi9  & pi128 ;
  assign n721 = ~n719 & ~n720;
  assign n722 = ~n717 & ~n718;
  assign n723 = pi129  & n717;
  assign n724 = pi129  & n718;
  assign n725 = ~n723 & ~n724;
  assign n726 = pi129  & n4630;
  assign n727 = pi12  & ~pi128 ;
  assign n728 = pi11  & pi128 ;
  assign n729 = ~pi11  & pi128 ;
  assign n730 = ~pi12  & ~pi128 ;
  assign n731 = ~n729 & ~n730;
  assign n732 = ~n727 & ~n728;
  assign n733 = ~pi129  & n727;
  assign n734 = ~pi129  & n728;
  assign n735 = ~n733 & ~n734;
  assign n736 = ~pi129  & n4632;
  assign n737 = pi129  & ~n4630;
  assign n738 = ~pi129  & ~n4632;
  assign n739 = ~n737 & ~n738;
  assign n740 = n4631 & n4633;
  assign n741 = n290 & n4634;
  assign n742 = ~n716 & ~n741;
  assign n743 = pi1  & pi128 ;
  assign n744 = pi2  & ~pi128 ;
  assign n745 = ~pi2  & ~pi128 ;
  assign n746 = ~pi1  & pi128 ;
  assign n747 = ~n745 & ~n746;
  assign n748 = ~n743 & ~n744;
  assign n749 = pi129  & n743;
  assign n750 = pi129  & n744;
  assign n751 = ~n749 & ~n750;
  assign n752 = pi129  & n4635;
  assign n753 = pi4  & ~pi128 ;
  assign n754 = pi3  & pi128 ;
  assign n755 = ~pi3  & pi128 ;
  assign n756 = ~pi4  & ~pi128 ;
  assign n757 = ~n755 & ~n756;
  assign n758 = ~n753 & ~n754;
  assign n759 = ~pi129  & n753;
  assign n760 = ~pi129  & n754;
  assign n761 = ~n759 & ~n760;
  assign n762 = ~pi129  & n4637;
  assign n763 = pi129  & ~n4635;
  assign n764 = ~pi129  & ~n4637;
  assign n765 = ~n763 & ~n764;
  assign n766 = n4636 & n4638;
  assign n767 = n317 & n4639;
  assign n768 = pi5  & pi128 ;
  assign n769 = pi6  & ~pi128 ;
  assign n770 = ~pi6  & ~pi128 ;
  assign n771 = ~pi5  & pi128 ;
  assign n772 = ~n770 & ~n771;
  assign n773 = ~n768 & ~n769;
  assign n774 = pi129  & n768;
  assign n775 = pi129  & n769;
  assign n776 = ~n774 & ~n775;
  assign n777 = pi129  & n4640;
  assign n778 = pi8  & ~pi128 ;
  assign n779 = pi7  & pi128 ;
  assign n780 = ~pi7  & pi128 ;
  assign n781 = ~pi8  & ~pi128 ;
  assign n782 = ~n780 & ~n781;
  assign n783 = ~n778 & ~n779;
  assign n784 = ~pi129  & n778;
  assign n785 = ~pi129  & n779;
  assign n786 = ~n784 & ~n785;
  assign n787 = ~pi129  & n4642;
  assign n788 = pi129  & ~n4640;
  assign n789 = ~pi129  & ~n4642;
  assign n790 = ~n788 & ~n789;
  assign n791 = n4641 & n4643;
  assign n792 = n343 & n4644;
  assign n793 = ~n767 & ~n792;
  assign n794 = n742 & n793;
  assign n795 = n371 & ~n794;
  assign n796 = pi29  & pi128 ;
  assign n797 = pi30  & ~pi128 ;
  assign n798 = ~pi30  & ~pi128 ;
  assign n799 = ~pi29  & pi128 ;
  assign n800 = ~n798 & ~n799;
  assign n801 = ~n796 & ~n797;
  assign n802 = pi129  & n796;
  assign n803 = pi129  & n797;
  assign n804 = ~n802 & ~n803;
  assign n805 = pi129  & n4645;
  assign n806 = pi32  & ~pi128 ;
  assign n807 = pi31  & pi128 ;
  assign n808 = ~pi31  & pi128 ;
  assign n809 = ~pi32  & ~pi128 ;
  assign n810 = ~n808 & ~n809;
  assign n811 = ~n806 & ~n807;
  assign n812 = ~pi129  & n806;
  assign n813 = ~pi129  & n807;
  assign n814 = ~n812 & ~n813;
  assign n815 = ~pi129  & n4647;
  assign n816 = pi129  & ~n4645;
  assign n817 = ~pi129  & ~n4647;
  assign n818 = ~n816 & ~n817;
  assign n819 = n4646 & n4648;
  assign n820 = n264 & n4649;
  assign n821 = pi25  & pi128 ;
  assign n822 = pi26  & ~pi128 ;
  assign n823 = ~pi26  & ~pi128 ;
  assign n824 = ~pi25  & pi128 ;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~n821 & ~n822;
  assign n827 = pi129  & n821;
  assign n828 = pi129  & n822;
  assign n829 = ~n827 & ~n828;
  assign n830 = pi129  & n4650;
  assign n831 = pi28  & ~pi128 ;
  assign n832 = pi27  & pi128 ;
  assign n833 = ~pi27  & pi128 ;
  assign n834 = ~pi28  & ~pi128 ;
  assign n835 = ~n833 & ~n834;
  assign n836 = ~n831 & ~n832;
  assign n837 = ~pi129  & n831;
  assign n838 = ~pi129  & n832;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~pi129  & n4652;
  assign n841 = pi129  & ~n4650;
  assign n842 = ~pi129  & ~n4652;
  assign n843 = ~n841 & ~n842;
  assign n844 = n4651 & n4653;
  assign n845 = n290 & n4654;
  assign n846 = ~n820 & ~n845;
  assign n847 = pi17  & pi128 ;
  assign n848 = pi18  & ~pi128 ;
  assign n849 = ~pi18  & ~pi128 ;
  assign n850 = ~pi17  & pi128 ;
  assign n851 = ~n849 & ~n850;
  assign n852 = ~n847 & ~n848;
  assign n853 = pi129  & n847;
  assign n854 = pi129  & n848;
  assign n855 = ~n853 & ~n854;
  assign n856 = pi129  & n4655;
  assign n857 = pi20  & ~pi128 ;
  assign n858 = pi19  & pi128 ;
  assign n859 = ~pi19  & pi128 ;
  assign n860 = ~pi20  & ~pi128 ;
  assign n861 = ~n859 & ~n860;
  assign n862 = ~n857 & ~n858;
  assign n863 = ~pi129  & n857;
  assign n864 = ~pi129  & n858;
  assign n865 = ~n863 & ~n864;
  assign n866 = ~pi129  & n4657;
  assign n867 = pi129  & ~n4655;
  assign n868 = ~pi129  & ~n4657;
  assign n869 = ~n867 & ~n868;
  assign n870 = n4656 & n4658;
  assign n871 = n317 & n4659;
  assign n872 = pi21  & pi128 ;
  assign n873 = pi22  & ~pi128 ;
  assign n874 = ~pi22  & ~pi128 ;
  assign n875 = ~pi21  & pi128 ;
  assign n876 = ~n874 & ~n875;
  assign n877 = ~n872 & ~n873;
  assign n878 = pi129  & n872;
  assign n879 = pi129  & n873;
  assign n880 = ~n878 & ~n879;
  assign n881 = pi129  & n4660;
  assign n882 = pi24  & ~pi128 ;
  assign n883 = pi23  & pi128 ;
  assign n884 = ~pi23  & pi128 ;
  assign n885 = ~pi24  & ~pi128 ;
  assign n886 = ~n884 & ~n885;
  assign n887 = ~n882 & ~n883;
  assign n888 = ~pi129  & n882;
  assign n889 = ~pi129  & n883;
  assign n890 = ~n888 & ~n889;
  assign n891 = ~pi129  & n4662;
  assign n892 = pi129  & ~n4660;
  assign n893 = ~pi129  & ~n4662;
  assign n894 = ~n892 & ~n893;
  assign n895 = n4661 & n4663;
  assign n896 = n343 & n4664;
  assign n897 = ~n871 & ~n896;
  assign n898 = n846 & n897;
  assign n899 = n476 & ~n898;
  assign n900 = ~n795 & ~n899;
  assign n901 = pi61  & pi128 ;
  assign n902 = pi62  & ~pi128 ;
  assign n903 = ~pi62  & ~pi128 ;
  assign n904 = ~pi61  & pi128 ;
  assign n905 = ~n903 & ~n904;
  assign n906 = ~n901 & ~n902;
  assign n907 = pi129  & n901;
  assign n908 = pi129  & n902;
  assign n909 = ~n907 & ~n908;
  assign n910 = pi129  & n4665;
  assign n911 = pi64  & ~pi128 ;
  assign n912 = pi63  & pi128 ;
  assign n913 = ~pi63  & pi128 ;
  assign n914 = ~pi64  & ~pi128 ;
  assign n915 = ~n913 & ~n914;
  assign n916 = ~n911 & ~n912;
  assign n917 = ~pi129  & n911;
  assign n918 = ~pi129  & n912;
  assign n919 = ~n917 & ~n918;
  assign n920 = ~pi129  & n4667;
  assign n921 = pi129  & ~n4665;
  assign n922 = ~pi129  & ~n4667;
  assign n923 = ~n921 & ~n922;
  assign n924 = n4666 & n4668;
  assign n925 = n264 & n4669;
  assign n926 = pi57  & pi128 ;
  assign n927 = pi58  & ~pi128 ;
  assign n928 = ~pi58  & ~pi128 ;
  assign n929 = ~pi57  & pi128 ;
  assign n930 = ~n928 & ~n929;
  assign n931 = ~n926 & ~n927;
  assign n932 = pi129  & n926;
  assign n933 = pi129  & n927;
  assign n934 = ~n932 & ~n933;
  assign n935 = pi129  & n4670;
  assign n936 = pi60  & ~pi128 ;
  assign n937 = pi59  & pi128 ;
  assign n938 = ~pi59  & pi128 ;
  assign n939 = ~pi60  & ~pi128 ;
  assign n940 = ~n938 & ~n939;
  assign n941 = ~n936 & ~n937;
  assign n942 = ~pi129  & n936;
  assign n943 = ~pi129  & n937;
  assign n944 = ~n942 & ~n943;
  assign n945 = ~pi129  & n4672;
  assign n946 = pi129  & ~n4670;
  assign n947 = ~pi129  & ~n4672;
  assign n948 = ~n946 & ~n947;
  assign n949 = n4671 & n4673;
  assign n950 = n290 & n4674;
  assign n951 = ~n925 & ~n950;
  assign n952 = pi49  & pi128 ;
  assign n953 = pi50  & ~pi128 ;
  assign n954 = ~pi50  & ~pi128 ;
  assign n955 = ~pi49  & pi128 ;
  assign n956 = ~n954 & ~n955;
  assign n957 = ~n952 & ~n953;
  assign n958 = pi129  & n952;
  assign n959 = pi129  & n953;
  assign n960 = ~n958 & ~n959;
  assign n961 = pi129  & n4675;
  assign n962 = pi52  & ~pi128 ;
  assign n963 = pi51  & pi128 ;
  assign n964 = ~pi51  & pi128 ;
  assign n965 = ~pi52  & ~pi128 ;
  assign n966 = ~n964 & ~n965;
  assign n967 = ~n962 & ~n963;
  assign n968 = ~pi129  & n962;
  assign n969 = ~pi129  & n963;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~pi129  & n4677;
  assign n972 = pi129  & ~n4675;
  assign n973 = ~pi129  & ~n4677;
  assign n974 = ~n972 & ~n973;
  assign n975 = n4676 & n4678;
  assign n976 = n317 & n4679;
  assign n977 = pi53  & pi128 ;
  assign n978 = pi54  & ~pi128 ;
  assign n979 = ~pi54  & ~pi128 ;
  assign n980 = ~pi53  & pi128 ;
  assign n981 = ~n979 & ~n980;
  assign n982 = ~n977 & ~n978;
  assign n983 = pi129  & n977;
  assign n984 = pi129  & n978;
  assign n985 = ~n983 & ~n984;
  assign n986 = pi129  & n4680;
  assign n987 = pi56  & ~pi128 ;
  assign n988 = pi55  & pi128 ;
  assign n989 = ~pi55  & pi128 ;
  assign n990 = ~pi56  & ~pi128 ;
  assign n991 = ~n989 & ~n990;
  assign n992 = ~n987 & ~n988;
  assign n993 = ~pi129  & n987;
  assign n994 = ~pi129  & n988;
  assign n995 = ~n993 & ~n994;
  assign n996 = ~pi129  & n4682;
  assign n997 = pi129  & ~n4680;
  assign n998 = ~pi129  & ~n4682;
  assign n999 = ~n997 & ~n998;
  assign n1000 = n4681 & n4683;
  assign n1001 = n343 & n4684;
  assign n1002 = ~n976 & ~n1001;
  assign n1003 = n951 & n1002;
  assign n1004 = n582 & ~n1003;
  assign n1005 = pi45  & pi128 ;
  assign n1006 = pi46  & ~pi128 ;
  assign n1007 = ~pi46  & ~pi128 ;
  assign n1008 = ~pi45  & pi128 ;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = ~n1005 & ~n1006;
  assign n1011 = pi129  & n1005;
  assign n1012 = pi129  & n1006;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = pi129  & n4685;
  assign n1015 = pi48  & ~pi128 ;
  assign n1016 = pi47  & pi128 ;
  assign n1017 = ~pi47  & pi128 ;
  assign n1018 = ~pi48  & ~pi128 ;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = ~n1015 & ~n1016;
  assign n1021 = ~pi129  & n1015;
  assign n1022 = ~pi129  & n1016;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = ~pi129  & n4687;
  assign n1025 = pi129  & ~n4685;
  assign n1026 = ~pi129  & ~n4687;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = n4686 & n4688;
  assign n1029 = n264 & n4689;
  assign n1030 = pi41  & pi128 ;
  assign n1031 = pi42  & ~pi128 ;
  assign n1032 = ~pi42  & ~pi128 ;
  assign n1033 = ~pi41  & pi128 ;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = ~n1030 & ~n1031;
  assign n1036 = pi129  & n1030;
  assign n1037 = pi129  & n1031;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = pi129  & n4690;
  assign n1040 = pi44  & ~pi128 ;
  assign n1041 = pi43  & pi128 ;
  assign n1042 = ~pi43  & pi128 ;
  assign n1043 = ~pi44  & ~pi128 ;
  assign n1044 = ~n1042 & ~n1043;
  assign n1045 = ~n1040 & ~n1041;
  assign n1046 = ~pi129  & n1040;
  assign n1047 = ~pi129  & n1041;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~pi129  & n4692;
  assign n1050 = pi129  & ~n4690;
  assign n1051 = ~pi129  & ~n4692;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = n4691 & n4693;
  assign n1054 = n290 & n4694;
  assign n1055 = ~n1029 & ~n1054;
  assign n1056 = pi33  & pi128 ;
  assign n1057 = pi34  & ~pi128 ;
  assign n1058 = ~pi34  & ~pi128 ;
  assign n1059 = ~pi33  & pi128 ;
  assign n1060 = ~n1058 & ~n1059;
  assign n1061 = ~n1056 & ~n1057;
  assign n1062 = pi129  & n1056;
  assign n1063 = pi129  & n1057;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = pi129  & n4695;
  assign n1066 = pi36  & ~pi128 ;
  assign n1067 = pi35  & pi128 ;
  assign n1068 = ~pi35  & pi128 ;
  assign n1069 = ~pi36  & ~pi128 ;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = ~n1066 & ~n1067;
  assign n1072 = ~pi129  & n1066;
  assign n1073 = ~pi129  & n1067;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = ~pi129  & n4697;
  assign n1076 = pi129  & ~n4695;
  assign n1077 = ~pi129  & ~n4697;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = n4696 & n4698;
  assign n1080 = n317 & n4699;
  assign n1081 = pi40  & ~pi128 ;
  assign n1082 = ~pi129  & ~n1081;
  assign n1083 = pi37  & pi128 ;
  assign n1084 = pi129  & ~n1083;
  assign n1085 = ~pi129  & n1081;
  assign n1086 = pi129  & n1083;
  assign n1087 = ~n1085 & ~n1086;
  assign n1088 = ~n1082 & ~n1084;
  assign n1089 = pi38  & ~pi128 ;
  assign n1090 = pi129  & n1089;
  assign n1091 = pi39  & pi128 ;
  assign n1092 = ~pi129  & n1091;
  assign n1093 = ~pi129  & ~n1091;
  assign n1094 = pi129  & ~n1089;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = ~n1090 & ~n1092;
  assign n1097 = n4700 & ~n4701;
  assign n1098 = n343 & ~n1097;
  assign n1099 = ~n1080 & ~n1098;
  assign n1100 = n1055 & n1099;
  assign n1101 = n687 & ~n1100;
  assign n1102 = ~n1004 & ~n1101;
  assign n1103 = n900 & n1102;
  assign n1104 = pi134  & ~n1103;
  assign n1105 = ~n691 & ~n1104;
  assign n1106 = pi81  & ~pi128 ;
  assign n1107 = ~pi129  & ~n1106;
  assign n1108 = pi78  & pi128 ;
  assign n1109 = pi129  & ~n1108;
  assign n1110 = ~pi129  & n1106;
  assign n1111 = pi129  & n1108;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = ~n1107 & ~n1109;
  assign n1114 = pi79  & ~pi128 ;
  assign n1115 = pi129  & n1114;
  assign n1116 = pi80  & pi128 ;
  assign n1117 = ~pi129  & n1116;
  assign n1118 = ~pi129  & ~n1116;
  assign n1119 = pi129  & ~n1114;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = ~n1115 & ~n1117;
  assign n1122 = n4702 & ~n4703;
  assign n1123 = n264 & ~n1122;
  assign n1124 = pi77  & ~pi128 ;
  assign n1125 = ~pi129  & ~n1124;
  assign n1126 = pi74  & pi128 ;
  assign n1127 = pi129  & ~n1126;
  assign n1128 = ~pi129  & n1124;
  assign n1129 = pi129  & n1126;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = ~n1125 & ~n1127;
  assign n1132 = pi75  & ~pi128 ;
  assign n1133 = pi129  & n1132;
  assign n1134 = pi76  & pi128 ;
  assign n1135 = ~pi129  & n1134;
  assign n1136 = ~pi129  & ~n1134;
  assign n1137 = pi129  & ~n1132;
  assign n1138 = ~n1136 & ~n1137;
  assign n1139 = ~n1133 & ~n1135;
  assign n1140 = n4704 & ~n4705;
  assign n1141 = n290 & ~n1140;
  assign n1142 = ~n1123 & ~n1141;
  assign n1143 = pi69  & ~pi128 ;
  assign n1144 = ~pi129  & ~n1143;
  assign n1145 = pi66  & pi128 ;
  assign n1146 = pi129  & ~n1145;
  assign n1147 = ~pi129  & n1143;
  assign n1148 = pi129  & n1145;
  assign n1149 = ~n1147 & ~n1148;
  assign n1150 = ~n1144 & ~n1146;
  assign n1151 = pi67  & ~pi128 ;
  assign n1152 = pi129  & n1151;
  assign n1153 = pi68  & pi128 ;
  assign n1154 = ~pi129  & n1153;
  assign n1155 = ~pi129  & ~n1153;
  assign n1156 = pi129  & ~n1151;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~n1152 & ~n1154;
  assign n1159 = n4706 & ~n4707;
  assign n1160 = n317 & ~n1159;
  assign n1161 = pi73  & ~pi128 ;
  assign n1162 = ~pi129  & ~n1161;
  assign n1163 = pi70  & pi128 ;
  assign n1164 = pi129  & ~n1163;
  assign n1165 = ~pi129  & n1161;
  assign n1166 = pi129  & n1163;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~n1162 & ~n1164;
  assign n1169 = pi71  & ~pi128 ;
  assign n1170 = pi129  & n1169;
  assign n1171 = pi72  & pi128 ;
  assign n1172 = ~pi129  & n1171;
  assign n1173 = ~pi129  & ~n1171;
  assign n1174 = pi129  & ~n1169;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = ~n1170 & ~n1172;
  assign n1177 = n4708 & ~n4709;
  assign n1178 = n343 & ~n1177;
  assign n1179 = ~n1160 & ~n1178;
  assign n1180 = n1142 & n1179;
  assign n1181 = n371 & ~n1180;
  assign n1182 = pi97  & ~pi128 ;
  assign n1183 = ~pi129  & ~n1182;
  assign n1184 = pi94  & pi128 ;
  assign n1185 = pi129  & ~n1184;
  assign n1186 = ~pi129  & n1182;
  assign n1187 = pi129  & n1184;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = ~n1183 & ~n1185;
  assign n1190 = pi95  & ~pi128 ;
  assign n1191 = pi129  & n1190;
  assign n1192 = pi96  & pi128 ;
  assign n1193 = ~pi129  & n1192;
  assign n1194 = ~pi129  & ~n1192;
  assign n1195 = pi129  & ~n1190;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = ~n1191 & ~n1193;
  assign n1198 = n4710 & ~n4711;
  assign n1199 = n264 & ~n1198;
  assign n1200 = pi93  & ~pi128 ;
  assign n1201 = ~pi129  & ~n1200;
  assign n1202 = pi90  & pi128 ;
  assign n1203 = pi129  & ~n1202;
  assign n1204 = ~pi129  & n1200;
  assign n1205 = pi129  & n1202;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = ~n1201 & ~n1203;
  assign n1208 = pi91  & ~pi128 ;
  assign n1209 = pi129  & n1208;
  assign n1210 = pi92  & pi128 ;
  assign n1211 = ~pi129  & n1210;
  assign n1212 = ~pi129  & ~n1210;
  assign n1213 = pi129  & ~n1208;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = ~n1209 & ~n1211;
  assign n1216 = n4712 & ~n4713;
  assign n1217 = n290 & ~n1216;
  assign n1218 = ~n1199 & ~n1217;
  assign n1219 = pi85  & ~pi128 ;
  assign n1220 = ~pi129  & ~n1219;
  assign n1221 = pi82  & pi128 ;
  assign n1222 = pi129  & ~n1221;
  assign n1223 = ~pi129  & n1219;
  assign n1224 = pi129  & n1221;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = ~n1220 & ~n1222;
  assign n1227 = pi83  & ~pi128 ;
  assign n1228 = pi129  & n1227;
  assign n1229 = pi84  & pi128 ;
  assign n1230 = ~pi129  & n1229;
  assign n1231 = ~pi129  & ~n1229;
  assign n1232 = pi129  & ~n1227;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = ~n1228 & ~n1230;
  assign n1235 = n4714 & ~n4715;
  assign n1236 = n317 & ~n1235;
  assign n1237 = pi89  & ~pi128 ;
  assign n1238 = ~pi129  & ~n1237;
  assign n1239 = pi86  & pi128 ;
  assign n1240 = pi129  & ~n1239;
  assign n1241 = ~pi129  & n1237;
  assign n1242 = pi129  & n1239;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = ~n1238 & ~n1240;
  assign n1245 = pi87  & ~pi128 ;
  assign n1246 = pi129  & n1245;
  assign n1247 = pi88  & pi128 ;
  assign n1248 = ~pi129  & n1247;
  assign n1249 = ~pi129  & ~n1247;
  assign n1250 = pi129  & ~n1245;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = ~n1246 & ~n1248;
  assign n1253 = n4716 & ~n4717;
  assign n1254 = n343 & ~n1253;
  assign n1255 = ~n1236 & ~n1254;
  assign n1256 = n1218 & n1255;
  assign n1257 = n476 & ~n1256;
  assign n1258 = ~n1181 & ~n1257;
  assign n1259 = pi1  & ~pi128 ;
  assign n1260 = ~pi129  & ~n1259;
  assign n1261 = pi126  & pi128 ;
  assign n1262 = pi129  & ~n1261;
  assign n1263 = ~pi129  & n1259;
  assign n1264 = pi129  & n1261;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = ~n1260 & ~n1262;
  assign n1267 = pi127  & ~pi128 ;
  assign n1268 = pi129  & n1267;
  assign n1269 = pi0  & pi128 ;
  assign n1270 = ~pi129  & n1269;
  assign n1271 = ~pi129  & ~n1269;
  assign n1272 = pi129  & ~n1267;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = ~n1268 & ~n1270;
  assign n1275 = n4718 & ~n4719;
  assign n1276 = n264 & ~n1275;
  assign n1277 = pi125  & ~pi128 ;
  assign n1278 = ~pi129  & ~n1277;
  assign n1279 = pi122  & pi128 ;
  assign n1280 = pi129  & ~n1279;
  assign n1281 = ~pi129  & n1277;
  assign n1282 = pi129  & n1279;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = ~n1278 & ~n1280;
  assign n1285 = pi123  & ~pi128 ;
  assign n1286 = pi129  & n1285;
  assign n1287 = pi124  & pi128 ;
  assign n1288 = ~pi129  & n1287;
  assign n1289 = ~pi129  & ~n1287;
  assign n1290 = pi129  & ~n1285;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292 = ~n1286 & ~n1288;
  assign n1293 = n4720 & ~n4721;
  assign n1294 = n290 & ~n1293;
  assign n1295 = ~n1276 & ~n1294;
  assign n1296 = pi117  & ~pi128 ;
  assign n1297 = ~pi129  & ~n1296;
  assign n1298 = pi114  & pi128 ;
  assign n1299 = pi129  & ~n1298;
  assign n1300 = ~pi129  & n1296;
  assign n1301 = pi129  & n1298;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = ~n1297 & ~n1299;
  assign n1304 = pi115  & ~pi128 ;
  assign n1305 = pi129  & n1304;
  assign n1306 = pi116  & pi128 ;
  assign n1307 = ~pi129  & n1306;
  assign n1308 = ~pi129  & ~n1306;
  assign n1309 = pi129  & ~n1304;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~n1305 & ~n1307;
  assign n1312 = n4722 & ~n4723;
  assign n1313 = n317 & ~n1312;
  assign n1314 = pi121  & ~pi128 ;
  assign n1315 = ~pi129  & ~n1314;
  assign n1316 = pi118  & pi128 ;
  assign n1317 = pi129  & ~n1316;
  assign n1318 = ~pi129  & n1314;
  assign n1319 = pi129  & n1316;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321 = ~n1315 & ~n1317;
  assign n1322 = pi119  & ~pi128 ;
  assign n1323 = pi129  & n1322;
  assign n1324 = pi120  & pi128 ;
  assign n1325 = ~pi129  & n1324;
  assign n1326 = ~pi129  & ~n1324;
  assign n1327 = pi129  & ~n1322;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1323 & ~n1325;
  assign n1330 = n4724 & ~n4725;
  assign n1331 = n343 & ~n1330;
  assign n1332 = ~n1313 & ~n1331;
  assign n1333 = n1295 & n1332;
  assign n1334 = n582 & ~n1333;
  assign n1335 = pi113  & ~pi128 ;
  assign n1336 = ~pi129  & ~n1335;
  assign n1337 = pi110  & pi128 ;
  assign n1338 = pi129  & ~n1337;
  assign n1339 = ~pi129  & n1335;
  assign n1340 = pi129  & n1337;
  assign n1341 = ~n1339 & ~n1340;
  assign n1342 = ~n1336 & ~n1338;
  assign n1343 = pi111  & ~pi128 ;
  assign n1344 = pi129  & n1343;
  assign n1345 = pi112  & pi128 ;
  assign n1346 = ~pi129  & n1345;
  assign n1347 = ~pi129  & ~n1345;
  assign n1348 = pi129  & ~n1343;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = ~n1344 & ~n1346;
  assign n1351 = n4726 & ~n4727;
  assign n1352 = n264 & ~n1351;
  assign n1353 = pi109  & ~pi128 ;
  assign n1354 = ~pi129  & ~n1353;
  assign n1355 = pi106  & pi128 ;
  assign n1356 = pi129  & ~n1355;
  assign n1357 = ~pi129  & n1353;
  assign n1358 = pi129  & n1355;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = ~n1354 & ~n1356;
  assign n1361 = pi107  & ~pi128 ;
  assign n1362 = pi129  & n1361;
  assign n1363 = pi108  & pi128 ;
  assign n1364 = ~pi129  & n1363;
  assign n1365 = ~pi129  & ~n1363;
  assign n1366 = pi129  & ~n1361;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = ~n1362 & ~n1364;
  assign n1369 = n4728 & ~n4729;
  assign n1370 = n290 & ~n1369;
  assign n1371 = ~n1352 & ~n1370;
  assign n1372 = pi101  & ~pi128 ;
  assign n1373 = ~pi129  & ~n1372;
  assign n1374 = pi98  & pi128 ;
  assign n1375 = pi129  & ~n1374;
  assign n1376 = ~pi129  & n1372;
  assign n1377 = pi129  & n1374;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = ~n1373 & ~n1375;
  assign n1380 = pi99  & ~pi128 ;
  assign n1381 = pi129  & n1380;
  assign n1382 = pi100  & pi128 ;
  assign n1383 = ~pi129  & n1382;
  assign n1384 = ~pi129  & ~n1382;
  assign n1385 = pi129  & ~n1380;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = ~n1381 & ~n1383;
  assign n1388 = n4730 & ~n4731;
  assign n1389 = n317 & ~n1388;
  assign n1390 = pi105  & ~pi128 ;
  assign n1391 = ~pi129  & ~n1390;
  assign n1392 = pi102  & pi128 ;
  assign n1393 = pi129  & ~n1392;
  assign n1394 = ~pi129  & n1390;
  assign n1395 = pi129  & n1392;
  assign n1396 = ~n1394 & ~n1395;
  assign n1397 = ~n1391 & ~n1393;
  assign n1398 = pi103  & ~pi128 ;
  assign n1399 = pi129  & n1398;
  assign n1400 = pi104  & pi128 ;
  assign n1401 = ~pi129  & n1400;
  assign n1402 = ~pi129  & ~n1400;
  assign n1403 = pi129  & ~n1398;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~n1399 & ~n1401;
  assign n1406 = n4732 & ~n4733;
  assign n1407 = n343 & ~n1406;
  assign n1408 = ~n1389 & ~n1407;
  assign n1409 = n1371 & n1408;
  assign n1410 = n687 & ~n1409;
  assign n1411 = ~n1334 & ~n1410;
  assign n1412 = n1258 & n1411;
  assign n1413 = ~pi134  & ~n1412;
  assign n1414 = pi65  & ~pi128 ;
  assign n1415 = ~pi129  & ~n1414;
  assign n1416 = pi62  & pi128 ;
  assign n1417 = pi129  & ~n1416;
  assign n1418 = ~pi129  & n1414;
  assign n1419 = pi129  & n1416;
  assign n1420 = ~n1418 & ~n1419;
  assign n1421 = ~n1415 & ~n1417;
  assign n1422 = pi63  & ~pi128 ;
  assign n1423 = pi129  & n1422;
  assign n1424 = pi64  & pi128 ;
  assign n1425 = ~pi129  & n1424;
  assign n1426 = ~pi129  & ~n1424;
  assign n1427 = pi129  & ~n1422;
  assign n1428 = ~n1426 & ~n1427;
  assign n1429 = ~n1423 & ~n1425;
  assign n1430 = n4734 & ~n4735;
  assign n1431 = n264 & ~n1430;
  assign n1432 = pi61  & ~pi128 ;
  assign n1433 = ~pi129  & ~n1432;
  assign n1434 = pi58  & pi128 ;
  assign n1435 = pi129  & ~n1434;
  assign n1436 = ~pi129  & n1432;
  assign n1437 = pi129  & n1434;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = ~n1433 & ~n1435;
  assign n1440 = pi59  & ~pi128 ;
  assign n1441 = pi129  & n1440;
  assign n1442 = pi60  & pi128 ;
  assign n1443 = ~pi129  & n1442;
  assign n1444 = ~pi129  & ~n1442;
  assign n1445 = pi129  & ~n1440;
  assign n1446 = ~n1444 & ~n1445;
  assign n1447 = ~n1441 & ~n1443;
  assign n1448 = n4736 & ~n4737;
  assign n1449 = n290 & ~n1448;
  assign n1450 = ~n1431 & ~n1449;
  assign n1451 = pi53  & ~pi128 ;
  assign n1452 = ~pi129  & ~n1451;
  assign n1453 = pi50  & pi128 ;
  assign n1454 = pi129  & ~n1453;
  assign n1455 = ~pi129  & n1451;
  assign n1456 = pi129  & n1453;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = ~n1452 & ~n1454;
  assign n1459 = pi51  & ~pi128 ;
  assign n1460 = pi129  & n1459;
  assign n1461 = pi52  & pi128 ;
  assign n1462 = ~pi129  & n1461;
  assign n1463 = ~pi129  & ~n1461;
  assign n1464 = pi129  & ~n1459;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = ~n1460 & ~n1462;
  assign n1467 = n4738 & ~n4739;
  assign n1468 = n317 & ~n1467;
  assign n1469 = pi57  & ~pi128 ;
  assign n1470 = ~pi129  & ~n1469;
  assign n1471 = pi54  & pi128 ;
  assign n1472 = pi129  & ~n1471;
  assign n1473 = ~pi129  & n1469;
  assign n1474 = pi129  & n1471;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = ~n1470 & ~n1472;
  assign n1477 = pi55  & ~pi128 ;
  assign n1478 = pi129  & n1477;
  assign n1479 = pi56  & pi128 ;
  assign n1480 = ~pi129  & n1479;
  assign n1481 = ~pi129  & ~n1479;
  assign n1482 = pi129  & ~n1477;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = ~n1478 & ~n1480;
  assign n1485 = n4740 & ~n4741;
  assign n1486 = n343 & ~n1485;
  assign n1487 = ~n1468 & ~n1486;
  assign n1488 = n1450 & n1487;
  assign n1489 = n582 & ~n1488;
  assign n1490 = pi17  & ~pi128 ;
  assign n1491 = ~pi129  & ~n1490;
  assign n1492 = pi14  & pi128 ;
  assign n1493 = pi129  & ~n1492;
  assign n1494 = ~pi129  & n1490;
  assign n1495 = pi129  & n1492;
  assign n1496 = ~n1494 & ~n1495;
  assign n1497 = ~n1491 & ~n1493;
  assign n1498 = pi15  & ~pi128 ;
  assign n1499 = pi129  & n1498;
  assign n1500 = pi16  & pi128 ;
  assign n1501 = ~pi129  & n1500;
  assign n1502 = ~pi129  & ~n1500;
  assign n1503 = pi129  & ~n1498;
  assign n1504 = ~n1502 & ~n1503;
  assign n1505 = ~n1499 & ~n1501;
  assign n1506 = n4742 & ~n4743;
  assign n1507 = n264 & ~n1506;
  assign n1508 = pi13  & ~pi128 ;
  assign n1509 = ~pi129  & ~n1508;
  assign n1510 = pi10  & pi128 ;
  assign n1511 = pi129  & ~n1510;
  assign n1512 = ~pi129  & n1508;
  assign n1513 = pi129  & n1510;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = ~n1509 & ~n1511;
  assign n1516 = pi11  & ~pi128 ;
  assign n1517 = pi129  & n1516;
  assign n1518 = pi12  & pi128 ;
  assign n1519 = ~pi129  & n1518;
  assign n1520 = ~pi129  & ~n1518;
  assign n1521 = pi129  & ~n1516;
  assign n1522 = ~n1520 & ~n1521;
  assign n1523 = ~n1517 & ~n1519;
  assign n1524 = n4744 & ~n4745;
  assign n1525 = n290 & ~n1524;
  assign n1526 = ~n1507 & ~n1525;
  assign n1527 = pi5  & ~pi128 ;
  assign n1528 = ~pi129  & ~n1527;
  assign n1529 = pi2  & pi128 ;
  assign n1530 = pi129  & ~n1529;
  assign n1531 = ~pi129  & n1527;
  assign n1532 = pi129  & n1529;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = ~n1528 & ~n1530;
  assign n1535 = pi3  & ~pi128 ;
  assign n1536 = pi129  & n1535;
  assign n1537 = pi4  & pi128 ;
  assign n1538 = ~pi129  & n1537;
  assign n1539 = ~pi129  & ~n1537;
  assign n1540 = pi129  & ~n1535;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = ~n1536 & ~n1538;
  assign n1543 = n4746 & ~n4747;
  assign n1544 = n317 & ~n1543;
  assign n1545 = pi9  & ~pi128 ;
  assign n1546 = ~pi129  & ~n1545;
  assign n1547 = pi6  & pi128 ;
  assign n1548 = pi129  & ~n1547;
  assign n1549 = ~pi129  & n1545;
  assign n1550 = pi129  & n1547;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = ~n1546 & ~n1548;
  assign n1553 = pi7  & ~pi128 ;
  assign n1554 = pi129  & n1553;
  assign n1555 = pi8  & pi128 ;
  assign n1556 = ~pi129  & n1555;
  assign n1557 = ~pi129  & ~n1555;
  assign n1558 = pi129  & ~n1553;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = ~n1554 & ~n1556;
  assign n1561 = n4748 & ~n4749;
  assign n1562 = n343 & ~n1561;
  assign n1563 = ~n1544 & ~n1562;
  assign n1564 = n1526 & n1563;
  assign n1565 = n371 & ~n1564;
  assign n1566 = ~n1489 & ~n1565;
  assign n1567 = pi49  & ~pi128 ;
  assign n1568 = ~pi129  & ~n1567;
  assign n1569 = pi46  & pi128 ;
  assign n1570 = pi129  & ~n1569;
  assign n1571 = ~pi129  & n1567;
  assign n1572 = pi129  & n1569;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = ~n1568 & ~n1570;
  assign n1575 = pi47  & ~pi128 ;
  assign n1576 = pi129  & n1575;
  assign n1577 = pi48  & pi128 ;
  assign n1578 = ~pi129  & n1577;
  assign n1579 = ~pi129  & ~n1577;
  assign n1580 = pi129  & ~n1575;
  assign n1581 = ~n1579 & ~n1580;
  assign n1582 = ~n1576 & ~n1578;
  assign n1583 = n4750 & ~n4751;
  assign n1584 = n264 & ~n1583;
  assign n1585 = pi42  & pi128 ;
  assign n1586 = pi43  & ~pi128 ;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = pi129  & n1585;
  assign n1589 = pi129  & n1586;
  assign n1590 = ~n1588 & ~n1589;
  assign n1591 = pi129  & ~n1587;
  assign n1592 = pi45  & ~pi128 ;
  assign n1593 = pi44  & pi128 ;
  assign n1594 = ~pi44  & pi128 ;
  assign n1595 = ~pi45  & ~pi128 ;
  assign n1596 = ~n1594 & ~n1595;
  assign n1597 = ~n1592 & ~n1593;
  assign n1598 = ~pi129  & n1592;
  assign n1599 = ~pi129  & n1593;
  assign n1600 = ~n1598 & ~n1599;
  assign n1601 = ~pi129  & n4753;
  assign n1602 = n4752 & n4754;
  assign n1603 = n290 & ~n1602;
  assign n1604 = ~n1584 & ~n1603;
  assign n1605 = pi37  & ~pi128 ;
  assign n1606 = ~pi129  & ~n1605;
  assign n1607 = pi34  & pi128 ;
  assign n1608 = pi129  & ~n1607;
  assign n1609 = ~pi129  & n1605;
  assign n1610 = pi129  & n1607;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = ~n1606 & ~n1608;
  assign n1613 = pi35  & ~pi128 ;
  assign n1614 = pi129  & n1613;
  assign n1615 = pi36  & pi128 ;
  assign n1616 = ~pi129  & n1615;
  assign n1617 = ~pi129  & ~n1615;
  assign n1618 = pi129  & ~n1613;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = ~n1614 & ~n1616;
  assign n1621 = n4755 & ~n4756;
  assign n1622 = n317 & ~n1621;
  assign n1623 = pi41  & ~pi128 ;
  assign n1624 = pi40  & pi128 ;
  assign n1625 = ~n1623 & ~n1624;
  assign n1626 = ~pi129  & n1623;
  assign n1627 = ~pi129  & n1624;
  assign n1628 = ~n1626 & ~n1627;
  assign n1629 = ~pi129  & ~n1625;
  assign n1630 = pi39  & ~pi128 ;
  assign n1631 = pi38  & pi128 ;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = pi129  & n1630;
  assign n1634 = pi129  & n1631;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = pi129  & ~n1632;
  assign n1637 = n4757 & n4758;
  assign n1638 = n343 & ~n1637;
  assign n1639 = ~n1622 & ~n1638;
  assign n1640 = n1604 & n1639;
  assign n1641 = n687 & ~n1640;
  assign n1642 = pi33  & ~pi128 ;
  assign n1643 = ~pi129  & ~n1642;
  assign n1644 = pi30  & pi128 ;
  assign n1645 = pi129  & ~n1644;
  assign n1646 = ~pi129  & n1642;
  assign n1647 = pi129  & n1644;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = ~n1643 & ~n1645;
  assign n1650 = pi31  & ~pi128 ;
  assign n1651 = pi129  & n1650;
  assign n1652 = pi32  & pi128 ;
  assign n1653 = ~pi129  & n1652;
  assign n1654 = ~pi129  & ~n1652;
  assign n1655 = pi129  & ~n1650;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = ~n1651 & ~n1653;
  assign n1658 = n4759 & ~n4760;
  assign n1659 = n264 & ~n1658;
  assign n1660 = pi29  & ~pi128 ;
  assign n1661 = ~pi129  & ~n1660;
  assign n1662 = pi26  & pi128 ;
  assign n1663 = pi129  & ~n1662;
  assign n1664 = ~pi129  & n1660;
  assign n1665 = pi129  & n1662;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = ~n1661 & ~n1663;
  assign n1668 = pi27  & ~pi128 ;
  assign n1669 = pi129  & n1668;
  assign n1670 = pi28  & pi128 ;
  assign n1671 = ~pi129  & n1670;
  assign n1672 = ~pi129  & ~n1670;
  assign n1673 = pi129  & ~n1668;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = ~n1669 & ~n1671;
  assign n1676 = n4761 & ~n4762;
  assign n1677 = n290 & ~n1676;
  assign n1678 = ~n1659 & ~n1677;
  assign n1679 = pi21  & ~pi128 ;
  assign n1680 = ~pi129  & ~n1679;
  assign n1681 = pi18  & pi128 ;
  assign n1682 = pi129  & ~n1681;
  assign n1683 = ~pi129  & n1679;
  assign n1684 = pi129  & n1681;
  assign n1685 = ~n1683 & ~n1684;
  assign n1686 = ~n1680 & ~n1682;
  assign n1687 = pi19  & ~pi128 ;
  assign n1688 = pi129  & n1687;
  assign n1689 = pi20  & pi128 ;
  assign n1690 = ~pi129  & n1689;
  assign n1691 = ~pi129  & ~n1689;
  assign n1692 = pi129  & ~n1687;
  assign n1693 = ~n1691 & ~n1692;
  assign n1694 = ~n1688 & ~n1690;
  assign n1695 = n4763 & ~n4764;
  assign n1696 = n317 & ~n1695;
  assign n1697 = pi25  & ~pi128 ;
  assign n1698 = ~pi129  & ~n1697;
  assign n1699 = pi22  & pi128 ;
  assign n1700 = pi129  & ~n1699;
  assign n1701 = ~pi129  & n1697;
  assign n1702 = pi129  & n1699;
  assign n1703 = ~n1701 & ~n1702;
  assign n1704 = ~n1698 & ~n1700;
  assign n1705 = pi23  & ~pi128 ;
  assign n1706 = pi129  & n1705;
  assign n1707 = pi24  & pi128 ;
  assign n1708 = ~pi129  & n1707;
  assign n1709 = ~pi129  & ~n1707;
  assign n1710 = pi129  & ~n1705;
  assign n1711 = ~n1709 & ~n1710;
  assign n1712 = ~n1706 & ~n1708;
  assign n1713 = n4765 & ~n4766;
  assign n1714 = n343 & ~n1713;
  assign n1715 = ~n1696 & ~n1714;
  assign n1716 = n1678 & n1715;
  assign n1717 = n476 & ~n1716;
  assign n1718 = ~n1641 & ~n1717;
  assign n1719 = n1566 & n1718;
  assign n1720 = pi134  & ~n1719;
  assign n1721 = ~n1413 & ~n1720;
  assign n1722 = pi129  & n275;
  assign n1723 = pi129  & n276;
  assign n1724 = ~n1722 & ~n1723;
  assign n1725 = pi129  & n4547;
  assign n1726 = ~pi129  & n424;
  assign n1727 = ~pi129  & n425;
  assign n1728 = ~n1726 & ~n1727;
  assign n1729 = ~pi129  & n4575;
  assign n1730 = pi129  & ~n4547;
  assign n1731 = ~pi129  & ~n4575;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = n4767 & n4768;
  assign n1734 = n264 & n4769;
  assign n1735 = pi129  & n301;
  assign n1736 = pi129  & n302;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = pi129  & n4552;
  assign n1739 = ~pi129  & n265;
  assign n1740 = ~pi129  & n266;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = ~pi129  & n4545;
  assign n1743 = pi129  & ~n4552;
  assign n1744 = ~pi129  & ~n4545;
  assign n1745 = ~n1743 & ~n1744;
  assign n1746 = n4770 & n4771;
  assign n1747 = n290 & n4772;
  assign n1748 = ~n1734 & ~n1747;
  assign n1749 = pi129  & n328;
  assign n1750 = pi129  & n329;
  assign n1751 = ~n1749 & ~n1750;
  assign n1752 = pi129  & n4557;
  assign n1753 = ~pi129  & n344;
  assign n1754 = ~pi129  & n345;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = ~pi129  & n4560;
  assign n1757 = pi129  & ~n4557;
  assign n1758 = ~pi129  & ~n4560;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = n4773 & n4774;
  assign n1761 = n317 & n4775;
  assign n1762 = pi129  & n354;
  assign n1763 = pi129  & n355;
  assign n1764 = ~n1762 & ~n1763;
  assign n1765 = pi129  & n4562;
  assign n1766 = ~pi129  & n291;
  assign n1767 = ~pi129  & n292;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = ~pi129  & n4550;
  assign n1770 = pi129  & ~n4562;
  assign n1771 = ~pi129  & ~n4550;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = n4776 & n4777;
  assign n1774 = n343 & n4778;
  assign n1775 = ~n1761 & ~n1774;
  assign n1776 = n1748 & n1775;
  assign n1777 = n371 & ~n1776;
  assign n1778 = pi129  & n383;
  assign n1779 = pi129  & n384;
  assign n1780 = ~n1778 & ~n1779;
  assign n1781 = pi129  & n4567;
  assign n1782 = ~pi129  & n635;
  assign n1783 = ~pi129  & n636;
  assign n1784 = ~n1782 & ~n1783;
  assign n1785 = ~pi129  & n4615;
  assign n1786 = pi129  & ~n4567;
  assign n1787 = ~pi129  & ~n4615;
  assign n1788 = ~n1786 & ~n1787;
  assign n1789 = n4779 & n4780;
  assign n1790 = n264 & n4781;
  assign n1791 = pi129  & n408;
  assign n1792 = pi129  & n409;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = pi129  & n4572;
  assign n1795 = ~pi129  & n373;
  assign n1796 = ~pi129  & n374;
  assign n1797 = ~n1795 & ~n1796;
  assign n1798 = ~pi129  & n4565;
  assign n1799 = pi129  & ~n4572;
  assign n1800 = ~pi129  & ~n4565;
  assign n1801 = ~n1799 & ~n1800;
  assign n1802 = n4782 & n4783;
  assign n1803 = n290 & n4784;
  assign n1804 = ~n1790 & ~n1803;
  assign n1805 = pi129  & n434;
  assign n1806 = pi129  & n435;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = pi129  & n4577;
  assign n1809 = ~pi129  & n449;
  assign n1810 = ~pi129  & n450;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = ~pi129  & n4580;
  assign n1813 = pi129  & ~n4577;
  assign n1814 = ~pi129  & ~n4580;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = n4785 & n4786;
  assign n1817 = n317 & n4787;
  assign n1818 = pi129  & n459;
  assign n1819 = pi129  & n460;
  assign n1820 = ~n1818 & ~n1819;
  assign n1821 = pi129  & n4582;
  assign n1822 = ~pi129  & n398;
  assign n1823 = ~pi129  & n399;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = ~pi129  & n4570;
  assign n1826 = pi129  & ~n4582;
  assign n1827 = ~pi129  & ~n4570;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = n4788 & n4789;
  assign n1830 = n343 & n4790;
  assign n1831 = ~n1817 & ~n1830;
  assign n1832 = n1804 & n1831;
  assign n1833 = n476 & ~n1832;
  assign n1834 = ~n1777 & ~n1833;
  assign n1835 = pi129  & n489;
  assign n1836 = pi129  & n490;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = pi129  & n4587;
  assign n1839 = ~pi129  & n743;
  assign n1840 = ~pi129  & n744;
  assign n1841 = ~n1839 & ~n1840;
  assign n1842 = ~pi129  & n4635;
  assign n1843 = pi129  & ~n4587;
  assign n1844 = ~pi129  & ~n4635;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = n4791 & n4792;
  assign n1847 = n264 & n4793;
  assign n1848 = pi129  & n514;
  assign n1849 = pi129  & n515;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = pi129  & n4592;
  assign n1852 = ~pi129  & n479;
  assign n1853 = ~pi129  & n480;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = ~pi129  & n4585;
  assign n1856 = pi129  & ~n4592;
  assign n1857 = ~pi129  & ~n4585;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = n4794 & n4795;
  assign n1860 = n290 & n4796;
  assign n1861 = ~n1847 & ~n1860;
  assign n1862 = pi129  & n540;
  assign n1863 = pi129  & n541;
  assign n1864 = ~n1862 & ~n1863;
  assign n1865 = pi129  & n4597;
  assign n1866 = ~pi129  & n555;
  assign n1867 = ~pi129  & n556;
  assign n1868 = ~n1866 & ~n1867;
  assign n1869 = ~pi129  & n4600;
  assign n1870 = pi129  & ~n4597;
  assign n1871 = ~pi129  & ~n4600;
  assign n1872 = ~n1870 & ~n1871;
  assign n1873 = n4797 & n4798;
  assign n1874 = n317 & n4799;
  assign n1875 = pi129  & n565;
  assign n1876 = pi129  & n566;
  assign n1877 = ~n1875 & ~n1876;
  assign n1878 = pi129  & n4602;
  assign n1879 = ~pi129  & n504;
  assign n1880 = ~pi129  & n505;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = ~pi129  & n4590;
  assign n1883 = pi129  & ~n4602;
  assign n1884 = ~pi129  & ~n4590;
  assign n1885 = ~n1883 & ~n1884;
  assign n1886 = n4800 & n4801;
  assign n1887 = n343 & n4802;
  assign n1888 = ~n1874 & ~n1887;
  assign n1889 = n1861 & n1888;
  assign n1890 = n582 & ~n1889;
  assign n1891 = pi129  & n594;
  assign n1892 = pi129  & n595;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = pi129  & n4607;
  assign n1895 = ~pi129  & n530;
  assign n1896 = ~pi129  & n531;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = ~pi129  & n4595;
  assign n1899 = pi129  & ~n4607;
  assign n1900 = ~pi129  & ~n4595;
  assign n1901 = ~n1899 & ~n1900;
  assign n1902 = n4803 & n4804;
  assign n1903 = n264 & n4805;
  assign n1904 = pi129  & n619;
  assign n1905 = pi129  & n620;
  assign n1906 = ~n1904 & ~n1905;
  assign n1907 = pi129  & n4612;
  assign n1908 = ~pi129  & n584;
  assign n1909 = ~pi129  & n585;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = ~pi129  & n4605;
  assign n1912 = pi129  & ~n4612;
  assign n1913 = ~pi129  & ~n4605;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = n4806 & n4807;
  assign n1916 = n290 & n4808;
  assign n1917 = ~n1903 & ~n1916;
  assign n1918 = pi129  & n645;
  assign n1919 = pi129  & n646;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = pi129  & n4617;
  assign n1922 = ~pi129  & n660;
  assign n1923 = ~pi129  & n661;
  assign n1924 = ~n1922 & ~n1923;
  assign n1925 = ~pi129  & n4620;
  assign n1926 = pi129  & ~n4617;
  assign n1927 = ~pi129  & ~n4620;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = n4809 & n4810;
  assign n1930 = n317 & n4811;
  assign n1931 = pi129  & n670;
  assign n1932 = pi129  & n671;
  assign n1933 = ~n1931 & ~n1932;
  assign n1934 = pi129  & n4622;
  assign n1935 = ~pi129  & n609;
  assign n1936 = ~pi129  & n610;
  assign n1937 = ~n1935 & ~n1936;
  assign n1938 = ~pi129  & n4610;
  assign n1939 = pi129  & ~n4622;
  assign n1940 = ~pi129  & ~n4610;
  assign n1941 = ~n1939 & ~n1940;
  assign n1942 = n4812 & n4813;
  assign n1943 = n343 & n4814;
  assign n1944 = ~n1930 & ~n1943;
  assign n1945 = n1917 & n1944;
  assign n1946 = n687 & ~n1945;
  assign n1947 = ~n1890 & ~n1946;
  assign n1948 = n1834 & n1947;
  assign n1949 = ~pi134  & ~n1948;
  assign n1950 = pi129  & n911;
  assign n1951 = pi129  & n912;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = pi129  & n4667;
  assign n1954 = ~pi129  & n318;
  assign n1955 = ~pi129  & n319;
  assign n1956 = ~n1954 & ~n1955;
  assign n1957 = ~pi129  & n4555;
  assign n1958 = pi129  & ~n4667;
  assign n1959 = ~pi129  & ~n4555;
  assign n1960 = ~n1958 & ~n1959;
  assign n1961 = n4815 & n4816;
  assign n1962 = n264 & n4817;
  assign n1963 = pi129  & n936;
  assign n1964 = pi129  & n937;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = pi129  & n4672;
  assign n1967 = ~pi129  & n901;
  assign n1968 = ~pi129  & n902;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = ~pi129  & n4665;
  assign n1971 = pi129  & ~n4672;
  assign n1972 = ~pi129  & ~n4665;
  assign n1973 = ~n1971 & ~n1972;
  assign n1974 = n4818 & n4819;
  assign n1975 = n290 & n4820;
  assign n1976 = ~n1962 & ~n1975;
  assign n1977 = pi129  & n962;
  assign n1978 = pi129  & n963;
  assign n1979 = ~n1977 & ~n1978;
  assign n1980 = pi129  & n4677;
  assign n1981 = ~pi129  & n977;
  assign n1982 = ~pi129  & n978;
  assign n1983 = ~n1981 & ~n1982;
  assign n1984 = ~pi129  & n4680;
  assign n1985 = pi129  & ~n4677;
  assign n1986 = ~pi129  & ~n4680;
  assign n1987 = ~n1985 & ~n1986;
  assign n1988 = n4821 & n4822;
  assign n1989 = n317 & n4823;
  assign n1990 = pi129  & n987;
  assign n1991 = pi129  & n988;
  assign n1992 = ~n1990 & ~n1991;
  assign n1993 = pi129  & n4682;
  assign n1994 = ~pi129  & n926;
  assign n1995 = ~pi129  & n927;
  assign n1996 = ~n1994 & ~n1995;
  assign n1997 = ~pi129  & n4670;
  assign n1998 = pi129  & ~n4682;
  assign n1999 = ~pi129  & ~n4670;
  assign n2000 = ~n1998 & ~n1999;
  assign n2001 = n4824 & n4825;
  assign n2002 = n343 & n4826;
  assign n2003 = ~n1989 & ~n2002;
  assign n2004 = n1976 & n2003;
  assign n2005 = n582 & ~n2004;
  assign n2006 = pi129  & n702;
  assign n2007 = pi129  & n703;
  assign n2008 = ~n2006 & ~n2007;
  assign n2009 = pi129  & n4627;
  assign n2010 = ~pi129  & n847;
  assign n2011 = ~pi129  & n848;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = ~pi129  & n4655;
  assign n2014 = pi129  & ~n4627;
  assign n2015 = ~pi129  & ~n4655;
  assign n2016 = ~n2014 & ~n2015;
  assign n2017 = n4827 & n4828;
  assign n2018 = n264 & n4829;
  assign n2019 = pi129  & n727;
  assign n2020 = pi129  & n728;
  assign n2021 = ~n2019 & ~n2020;
  assign n2022 = pi129  & n4632;
  assign n2023 = ~pi129  & n692;
  assign n2024 = ~pi129  & n693;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = ~pi129  & n4625;
  assign n2027 = pi129  & ~n4632;
  assign n2028 = ~pi129  & ~n4625;
  assign n2029 = ~n2027 & ~n2028;
  assign n2030 = n4830 & n4831;
  assign n2031 = n290 & n4832;
  assign n2032 = ~n2018 & ~n2031;
  assign n2033 = pi129  & n753;
  assign n2034 = pi129  & n754;
  assign n2035 = ~n2033 & ~n2034;
  assign n2036 = pi129  & n4637;
  assign n2037 = ~pi129  & n768;
  assign n2038 = ~pi129  & n769;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = ~pi129  & n4640;
  assign n2041 = pi129  & ~n4637;
  assign n2042 = ~pi129  & ~n4640;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = n4833 & n4834;
  assign n2045 = n317 & n4835;
  assign n2046 = pi129  & n778;
  assign n2047 = pi129  & n779;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = pi129  & n4642;
  assign n2050 = ~pi129  & n717;
  assign n2051 = ~pi129  & n718;
  assign n2052 = ~n2050 & ~n2051;
  assign n2053 = ~pi129  & n4630;
  assign n2054 = pi129  & ~n4642;
  assign n2055 = ~pi129  & ~n4630;
  assign n2056 = ~n2054 & ~n2055;
  assign n2057 = n4836 & n4837;
  assign n2058 = n343 & n4838;
  assign n2059 = ~n2045 & ~n2058;
  assign n2060 = n2032 & n2059;
  assign n2061 = n371 & ~n2060;
  assign n2062 = ~n2005 & ~n2061;
  assign n2063 = pi129  & n1015;
  assign n2064 = pi129  & n1016;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = pi129  & n4687;
  assign n2067 = ~pi129  & n952;
  assign n2068 = ~pi129  & n953;
  assign n2069 = ~n2067 & ~n2068;
  assign n2070 = ~pi129  & n4675;
  assign n2071 = pi129  & ~n4687;
  assign n2072 = ~pi129  & ~n4675;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = n4839 & n4840;
  assign n2075 = n264 & n4841;
  assign n2076 = pi129  & n1041;
  assign n2077 = pi129  & n1040;
  assign n2078 = ~n2076 & ~n2077;
  assign n2079 = pi129  & n4692;
  assign n2080 = ~pi129  & n1006;
  assign n2081 = ~pi129  & n1005;
  assign n2082 = ~n2080 & ~n2081;
  assign n2083 = ~pi129  & n4685;
  assign n2084 = pi129  & ~n4692;
  assign n2085 = ~pi129  & ~n4685;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = n4842 & n4843;
  assign n2088 = n290 & n4844;
  assign n2089 = ~n2075 & ~n2088;
  assign n2090 = ~n1083 & ~n1089;
  assign n2091 = ~pi129  & n1083;
  assign n2092 = ~pi129  & n1089;
  assign n2093 = ~n2091 & ~n2092;
  assign n2094 = ~pi129  & ~n2090;
  assign n2095 = pi129  & n1066;
  assign n2096 = pi129  & n1067;
  assign n2097 = ~n2095 & ~n2096;
  assign n2098 = pi129  & n4697;
  assign n2099 = n4845 & n4846;
  assign n2100 = n317 & ~n2099;
  assign n2101 = ~pi129  & n1030;
  assign n2102 = ~pi129  & n1031;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = ~pi129  & n4690;
  assign n2105 = ~n1081 & ~n1091;
  assign n2106 = pi129  & n1091;
  assign n2107 = pi129  & n1081;
  assign n2108 = ~n2106 & ~n2107;
  assign n2109 = pi129  & ~n2105;
  assign n2110 = n4847 & n4848;
  assign n2111 = n343 & ~n2110;
  assign n2112 = ~n2100 & ~n2111;
  assign n2113 = n2089 & n2112;
  assign n2114 = n687 & ~n2113;
  assign n2115 = pi129  & n806;
  assign n2116 = pi129  & n807;
  assign n2117 = ~n2115 & ~n2116;
  assign n2118 = pi129  & n4647;
  assign n2119 = ~pi129  & n1056;
  assign n2120 = ~pi129  & n1057;
  assign n2121 = ~n2119 & ~n2120;
  assign n2122 = ~pi129  & n4695;
  assign n2123 = pi129  & ~n4647;
  assign n2124 = ~pi129  & ~n4695;
  assign n2125 = ~n2123 & ~n2124;
  assign n2126 = n4849 & n4850;
  assign n2127 = n264 & n4851;
  assign n2128 = pi129  & n831;
  assign n2129 = pi129  & n832;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = pi129  & n4652;
  assign n2132 = ~pi129  & n796;
  assign n2133 = ~pi129  & n797;
  assign n2134 = ~n2132 & ~n2133;
  assign n2135 = ~pi129  & n4645;
  assign n2136 = pi129  & ~n4652;
  assign n2137 = ~pi129  & ~n4645;
  assign n2138 = ~n2136 & ~n2137;
  assign n2139 = n4852 & n4853;
  assign n2140 = n290 & n4854;
  assign n2141 = ~n2127 & ~n2140;
  assign n2142 = pi129  & n857;
  assign n2143 = pi129  & n858;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = pi129  & n4657;
  assign n2146 = ~pi129  & n872;
  assign n2147 = ~pi129  & n873;
  assign n2148 = ~n2146 & ~n2147;
  assign n2149 = ~pi129  & n4660;
  assign n2150 = pi129  & ~n4657;
  assign n2151 = ~pi129  & ~n4660;
  assign n2152 = ~n2150 & ~n2151;
  assign n2153 = n4855 & n4856;
  assign n2154 = n317 & n4857;
  assign n2155 = pi129  & n882;
  assign n2156 = pi129  & n883;
  assign n2157 = ~n2155 & ~n2156;
  assign n2158 = pi129  & n4662;
  assign n2159 = ~pi129  & n821;
  assign n2160 = ~pi129  & n822;
  assign n2161 = ~n2159 & ~n2160;
  assign n2162 = ~pi129  & n4650;
  assign n2163 = pi129  & ~n4662;
  assign n2164 = ~pi129  & ~n4650;
  assign n2165 = ~n2163 & ~n2164;
  assign n2166 = n4858 & n4859;
  assign n2167 = n343 & n4860;
  assign n2168 = ~n2154 & ~n2167;
  assign n2169 = n2141 & n2168;
  assign n2170 = n476 & ~n2169;
  assign n2171 = ~n2114 & ~n2170;
  assign n2172 = n2062 & n2171;
  assign n2173 = pi134  & ~n2172;
  assign n2174 = ~n1949 & ~n2173;
  assign n2175 = ~pi129  & ~n1298;
  assign n2176 = pi129  & ~n1335;
  assign n2177 = pi129  & n1335;
  assign n2178 = ~pi129  & n1298;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = ~n2175 & ~n2176;
  assign n2181 = pi129  & n1345;
  assign n2182 = ~pi129  & n1304;
  assign n2183 = ~pi129  & ~n1304;
  assign n2184 = pi129  & ~n1345;
  assign n2185 = ~n2183 & ~n2184;
  assign n2186 = ~n2181 & ~n2182;
  assign n2187 = n4861 & ~n4862;
  assign n2188 = n264 & ~n2187;
  assign n2189 = ~pi129  & ~n1337;
  assign n2190 = pi129  & ~n1353;
  assign n2191 = pi129  & n1353;
  assign n2192 = ~pi129  & n1337;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = ~n2189 & ~n2190;
  assign n2195 = pi129  & n1363;
  assign n2196 = ~pi129  & n1343;
  assign n2197 = ~pi129  & ~n1343;
  assign n2198 = pi129  & ~n1363;
  assign n2199 = ~n2197 & ~n2198;
  assign n2200 = ~n2195 & ~n2196;
  assign n2201 = n4863 & ~n4864;
  assign n2202 = n290 & ~n2201;
  assign n2203 = ~n2188 & ~n2202;
  assign n2204 = ~pi129  & ~n1392;
  assign n2205 = pi129  & ~n1372;
  assign n2206 = pi129  & n1372;
  assign n2207 = ~pi129  & n1392;
  assign n2208 = ~n2206 & ~n2207;
  assign n2209 = ~n2204 & ~n2205;
  assign n2210 = pi129  & n1382;
  assign n2211 = ~pi129  & n1398;
  assign n2212 = ~pi129  & ~n1398;
  assign n2213 = pi129  & ~n1382;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = ~n2210 & ~n2211;
  assign n2216 = n4865 & ~n4866;
  assign n2217 = n317 & ~n2216;
  assign n2218 = ~pi129  & ~n1355;
  assign n2219 = pi129  & ~n1390;
  assign n2220 = pi129  & n1390;
  assign n2221 = ~pi129  & n1355;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = ~n2218 & ~n2219;
  assign n2224 = pi129  & n1400;
  assign n2225 = ~pi129  & n1361;
  assign n2226 = ~pi129  & ~n1361;
  assign n2227 = pi129  & ~n1400;
  assign n2228 = ~n2226 & ~n2227;
  assign n2229 = ~n2224 & ~n2225;
  assign n2230 = n4867 & ~n4868;
  assign n2231 = n343 & ~n2230;
  assign n2232 = ~n2217 & ~n2231;
  assign n2233 = n2203 & n2232;
  assign n2234 = n687 & ~n2233;
  assign n2235 = ~pi129  & ~n1374;
  assign n2236 = pi129  & ~n1182;
  assign n2237 = pi129  & n1182;
  assign n2238 = ~pi129  & n1374;
  assign n2239 = ~n2237 & ~n2238;
  assign n2240 = ~n2235 & ~n2236;
  assign n2241 = pi129  & n1192;
  assign n2242 = ~pi129  & n1380;
  assign n2243 = ~pi129  & ~n1380;
  assign n2244 = pi129  & ~n1192;
  assign n2245 = ~n2243 & ~n2244;
  assign n2246 = ~n2241 & ~n2242;
  assign n2247 = n4869 & ~n4870;
  assign n2248 = n264 & ~n2247;
  assign n2249 = ~pi129  & ~n1184;
  assign n2250 = pi129  & ~n1200;
  assign n2251 = pi129  & n1200;
  assign n2252 = ~pi129  & n1184;
  assign n2253 = ~n2251 & ~n2252;
  assign n2254 = ~n2249 & ~n2250;
  assign n2255 = pi129  & n1210;
  assign n2256 = ~pi129  & n1190;
  assign n2257 = ~pi129  & ~n1190;
  assign n2258 = pi129  & ~n1210;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = ~n2255 & ~n2256;
  assign n2261 = n4871 & ~n4872;
  assign n2262 = n290 & ~n2261;
  assign n2263 = ~n2248 & ~n2262;
  assign n2264 = ~pi129  & ~n1239;
  assign n2265 = pi129  & ~n1219;
  assign n2266 = pi129  & n1219;
  assign n2267 = ~pi129  & n1239;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = ~n2264 & ~n2265;
  assign n2270 = pi129  & n1229;
  assign n2271 = ~pi129  & n1245;
  assign n2272 = ~pi129  & ~n1245;
  assign n2273 = pi129  & ~n1229;
  assign n2274 = ~n2272 & ~n2273;
  assign n2275 = ~n2270 & ~n2271;
  assign n2276 = n4873 & ~n4874;
  assign n2277 = n317 & ~n2276;
  assign n2278 = ~pi129  & ~n1202;
  assign n2279 = pi129  & ~n1237;
  assign n2280 = pi129  & n1237;
  assign n2281 = ~pi129  & n1202;
  assign n2282 = ~n2280 & ~n2281;
  assign n2283 = ~n2278 & ~n2279;
  assign n2284 = pi129  & n1247;
  assign n2285 = ~pi129  & n1208;
  assign n2286 = ~pi129  & ~n1208;
  assign n2287 = pi129  & ~n1247;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = ~n2284 & ~n2285;
  assign n2290 = n4875 & ~n4876;
  assign n2291 = n343 & ~n2290;
  assign n2292 = ~n2277 & ~n2291;
  assign n2293 = n2263 & n2292;
  assign n2294 = n476 & ~n2293;
  assign n2295 = ~n2234 & ~n2294;
  assign n2296 = ~pi129  & ~n1529;
  assign n2297 = pi129  & ~n1259;
  assign n2298 = pi129  & n1259;
  assign n2299 = ~pi129  & n1529;
  assign n2300 = ~n2298 & ~n2299;
  assign n2301 = ~n2296 & ~n2297;
  assign n2302 = pi129  & n1269;
  assign n2303 = ~pi129  & n1535;
  assign n2304 = ~pi129  & ~n1535;
  assign n2305 = pi129  & ~n1269;
  assign n2306 = ~n2304 & ~n2305;
  assign n2307 = ~n2302 & ~n2303;
  assign n2308 = n4877 & ~n4878;
  assign n2309 = n264 & ~n2308;
  assign n2310 = ~pi129  & ~n1261;
  assign n2311 = pi129  & ~n1277;
  assign n2312 = pi129  & n1277;
  assign n2313 = ~pi129  & n1261;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = ~n2310 & ~n2311;
  assign n2316 = pi129  & n1287;
  assign n2317 = ~pi129  & n1267;
  assign n2318 = ~pi129  & ~n1267;
  assign n2319 = pi129  & ~n1287;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = ~n2316 & ~n2317;
  assign n2322 = n4879 & ~n4880;
  assign n2323 = n290 & ~n2322;
  assign n2324 = ~n2309 & ~n2323;
  assign n2325 = ~pi129  & ~n1316;
  assign n2326 = pi129  & ~n1296;
  assign n2327 = pi129  & n1296;
  assign n2328 = ~pi129  & n1316;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = ~n2325 & ~n2326;
  assign n2331 = pi129  & n1306;
  assign n2332 = ~pi129  & n1322;
  assign n2333 = ~pi129  & ~n1322;
  assign n2334 = pi129  & ~n1306;
  assign n2335 = ~n2333 & ~n2334;
  assign n2336 = ~n2331 & ~n2332;
  assign n2337 = n4881 & ~n4882;
  assign n2338 = n317 & ~n2337;
  assign n2339 = ~pi129  & ~n1279;
  assign n2340 = pi129  & ~n1314;
  assign n2341 = pi129  & n1314;
  assign n2342 = ~pi129  & n1279;
  assign n2343 = ~n2341 & ~n2342;
  assign n2344 = ~n2339 & ~n2340;
  assign n2345 = pi129  & n1324;
  assign n2346 = ~pi129  & n1285;
  assign n2347 = ~pi129  & ~n1285;
  assign n2348 = pi129  & ~n1324;
  assign n2349 = ~n2347 & ~n2348;
  assign n2350 = ~n2345 & ~n2346;
  assign n2351 = n4883 & ~n4884;
  assign n2352 = n343 & ~n2351;
  assign n2353 = ~n2338 & ~n2352;
  assign n2354 = n2324 & n2353;
  assign n2355 = n582 & ~n2354;
  assign n2356 = ~pi129  & ~n1221;
  assign n2357 = pi129  & ~n1106;
  assign n2358 = pi129  & n1106;
  assign n2359 = ~pi129  & n1221;
  assign n2360 = ~n2358 & ~n2359;
  assign n2361 = ~n2356 & ~n2357;
  assign n2362 = pi129  & n1116;
  assign n2363 = ~pi129  & n1227;
  assign n2364 = ~pi129  & ~n1227;
  assign n2365 = pi129  & ~n1116;
  assign n2366 = ~n2364 & ~n2365;
  assign n2367 = ~n2362 & ~n2363;
  assign n2368 = n4885 & ~n4886;
  assign n2369 = n264 & ~n2368;
  assign n2370 = ~pi129  & ~n1108;
  assign n2371 = pi129  & ~n1124;
  assign n2372 = pi129  & n1124;
  assign n2373 = ~pi129  & n1108;
  assign n2374 = ~n2372 & ~n2373;
  assign n2375 = ~n2370 & ~n2371;
  assign n2376 = pi129  & n1134;
  assign n2377 = ~pi129  & n1114;
  assign n2378 = ~pi129  & ~n1114;
  assign n2379 = pi129  & ~n1134;
  assign n2380 = ~n2378 & ~n2379;
  assign n2381 = ~n2376 & ~n2377;
  assign n2382 = n4887 & ~n4888;
  assign n2383 = n290 & ~n2382;
  assign n2384 = ~n2369 & ~n2383;
  assign n2385 = ~pi129  & ~n1163;
  assign n2386 = pi129  & ~n1143;
  assign n2387 = pi129  & n1143;
  assign n2388 = ~pi129  & n1163;
  assign n2389 = ~n2387 & ~n2388;
  assign n2390 = ~n2385 & ~n2386;
  assign n2391 = pi129  & n1153;
  assign n2392 = ~pi129  & n1169;
  assign n2393 = ~pi129  & ~n1169;
  assign n2394 = pi129  & ~n1153;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = ~n2391 & ~n2392;
  assign n2397 = n4889 & ~n4890;
  assign n2398 = n317 & ~n2397;
  assign n2399 = ~pi129  & ~n1126;
  assign n2400 = pi129  & ~n1161;
  assign n2401 = pi129  & n1161;
  assign n2402 = ~pi129  & n1126;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = ~n2399 & ~n2400;
  assign n2405 = pi129  & n1171;
  assign n2406 = ~pi129  & n1132;
  assign n2407 = ~pi129  & ~n1132;
  assign n2408 = pi129  & ~n1171;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410 = ~n2405 & ~n2406;
  assign n2411 = n4891 & ~n4892;
  assign n2412 = n343 & ~n2411;
  assign n2413 = ~n2398 & ~n2412;
  assign n2414 = n2384 & n2413;
  assign n2415 = n371 & ~n2414;
  assign n2416 = ~n2355 & ~n2415;
  assign n2417 = n2295 & n2416;
  assign n2418 = ~pi134  & ~n2417;
  assign n2419 = ~pi129  & ~n1145;
  assign n2420 = pi129  & ~n1414;
  assign n2421 = pi129  & n1414;
  assign n2422 = ~pi129  & n1145;
  assign n2423 = ~n2421 & ~n2422;
  assign n2424 = ~n2419 & ~n2420;
  assign n2425 = pi129  & n1424;
  assign n2426 = ~pi129  & n1151;
  assign n2427 = ~pi129  & ~n1151;
  assign n2428 = pi129  & ~n1424;
  assign n2429 = ~n2427 & ~n2428;
  assign n2430 = ~n2425 & ~n2426;
  assign n2431 = n4893 & ~n4894;
  assign n2432 = n264 & ~n2431;
  assign n2433 = ~pi129  & ~n1416;
  assign n2434 = pi129  & ~n1432;
  assign n2435 = pi129  & n1432;
  assign n2436 = ~pi129  & n1416;
  assign n2437 = ~n2435 & ~n2436;
  assign n2438 = ~n2433 & ~n2434;
  assign n2439 = pi129  & n1442;
  assign n2440 = ~pi129  & n1422;
  assign n2441 = ~pi129  & ~n1422;
  assign n2442 = pi129  & ~n1442;
  assign n2443 = ~n2441 & ~n2442;
  assign n2444 = ~n2439 & ~n2440;
  assign n2445 = n4895 & ~n4896;
  assign n2446 = n290 & ~n2445;
  assign n2447 = ~n2432 & ~n2446;
  assign n2448 = ~pi129  & ~n1471;
  assign n2449 = pi129  & ~n1451;
  assign n2450 = pi129  & n1451;
  assign n2451 = ~pi129  & n1471;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = ~n2448 & ~n2449;
  assign n2454 = pi129  & n1461;
  assign n2455 = ~pi129  & n1477;
  assign n2456 = ~pi129  & ~n1477;
  assign n2457 = pi129  & ~n1461;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = ~n2454 & ~n2455;
  assign n2460 = n4897 & ~n4898;
  assign n2461 = n317 & ~n2460;
  assign n2462 = ~pi129  & ~n1434;
  assign n2463 = pi129  & ~n1469;
  assign n2464 = pi129  & n1469;
  assign n2465 = ~pi129  & n1434;
  assign n2466 = ~n2464 & ~n2465;
  assign n2467 = ~n2462 & ~n2463;
  assign n2468 = pi129  & n1479;
  assign n2469 = ~pi129  & n1440;
  assign n2470 = ~pi129  & ~n1440;
  assign n2471 = pi129  & ~n1479;
  assign n2472 = ~n2470 & ~n2471;
  assign n2473 = ~n2468 & ~n2469;
  assign n2474 = n4899 & ~n4900;
  assign n2475 = n343 & ~n2474;
  assign n2476 = ~n2461 & ~n2475;
  assign n2477 = n2447 & n2476;
  assign n2478 = n582 & ~n2477;
  assign n2479 = ~pi129  & ~n1453;
  assign n2480 = pi129  & ~n1567;
  assign n2481 = pi129  & n1567;
  assign n2482 = ~pi129  & n1453;
  assign n2483 = ~n2481 & ~n2482;
  assign n2484 = ~n2479 & ~n2480;
  assign n2485 = pi129  & n1577;
  assign n2486 = ~pi129  & n1459;
  assign n2487 = ~pi129  & ~n1459;
  assign n2488 = pi129  & ~n1577;
  assign n2489 = ~n2487 & ~n2488;
  assign n2490 = ~n2485 & ~n2486;
  assign n2491 = n4901 & ~n4902;
  assign n2492 = n264 & ~n2491;
  assign n2493 = pi129  & n1593;
  assign n2494 = pi129  & n1592;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = pi129  & n4753;
  assign n2497 = ~n1569 & ~n1575;
  assign n2498 = ~pi129  & n1575;
  assign n2499 = ~pi129  & n1569;
  assign n2500 = ~n2498 & ~n2499;
  assign n2501 = ~pi129  & ~n2497;
  assign n2502 = n4903 & n4904;
  assign n2503 = n290 & ~n2502;
  assign n2504 = ~n2492 & ~n2503;
  assign n2505 = ~pi129  & ~n1631;
  assign n2506 = pi129  & ~n1605;
  assign n2507 = pi129  & n1605;
  assign n2508 = ~pi129  & n1631;
  assign n2509 = ~n2507 & ~n2508;
  assign n2510 = ~n2505 & ~n2506;
  assign n2511 = pi129  & n1615;
  assign n2512 = ~pi129  & n1630;
  assign n2513 = ~pi129  & ~n1630;
  assign n2514 = pi129  & ~n1615;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = ~n2511 & ~n2512;
  assign n2517 = n4905 & ~n4906;
  assign n2518 = n317 & ~n2517;
  assign n2519 = ~pi129  & ~n1585;
  assign n2520 = pi129  & ~n1623;
  assign n2521 = pi129  & n1623;
  assign n2522 = ~pi129  & n1585;
  assign n2523 = ~n2521 & ~n2522;
  assign n2524 = ~n2519 & ~n2520;
  assign n2525 = pi129  & n1624;
  assign n2526 = ~pi129  & n1586;
  assign n2527 = ~pi129  & ~n1586;
  assign n2528 = pi129  & ~n1624;
  assign n2529 = ~n2527 & ~n2528;
  assign n2530 = ~n2525 & ~n2526;
  assign n2531 = n4907 & ~n4908;
  assign n2532 = n343 & ~n2531;
  assign n2533 = ~n2518 & ~n2532;
  assign n2534 = n2504 & n2533;
  assign n2535 = n687 & ~n2534;
  assign n2536 = ~n2478 & ~n2535;
  assign n2537 = ~pi129  & ~n1681;
  assign n2538 = pi129  & ~n1490;
  assign n2539 = pi129  & n1490;
  assign n2540 = ~pi129  & n1681;
  assign n2541 = ~n2539 & ~n2540;
  assign n2542 = ~n2537 & ~n2538;
  assign n2543 = pi129  & n1500;
  assign n2544 = ~pi129  & n1687;
  assign n2545 = ~pi129  & ~n1687;
  assign n2546 = pi129  & ~n1500;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = ~n2543 & ~n2544;
  assign n2549 = n4909 & ~n4910;
  assign n2550 = n264 & ~n2549;
  assign n2551 = ~pi129  & ~n1492;
  assign n2552 = pi129  & ~n1508;
  assign n2553 = pi129  & n1508;
  assign n2554 = ~pi129  & n1492;
  assign n2555 = ~n2553 & ~n2554;
  assign n2556 = ~n2551 & ~n2552;
  assign n2557 = pi129  & n1518;
  assign n2558 = ~pi129  & n1498;
  assign n2559 = ~pi129  & ~n1498;
  assign n2560 = pi129  & ~n1518;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = ~n2557 & ~n2558;
  assign n2563 = n4911 & ~n4912;
  assign n2564 = n290 & ~n2563;
  assign n2565 = ~n2550 & ~n2564;
  assign n2566 = ~pi129  & ~n1547;
  assign n2567 = pi129  & ~n1527;
  assign n2568 = pi129  & n1527;
  assign n2569 = ~pi129  & n1547;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = ~n2566 & ~n2567;
  assign n2572 = pi129  & n1537;
  assign n2573 = ~pi129  & n1553;
  assign n2574 = ~pi129  & ~n1553;
  assign n2575 = pi129  & ~n1537;
  assign n2576 = ~n2574 & ~n2575;
  assign n2577 = ~n2572 & ~n2573;
  assign n2578 = n4913 & ~n4914;
  assign n2579 = n317 & ~n2578;
  assign n2580 = ~pi129  & ~n1510;
  assign n2581 = pi129  & ~n1545;
  assign n2582 = pi129  & n1545;
  assign n2583 = ~pi129  & n1510;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = ~n2580 & ~n2581;
  assign n2586 = pi129  & n1555;
  assign n2587 = ~pi129  & n1516;
  assign n2588 = ~pi129  & ~n1516;
  assign n2589 = pi129  & ~n1555;
  assign n2590 = ~n2588 & ~n2589;
  assign n2591 = ~n2586 & ~n2587;
  assign n2592 = n4915 & ~n4916;
  assign n2593 = n343 & ~n2592;
  assign n2594 = ~n2579 & ~n2593;
  assign n2595 = n2565 & n2594;
  assign n2596 = n371 & ~n2595;
  assign n2597 = ~pi129  & ~n1607;
  assign n2598 = pi129  & ~n1642;
  assign n2599 = pi129  & n1642;
  assign n2600 = ~pi129  & n1607;
  assign n2601 = ~n2599 & ~n2600;
  assign n2602 = ~n2597 & ~n2598;
  assign n2603 = pi129  & n1652;
  assign n2604 = ~pi129  & n1613;
  assign n2605 = ~pi129  & ~n1613;
  assign n2606 = pi129  & ~n1652;
  assign n2607 = ~n2605 & ~n2606;
  assign n2608 = ~n2603 & ~n2604;
  assign n2609 = n4917 & ~n4918;
  assign n2610 = n264 & ~n2609;
  assign n2611 = ~pi129  & ~n1644;
  assign n2612 = pi129  & ~n1660;
  assign n2613 = pi129  & n1660;
  assign n2614 = ~pi129  & n1644;
  assign n2615 = ~n2613 & ~n2614;
  assign n2616 = ~n2611 & ~n2612;
  assign n2617 = pi129  & n1670;
  assign n2618 = ~pi129  & n1650;
  assign n2619 = ~pi129  & ~n1650;
  assign n2620 = pi129  & ~n1670;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = ~n2617 & ~n2618;
  assign n2623 = n4919 & ~n4920;
  assign n2624 = n290 & ~n2623;
  assign n2625 = ~n2610 & ~n2624;
  assign n2626 = ~pi129  & ~n1699;
  assign n2627 = pi129  & ~n1679;
  assign n2628 = pi129  & n1679;
  assign n2629 = ~pi129  & n1699;
  assign n2630 = ~n2628 & ~n2629;
  assign n2631 = ~n2626 & ~n2627;
  assign n2632 = pi129  & n1689;
  assign n2633 = ~pi129  & n1705;
  assign n2634 = ~pi129  & ~n1705;
  assign n2635 = pi129  & ~n1689;
  assign n2636 = ~n2634 & ~n2635;
  assign n2637 = ~n2632 & ~n2633;
  assign n2638 = n4921 & ~n4922;
  assign n2639 = n317 & ~n2638;
  assign n2640 = ~pi129  & ~n1662;
  assign n2641 = pi129  & ~n1697;
  assign n2642 = pi129  & n1697;
  assign n2643 = ~pi129  & n1662;
  assign n2644 = ~n2642 & ~n2643;
  assign n2645 = ~n2640 & ~n2641;
  assign n2646 = pi129  & n1707;
  assign n2647 = ~pi129  & n1668;
  assign n2648 = ~pi129  & ~n1668;
  assign n2649 = pi129  & ~n1707;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = ~n2646 & ~n2647;
  assign n2652 = n4923 & ~n4924;
  assign n2653 = n343 & ~n2652;
  assign n2654 = ~n2639 & ~n2653;
  assign n2655 = n2625 & n2654;
  assign n2656 = n476 & ~n2655;
  assign n2657 = ~n2596 & ~n2656;
  assign n2658 = n2536 & n2657;
  assign n2659 = pi134  & ~n2658;
  assign n2660 = ~n2418 & ~n2659;
  assign n2661 = n264 & n4579;
  assign n2662 = n4549 & n290;
  assign n2663 = ~n2661 & ~n2662;
  assign n2664 = n317 & n4564;
  assign n2665 = n4554 & n343;
  assign n2666 = ~n2664 & ~n2665;
  assign n2667 = n2663 & n2666;
  assign n2668 = n371 & ~n2667;
  assign n2669 = n264 & n4619;
  assign n2670 = n290 & n4569;
  assign n2671 = ~n2669 & ~n2670;
  assign n2672 = n317 & n4584;
  assign n2673 = n343 & n4574;
  assign n2674 = ~n2672 & ~n2673;
  assign n2675 = n2671 & n2674;
  assign n2676 = n476 & ~n2675;
  assign n2677 = ~n2668 & ~n2676;
  assign n2678 = n264 & n4639;
  assign n2679 = n290 & n4589;
  assign n2680 = ~n2678 & ~n2679;
  assign n2681 = n317 & n4604;
  assign n2682 = n343 & n4594;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = n2680 & n2683;
  assign n2685 = n582 & ~n2684;
  assign n2686 = n264 & n4599;
  assign n2687 = n290 & n4609;
  assign n2688 = ~n2686 & ~n2687;
  assign n2689 = n317 & n4624;
  assign n2690 = n343 & n4614;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = n2688 & n2691;
  assign n2693 = n687 & ~n2692;
  assign n2694 = ~n2685 & ~n2693;
  assign n2695 = n2677 & n2694;
  assign n2696 = ~pi134  & ~n2695;
  assign n2697 = n264 & n4679;
  assign n2698 = n290 & n4689;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = n317 & ~n1097;
  assign n2701 = n343 & n4694;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = n2699 & n2702;
  assign n2704 = n687 & ~n2703;
  assign n2705 = n264 & n4559;
  assign n2706 = n290 & n4669;
  assign n2707 = ~n2705 & ~n2706;
  assign n2708 = n317 & n4684;
  assign n2709 = n343 & n4674;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = n2707 & n2710;
  assign n2712 = n582 & ~n2711;
  assign n2713 = ~n2704 & ~n2712;
  assign n2714 = n264 & n4699;
  assign n2715 = n290 & n4649;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = n317 & n4664;
  assign n2718 = n343 & n4654;
  assign n2719 = ~n2717 & ~n2718;
  assign n2720 = n2716 & n2719;
  assign n2721 = n476 & ~n2720;
  assign n2722 = n264 & n4659;
  assign n2723 = n290 & n4629;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = n317 & n4644;
  assign n2726 = n343 & n4634;
  assign n2727 = ~n2725 & ~n2726;
  assign n2728 = n2724 & n2727;
  assign n2729 = n371 & ~n2728;
  assign n2730 = ~n2721 & ~n2729;
  assign n2731 = n2713 & n2730;
  assign n2732 = pi134  & ~n2731;
  assign n2733 = ~n2696 & ~n2732;
  assign n2734 = n264 & ~n1235;
  assign n2735 = n290 & ~n1122;
  assign n2736 = ~n2734 & ~n2735;
  assign n2737 = n317 & ~n1177;
  assign n2738 = n343 & ~n1140;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = n2736 & n2739;
  assign n2741 = n371 & ~n2740;
  assign n2742 = n264 & ~n1388;
  assign n2743 = n290 & ~n1198;
  assign n2744 = ~n2742 & ~n2743;
  assign n2745 = n317 & ~n1253;
  assign n2746 = n343 & ~n1216;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = n2744 & n2747;
  assign n2749 = n476 & ~n2748;
  assign n2750 = ~n2741 & ~n2749;
  assign n2751 = n264 & ~n1543;
  assign n2752 = n290 & ~n1275;
  assign n2753 = ~n2751 & ~n2752;
  assign n2754 = n317 & ~n1330;
  assign n2755 = n343 & ~n1293;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = n2753 & n2756;
  assign n2758 = n582 & ~n2757;
  assign n2759 = n264 & ~n1312;
  assign n2760 = n290 & ~n1351;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = n317 & ~n1406;
  assign n2763 = n343 & ~n1369;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = n2761 & n2764;
  assign n2766 = n687 & ~n2765;
  assign n2767 = ~n2758 & ~n2766;
  assign n2768 = n2750 & n2767;
  assign n2769 = ~pi134  & ~n2768;
  assign n2770 = n264 & ~n1467;
  assign n2771 = n290 & ~n1583;
  assign n2772 = ~n2770 & ~n2771;
  assign n2773 = n317 & ~n1637;
  assign n2774 = n343 & ~n1602;
  assign n2775 = ~n2773 & ~n2774;
  assign n2776 = n2772 & n2775;
  assign n2777 = n687 & ~n2776;
  assign n2778 = n264 & ~n1159;
  assign n2779 = n290 & ~n1430;
  assign n2780 = ~n2778 & ~n2779;
  assign n2781 = n317 & ~n1485;
  assign n2782 = n343 & ~n1448;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = n2780 & n2783;
  assign n2785 = n582 & ~n2784;
  assign n2786 = ~n2777 & ~n2785;
  assign n2787 = n264 & ~n1621;
  assign n2788 = n290 & ~n1658;
  assign n2789 = ~n2787 & ~n2788;
  assign n2790 = n317 & ~n1713;
  assign n2791 = n343 & ~n1676;
  assign n2792 = ~n2790 & ~n2791;
  assign n2793 = n2789 & n2792;
  assign n2794 = n476 & ~n2793;
  assign n2795 = n264 & ~n1695;
  assign n2796 = n290 & ~n1506;
  assign n2797 = ~n2795 & ~n2796;
  assign n2798 = n317 & ~n1561;
  assign n2799 = n343 & ~n1524;
  assign n2800 = ~n2798 & ~n2799;
  assign n2801 = n2797 & n2800;
  assign n2802 = n371 & ~n2801;
  assign n2803 = ~n2794 & ~n2802;
  assign n2804 = n2786 & n2803;
  assign n2805 = pi134  & ~n2804;
  assign n2806 = ~n2769 & ~n2805;
  assign n2807 = n264 & n4787;
  assign n2808 = n290 & n4769;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = n317 & n4778;
  assign n2811 = n343 & n4772;
  assign n2812 = ~n2810 & ~n2811;
  assign n2813 = n2809 & n2812;
  assign n2814 = n371 & ~n2813;
  assign n2815 = n264 & n4811;
  assign n2816 = n290 & n4781;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = n317 & n4790;
  assign n2819 = n343 & n4784;
  assign n2820 = ~n2818 & ~n2819;
  assign n2821 = n2817 & n2820;
  assign n2822 = n476 & ~n2821;
  assign n2823 = ~n2814 & ~n2822;
  assign n2824 = n264 & n4835;
  assign n2825 = n290 & n4793;
  assign n2826 = ~n2824 & ~n2825;
  assign n2827 = n317 & n4802;
  assign n2828 = n343 & n4796;
  assign n2829 = ~n2827 & ~n2828;
  assign n2830 = n2826 & n2829;
  assign n2831 = n582 & ~n2830;
  assign n2832 = n264 & n4799;
  assign n2833 = n290 & n4805;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = n317 & n4814;
  assign n2836 = n343 & n4808;
  assign n2837 = ~n2835 & ~n2836;
  assign n2838 = n2834 & n2837;
  assign n2839 = n687 & ~n2838;
  assign n2840 = ~n2831 & ~n2839;
  assign n2841 = n2823 & n2840;
  assign n2842 = ~pi134  & ~n2841;
  assign n2843 = n264 & n4823;
  assign n2844 = n290 & n4841;
  assign n2845 = ~n2843 & ~n2844;
  assign n2846 = n317 & ~n2110;
  assign n2847 = n343 & n4844;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = n2845 & n2848;
  assign n2850 = n687 & ~n2849;
  assign n2851 = n264 & n4775;
  assign n2852 = n290 & n4817;
  assign n2853 = ~n2851 & ~n2852;
  assign n2854 = n317 & n4826;
  assign n2855 = n343 & n4820;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857 = n2853 & n2856;
  assign n2858 = n582 & ~n2857;
  assign n2859 = ~n2850 & ~n2858;
  assign n2860 = n264 & ~n2099;
  assign n2861 = n290 & n4851;
  assign n2862 = ~n2860 & ~n2861;
  assign n2863 = n317 & n4860;
  assign n2864 = n343 & n4854;
  assign n2865 = ~n2863 & ~n2864;
  assign n2866 = n2862 & n2865;
  assign n2867 = n476 & ~n2866;
  assign n2868 = n264 & n4857;
  assign n2869 = n290 & n4829;
  assign n2870 = ~n2868 & ~n2869;
  assign n2871 = n317 & n4838;
  assign n2872 = n343 & n4832;
  assign n2873 = ~n2871 & ~n2872;
  assign n2874 = n2870 & n2873;
  assign n2875 = n371 & ~n2874;
  assign n2876 = ~n2867 & ~n2875;
  assign n2877 = n2859 & n2876;
  assign n2878 = pi134  & ~n2877;
  assign n2879 = ~n2842 & ~n2878;
  assign n2880 = n264 & ~n2276;
  assign n2881 = n290 & ~n2368;
  assign n2882 = ~n2880 & ~n2881;
  assign n2883 = n317 & ~n2411;
  assign n2884 = n343 & ~n2382;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = n2882 & n2885;
  assign n2887 = n371 & ~n2886;
  assign n2888 = n264 & ~n2216;
  assign n2889 = n290 & ~n2247;
  assign n2890 = ~n2888 & ~n2889;
  assign n2891 = n317 & ~n2290;
  assign n2892 = n343 & ~n2261;
  assign n2893 = ~n2891 & ~n2892;
  assign n2894 = n2890 & n2893;
  assign n2895 = n476 & ~n2894;
  assign n2896 = ~n2887 & ~n2895;
  assign n2897 = n264 & ~n2578;
  assign n2898 = n290 & ~n2308;
  assign n2899 = ~n2897 & ~n2898;
  assign n2900 = n317 & ~n2351;
  assign n2901 = n343 & ~n2322;
  assign n2902 = ~n2900 & ~n2901;
  assign n2903 = n2899 & n2902;
  assign n2904 = n582 & ~n2903;
  assign n2905 = n264 & ~n2337;
  assign n2906 = n290 & ~n2187;
  assign n2907 = ~n2905 & ~n2906;
  assign n2908 = n317 & ~n2230;
  assign n2909 = n343 & ~n2201;
  assign n2910 = ~n2908 & ~n2909;
  assign n2911 = n2907 & n2910;
  assign n2912 = n687 & ~n2911;
  assign n2913 = ~n2904 & ~n2912;
  assign n2914 = n2896 & n2913;
  assign n2915 = ~pi134  & ~n2914;
  assign n2916 = n290 & ~n2491;
  assign n2917 = n343 & ~n2502;
  assign n2918 = ~n2916 & ~n2917;
  assign n2919 = n317 & ~n2531;
  assign n2920 = n264 & ~n2460;
  assign n2921 = ~n2919 & ~n2920;
  assign n2922 = n2918 & n2921;
  assign n2923 = n687 & ~n2922;
  assign n2924 = n264 & ~n2397;
  assign n2925 = n290 & ~n2431;
  assign n2926 = ~n2924 & ~n2925;
  assign n2927 = n317 & ~n2474;
  assign n2928 = n343 & ~n2445;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = n2926 & n2929;
  assign n2931 = n582 & ~n2930;
  assign n2932 = ~n2923 & ~n2931;
  assign n2933 = n264 & ~n2517;
  assign n2934 = n290 & ~n2609;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = n317 & ~n2652;
  assign n2937 = n343 & ~n2623;
  assign n2938 = ~n2936 & ~n2937;
  assign n2939 = n2935 & n2938;
  assign n2940 = n476 & ~n2939;
  assign n2941 = n264 & ~n2638;
  assign n2942 = n290 & ~n2549;
  assign n2943 = ~n2941 & ~n2942;
  assign n2944 = n317 & ~n2592;
  assign n2945 = n343 & ~n2563;
  assign n2946 = ~n2944 & ~n2945;
  assign n2947 = n2943 & n2946;
  assign n2948 = n371 & ~n2947;
  assign n2949 = ~n2940 & ~n2948;
  assign n2950 = n2932 & n2949;
  assign n2951 = pi134  & ~n2950;
  assign n2952 = ~n2915 & ~n2951;
  assign n2953 = n264 & n4584;
  assign n2954 = n290 & n4579;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = n4554 & n317;
  assign n2957 = n4549 & n343;
  assign n2958 = ~n2956 & ~n2957;
  assign n2959 = n2955 & n2958;
  assign n2960 = n371 & ~n2959;
  assign n2961 = n264 & n4624;
  assign n2962 = n290 & n4619;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = n317 & n4574;
  assign n2965 = n343 & n4569;
  assign n2966 = ~n2964 & ~n2965;
  assign n2967 = n2963 & n2966;
  assign n2968 = n476 & ~n2967;
  assign n2969 = ~n2960 & ~n2968;
  assign n2970 = n264 & n4644;
  assign n2971 = n290 & n4639;
  assign n2972 = ~n2970 & ~n2971;
  assign n2973 = n317 & n4594;
  assign n2974 = n343 & n4589;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = n2972 & n2975;
  assign n2977 = n582 & ~n2976;
  assign n2978 = n264 & n4604;
  assign n2979 = n290 & n4599;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = n317 & n4614;
  assign n2982 = n343 & n4609;
  assign n2983 = ~n2981 & ~n2982;
  assign n2984 = n2980 & n2983;
  assign n2985 = n687 & ~n2984;
  assign n2986 = ~n2977 & ~n2985;
  assign n2987 = n2969 & n2986;
  assign n2988 = ~pi134  & ~n2987;
  assign n2989 = n264 & n4684;
  assign n2990 = n290 & n4679;
  assign n2991 = ~n2989 & ~n2990;
  assign n2992 = n317 & n4694;
  assign n2993 = n343 & n4689;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = n2991 & n2994;
  assign n2996 = n687 & ~n2995;
  assign n2997 = n264 & n4564;
  assign n2998 = n290 & n4559;
  assign n2999 = ~n2997 & ~n2998;
  assign n3000 = n317 & n4674;
  assign n3001 = n343 & n4669;
  assign n3002 = ~n3000 & ~n3001;
  assign n3003 = n2999 & n3002;
  assign n3004 = n582 & ~n3003;
  assign n3005 = ~n2996 & ~n3004;
  assign n3006 = n264 & ~n1097;
  assign n3007 = n290 & n4699;
  assign n3008 = ~n3006 & ~n3007;
  assign n3009 = n317 & n4654;
  assign n3010 = n343 & n4649;
  assign n3011 = ~n3009 & ~n3010;
  assign n3012 = n3008 & n3011;
  assign n3013 = n476 & ~n3012;
  assign n3014 = n264 & n4664;
  assign n3015 = n290 & n4659;
  assign n3016 = ~n3014 & ~n3015;
  assign n3017 = n317 & n4634;
  assign n3018 = n343 & n4629;
  assign n3019 = ~n3017 & ~n3018;
  assign n3020 = n3016 & n3019;
  assign n3021 = n371 & ~n3020;
  assign n3022 = ~n3013 & ~n3021;
  assign n3023 = n3005 & n3022;
  assign n3024 = pi134  & ~n3023;
  assign n3025 = ~n2988 & ~n3024;
  assign n3026 = n264 & ~n1253;
  assign n3027 = n290 & ~n1235;
  assign n3028 = ~n3026 & ~n3027;
  assign n3029 = n317 & ~n1140;
  assign n3030 = n343 & ~n1122;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = n3028 & n3031;
  assign n3033 = n371 & ~n3032;
  assign n3034 = n264 & ~n1406;
  assign n3035 = n290 & ~n1388;
  assign n3036 = ~n3034 & ~n3035;
  assign n3037 = n317 & ~n1216;
  assign n3038 = n343 & ~n1198;
  assign n3039 = ~n3037 & ~n3038;
  assign n3040 = n3036 & n3039;
  assign n3041 = n476 & ~n3040;
  assign n3042 = ~n3033 & ~n3041;
  assign n3043 = n264 & ~n1561;
  assign n3044 = n290 & ~n1543;
  assign n3045 = ~n3043 & ~n3044;
  assign n3046 = n317 & ~n1293;
  assign n3047 = n343 & ~n1275;
  assign n3048 = ~n3046 & ~n3047;
  assign n3049 = n3045 & n3048;
  assign n3050 = n582 & ~n3049;
  assign n3051 = n264 & ~n1330;
  assign n3052 = n290 & ~n1312;
  assign n3053 = ~n3051 & ~n3052;
  assign n3054 = n317 & ~n1369;
  assign n3055 = n343 & ~n1351;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = n3053 & n3056;
  assign n3058 = n687 & ~n3057;
  assign n3059 = ~n3050 & ~n3058;
  assign n3060 = n3042 & n3059;
  assign n3061 = ~pi134  & ~n3060;
  assign n3062 = n264 & ~n1485;
  assign n3063 = n290 & ~n1467;
  assign n3064 = ~n3062 & ~n3063;
  assign n3065 = n317 & ~n1602;
  assign n3066 = n343 & ~n1583;
  assign n3067 = ~n3065 & ~n3066;
  assign n3068 = n3064 & n3067;
  assign n3069 = n687 & ~n3068;
  assign n3070 = n264 & ~n1177;
  assign n3071 = n290 & ~n1159;
  assign n3072 = ~n3070 & ~n3071;
  assign n3073 = n317 & ~n1448;
  assign n3074 = n343 & ~n1430;
  assign n3075 = ~n3073 & ~n3074;
  assign n3076 = n3072 & n3075;
  assign n3077 = n582 & ~n3076;
  assign n3078 = ~n3069 & ~n3077;
  assign n3079 = n264 & ~n1637;
  assign n3080 = n290 & ~n1621;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = n317 & ~n1676;
  assign n3083 = n343 & ~n1658;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = n3081 & n3084;
  assign n3086 = n476 & ~n3085;
  assign n3087 = n264 & ~n1713;
  assign n3088 = n290 & ~n1695;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090 = n317 & ~n1524;
  assign n3091 = n343 & ~n1506;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = n3089 & n3092;
  assign n3094 = n371 & ~n3093;
  assign n3095 = ~n3086 & ~n3094;
  assign n3096 = n3078 & n3095;
  assign n3097 = pi134  & ~n3096;
  assign n3098 = ~n3061 & ~n3097;
  assign n3099 = n264 & n4790;
  assign n3100 = n290 & n4787;
  assign n3101 = ~n3099 & ~n3100;
  assign n3102 = n317 & n4772;
  assign n3103 = n343 & n4769;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = n3101 & n3104;
  assign n3106 = n371 & ~n3105;
  assign n3107 = n264 & n4814;
  assign n3108 = n290 & n4811;
  assign n3109 = ~n3107 & ~n3108;
  assign n3110 = n317 & n4784;
  assign n3111 = n343 & n4781;
  assign n3112 = ~n3110 & ~n3111;
  assign n3113 = n3109 & n3112;
  assign n3114 = n476 & ~n3113;
  assign n3115 = ~n3106 & ~n3114;
  assign n3116 = n264 & n4838;
  assign n3117 = n290 & n4835;
  assign n3118 = ~n3116 & ~n3117;
  assign n3119 = n317 & n4796;
  assign n3120 = n343 & n4793;
  assign n3121 = ~n3119 & ~n3120;
  assign n3122 = n3118 & n3121;
  assign n3123 = n582 & ~n3122;
  assign n3124 = n264 & n4802;
  assign n3125 = n290 & n4799;
  assign n3126 = ~n3124 & ~n3125;
  assign n3127 = n317 & n4808;
  assign n3128 = n343 & n4805;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130 = n3126 & n3129;
  assign n3131 = n687 & ~n3130;
  assign n3132 = ~n3123 & ~n3131;
  assign n3133 = n3115 & n3132;
  assign n3134 = ~pi134  & ~n3133;
  assign n3135 = n264 & n4826;
  assign n3136 = n290 & n4823;
  assign n3137 = ~n3135 & ~n3136;
  assign n3138 = n317 & n4844;
  assign n3139 = n343 & n4841;
  assign n3140 = ~n3138 & ~n3139;
  assign n3141 = n3137 & n3140;
  assign n3142 = n687 & ~n3141;
  assign n3143 = n264 & n4778;
  assign n3144 = n290 & n4775;
  assign n3145 = ~n3143 & ~n3144;
  assign n3146 = n317 & n4820;
  assign n3147 = n343 & n4817;
  assign n3148 = ~n3146 & ~n3147;
  assign n3149 = n3145 & n3148;
  assign n3150 = n582 & ~n3149;
  assign n3151 = ~n3142 & ~n3150;
  assign n3152 = n264 & ~n2110;
  assign n3153 = n290 & ~n2099;
  assign n3154 = ~n3152 & ~n3153;
  assign n3155 = n317 & n4854;
  assign n3156 = n343 & n4851;
  assign n3157 = ~n3155 & ~n3156;
  assign n3158 = n3154 & n3157;
  assign n3159 = n476 & ~n3158;
  assign n3160 = n264 & n4860;
  assign n3161 = n290 & n4857;
  assign n3162 = ~n3160 & ~n3161;
  assign n3163 = n317 & n4832;
  assign n3164 = n343 & n4829;
  assign n3165 = ~n3163 & ~n3164;
  assign n3166 = n3162 & n3165;
  assign n3167 = n371 & ~n3166;
  assign n3168 = ~n3159 & ~n3167;
  assign n3169 = n3151 & n3168;
  assign n3170 = pi134  & ~n3169;
  assign n3171 = ~n3134 & ~n3170;
  assign n3172 = n264 & ~n2290;
  assign n3173 = n290 & ~n2276;
  assign n3174 = ~n3172 & ~n3173;
  assign n3175 = n317 & ~n2382;
  assign n3176 = n343 & ~n2368;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = n3174 & n3177;
  assign n3179 = n371 & ~n3178;
  assign n3180 = n264 & ~n2230;
  assign n3181 = n290 & ~n2216;
  assign n3182 = ~n3180 & ~n3181;
  assign n3183 = n317 & ~n2261;
  assign n3184 = n343 & ~n2247;
  assign n3185 = ~n3183 & ~n3184;
  assign n3186 = n3182 & n3185;
  assign n3187 = n476 & ~n3186;
  assign n3188 = ~n3179 & ~n3187;
  assign n3189 = n264 & ~n2592;
  assign n3190 = n290 & ~n2578;
  assign n3191 = ~n3189 & ~n3190;
  assign n3192 = n317 & ~n2322;
  assign n3193 = n343 & ~n2308;
  assign n3194 = ~n3192 & ~n3193;
  assign n3195 = n3191 & n3194;
  assign n3196 = n582 & ~n3195;
  assign n3197 = n264 & ~n2351;
  assign n3198 = n290 & ~n2337;
  assign n3199 = ~n3197 & ~n3198;
  assign n3200 = n317 & ~n2201;
  assign n3201 = n343 & ~n2187;
  assign n3202 = ~n3200 & ~n3201;
  assign n3203 = n3199 & n3202;
  assign n3204 = n687 & ~n3203;
  assign n3205 = ~n3196 & ~n3204;
  assign n3206 = n3188 & n3205;
  assign n3207 = ~pi134  & ~n3206;
  assign n3208 = n264 & ~n2474;
  assign n3209 = n343 & ~n2491;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = n317 & ~n2502;
  assign n3212 = n290 & ~n2460;
  assign n3213 = ~n3211 & ~n3212;
  assign n3214 = n3210 & n3213;
  assign n3215 = n687 & ~n3214;
  assign n3216 = n264 & ~n2411;
  assign n3217 = n290 & ~n2397;
  assign n3218 = ~n3216 & ~n3217;
  assign n3219 = n317 & ~n2445;
  assign n3220 = n343 & ~n2431;
  assign n3221 = ~n3219 & ~n3220;
  assign n3222 = n3218 & n3221;
  assign n3223 = n582 & ~n3222;
  assign n3224 = ~n3215 & ~n3223;
  assign n3225 = n264 & ~n2531;
  assign n3226 = n290 & ~n2517;
  assign n3227 = ~n3225 & ~n3226;
  assign n3228 = n317 & ~n2623;
  assign n3229 = n343 & ~n2609;
  assign n3230 = ~n3228 & ~n3229;
  assign n3231 = n3227 & n3230;
  assign n3232 = n476 & ~n3231;
  assign n3233 = n264 & ~n2652;
  assign n3234 = n290 & ~n2638;
  assign n3235 = ~n3233 & ~n3234;
  assign n3236 = n317 & ~n2563;
  assign n3237 = n343 & ~n2549;
  assign n3238 = ~n3236 & ~n3237;
  assign n3239 = n3235 & n3238;
  assign n3240 = n371 & ~n3239;
  assign n3241 = ~n3232 & ~n3240;
  assign n3242 = n3224 & n3241;
  assign n3243 = pi134  & ~n3242;
  assign n3244 = ~n3207 & ~n3243;
  assign n3245 = n264 & n4574;
  assign n3246 = n290 & n4584;
  assign n3247 = ~n3245 & ~n3246;
  assign n3248 = n4549 & n317;
  assign n3249 = n343 & n4579;
  assign n3250 = ~n3248 & ~n3249;
  assign n3251 = n3247 & n3250;
  assign n3252 = n371 & ~n3251;
  assign n3253 = n264 & n4614;
  assign n3254 = n290 & n4624;
  assign n3255 = ~n3253 & ~n3254;
  assign n3256 = n317 & n4569;
  assign n3257 = n343 & n4619;
  assign n3258 = ~n3256 & ~n3257;
  assign n3259 = n3255 & n3258;
  assign n3260 = n476 & ~n3259;
  assign n3261 = ~n3252 & ~n3260;
  assign n3262 = n264 & n4634;
  assign n3263 = n290 & n4644;
  assign n3264 = ~n3262 & ~n3263;
  assign n3265 = n317 & n4589;
  assign n3266 = n343 & n4639;
  assign n3267 = ~n3265 & ~n3266;
  assign n3268 = n3264 & n3267;
  assign n3269 = n582 & ~n3268;
  assign n3270 = n264 & n4594;
  assign n3271 = n290 & n4604;
  assign n3272 = ~n3270 & ~n3271;
  assign n3273 = n317 & n4609;
  assign n3274 = n343 & n4599;
  assign n3275 = ~n3273 & ~n3274;
  assign n3276 = n3272 & n3275;
  assign n3277 = n687 & ~n3276;
  assign n3278 = ~n3269 & ~n3277;
  assign n3279 = n3261 & n3278;
  assign n3280 = ~pi134  & ~n3279;
  assign n3281 = n264 & n4674;
  assign n3282 = n290 & n4684;
  assign n3283 = ~n3281 & ~n3282;
  assign n3284 = n317 & n4689;
  assign n3285 = n343 & n4679;
  assign n3286 = ~n3284 & ~n3285;
  assign n3287 = n3283 & n3286;
  assign n3288 = n687 & ~n3287;
  assign n3289 = n264 & n4554;
  assign n3290 = n290 & n4564;
  assign n3291 = ~n3289 & ~n3290;
  assign n3292 = n317 & n4669;
  assign n3293 = n4559 & n343;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = n3291 & n3294;
  assign n3296 = n582 & ~n3295;
  assign n3297 = ~n3288 & ~n3296;
  assign n3298 = n264 & n4694;
  assign n3299 = n290 & ~n1097;
  assign n3300 = ~n3298 & ~n3299;
  assign n3301 = n317 & n4649;
  assign n3302 = n343 & n4699;
  assign n3303 = ~n3301 & ~n3302;
  assign n3304 = n3300 & n3303;
  assign n3305 = n476 & ~n3304;
  assign n3306 = n264 & n4654;
  assign n3307 = n290 & n4664;
  assign n3308 = ~n3306 & ~n3307;
  assign n3309 = n317 & n4629;
  assign n3310 = n343 & n4659;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = n3308 & n3311;
  assign n3313 = n371 & ~n3312;
  assign n3314 = ~n3305 & ~n3313;
  assign n3315 = n3297 & n3314;
  assign n3316 = pi134  & ~n3315;
  assign n3317 = ~n3280 & ~n3316;
  assign n3318 = n264 & ~n1216;
  assign n3319 = n290 & ~n1253;
  assign n3320 = ~n3318 & ~n3319;
  assign n3321 = n317 & ~n1122;
  assign n3322 = n343 & ~n1235;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = n3320 & n3323;
  assign n3325 = n371 & ~n3324;
  assign n3326 = n264 & ~n1369;
  assign n3327 = n290 & ~n1406;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = n317 & ~n1198;
  assign n3330 = n343 & ~n1388;
  assign n3331 = ~n3329 & ~n3330;
  assign n3332 = n3328 & n3331;
  assign n3333 = n476 & ~n3332;
  assign n3334 = ~n3325 & ~n3333;
  assign n3335 = n264 & ~n1524;
  assign n3336 = n290 & ~n1561;
  assign n3337 = ~n3335 & ~n3336;
  assign n3338 = n317 & ~n1275;
  assign n3339 = n343 & ~n1543;
  assign n3340 = ~n3338 & ~n3339;
  assign n3341 = n3337 & n3340;
  assign n3342 = n582 & ~n3341;
  assign n3343 = n264 & ~n1293;
  assign n3344 = n290 & ~n1330;
  assign n3345 = ~n3343 & ~n3344;
  assign n3346 = n317 & ~n1351;
  assign n3347 = n343 & ~n1312;
  assign n3348 = ~n3346 & ~n3347;
  assign n3349 = n3345 & n3348;
  assign n3350 = n687 & ~n3349;
  assign n3351 = ~n3342 & ~n3350;
  assign n3352 = n3334 & n3351;
  assign n3353 = ~pi134  & ~n3352;
  assign n3354 = n264 & ~n1448;
  assign n3355 = n290 & ~n1485;
  assign n3356 = ~n3354 & ~n3355;
  assign n3357 = n317 & ~n1583;
  assign n3358 = n343 & ~n1467;
  assign n3359 = ~n3357 & ~n3358;
  assign n3360 = n3356 & n3359;
  assign n3361 = n687 & ~n3360;
  assign n3362 = n264 & ~n1140;
  assign n3363 = n290 & ~n1177;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = n317 & ~n1430;
  assign n3366 = n343 & ~n1159;
  assign n3367 = ~n3365 & ~n3366;
  assign n3368 = n3364 & n3367;
  assign n3369 = n582 & ~n3368;
  assign n3370 = ~n3361 & ~n3369;
  assign n3371 = n264 & ~n1602;
  assign n3372 = n290 & ~n1637;
  assign n3373 = ~n3371 & ~n3372;
  assign n3374 = n317 & ~n1658;
  assign n3375 = n343 & ~n1621;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = n3373 & n3376;
  assign n3378 = n476 & ~n3377;
  assign n3379 = n264 & ~n1676;
  assign n3380 = n290 & ~n1713;
  assign n3381 = ~n3379 & ~n3380;
  assign n3382 = n317 & ~n1506;
  assign n3383 = n343 & ~n1695;
  assign n3384 = ~n3382 & ~n3383;
  assign n3385 = n3381 & n3384;
  assign n3386 = n371 & ~n3385;
  assign n3387 = ~n3378 & ~n3386;
  assign n3388 = n3370 & n3387;
  assign n3389 = pi134  & ~n3388;
  assign n3390 = ~n3353 & ~n3389;
  assign n3391 = n264 & n4784;
  assign n3392 = n290 & n4790;
  assign n3393 = ~n3391 & ~n3392;
  assign n3394 = n317 & n4769;
  assign n3395 = n343 & n4787;
  assign n3396 = ~n3394 & ~n3395;
  assign n3397 = n3393 & n3396;
  assign n3398 = n371 & ~n3397;
  assign n3399 = n264 & n4808;
  assign n3400 = n290 & n4814;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = n317 & n4781;
  assign n3403 = n343 & n4811;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = n3401 & n3404;
  assign n3406 = n476 & ~n3405;
  assign n3407 = ~n3398 & ~n3406;
  assign n3408 = n264 & n4832;
  assign n3409 = n290 & n4838;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = n317 & n4793;
  assign n3412 = n343 & n4835;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = n3410 & n3413;
  assign n3415 = n582 & ~n3414;
  assign n3416 = n264 & n4796;
  assign n3417 = n290 & n4802;
  assign n3418 = ~n3416 & ~n3417;
  assign n3419 = n317 & n4805;
  assign n3420 = n343 & n4799;
  assign n3421 = ~n3419 & ~n3420;
  assign n3422 = n3418 & n3421;
  assign n3423 = n687 & ~n3422;
  assign n3424 = ~n3415 & ~n3423;
  assign n3425 = n3407 & n3424;
  assign n3426 = ~pi134  & ~n3425;
  assign n3427 = n264 & n4820;
  assign n3428 = n290 & n4826;
  assign n3429 = ~n3427 & ~n3428;
  assign n3430 = n317 & n4841;
  assign n3431 = n343 & n4823;
  assign n3432 = ~n3430 & ~n3431;
  assign n3433 = n3429 & n3432;
  assign n3434 = n687 & ~n3433;
  assign n3435 = n264 & n4772;
  assign n3436 = n290 & n4778;
  assign n3437 = ~n3435 & ~n3436;
  assign n3438 = n317 & n4817;
  assign n3439 = n343 & n4775;
  assign n3440 = ~n3438 & ~n3439;
  assign n3441 = n3437 & n3440;
  assign n3442 = n582 & ~n3441;
  assign n3443 = ~n3434 & ~n3442;
  assign n3444 = n264 & n4844;
  assign n3445 = n290 & ~n2110;
  assign n3446 = ~n3444 & ~n3445;
  assign n3447 = n317 & n4851;
  assign n3448 = n343 & ~n2099;
  assign n3449 = ~n3447 & ~n3448;
  assign n3450 = n3446 & n3449;
  assign n3451 = n476 & ~n3450;
  assign n3452 = n264 & n4854;
  assign n3453 = n290 & n4860;
  assign n3454 = ~n3452 & ~n3453;
  assign n3455 = n317 & n4829;
  assign n3456 = n343 & n4857;
  assign n3457 = ~n3455 & ~n3456;
  assign n3458 = n3454 & n3457;
  assign n3459 = n371 & ~n3458;
  assign n3460 = ~n3451 & ~n3459;
  assign n3461 = n3443 & n3460;
  assign n3462 = pi134  & ~n3461;
  assign n3463 = ~n3426 & ~n3462;
  assign n3464 = n264 & ~n2261;
  assign n3465 = n290 & ~n2290;
  assign n3466 = ~n3464 & ~n3465;
  assign n3467 = n317 & ~n2368;
  assign n3468 = n343 & ~n2276;
  assign n3469 = ~n3467 & ~n3468;
  assign n3470 = n3466 & n3469;
  assign n3471 = n371 & ~n3470;
  assign n3472 = n264 & ~n2201;
  assign n3473 = n290 & ~n2230;
  assign n3474 = ~n3472 & ~n3473;
  assign n3475 = n317 & ~n2247;
  assign n3476 = n343 & ~n2216;
  assign n3477 = ~n3475 & ~n3476;
  assign n3478 = n3474 & n3477;
  assign n3479 = n476 & ~n3478;
  assign n3480 = ~n3471 & ~n3479;
  assign n3481 = n264 & ~n2563;
  assign n3482 = n290 & ~n2592;
  assign n3483 = ~n3481 & ~n3482;
  assign n3484 = n317 & ~n2308;
  assign n3485 = n343 & ~n2578;
  assign n3486 = ~n3484 & ~n3485;
  assign n3487 = n3483 & n3486;
  assign n3488 = n582 & ~n3487;
  assign n3489 = n264 & ~n2322;
  assign n3490 = n290 & ~n2351;
  assign n3491 = ~n3489 & ~n3490;
  assign n3492 = n317 & ~n2187;
  assign n3493 = n343 & ~n2337;
  assign n3494 = ~n3492 & ~n3493;
  assign n3495 = n3491 & n3494;
  assign n3496 = n687 & ~n3495;
  assign n3497 = ~n3488 & ~n3496;
  assign n3498 = n3480 & n3497;
  assign n3499 = ~pi134  & ~n3498;
  assign n3500 = n264 & ~n2445;
  assign n3501 = n290 & ~n2474;
  assign n3502 = ~n3500 & ~n3501;
  assign n3503 = n317 & ~n2491;
  assign n3504 = n343 & ~n2460;
  assign n3505 = ~n3503 & ~n3504;
  assign n3506 = n3502 & n3505;
  assign n3507 = n687 & ~n3506;
  assign n3508 = n264 & ~n2382;
  assign n3509 = n290 & ~n2411;
  assign n3510 = ~n3508 & ~n3509;
  assign n3511 = n317 & ~n2431;
  assign n3512 = n343 & ~n2397;
  assign n3513 = ~n3511 & ~n3512;
  assign n3514 = n3510 & n3513;
  assign n3515 = n582 & ~n3514;
  assign n3516 = ~n3507 & ~n3515;
  assign n3517 = n264 & ~n2502;
  assign n3518 = n290 & ~n2531;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520 = n317 & ~n2609;
  assign n3521 = n343 & ~n2517;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = n3519 & n3522;
  assign n3524 = n476 & ~n3523;
  assign n3525 = n264 & ~n2623;
  assign n3526 = n290 & ~n2652;
  assign n3527 = ~n3525 & ~n3526;
  assign n3528 = n317 & ~n2549;
  assign n3529 = n343 & ~n2638;
  assign n3530 = ~n3528 & ~n3529;
  assign n3531 = n3527 & n3530;
  assign n3532 = n371 & ~n3531;
  assign n3533 = ~n3524 & ~n3532;
  assign n3534 = n3516 & n3533;
  assign n3535 = pi134  & ~n3534;
  assign n3536 = ~n3499 & ~n3535;
  assign n3537 = n371 & ~n475;
  assign n3538 = n476 & ~n686;
  assign n3539 = ~n3537 & ~n3538;
  assign n3540 = n582 & ~n794;
  assign n3541 = ~n581 & n687;
  assign n3542 = ~n3540 & ~n3541;
  assign n3543 = n3539 & n3542;
  assign n3544 = ~pi134  & ~n3543;
  assign n3545 = ~n370 & n582;
  assign n3546 = n371 & ~n898;
  assign n3547 = ~n3545 & ~n3546;
  assign n3548 = n687 & ~n1003;
  assign n3549 = n476 & ~n1100;
  assign n3550 = ~n3548 & ~n3549;
  assign n3551 = n3547 & n3550;
  assign n3552 = pi134  & ~n3551;
  assign n3553 = ~n3544 & ~n3552;
  assign n3554 = n371 & ~n1256;
  assign n3555 = n476 & ~n1409;
  assign n3556 = ~n3554 & ~n3555;
  assign n3557 = n582 & ~n1564;
  assign n3558 = n687 & ~n1333;
  assign n3559 = ~n3557 & ~n3558;
  assign n3560 = n3556 & n3559;
  assign n3561 = ~pi134  & ~n3560;
  assign n3562 = n687 & ~n1488;
  assign n3563 = n582 & ~n1180;
  assign n3564 = ~n3562 & ~n3563;
  assign n3565 = n476 & ~n1640;
  assign n3566 = n371 & ~n1716;
  assign n3567 = ~n3565 & ~n3566;
  assign n3568 = n3564 & n3567;
  assign n3569 = pi134  & ~n3568;
  assign n3570 = ~n3561 & ~n3569;
  assign n3571 = n371 & ~n1832;
  assign n3572 = n476 & ~n1945;
  assign n3573 = ~n3571 & ~n3572;
  assign n3574 = n582 & ~n2060;
  assign n3575 = n687 & ~n1889;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = n3573 & n3576;
  assign n3578 = ~pi134  & ~n3577;
  assign n3579 = n687 & ~n2004;
  assign n3580 = n582 & ~n1776;
  assign n3581 = ~n3579 & ~n3580;
  assign n3582 = n476 & ~n2113;
  assign n3583 = n371 & ~n2169;
  assign n3584 = ~n3582 & ~n3583;
  assign n3585 = n3581 & n3584;
  assign n3586 = pi134  & ~n3585;
  assign n3587 = ~n3578 & ~n3586;
  assign n3588 = n476 & ~n2233;
  assign n3589 = n371 & ~n2293;
  assign n3590 = ~n3588 & ~n3589;
  assign n3591 = n687 & ~n2354;
  assign n3592 = n582 & ~n2595;
  assign n3593 = ~n3591 & ~n3592;
  assign n3594 = n3590 & n3593;
  assign n3595 = ~pi134  & ~n3594;
  assign n3596 = n687 & ~n2477;
  assign n3597 = n582 & ~n2414;
  assign n3598 = ~n3596 & ~n3597;
  assign n3599 = n371 & ~n2655;
  assign n3600 = n476 & ~n2534;
  assign n3601 = ~n3599 & ~n3600;
  assign n3602 = n3598 & n3601;
  assign n3603 = pi134  & ~n3602;
  assign n3604 = ~n3595 & ~n3603;
  assign n3605 = n371 & ~n2675;
  assign n3606 = n476 & ~n2692;
  assign n3607 = ~n3605 & ~n3606;
  assign n3608 = n582 & ~n2728;
  assign n3609 = n687 & ~n2684;
  assign n3610 = ~n3608 & ~n3609;
  assign n3611 = n3607 & n3610;
  assign n3612 = ~pi134  & ~n3611;
  assign n3613 = n582 & ~n2667;
  assign n3614 = n476 & ~n2703;
  assign n3615 = ~n3613 & ~n3614;
  assign n3616 = n371 & ~n2720;
  assign n3617 = n687 & ~n2711;
  assign n3618 = ~n3616 & ~n3617;
  assign n3619 = n3615 & n3618;
  assign n3620 = pi134  & ~n3619;
  assign n3621 = ~n3612 & ~n3620;
  assign n3622 = n371 & ~n2748;
  assign n3623 = n476 & ~n2765;
  assign n3624 = ~n3622 & ~n3623;
  assign n3625 = n582 & ~n2801;
  assign n3626 = n687 & ~n2757;
  assign n3627 = ~n3625 & ~n3626;
  assign n3628 = n3624 & n3627;
  assign n3629 = ~pi134  & ~n3628;
  assign n3630 = n582 & ~n2740;
  assign n3631 = n476 & ~n2776;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = n371 & ~n2793;
  assign n3634 = n687 & ~n2784;
  assign n3635 = ~n3633 & ~n3634;
  assign n3636 = n3632 & n3635;
  assign n3637 = pi134  & ~n3636;
  assign n3638 = ~n3629 & ~n3637;
  assign n3639 = n371 & ~n2821;
  assign n3640 = n476 & ~n2838;
  assign n3641 = ~n3639 & ~n3640;
  assign n3642 = n582 & ~n2874;
  assign n3643 = n687 & ~n2830;
  assign n3644 = ~n3642 & ~n3643;
  assign n3645 = n3641 & n3644;
  assign n3646 = ~pi134  & ~n3645;
  assign n3647 = n582 & ~n2813;
  assign n3648 = n476 & ~n2849;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = n371 & ~n2866;
  assign n3651 = n687 & ~n2857;
  assign n3652 = ~n3650 & ~n3651;
  assign n3653 = n3649 & n3652;
  assign n3654 = pi134  & ~n3653;
  assign n3655 = ~n3646 & ~n3654;
  assign n3656 = n371 & ~n2894;
  assign n3657 = n582 & ~n2947;
  assign n3658 = ~n3656 & ~n3657;
  assign n3659 = n687 & ~n2903;
  assign n3660 = n476 & ~n2911;
  assign n3661 = ~n3659 & ~n3660;
  assign n3662 = n3658 & n3661;
  assign n3663 = ~pi134  & ~n3662;
  assign n3664 = n476 & ~n2922;
  assign n3665 = n687 & ~n2930;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = n371 & ~n2939;
  assign n3668 = n582 & ~n2886;
  assign n3669 = ~n3667 & ~n3668;
  assign n3670 = n3666 & n3669;
  assign n3671 = pi134  & ~n3670;
  assign n3672 = ~n3663 & ~n3671;
  assign n3673 = n371 & ~n2967;
  assign n3674 = n582 & ~n3020;
  assign n3675 = ~n3673 & ~n3674;
  assign n3676 = n687 & ~n2976;
  assign n3677 = n476 & ~n2984;
  assign n3678 = ~n3676 & ~n3677;
  assign n3679 = n3675 & n3678;
  assign n3680 = ~pi134  & ~n3679;
  assign n3681 = n476 & ~n2995;
  assign n3682 = n687 & ~n3003;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = n371 & ~n3012;
  assign n3685 = n582 & ~n2959;
  assign n3686 = ~n3684 & ~n3685;
  assign n3687 = n3683 & n3686;
  assign n3688 = pi134  & ~n3687;
  assign n3689 = ~n3680 & ~n3688;
  assign n3690 = n371 & ~n3040;
  assign n3691 = n582 & ~n3093;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = n687 & ~n3049;
  assign n3694 = n476 & ~n3057;
  assign n3695 = ~n3693 & ~n3694;
  assign n3696 = n3692 & n3695;
  assign n3697 = ~pi134  & ~n3696;
  assign n3698 = n476 & ~n3068;
  assign n3699 = n687 & ~n3076;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = n371 & ~n3085;
  assign n3702 = n582 & ~n3032;
  assign n3703 = ~n3701 & ~n3702;
  assign n3704 = n3700 & n3703;
  assign n3705 = pi134  & ~n3704;
  assign n3706 = ~n3697 & ~n3705;
  assign n3707 = n371 & ~n3113;
  assign n3708 = n476 & ~n3130;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = n582 & ~n3166;
  assign n3711 = n687 & ~n3122;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = n3709 & n3712;
  assign n3714 = ~pi134  & ~n3713;
  assign n3715 = n476 & ~n3141;
  assign n3716 = n687 & ~n3149;
  assign n3717 = ~n3715 & ~n3716;
  assign n3718 = n371 & ~n3158;
  assign n3719 = n582 & ~n3105;
  assign n3720 = ~n3718 & ~n3719;
  assign n3721 = n3717 & n3720;
  assign n3722 = pi134  & ~n3721;
  assign n3723 = ~n3714 & ~n3722;
  assign n3724 = n371 & ~n3186;
  assign n3725 = n476 & ~n3203;
  assign n3726 = ~n3724 & ~n3725;
  assign n3727 = n582 & ~n3239;
  assign n3728 = n687 & ~n3195;
  assign n3729 = ~n3727 & ~n3728;
  assign n3730 = n3726 & n3729;
  assign n3731 = ~pi134  & ~n3730;
  assign n3732 = n476 & ~n3214;
  assign n3733 = n687 & ~n3222;
  assign n3734 = ~n3732 & ~n3733;
  assign n3735 = n371 & ~n3231;
  assign n3736 = n582 & ~n3178;
  assign n3737 = ~n3735 & ~n3736;
  assign n3738 = n3734 & n3737;
  assign n3739 = pi134  & ~n3738;
  assign n3740 = ~n3731 & ~n3739;
  assign n3741 = n371 & ~n3259;
  assign n3742 = n476 & ~n3276;
  assign n3743 = ~n3741 & ~n3742;
  assign n3744 = n582 & ~n3312;
  assign n3745 = n687 & ~n3268;
  assign n3746 = ~n3744 & ~n3745;
  assign n3747 = n3743 & n3746;
  assign n3748 = ~pi134  & ~n3747;
  assign n3749 = n476 & ~n3287;
  assign n3750 = n687 & ~n3295;
  assign n3751 = ~n3749 & ~n3750;
  assign n3752 = n371 & ~n3304;
  assign n3753 = n582 & ~n3251;
  assign n3754 = ~n3752 & ~n3753;
  assign n3755 = n3751 & n3754;
  assign n3756 = pi134  & ~n3755;
  assign n3757 = ~n3748 & ~n3756;
  assign n3758 = n371 & ~n3332;
  assign n3759 = n476 & ~n3349;
  assign n3760 = ~n3758 & ~n3759;
  assign n3761 = n582 & ~n3385;
  assign n3762 = n687 & ~n3341;
  assign n3763 = ~n3761 & ~n3762;
  assign n3764 = n3760 & n3763;
  assign n3765 = ~pi134  & ~n3764;
  assign n3766 = n476 & ~n3360;
  assign n3767 = n687 & ~n3368;
  assign n3768 = ~n3766 & ~n3767;
  assign n3769 = n371 & ~n3377;
  assign n3770 = n582 & ~n3324;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = n3768 & n3771;
  assign n3773 = pi134  & ~n3772;
  assign n3774 = ~n3765 & ~n3773;
  assign n3775 = n371 & ~n3405;
  assign n3776 = n476 & ~n3422;
  assign n3777 = ~n3775 & ~n3776;
  assign n3778 = n582 & ~n3458;
  assign n3779 = n687 & ~n3414;
  assign n3780 = ~n3778 & ~n3779;
  assign n3781 = n3777 & n3780;
  assign n3782 = ~pi134  & ~n3781;
  assign n3783 = n476 & ~n3433;
  assign n3784 = n687 & ~n3441;
  assign n3785 = ~n3783 & ~n3784;
  assign n3786 = n371 & ~n3450;
  assign n3787 = n582 & ~n3397;
  assign n3788 = ~n3786 & ~n3787;
  assign n3789 = n3785 & n3788;
  assign n3790 = pi134  & ~n3789;
  assign n3791 = ~n3782 & ~n3790;
  assign n3792 = n371 & ~n3478;
  assign n3793 = n476 & ~n3495;
  assign n3794 = ~n3792 & ~n3793;
  assign n3795 = n582 & ~n3531;
  assign n3796 = n687 & ~n3487;
  assign n3797 = ~n3795 & ~n3796;
  assign n3798 = n3794 & n3797;
  assign n3799 = ~pi134  & ~n3798;
  assign n3800 = n476 & ~n3506;
  assign n3801 = n687 & ~n3514;
  assign n3802 = ~n3800 & ~n3801;
  assign n3803 = n371 & ~n3523;
  assign n3804 = n582 & ~n3470;
  assign n3805 = ~n3803 & ~n3804;
  assign n3806 = n3802 & n3805;
  assign n3807 = pi134  & ~n3806;
  assign n3808 = ~n3799 & ~n3807;
  assign n3809 = n371 & ~n686;
  assign n3810 = n476 & ~n581;
  assign n3811 = ~n3809 & ~n3810;
  assign n3812 = n582 & ~n898;
  assign n3813 = n687 & ~n794;
  assign n3814 = ~n3812 & ~n3813;
  assign n3815 = n3811 & n3814;
  assign n3816 = ~pi134  & ~n3815;
  assign n3817 = ~n370 & n687;
  assign n3818 = ~n475 & n582;
  assign n3819 = ~n3817 & ~n3818;
  assign n3820 = n476 & ~n1003;
  assign n3821 = n371 & ~n1100;
  assign n3822 = ~n3820 & ~n3821;
  assign n3823 = n3819 & n3822;
  assign n3824 = pi134  & ~n3823;
  assign n3825 = ~n3816 & ~n3824;
  assign n3826 = n371 & ~n1409;
  assign n3827 = n476 & ~n1333;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = n582 & ~n1716;
  assign n3830 = n687 & ~n1564;
  assign n3831 = ~n3829 & ~n3830;
  assign n3832 = n3828 & n3831;
  assign n3833 = ~pi134  & ~n3832;
  assign n3834 = n476 & ~n1488;
  assign n3835 = n687 & ~n1180;
  assign n3836 = ~n3834 & ~n3835;
  assign n3837 = n371 & ~n1640;
  assign n3838 = n582 & ~n1256;
  assign n3839 = ~n3837 & ~n3838;
  assign n3840 = n3836 & n3839;
  assign n3841 = pi134  & ~n3840;
  assign n3842 = ~n3833 & ~n3841;
  assign n3843 = n371 & ~n1945;
  assign n3844 = n476 & ~n1889;
  assign n3845 = ~n3843 & ~n3844;
  assign n3846 = n582 & ~n2169;
  assign n3847 = n687 & ~n2060;
  assign n3848 = ~n3846 & ~n3847;
  assign n3849 = n3845 & n3848;
  assign n3850 = ~pi134  & ~n3849;
  assign n3851 = n476 & ~n2004;
  assign n3852 = n687 & ~n1776;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = n371 & ~n2113;
  assign n3855 = n582 & ~n1832;
  assign n3856 = ~n3854 & ~n3855;
  assign n3857 = n3853 & n3856;
  assign n3858 = pi134  & ~n3857;
  assign n3859 = ~n3850 & ~n3858;
  assign n3860 = n371 & ~n2233;
  assign n3861 = n582 & ~n2655;
  assign n3862 = ~n3860 & ~n3861;
  assign n3863 = n476 & ~n2354;
  assign n3864 = n687 & ~n2595;
  assign n3865 = ~n3863 & ~n3864;
  assign n3866 = n3862 & n3865;
  assign n3867 = ~pi134  & ~n3866;
  assign n3868 = n476 & ~n2477;
  assign n3869 = n582 & ~n2293;
  assign n3870 = ~n3868 & ~n3869;
  assign n3871 = n371 & ~n2534;
  assign n3872 = n687 & ~n2414;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = n3870 & n3873;
  assign n3875 = pi134  & ~n3874;
  assign n3876 = ~n3867 & ~n3875;
  assign n3877 = n371 & ~n2692;
  assign n3878 = n476 & ~n2684;
  assign n3879 = ~n3877 & ~n3878;
  assign n3880 = n582 & ~n2720;
  assign n3881 = n687 & ~n2728;
  assign n3882 = ~n3880 & ~n3881;
  assign n3883 = n3879 & n3882;
  assign n3884 = ~pi134  & ~n3883;
  assign n3885 = n687 & ~n2667;
  assign n3886 = n582 & ~n2675;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = n476 & ~n2711;
  assign n3889 = n371 & ~n2703;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = n3887 & n3890;
  assign n3892 = pi134  & ~n3891;
  assign n3893 = ~n3884 & ~n3892;
  assign n3894 = n371 & ~n2765;
  assign n3895 = n476 & ~n2757;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = n582 & ~n2793;
  assign n3898 = n687 & ~n2801;
  assign n3899 = ~n3897 & ~n3898;
  assign n3900 = n3896 & n3899;
  assign n3901 = ~pi134  & ~n3900;
  assign n3902 = n687 & ~n2740;
  assign n3903 = n582 & ~n2748;
  assign n3904 = ~n3902 & ~n3903;
  assign n3905 = n476 & ~n2784;
  assign n3906 = n371 & ~n2776;
  assign n3907 = ~n3905 & ~n3906;
  assign n3908 = n3904 & n3907;
  assign n3909 = pi134  & ~n3908;
  assign n3910 = ~n3901 & ~n3909;
  assign n3911 = n371 & ~n2838;
  assign n3912 = n476 & ~n2830;
  assign n3913 = ~n3911 & ~n3912;
  assign n3914 = n582 & ~n2866;
  assign n3915 = n687 & ~n2874;
  assign n3916 = ~n3914 & ~n3915;
  assign n3917 = n3913 & n3916;
  assign n3918 = ~pi134  & ~n3917;
  assign n3919 = n687 & ~n2813;
  assign n3920 = n582 & ~n2821;
  assign n3921 = ~n3919 & ~n3920;
  assign n3922 = n476 & ~n2857;
  assign n3923 = n371 & ~n2849;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = n3921 & n3924;
  assign n3926 = pi134  & ~n3925;
  assign n3927 = ~n3918 & ~n3926;
  assign n3928 = n687 & ~n2947;
  assign n3929 = n582 & ~n2939;
  assign n3930 = ~n3928 & ~n3929;
  assign n3931 = n476 & ~n2903;
  assign n3932 = n371 & ~n2911;
  assign n3933 = ~n3931 & ~n3932;
  assign n3934 = n3930 & n3933;
  assign n3935 = ~pi134  & ~n3934;
  assign n3936 = n371 & ~n2922;
  assign n3937 = n476 & ~n2930;
  assign n3938 = ~n3936 & ~n3937;
  assign n3939 = n582 & ~n2894;
  assign n3940 = n687 & ~n2886;
  assign n3941 = ~n3939 & ~n3940;
  assign n3942 = n3938 & n3941;
  assign n3943 = pi134  & ~n3942;
  assign n3944 = ~n3935 & ~n3943;
  assign n3945 = n687 & ~n3020;
  assign n3946 = n582 & ~n3012;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = n476 & ~n2976;
  assign n3949 = n371 & ~n2984;
  assign n3950 = ~n3948 & ~n3949;
  assign n3951 = n3947 & n3950;
  assign n3952 = ~pi134  & ~n3951;
  assign n3953 = n371 & ~n2995;
  assign n3954 = n476 & ~n3003;
  assign n3955 = ~n3953 & ~n3954;
  assign n3956 = n582 & ~n2967;
  assign n3957 = n687 & ~n2959;
  assign n3958 = ~n3956 & ~n3957;
  assign n3959 = n3955 & n3958;
  assign n3960 = pi134  & ~n3959;
  assign n3961 = ~n3952 & ~n3960;
  assign n3962 = n687 & ~n3093;
  assign n3963 = n582 & ~n3085;
  assign n3964 = ~n3962 & ~n3963;
  assign n3965 = n476 & ~n3049;
  assign n3966 = n371 & ~n3057;
  assign n3967 = ~n3965 & ~n3966;
  assign n3968 = n3964 & n3967;
  assign n3969 = ~pi134  & ~n3968;
  assign n3970 = n371 & ~n3068;
  assign n3971 = n476 & ~n3076;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = n582 & ~n3040;
  assign n3974 = n687 & ~n3032;
  assign n3975 = ~n3973 & ~n3974;
  assign n3976 = n3972 & n3975;
  assign n3977 = pi134  & ~n3976;
  assign n3978 = ~n3969 & ~n3977;
  assign n3979 = n371 & ~n3130;
  assign n3980 = n476 & ~n3122;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = n582 & ~n3158;
  assign n3983 = n687 & ~n3166;
  assign n3984 = ~n3982 & ~n3983;
  assign n3985 = n3981 & n3984;
  assign n3986 = ~pi134  & ~n3985;
  assign n3987 = n371 & ~n3141;
  assign n3988 = n476 & ~n3149;
  assign n3989 = ~n3987 & ~n3988;
  assign n3990 = n582 & ~n3113;
  assign n3991 = n687 & ~n3105;
  assign n3992 = ~n3990 & ~n3991;
  assign n3993 = n3989 & n3992;
  assign n3994 = pi134  & ~n3993;
  assign n3995 = ~n3986 & ~n3994;
  assign n3996 = n371 & ~n3203;
  assign n3997 = n476 & ~n3195;
  assign n3998 = ~n3996 & ~n3997;
  assign n3999 = n582 & ~n3231;
  assign n4000 = n687 & ~n3239;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = n3998 & n4001;
  assign n4003 = ~pi134  & ~n4002;
  assign n4004 = n371 & ~n3214;
  assign n4005 = n476 & ~n3222;
  assign n4006 = ~n4004 & ~n4005;
  assign n4007 = n582 & ~n3186;
  assign n4008 = n687 & ~n3178;
  assign n4009 = ~n4007 & ~n4008;
  assign n4010 = n4006 & n4009;
  assign n4011 = pi134  & ~n4010;
  assign n4012 = ~n4003 & ~n4011;
  assign n4013 = n371 & ~n3276;
  assign n4014 = n476 & ~n3268;
  assign n4015 = ~n4013 & ~n4014;
  assign n4016 = n582 & ~n3304;
  assign n4017 = n687 & ~n3312;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = n4015 & n4018;
  assign n4020 = ~pi134  & ~n4019;
  assign n4021 = n371 & ~n3287;
  assign n4022 = n476 & ~n3295;
  assign n4023 = ~n4021 & ~n4022;
  assign n4024 = n582 & ~n3259;
  assign n4025 = n687 & ~n3251;
  assign n4026 = ~n4024 & ~n4025;
  assign n4027 = n4023 & n4026;
  assign n4028 = pi134  & ~n4027;
  assign n4029 = ~n4020 & ~n4028;
  assign n4030 = n371 & ~n3349;
  assign n4031 = n476 & ~n3341;
  assign n4032 = ~n4030 & ~n4031;
  assign n4033 = n582 & ~n3377;
  assign n4034 = n687 & ~n3385;
  assign n4035 = ~n4033 & ~n4034;
  assign n4036 = n4032 & n4035;
  assign n4037 = ~pi134  & ~n4036;
  assign n4038 = n371 & ~n3360;
  assign n4039 = n476 & ~n3368;
  assign n4040 = ~n4038 & ~n4039;
  assign n4041 = n582 & ~n3332;
  assign n4042 = n687 & ~n3324;
  assign n4043 = ~n4041 & ~n4042;
  assign n4044 = n4040 & n4043;
  assign n4045 = pi134  & ~n4044;
  assign n4046 = ~n4037 & ~n4045;
  assign n4047 = n371 & ~n3422;
  assign n4048 = n476 & ~n3414;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = n582 & ~n3450;
  assign n4051 = n687 & ~n3458;
  assign n4052 = ~n4050 & ~n4051;
  assign n4053 = n4049 & n4052;
  assign n4054 = ~pi134  & ~n4053;
  assign n4055 = n371 & ~n3433;
  assign n4056 = n476 & ~n3441;
  assign n4057 = ~n4055 & ~n4056;
  assign n4058 = n582 & ~n3405;
  assign n4059 = n687 & ~n3397;
  assign n4060 = ~n4058 & ~n4059;
  assign n4061 = n4057 & n4060;
  assign n4062 = pi134  & ~n4061;
  assign n4063 = ~n4054 & ~n4062;
  assign n4064 = n371 & ~n3495;
  assign n4065 = n476 & ~n3487;
  assign n4066 = ~n4064 & ~n4065;
  assign n4067 = n582 & ~n3523;
  assign n4068 = n687 & ~n3531;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = n4066 & n4069;
  assign n4071 = ~pi134  & ~n4070;
  assign n4072 = n371 & ~n3506;
  assign n4073 = n476 & ~n3514;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = n582 & ~n3478;
  assign n4076 = n687 & ~n3470;
  assign n4077 = ~n4075 & ~n4076;
  assign n4078 = n4074 & n4077;
  assign n4079 = pi134  & ~n4078;
  assign n4080 = ~n4071 & ~n4079;
  assign n4081 = n371 & ~n581;
  assign n4082 = n476 & ~n794;
  assign n4083 = ~n4081 & ~n4082;
  assign n4084 = n582 & ~n1100;
  assign n4085 = n687 & ~n898;
  assign n4086 = ~n4084 & ~n4085;
  assign n4087 = n4083 & n4086;
  assign n4088 = ~pi134  & ~n4087;
  assign n4089 = ~n370 & n476;
  assign n4090 = ~n475 & n687;
  assign n4091 = ~n4089 & ~n4090;
  assign n4092 = n371 & ~n1003;
  assign n4093 = n582 & ~n686;
  assign n4094 = ~n4092 & ~n4093;
  assign n4095 = n4091 & n4094;
  assign n4096 = pi134  & ~n4095;
  assign n4097 = ~n4088 & ~n4096;
  assign n4098 = n371 & ~n1333;
  assign n4099 = n476 & ~n1564;
  assign n4100 = ~n4098 & ~n4099;
  assign n4101 = n582 & ~n1640;
  assign n4102 = n687 & ~n1716;
  assign n4103 = ~n4101 & ~n4102;
  assign n4104 = n4100 & n4103;
  assign n4105 = ~pi134  & ~n4104;
  assign n4106 = n371 & ~n1488;
  assign n4107 = n476 & ~n1180;
  assign n4108 = ~n4106 & ~n4107;
  assign n4109 = n582 & ~n1409;
  assign n4110 = n687 & ~n1256;
  assign n4111 = ~n4109 & ~n4110;
  assign n4112 = n4108 & n4111;
  assign n4113 = pi134  & ~n4112;
  assign n4114 = ~n4105 & ~n4113;
  assign n4115 = n371 & ~n1889;
  assign n4116 = n476 & ~n2060;
  assign n4117 = ~n4115 & ~n4116;
  assign n4118 = n582 & ~n2113;
  assign n4119 = n687 & ~n2169;
  assign n4120 = ~n4118 & ~n4119;
  assign n4121 = n4117 & n4120;
  assign n4122 = ~pi134  & ~n4121;
  assign n4123 = n371 & ~n2004;
  assign n4124 = n476 & ~n1776;
  assign n4125 = ~n4123 & ~n4124;
  assign n4126 = n582 & ~n1945;
  assign n4127 = n687 & ~n1832;
  assign n4128 = ~n4126 & ~n4127;
  assign n4129 = n4125 & n4128;
  assign n4130 = pi134  & ~n4129;
  assign n4131 = ~n4122 & ~n4130;
  assign n4132 = n582 & ~n2534;
  assign n4133 = n687 & ~n2655;
  assign n4134 = ~n4132 & ~n4133;
  assign n4135 = n371 & ~n2354;
  assign n4136 = n476 & ~n2595;
  assign n4137 = ~n4135 & ~n4136;
  assign n4138 = n4134 & n4137;
  assign n4139 = ~pi134  & ~n4138;
  assign n4140 = n371 & ~n2477;
  assign n4141 = n582 & ~n2233;
  assign n4142 = ~n4140 & ~n4141;
  assign n4143 = n476 & ~n2414;
  assign n4144 = n687 & ~n2293;
  assign n4145 = ~n4143 & ~n4144;
  assign n4146 = n4142 & n4145;
  assign n4147 = pi134  & ~n4146;
  assign n4148 = ~n4139 & ~n4147;
  assign n4149 = n582 & ~n2703;
  assign n4150 = n371 & ~n2684;
  assign n4151 = ~n4149 & ~n4150;
  assign n4152 = n687 & ~n2720;
  assign n4153 = n476 & ~n2728;
  assign n4154 = ~n4152 & ~n4153;
  assign n4155 = n4151 & n4154;
  assign n4156 = ~pi134  & ~n4155;
  assign n4157 = n476 & ~n2667;
  assign n4158 = n687 & ~n2675;
  assign n4159 = ~n4157 & ~n4158;
  assign n4160 = n582 & ~n2692;
  assign n4161 = n371 & ~n2711;
  assign n4162 = ~n4160 & ~n4161;
  assign n4163 = n4159 & n4162;
  assign n4164 = pi134  & ~n4163;
  assign n4165 = ~n4156 & ~n4164;
  assign n4166 = n582 & ~n2776;
  assign n4167 = n371 & ~n2757;
  assign n4168 = ~n4166 & ~n4167;
  assign n4169 = n687 & ~n2793;
  assign n4170 = n476 & ~n2801;
  assign n4171 = ~n4169 & ~n4170;
  assign n4172 = n4168 & n4171;
  assign n4173 = ~pi134  & ~n4172;
  assign n4174 = n476 & ~n2740;
  assign n4175 = n687 & ~n2748;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = n582 & ~n2765;
  assign n4178 = n371 & ~n2784;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180 = n4176 & n4179;
  assign n4181 = pi134  & ~n4180;
  assign n4182 = ~n4173 & ~n4181;
  assign n4183 = n582 & ~n2849;
  assign n4184 = n371 & ~n2830;
  assign n4185 = ~n4183 & ~n4184;
  assign n4186 = n687 & ~n2866;
  assign n4187 = n476 & ~n2874;
  assign n4188 = ~n4186 & ~n4187;
  assign n4189 = n4185 & n4188;
  assign n4190 = ~pi134  & ~n4189;
  assign n4191 = n476 & ~n2813;
  assign n4192 = n687 & ~n2821;
  assign n4193 = ~n4191 & ~n4192;
  assign n4194 = n582 & ~n2838;
  assign n4195 = n371 & ~n2857;
  assign n4196 = ~n4194 & ~n4195;
  assign n4197 = n4193 & n4196;
  assign n4198 = pi134  & ~n4197;
  assign n4199 = ~n4190 & ~n4198;
  assign n4200 = n582 & ~n2922;
  assign n4201 = n476 & ~n2947;
  assign n4202 = ~n4200 & ~n4201;
  assign n4203 = n371 & ~n2903;
  assign n4204 = n687 & ~n2939;
  assign n4205 = ~n4203 & ~n4204;
  assign n4206 = n4202 & n4205;
  assign n4207 = ~pi134  & ~n4206;
  assign n4208 = n371 & ~n2930;
  assign n4209 = n476 & ~n2886;
  assign n4210 = ~n4208 & ~n4209;
  assign n4211 = n582 & ~n2911;
  assign n4212 = n687 & ~n2894;
  assign n4213 = ~n4211 & ~n4212;
  assign n4214 = n4210 & n4213;
  assign n4215 = pi134  & ~n4214;
  assign n4216 = ~n4207 & ~n4215;
  assign n4217 = n582 & ~n2995;
  assign n4218 = n476 & ~n3020;
  assign n4219 = ~n4217 & ~n4218;
  assign n4220 = n371 & ~n2976;
  assign n4221 = n687 & ~n3012;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = n4219 & n4222;
  assign n4224 = ~pi134  & ~n4223;
  assign n4225 = n371 & ~n3003;
  assign n4226 = n476 & ~n2959;
  assign n4227 = ~n4225 & ~n4226;
  assign n4228 = n582 & ~n2984;
  assign n4229 = n687 & ~n2967;
  assign n4230 = ~n4228 & ~n4229;
  assign n4231 = n4227 & n4230;
  assign n4232 = pi134  & ~n4231;
  assign n4233 = ~n4224 & ~n4232;
  assign n4234 = n582 & ~n3068;
  assign n4235 = n476 & ~n3093;
  assign n4236 = ~n4234 & ~n4235;
  assign n4237 = n371 & ~n3049;
  assign n4238 = n687 & ~n3085;
  assign n4239 = ~n4237 & ~n4238;
  assign n4240 = n4236 & n4239;
  assign n4241 = ~pi134  & ~n4240;
  assign n4242 = n371 & ~n3076;
  assign n4243 = n476 & ~n3032;
  assign n4244 = ~n4242 & ~n4243;
  assign n4245 = n582 & ~n3057;
  assign n4246 = n687 & ~n3040;
  assign n4247 = ~n4245 & ~n4246;
  assign n4248 = n4244 & n4247;
  assign n4249 = pi134  & ~n4248;
  assign n4250 = ~n4241 & ~n4249;
  assign n4251 = n582 & ~n3141;
  assign n4252 = n371 & ~n3122;
  assign n4253 = ~n4251 & ~n4252;
  assign n4254 = n687 & ~n3158;
  assign n4255 = n476 & ~n3166;
  assign n4256 = ~n4254 & ~n4255;
  assign n4257 = n4253 & n4256;
  assign n4258 = ~pi134  & ~n4257;
  assign n4259 = n371 & ~n3149;
  assign n4260 = n476 & ~n3105;
  assign n4261 = ~n4259 & ~n4260;
  assign n4262 = n582 & ~n3130;
  assign n4263 = n687 & ~n3113;
  assign n4264 = ~n4262 & ~n4263;
  assign n4265 = n4261 & n4264;
  assign n4266 = pi134  & ~n4265;
  assign n4267 = ~n4258 & ~n4266;
  assign n4268 = n582 & ~n3214;
  assign n4269 = n371 & ~n3195;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = n687 & ~n3231;
  assign n4272 = n476 & ~n3239;
  assign n4273 = ~n4271 & ~n4272;
  assign n4274 = n4270 & n4273;
  assign n4275 = ~pi134  & ~n4274;
  assign n4276 = n371 & ~n3222;
  assign n4277 = n476 & ~n3178;
  assign n4278 = ~n4276 & ~n4277;
  assign n4279 = n582 & ~n3203;
  assign n4280 = n687 & ~n3186;
  assign n4281 = ~n4279 & ~n4280;
  assign n4282 = n4278 & n4281;
  assign n4283 = pi134  & ~n4282;
  assign n4284 = ~n4275 & ~n4283;
  assign n4285 = n582 & ~n3287;
  assign n4286 = n371 & ~n3268;
  assign n4287 = ~n4285 & ~n4286;
  assign n4288 = n687 & ~n3304;
  assign n4289 = n476 & ~n3312;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = n4287 & n4290;
  assign n4292 = ~pi134  & ~n4291;
  assign n4293 = n371 & ~n3295;
  assign n4294 = n476 & ~n3251;
  assign n4295 = ~n4293 & ~n4294;
  assign n4296 = n582 & ~n3276;
  assign n4297 = n687 & ~n3259;
  assign n4298 = ~n4296 & ~n4297;
  assign n4299 = n4295 & n4298;
  assign n4300 = pi134  & ~n4299;
  assign n4301 = ~n4292 & ~n4300;
  assign n4302 = n582 & ~n3360;
  assign n4303 = n371 & ~n3341;
  assign n4304 = ~n4302 & ~n4303;
  assign n4305 = n687 & ~n3377;
  assign n4306 = n476 & ~n3385;
  assign n4307 = ~n4305 & ~n4306;
  assign n4308 = n4304 & n4307;
  assign n4309 = ~pi134  & ~n4308;
  assign n4310 = n371 & ~n3368;
  assign n4311 = n476 & ~n3324;
  assign n4312 = ~n4310 & ~n4311;
  assign n4313 = n582 & ~n3349;
  assign n4314 = n687 & ~n3332;
  assign n4315 = ~n4313 & ~n4314;
  assign n4316 = n4312 & n4315;
  assign n4317 = pi134  & ~n4316;
  assign n4318 = ~n4309 & ~n4317;
  assign n4319 = n582 & ~n3433;
  assign n4320 = n371 & ~n3414;
  assign n4321 = ~n4319 & ~n4320;
  assign n4322 = n687 & ~n3450;
  assign n4323 = n476 & ~n3458;
  assign n4324 = ~n4322 & ~n4323;
  assign n4325 = n4321 & n4324;
  assign n4326 = ~pi134  & ~n4325;
  assign n4327 = n371 & ~n3441;
  assign n4328 = n476 & ~n3397;
  assign n4329 = ~n4327 & ~n4328;
  assign n4330 = n582 & ~n3422;
  assign n4331 = n687 & ~n3405;
  assign n4332 = ~n4330 & ~n4331;
  assign n4333 = n4329 & n4332;
  assign n4334 = pi134  & ~n4333;
  assign n4335 = ~n4326 & ~n4334;
  assign n4336 = n582 & ~n3506;
  assign n4337 = n371 & ~n3487;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = n687 & ~n3523;
  assign n4340 = n476 & ~n3531;
  assign n4341 = ~n4339 & ~n4340;
  assign n4342 = n4338 & n4341;
  assign n4343 = ~pi134  & ~n4342;
  assign n4344 = n371 & ~n3514;
  assign n4345 = n476 & ~n3470;
  assign n4346 = ~n4344 & ~n4345;
  assign n4347 = n582 & ~n3495;
  assign n4348 = n687 & ~n3478;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = n4346 & n4349;
  assign n4351 = pi134  & ~n4350;
  assign n4352 = ~n4343 & ~n4351;
  assign n4353 = ~pi134  & ~n1103;
  assign n4354 = pi134  & ~n690;
  assign n4355 = ~n4353 & ~n4354;
  assign n4356 = ~pi134  & ~n1719;
  assign n4357 = pi134  & ~n1412;
  assign n4358 = ~n4356 & ~n4357;
  assign n4359 = ~pi134  & ~n2172;
  assign n4360 = pi134  & ~n1948;
  assign n4361 = ~n4359 & ~n4360;
  assign n4362 = ~pi134  & ~n2658;
  assign n4363 = pi134  & ~n2417;
  assign n4364 = ~n4362 & ~n4363;
  assign n4365 = ~pi134  & ~n2731;
  assign n4366 = pi134  & ~n2695;
  assign n4367 = ~n4365 & ~n4366;
  assign n4368 = ~pi134  & ~n2804;
  assign n4369 = pi134  & ~n2768;
  assign n4370 = ~n4368 & ~n4369;
  assign n4371 = ~pi134  & ~n2877;
  assign n4372 = pi134  & ~n2841;
  assign n4373 = ~n4371 & ~n4372;
  assign n4374 = ~pi134  & ~n2950;
  assign n4375 = pi134  & ~n2914;
  assign n4376 = ~n4374 & ~n4375;
  assign n4377 = ~pi134  & ~n3023;
  assign n4378 = pi134  & ~n2987;
  assign n4379 = ~n4377 & ~n4378;
  assign n4380 = ~pi134  & ~n3096;
  assign n4381 = pi134  & ~n3060;
  assign n4382 = ~n4380 & ~n4381;
  assign n4383 = ~pi134  & ~n3169;
  assign n4384 = pi134  & ~n3133;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = ~pi134  & ~n3242;
  assign n4387 = pi134  & ~n3206;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = ~pi134  & ~n3315;
  assign n4390 = pi134  & ~n3279;
  assign n4391 = ~n4389 & ~n4390;
  assign n4392 = ~pi134  & ~n3388;
  assign n4393 = pi134  & ~n3352;
  assign n4394 = ~n4392 & ~n4393;
  assign n4395 = ~pi134  & ~n3461;
  assign n4396 = pi134  & ~n3425;
  assign n4397 = ~n4395 & ~n4396;
  assign n4398 = ~pi134  & ~n3534;
  assign n4399 = pi134  & ~n3498;
  assign n4400 = ~n4398 & ~n4399;
  assign n4401 = ~pi134  & ~n3551;
  assign n4402 = pi134  & ~n3543;
  assign n4403 = ~n4401 & ~n4402;
  assign n4404 = ~pi134  & ~n3568;
  assign n4405 = pi134  & ~n3560;
  assign n4406 = ~n4404 & ~n4405;
  assign n4407 = ~pi134  & ~n3585;
  assign n4408 = pi134  & ~n3577;
  assign n4409 = ~n4407 & ~n4408;
  assign n4410 = ~pi134  & ~n3602;
  assign n4411 = pi134  & ~n3594;
  assign n4412 = ~n4410 & ~n4411;
  assign n4413 = ~pi134  & ~n3619;
  assign n4414 = pi134  & ~n3611;
  assign n4415 = ~n4413 & ~n4414;
  assign n4416 = ~pi134  & ~n3636;
  assign n4417 = pi134  & ~n3628;
  assign n4418 = ~n4416 & ~n4417;
  assign n4419 = ~pi134  & ~n3653;
  assign n4420 = pi134  & ~n3645;
  assign n4421 = ~n4419 & ~n4420;
  assign n4422 = ~pi134  & ~n3670;
  assign n4423 = pi134  & ~n3662;
  assign n4424 = ~n4422 & ~n4423;
  assign n4425 = ~pi134  & ~n3687;
  assign n4426 = pi134  & ~n3679;
  assign n4427 = ~n4425 & ~n4426;
  assign n4428 = ~pi134  & ~n3704;
  assign n4429 = pi134  & ~n3696;
  assign n4430 = ~n4428 & ~n4429;
  assign n4431 = ~pi134  & ~n3721;
  assign n4432 = pi134  & ~n3713;
  assign n4433 = ~n4431 & ~n4432;
  assign n4434 = ~pi134  & ~n3738;
  assign n4435 = pi134  & ~n3730;
  assign n4436 = ~n4434 & ~n4435;
  assign n4437 = ~pi134  & ~n3755;
  assign n4438 = pi134  & ~n3747;
  assign n4439 = ~n4437 & ~n4438;
  assign n4440 = ~pi134  & ~n3772;
  assign n4441 = pi134  & ~n3764;
  assign n4442 = ~n4440 & ~n4441;
  assign n4443 = ~pi134  & ~n3789;
  assign n4444 = pi134  & ~n3781;
  assign n4445 = ~n4443 & ~n4444;
  assign n4446 = ~pi134  & ~n3806;
  assign n4447 = pi134  & ~n3798;
  assign n4448 = ~n4446 & ~n4447;
  assign n4449 = ~pi134  & ~n3823;
  assign n4450 = pi134  & ~n3815;
  assign n4451 = ~n4449 & ~n4450;
  assign n4452 = ~pi134  & ~n3840;
  assign n4453 = pi134  & ~n3832;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = ~pi134  & ~n3857;
  assign n4456 = pi134  & ~n3849;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = ~pi134  & ~n3874;
  assign n4459 = pi134  & ~n3866;
  assign n4460 = ~n4458 & ~n4459;
  assign n4461 = ~pi134  & ~n3891;
  assign n4462 = pi134  & ~n3883;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = ~pi134  & ~n3908;
  assign n4465 = pi134  & ~n3900;
  assign n4466 = ~n4464 & ~n4465;
  assign n4467 = ~pi134  & ~n3925;
  assign n4468 = pi134  & ~n3917;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = ~pi134  & ~n3942;
  assign n4471 = pi134  & ~n3934;
  assign n4472 = ~n4470 & ~n4471;
  assign n4473 = ~pi134  & ~n3959;
  assign n4474 = pi134  & ~n3951;
  assign n4475 = ~n4473 & ~n4474;
  assign n4476 = ~pi134  & ~n3976;
  assign n4477 = pi134  & ~n3968;
  assign n4478 = ~n4476 & ~n4477;
  assign n4479 = ~pi134  & ~n3993;
  assign n4480 = pi134  & ~n3985;
  assign n4481 = ~n4479 & ~n4480;
  assign n4482 = ~pi134  & ~n4010;
  assign n4483 = pi134  & ~n4002;
  assign n4484 = ~n4482 & ~n4483;
  assign n4485 = ~pi134  & ~n4027;
  assign n4486 = pi134  & ~n4019;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = ~pi134  & ~n4044;
  assign n4489 = pi134  & ~n4036;
  assign n4490 = ~n4488 & ~n4489;
  assign n4491 = ~pi134  & ~n4061;
  assign n4492 = pi134  & ~n4053;
  assign n4493 = ~n4491 & ~n4492;
  assign n4494 = ~pi134  & ~n4078;
  assign n4495 = pi134  & ~n4070;
  assign n4496 = ~n4494 & ~n4495;
  assign n4497 = ~pi134  & ~n4095;
  assign n4498 = pi134  & ~n4087;
  assign n4499 = ~n4497 & ~n4498;
  assign n4500 = ~pi134  & ~n4112;
  assign n4501 = pi134  & ~n4104;
  assign n4502 = ~n4500 & ~n4501;
  assign n4503 = ~pi134  & ~n4129;
  assign n4504 = pi134  & ~n4121;
  assign n4505 = ~n4503 & ~n4504;
  assign n4506 = ~pi134  & ~n4146;
  assign n4507 = pi134  & ~n4138;
  assign n4508 = ~n4506 & ~n4507;
  assign n4509 = ~pi134  & ~n4163;
  assign n4510 = pi134  & ~n4155;
  assign n4511 = ~n4509 & ~n4510;
  assign n4512 = ~pi134  & ~n4180;
  assign n4513 = pi134  & ~n4172;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = ~pi134  & ~n4197;
  assign n4516 = pi134  & ~n4189;
  assign n4517 = ~n4515 & ~n4516;
  assign n4518 = ~pi134  & ~n4214;
  assign n4519 = pi134  & ~n4206;
  assign n4520 = ~n4518 & ~n4519;
  assign n4521 = ~pi134  & ~n4231;
  assign n4522 = pi134  & ~n4223;
  assign n4523 = ~n4521 & ~n4522;
  assign n4524 = ~pi134  & ~n4248;
  assign n4525 = pi134  & ~n4240;
  assign n4526 = ~n4524 & ~n4525;
  assign n4527 = ~pi134  & ~n4265;
  assign n4528 = pi134  & ~n4257;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = ~pi134  & ~n4282;
  assign n4531 = pi134  & ~n4274;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = ~pi134  & ~n4299;
  assign n4534 = pi134  & ~n4291;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = ~pi134  & ~n4316;
  assign n4537 = pi134  & ~n4308;
  assign n4538 = ~n4536 & ~n4537;
  assign n4539 = ~pi134  & ~n4333;
  assign n4540 = pi134  & ~n4325;
  assign n4541 = ~n4539 & ~n4540;
  assign n4542 = ~pi134  & ~n4350;
  assign n4543 = pi134  & ~n4342;
  assign n4544 = ~n4542 & ~n4543;
  assign n4545 = n269 | ~n270;
  assign n4546 = n273 | ~n274;
  assign n4547 = n279 | ~n280;
  assign n4548 = n283 | ~n284;
  assign n4549 = n287 | ~n288;
  assign n4550 = n295 | ~n296;
  assign n4551 = n299 | ~n300;
  assign n4552 = n305 | ~n306;
  assign n4553 = n309 | ~n310;
  assign n4554 = n313 | ~n314;
  assign n4555 = n322 | ~n323;
  assign n4556 = n326 | ~n327;
  assign n4557 = n332 | ~n333;
  assign n4558 = n336 | ~n337;
  assign n4559 = n340 | ~n341;
  assign n4560 = n348 | ~n349;
  assign n4561 = n352 | ~n353;
  assign n4562 = n358 | ~n359;
  assign n4563 = n362 | ~n363;
  assign n4564 = n366 | ~n367;
  assign n4565 = n377 | ~n378;
  assign n4566 = n381 | ~n382;
  assign n4567 = n387 | ~n388;
  assign n4568 = n391 | ~n392;
  assign n4569 = n395 | ~n396;
  assign n4570 = n402 | ~n403;
  assign n4571 = n406 | ~n407;
  assign n4572 = n412 | ~n413;
  assign n4573 = n416 | ~n417;
  assign n4574 = n420 | ~n421;
  assign n4575 = n428 | ~n429;
  assign n4576 = n432 | ~n433;
  assign n4577 = n438 | ~n439;
  assign n4578 = n442 | ~n443;
  assign n4579 = n446 | ~n447;
  assign n4580 = n453 | ~n454;
  assign n4581 = n457 | ~n458;
  assign n4582 = n463 | ~n464;
  assign n4583 = n467 | ~n468;
  assign n4584 = n471 | ~n472;
  assign n4585 = n483 | ~n484;
  assign n4586 = n487 | ~n488;
  assign n4587 = n493 | ~n494;
  assign n4588 = n497 | ~n498;
  assign n4589 = n501 | ~n502;
  assign n4590 = n508 | ~n509;
  assign n4591 = n512 | ~n513;
  assign n4592 = n518 | ~n519;
  assign n4593 = n522 | ~n523;
  assign n4594 = n526 | ~n527;
  assign n4595 = n534 | ~n535;
  assign n4596 = n538 | ~n539;
  assign n4597 = n544 | ~n545;
  assign n4598 = n548 | ~n549;
  assign n4599 = n552 | ~n553;
  assign n4600 = n559 | ~n560;
  assign n4601 = n563 | ~n564;
  assign n4602 = n569 | ~n570;
  assign n4603 = n573 | ~n574;
  assign n4604 = n577 | ~n578;
  assign n4605 = n588 | ~n589;
  assign n4606 = n592 | ~n593;
  assign n4607 = n598 | ~n599;
  assign n4608 = n602 | ~n603;
  assign n4609 = n606 | ~n607;
  assign n4610 = n613 | ~n614;
  assign n4611 = n617 | ~n618;
  assign n4612 = n623 | ~n624;
  assign n4613 = n627 | ~n628;
  assign n4614 = n631 | ~n632;
  assign n4615 = n639 | ~n640;
  assign n4616 = n643 | ~n644;
  assign n4617 = n649 | ~n650;
  assign n4618 = n653 | ~n654;
  assign n4619 = n657 | ~n658;
  assign n4620 = n664 | ~n665;
  assign n4621 = n668 | ~n669;
  assign n4622 = n674 | ~n675;
  assign n4623 = n678 | ~n679;
  assign n4624 = n682 | ~n683;
  assign n4625 = n696 | ~n697;
  assign n4626 = n700 | ~n701;
  assign n4627 = n706 | ~n707;
  assign n4628 = n710 | ~n711;
  assign n4629 = n714 | ~n715;
  assign n4630 = n721 | ~n722;
  assign n4631 = n725 | ~n726;
  assign n4632 = n731 | ~n732;
  assign n4633 = n735 | ~n736;
  assign n4634 = n739 | ~n740;
  assign n4635 = n747 | ~n748;
  assign n4636 = n751 | ~n752;
  assign n4637 = n757 | ~n758;
  assign n4638 = n761 | ~n762;
  assign n4639 = n765 | ~n766;
  assign n4640 = n772 | ~n773;
  assign n4641 = n776 | ~n777;
  assign n4642 = n782 | ~n783;
  assign n4643 = n786 | ~n787;
  assign n4644 = n790 | ~n791;
  assign n4645 = n800 | ~n801;
  assign n4646 = n804 | ~n805;
  assign n4647 = n810 | ~n811;
  assign n4648 = n814 | ~n815;
  assign n4649 = n818 | ~n819;
  assign n4650 = n825 | ~n826;
  assign n4651 = n829 | ~n830;
  assign n4652 = n835 | ~n836;
  assign n4653 = n839 | ~n840;
  assign n4654 = n843 | ~n844;
  assign n4655 = n851 | ~n852;
  assign n4656 = n855 | ~n856;
  assign n4657 = n861 | ~n862;
  assign n4658 = n865 | ~n866;
  assign n4659 = n869 | ~n870;
  assign n4660 = n876 | ~n877;
  assign n4661 = n880 | ~n881;
  assign n4662 = n886 | ~n887;
  assign n4663 = n890 | ~n891;
  assign n4664 = n894 | ~n895;
  assign n4665 = n905 | ~n906;
  assign n4666 = n909 | ~n910;
  assign n4667 = n915 | ~n916;
  assign n4668 = n919 | ~n920;
  assign n4669 = n923 | ~n924;
  assign n4670 = n930 | ~n931;
  assign n4671 = n934 | ~n935;
  assign n4672 = n940 | ~n941;
  assign n4673 = n944 | ~n945;
  assign n4674 = n948 | ~n949;
  assign n4675 = n956 | ~n957;
  assign n4676 = n960 | ~n961;
  assign n4677 = n966 | ~n967;
  assign n4678 = n970 | ~n971;
  assign n4679 = n974 | ~n975;
  assign n4680 = n981 | ~n982;
  assign n4681 = n985 | ~n986;
  assign n4682 = n991 | ~n992;
  assign n4683 = n995 | ~n996;
  assign n4684 = n999 | ~n1000;
  assign n4685 = n1009 | ~n1010;
  assign n4686 = n1013 | ~n1014;
  assign n4687 = n1019 | ~n1020;
  assign n4688 = n1023 | ~n1024;
  assign n4689 = n1027 | ~n1028;
  assign n4690 = n1034 | ~n1035;
  assign n4691 = n1038 | ~n1039;
  assign n4692 = n1044 | ~n1045;
  assign n4693 = n1048 | ~n1049;
  assign n4694 = n1052 | ~n1053;
  assign n4695 = n1060 | ~n1061;
  assign n4696 = n1064 | ~n1065;
  assign n4697 = n1070 | ~n1071;
  assign n4698 = n1074 | ~n1075;
  assign n4699 = n1078 | ~n1079;
  assign n4700 = n1087 | ~n1088;
  assign n4701 = n1095 | ~n1096;
  assign n4702 = n1112 | ~n1113;
  assign n4703 = n1120 | ~n1121;
  assign n4704 = n1130 | ~n1131;
  assign n4705 = n1138 | ~n1139;
  assign n4706 = n1149 | ~n1150;
  assign n4707 = n1157 | ~n1158;
  assign n4708 = n1167 | ~n1168;
  assign n4709 = n1175 | ~n1176;
  assign n4710 = n1188 | ~n1189;
  assign n4711 = n1196 | ~n1197;
  assign n4712 = n1206 | ~n1207;
  assign n4713 = n1214 | ~n1215;
  assign n4714 = n1225 | ~n1226;
  assign n4715 = n1233 | ~n1234;
  assign n4716 = n1243 | ~n1244;
  assign n4717 = n1251 | ~n1252;
  assign n4718 = n1265 | ~n1266;
  assign n4719 = n1273 | ~n1274;
  assign n4720 = n1283 | ~n1284;
  assign n4721 = n1291 | ~n1292;
  assign n4722 = n1302 | ~n1303;
  assign n4723 = n1310 | ~n1311;
  assign n4724 = n1320 | ~n1321;
  assign n4725 = n1328 | ~n1329;
  assign n4726 = n1341 | ~n1342;
  assign n4727 = n1349 | ~n1350;
  assign n4728 = n1359 | ~n1360;
  assign n4729 = n1367 | ~n1368;
  assign n4730 = n1378 | ~n1379;
  assign n4731 = n1386 | ~n1387;
  assign n4732 = n1396 | ~n1397;
  assign n4733 = n1404 | ~n1405;
  assign n4734 = n1420 | ~n1421;
  assign n4735 = n1428 | ~n1429;
  assign n4736 = n1438 | ~n1439;
  assign n4737 = n1446 | ~n1447;
  assign n4738 = n1457 | ~n1458;
  assign n4739 = n1465 | ~n1466;
  assign n4740 = n1475 | ~n1476;
  assign n4741 = n1483 | ~n1484;
  assign n4742 = n1496 | ~n1497;
  assign n4743 = n1504 | ~n1505;
  assign n4744 = n1514 | ~n1515;
  assign n4745 = n1522 | ~n1523;
  assign n4746 = n1533 | ~n1534;
  assign n4747 = n1541 | ~n1542;
  assign n4748 = n1551 | ~n1552;
  assign n4749 = n1559 | ~n1560;
  assign n4750 = n1573 | ~n1574;
  assign n4751 = n1581 | ~n1582;
  assign n4752 = n1590 | ~n1591;
  assign n4753 = n1596 | ~n1597;
  assign n4754 = n1600 | ~n1601;
  assign n4755 = n1611 | ~n1612;
  assign n4756 = n1619 | ~n1620;
  assign n4757 = n1628 | ~n1629;
  assign n4758 = n1635 | ~n1636;
  assign n4759 = n1648 | ~n1649;
  assign n4760 = n1656 | ~n1657;
  assign n4761 = n1666 | ~n1667;
  assign n4762 = n1674 | ~n1675;
  assign n4763 = n1685 | ~n1686;
  assign n4764 = n1693 | ~n1694;
  assign n4765 = n1703 | ~n1704;
  assign n4766 = n1711 | ~n1712;
  assign n4767 = n1724 | ~n1725;
  assign n4768 = n1728 | ~n1729;
  assign n4769 = n1732 | ~n1733;
  assign n4770 = n1737 | ~n1738;
  assign n4771 = n1741 | ~n1742;
  assign n4772 = n1745 | ~n1746;
  assign n4773 = n1751 | ~n1752;
  assign n4774 = n1755 | ~n1756;
  assign n4775 = n1759 | ~n1760;
  assign n4776 = n1764 | ~n1765;
  assign n4777 = n1768 | ~n1769;
  assign n4778 = n1772 | ~n1773;
  assign n4779 = n1780 | ~n1781;
  assign n4780 = n1784 | ~n1785;
  assign n4781 = n1788 | ~n1789;
  assign n4782 = n1793 | ~n1794;
  assign n4783 = n1797 | ~n1798;
  assign n4784 = n1801 | ~n1802;
  assign n4785 = n1807 | ~n1808;
  assign n4786 = n1811 | ~n1812;
  assign n4787 = n1815 | ~n1816;
  assign n4788 = n1820 | ~n1821;
  assign n4789 = n1824 | ~n1825;
  assign n4790 = n1828 | ~n1829;
  assign n4791 = n1837 | ~n1838;
  assign n4792 = n1841 | ~n1842;
  assign n4793 = n1845 | ~n1846;
  assign n4794 = n1850 | ~n1851;
  assign n4795 = n1854 | ~n1855;
  assign n4796 = n1858 | ~n1859;
  assign n4797 = n1864 | ~n1865;
  assign n4798 = n1868 | ~n1869;
  assign n4799 = n1872 | ~n1873;
  assign n4800 = n1877 | ~n1878;
  assign n4801 = n1881 | ~n1882;
  assign n4802 = n1885 | ~n1886;
  assign n4803 = n1893 | ~n1894;
  assign n4804 = n1897 | ~n1898;
  assign n4805 = n1901 | ~n1902;
  assign n4806 = n1906 | ~n1907;
  assign n4807 = n1910 | ~n1911;
  assign n4808 = n1914 | ~n1915;
  assign n4809 = n1920 | ~n1921;
  assign n4810 = n1924 | ~n1925;
  assign n4811 = n1928 | ~n1929;
  assign n4812 = n1933 | ~n1934;
  assign n4813 = n1937 | ~n1938;
  assign n4814 = n1941 | ~n1942;
  assign n4815 = n1952 | ~n1953;
  assign n4816 = n1956 | ~n1957;
  assign n4817 = n1960 | ~n1961;
  assign n4818 = n1965 | ~n1966;
  assign n4819 = n1969 | ~n1970;
  assign n4820 = n1973 | ~n1974;
  assign n4821 = n1979 | ~n1980;
  assign n4822 = n1983 | ~n1984;
  assign n4823 = n1987 | ~n1988;
  assign n4824 = n1992 | ~n1993;
  assign n4825 = n1996 | ~n1997;
  assign n4826 = n2000 | ~n2001;
  assign n4827 = n2008 | ~n2009;
  assign n4828 = n2012 | ~n2013;
  assign n4829 = n2016 | ~n2017;
  assign n4830 = n2021 | ~n2022;
  assign n4831 = n2025 | ~n2026;
  assign n4832 = n2029 | ~n2030;
  assign n4833 = n2035 | ~n2036;
  assign n4834 = n2039 | ~n2040;
  assign n4835 = n2043 | ~n2044;
  assign n4836 = n2048 | ~n2049;
  assign n4837 = n2052 | ~n2053;
  assign n4838 = n2056 | ~n2057;
  assign n4839 = n2065 | ~n2066;
  assign n4840 = n2069 | ~n2070;
  assign n4841 = n2073 | ~n2074;
  assign n4842 = n2078 | ~n2079;
  assign n4843 = n2082 | ~n2083;
  assign n4844 = n2086 | ~n2087;
  assign n4845 = n2093 | ~n2094;
  assign n4846 = n2097 | ~n2098;
  assign n4847 = n2103 | ~n2104;
  assign n4848 = n2108 | ~n2109;
  assign n4849 = n2117 | ~n2118;
  assign n4850 = n2121 | ~n2122;
  assign n4851 = n2125 | ~n2126;
  assign n4852 = n2130 | ~n2131;
  assign n4853 = n2134 | ~n2135;
  assign n4854 = n2138 | ~n2139;
  assign n4855 = n2144 | ~n2145;
  assign n4856 = n2148 | ~n2149;
  assign n4857 = n2152 | ~n2153;
  assign n4858 = n2157 | ~n2158;
  assign n4859 = n2161 | ~n2162;
  assign n4860 = n2165 | ~n2166;
  assign n4861 = n2179 | ~n2180;
  assign n4862 = n2185 | ~n2186;
  assign n4863 = n2193 | ~n2194;
  assign n4864 = n2199 | ~n2200;
  assign n4865 = n2208 | ~n2209;
  assign n4866 = n2214 | ~n2215;
  assign n4867 = n2222 | ~n2223;
  assign n4868 = n2228 | ~n2229;
  assign n4869 = n2239 | ~n2240;
  assign n4870 = n2245 | ~n2246;
  assign n4871 = n2253 | ~n2254;
  assign n4872 = n2259 | ~n2260;
  assign n4873 = n2268 | ~n2269;
  assign n4874 = n2274 | ~n2275;
  assign n4875 = n2282 | ~n2283;
  assign n4876 = n2288 | ~n2289;
  assign n4877 = n2300 | ~n2301;
  assign n4878 = n2306 | ~n2307;
  assign n4879 = n2314 | ~n2315;
  assign n4880 = n2320 | ~n2321;
  assign n4881 = n2329 | ~n2330;
  assign n4882 = n2335 | ~n2336;
  assign n4883 = n2343 | ~n2344;
  assign n4884 = n2349 | ~n2350;
  assign n4885 = n2360 | ~n2361;
  assign n4886 = n2366 | ~n2367;
  assign n4887 = n2374 | ~n2375;
  assign n4888 = n2380 | ~n2381;
  assign n4889 = n2389 | ~n2390;
  assign n4890 = n2395 | ~n2396;
  assign n4891 = n2403 | ~n2404;
  assign n4892 = n2409 | ~n2410;
  assign n4893 = n2423 | ~n2424;
  assign n4894 = n2429 | ~n2430;
  assign n4895 = n2437 | ~n2438;
  assign n4896 = n2443 | ~n2444;
  assign n4897 = n2452 | ~n2453;
  assign n4898 = n2458 | ~n2459;
  assign n4899 = n2466 | ~n2467;
  assign n4900 = n2472 | ~n2473;
  assign n4901 = n2483 | ~n2484;
  assign n4902 = n2489 | ~n2490;
  assign n4903 = n2495 | ~n2496;
  assign n4904 = n2500 | ~n2501;
  assign n4905 = n2509 | ~n2510;
  assign n4906 = n2515 | ~n2516;
  assign n4907 = n2523 | ~n2524;
  assign n4908 = n2529 | ~n2530;
  assign n4909 = n2541 | ~n2542;
  assign n4910 = n2547 | ~n2548;
  assign n4911 = n2555 | ~n2556;
  assign n4912 = n2561 | ~n2562;
  assign n4913 = n2570 | ~n2571;
  assign n4914 = n2576 | ~n2577;
  assign n4915 = n2584 | ~n2585;
  assign n4916 = n2590 | ~n2591;
  assign n4917 = n2601 | ~n2602;
  assign n4918 = n2607 | ~n2608;
  assign n4919 = n2615 | ~n2616;
  assign n4920 = n2621 | ~n2622;
  assign n4921 = n2630 | ~n2631;
  assign n4922 = n2636 | ~n2637;
  assign n4923 = n2644 | ~n2645;
  assign n4924 = n2650 | ~n2651;
  assign po0  = ~n1105;
  assign po1  = ~n1721;
  assign po2  = ~n2174;
  assign po3  = ~n2660;
  assign po4  = ~n2733;
  assign po5  = ~n2806;
  assign po6  = ~n2879;
  assign po7  = ~n2952;
  assign po8  = ~n3025;
  assign po9  = ~n3098;
  assign po10  = ~n3171;
  assign po11  = ~n3244;
  assign po12  = ~n3317;
  assign po13  = ~n3390;
  assign po14  = ~n3463;
  assign po15  = ~n3536;
  assign po16  = ~n3553;
  assign po17  = ~n3570;
  assign po18  = ~n3587;
  assign po19  = ~n3604;
  assign po20  = ~n3621;
  assign po21  = ~n3638;
  assign po22  = ~n3655;
  assign po23  = ~n3672;
  assign po24  = ~n3689;
  assign po25  = ~n3706;
  assign po26  = ~n3723;
  assign po27  = ~n3740;
  assign po28  = ~n3757;
  assign po29  = ~n3774;
  assign po30  = ~n3791;
  assign po31  = ~n3808;
  assign po32  = ~n3825;
  assign po33  = ~n3842;
  assign po34  = ~n3859;
  assign po35  = ~n3876;
  assign po36  = ~n3893;
  assign po37  = ~n3910;
  assign po38  = ~n3927;
  assign po39  = ~n3944;
  assign po40  = ~n3961;
  assign po41  = ~n3978;
  assign po42  = ~n3995;
  assign po43  = ~n4012;
  assign po44  = ~n4029;
  assign po45  = ~n4046;
  assign po46  = ~n4063;
  assign po47  = ~n4080;
  assign po48  = ~n4097;
  assign po49  = ~n4114;
  assign po50  = ~n4131;
  assign po51  = ~n4148;
  assign po52  = ~n4165;
  assign po53  = ~n4182;
  assign po54  = ~n4199;
  assign po55  = ~n4216;
  assign po56  = ~n4233;
  assign po57  = ~n4250;
  assign po58  = ~n4267;
  assign po59  = ~n4284;
  assign po60  = ~n4301;
  assign po61  = ~n4318;
  assign po62  = ~n4335;
  assign po63  = ~n4352;
  assign po64  = ~n4355;
  assign po65  = ~n4358;
  assign po66  = ~n4361;
  assign po67  = ~n4364;
  assign po68  = ~n4367;
  assign po69  = ~n4370;
  assign po70  = ~n4373;
  assign po71  = ~n4376;
  assign po72  = ~n4379;
  assign po73  = ~n4382;
  assign po74  = ~n4385;
  assign po75  = ~n4388;
  assign po76  = ~n4391;
  assign po77  = ~n4394;
  assign po78  = ~n4397;
  assign po79  = ~n4400;
  assign po80  = ~n4403;
  assign po81  = ~n4406;
  assign po82  = ~n4409;
  assign po83  = ~n4412;
  assign po84  = ~n4415;
  assign po85  = ~n4418;
  assign po86  = ~n4421;
  assign po87  = ~n4424;
  assign po88  = ~n4427;
  assign po89  = ~n4430;
  assign po90  = ~n4433;
  assign po91  = ~n4436;
  assign po92  = ~n4439;
  assign po93  = ~n4442;
  assign po94  = ~n4445;
  assign po95  = ~n4448;
  assign po96  = ~n4451;
  assign po97  = ~n4454;
  assign po98  = ~n4457;
  assign po99  = ~n4460;
  assign po100  = ~n4463;
  assign po101  = ~n4466;
  assign po102  = ~n4469;
  assign po103  = ~n4472;
  assign po104  = ~n4475;
  assign po105  = ~n4478;
  assign po106  = ~n4481;
  assign po107  = ~n4484;
  assign po108  = ~n4487;
  assign po109  = ~n4490;
  assign po110  = ~n4493;
  assign po111  = ~n4496;
  assign po112  = ~n4499;
  assign po113  = ~n4502;
  assign po114  = ~n4505;
  assign po115  = ~n4508;
  assign po116  = ~n4511;
  assign po117  = ~n4514;
  assign po118  = ~n4517;
  assign po119  = ~n4520;
  assign po120  = ~n4523;
  assign po121  = ~n4526;
  assign po122  = ~n4529;
  assign po123  = ~n4532;
  assign po124  = ~n4535;
  assign po125  = ~n4538;
  assign po126  = ~n4541;
  assign po127  = ~n4544;
endmodule
