module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 ;
  wire n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102,
    n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396,
    n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426,
    n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894,
    n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924,
    n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170,
    n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182,
    n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200,
    n3201, n3202, n3203, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212,
    n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242,
    n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272,
    n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302,
    n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332,
    n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362,
    n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3390, n3391, n3392,
    n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416,
    n3417, n3418, n3419, n3420, n3421, n3422,
    n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3439, n3440,
    n3441, n3442, n3443, n3444, n3445, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476,
    n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722,
    n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782,
    n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052,
    n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292,
    n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334,
    n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346,
    n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382,
    n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412,
    n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430,
    n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442,
    n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466,
    n4467, n4468, n4469, n4470, n4471, n4472,
    n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496,
    n4497, n4498, n4499, n4500, n4501, n4502,
    n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526,
    n4527, n4528, n4529, n4530, n4531, n4532,
    n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562,
    n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586,
    n4587, n4588, n4589, n4590, n4591, n4592,
    n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622,
    n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700,
    n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708, n4709, n4710, n4711, n4712,
    n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5040, n5041, n5042,
    n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072,
    n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372,
    n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390,
    n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402,
    n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414,
    n5415, n5416, n5417, n5418, n5419, n5420,
    n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5436, n5437, n5438,
    n5439, n5440, n5441, n5442, n5443, n5444,
    n5445, n5446, n5447, n5448, n5449, n5450,
    n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5460, n5461, n5462,
    n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5470, n5471, n5472, n5473, n5474,
    n5475, n5476, n5477, n5478, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528,
    n5529, n5530, n5531, n5532, n5533, n5534,
    n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5542, n5543, n5544, n5545, n5546,
    n5547, n5548, n5549, n5550, n5551, n5552,
    n5553, n5554, n5555, n5556, n5557, n5558,
    n5559, n5560, n5561, n5562, n5563, n5564,
    n5565, n5566, n5567, n5568, n5569, n5570,
    n5571, n5572, n5573, n5574, n5575, n5576,
    n5577, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588,
    n5589, n5590, n5591, n5592, n5593, n5594,
    n5595, n5596, n5597, n5598, n5599, n5600,
    n5601, n5602, n5603, n5604, n5605, n5606,
    n5607, n5608, n5609, n5610, n5611, n5612,
    n5613, n5614, n5615, n5616, n5617, n5618,
    n5619, n5620, n5621, n5622, n5623, n5624,
    n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636,
    n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648,
    n5649, n5650, n5651, n5652, n5653, n5654,
    n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678,
    n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708,
    n5709, n5710, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5718, n5719, n5720,
    n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732,
    n5733, n5734, n5735, n5736, n5737, n5738,
    n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750,
    n5751, n5752, n5753, n5754, n5755, n5756,
    n5757, n5758, n5759, n5760, n5761, n5762,
    n5763, n5764, n5765, n5766, n5767, n5768,
    n5769, n5770, n5771, n5772, n5773, n5774,
    n5775, n5776, n5777, n5778, n5779, n5780,
    n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792,
    n5793, n5794, n5795, n5796, n5797, n5798,
    n5799, n5800, n5801, n5802, n5803, n5804,
    n5805, n5806, n5807, n5808, n5809, n5810,
    n5811, n5812, n5813, n5814, n5815, n5816,
    n5817, n5818, n5819, n5820, n5821, n5822,
    n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5834,
    n5835, n5836, n5837, n5838, n5839, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846,
    n5847, n5848, n5849, n5850, n5851, n5852,
    n5853, n5854, n5855, n5856, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864,
    n5865, n5866, n5867, n5868, n5869, n5870,
    n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882,
    n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894,
    n5895, n5896, n5897, n5898, n5899, n5900,
    n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912,
    n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924,
    n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954,
    n5955, n5956, n5957, n5958, n5959, n5960,
    n5961, n5962, n5963, n5964, n5965, n5966,
    n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5986, n5987, n5988, n5989, n5990,
    n5991, n5992, n5993, n5994, n5995, n5996,
    n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020,
    n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050,
    n6051, n6052, n6053, n6054, n6055, n6056,
    n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074,
    n6075, n6076, n6077, n6078, n6079, n6080,
    n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110,
    n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122,
    n6123, n6124, n6125, n6126, n6127, n6128,
    n6129, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140,
    n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236,
    n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266,
    n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278,
    n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296,
    n6297, n6298, n6299, n6300, n6301, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326,
    n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362,
    n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386,
    n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398,
    n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416,
    n6417, n6418, n6419, n6420, n6421, n6422,
    n6423, n6424, n6425, n6426, n6427, n6428,
    n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446,
    n6447, n6448, n6449, n6450, n6451, n6452,
    n6453, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470,
    n6471, n6472, n6473, n6474, n6475, n6476,
    n6477, n6478, n6479, n6480, n6481, n6482,
    n6483, n6484, n6485, n6486, n6487, n6488,
    n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500,
    n6501, n6502, n6503, n6504, n6505, n6506,
    n6507, n6508, n6509, n6510, n6511, n6512,
    n6513, n6514, n6515, n6516, n6517, n6518,
    n6519, n6520, n6521, n6522, n6523, n6524,
    n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6533, n6534, n6535, n6536,
    n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548,
    n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566,
    n6567, n6568, n6569, n6570, n6571, n6572,
    n6573, n6574, n6575, n6576, n6577, n6578,
    n6579, n6580, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6588, n6589, n6590,
    n6591, n6592, n6593, n6594, n6595, n6596,
    n6597, n6598, n6599, n6600, n6601, n6602,
    n6603, n6604, n6605, n6606, n6607, n6608,
    n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620,
    n6621, n6622, n6623, n6624, n6625, n6626,
    n6627, n6628, n6629, n6630, n6631, n6632,
    n6633, n6634, n6635, n6636, n6637, n6638,
    n6639, n6640, n6641, n6642, n6643, n6644,
    n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902,
    n6903, n6904, n6905, n6906, n6907, n6908,
    n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6937, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962,
    n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992,
    n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112,
    n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136,
    n7137, n7138, n7139, n7140, n7141, n7142,
    n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154,
    n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172,
    n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214,
    n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370,
    n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400,
    n7401, n7402, n7403, n7404, n7405, n7406,
    n7407, n7408, n7409, n7410, n7411, n7412,
    n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430,
    n7431, n7432, n7433, n7434, n7435, n7436,
    n7437, n7438, n7439, n7440, n7441, n7442,
    n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472,
    n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496,
    n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562,
    n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580,
    n7581, n7582, n7583, n7584, n7585, n7586,
    n7587, n7588, n7589, n7590, n7591, n7592,
    n7593, n7594, n7595, n7596, n7597, n7598,
    n7599, n7600, n7601, n7602, n7603, n7604,
    n7605, n7606, n7607, n7608, n7609, n7610,
    n7611, n7612, n7613, n7614, n7615, n7616,
    n7617, n7618, n7619, n7620, n7621, n7622,
    n7623, n7624, n7625, n7626, n7627, n7628,
    n7629, n7630, n7631, n7632, n7633, n7634,
    n7635, n7636, n7637, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7645, n7646,
    n7647, n7648, n7649, n7650, n7651, n7652,
    n7653, n7654, n7655, n7656, n7657, n7658,
    n7659, n7660, n7661, n7662, n7663, n7664,
    n7665, n7666, n7667, n7668, n7669, n7670,
    n7671, n7672, n7673, n7674, n7675, n7676,
    n7677, n7678, n7679, n7680, n7681, n7682,
    n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694,
    n7695, n7696, n7697, n7698, n7699, n7700,
    n7701, n7702, n7703, n7704, n7705, n7706,
    n7707, n7708, n7709, n7710, n7711, n7712,
    n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724,
    n7725, n7726, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7735, n7736,
    n7737, n7738, n7739, n7740, n7741, n7742,
    n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7760,
    n7761, n7762, n7763, n7764, n7765, n7766,
    n7767, n7768, n7769, n7770, n7771, n7772,
    n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790,
    n7791, n7792, n7793, n7794, n7795, n7796,
    n7797, n7798, n7799, n7800, n7801, n7802,
    n7803, n7804, n7805, n7806, n7807, n7808,
    n7809, n7810, n7811, n7812, n7813, n7814,
    n7815, n7816, n7817, n7818, n7819, n7820,
    n7821, n7822, n7823, n7824, n7825, n7826,
    n7827, n7828, n7829, n7830, n7831, n7832,
    n7833, n7834, n7835, n7836, n7837, n7838,
    n7839, n7840, n7841, n7842, n7843, n7844,
    n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7854, n7855, n7856,
    n7857, n7858, n7859, n7860, n7861, n7862,
    n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886,
    n7887, n7888, n7889, n7890, n7891, n7892,
    n7893, n7894, n7895, n7896, n7897, n7898,
    n7899, n7900, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922,
    n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7948, n7949, n7950, n7951, n7952,
    n7953, n7954, n7955, n7956, n7957, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976,
    n7977, n7978, n7979, n7980, n7981, n7982,
    n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012,
    n8013, n8014, n8015, n8016, n8017, n8018,
    n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042,
    n8043, n8044, n8045, n8046, n8047, n8048,
    n8049, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066,
    n8067, n8068, n8069, n8070, n8071, n8072,
    n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084,
    n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102,
    n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114,
    n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126,
    n8127, n8128, n8129, n8130, n8131, n8132,
    n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144,
    n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156,
    n8157, n8158, n8159, n8160, n8161, n8162,
    n8163, n8164, n8165, n8166, n8167, n8168,
    n8169, n8170, n8171, n8172, n8173, n8174,
    n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186,
    n8187, n8188, n8189, n8190, n8191, n8192,
    n8193, n8194, n8195, n8196, n8197, n8198,
    n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8219, n8220, n8221, n8222,
    n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246,
    n8247, n8248, n8249, n8250, n8251, n8252,
    n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8278, n8279, n8280, n8281, n8282,
    n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8290, n8291, n8292, n8293, n8294,
    n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306,
    n8307, n8308, n8309, n8310, n8311, n8312,
    n8313, n8314, n8315, n8316, n8317, n8318,
    n8319, n8320, n8321, n8322, n8323, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336,
    n8337, n8338, n8339, n8340, n8341, n8342,
    n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366,
    n8367, n8368, n8369, n8370, n8371, n8372,
    n8373, n8374, n8375, n8376, n8377, n8378,
    n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396,
    n8397, n8398, n8399, n8400, n8401, n8402,
    n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456,
    n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486,
    n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564,
    n8565, n8566, n8567, n8568, n8569, n8570,
    n8571, n8572, n8573, n8574, n8575, n8576,
    n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8593, n8594,
    n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606,
    n8607, n8608, n8609, n8610, n8611, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618,
    n8619, n8620, n8621, n8622, n8623, n8624,
    n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648,
    n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678,
    n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708,
    n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726,
    n8727, n8728, n8729, n8730, n8731, n8732,
    n8733, n8734, n8735, n8736, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756,
    n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768,
    n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786,
    n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816,
    n8817, n8818, n8819, n8820, n8821, n8822,
    n8823, n8824, n8825, n8826, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8834,
    n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846,
    n8847, n8848, n8849, n8850, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864,
    n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876,
    n8877, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888,
    n8889, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8902, n8903, n8904, n8905, n8906,
    n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936,
    n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966,
    n8967, n8968, n8969, n8970, n8971, n8972,
    n8973, n8974, n8975, n8976, n8977, n8978,
    n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n8993, n8994, n8995, n8996,
    n8997, n8998, n8999, n9000, n9001, n9002,
    n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9026,
    n9027, n9028, n9029, n9030, n9031, n9032,
    n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050,
    n9051, n9052, n9053, n9054, n9055, n9056,
    n9057, n9058, n9059, n9060, n9061, n9062,
    n9063, n9064, n9065, n9066, n9067, n9068,
    n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9080,
    n9081, n9082, n9083, n9084, n9085, n9086,
    n9087, n9088, n9089, n9090, n9091, n9092,
    n9093, n9094, n9095, n9096, n9097, n9098,
    n9099, n9100, n9101, n9102, n9103, n9104,
    n9105, n9106, n9107, n9108, n9109, n9110,
    n9111, n9112, n9113, n9114, n9115, n9116,
    n9117, n9118, n9119, n9120, n9121, n9122,
    n9123, n9124, n9125, n9126, n9127, n9128,
    n9129, n9130, n9131, n9132, n9133, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140,
    n9141, n9142, n9143, n9144, n9145, n9146,
    n9147, n9148, n9149, n9150, n9151, n9152,
    n9153, n9154, n9155, n9156, n9157, n9158,
    n9159, n9160, n9161, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170,
    n9171, n9172, n9173, n9174, n9175, n9176,
    n9177, n9178, n9179, n9180, n9181, n9182,
    n9183, n9184, n9185, n9186, n9187, n9188,
    n9189, n9190, n9191, n9192, n9193, n9194,
    n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206,
    n9207, n9208, n9209, n9210, n9211, n9212,
    n9213, n9214, n9215, n9216, n9217, n9218,
    n9219, n9220, n9221, n9222, n9223, n9224,
    n9225, n9226, n9227, n9228, n9229, n9230,
    n9231, n9232, n9233, n9234, n9235, n9236,
    n9237, n9238, n9239, n9240, n9241, n9242,
    n9243, n9244, n9245, n9246, n9247, n9248,
    n9249, n9250, n9251, n9252, n9253, n9254,
    n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266,
    n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296,
    n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326,
    n9327, n9328, n9329, n9330, n9331, n9332,
    n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386,
    n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416,
    n9417, n9418, n9419, n9420, n9421, n9422,
    n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446,
    n9447, n9448, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052,
    n10053, n10054, n10055, n10056, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064,
    n10065, n10066, n10067, n10068, n10069, n10070,
    n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10082,
    n10083, n10084, n10085, n10086, n10087, n10088,
    n10089, n10090, n10091, n10092, n10093, n10094,
    n10095, n10096, n10097, n10098, n10099, n10100,
    n10101, n10102, n10103, n10104, n10105, n10106,
    n10107, n10108, n10109, n10110, n10111, n10112,
    n10113, n10114, n10115, n10116, n10117, n10118,
    n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10128, n10129, n10130,
    n10131, n10132, n10133, n10134, n10135, n10136,
    n10137, n10138, n10139, n10140, n10141, n10142,
    n10143, n10144, n10145, n10146, n10147, n10148,
    n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10158, n10159, n10160,
    n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10169, n10170, n10171, n10172,
    n10173, n10174, n10175, n10176, n10177, n10178,
    n10179, n10180, n10181, n10182, n10183, n10184,
    n10185, n10186, n10187, n10188, n10189, n10190,
    n10191, n10192, n10193, n10194, n10195, n10196,
    n10197, n10198, n10199, n10200, n10201, n10202,
    n10203, n10204, n10205, n10206, n10207, n10208,
    n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10222, n10223, n10224, n10225, n10226,
    n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238,
    n10239, n10240, n10241, n10242, n10243, n10244,
    n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256,
    n10257, n10258, n10259, n10260, n10261, n10262,
    n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292,
    n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328,
    n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10370,
    n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382,
    n10383, n10384, n10385, n10386, n10387, n10388,
    n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406,
    n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424,
    n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442,
    n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460,
    n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472,
    n10473, n10474, n10475, n10476, n10477, n10478,
    n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490,
    n10491, n10492, n10493, n10494, n10495, n10496,
    n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514,
    n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532,
    n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10546, n10547, n10548, n10549, n10550,
    n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562,
    n10563, n10564, n10565, n10566, n10567, n10568,
    n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580,
    n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598,
    n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10651, n10652,
    n10653, n10654, n10655, n10656, n10657, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664,
    n10665, n10666, n10667, n10668, n10669, n10670,
    n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706,
    n10707, n10708, n10709, n10710, n10711, n10712,
    n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724,
    n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742,
    n10743, n10744, n10745, n10746, n10747, n10748,
    n10749, n10750, n10751, n10752, n10753, n10754,
    n10755, n10756, n10757, n10758, n10759, n10760,
    n10761, n10762, n10763, n10764, n10765, n10766,
    n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778,
    n10779, n10780, n10781, n10782, n10783, n10784,
    n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868,
    n10869, n10870, n10871, n10872, n10873, n10874,
    n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892,
    n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904,
    n10905, n10906, n10907, n10908, n10909, n10910,
    n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922,
    n10923, n10924, n10925, n10926, n10927, n10928,
    n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940,
    n10941, n10942, n10943, n10944, n10945, n10946,
    n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054,
    n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066,
    n11067, n11068, n11069, n11070, n11071, n11072,
    n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084,
    n11085, n11086, n11087, n11088, n11089, n11090,
    n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108,
    n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126,
    n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144,
    n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156,
    n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174,
    n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11189, n11190, n11191, n11192,
    n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204,
    n11205, n11206, n11207, n11208, n11209, n11210,
    n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222,
    n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11242, n11243, n11244, n11245, n11246,
    n11247, n11248, n11249, n11250, n11251, n11252,
    n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264,
    n11265, n11266, n11267, n11268, n11269, n11270,
    n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282,
    n11283, n11284, n11285, n11286, n11287, n11288,
    n11289, n11290, n11291, n11292, n11293, n11294,
    n11295, n11296, n11297, n11298, n11299, n11300,
    n11301, n11302, n11303, n11304, n11305, n11306,
    n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318,
    n11319, n11320, n11321, n11322, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336,
    n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354,
    n11355, n11356, n11357, n11358, n11359, n11360,
    n11361, n11362, n11363, n11364, n11365, n11366,
    n11367, n11368, n11369, n11370, n11371, n11372,
    n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11394, n11395, n11396,
    n11397, n11398, n11399, n11400, n11401, n11402,
    n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414,
    n11415, n11416, n11417, n11418, n11419, n11420,
    n11421, n11422, n11423, n11424, n11425, n11426,
    n11427, n11428, n11429, n11430, n11431, n11432,
    n11433, n11434, n11435, n11436, n11437, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444,
    n11445, n11446, n11447, n11448, n11449, n11450,
    n11451, n11452, n11453, n11454, n11455, n11456,
    n11457, n11458, n11459, n11460, n11461, n11462,
    n11463, n11464, n11465, n11466, n11467, n11468,
    n11469, n11470, n11471, n11472, n11473, n11474,
    n11475, n11476, n11477, n11478, n11479, n11480,
    n11481, n11482, n11483, n11484, n11485, n11486,
    n11487, n11488, n11489, n11490, n11491, n11492,
    n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504,
    n11505, n11506, n11507, n11508, n11509, n11510,
    n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11520, n11521, n11522,
    n11523, n11524, n11525, n11526, n11527, n11528,
    n11529, n11530, n11531, n11532, n11533, n11534,
    n11535, n11536, n11537, n11538, n11539, n11540,
    n11541, n11542, n11543, n11544, n11545, n11546,
    n11547, n11548, n11549, n11550, n11551, n11552,
    n11553, n11554, n11555, n11556, n11557, n11558,
    n11559, n11560, n11561, n11562, n11563, n11564,
    n11565, n11566, n11567, n11568, n11569, n11570,
    n11571, n11572, n11573, n11574, n11575, n11576,
    n11577, n11578, n11579, n11580, n11581, n11582,
    n11583, n11584, n11585, n11586, n11587, n11588,
    n11589, n11590, n11591, n11592, n11593, n11594,
    n11595, n11596, n11597, n11598, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618,
    n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630,
    n11631, n11632, n11633, n11634, n11635, n11636,
    n11637, n11638, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11648,
    n11649, n11650, n11651, n11652, n11653, n11654,
    n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666,
    n11667, n11668, n11669, n11670, n11671, n11672,
    n11673, n11674, n11675, n11676, n11677, n11678,
    n11679, n11680, n11681, n11682, n11683, n11684,
    n11685, n11686, n11687, n11688, n11689, n11690,
    n11691, n11692, n11693, n11694, n11695, n11696,
    n11697, n11698, n11699, n11700, n11701, n11702,
    n11703, n11704, n11705, n11706, n11707, n11708,
    n11709, n11710, n11711, n11712, n11713, n11714,
    n11715, n11716, n11717, n11718, n11719, n11720,
    n11721, n11722, n11723, n11724, n11725, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756,
    n11757, n11758, n11759, n11760, n11761, n11762,
    n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774,
    n11775, n11776, n11777, n11778, n11779, n11780,
    n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792,
    n11793, n11794, n11795, n11796, n11797, n11798,
    n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810,
    n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218,
    n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236,
    n12237, n12238, n12239, n12240, n12241, n12242,
    n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254,
    n12255, n12256, n12257, n12258, n12259, n12260,
    n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272,
    n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290,
    n12291, n12292, n12293, n12294, n12295, n12296,
    n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314,
    n12315, n12316, n12317, n12318, n12319, n12320,
    n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12340, n12341, n12342, n12343, n12344,
    n12345, n12346, n12347, n12348, n12349, n12350,
    n12351, n12352, n12353, n12354, n12355, n12356,
    n12357, n12358, n12359, n12360, n12361, n12362,
    n12363, n12364, n12365, n12366, n12367, n12368,
    n12369, n12370, n12371, n12372, n12373, n12374,
    n12375, n12376, n12377, n12378, n12379, n12380,
    n12381, n12382, n12383, n12384, n12385, n12386,
    n12387, n12388, n12389, n12390, n12391, n12392,
    n12393, n12394, n12395, n12396, n12397, n12398,
    n12399, n12400, n12401, n12402, n12403, n12404,
    n12405, n12406, n12407, n12408, n12409, n12410,
    n12411, n12412, n12413, n12414, n12415, n12416,
    n12417, n12418, n12419, n12420, n12421, n12422,
    n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434,
    n12435, n12436, n12437, n12438, n12439, n12440,
    n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452,
    n12453, n12454, n12455, n12456, n12457, n12458,
    n12459, n12460, n12461, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470,
    n12471, n12472, n12473, n12474, n12475, n12476,
    n12477, n12478, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488,
    n12489, n12490, n12491, n12492, n12493, n12494,
    n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506,
    n12507, n12508, n12509, n12510, n12511, n12512,
    n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524,
    n12525, n12526, n12527, n12528, n12529, n12530,
    n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542,
    n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560,
    n12561, n12562, n12563, n12564, n12565, n12566,
    n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578,
    n12579, n12580, n12581, n12582, n12583, n12584,
    n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596,
    n12597, n12598, n12599, n12600, n12601, n12602,
    n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614,
    n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632,
    n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650,
    n12651, n12652, n12653, n12654, n12655, n12656,
    n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668,
    n12669, n12670, n12671, n12672, n12673, n12674,
    n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12691, n12692,
    n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704,
    n12705, n12706, n12707, n12708, n12709, n12710,
    n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722,
    n12723, n12724, n12725, n12726, n12727, n12728,
    n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740,
    n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758,
    n12759, n12760, n12761, n12762, n12763, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776,
    n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794,
    n12795, n12796, n12797, n12798, n12799, n12800,
    n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812,
    n12813, n12814, n12815, n12816, n12817, n12818,
    n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12830,
    n12831, n12832, n12833, n12834, n12835, n12836,
    n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848,
    n12849, n12850, n12851, n12852, n12853, n12854,
    n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866,
    n12867, n12868, n12869, n12870, n12871, n12872,
    n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884,
    n12885, n12886, n12887, n12888, n12889, n12890,
    n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902,
    n12903, n12904, n12905, n12906, n12907, n12908,
    n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920,
    n12921, n12922, n12923, n12924, n12925, n12926,
    n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938,
    n12939, n12940, n12941, n12942, n12943, n12944,
    n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956,
    n12957, n12958, n12959, n12960, n12961, n12962,
    n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974,
    n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010,
    n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028,
    n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046,
    n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058,
    n13059, n13060, n13061, n13062, n13063, n13064,
    n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13073, n13074, n13075, n13076,
    n13077, n13078, n13079, n13080, n13081, n13082,
    n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100,
    n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112,
    n13113, n13114, n13115, n13116, n13117, n13118,
    n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130,
    n13131, n13132, n13133, n13134, n13135, n13136,
    n13137, n13138, n13139, n13140, n13141, n13142,
    n13143, n13144, n13145, n13146, n13147, n13148,
    n13149, n13150, n13151, n13152, n13153, n13154,
    n13155, n13156, n13157, n13158, n13159, n13160,
    n13161, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232,
    n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322,
    n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13354, n13355, n13356, n13357, n13358,
    n13359, n13360, n13361, n13362, n13363, n13364,
    n13365, n13366, n13367, n13368, n13369, n13370,
    n13371, n13372, n13373, n13374, n13375, n13376,
    n13377, n13378, n13379, n13380, n13381, n13382,
    n13383, n13384, n13385, n13386, n13387, n13388,
    n13389, n13390, n13391, n13392, n13393, n13394,
    n13395, n13396, n13397, n13398, n13399, n13400,
    n13401, n13402, n13403, n13404, n13405, n13406,
    n13407, n13408, n13409, n13410, n13411, n13412,
    n13413, n13414, n13415, n13416, n13417, n13418,
    n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430,
    n13431, n13432, n13433, n13434, n13435, n13436,
    n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448,
    n13449, n13450, n13451, n13452, n13453, n13454,
    n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13464, n13465, n13466,
    n13467, n13468, n13469, n13470, n13471, n13472,
    n13473, n13474, n13475, n13476, n13477, n13478,
    n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13486, n13487, n13488, n13489, n13490,
    n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502,
    n13503, n13504, n13505, n13506, n13507, n13508,
    n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13516, n13517, n13518, n13519, n13520,
    n13521, n13522, n13523, n13524, n13525, n13526,
    n13527, n13528, n13529, n13530, n13531, n13532,
    n13533, n13534, n13535, n13536, n13537, n13538,
    n13539, n13540, n13541, n13542, n13543, n13544,
    n13545, n13546, n13547, n13548, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562,
    n13563, n13564, n13565, n13566, n13567, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580,
    n13581, n13582, n13583, n13584, n13585, n13586,
    n13587, n13588, n13589, n13590, n13591, n13592,
    n13593, n13594, n13595, n13596, n13597, n13598,
    n13599, n13600, n13601, n13602, n13603, n13604,
    n13605, n13606, n13607, n13608, n13609, n13610,
    n13611, n13612, n13613, n13614, n13615, n13616,
    n13617, n13618, n13619, n13620, n13621, n13622,
    n13623, n13624, n13625, n13626, n13627, n13628,
    n13629, n13630, n13631, n13632, n13633, n13634,
    n13635, n13636, n13637, n13638, n13639, n13640,
    n13641, n13642, n13643, n13644, n13645, n13646,
    n13647, n13648, n13649, n13650, n13651, n13652,
    n13653, n13654, n13655, n13656, n13657, n13658,
    n13659, n13660, n13661, n13662, n13663, n13664,
    n13665, n13666, n13667, n13668, n13669, n13670,
    n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682,
    n13683, n13684, n13685, n13686, n13687, n13688,
    n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700,
    n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718,
    n13719, n13720, n13721, n13722, n13723, n13724,
    n13725, n13726, n13727, n13728, n13729, n13730,
    n13731, n13732, n13733, n13734, n13735, n13736,
    n13737, n13738, n13739, n13740, n13741, n13742,
    n13743, n13744, n13745, n13746, n13747, n13748,
    n13749, n13750, n13751, n13752, n13753, n13754,
    n13755, n13756, n13757, n13758, n13759, n13760,
    n13761, n13762, n13763, n13764, n13765, n13766,
    n13767, n13768, n13769, n13770, n13771, n13772,
    n13773, n13774, n13775, n13776, n13777, n13778,
    n13779, n13780, n13781, n13782, n13783, n13784,
    n13785, n13786, n13787, n13788, n13789, n13790,
    n13791, n13792, n13793, n13794, n13795, n13796,
    n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808,
    n13809, n13810, n13811, n13812, n13813, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826,
    n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844,
    n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862,
    n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880,
    n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898,
    n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916,
    n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934,
    n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952,
    n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970,
    n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988,
    n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006,
    n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060,
    n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078,
    n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144,
    n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330,
    n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348,
    n14349, n14350, n14351, n14352, n14353, n14354,
    n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372,
    n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14381, n14382, n14383, n14384,
    n14385, n14386, n14387, n14388, n14389, n14390,
    n14391, n14392, n14393, n14394, n14395, n14396,
    n14397, n14398, n14399, n14400, n14401, n14402,
    n14403, n14404, n14405, n14406, n14407, n14408,
    n14409, n14410, n14411, n14412, n14413, n14414,
    n14415, n14416, n14417, n14418, n14419, n14420,
    n14421, n14422, n14423, n14424, n14425, n14426,
    n14427, n14428, n14429, n14430, n14431, n14432,
    n14433, n14434, n14435, n14436, n14437, n14438,
    n14439, n14440, n14441, n14442, n14443, n14444,
    n14445, n14446, n14447, n14448, n14449, n14450,
    n14451, n14452, n14453, n14454, n14455, n14456,
    n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468,
    n14469, n14470, n14471, n14472, n14473, n14474,
    n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486,
    n14487, n14488, n14489, n14490, n14491, n14492,
    n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504,
    n14505, n14506, n14507, n14508, n14509, n14510,
    n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522,
    n14523, n14524, n14525, n14526, n14527, n14528,
    n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540,
    n14541, n14542, n14543, n14544, n14545, n14546,
    n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558,
    n14559, n14560, n14561, n14562, n14563, n14564,
    n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576,
    n14577, n14578, n14579, n14580, n14581, n14582,
    n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594,
    n14595, n14596, n14597, n14598, n14599, n14600,
    n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612,
    n14613, n14614, n14615, n14616, n14617, n14618,
    n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630,
    n14631, n14632, n14633, n14634, n14635, n14636,
    n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648,
    n14649, n14650, n14651, n14652, n14653, n14654,
    n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666,
    n14667, n14668, n14669, n14670, n14671, n14672,
    n14673, n14674, n14675, n14676, n14677, n14678,
    n14679, n14680, n14681, n14682, n14683, n14684,
    n14685, n14686, n14687, n14688, n14689, n14690,
    n14691, n14692, n14693, n14694, n14695, n14696,
    n14697, n14698, n14699, n14700, n14701, n14702,
    n14703, n14704, n14705, n14706, n14707, n14708,
    n14709, n14710, n14711, n14712, n14713, n14714,
    n14715, n14716, n14717, n14718, n14719, n14720,
    n14721, n14722, n14723, n14724, n14725, n14726,
    n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738,
    n14739, n14740, n14741, n14742, n14743, n14744,
    n14745, n14746, n14747, n14748, n14749, n14750,
    n14751, n14752, n14753, n14754, n14755, n14756,
    n14757, n14758, n14759, n14760, n14761, n14762,
    n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816,
    n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834,
    n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846,
    n14847, n14848, n14849, n14850, n14851, n14852,
    n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864,
    n14865, n14866, n14867, n14868, n14869, n14870,
    n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882,
    n14883, n14884, n14885, n14886, n14887, n14888,
    n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906,
    n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924,
    n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942,
    n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978,
    n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996,
    n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014,
    n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032,
    n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050,
    n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068,
    n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086,
    n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122,
    n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194,
    n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230,
    n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248,
    n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15281, n15282, n15283, n15284,
    n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302,
    n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314,
    n15315, n15316, n15317, n15318, n15319, n15320,
    n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338,
    n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15355, n15356,
    n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368,
    n15369, n15370, n15371, n15372, n15373, n15374,
    n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392,
    n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404,
    n15405, n15406, n15407, n15408, n15409, n15410,
    n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422,
    n15423, n15424, n15425, n15426, n15427, n15428,
    n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440,
    n15441, n15442, n15443, n15444, n15445, n15446,
    n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458,
    n15459, n15460, n15461, n15462, n15463, n15464,
    n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476,
    n15477, n15478, n15479, n15480, n15481, n15482,
    n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494,
    n15495, n15496, n15497, n15498, n15499, n15500,
    n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512,
    n15513, n15514, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530,
    n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15768, n15769, n15770,
    n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782,
    n15783, n15784, n15785, n15786, n15787, n15788,
    n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800,
    n15801, n15802, n15803, n15804, n15805, n15806,
    n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824,
    n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854,
    n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872,
    n15873, n15874, n15875, n15876, n15877, n15878,
    n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890,
    n15891, n15892, n15893, n15894, n15895, n15896,
    n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908,
    n15909, n15910, n15911, n15912, n15913, n15914,
    n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926,
    n15927, n15928, n15929, n15930, n15931, n15932,
    n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944,
    n15945, n15946, n15947, n15948, n15949, n15950,
    n15951, n15952, n15953, n15954, n15955, n15956,
    n15957, n15958, n15959, n15960, n15961, n15962,
    n15963, n15964, n15965, n15966, n15967, n15968,
    n15969, n15970, n15971, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980,
    n15981, n15982, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998,
    n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016,
    n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034,
    n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106,
    n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178,
    n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196,
    n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214,
    n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232,
    n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250,
    n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262,
    n16263, n16264, n16265, n16266, n16267, n16268,
    n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280,
    n16281, n16282, n16283, n16284, n16285, n16286,
    n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16302, n16303, n16304,
    n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316,
    n16317, n16318, n16319, n16320, n16321, n16322,
    n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334,
    n16335, n16336, n16337, n16338, n16339, n16340,
    n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352,
    n16353, n16354, n16355, n16356, n16357, n16358,
    n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370,
    n16371, n16372, n16373, n16374, n16375, n16376,
    n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388,
    n16389, n16390, n16391, n16392, n16393, n16394,
    n16395, n16396, n16397, n16398, n16399, n16400,
    n16401, n16402, n16403, n16404, n16405, n16406,
    n16407, n16408, n16409, n16410, n16411, n16412,
    n16413, n16414, n16415, n16416, n16417, n16418,
    n16419, n16420, n16421, n16422, n16423, n16424,
    n16425, n16426, n16427, n16428, n16429, n16430,
    n16431, n16432, n16433, n16434, n16435, n16436,
    n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448,
    n16449, n16450, n16451, n16452, n16453, n16454,
    n16455, n16456, n16457, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466,
    n16467, n16468, n16469, n16470, n16471, n16472,
    n16473, n16474, n16475, n16476, n16477, n16478,
    n16479, n16480, n16481, n16482, n16483, n16484,
    n16485, n16486, n16487, n16488, n16489, n16490,
    n16491, n16492, n16493, n16494, n16495, n16496,
    n16497, n16498, n16499, n16500, n16501, n16502,
    n16503, n16504, n16505, n16506, n16507, n16508,
    n16509, n16510, n16511, n16512, n16513, n16514,
    n16515, n16516, n16517, n16518, n16519, n16520,
    n16521, n16522, n16523, n16524, n16525, n16526,
    n16527, n16528, n16529, n16530, n16531, n16532,
    n16533, n16534, n16535, n16536, n16537, n16538,
    n16539, n16540, n16541, n16542, n16543, n16544,
    n16545, n16546, n16547, n16548, n16549, n16550,
    n16551, n16552, n16553, n16554, n16555, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562,
    n16563, n16564, n16565, n16566, n16567, n16568,
    n16569, n16570, n16571, n16572, n16573, n16574,
    n16575, n16576, n16577, n16578, n16579, n16580,
    n16581, n16582, n16583, n16584, n16585, n16586,
    n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598,
    n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652,
    n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670,
    n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16687, n16688,
    n16689, n16690, n16691, n16692, n16693, n16694,
    n16695, n16696, n16697, n16698, n16699, n16700,
    n16701, n16702, n16703, n16704, n16705, n16706,
    n16707, n16708, n16709, n16710, n16711, n16712,
    n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724,
    n16725, n16726, n16727, n16728, n16729, n16730,
    n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742,
    n16743, n16744, n16745, n16746, n16747, n16748,
    n16749, n16750, n16751, n16752, n16753, n16754,
    n16755, n16756, n16757, n16758, n16759, n16760,
    n16761, n16762, n16763, n16764, n16765, n16766,
    n16767, n16768, n16769, n16770, n16771, n16772,
    n16773, n16774, n16775, n16776, n16777, n16778,
    n16779, n16780, n16781, n16782, n16783, n16784,
    n16785, n16786, n16787, n16788, n16789, n16790,
    n16791, n16792, n16793, n16794, n16795, n16796,
    n16797, n16798, n16799, n16800, n16801, n16802,
    n16803, n16804, n16805, n16806, n16807, n16808,
    n16809, n16810, n16811, n16812, n16813, n16814,
    n16815, n16816, n16817, n16818, n16819, n16820,
    n16821, n16822, n16823, n16824, n16825, n16826,
    n16827, n16828, n16829, n16830, n16831, n16832,
    n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844,
    n16845, n16846, n16847, n16848, n16849, n16850,
    n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16868,
    n16869, n16870, n16871, n16872, n16873, n16874,
    n16875, n16876, n16877, n16878, n16879, n16880,
    n16881, n16882, n16883, n16884, n16885, n16886,
    n16887, n16888, n16889, n16890, n16891, n16892,
    n16893, n16894, n16895, n16896, n16897, n16898,
    n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16906, n16907, n16908, n16909, n16910,
    n16911, n16912, n16913, n16914, n16915, n16916,
    n16917, n16918, n16919, n16920, n16921, n16922,
    n16923, n16924, n16925, n16926, n16927, n16928,
    n16929, n16930, n16931, n16932, n16933, n16934,
    n16935, n16936, n16937, n16938, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16952,
    n16953, n16954, n16955, n16956, n16957, n16958,
    n16959, n16960, n16961, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976,
    n16977, n16978, n16979, n16980, n16981, n16982,
    n16983, n16984, n16985, n16986, n16987, n16988,
    n16989, n16990, n16991, n16992, n16993, n16994,
    n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17004, n17005, n17006,
    n17007, n17008, n17009, n17010, n17011, n17012,
    n17013, n17014, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024,
    n17025, n17026, n17027, n17028, n17029, n17030,
    n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042,
    n17043, n17044, n17045, n17046, n17047, n17048,
    n17049, n17050, n17051, n17052, n17053, n17054,
    n17055, n17056, n17057, n17058, n17059, n17060,
    n17061, n17062, n17063, n17064, n17065, n17066,
    n17067, n17068, n17069, n17070, n17071, n17072,
    n17073, n17074, n17075, n17076, n17077, n17078,
    n17079, n17080, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090,
    n17091, n17092, n17093, n17094, n17095, n17096,
    n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17114,
    n17115, n17116, n17117, n17118, n17119, n17120,
    n17121, n17122, n17123, n17124, n17125, n17126,
    n17127, n17128, n17129, n17130, n17131, n17132,
    n17133, n17134, n17135, n17136, n17137, n17138,
    n17139, n17140, n17141, n17142, n17143, n17144,
    n17145, n17146, n17147, n17148, n17149, n17150,
    n17151, n17152, n17153, n17154, n17155, n17156,
    n17157, n17158, n17159, n17160, n17161, n17162,
    n17163, n17164, n17165, n17166, n17167, n17168,
    n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180,
    n17181, n17182, n17183, n17184, n17185, n17186,
    n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204,
    n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222,
    n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240,
    n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258,
    n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276,
    n17277, n17278, n17279, n17280, n17281, n17282,
    n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294,
    n17295, n17296, n17297, n17298, n17299, n17300,
    n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312,
    n17313, n17314, n17315, n17316, n17317, n17318,
    n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330,
    n17331, n17332, n17333, n17334, n17335, n17336,
    n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348,
    n17349, n17350, n17351, n17352, n17353, n17354,
    n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366,
    n17367, n17368, n17369, n17370, n17371, n17372,
    n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384,
    n17385, n17386, n17387, n17388, n17389, n17390,
    n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402,
    n17403, n17404, n17405, n17406, n17407, n17408,
    n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420,
    n17421, n17422, n17423, n17424, n17425, n17426,
    n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438,
    n17439, n17440, n17441, n17442, n17443, n17444,
    n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456,
    n17457, n17458, n17459, n17460, n17461, n17462,
    n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474,
    n17475, n17476, n17477, n17478, n17479, n17480,
    n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492,
    n17493, n17494, n17495, n17496, n17497, n17498,
    n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510,
    n17511, n17512, n17513, n17514, n17515, n17516,
    n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528,
    n17529, n17530, n17531, n17532, n17533, n17534,
    n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546,
    n17547, n17548, n17549, n17550, n17551, n17552,
    n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564,
    n17565, n17566, n17567, n17568, n17569, n17570,
    n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582,
    n17583, n17584, n17585, n17586, n17587, n17588,
    n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624,
    n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672,
    n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696,
    n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708,
    n17709, n17710, n17711, n17712, n17713, n17714,
    n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726,
    n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744,
    n17745, n17746, n17747, n17748, n17749, n17750,
    n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762,
    n17763, n17764, n17765, n17766, n17767, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780,
    n17781, n17782, n17783, n17784, n17785, n17786,
    n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798,
    n17799, n17800, n17801, n17802, n17803, n17804,
    n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816,
    n17817, n17818, n17819, n17820, n17821, n17822,
    n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834,
    n17835, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852,
    n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888,
    n17889, n17890, n17891, n17892, n17893, n17894,
    n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906,
    n17907, n17908, n17909, n17910, n17911, n17912,
    n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17923, n17924,
    n17925, n17926, n17927, n17928, n17929, n17930,
    n17931, n17932, n17933, n17934, n17935, n17936,
    n17937, n17938, n17939, n17940, n17941, n17942,
    n17943, n17944, n17945, n17946, n17947, n17948,
    n17949, n17950, n17951, n17952, n17953, n17954,
    n17955, n17956, n17957, n17958, n17959, n17960,
    n17961, n17962, n17963, n17964, n17965, n17966,
    n17967, n17968, n17969, n17970, n17971, n17972,
    n17973, n17974, n17975, n17976, n17977, n17978,
    n17979, n17980, n17981, n17982, n17983, n17984,
    n17985, n17986, n17987, n17988, n17989, n17990,
    n17991, n17992, n17993, n17994, n17995, n17996,
    n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014,
    n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032,
    n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050,
    n18051, n18052, n18053, n18054, n18055, n18056,
    n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068,
    n18069, n18070, n18071, n18072, n18073, n18074,
    n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086,
    n18087, n18088, n18089, n18090, n18091, n18092,
    n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104,
    n18105, n18106, n18107, n18108, n18109, n18110,
    n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122,
    n18123, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140,
    n18141, n18142, n18143, n18144, n18145, n18146,
    n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158,
    n18159, n18160, n18161, n18162, n18163, n18164,
    n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176,
    n18177, n18178, n18179, n18180, n18181, n18182,
    n18183, n18184, n18185, n18186, n18187, n18188,
    n18189, n18190, n18191, n18192, n18193, n18194,
    n18195, n18196, n18197, n18198, n18199, n18200,
    n18201, n18202, n18203, n18204, n18205, n18206,
    n18207, n18208, n18209, n18210, n18211, n18212,
    n18213, n18214, n18215, n18216, n18217, n18218,
    n18219, n18220, n18221, n18222, n18223, n18224,
    n18225, n18226, n18227, n18228, n18229, n18230,
    n18231, n18232, n18233, n18234, n18235, n18236,
    n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18248,
    n18249, n18250, n18251, n18252, n18253, n18254,
    n18255, n18256, n18257, n18258, n18259, n18260,
    n18261, n18262, n18263, n18264, n18265, n18266,
    n18267, n18268, n18269, n18270, n18271, n18272,
    n18273, n18274, n18275, n18276, n18277, n18278,
    n18279, n18280, n18281, n18282, n18283, n18284,
    n18285, n18286, n18287, n18288, n18289, n18290,
    n18291, n18292, n18293, n18294, n18295, n18296,
    n18297, n18298, n18299, n18300, n18301, n18302,
    n18303, n18304, n18305, n18306, n18307, n18308,
    n18309, n18310, n18311, n18312, n18313, n18314,
    n18315, n18316, n18317, n18318, n18319, n18320,
    n18321, n18322, n18323, n18324, n18325, n18326,
    n18327, n18328, n18329, n18330, n18331, n18332,
    n18333, n18334, n18335, n18336, n18337, n18338,
    n18339, n18340, n18341, n18342, n18343, n18344,
    n18345, n18346, n18347, n18348, n18349, n18350,
    n18351, n18352, n18353, n18354, n18355, n18356,
    n18357, n18358, n18359, n18360, n18361, n18362,
    n18363, n18364, n18365, n18366, n18367, n18368,
    n18369, n18370, n18371, n18372, n18373, n18374,
    n18375, n18376, n18377, n18378, n18379, n18380,
    n18381, n18382, n18383, n18384, n18385, n18386,
    n18387, n18388, n18389, n18390, n18391, n18392,
    n18393, n18394, n18395, n18396, n18397, n18398,
    n18399, n18400, n18401, n18402, n18403, n18404,
    n18405, n18406, n18407, n18408, n18409, n18410,
    n18411, n18412, n18413, n18414, n18415, n18416,
    n18417, n18418, n18419, n18420, n18421, n18422,
    n18423, n18424, n18425, n18426, n18427, n18428,
    n18429, n18430, n18431, n18432, n18433, n18434,
    n18435, n18436, n18437, n18438, n18439, n18440,
    n18441, n18442, n18443, n18444, n18445, n18446,
    n18447, n18448, n18449, n18450, n18451, n18452,
    n18453, n18454, n18455, n18456, n18457, n18458,
    n18459, n18460, n18461, n18462, n18463, n18464,
    n18465, n18466, n18467, n18468, n18469, n18470,
    n18471, n18472, n18473, n18474, n18475, n18476,
    n18477, n18478, n18479, n18480, n18481, n18482,
    n18483, n18484, n18485, n18486, n18487, n18488,
    n18489, n18490, n18491, n18492, n18493, n18494,
    n18495, n18496, n18497, n18498, n18499, n18500,
    n18501, n18502, n18503, n18504, n18505, n18506,
    n18507, n18508, n18509, n18510, n18511, n18512,
    n18513, n18514, n18515, n18516, n18517, n18518,
    n18519, n18520, n18521, n18522, n18523, n18524,
    n18525, n18526, n18527, n18528, n18529, n18530,
    n18531, n18532, n18533, n18534, n18535, n18536,
    n18537, n18538, n18539, n18540, n18541, n18542,
    n18543, n18544, n18545, n18546, n18547, n18548,
    n18549, n18550, n18551, n18552, n18553, n18554,
    n18555, n18556, n18557, n18558, n18559, n18560,
    n18561, n18562, n18563, n18564, n18565, n18566,
    n18567, n18568, n18569, n18570, n18571, n18572,
    n18573, n18574, n18575, n18576, n18577, n18578,
    n18579, n18580, n18581, n18582, n18583, n18584,
    n18585, n18586, n18587, n18588, n18589, n18590,
    n18591, n18592, n18593, n18594, n18595, n18596,
    n18597, n18598, n18599, n18600, n18601, n18602,
    n18603, n18604, n18605, n18606, n18607, n18608,
    n18609, n18610, n18611, n18612, n18613, n18614,
    n18615, n18616, n18617, n18618, n18619, n18620,
    n18621, n18622, n18623, n18624, n18625, n18626,
    n18627, n18628, n18629, n18630, n18631, n18632,
    n18633, n18634, n18635, n18636, n18637, n18638,
    n18639, n18640, n18641, n18642, n18643, n18644,
    n18645, n18646, n18647, n18648, n18649, n18650,
    n18651, n18652, n18653, n18654, n18655, n18656,
    n18657, n18658, n18659, n18660, n18661, n18662,
    n18663, n18664, n18665, n18666, n18667, n18668,
    n18669, n18670, n18671, n18672, n18673, n18674,
    n18675, n18676, n18677, n18678, n18679, n18680,
    n18681, n18682, n18683, n18684, n18685, n18686,
    n18687, n18688, n18689, n18690, n18691, n18692,
    n18693, n18694, n18695, n18696, n18697, n18698,
    n18699, n18700, n18701, n18702, n18703, n18704,
    n18705, n18706, n18707, n18708, n18709, n18710,
    n18711, n18712, n18713, n18714, n18715, n18716,
    n18717, n18718, n18719, n18720, n18721, n18722,
    n18723, n18724, n18725, n18726, n18727, n18728,
    n18729, n18730, n18731, n18732, n18733, n18734,
    n18735, n18736, n18737, n18738, n18739, n18740,
    n18741, n18742, n18743, n18744, n18745, n18746,
    n18747, n18748, n18749, n18750, n18751, n18752,
    n18753, n18754, n18755, n18756, n18757, n18758,
    n18759, n18760, n18761, n18762, n18763, n18764,
    n18765, n18766, n18767, n18768, n18769, n18770,
    n18771, n18772, n18773, n18774, n18775, n18776,
    n18777, n18778, n18779, n18780, n18781, n18782,
    n18783, n18784, n18785, n18786, n18787, n18788,
    n18789, n18790, n18791, n18792, n18793, n18794,
    n18795, n18796, n18797, n18798, n18799, n18800,
    n18801, n18802, n18803, n18804, n18805, n18806,
    n18807, n18808, n18809, n18810, n18811, n18812,
    n18813, n18814, n18815, n18816, n18817, n18818,
    n18819, n18820, n18821, n18822, n18823, n18824,
    n18825, n18826, n18827, n18828, n18829, n18830,
    n18831, n18832, n18833, n18834, n18835, n18836,
    n18837, n18838, n18839, n18840, n18841, n18842,
    n18843, n18844, n18845, n18846, n18847, n18848,
    n18849, n18850, n18851, n18852, n18853, n18854,
    n18855, n18856, n18857, n18858, n18859, n18860,
    n18861, n18862, n18863, n18864, n18865, n18866,
    n18867, n18868, n18869, n18870, n18871, n18872,
    n18873, n18874, n18875, n18876, n18877, n18878,
    n18879, n18880, n18881, n18882, n18883, n18884,
    n18885, n18886, n18887, n18888, n18889, n18890,
    n18891, n18892, n18893, n18894, n18895, n18896,
    n18897, n18898, n18899, n18900, n18901, n18902,
    n18903, n18904, n18905, n18906, n18907, n18908,
    n18909, n18910, n18911, n18912, n18913, n18914,
    n18915, n18916, n18917, n18918, n18919, n18920,
    n18921, n18922, n18923, n18924, n18925, n18926,
    n18927, n18928, n18929, n18930, n18931, n18932,
    n18933, n18934, n18935, n18936, n18937, n18938,
    n18939, n18940, n18941, n18942, n18943, n18944,
    n18945, n18946, n18947, n18948, n18949, n18950,
    n18951, n18952, n18953, n18954, n18955, n18956,
    n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968,
    n18969, n18970, n18971, n18972, n18973, n18974,
    n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986,
    n18987, n18988, n18989, n18990, n18991, n18992,
    n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004,
    n19005, n19006, n19007, n19008, n19009, n19010,
    n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022,
    n19023, n19024, n19025, n19026, n19027, n19028,
    n19029, n19030, n19031, n19032, n19033, n19034,
    n19035, n19036, n19037, n19038, n19039, n19040,
    n19041, n19042, n19043, n19044, n19045, n19046,
    n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058,
    n19059, n19060, n19061, n19062, n19063, n19064,
    n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076,
    n19077, n19078, n19079, n19080, n19081, n19082,
    n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094,
    n19095, n19096, n19097, n19098, n19099, n19100,
    n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112,
    n19113, n19114, n19115, n19116, n19117, n19118,
    n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130,
    n19131, n19132, n19133, n19134, n19135, n19136,
    n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148,
    n19149, n19150, n19151, n19152, n19153, n19154,
    n19155, n19156, n19157, n19158, n19159, n19160,
    n19161, n19162, n19163, n19164, n19165, n19166,
    n19167, n19168, n19169, n19170, n19171, n19172,
    n19173, n19174, n19175, n19176, n19177, n19178,
    n19179, n19180, n19181, n19182, n19183, n19184,
    n19185, n19186, n19187, n19188, n19189, n19190,
    n19191, n19192, n19193, n19194, n19195, n19196,
    n19197, n19198, n19199, n19200, n19201, n19202,
    n19203, n19204, n19205, n19206, n19207, n19208,
    n19209, n19210, n19211, n19212, n19213, n19214,
    n19215, n19216, n19217, n19218, n19219, n19220,
    n19221, n19222, n19223, n19224, n19225, n19226,
    n19227, n19228, n19229, n19230, n19231, n19232,
    n19233, n19234, n19235, n19236, n19237, n19238,
    n19239, n19240, n19241, n19242, n19243, n19244,
    n19245, n19246, n19247, n19248, n19249, n19250,
    n19251, n19252, n19253, n19254, n19255, n19256,
    n19257, n19258, n19259, n19260, n19261, n19262,
    n19263, n19264, n19265, n19266, n19267, n19268,
    n19269, n19270, n19271, n19272, n19273, n19274,
    n19275, n19276, n19277, n19278, n19279, n19280,
    n19281, n19282, n19283, n19284, n19285, n19286,
    n19287, n19288, n19289, n19290, n19291, n19292,
    n19293, n19294, n19295, n19296, n19297, n19298,
    n19299, n19300, n19301, n19302, n19303, n19304,
    n19305, n19306, n19307, n19308, n19309, n19310,
    n19311, n19312, n19313, n19314, n19315, n19316,
    n19317, n19318, n19319, n19320, n19321, n19322,
    n19323, n19324, n19325, n19326, n19327, n19328,
    n19329, n19330, n19331, n19332, n19333, n19334,
    n19335, n19336, n19337, n19338, n19339, n19340,
    n19341, n19342, n19343, n19344, n19345, n19346,
    n19347, n19348, n19349, n19350, n19351, n19352,
    n19353, n19354, n19355, n19356, n19357, n19358,
    n19359, n19360, n19361, n19362, n19363, n19364,
    n19365, n19366, n19367, n19368, n19369, n19370,
    n19371, n19372, n19373, n19374, n19375, n19376,
    n19377, n19378, n19379, n19380, n19381, n19382,
    n19383, n19384, n19385, n19386, n19387, n19388,
    n19389, n19390, n19391, n19392, n19393, n19394,
    n19395, n19396, n19397, n19398, n19399, n19400,
    n19401, n19402, n19403, n19404, n19405, n19406,
    n19407, n19408, n19409, n19410, n19411, n19412,
    n19413, n19414, n19415, n19416, n19417, n19418,
    n19419, n19420, n19421, n19422, n19423, n19424,
    n19425, n19426, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19435, n19436,
    n19437, n19438, n19439, n19440, n19441, n19442,
    n19443, n19444, n19445, n19446, n19447, n19448,
    n19449, n19450, n19451, n19452, n19453, n19454,
    n19455, n19456, n19457, n19458, n19459, n19460,
    n19461, n19462, n19463, n19464, n19465, n19466,
    n19467, n19468, n19469, n19470, n19471, n19472,
    n19473, n19474, n19475, n19476, n19477, n19478,
    n19479, n19480, n19481, n19482, n19483, n19484,
    n19485, n19486, n19487, n19488, n19489, n19490,
    n19491, n19492, n19493, n19494, n19495, n19496,
    n19497, n19498, n19499, n19500, n19501, n19502,
    n19503, n19504, n19505, n19506, n19507, n19508,
    n19509, n19510, n19511, n19512, n19513, n19514,
    n19515, n19516, n19517, n19518, n19519, n19520,
    n19521, n19522, n19523, n19524, n19525, n19526,
    n19527, n19528, n19529, n19530, n19531, n19532,
    n19533, n19534, n19535, n19536, n19537, n19538,
    n19539, n19540, n19541, n19542, n19543, n19544,
    n19545, n19546, n19547, n19548, n19549, n19550,
    n19551, n19552, n19553, n19554, n19555, n19556,
    n19557, n19558, n19559, n19560, n19561, n19562,
    n19563, n19564, n19565, n19566, n19567, n19568,
    n19569, n19570, n19571, n19572, n19573, n19574,
    n19575, n19576, n19577, n19578, n19579, n19580,
    n19581, n19582, n19583, n19584, n19585, n19586,
    n19587, n19588, n19589, n19590, n19591, n19592,
    n19593, n19594, n19595, n19596, n19597, n19598,
    n19599, n19600, n19601, n19602, n19603, n19604,
    n19605, n19606, n19607, n19608, n19609, n19610,
    n19611, n19612, n19613, n19614, n19615, n19616,
    n19617, n19618, n19619, n19620, n19621, n19622,
    n19623, n19624, n19625, n19626, n19627, n19628,
    n19629, n19630, n19631, n19632, n19633, n19634,
    n19635, n19636, n19637, n19638, n19639, n19640,
    n19641, n19642, n19643, n19644, n19645, n19646,
    n19647, n19648, n19649, n19650, n19651, n19652,
    n19653, n19654, n19655, n19656, n19657, n19658,
    n19659, n19660, n19661, n19662, n19663, n19664,
    n19665, n19666, n19667, n19668, n19669, n19670,
    n19671, n19672, n19673, n19674, n19675, n19676,
    n19677, n19678, n19679, n19680, n19681, n19682,
    n19683, n19684, n19685, n19686, n19687, n19688,
    n19689, n19690, n19691, n19692, n19693, n19694,
    n19695, n19696, n19697, n19698, n19699, n19700,
    n19701, n19702, n19703, n19704, n19705, n19706,
    n19707, n19708, n19709, n19710, n19711, n19712,
    n19713, n19714, n19715, n19716, n19717, n19718,
    n19719, n19720, n19721, n19722, n19723, n19724,
    n19725, n19726, n19727, n19728, n19729, n19730,
    n19731, n19732, n19733, n19734, n19735, n19736,
    n19737, n19738, n19739, n19740, n19741, n19742,
    n19743, n19744, n19745, n19746, n19747, n19748,
    n19749, n19750, n19751, n19752, n19753, n19754,
    n19755, n19756, n19757, n19758, n19759, n19760,
    n19761, n19762, n19763, n19764, n19765, n19766,
    n19767, n19768, n19769, n19770, n19771, n19772,
    n19773, n19774, n19775, n19776, n19777, n19778,
    n19779, n19780, n19781, n19782, n19783, n19784,
    n19785, n19786, n19787, n19788, n19789, n19790,
    n19791, n19792, n19793, n19794, n19795, n19796,
    n19797, n19798, n19799, n19800, n19801, n19802,
    n19803, n19804, n19805, n19806, n19807, n19808,
    n19809, n19810, n19811, n19812, n19813, n19814,
    n19815, n19816, n19817, n19818, n19819, n19820,
    n19821, n19822, n19823, n19824, n19825, n19826,
    n19827, n19828, n19829, n19830, n19831, n19832,
    n19833, n19834, n19835, n19836, n19837, n19838,
    n19839, n19840, n19841, n19842, n19843, n19844,
    n19845, n19846, n19847, n19848, n19849, n19850,
    n19851, n19852, n19853, n19854, n19855, n19856,
    n19857, n19858, n19859, n19860, n19861, n19862,
    n19863, n19864, n19865, n19866, n19867, n19868,
    n19869, n19870, n19871, n19872, n19873, n19874,
    n19875, n19876, n19877, n19878, n19879, n19880,
    n19881, n19882, n19883, n19884, n19885, n19886,
    n19887, n19888, n19889, n19890, n19891, n19892,
    n19893, n19894, n19895, n19896, n19897, n19898,
    n19899, n19900, n19901, n19902, n19903, n19904,
    n19905, n19906, n19907, n19908, n19909, n19910,
    n19911, n19912, n19913, n19914, n19915, n19916,
    n19917, n19918, n19919, n19920, n19921, n19922,
    n19923, n19924, n19925, n19926, n19927, n19928,
    n19929, n19930, n19931, n19932, n19933, n19934,
    n19935, n19936, n19937, n19938, n19939, n19940,
    n19941, n19942, n19943, n19944, n19945, n19946,
    n19947, n19948, n19949, n19950, n19951, n19952,
    n19953, n19954, n19955, n19956, n19957, n19958,
    n19959, n19960, n19961, n19962, n19963, n19964,
    n19965, n19966, n19967, n19968, n19969, n19970,
    n19971, n19972, n19973, n19974, n19975, n19976,
    n19977, n19978, n19979, n19980, n19981, n19982,
    n19983, n19984, n19985, n19986, n19987, n19988,
    n19989, n19990, n19991, n19992, n19993, n19994,
    n19995, n19996, n19997, n19998, n19999, n20000,
    n20001, n20002, n20003, n20004, n20005, n20006,
    n20007, n20008, n20009, n20010, n20011, n20012,
    n20013, n20014, n20015, n20016, n20017, n20018,
    n20019, n20020, n20021, n20022, n20023, n20024,
    n20025, n20026, n20027, n20028, n20029, n20030,
    n20031, n20032, n20033, n20034, n20035, n20036,
    n20037, n20038, n20039, n20040, n20041, n20042,
    n20043, n20044, n20045, n20046, n20047, n20048,
    n20049, n20050, n20051, n20052, n20053, n20054,
    n20055, n20056, n20057, n20058, n20059, n20060,
    n20061, n20062, n20063, n20064, n20065, n20066,
    n20067, n20068, n20069, n20070, n20071, n20072,
    n20073, n20074, n20075, n20076, n20077, n20078,
    n20079, n20080, n20081, n20082, n20083, n20084,
    n20085, n20086, n20087, n20088, n20089, n20090,
    n20091, n20092, n20093, n20094, n20095, n20096,
    n20097, n20098, n20099, n20100, n20101, n20102,
    n20103, n20104, n20105, n20106, n20107, n20108,
    n20109, n20110, n20111, n20112, n20113, n20114,
    n20115, n20116, n20117, n20118, n20119, n20120,
    n20121, n20122, n20123, n20124, n20125, n20126,
    n20127, n20128, n20129, n20130, n20131, n20132,
    n20133, n20134, n20135, n20136, n20137, n20138,
    n20139, n20140, n20141, n20142, n20143, n20144,
    n20145, n20146, n20147, n20148, n20149, n20150,
    n20151, n20152, n20153, n20154, n20155, n20156,
    n20157, n20158, n20159, n20160, n20161, n20162,
    n20163, n20164, n20165, n20166, n20167, n20168,
    n20169, n20170, n20171, n20172, n20173, n20174,
    n20175, n20176, n20177, n20178, n20179, n20180,
    n20181, n20182, n20183, n20184, n20185, n20186,
    n20187, n20188, n20189, n20190, n20191, n20192,
    n20193, n20194, n20195, n20196, n20197, n20198,
    n20199, n20200, n20201, n20202, n20203, n20204,
    n20205, n20206, n20207, n20208, n20209, n20210,
    n20211, n20212, n20213, n20214, n20215, n20216,
    n20217, n20218, n20219, n20220, n20221, n20222,
    n20223, n20224, n20225, n20226, n20227, n20228,
    n20229, n20230, n20231, n20232, n20233, n20234,
    n20235, n20236, n20237, n20238, n20239, n20240,
    n20241, n20242, n20243, n20244, n20245, n20246,
    n20247, n20248, n20249, n20250, n20251, n20252,
    n20253, n20254, n20255, n20256, n20257, n20258,
    n20259, n20260, n20261, n20262, n20263, n20264,
    n20265, n20266, n20267, n20268, n20269, n20270,
    n20271, n20272, n20273, n20274, n20275, n20276,
    n20277, n20278, n20279, n20280, n20281, n20282,
    n20283, n20284, n20285, n20286, n20287, n20288,
    n20289, n20290, n20291, n20292, n20293, n20294,
    n20295, n20296, n20297, n20298, n20299, n20300,
    n20301, n20302, n20303, n20304, n20305, n20306,
    n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318,
    n20319, n20320, n20321, n20322, n20323, n20324,
    n20325, n20326, n20327, n20328, n20329, n20330,
    n20331, n20332, n20333, n20334, n20335, n20336,
    n20337, n20338, n20339, n20340, n20341, n20342,
    n20343, n20344, n20345, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354,
    n20355, n20356, n20357, n20358, n20359, n20360,
    n20361, n20362, n20363, n20364, n20365, n20366,
    n20367, n20368, n20369, n20370, n20371, n20372,
    n20373, n20374, n20375, n20376, n20377, n20378,
    n20379, n20380, n20381, n20382, n20383, n20384,
    n20385, n20386, n20387, n20388, n20389, n20390,
    n20391, n20392, n20393, n20394, n20395, n20396,
    n20397, n20398, n20399, n20400, n20401, n20402,
    n20403, n20404, n20405, n20406, n20407, n20408,
    n20409, n20410, n20411, n20412, n20413, n20414,
    n20415, n20416, n20417, n20418, n20419, n20420,
    n20421, n20422, n20423, n20424, n20425, n20426,
    n20427, n20428, n20429, n20430, n20431, n20432,
    n20433, n20434, n20435, n20436, n20437, n20438,
    n20439, n20440, n20441, n20442, n20443, n20444,
    n20445, n20446, n20447, n20448, n20449, n20450,
    n20451, n20452, n20453, n20454, n20455, n20456,
    n20457, n20458, n20459, n20460, n20461, n20462,
    n20463, n20464, n20465, n20466, n20467, n20468,
    n20469, n20470, n20471, n20472, n20473, n20474,
    n20475, n20476, n20477, n20478, n20479, n20480,
    n20481, n20482, n20483, n20484, n20485, n20486,
    n20487, n20488, n20489, n20490, n20491, n20492,
    n20493, n20494, n20495, n20496, n20497, n20498,
    n20499, n20500, n20501, n20502, n20503, n20504,
    n20505, n20506, n20507, n20508, n20509, n20510,
    n20511, n20512, n20513, n20514, n20515, n20516,
    n20517, n20518, n20519, n20520, n20521, n20522,
    n20523, n20524, n20525, n20526, n20527, n20528,
    n20529, n20530, n20531, n20532, n20533, n20534,
    n20535, n20536, n20537, n20538, n20539, n20540,
    n20541, n20542, n20543, n20544, n20545, n20546,
    n20547, n20548, n20549, n20550, n20551, n20552,
    n20553, n20554, n20555, n20556, n20557, n20558,
    n20559, n20560, n20561, n20562, n20563, n20564,
    n20565, n20566, n20567, n20568, n20569, n20570,
    n20571, n20572, n20573, n20574, n20575, n20576,
    n20577, n20578, n20579, n20580, n20581, n20582,
    n20583, n20584, n20585, n20586, n20587, n20588,
    n20589, n20590, n20591, n20592, n20593, n20594,
    n20595, n20596, n20597, n20598, n20599, n20600,
    n20601, n20602, n20603, n20604, n20605, n20606,
    n20607, n20608, n20609, n20610, n20611, n20612,
    n20613, n20614, n20615, n20616, n20617, n20618,
    n20619, n20620, n20621, n20622, n20623, n20624,
    n20625, n20626, n20627, n20628, n20629, n20630,
    n20631, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20645, n20646, n20647, n20648,
    n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660,
    n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20675, n20676, n20677, n20678,
    n20679, n20680, n20681, n20682, n20683, n20684,
    n20685, n20686, n20687, n20688, n20689, n20690,
    n20691, n20692, n20693, n20694, n20695, n20696,
    n20697, n20698, n20699, n20700, n20701, n20702,
    n20703, n20704, n20705, n20706, n20707, n20708,
    n20709, n20710, n20711, n20712, n20713, n20714,
    n20715, n20716, n20717, n20718, n20719, n20720,
    n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732,
    n20733, n20734, n20735, n20736, n20737, n20738,
    n20739, n20740, n20741, n20742, n20743, n20744,
    n20745, n20746, n20747, n20748, n20749, n20750,
    n20751, n20752, n20753, n20754, n20755, n20756,
    n20757, n20758, n20759, n20760, n20761, n20762,
    n20763, n20764, n20765, n20766, n20767, n20768,
    n20769, n20770, n20771, n20772, n20773, n20774,
    n20775, n20776, n20777, n20778, n20779, n20780,
    n20781, n20782, n20783, n20784, n20785, n20786,
    n20787, n20788, n20789, n20790, n20791, n20792,
    n20793, n20794, n20795, n20796, n20797, n20798,
    n20799, n20800, n20801, n20802, n20803, n20804,
    n20805, n20806, n20807, n20808, n20809, n20810,
    n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822,
    n20823, n20824, n20825, n20826, n20827, n20828,
    n20829, n20830, n20831, n20832, n20833, n20834,
    n20835, n20836, n20837, n20838, n20839, n20840,
    n20841, n20842, n20843, n20844, n20845, n20846,
    n20847, n20848, n20849, n20850, n20851, n20852,
    n20853, n20854, n20855, n20856, n20857, n20858,
    n20859, n20860, n20861, n20862, n20863, n20864,
    n20865, n20866, n20867, n20868, n20869, n20870,
    n20871, n20872, n20873, n20874, n20875, n20876,
    n20877, n20878, n20879, n20880, n20881, n20882,
    n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20892, n20893, n20894,
    n20895, n20896, n20897, n20898, n20899, n20900,
    n20901, n20902, n20903, n20904, n20905, n20906,
    n20907, n20908, n20909, n20910, n20911, n20912,
    n20913, n20914, n20915, n20916, n20917, n20918,
    n20919, n20920, n20921, n20922, n20923, n20924,
    n20925, n20926, n20927, n20928, n20929, n20930,
    n20931, n20932, n20933, n20934, n20935, n20936,
    n20937, n20938, n20939, n20940, n20941, n20942,
    n20943, n20944, n20945, n20946, n20947, n20948,
    n20949, n20950, n20951, n20952, n20953, n20954,
    n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972,
    n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984,
    n20985, n20986, n20987, n20988, n20989, n20990,
    n20991, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008,
    n21009, n21010, n21011, n21012, n21013, n21014,
    n21015, n21016, n21017, n21018, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026,
    n21027, n21028, n21029, n21030, n21031, n21032,
    n21033, n21034, n21035, n21036, n21037, n21038,
    n21039, n21040, n21041, n21042, n21043, n21044,
    n21045, n21046, n21047, n21048, n21049, n21050,
    n21051, n21052, n21053, n21054, n21055, n21056,
    n21057, n21058, n21059, n21060, n21061, n21062,
    n21063, n21064, n21065, n21066, n21067, n21068,
    n21069, n21070, n21071, n21072, n21073, n21074,
    n21075, n21076, n21077, n21078, n21079, n21080,
    n21081, n21082, n21083, n21084, n21085, n21086,
    n21087, n21088, n21089, n21090, n21091, n21092,
    n21093, n21094, n21095, n21096, n21097, n21098,
    n21099, n21100, n21101, n21102, n21103, n21104,
    n21105, n21106, n21107, n21108, n21109, n21110,
    n21111, n21112, n21113, n21114, n21115, n21116,
    n21117, n21118, n21119, n21120, n21121, n21122,
    n21123, n21124, n21125, n21126, n21127, n21128,
    n21129, n21130, n21131, n21132, n21133, n21134,
    n21135, n21136, n21137, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21145, n21146,
    n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158,
    n21159, n21160, n21161, n21162, n21163, n21164,
    n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176,
    n21177, n21178, n21179, n21180, n21181, n21182,
    n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200,
    n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218,
    n21219, n21220, n21221, n21222, n21223, n21224,
    n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236,
    n21237, n21238, n21239, n21240, n21241, n21242,
    n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260,
    n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21278,
    n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290,
    n21291, n21292, n21293, n21294, n21295, n21296,
    n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314,
    n21315, n21316, n21317, n21318, n21319, n21320,
    n21321, n21322, n21323, n21324, n21325, n21326,
    n21327, n21328, n21329, n21330, n21331, n21332,
    n21333, n21334, n21335, n21336, n21337, n21338,
    n21339, n21340, n21341, n21342, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350,
    n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368,
    n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428,
    n21429, n21430, n21431, n21432, n21433, n21434,
    n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21446,
    n21447, n21448, n21449, n21450, n21451, n21452,
    n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464,
    n21465, n21466, n21467, n21468, n21469, n21470,
    n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482,
    n21483, n21484, n21485, n21486, n21487, n21488,
    n21489, n21490, n21491, n21492, n21493, n21494,
    n21495, n21496, n21497, n21498, n21499, n21500,
    n21501, n21502, n21503, n21504, n21505, n21506,
    n21507, n21508, n21509, n21510, n21511, n21512,
    n21513, n21514, n21515, n21516, n21517, n21518,
    n21519, n21520, n21521, n21522, n21523, n21524,
    n21525, n21526, n21527, n21528, n21529, n21530,
    n21531, n21532, n21533, n21534, n21535, n21536,
    n21537, n21538, n21539, n21540, n21541, n21542,
    n21543, n21544, n21545, n21546, n21547, n21548,
    n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560,
    n21561, n21562, n21563, n21564, n21565, n21566,
    n21567, n21568, n21569, n21570, n21571, n21572,
    n21573, n21574, n21575, n21576, n21577, n21578,
    n21579, n21580, n21581, n21582, n21583, n21584,
    n21585, n21586, n21587, n21588, n21589, n21590,
    n21591, n21592, n21593, n21594, n21595, n21596,
    n21597, n21598, n21599, n21600, n21601, n21602,
    n21603, n21604, n21605, n21606, n21607, n21608,
    n21609, n21610, n21611, n21612, n21613, n21614,
    n21615, n21616, n21617, n21618, n21619, n21620,
    n21621, n21622, n21623, n21624, n21625, n21626,
    n21627, n21628, n21629, n21630, n21631, n21632,
    n21633, n21634, n21635, n21636, n21637, n21638,
    n21639, n21640, n21641, n21642, n21643, n21644,
    n21645, n21646, n21647, n21648, n21649, n21650,
    n21651, n21652, n21653, n21654, n21655, n21656,
    n21657, n21658, n21659, n21660, n21661, n21662,
    n21663, n21664, n21665, n21666, n21667, n21668,
    n21669, n21670, n21671, n21672, n21673, n21674,
    n21675, n21676, n21677, n21678, n21679, n21680,
    n21681, n21682, n21683, n21684, n21685, n21686,
    n21687, n21688, n21689, n21690, n21691, n21692,
    n21693, n21694, n21695, n21696, n21697, n21698,
    n21699, n21700, n21701, n21702, n21703, n21704,
    n21705, n21706, n21707, n21708, n21709, n21710,
    n21711, n21712, n21713, n21714, n21715, n21716,
    n21717, n21718, n21719, n21720, n21721, n21722,
    n21723, n21724, n21725, n21726, n21727, n21728,
    n21729, n21730, n21731, n21732, n21733, n21734,
    n21735, n21736, n21737, n21738, n21739, n21740,
    n21741, n21742, n21743, n21744, n21745, n21746,
    n21747, n21748, n21749, n21750, n21751, n21752,
    n21753, n21754, n21755, n21756, n21757, n21758,
    n21759, n21760, n21761, n21762, n21763, n21764,
    n21765, n21766, n21767, n21768, n21769, n21770,
    n21771, n21772, n21773, n21774, n21775, n21776,
    n21777, n21778, n21779, n21780, n21781, n21782,
    n21783, n21784, n21785, n21786, n21787, n21788,
    n21789, n21790, n21791, n21792, n21793, n21794,
    n21795, n21796, n21797, n21798, n21799, n21800,
    n21801, n21802, n21803, n21804, n21805, n21806,
    n21807, n21808, n21809, n21810, n21811, n21812,
    n21813, n21814, n21815, n21816, n21817, n21818,
    n21819, n21820, n21821, n21822, n21823, n21824,
    n21825, n21826, n21827, n21828, n21829, n21830,
    n21831, n21832, n21833, n21834, n21835, n21836,
    n21837, n21838, n21839, n21840, n21841, n21842,
    n21843, n21844, n21845, n21846, n21847, n21848,
    n21849, n21850, n21851, n21852, n21853, n21854,
    n21855, n21856, n21857, n21858, n21859, n21860,
    n21861, n21862, n21863, n21864, n21865, n21866,
    n21867, n21868, n21869, n21870, n21871, n21872,
    n21873, n21874, n21875, n21876, n21877, n21878,
    n21879, n21880, n21881, n21882, n21883, n21884,
    n21885, n21886, n21887, n21888, n21889, n21890,
    n21891, n21892, n21893, n21894, n21895, n21896,
    n21897, n21898, n21899, n21900, n21901, n21902,
    n21903, n21904, n21905, n21906, n21907, n21908,
    n21909, n21910, n21911, n21912, n21913, n21914,
    n21915, n21916, n21917, n21918, n21919, n21920,
    n21921, n21922, n21923, n21924, n21925, n21926,
    n21927, n21928, n21929, n21930, n21931, n21932,
    n21933, n21934, n21935, n21936, n21937, n21938,
    n21939, n21940, n21941, n21942, n21943, n21944,
    n21945, n21946, n21947, n21948, n21949, n21950,
    n21951, n21952, n21953, n21954, n21955, n21956,
    n21957, n21958, n21959, n21960, n21961, n21962,
    n21963, n21964, n21965, n21966, n21967, n21968,
    n21969, n21970, n21971, n21972, n21973, n21974,
    n21975, n21976, n21977, n21978, n21979, n21980,
    n21981, n21982, n21983, n21984, n21985, n21986,
    n21987, n21988, n21989, n21990, n21991, n21992,
    n21993, n21994, n21995, n21996, n21997, n21998,
    n21999, n22000, n22001, n22002, n22003, n22004,
    n22005, n22006, n22007, n22008, n22009, n22010,
    n22011, n22012, n22013, n22014, n22015, n22016,
    n22017, n22018, n22019, n22020, n22021, n22022,
    n22023, n22024, n22025, n22026, n22027, n22028,
    n22029, n22030, n22031, n22032, n22033, n22034,
    n22035, n22036, n22037, n22038, n22039, n22040,
    n22041, n22042, n22043, n22044, n22045, n22046,
    n22047, n22048, n22049, n22050, n22051, n22052,
    n22053, n22054, n22055, n22056, n22057, n22058,
    n22059, n22060, n22061, n22062, n22063, n22064,
    n22065, n22066, n22067, n22068, n22069, n22070,
    n22071, n22072, n22073, n22074, n22075, n22076,
    n22077, n22078, n22079, n22080, n22081, n22082,
    n22083, n22084, n22085, n22086, n22087, n22088,
    n22089, n22090, n22091, n22092, n22093, n22094,
    n22095, n22096, n22097, n22098, n22099, n22100,
    n22101, n22102, n22103, n22104, n22105, n22106,
    n22107, n22108, n22109, n22110, n22111, n22112,
    n22113, n22114, n22115, n22116, n22117, n22118,
    n22119, n22120, n22121, n22122, n22123, n22124,
    n22125, n22126, n22127, n22128, n22129, n22130,
    n22131, n22132, n22133, n22134, n22135, n22136,
    n22137, n22138, n22139, n22140, n22141, n22142,
    n22143, n22144, n22145, n22146, n22147, n22148,
    n22149, n22150, n22151, n22152, n22153, n22154,
    n22155, n22156, n22157, n22158, n22159, n22160,
    n22161, n22162, n22163, n22164, n22165, n22166,
    n22167, n22168, n22169, n22170, n22171, n22172,
    n22173, n22174, n22175, n22176, n22177, n22178,
    n22179, n22180, n22181, n22182, n22183, n22184,
    n22185, n22186, n22187, n22188, n22189, n22190,
    n22191, n22192, n22193, n22194, n22195, n22196,
    n22197, n22198, n22199, n22200, n22201, n22202,
    n22203, n22204, n22205, n22206, n22207, n22208,
    n22209, n22210, n22211, n22212, n22213, n22214,
    n22215, n22216, n22217, n22218, n22219, n22220,
    n22221, n22222, n22223, n22224, n22225, n22226,
    n22227, n22228, n22229, n22230, n22231, n22232,
    n22233, n22234, n22235, n22236, n22237, n22238,
    n22239, n22240, n22241, n22242, n22243, n22244,
    n22245, n22246, n22247, n22248, n22249, n22250,
    n22251, n22252, n22253, n22254, n22255, n22256,
    n22257, n22258, n22259, n22260, n22261, n22262,
    n22263, n22264, n22265, n22266, n22267, n22268,
    n22269, n22270, n22271, n22272, n22273, n22274,
    n22275, n22276, n22277, n22278, n22279, n22280,
    n22281, n22282, n22283, n22284, n22285, n22286,
    n22287, n22288, n22289, n22290, n22291, n22292,
    n22293, n22294, n22295, n22296, n22297, n22298,
    n22299, n22300, n22301, n22302, n22303, n22304,
    n22305, n22306, n22307, n22308, n22309, n22310,
    n22311, n22312, n22313, n22314, n22315, n22316,
    n22317, n22318, n22319, n22320, n22321, n22322,
    n22323, n22324, n22325, n22326, n22327, n22328,
    n22329, n22330, n22331, n22332, n22333, n22334,
    n22335, n22336, n22337, n22338, n22339, n22340,
    n22341, n22342, n22343, n22344, n22345, n22346,
    n22347, n22348, n22349, n22350, n22351, n22352,
    n22353, n22354, n22355, n22356, n22357, n22358,
    n22359, n22360, n22361, n22362, n22363, n22364,
    n22365, n22366, n22367, n22368, n22369, n22370,
    n22371, n22372, n22373, n22374, n22375, n22376,
    n22377, n22378, n22379, n22380, n22381, n22382,
    n22383, n22384, n22385, n22386, n22387, n22388,
    n22389, n22390, n22391, n22392, n22393, n22394,
    n22395, n22396, n22397, n22398, n22399, n22400,
    n22401, n22402, n22403, n22404, n22405, n22406,
    n22407, n22408, n22409, n22410, n22411, n22412,
    n22413, n22414, n22415, n22416, n22417, n22418,
    n22419, n22420, n22421, n22422, n22423, n22424,
    n22425, n22426, n22427, n22428, n22429, n22430,
    n22431, n22432, n22433, n22434, n22435, n22436,
    n22437, n22438, n22439, n22440, n22441, n22442,
    n22443, n22444, n22445, n22446, n22447, n22448,
    n22449, n22450, n22451, n22452, n22453, n22454,
    n22455, n22456, n22457, n22458, n22459, n22460,
    n22461, n22462, n22463, n22464, n22465, n22466,
    n22467, n22468, n22469, n22470, n22471, n22472,
    n22473, n22474, n22475, n22476, n22477, n22478,
    n22479, n22480, n22481, n22482, n22483, n22484,
    n22485, n22486, n22487, n22488, n22489, n22490,
    n22491, n22492, n22493, n22494, n22495, n22496,
    n22497, n22498, n22499, n22500, n22501, n22502,
    n22503, n22504, n22505, n22506, n22507, n22508,
    n22509, n22510, n22511, n22512, n22513, n22514,
    n22515, n22516, n22517, n22518, n22519, n22520,
    n22521, n22522, n22523, n22524, n22525, n22526,
    n22527, n22528, n22529, n22530, n22531, n22532,
    n22533, n22534, n22535, n22536, n22537, n22538,
    n22539, n22540, n22541, n22542, n22543, n22544,
    n22545, n22546, n22547, n22548, n22549, n22550,
    n22551, n22552, n22553, n22554, n22555, n22556,
    n22557, n22558, n22559, n22560, n22561, n22562,
    n22563, n22564, n22565, n22566, n22567, n22568,
    n22569, n22570, n22571, n22572, n22573, n22574,
    n22575, n22576, n22577, n22578, n22579, n22580,
    n22581, n22582, n22583, n22584, n22585, n22586,
    n22587, n22588, n22589, n22590, n22591, n22592,
    n22593, n22594, n22595, n22596, n22597, n22598,
    n22599, n22600, n22601, n22602, n22603, n22604,
    n22605, n22606, n22607, n22608, n22609, n22610,
    n22611, n22612, n22613, n22614, n22615, n22616,
    n22617, n22618, n22619, n22620, n22621, n22622,
    n22623, n22624, n22625, n22626, n22627, n22628,
    n22629, n22630, n22631, n22632, n22633, n22634,
    n22635, n22636, n22637, n22638, n22639, n22640,
    n22641, n22642, n22643, n22644, n22645, n22646,
    n22647, n22648, n22649, n22650, n22651, n22652,
    n22653, n22654, n22655, n22656, n22657, n22658,
    n22659, n22660, n22661, n22662, n22663, n22664,
    n22665, n22666, n22667, n22668, n22669, n22670,
    n22671, n22672, n22673, n22674, n22675, n22676,
    n22677, n22678, n22679, n22680, n22681, n22682,
    n22683, n22684, n22685, n22686, n22687, n22688,
    n22689, n22690, n22691, n22692, n22693, n22694,
    n22695, n22696, n22697, n22698, n22699, n22700,
    n22701, n22702, n22703, n22704, n22705, n22706,
    n22707, n22708, n22709, n22710, n22711, n22712,
    n22713, n22714, n22715, n22716, n22717, n22718,
    n22719, n22720, n22721, n22722, n22723, n22724,
    n22725, n22726, n22727, n22728, n22729, n22730,
    n22731, n22732, n22733, n22734, n22735, n22736,
    n22737, n22738, n22739, n22740, n22741, n22742,
    n22743, n22744, n22745, n22746, n22747, n22748,
    n22749, n22750, n22751, n22752, n22753, n22754,
    n22755, n22756, n22757, n22758, n22759, n22760,
    n22761, n22762, n22763, n22764, n22765, n22766,
    n22767, n22768, n22769, n22770, n22771, n22772,
    n22773, n22774, n22775, n22776, n22777, n22778,
    n22779, n22780, n22781, n22782, n22783, n22784,
    n22785, n22786, n22787, n22788, n22789, n22790,
    n22791, n22792, n22793, n22794, n22795, n22796,
    n22797, n22798, n22799, n22800, n22801, n22802,
    n22803, n22804, n22805, n22806, n22807, n22808,
    n22809, n22810, n22811, n22812, n22813, n22814,
    n22815, n22816, n22817, n22818, n22819, n22820,
    n22821, n22822, n22823, n22824, n22825, n22826,
    n22827, n22828, n22829, n22830, n22831, n22832,
    n22833, n22834, n22835, n22836, n22837, n22838,
    n22839, n22840, n22841, n22842, n22843, n22844,
    n22845, n22846, n22847, n22848, n22849, n22850,
    n22851, n22852, n22853, n22854, n22855, n22856,
    n22857, n22858, n22859, n22860, n22861, n22862,
    n22863, n22864, n22865, n22866, n22867, n22868,
    n22869, n22870, n22871, n22872, n22873, n22874,
    n22875, n22876, n22877, n22878, n22879, n22880,
    n22881, n22882, n22883, n22884, n22885, n22886,
    n22887, n22888, n22889, n22890, n22891, n22892,
    n22893, n22894, n22895, n22896, n22897, n22898,
    n22899, n22900, n22901, n22902, n22903, n22904,
    n22905, n22906, n22907, n22908, n22909, n22910,
    n22911, n22912, n22913, n22914, n22915, n22916,
    n22917, n22918, n22919, n22920, n22921, n22922,
    n22923, n22924, n22925, n22926, n22927, n22928,
    n22929, n22930, n22931, n22932, n22933, n22934,
    n22935, n22936, n22937, n22938, n22939, n22940,
    n22941, n22942, n22943, n22944, n22945, n22946,
    n22947, n22948, n22949, n22950, n22951, n22952,
    n22953, n22954, n22955, n22956, n22957, n22958,
    n22959, n22960, n22961, n22962, n22963, n22964,
    n22965, n22966, n22967, n22968, n22969, n22970,
    n22971, n22972, n22973, n22974, n22975, n22976,
    n22977, n22978, n22979, n22980, n22981, n22982,
    n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994,
    n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012,
    n23013, n23014, n23015, n23016, n23017, n23018,
    n23019, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n23028, n23029, n23030,
    n23031, n23032, n23033, n23034, n23035, n23036,
    n23037, n23038, n23039, n23040, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048,
    n23049, n23050, n23051, n23052, n23053, n23054,
    n23055, n23056, n23057, n23058, n23059, n23060,
    n23061, n23062, n23063, n23064, n23065, n23066,
    n23067, n23068, n23069, n23070, n23071, n23072,
    n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084,
    n23085, n23086, n23087, n23088, n23089, n23090,
    n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102,
    n23103, n23104, n23105, n23106, n23107, n23108,
    n23109, n23110, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120,
    n23121, n23122, n23123, n23124, n23125, n23126,
    n23127, n23128, n23129, n23130, n23131, n23132,
    n23133, n23134, n23135, n23136, n23137, n23138,
    n23139, n23140, n23141, n23142, n23143, n23144,
    n23145, n23146, n23147, n23148, n23149, n23150,
    n23151, n23152, n23153, n23154, n23155, n23156,
    n23157, n23158, n23159, n23160, n23161, n23162,
    n23163, n23164, n23165, n23166, n23167, n23168,
    n23169, n23170, n23171, n23172, n23173, n23174,
    n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186,
    n23187, n23188, n23189, n23190, n23191, n23192,
    n23193, n23194, n23195, n23196, n23197, n23198,
    n23199, n23200, n23201, n23202, n23203, n23204,
    n23205, n23206, n23207, n23208, n23209, n23210,
    n23211, n23212, n23213, n23214, n23215, n23216,
    n23217, n23218, n23219, n23220, n23221, n23222,
    n23223, n23224, n23225, n23226, n23227, n23228,
    n23229, n23230, n23231, n23232, n23233, n23234,
    n23235, n23236, n23237, n23238, n23239, n23240,
    n23241, n23242, n23243, n23244, n23245, n23246,
    n23247, n23248, n23249, n23250, n23251, n23252,
    n23253, n23254, n23255, n23256, n23257, n23258,
    n23259, n23260, n23261, n23262, n23263, n23264,
    n23265, n23266, n23267, n23268, n23269, n23270,
    n23271, n23272, n23273, n23274, n23275, n23276,
    n23277, n23278, n23279, n23280, n23281, n23282,
    n23283, n23284, n23285, n23286, n23287, n23288,
    n23289, n23290, n23291, n23292, n23293, n23294,
    n23295, n23296, n23297, n23298, n23299, n23300,
    n23301, n23302, n23303, n23304, n23305, n23306,
    n23307, n23308, n23309, n23310, n23311, n23312,
    n23313, n23314, n23315, n23316, n23317, n23318,
    n23319, n23320, n23321, n23322, n23323, n23324,
    n23325, n23326, n23327, n23328, n23329, n23330,
    n23331, n23332, n23333, n23334, n23335, n23336,
    n23337, n23338, n23339, n23340, n23341, n23342,
    n23343, n23344, n23345, n23346, n23347, n23348,
    n23349, n23350, n23351, n23352, n23353, n23354,
    n23355, n23356, n23357, n23358, n23359, n23360,
    n23361, n23362, n23363, n23364, n23365, n23366,
    n23367, n23368, n23369, n23370, n23371, n23372,
    n23373, n23374, n23375, n23376, n23377, n23378,
    n23379, n23380, n23381, n23382, n23383, n23384,
    n23385, n23386, n23387, n23388, n23389, n23390,
    n23391, n23392, n23393, n23394, n23395, n23396,
    n23397, n23398, n23399, n23400, n23401, n23402,
    n23403, n23404, n23405, n23406, n23407, n23408,
    n23409, n23410, n23411, n23412, n23413, n23414,
    n23415, n23416, n23417, n23418, n23419, n23420,
    n23421, n23422, n23423, n23424, n23425, n23426,
    n23427, n23428, n23429, n23430, n23431, n23432,
    n23433, n23434, n23435, n23436, n23437, n23438,
    n23439, n23440, n23441, n23442, n23443, n23444,
    n23445, n23446, n23447, n23448, n23449, n23450,
    n23451, n23452, n23453, n23454, n23455, n23456,
    n23457, n23458, n23459, n23460, n23461, n23462,
    n23463, n23464, n23465, n23466, n23467, n23468,
    n23469, n23470, n23471, n23472, n23473, n23474,
    n23475, n23476, n23477, n23478, n23479, n23480,
    n23481, n23482, n23483, n23484, n23485, n23486,
    n23487, n23488, n23489, n23490, n23491, n23492,
    n23493, n23494, n23495, n23496, n23497, n23498,
    n23499, n23500, n23501, n23502, n23503, n23504,
    n23505, n23506, n23507, n23508, n23509, n23510,
    n23511, n23512, n23513, n23514, n23515, n23516,
    n23517, n23518, n23519, n23520, n23521, n23522,
    n23523, n23524, n23525, n23526, n23527, n23528,
    n23529, n23530, n23531, n23532, n23533, n23534,
    n23535, n23536, n23537, n23538, n23539, n23540,
    n23541, n23542, n23543, n23544, n23545, n23546,
    n23547, n23548, n23549, n23550, n23551, n23552,
    n23553, n23554, n23555, n23556, n23557, n23558,
    n23559, n23560, n23561, n23562, n23563, n23564,
    n23565, n23566, n23567, n23568, n23569, n23570,
    n23571, n23572, n23573, n23574, n23575, n23576,
    n23577, n23578, n23579, n23580, n23581, n23582,
    n23583, n23584, n23585, n23586, n23587, n23588,
    n23589, n23590, n23591, n23592, n23593, n23594,
    n23595, n23596, n23597, n23598, n23599, n23600,
    n23601, n23602, n23603, n23604, n23605, n23606,
    n23607, n23608, n23609, n23610, n23611, n23612,
    n23613, n23614, n23615, n23616, n23617, n23618,
    n23619, n23620, n23621, n23622, n23623, n23624,
    n23625, n23626, n23627, n23628, n23629, n23630,
    n23631, n23632, n23633, n23634, n23635, n23636,
    n23637, n23638, n23639, n23640, n23641, n23642,
    n23643, n23644, n23645, n23646, n23647, n23648,
    n23649, n23650, n23651, n23652, n23653, n23654,
    n23655, n23656, n23657, n23658, n23659, n23660,
    n23661, n23662, n23663, n23664, n23665, n23666,
    n23667, n23668, n23669, n23670, n23671, n23672,
    n23673, n23674, n23675, n23676, n23677, n23678,
    n23679, n23680, n23681, n23682, n23683, n23684,
    n23685, n23686, n23687, n23688, n23689, n23690,
    n23691, n23692, n23693, n23694, n23695, n23696,
    n23697, n23698, n23699, n23700, n23701, n23702,
    n23703, n23704, n23705, n23706, n23707, n23708,
    n23709, n23710, n23711, n23712, n23713, n23714,
    n23715, n23716, n23717, n23718, n23719, n23720,
    n23721, n23722, n23723, n23724, n23725, n23726,
    n23727, n23728, n23729, n23730, n23731, n23732,
    n23733, n23734, n23735, n23736, n23737, n23738,
    n23739, n23740, n23741, n23742, n23743, n23744,
    n23745, n23746, n23747, n23748, n23749, n23750,
    n23751, n23752, n23753, n23754, n23755, n23756,
    n23757, n23758, n23759, n23760, n23761, n23762,
    n23763, n23764, n23765, n23766, n23767, n23768,
    n23769, n23770, n23771, n23772, n23773, n23774,
    n23775, n23776, n23777, n23778, n23779, n23780,
    n23781, n23782, n23783, n23784, n23785, n23786,
    n23787, n23788, n23789, n23790, n23791, n23792,
    n23793, n23794, n23795, n23796, n23797, n23798,
    n23799, n23800, n23801, n23802, n23803, n23804,
    n23805, n23806, n23807, n23808, n23809, n23810,
    n23811, n23812, n23813, n23814, n23815, n23816,
    n23817, n23818, n23819, n23820, n23821, n23822,
    n23823, n23824, n23825, n23826, n23827, n23828,
    n23829, n23830, n23831, n23832, n23833, n23834,
    n23835, n23836, n23837, n23838, n23839, n23840,
    n23841, n23842, n23843, n23844, n23845, n23846,
    n23847, n23848, n23849, n23850, n23851, n23852,
    n23853, n23854, n23855, n23856, n23857, n23858,
    n23859, n23860, n23861, n23862, n23863, n23864,
    n23865, n23866, n23867, n23868, n23869, n23870,
    n23871, n23872, n23873, n23874, n23875, n23876,
    n23877, n23878, n23879, n23880, n23881, n23882,
    n23883, n23884, n23885, n23886, n23887, n23888,
    n23889, n23890, n23891, n23892, n23893, n23894,
    n23895, n23896, n23897, n23898, n23899, n23900,
    n23901, n23902, n23903, n23904, n23905, n23906,
    n23907, n23908, n23909, n23910, n23911, n23912,
    n23913, n23914, n23915, n23916, n23917, n23918,
    n23919, n23920, n23921, n23922, n23923, n23924,
    n23925, n23926, n23927, n23928, n23929, n23930,
    n23931, n23932, n23933, n23934, n23935, n23936,
    n23937, n23938, n23939, n23940, n23941, n23942,
    n23943, n23944, n23945, n23946, n23947, n23948,
    n23949, n23950, n23951, n23952, n23953, n23954,
    n23955, n23956, n23957, n23958, n23959, n23960,
    n23961, n23962, n23963, n23964, n23965, n23966,
    n23967, n23968, n23969, n23970, n23971, n23972,
    n23973, n23974, n23975, n23976, n23977, n23978,
    n23979, n23980, n23981, n23982, n23983, n23984,
    n23985, n23986, n23987, n23988, n23989, n23990,
    n23991, n23992, n23993, n23994, n23995, n23996,
    n23997, n23998, n23999, n24000, n24001, n24002,
    n24003, n24004, n24005, n24006, n24007, n24008,
    n24009, n24010, n24011, n24012, n24013, n24014,
    n24015, n24016, n24017, n24018, n24019, n24020,
    n24021, n24022, n24023, n24024, n24025, n24026,
    n24027, n24028, n24029, n24030, n24031, n24032,
    n24033, n24034, n24035, n24036, n24037, n24038,
    n24039, n24040, n24041, n24042, n24043, n24044,
    n24045, n24046, n24047, n24048, n24049, n24050,
    n24051, n24052, n24053, n24054, n24055, n24056,
    n24057, n24058, n24059, n24060, n24061, n24062,
    n24063, n24064, n24065, n24066, n24067, n24068,
    n24069, n24070, n24071, n24072, n24073, n24074,
    n24075, n24076, n24077, n24078, n24079, n24080,
    n24081, n24082, n24083, n24084, n24085, n24086,
    n24087, n24088, n24089, n24090, n24091, n24092,
    n24093, n24094, n24095, n24096, n24097, n24098,
    n24099, n24100, n24101, n24102, n24103, n24104,
    n24105, n24106, n24107, n24108, n24109, n24110,
    n24111, n24112, n24113, n24114, n24115, n24116,
    n24117, n24118, n24119, n24120, n24121, n24122,
    n24123, n24124, n24125, n24126, n24127, n24128,
    n24129, n24130, n24131, n24132, n24133, n24134,
    n24135, n24136, n24137, n24138, n24139, n24140,
    n24141, n24142, n24143, n24144, n24145, n24146,
    n24147, n24148, n24149, n24150, n24151, n24152,
    n24153, n24154, n24155, n24156, n24157, n24158,
    n24159, n24160, n24161, n24162, n24163, n24164,
    n24165, n24166, n24167, n24168, n24169, n24170,
    n24171, n24172, n24173, n24174, n24175, n24176,
    n24177, n24178, n24179, n24180, n24181, n24182,
    n24183, n24184, n24185, n24186, n24187, n24188,
    n24189, n24190, n24191, n24192, n24193, n24194,
    n24195, n24196, n24197, n24198, n24199, n24200,
    n24201, n24202, n24203, n24204, n24205, n24206,
    n24207, n24208, n24209, n24210, n24211, n24212,
    n24213, n24214, n24215, n24216, n24217, n24218,
    n24219, n24220, n24221, n24222, n24223, n24224,
    n24225, n24226, n24227, n24228, n24229, n24230,
    n24231, n24232, n24233, n24234, n24235, n24236,
    n24237, n24238, n24239, n24240, n24241, n24242,
    n24243, n24244, n24245, n24246, n24247, n24248,
    n24249, n24250, n24251, n24252, n24253, n24254,
    n24255, n24256, n24257, n24258, n24259, n24260,
    n24261, n24262, n24263, n24264, n24265, n24266,
    n24267, n24268, n24269, n24270, n24271, n24272,
    n24273, n24274, n24275, n24276, n24277, n24278,
    n24279, n24280, n24281, n24282, n24283, n24284,
    n24285, n24286, n24287, n24288, n24289, n24290,
    n24291, n24292, n24293, n24294, n24295, n24296,
    n24297, n24298, n24299, n24300, n24301, n24302,
    n24303, n24304, n24305, n24306, n24307, n24308,
    n24309, n24310, n24311, n24312, n24313, n24314,
    n24315, n24316, n24317, n24318, n24319, n24320,
    n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332,
    n24333, n24334, n24335, n24336, n24337, n24338,
    n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350,
    n24351, n24352, n24353, n24354, n24355, n24356,
    n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368,
    n24369, n24370, n24371, n24372, n24373, n24374,
    n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386,
    n24387, n24388, n24389, n24390, n24391, n24392,
    n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404,
    n24405, n24406, n24407, n24408, n24409, n24410,
    n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422,
    n24423, n24424, n24425, n24426, n24427, n24428,
    n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440,
    n24441, n24442, n24443, n24444, n24445, n24446,
    n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24458,
    n24459, n24460, n24461, n24462, n24463, n24464,
    n24465, n24466, n24467, n24468, n24469, n24470,
    n24471, n24472, n24473, n24474, n24475, n24476,
    n24477, n24478, n24479, n24480, n24481, n24482,
    n24483, n24484, n24485, n24486, n24487, n24488,
    n24489, n24490, n24491, n24492, n24493, n24494,
    n24495, n24496, n24497, n24498, n24499, n24500,
    n24501, n24502, n24503, n24504, n24505, n24506,
    n24507, n24508, n24509, n24510, n24511, n24512,
    n24513, n24514, n24515, n24516, n24517, n24518,
    n24519, n24520, n24521, n24522, n24523, n24524,
    n24525, n24526, n24527, n24528, n24529, n24530,
    n24531, n24532, n24533, n24534, n24535, n24536,
    n24537, n24538, n24539, n24540, n24541, n24542,
    n24543, n24544, n24545, n24546, n24547, n24548,
    n24549, n24550, n24551, n24552, n24553, n24554,
    n24555, n24556, n24557, n24558, n24559, n24560,
    n24561, n24562, n24563, n24564, n24565, n24566,
    n24567, n24568, n24569, n24570, n24571, n24572,
    n24573, n24574, n24575, n24576, n24577, n24578,
    n24579, n24580, n24581, n24582, n24583, n24584,
    n24585, n24586, n24587, n24588, n24589, n24590,
    n24591, n24592, n24593, n24594, n24595, n24596,
    n24597, n24598, n24599, n24600, n24601, n24602,
    n24603, n24604, n24605, n24606, n24607, n24608,
    n24609, n24610, n24611, n24612, n24613, n24614,
    n24615, n24616, n24617, n24618, n24619, n24620,
    n24621, n24622, n24623, n24624, n24625, n24626,
    n24627, n24628, n24629, n24630, n24631, n24632,
    n24633, n24634, n24635, n24636, n24637, n24638,
    n24639, n24640, n24641, n24642, n24643, n24644,
    n24645, n24646, n24647, n24648, n24649, n24650,
    n24651, n24652, n24653, n24654, n24655, n24656,
    n24657, n24658, n24659, n24660, n24661, n24662,
    n24663, n24664, n24665, n24666, n24667, n24668,
    n24669, n24670, n24671, n24672, n24673, n24674,
    n24675, n24676, n24677, n24678, n24679, n24680,
    n24681, n24682, n24683, n24684, n24685, n24686,
    n24687, n24688, n24689, n24690, n24691, n24692,
    n24693, n24694, n24695, n24696, n24697, n24698,
    n24699, n24700, n24701, n24702, n24703, n24704,
    n24705, n24706, n24707, n24708, n24709, n24710,
    n24711, n24712, n24713, n24714, n24715, n24716,
    n24717, n24718, n24719, n24720, n24721, n24722,
    n24723, n24724, n24725, n24726, n24727, n24728,
    n24729, n24730, n24731, n24732, n24733, n24734,
    n24735, n24736, n24737, n24738, n24739, n24740,
    n24741, n24742, n24743, n24744, n24745, n24746,
    n24747, n24748, n24749, n24750, n24751, n24752,
    n24753, n24754, n24755, n24756, n24757, n24758,
    n24759, n24760, n24761, n24762, n24763, n24764,
    n24765, n24766, n24767, n24768, n24769, n24770,
    n24771, n24772, n24773, n24774, n24775, n24776,
    n24777, n24778, n24779, n24780, n24781, n24782,
    n24783, n24784, n24785, n24786, n24787, n24788,
    n24789, n24790, n24791, n24792, n24793, n24794,
    n24795, n24796, n24797, n24798, n24799, n24800,
    n24801, n24802, n24803, n24804, n24805, n24806,
    n24807, n24808, n24809, n24810, n24811, n24812,
    n24813, n24814, n24815, n24816, n24817, n24818,
    n24819, n24820, n24821, n24822, n24823, n24824,
    n24825, n24826, n24827, n24828, n24829, n24830,
    n24831, n24832, n24833, n24834, n24835, n24836,
    n24837, n24838, n24839, n24840, n24841, n24842,
    n24843, n24844, n24845, n24846, n24847, n24848,
    n24849, n24850, n24851, n24852, n24853, n24854,
    n24855, n24856, n24857, n24858, n24859, n24860,
    n24861, n24862, n24863, n24864, n24865, n24866,
    n24867, n24868, n24869, n24870, n24871, n24872,
    n24873, n24874, n24875, n24876, n24877, n24878,
    n24879, n24880, n24881, n24882, n24883, n24884,
    n24885, n24886, n24887, n24888, n24889, n24890,
    n24891, n24892, n24893, n24894, n24895, n24896,
    n24897, n24898, n24899, n24900, n24901, n24902,
    n24903, n24904, n24905, n24906, n24907, n24908,
    n24909, n24910, n24911, n24912, n24913, n24914,
    n24915, n24916, n24917, n24918, n24919, n24920,
    n24921, n24922, n24923, n24924, n24925, n24926,
    n24927, n24928, n24929, n24930, n24931, n24932,
    n24933, n24934, n24935, n24936, n24937, n24938,
    n24939, n24940, n24941, n24942, n24943, n24944,
    n24945, n24946, n24947, n24948, n24949, n24950,
    n24951, n24952, n24953, n24954, n24955, n24956,
    n24957, n24958, n24959, n24960, n24961, n24962,
    n24963, n24964, n24965, n24966, n24967, n24968,
    n24969, n24970, n24971, n24972, n24973, n24974,
    n24975, n24976, n24977, n24978, n24979, n24980,
    n24981, n24982, n24983, n24984, n24985, n24986,
    n24987, n24988, n24989, n24990, n24991, n24992,
    n24993, n24994, n24995, n24996, n24997, n24998,
    n24999, n25000, n25001, n25002, n25003, n25004,
    n25005, n25006, n25007, n25008, n25009, n25010,
    n25011, n25012, n25013, n25014, n25015, n25016,
    n25017, n25018, n25019, n25020, n25021, n25022,
    n25023, n25024, n25025, n25026, n25027, n25028,
    n25029, n25030, n25031, n25032, n25033, n25034,
    n25035, n25036, n25037, n25038, n25039, n25040,
    n25041, n25042, n25043, n25044, n25045, n25046,
    n25047, n25048, n25049, n25050, n25051, n25052,
    n25053, n25054, n25055, n25056, n25057, n25058,
    n25059, n25060, n25061, n25062, n25063, n25064,
    n25065, n25066, n25067, n25068, n25069, n25070,
    n25071, n25072, n25073, n25074, n25075, n25076,
    n25077, n25078, n25079, n25080, n25081, n25082,
    n25083, n25084, n25085, n25086, n25087, n25088,
    n25089, n25090, n25091, n25092, n25093, n25094,
    n25095, n25096, n25097, n25098, n25099, n25100,
    n25101, n25102, n25103, n25104, n25105, n25106,
    n25107, n25108, n25109, n25110, n25111, n25112,
    n25113, n25114, n25115, n25116, n25117, n25118,
    n25119, n25120, n25121, n25122, n25123, n25124,
    n25125, n25126, n25127, n25128, n25129, n25130,
    n25131, n25132, n25133, n25134, n25135, n25136,
    n25137, n25138, n25139, n25140, n25141, n25142,
    n25143, n25144, n25145, n25146, n25147, n25148,
    n25149, n25150, n25151, n25152, n25153, n25154,
    n25155, n25156, n25157, n25158, n25159, n25160,
    n25161, n25162, n25163, n25164, n25165, n25166,
    n25167, n25168, n25169, n25170, n25171, n25172,
    n25173, n25174, n25175, n25176, n25177, n25178,
    n25179, n25180, n25181, n25182, n25183, n25184,
    n25185, n25186, n25187, n25188, n25189, n25190,
    n25191, n25192, n25193, n25194, n25195, n25196,
    n25197, n25198, n25199, n25200, n25201, n25202,
    n25203, n25204, n25205, n25206, n25207, n25208,
    n25209, n25210, n25211, n25212, n25213, n25214,
    n25215, n25216, n25217, n25218, n25219, n25220,
    n25221, n25222, n25223, n25224, n25225, n25226,
    n25227, n25228, n25229, n25230, n25231, n25232,
    n25233, n25234, n25235, n25236, n25237, n25238,
    n25239, n25240, n25241, n25242, n25243, n25244,
    n25245, n25246, n25247, n25248, n25249, n25250,
    n25251, n25252, n25253, n25254, n25255, n25256,
    n25257, n25258, n25259, n25260, n25261, n25262,
    n25263, n25264, n25265, n25266, n25267, n25268,
    n25269, n25270, n25271, n25272, n25273, n25274,
    n25275, n25276, n25277, n25278, n25279, n25280,
    n25281, n25282, n25283, n25284, n25285, n25286,
    n25287, n25288, n25289, n25290, n25291, n25292,
    n25293, n25294, n25295, n25296, n25297, n25298,
    n25299, n25300, n25301, n25302, n25303, n25304,
    n25305, n25306, n25307, n25308, n25309, n25310,
    n25311, n25312, n25313, n25314, n25315, n25316,
    n25317, n25318, n25319, n25320, n25321, n25322,
    n25323, n25324, n25325, n25326, n25327, n25328,
    n25329, n25330, n25331, n25332, n25333, n25334,
    n25335, n25336, n25337, n25338, n25339, n25340,
    n25341, n25342, n25343, n25344, n25345, n25346,
    n25347, n25348, n25349, n25350, n25351, n25352,
    n25353, n25354, n25355, n25356, n25357, n25358,
    n25359, n25360, n25361, n25362, n25363, n25364,
    n25365, n25366, n25367, n25368, n25369, n25370,
    n25371, n25372, n25373, n25374, n25375, n25376,
    n25377, n25378, n25379, n25380, n25381, n25382,
    n25383, n25384, n25385, n25386, n25387, n25388,
    n25389, n25390, n25391, n25392, n25393, n25394,
    n25395, n25396, n25397, n25398, n25399, n25400,
    n25401, n25402, n25403, n25404, n25405, n25406,
    n25407, n25408, n25409, n25410, n25411, n25412,
    n25413, n25414, n25415, n25416, n25417, n25418,
    n25419, n25420, n25421, n25422, n25423, n25424,
    n25425, n25426, n25427, n25428, n25429, n25430,
    n25431, n25432, n25433, n25434, n25435, n25436,
    n25437, n25438, n25439, n25440, n25441, n25442,
    n25443, n25444, n25445, n25446, n25447, n25448,
    n25449, n25450, n25451, n25452, n25453, n25454,
    n25455, n25456, n25457, n25458, n25459, n25460,
    n25461, n25462, n25463, n25464, n25465, n25466,
    n25467, n25468, n25469, n25470, n25471, n25472,
    n25473, n25474, n25475, n25476, n25477, n25478,
    n25479, n25480, n25481, n25482, n25483, n25484,
    n25485, n25486, n25487, n25488, n25489, n25490,
    n25491, n25492, n25493, n25494, n25495, n25496,
    n25497, n25498, n25499, n25500, n25501, n25502,
    n25503, n25504, n25505, n25506, n25507, n25508,
    n25509, n25510, n25511, n25512, n25513, n25514,
    n25515, n25516, n25517, n25518, n25519, n25520,
    n25521, n25522, n25523, n25524, n25525, n25526,
    n25527, n25528, n25529, n25530, n25531, n25532,
    n25533, n25534, n25535, n25536, n25537, n25538,
    n25539, n25540, n25541, n25542, n25543, n25544,
    n25545, n25546, n25547, n25548, n25550, n25551,
    n25552, n25553, n25554, n25555, n25556, n25557,
    n25558, n25559, n25560, n25561, n25562, n25563,
    n25564, n25565, n25566, n25567, n25568, n25569,
    n25570, n25571, n25572, n25573, n25574, n25575,
    n25576, n25577, n25578, n25579, n25580, n25581,
    n25582, n25583, n25584, n25585, n25586, n25587,
    n25588, n25589, n25590, n25591, n25592, n25593,
    n25594, n25595, n25596, n25597, n25598, n25599,
    n25600, n25601, n25602, n25603, n25604, n25605,
    n25606, n25607, n25608, n25609, n25610, n25611,
    n25612, n25613, n25614, n25615, n25616, n25617,
    n25618, n25619, n25620, n25621, n25622, n25623,
    n25624, n25625, n25626, n25627, n25628, n25629,
    n25630, n25631, n25632, n25633, n25634, n25635,
    n25636, n25637, n25638, n25639, n25640, n25641,
    n25642, n25643, n25644, n25645, n25646, n25647,
    n25648, n25649, n25650, n25651, n25652, n25653,
    n25654, n25655, n25656, n25657, n25658, n25659,
    n25660, n25661, n25662, n25663, n25664, n25665,
    n25666, n25667, n25668, n25669, n25670, n25671,
    n25672, n25673, n25674, n25675, n25676, n25677,
    n25678, n25679, n25680, n25681, n25682, n25683,
    n25684, n25685, n25686, n25687, n25688, n25689,
    n25690, n25691, n25692, n25693, n25694, n25695,
    n25696, n25697, n25698, n25699, n25700, n25701,
    n25702, n25703, n25704, n25705, n25706, n25707,
    n25708, n25709, n25710, n25711, n25712, n25713,
    n25714, n25715, n25716, n25717, n25718, n25719,
    n25720, n25721, n25722, n25723, n25724, n25725,
    n25726, n25727, n25728, n25729, n25730, n25731,
    n25732, n25733, n25734, n25735, n25736, n25737,
    n25738, n25739, n25740, n25741, n25742, n25743,
    n25744, n25745, n25746, n25747, n25748, n25749,
    n25750, n25751, n25752, n25753, n25754, n25755,
    n25756, n25757, n25758, n25759, n25760, n25761,
    n25762, n25763, n25764, n25765, n25766, n25767,
    n25768, n25769, n25770, n25771, n25772, n25773,
    n25774, n25775, n25776, n25777, n25778, n25779,
    n25780, n25781, n25782, n25783, n25784, n25785,
    n25786, n25787, n25788, n25789, n25790, n25791,
    n25792, n25793, n25794, n25795, n25796, n25797,
    n25798, n25799, n25800, n25801, n25802, n25803,
    n25804, n25805, n25806, n25807, n25808, n25809,
    n25811, n25812, n25813, n25814, n25815, n25816,
    n25817, n25818, n25819, n25820, n25821, n25822,
    n25823, n25824, n25825, n25826, n25827, n25828,
    n25829, n25830, n25831, n25832, n25833, n25834,
    n25835, n25836, n25837, n25838, n25839, n25840,
    n25841, n25842, n25843, n25844, n25845, n25846,
    n25847, n25848, n25849, n25850, n25851, n25852,
    n25853, n25854, n25855, n25856, n25857, n25858,
    n25859, n25860, n25861, n25862, n25863, n25864,
    n25865, n25866, n25867, n25868, n25869, n25870,
    n25871, n25872, n25873, n25874, n25875, n25876,
    n25877, n25878, n25879, n25880, n25881, n25882,
    n25883, n25884, n25885, n25886, n25887, n25888,
    n25889, n25890, n25891, n25892, n25893, n25894,
    n25895, n25896, n25897, n25898, n25899, n25900,
    n25901, n25902, n25903, n25904, n25905, n25906,
    n25907, n25908, n25909, n25910, n25911, n25912,
    n25913, n25914, n25915, n25916, n25917, n25918,
    n25919, n25920, n25921, n25922, n25923, n25924,
    n25925, n25926, n25927, n25928, n25929, n25930,
    n25931, n25932, n25933, n25934, n25935, n25936,
    n25937, n25938, n25939, n25940, n25941, n25942,
    n25943, n25944, n25945, n25946, n25947, n25948,
    n25949, n25950, n25951, n25952, n25953, n25954,
    n25955, n25956, n25957, n25958, n25959, n25960,
    n25961, n25962, n25963, n25964, n25965, n25966,
    n25967, n25968, n25969, n25970, n25971, n25972,
    n25973, n25974, n25975, n25976, n25977, n25978,
    n25979, n25980, n25981, n25982, n25983, n25984,
    n25985, n25986, n25987, n25988, n25989, n25990,
    n25991, n25992, n25993, n25994, n25995, n25996,
    n25997, n25998, n25999, n26000, n26001, n26002,
    n26003, n26004, n26005, n26006, n26007, n26008,
    n26009, n26010, n26011, n26012, n26013, n26014,
    n26015, n26016, n26017, n26018, n26019, n26020,
    n26021, n26022, n26023, n26024, n26025, n26026,
    n26027, n26028, n26029, n26030, n26031, n26032,
    n26033, n26034, n26035, n26036, n26037, n26038,
    n26039, n26040, n26041, n26042, n26043, n26044,
    n26045, n26046, n26047, n26048, n26049, n26050,
    n26051, n26052, n26053, n26054, n26055, n26056,
    n26057, n26058, n26059, n26060, n26061, n26062,
    n26063, n26064, n26065, n26067, n26068, n26069,
    n26070, n26071, n26072, n26073, n26074, n26075,
    n26076, n26077, n26078, n26079, n26080, n26081,
    n26082, n26083, n26084, n26085, n26086, n26087,
    n26088, n26089, n26090, n26091, n26092, n26093,
    n26094, n26095, n26096, n26097, n26098, n26099,
    n26100, n26101, n26102, n26103, n26104, n26105,
    n26106, n26107, n26108, n26109, n26110, n26111,
    n26112, n26113, n26114, n26115, n26116, n26117,
    n26118, n26119, n26120, n26121, n26122, n26123,
    n26124, n26125, n26126, n26127, n26128, n26129,
    n26130, n26131, n26132, n26133, n26134, n26135,
    n26136, n26137, n26138, n26139, n26140, n26141,
    n26142, n26143, n26144, n26145, n26146, n26147,
    n26148, n26149, n26150, n26151, n26152, n26153,
    n26154, n26155, n26156, n26157, n26158, n26159,
    n26160, n26161, n26162, n26163, n26164, n26165,
    n26166, n26167, n26168, n26169, n26170, n26171,
    n26172, n26173, n26174, n26175, n26176, n26177,
    n26178, n26179, n26180, n26181, n26182, n26183,
    n26184, n26185, n26186, n26187, n26188, n26189,
    n26190, n26191, n26192, n26193, n26194, n26195,
    n26196, n26197, n26198, n26199, n26200, n26201,
    n26202, n26203, n26204, n26205, n26206, n26207,
    n26208, n26209, n26210, n26211, n26212, n26213,
    n26214, n26215, n26216, n26217, n26218, n26219,
    n26220, n26221, n26222, n26223, n26224, n26225,
    n26226, n26227, n26228, n26229, n26230, n26231,
    n26232, n26233, n26234, n26235, n26236, n26237,
    n26238, n26239, n26240, n26241, n26242, n26243,
    n26244, n26245, n26246, n26247, n26248, n26249,
    n26250, n26251, n26252, n26253, n26254, n26255,
    n26256, n26257, n26258, n26259, n26260, n26261,
    n26262, n26263, n26264, n26265, n26266, n26267,
    n26268, n26269, n26270, n26271, n26272, n26273,
    n26274, n26275, n26276, n26277, n26278, n26279,
    n26280, n26281, n26282, n26283, n26284, n26285,
    n26286, n26287, n26288, n26289, n26290, n26291,
    n26292, n26293, n26294, n26295, n26296, n26297,
    n26298, n26299, n26300, n26301, n26302, n26303,
    n26304, n26305, n26306, n26308, n26309, n26310,
    n26311, n26312, n26313, n26314, n26315, n26316,
    n26317, n26318, n26319, n26320, n26321, n26322,
    n26323, n26324, n26325, n26326, n26327, n26328,
    n26329, n26330, n26331, n26332, n26333, n26334,
    n26335, n26336, n26337, n26338, n26339, n26340,
    n26341, n26342, n26343, n26344, n26345, n26346,
    n26347, n26348, n26349, n26350, n26351, n26352,
    n26353, n26354, n26355, n26356, n26357, n26358,
    n26359, n26360, n26361, n26362, n26363, n26364,
    n26365, n26366, n26367, n26368, n26369, n26370,
    n26371, n26372, n26373, n26374, n26375, n26376,
    n26377, n26378, n26379, n26380, n26381, n26382,
    n26383, n26384, n26385, n26386, n26387, n26388,
    n26389, n26390, n26391, n26392, n26393, n26394,
    n26395, n26396, n26397, n26398, n26399, n26400,
    n26401, n26402, n26403, n26404, n26405, n26406,
    n26407, n26408, n26409, n26410, n26411, n26412,
    n26413, n26414, n26415, n26416, n26417, n26418,
    n26419, n26420, n26421, n26422, n26423, n26424,
    n26425, n26426, n26427, n26428, n26429, n26430,
    n26431, n26432, n26433, n26434, n26435, n26436,
    n26437, n26438, n26439, n26440, n26441, n26442,
    n26443, n26444, n26445, n26446, n26447, n26448,
    n26449, n26450, n26451, n26452, n26453, n26454,
    n26455, n26456, n26457, n26458, n26459, n26460,
    n26461, n26462, n26463, n26464, n26465, n26466,
    n26467, n26468, n26469, n26470, n26471, n26472,
    n26473, n26474, n26475, n26476, n26477, n26478,
    n26479, n26480, n26481, n26482, n26483, n26484,
    n26485, n26486, n26487, n26488, n26489, n26490,
    n26491, n26492, n26493, n26494, n26495, n26496,
    n26497, n26498, n26499, n26500, n26501, n26502,
    n26503, n26504, n26505, n26506, n26507, n26508,
    n26509, n26510, n26511, n26512, n26513, n26514,
    n26515, n26516, n26517, n26518, n26519, n26520,
    n26521, n26522, n26523, n26524, n26525, n26526,
    n26527, n26528, n26529, n26530, n26531, n26532,
    n26533, n26534, n26535, n26536, n26537, n26538,
    n26539, n26540, n26541, n26542, n26543, n26544,
    n26545, n26546, n26547, n26548, n26549, n26550,
    n26551, n26552, n26553, n26554, n26555, n26556,
    n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26571, n26572, n26573, n26574, n26575,
    n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587,
    n26588, n26589, n26590, n26591, n26592, n26593,
    n26594, n26595, n26596, n26597, n26598, n26599,
    n26600, n26601, n26602, n26603, n26604, n26605,
    n26606, n26607, n26608, n26609, n26610, n26611,
    n26612, n26613, n26614, n26615, n26616, n26617,
    n26618, n26619, n26620, n26621, n26622, n26623,
    n26624, n26625, n26626, n26627, n26628, n26629,
    n26630, n26631, n26632, n26633, n26634, n26635,
    n26636, n26637, n26638, n26639, n26640, n26641,
    n26642, n26643, n26644, n26645, n26646, n26647,
    n26648, n26649, n26650, n26651, n26652, n26653,
    n26654, n26655, n26656, n26657, n26658, n26659,
    n26660, n26661, n26662, n26663, n26664, n26665,
    n26666, n26667, n26668, n26669, n26670, n26671,
    n26672, n26673, n26674, n26675, n26676, n26677,
    n26678, n26679, n26680, n26681, n26682, n26683,
    n26684, n26685, n26686, n26687, n26688, n26689,
    n26690, n26691, n26692, n26693, n26694, n26695,
    n26696, n26697, n26698, n26699, n26700, n26701,
    n26702, n26703, n26704, n26705, n26706, n26707,
    n26708, n26709, n26710, n26711, n26712, n26713,
    n26714, n26715, n26716, n26717, n26718, n26719,
    n26720, n26721, n26722, n26723, n26724, n26725,
    n26726, n26727, n26728, n26729, n26730, n26731,
    n26732, n26733, n26734, n26735, n26736, n26737,
    n26738, n26739, n26740, n26741, n26742, n26743,
    n26744, n26745, n26746, n26747, n26748, n26749,
    n26750, n26751, n26752, n26753, n26754, n26755,
    n26756, n26757, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767,
    n26768, n26769, n26770, n26771, n26772, n26773,
    n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785,
    n26786, n26788, n26789, n26790, n26791, n26792,
    n26793, n26794, n26795, n26796, n26797, n26798,
    n26799, n26800, n26801, n26802, n26803, n26804,
    n26805, n26806, n26807, n26808, n26809, n26810,
    n26811, n26812, n26813, n26814, n26815, n26816,
    n26817, n26818, n26819, n26820, n26821, n26822,
    n26823, n26824, n26825, n26826, n26827, n26828,
    n26829, n26830, n26831, n26832, n26833, n26834,
    n26835, n26836, n26837, n26838, n26839, n26840,
    n26841, n26842, n26843, n26844, n26845, n26846,
    n26847, n26848, n26849, n26850, n26851, n26852,
    n26853, n26854, n26855, n26856, n26857, n26858,
    n26859, n26860, n26861, n26862, n26863, n26864,
    n26865, n26866, n26867, n26868, n26869, n26870,
    n26871, n26872, n26873, n26874, n26875, n26876,
    n26877, n26878, n26879, n26880, n26881, n26882,
    n26883, n26884, n26885, n26886, n26887, n26888,
    n26889, n26890, n26891, n26892, n26893, n26894,
    n26895, n26896, n26897, n26898, n26899, n26900,
    n26901, n26902, n26903, n26904, n26905, n26906,
    n26907, n26908, n26909, n26910, n26911, n26912,
    n26913, n26914, n26915, n26916, n26917, n26918,
    n26919, n26920, n26921, n26922, n26923, n26924,
    n26925, n26926, n26927, n26928, n26929, n26930,
    n26931, n26932, n26933, n26934, n26935, n26936,
    n26937, n26938, n26939, n26940, n26941, n26942,
    n26943, n26944, n26945, n26946, n26947, n26948,
    n26949, n26950, n26951, n26952, n26953, n26954,
    n26955, n26956, n26957, n26958, n26959, n26960,
    n26961, n26962, n26963, n26964, n26965, n26966,
    n26967, n26968, n26969, n26970, n26971, n26972,
    n26973, n26974, n26975, n26976, n26977, n26978,
    n26979, n26980, n26981, n26982, n26983, n26984,
    n26985, n26986, n26987, n26988, n26989, n26990,
    n26991, n26992, n26993, n26994, n26995, n26996,
    n26997, n26998, n26999, n27000, n27001, n27002,
    n27003, n27004, n27005, n27006, n27007, n27009,
    n27010, n27011, n27012, n27013, n27014, n27015,
    n27016, n27017, n27018, n27019, n27020, n27021,
    n27022, n27023, n27024, n27025, n27026, n27027,
    n27028, n27029, n27030, n27031, n27032, n27033,
    n27034, n27035, n27036, n27037, n27038, n27039,
    n27040, n27041, n27042, n27043, n27044, n27045,
    n27046, n27047, n27048, n27049, n27050, n27051,
    n27052, n27053, n27054, n27055, n27056, n27057,
    n27058, n27059, n27060, n27061, n27062, n27063,
    n27064, n27065, n27066, n27067, n27068, n27069,
    n27070, n27071, n27072, n27073, n27074, n27075,
    n27076, n27077, n27078, n27079, n27080, n27081,
    n27082, n27083, n27084, n27085, n27086, n27087,
    n27088, n27089, n27090, n27091, n27092, n27093,
    n27094, n27095, n27096, n27097, n27098, n27099,
    n27100, n27101, n27102, n27103, n27104, n27105,
    n27106, n27107, n27108, n27109, n27110, n27111,
    n27112, n27113, n27114, n27115, n27116, n27117,
    n27118, n27119, n27120, n27121, n27122, n27123,
    n27124, n27125, n27126, n27127, n27128, n27129,
    n27130, n27131, n27132, n27133, n27134, n27135,
    n27136, n27137, n27138, n27139, n27140, n27141,
    n27142, n27143, n27144, n27145, n27146, n27147,
    n27148, n27149, n27150, n27151, n27152, n27153,
    n27154, n27155, n27156, n27157, n27158, n27159,
    n27160, n27161, n27162, n27163, n27164, n27165,
    n27166, n27167, n27168, n27169, n27170, n27171,
    n27172, n27173, n27174, n27175, n27176, n27177,
    n27178, n27179, n27180, n27181, n27182, n27183,
    n27184, n27185, n27186, n27187, n27188, n27189,
    n27190, n27191, n27192, n27193, n27194, n27195,
    n27196, n27197, n27198, n27199, n27200, n27201,
    n27202, n27203, n27204, n27205, n27206, n27207,
    n27208, n27209, n27210, n27212, n27213, n27214,
    n27215, n27216, n27217, n27218, n27219, n27220,
    n27221, n27222, n27223, n27224, n27225, n27226,
    n27227, n27228, n27229, n27230, n27231, n27232,
    n27233, n27234, n27235, n27236, n27237, n27238,
    n27239, n27240, n27241, n27242, n27243, n27244,
    n27245, n27246, n27247, n27248, n27249, n27250,
    n27251, n27252, n27253, n27254, n27255, n27256,
    n27257, n27258, n27259, n27260, n27261, n27262,
    n27263, n27264, n27265, n27266, n27267, n27268,
    n27269, n27270, n27271, n27272, n27273, n27274,
    n27275, n27276, n27277, n27278, n27279, n27280,
    n27281, n27282, n27283, n27284, n27285, n27286,
    n27287, n27288, n27289, n27290, n27291, n27292,
    n27293, n27294, n27295, n27296, n27297, n27298,
    n27299, n27300, n27301, n27302, n27303, n27304,
    n27305, n27306, n27307, n27308, n27309, n27310,
    n27311, n27312, n27313, n27314, n27315, n27316,
    n27317, n27318, n27319, n27320, n27321, n27322,
    n27323, n27324, n27325, n27326, n27327, n27328,
    n27329, n27330, n27331, n27332, n27333, n27334,
    n27335, n27336, n27337, n27338, n27339, n27340,
    n27341, n27342, n27343, n27344, n27345, n27346,
    n27347, n27348, n27349, n27350, n27351, n27352,
    n27353, n27354, n27355, n27356, n27357, n27358,
    n27359, n27360, n27361, n27362, n27363, n27364,
    n27365, n27366, n27367, n27368, n27369, n27370,
    n27371, n27372, n27373, n27374, n27375, n27376,
    n27377, n27378, n27379, n27380, n27381, n27382,
    n27383, n27384, n27385, n27386, n27387, n27388,
    n27389, n27390, n27391, n27392, n27393, n27394,
    n27395, n27396, n27397, n27398, n27399, n27400,
    n27401, n27402, n27403, n27404, n27405, n27406,
    n27407, n27408, n27409, n27410, n27411, n27412,
    n27413, n27414, n27415, n27416, n27417, n27418,
    n27420, n27421, n27422, n27423, n27424, n27425,
    n27426, n27427, n27428, n27429, n27430, n27431,
    n27432, n27433, n27434, n27435, n27436, n27437,
    n27438, n27439, n27440, n27441, n27442, n27443,
    n27444, n27445, n27446, n27447, n27448, n27449,
    n27450, n27451, n27452, n27453, n27454, n27455,
    n27456, n27457, n27458, n27459, n27460, n27461,
    n27462, n27463, n27464, n27465, n27466, n27467,
    n27468, n27469, n27470, n27471, n27472, n27473,
    n27474, n27475, n27476, n27477, n27478, n27479,
    n27480, n27481, n27482, n27483, n27484, n27485,
    n27486, n27487, n27488, n27489, n27490, n27491,
    n27492, n27493, n27494, n27495, n27496, n27497,
    n27498, n27499, n27500, n27501, n27502, n27503,
    n27504, n27505, n27506, n27507, n27508, n27509,
    n27510, n27511, n27512, n27513, n27514, n27515,
    n27516, n27517, n27518, n27519, n27520, n27521,
    n27522, n27523, n27524, n27525, n27526, n27527,
    n27528, n27529, n27530, n27531, n27532, n27533,
    n27534, n27535, n27536, n27537, n27538, n27539,
    n27540, n27541, n27542, n27543, n27544, n27545,
    n27546, n27547, n27548, n27549, n27550, n27551,
    n27552, n27553, n27554, n27555, n27556, n27557,
    n27558, n27559, n27560, n27561, n27562, n27563,
    n27564, n27565, n27566, n27567, n27568, n27569,
    n27570, n27571, n27572, n27573, n27574, n27575,
    n27576, n27577, n27578, n27579, n27580, n27581,
    n27582, n27583, n27584, n27585, n27586, n27587,
    n27588, n27589, n27590, n27591, n27592, n27593,
    n27594, n27595, n27596, n27597, n27598, n27599,
    n27600, n27601, n27602, n27603, n27604, n27605,
    n27606, n27607, n27608, n27609, n27610, n27611,
    n27612, n27613, n27614, n27615, n27616, n27617,
    n27618, n27619, n27620, n27622, n27623, n27624,
    n27625, n27626, n27627, n27628, n27629, n27630,
    n27631, n27632, n27633, n27634, n27635, n27636,
    n27637, n27638, n27639, n27640, n27641, n27642,
    n27643, n27644, n27645, n27646, n27647, n27648,
    n27649, n27650, n27651, n27652, n27653, n27654,
    n27655, n27656, n27657, n27658, n27659, n27660,
    n27661, n27662, n27663, n27664, n27665, n27666,
    n27667, n27668, n27669, n27670, n27671, n27672,
    n27673, n27674, n27675, n27676, n27677, n27678,
    n27679, n27680, n27681, n27682, n27683, n27684,
    n27685, n27686, n27687, n27688, n27689, n27690,
    n27691, n27692, n27693, n27694, n27695, n27696,
    n27697, n27698, n27699, n27700, n27701, n27702,
    n27703, n27704, n27705, n27706, n27707, n27708,
    n27709, n27710, n27711, n27712, n27713, n27714,
    n27715, n27716, n27717, n27718, n27719, n27720,
    n27721, n27722, n27723, n27724, n27725, n27726,
    n27727, n27728, n27729, n27730, n27731, n27732,
    n27733, n27734, n27735, n27736, n27737, n27738,
    n27739, n27740, n27741, n27742, n27743, n27744,
    n27745, n27746, n27747, n27748, n27749, n27750,
    n27751, n27752, n27753, n27754, n27755, n27756,
    n27757, n27758, n27759, n27760, n27761, n27762,
    n27763, n27764, n27765, n27766, n27767, n27768,
    n27769, n27770, n27771, n27772, n27773, n27774,
    n27775, n27776, n27777, n27778, n27779, n27780,
    n27781, n27782, n27783, n27784, n27785, n27786,
    n27787, n27788, n27789, n27790, n27791, n27792,
    n27793, n27794, n27795, n27796, n27797, n27798,
    n27799, n27800, n27801, n27802, n27803, n27804,
    n27805, n27806, n27807, n27808, n27809, n27810,
    n27811, n27812, n27813, n27814, n27815, n27816,
    n27817, n27819, n27820, n27821, n27822, n27823,
    n27824, n27825, n27826, n27827, n27828, n27829,
    n27830, n27831, n27832, n27833, n27834, n27835,
    n27836, n27837, n27838, n27839, n27840, n27841,
    n27842, n27843, n27844, n27845, n27846, n27847,
    n27848, n27849, n27850, n27851, n27852, n27853,
    n27854, n27855, n27856, n27857, n27858, n27859,
    n27860, n27861, n27862, n27863, n27864, n27865,
    n27866, n27867, n27868, n27869, n27870, n27871,
    n27872, n27873, n27874, n27875, n27876, n27877,
    n27878, n27879, n27880, n27881, n27882, n27883,
    n27884, n27885, n27886, n27887, n27888, n27889,
    n27890, n27891, n27892, n27893, n27894, n27895,
    n27896, n27897, n27898, n27899, n27900, n27901,
    n27902, n27903, n27904, n27905, n27906, n27907,
    n27908, n27909, n27910, n27911, n27912, n27913,
    n27914, n27915, n27916, n27917, n27918, n27919,
    n27920, n27921, n27922, n27923, n27924, n27925,
    n27926, n27927, n27928, n27929, n27930, n27931,
    n27932, n27933, n27934, n27935, n27936, n27937,
    n27938, n27939, n27940, n27941, n27942, n27943,
    n27944, n27945, n27946, n27947, n27948, n27949,
    n27950, n27951, n27952, n27953, n27954, n27955,
    n27956, n27957, n27958, n27959, n27960, n27961,
    n27962, n27963, n27964, n27965, n27966, n27967,
    n27968, n27969, n27970, n27971, n27972, n27973,
    n27974, n27975, n27976, n27977, n27978, n27979,
    n27980, n27981, n27982, n27983, n27984, n27985,
    n27986, n27987, n27988, n27989, n27990, n27991,
    n27992, n27993, n27994, n27995, n27996, n27997,
    n27998, n27999, n28000, n28001, n28002, n28003,
    n28004, n28005, n28006, n28007, n28008, n28009,
    n28010, n28011, n28012, n28013, n28014, n28015,
    n28016, n28018, n28019, n28020, n28021, n28022,
    n28023, n28024, n28025, n28026, n28027, n28028,
    n28029, n28030, n28031, n28032, n28033, n28034,
    n28035, n28036, n28037, n28038, n28039, n28040,
    n28041, n28042, n28043, n28044, n28045, n28046,
    n28047, n28048, n28049, n28050, n28051, n28052,
    n28053, n28054, n28055, n28056, n28057, n28058,
    n28059, n28060, n28061, n28062, n28063, n28064,
    n28065, n28066, n28067, n28068, n28069, n28070,
    n28071, n28072, n28073, n28074, n28075, n28076,
    n28077, n28078, n28079, n28080, n28081, n28082,
    n28083, n28084, n28085, n28086, n28087, n28088,
    n28089, n28090, n28091, n28092, n28093, n28094,
    n28095, n28096, n28097, n28098, n28099, n28100,
    n28101, n28102, n28103, n28104, n28105, n28106,
    n28107, n28108, n28109, n28110, n28111, n28112,
    n28113, n28114, n28115, n28116, n28117, n28118,
    n28119, n28120, n28121, n28122, n28123, n28124,
    n28125, n28126, n28127, n28128, n28129, n28130,
    n28131, n28132, n28133, n28134, n28135, n28136,
    n28137, n28138, n28139, n28140, n28141, n28142,
    n28143, n28144, n28145, n28146, n28147, n28148,
    n28149, n28150, n28151, n28152, n28153, n28154,
    n28155, n28156, n28157, n28158, n28159, n28160,
    n28161, n28162, n28163, n28164, n28165, n28166,
    n28167, n28168, n28169, n28170, n28171, n28172,
    n28173, n28174, n28175, n28176, n28177, n28178,
    n28179, n28180, n28181, n28182, n28183, n28184,
    n28185, n28186, n28187, n28188, n28189, n28190,
    n28191, n28192, n28193, n28194, n28195, n28196,
    n28197, n28198, n28199, n28200, n28201, n28202,
    n28203, n28204, n28205, n28206, n28207, n28208,
    n28209, n28210, n28211, n28212, n28213, n28214,
    n28215, n28216, n28218, n28219, n28220, n28221,
    n28222, n28223, n28224, n28225, n28226, n28227,
    n28228, n28229, n28230, n28231, n28232, n28233,
    n28234, n28235, n28236, n28237, n28238, n28239,
    n28240, n28241, n28242, n28243, n28244, n28245,
    n28246, n28247, n28248, n28249, n28250, n28251,
    n28252, n28253, n28254, n28255, n28256, n28257,
    n28258, n28259, n28260, n28261, n28262, n28263,
    n28264, n28265, n28266, n28267, n28268, n28269,
    n28270, n28271, n28272, n28273, n28274, n28275,
    n28276, n28277, n28278, n28279, n28280, n28281,
    n28282, n28283, n28284, n28285, n28286, n28287,
    n28288, n28289, n28290, n28291, n28292, n28293,
    n28294, n28295, n28296, n28297, n28298, n28299,
    n28300, n28301, n28302, n28303, n28304, n28305,
    n28306, n28307, n28308, n28309, n28310, n28311,
    n28312, n28313, n28314, n28315, n28316, n28317,
    n28318, n28319, n28320, n28321, n28322, n28323,
    n28324, n28325, n28326, n28327, n28328, n28329,
    n28330, n28331, n28332, n28333, n28334, n28335,
    n28336, n28337, n28338, n28339, n28340, n28341,
    n28342, n28343, n28344, n28345, n28346, n28347,
    n28348, n28349, n28350, n28351, n28352, n28353,
    n28354, n28355, n28356, n28357, n28358, n28359,
    n28360, n28361, n28362, n28363, n28364, n28365,
    n28366, n28367, n28368, n28369, n28370, n28371,
    n28372, n28373, n28374, n28375, n28376, n28377,
    n28378, n28379, n28380, n28381, n28382, n28383,
    n28384, n28385, n28386, n28387, n28388, n28389,
    n28390, n28391, n28392, n28394, n28395, n28396,
    n28397, n28398, n28399, n28400, n28401, n28402,
    n28403, n28404, n28405, n28406, n28407, n28408,
    n28409, n28410, n28411, n28412, n28413, n28414,
    n28415, n28416, n28417, n28418, n28419, n28420,
    n28421, n28422, n28423, n28424, n28425, n28426,
    n28427, n28428, n28429, n28430, n28431, n28432,
    n28433, n28434, n28435, n28436, n28437, n28438,
    n28439, n28440, n28441, n28442, n28443, n28444,
    n28445, n28446, n28447, n28448, n28449, n28450,
    n28451, n28452, n28453, n28454, n28455, n28456,
    n28457, n28458, n28459, n28460, n28461, n28462,
    n28463, n28464, n28465, n28466, n28467, n28468,
    n28469, n28470, n28471, n28472, n28473, n28474,
    n28475, n28476, n28477, n28478, n28479, n28480,
    n28481, n28482, n28483, n28484, n28485, n28486,
    n28487, n28488, n28489, n28490, n28491, n28492,
    n28493, n28494, n28495, n28496, n28497, n28498,
    n28499, n28500, n28501, n28502, n28503, n28504,
    n28505, n28506, n28507, n28508, n28509, n28510,
    n28511, n28512, n28513, n28514, n28515, n28516,
    n28517, n28518, n28519, n28520, n28521, n28522,
    n28523, n28524, n28525, n28526, n28527, n28528,
    n28529, n28530, n28531, n28532, n28533, n28534,
    n28535, n28536, n28537, n28538, n28539, n28540,
    n28541, n28542, n28543, n28544, n28545, n28546,
    n28547, n28548, n28549, n28550, n28551, n28552,
    n28553, n28554, n28555, n28556, n28557, n28558,
    n28560, n28561, n28562, n28563, n28564, n28565,
    n28566, n28567, n28568, n28569, n28570, n28571,
    n28572, n28573, n28574, n28575, n28576, n28577,
    n28578, n28579, n28580, n28581, n28582, n28583,
    n28584, n28585, n28586, n28587, n28588, n28589,
    n28590, n28591, n28592, n28593, n28594, n28595,
    n28596, n28597, n28598, n28599, n28600, n28601,
    n28602, n28603, n28604, n28605, n28606, n28607,
    n28608, n28609, n28610, n28611, n28612, n28613,
    n28614, n28615, n28616, n28617, n28618, n28619,
    n28620, n28621, n28622, n28623, n28624, n28625,
    n28626, n28627, n28628, n28629, n28630, n28631,
    n28632, n28633, n28634, n28635, n28636, n28637,
    n28638, n28639, n28640, n28641, n28642, n28643,
    n28644, n28645, n28646, n28647, n28648, n28649,
    n28650, n28651, n28652, n28653, n28654, n28655,
    n28656, n28657, n28658, n28659, n28660, n28661,
    n28662, n28663, n28664, n28665, n28666, n28667,
    n28668, n28669, n28670, n28671, n28672, n28673,
    n28674, n28675, n28676, n28677, n28678, n28679,
    n28680, n28681, n28682, n28683, n28684, n28685,
    n28686, n28687, n28688, n28689, n28690, n28691,
    n28692, n28693, n28694, n28695, n28696, n28697,
    n28698, n28699, n28700, n28701, n28702, n28703,
    n28704, n28705, n28706, n28707, n28708, n28709,
    n28710, n28711, n28712, n28713, n28714, n28715,
    n28716, n28717, n28718, n28719, n28720, n28721,
    n28722, n28723, n28724, n28726, n28727, n28728,
    n28729, n28730, n28731, n28732, n28733, n28734,
    n28735, n28736, n28737, n28738, n28739, n28740,
    n28741, n28742, n28743, n28744, n28745, n28746,
    n28747, n28748, n28749, n28750, n28751, n28752,
    n28753, n28754, n28755, n28756, n28757, n28758,
    n28759, n28760, n28761, n28762, n28763, n28764,
    n28765, n28766, n28767, n28768, n28769, n28770,
    n28771, n28772, n28773, n28774, n28775, n28776,
    n28777, n28778, n28779, n28780, n28781, n28782,
    n28783, n28784, n28785, n28786, n28787, n28788,
    n28789, n28790, n28791, n28792, n28793, n28794,
    n28795, n28796, n28797, n28798, n28799, n28800,
    n28801, n28802, n28803, n28804, n28805, n28806,
    n28807, n28808, n28809, n28810, n28811, n28812,
    n28813, n28814, n28815, n28816, n28817, n28818,
    n28819, n28820, n28821, n28822, n28823, n28824,
    n28825, n28826, n28827, n28828, n28829, n28830,
    n28831, n28832, n28833, n28834, n28835, n28836,
    n28837, n28838, n28839, n28840, n28841, n28842,
    n28843, n28844, n28845, n28846, n28847, n28848,
    n28849, n28850, n28851, n28852, n28853, n28854,
    n28855, n28856, n28857, n28858, n28859, n28860,
    n28861, n28862, n28863, n28864, n28865, n28866,
    n28867, n28868, n28869, n28870, n28871, n28872,
    n28873, n28874, n28875, n28876, n28877, n28878,
    n28879, n28880, n28881, n28882, n28883, n28884,
    n28886, n28887, n28888, n28889, n28890, n28891,
    n28892, n28893, n28894, n28895, n28896, n28897,
    n28898, n28899, n28900, n28901, n28902, n28903,
    n28904, n28905, n28906, n28907, n28908, n28909,
    n28910, n28911, n28912, n28913, n28914, n28915,
    n28916, n28917, n28918, n28919, n28920, n28921,
    n28922, n28923, n28924, n28925, n28926, n28927,
    n28928, n28929, n28930, n28931, n28932, n28933,
    n28934, n28935, n28936, n28937, n28938, n28939,
    n28940, n28941, n28942, n28943, n28944, n28945,
    n28946, n28947, n28948, n28949, n28950, n28951,
    n28952, n28953, n28954, n28955, n28956, n28957,
    n28958, n28959, n28960, n28961, n28962, n28963,
    n28964, n28965, n28966, n28967, n28968, n28969,
    n28970, n28971, n28972, n28973, n28974, n28975,
    n28976, n28977, n28978, n28979, n28980, n28981,
    n28982, n28983, n28984, n28985, n28986, n28987,
    n28988, n28989, n28990, n28991, n28992, n28993,
    n28994, n28995, n28996, n28997, n28998, n28999,
    n29000, n29001, n29002, n29003, n29004, n29005,
    n29006, n29007, n29008, n29009, n29010, n29011,
    n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023,
    n29024, n29025, n29026, n29027, n29028, n29029,
    n29030, n29031, n29032, n29034, n29035, n29036,
    n29037, n29038, n29039, n29040, n29041, n29042,
    n29043, n29044, n29045, n29046, n29047, n29048,
    n29049, n29050, n29051, n29052, n29053, n29054,
    n29055, n29056, n29057, n29058, n29059, n29060,
    n29061, n29062, n29063, n29064, n29065, n29066,
    n29067, n29068, n29069, n29070, n29071, n29072,
    n29073, n29074, n29075, n29076, n29077, n29078,
    n29079, n29080, n29081, n29082, n29083, n29084,
    n29085, n29086, n29087, n29088, n29089, n29090,
    n29091, n29092, n29093, n29094, n29095, n29096,
    n29097, n29098, n29099, n29100, n29101, n29102,
    n29103, n29104, n29105, n29106, n29107, n29108,
    n29109, n29110, n29111, n29112, n29113, n29114,
    n29115, n29116, n29117, n29118, n29119, n29120,
    n29121, n29122, n29123, n29124, n29125, n29126,
    n29127, n29128, n29129, n29130, n29131, n29132,
    n29133, n29134, n29135, n29136, n29137, n29138,
    n29139, n29140, n29141, n29142, n29143, n29144,
    n29145, n29146, n29147, n29148, n29149, n29150,
    n29151, n29152, n29153, n29154, n29155, n29156,
    n29157, n29158, n29159, n29160, n29161, n29162,
    n29163, n29164, n29165, n29166, n29167, n29168,
    n29169, n29170, n29171, n29172, n29173, n29174,
    n29175, n29176, n29177, n29178, n29179, n29181,
    n29182, n29183, n29184, n29185, n29186, n29187,
    n29188, n29189, n29190, n29191, n29192, n29193,
    n29194, n29195, n29196, n29197, n29198, n29199,
    n29200, n29201, n29202, n29203, n29204, n29205,
    n29206, n29207, n29208, n29209, n29210, n29211,
    n29212, n29213, n29214, n29215, n29216, n29217,
    n29218, n29219, n29220, n29221, n29222, n29223,
    n29224, n29225, n29226, n29227, n29228, n29229,
    n29230, n29231, n29232, n29233, n29234, n29235,
    n29236, n29237, n29238, n29239, n29240, n29241,
    n29242, n29243, n29244, n29245, n29246, n29247,
    n29248, n29249, n29250, n29251, n29252, n29253,
    n29254, n29255, n29256, n29257, n29258, n29259,
    n29260, n29261, n29262, n29263, n29264, n29265,
    n29266, n29267, n29268, n29269, n29270, n29271,
    n29272, n29273, n29274, n29275, n29276, n29277,
    n29278, n29279, n29280, n29281, n29282, n29283,
    n29284, n29285, n29286, n29287, n29288, n29289,
    n29290, n29291, n29292, n29293, n29294, n29295,
    n29296, n29297, n29298, n29299, n29300, n29301,
    n29302, n29303, n29304, n29305, n29306, n29307,
    n29308, n29309, n29310, n29311, n29312, n29313,
    n29314, n29315, n29316, n29317, n29319, n29320,
    n29321, n29322, n29323, n29324, n29325, n29326,
    n29327, n29328, n29329, n29330, n29331, n29332,
    n29333, n29334, n29335, n29336, n29337, n29338,
    n29339, n29340, n29341, n29342, n29343, n29344,
    n29345, n29346, n29347, n29348, n29349, n29350,
    n29351, n29352, n29353, n29354, n29355, n29356,
    n29357, n29358, n29359, n29360, n29361, n29362,
    n29363, n29364, n29365, n29366, n29367, n29368,
    n29369, n29370, n29371, n29372, n29373, n29374,
    n29375, n29376, n29377, n29378, n29379, n29380,
    n29381, n29382, n29383, n29384, n29385, n29386,
    n29387, n29388, n29389, n29390, n29391, n29392,
    n29393, n29394, n29395, n29396, n29397, n29398,
    n29399, n29400, n29401, n29402, n29403, n29404,
    n29405, n29406, n29407, n29408, n29409, n29410,
    n29411, n29412, n29413, n29414, n29415, n29416,
    n29417, n29418, n29419, n29420, n29421, n29422,
    n29423, n29424, n29425, n29426, n29427, n29428,
    n29429, n29430, n29431, n29432, n29433, n29434,
    n29435, n29436, n29437, n29438, n29439, n29440,
    n29441, n29442, n29443, n29444, n29445, n29446,
    n29447, n29448, n29450, n29451, n29452, n29453,
    n29454, n29455, n29456, n29457, n29458, n29459,
    n29460, n29461, n29462, n29463, n29464, n29465,
    n29466, n29467, n29468, n29469, n29470, n29471,
    n29472, n29473, n29474, n29475, n29476, n29477,
    n29478, n29479, n29480, n29481, n29482, n29483,
    n29484, n29485, n29486, n29487, n29488, n29489,
    n29490, n29491, n29492, n29493, n29494, n29495,
    n29496, n29497, n29498, n29499, n29500, n29501,
    n29502, n29503, n29504, n29505, n29506, n29507,
    n29508, n29509, n29510, n29511, n29512, n29513,
    n29514, n29515, n29516, n29517, n29518, n29519,
    n29520, n29521, n29522, n29523, n29524, n29525,
    n29526, n29527, n29528, n29529, n29530, n29531,
    n29532, n29533, n29534, n29535, n29536, n29537,
    n29538, n29539, n29540, n29541, n29542, n29543,
    n29544, n29545, n29546, n29547, n29548, n29549,
    n29550, n29551, n29552, n29553, n29554, n29555,
    n29556, n29557, n29558, n29559, n29560, n29561,
    n29562, n29563, n29564, n29565, n29566, n29567,
    n29568, n29569, n29570, n29571, n29572, n29573,
    n29574, n29575, n29576, n29577, n29579, n29580,
    n29581, n29582, n29583, n29584, n29585, n29586,
    n29587, n29588, n29589, n29590, n29591, n29592,
    n29593, n29594, n29595, n29596, n29597, n29598,
    n29599, n29600, n29601, n29602, n29603, n29604,
    n29605, n29606, n29607, n29608, n29609, n29610,
    n29611, n29612, n29613, n29614, n29615, n29616,
    n29617, n29618, n29619, n29620, n29621, n29622,
    n29623, n29624, n29625, n29626, n29627, n29628,
    n29629, n29630, n29631, n29632, n29633, n29634,
    n29635, n29636, n29637, n29638, n29639, n29640,
    n29641, n29642, n29643, n29644, n29645, n29646,
    n29647, n29648, n29649, n29650, n29651, n29652,
    n29653, n29654, n29655, n29656, n29657, n29658,
    n29659, n29660, n29661, n29662, n29663, n29664,
    n29665, n29666, n29667, n29668, n29669, n29670,
    n29671, n29672, n29673, n29674, n29675, n29676,
    n29677, n29678, n29679, n29680, n29681, n29682,
    n29683, n29684, n29685, n29686, n29687, n29688,
    n29689, n29690, n29691, n29692, n29693, n29694,
    n29695, n29696, n29697, n29698, n29700, n29701,
    n29702, n29703, n29704, n29705, n29706, n29707,
    n29708, n29709, n29710, n29711, n29712, n29713,
    n29714, n29715, n29716, n29717, n29718, n29719,
    n29720, n29721, n29722, n29723, n29724, n29725,
    n29726, n29727, n29728, n29729, n29730, n29731,
    n29732, n29733, n29734, n29735, n29736, n29737,
    n29738, n29739, n29740, n29741, n29742, n29743,
    n29744, n29745, n29746, n29747, n29748, n29749,
    n29750, n29751, n29752, n29753, n29754, n29755,
    n29756, n29757, n29758, n29759, n29760, n29761,
    n29762, n29763, n29764, n29765, n29766, n29767,
    n29768, n29769, n29770, n29771, n29772, n29773,
    n29774, n29775, n29776, n29777, n29778, n29779,
    n29780, n29781, n29782, n29783, n29784, n29785,
    n29786, n29787, n29788, n29789, n29790, n29791,
    n29792, n29793, n29794, n29795, n29796, n29797,
    n29798, n29799, n29800, n29801, n29802, n29803,
    n29804, n29805, n29806, n29807, n29808, n29809,
    n29810, n29812, n29813, n29814, n29815, n29816,
    n29817, n29818, n29819, n29820, n29821, n29822,
    n29823, n29824, n29825, n29826, n29827, n29828,
    n29829, n29830, n29831, n29832, n29833, n29834,
    n29835, n29836, n29837, n29838, n29839, n29840,
    n29841, n29842, n29843, n29844, n29845, n29846,
    n29847, n29848, n29849, n29850, n29851, n29852,
    n29853, n29854, n29855, n29856, n29857, n29858,
    n29859, n29860, n29861, n29862, n29863, n29864,
    n29865, n29866, n29867, n29868, n29869, n29870,
    n29871, n29872, n29873, n29874, n29875, n29876,
    n29877, n29878, n29879, n29880, n29881, n29882,
    n29883, n29884, n29885, n29886, n29887, n29888,
    n29889, n29890, n29891, n29892, n29893, n29894,
    n29895, n29896, n29897, n29898, n29899, n29900,
    n29901, n29902, n29903, n29904, n29905, n29906,
    n29907, n29908, n29909, n29910, n29911, n29912,
    n29913, n29914, n29915, n29916, n29917, n29918,
    n29920, n29921, n29922, n29923, n29924, n29925,
    n29926, n29927, n29928, n29929, n29930, n29931,
    n29932, n29933, n29934, n29935, n29936, n29937,
    n29938, n29939, n29940, n29941, n29942, n29943,
    n29944, n29945, n29946, n29947, n29948, n29949,
    n29950, n29951, n29952, n29953, n29954, n29955,
    n29956, n29957, n29958, n29959, n29960, n29961,
    n29962, n29963, n29964, n29965, n29966, n29967,
    n29968, n29969, n29970, n29971, n29972, n29973,
    n29974, n29975, n29976, n29977, n29978, n29979,
    n29980, n29981, n29982, n29983, n29984, n29985,
    n29986, n29987, n29988, n29989, n29990, n29991,
    n29992, n29993, n29994, n29995, n29996, n29997,
    n29998, n29999, n30000, n30001, n30002, n30003,
    n30004, n30005, n30006, n30007, n30008, n30009,
    n30010, n30011, n30012, n30013, n30014, n30015,
    n30016, n30017, n30018, n30019, n30020, n30021,
    n30022, n30023, n30024, n30026, n30027, n30028,
    n30029, n30030, n30031, n30032, n30033, n30034,
    n30035, n30036, n30037, n30038, n30039, n30040,
    n30041, n30042, n30043, n30044, n30045, n30046,
    n30047, n30048, n30049, n30050, n30051, n30052,
    n30053, n30054, n30055, n30056, n30057, n30058,
    n30059, n30060, n30061, n30062, n30063, n30064,
    n30065, n30066, n30067, n30068, n30069, n30070,
    n30071, n30072, n30073, n30074, n30075, n30076,
    n30077, n30078, n30079, n30080, n30081, n30082,
    n30083, n30084, n30085, n30086, n30087, n30088,
    n30089, n30090, n30091, n30092, n30093, n30094,
    n30095, n30096, n30097, n30098, n30099, n30100,
    n30101, n30102, n30103, n30104, n30105, n30106,
    n30107, n30108, n30109, n30110, n30111, n30112,
    n30113, n30114, n30115, n30116, n30117, n30118,
    n30119, n30121, n30122, n30123, n30124, n30125,
    n30126, n30127, n30128, n30129, n30130, n30131,
    n30132, n30133, n30134, n30135, n30136, n30137,
    n30138, n30139, n30140, n30141, n30142, n30143,
    n30144, n30145, n30146, n30147, n30148, n30149,
    n30150, n30151, n30152, n30153, n30154, n30155,
    n30156, n30157, n30158, n30159, n30160, n30161,
    n30162, n30163, n30164, n30165, n30166, n30167,
    n30168, n30169, n30170, n30171, n30172, n30173,
    n30174, n30175, n30176, n30177, n30178, n30179,
    n30180, n30181, n30182, n30183, n30184, n30185,
    n30186, n30187, n30188, n30189, n30190, n30191,
    n30192, n30193, n30194, n30195, n30196, n30197,
    n30198, n30199, n30200, n30201, n30202, n30203,
    n30204, n30205, n30206, n30207, n30208, n30209,
    n30210, n30211, n30213, n30214, n30215, n30216,
    n30217, n30218, n30219, n30220, n30221, n30222,
    n30223, n30224, n30225, n30226, n30227, n30228,
    n30229, n30230, n30231, n30232, n30233, n30234,
    n30235, n30236, n30237, n30238, n30239, n30240,
    n30241, n30242, n30243, n30244, n30245, n30246,
    n30247, n30248, n30249, n30250, n30251, n30252,
    n30253, n30254, n30255, n30256, n30257, n30258,
    n30259, n30260, n30261, n30262, n30263, n30264,
    n30265, n30266, n30267, n30268, n30269, n30270,
    n30271, n30272, n30273, n30274, n30275, n30276,
    n30277, n30278, n30279, n30280, n30281, n30282,
    n30283, n30284, n30285, n30286, n30287, n30288,
    n30289, n30290, n30291, n30292, n30293, n30294,
    n30295, n30296, n30297, n30299, n30300, n30301,
    n30302, n30303, n30304, n30305, n30306, n30307,
    n30308, n30309, n30310, n30311, n30312, n30313,
    n30314, n30315, n30316, n30317, n30318, n30319,
    n30320, n30321, n30322, n30323, n30324, n30325,
    n30326, n30327, n30328, n30329, n30330, n30331,
    n30332, n30333, n30334, n30335, n30336, n30337,
    n30338, n30339, n30340, n30341, n30342, n30343,
    n30344, n30345, n30346, n30347, n30348, n30349,
    n30350, n30351, n30352, n30353, n30354, n30355,
    n30356, n30357, n30358, n30359, n30360, n30361,
    n30362, n30363, n30364, n30365, n30366, n30367,
    n30368, n30369, n30370, n30371, n30372, n30373,
    n30374, n30375, n30377, n30378, n30379, n30380,
    n30381, n30382, n30383, n30384, n30385, n30386,
    n30387, n30388, n30389, n30390, n30391, n30392,
    n30393, n30394, n30395, n30396, n30397, n30398,
    n30399, n30400, n30401, n30402, n30403, n30404,
    n30405, n30406, n30407, n30408, n30409, n30410,
    n30411, n30412, n30413, n30414, n30415, n30416,
    n30417, n30418, n30419, n30420, n30421, n30422,
    n30423, n30424, n30425, n30426, n30427, n30428,
    n30429, n30430, n30431, n30432, n30433, n30434,
    n30435, n30436, n30437, n30438, n30439, n30440,
    n30442, n30443, n30444, n30445, n30446, n30447,
    n30448, n30449, n30450, n30451, n30452, n30453,
    n30454, n30455, n30456, n30457, n30458, n30459,
    n30460, n30461, n30462, n30463, n30464, n30465,
    n30466, n30467, n30468, n30469, n30470, n30471,
    n30472, n30473, n30474, n30475, n30476, n30477,
    n30478, n30479, n30480, n30481, n30482, n30483,
    n30484, n30485, n30486, n30487, n30488, n30489,
    n30490, n30491, n30492, n30493, n30494, n30495;
  assign n65 = ~pi21  & pi22 ;
  assign n66 = pi21  & ~pi22 ;
  assign n67 = ~n65 & ~n66;
  assign n68 = pi20  & ~pi21 ;
  assign n69 = ~pi20  & pi21 ;
  assign n70 = ~n68 & ~n69;
  assign n71 = ~n67 & n70;
  assign n72 = pi27  & pi28 ;
  assign n73 = ~pi29  & pi30 ;
  assign n74 = n72 & n73;
  assign n75 = pi23  & ~pi26 ;
  assign n76 = pi24  & pi25 ;
  assign n77 = n75 & n76;
  assign n78 = n74 & n77;
  assign n79 = ~pi23  & ~pi26 ;
  assign n80 = n76 & n79;
  assign n81 = n74 & n80;
  assign n82 = ~pi24  & ~pi25 ;
  assign n83 = ~pi23  & pi26 ;
  assign n84 = n82 & n83;
  assign n85 = n74 & n84;
  assign n86 = pi23  & pi26 ;
  assign n87 = n82 & n86;
  assign n88 = n74 & n87;
  assign n89 = ~n85 & ~n88;
  assign n90 = pi29  & ~pi30 ;
  assign n91 = n72 & n90;
  assign n92 = pi24  & ~pi25 ;
  assign n93 = n79 & n92;
  assign n94 = n91 & n93;
  assign n95 = ~pi29  & ~pi30 ;
  assign n96 = ~pi27  & ~pi28 ;
  assign n97 = n95 & n96;
  assign n98 = n77 & n97;
  assign n99 = n75 & n82;
  assign n100 = n91 & n99;
  assign n101 = ~n98 & ~n100;
  assign n102 = pi29  & pi30 ;
  assign n103 = n72 & n102;
  assign n104 = n80 & n103;
  assign n105 = n75 & n92;
  assign n106 = n91 & n105;
  assign n107 = ~n104 & ~n106;
  assign n108 = n101 & n107;
  assign n109 = ~n94 & n108;
  assign n110 = ~pi27  & pi28 ;
  assign n111 = n95 & n110;
  assign n112 = n77 & n111;
  assign n113 = n79 & n82;
  assign n114 = n103 & n113;
  assign n115 = n77 & n103;
  assign n116 = n103 & n105;
  assign n117 = n84 & n103;
  assign n118 = ~n116 & ~n117;
  assign n119 = ~n115 & n118;
  assign n120 = ~pi24  & pi25 ;
  assign n121 = n75 & n120;
  assign n122 = n103 & n121;
  assign n123 = n99 & n103;
  assign n124 = ~n122 & ~n123;
  assign n125 = n119 & n124;
  assign n126 = ~n114 & n125;
  assign n127 = n102 & n110;
  assign n128 = n76 & n86;
  assign n129 = n127 & n128;
  assign n130 = n79 & n120;
  assign n131 = n103 & n130;
  assign n132 = n93 & n103;
  assign n133 = n86 & n120;
  assign n134 = n127 & n133;
  assign n135 = ~n132 & ~n134;
  assign n136 = ~n131 & n135;
  assign n137 = ~n129 & n136;
  assign n138 = n126 & n137;
  assign n139 = ~n112 & n138;
  assign n140 = n109 & n139;
  assign n141 = n89 & n140;
  assign n142 = ~n81 & n141;
  assign n143 = ~n78 & n142;
  assign n144 = n74 & n130;
  assign n145 = pi27  & ~pi28 ;
  assign n146 = n90 & n145;
  assign n147 = n128 & n146;
  assign n148 = ~n144 & ~n147;
  assign n149 = n111 & n121;
  assign n150 = n87 & n111;
  assign n151 = n72 & n95;
  assign n152 = n93 & n151;
  assign n153 = n95 & n145;
  assign n154 = n128 & n153;
  assign n155 = n111 & n113;
  assign n156 = ~n154 & ~n155;
  assign n157 = ~n152 & n156;
  assign n158 = ~n150 & n157;
  assign n159 = ~n149 & n158;
  assign n160 = n93 & n111;
  assign n161 = n111 & n128;
  assign n162 = ~n160 & ~n161;
  assign n163 = n84 & n111;
  assign n164 = n76 & n83;
  assign n165 = n111 & n164;
  assign n166 = n133 & n153;
  assign n167 = ~n165 & ~n166;
  assign n168 = ~n163 & n167;
  assign n169 = n83 & n120;
  assign n170 = n111 & n169;
  assign n171 = n113 & n151;
  assign n172 = n111 & n130;
  assign n173 = n80 & n111;
  assign n174 = ~n172 & ~n173;
  assign n175 = ~n171 & n174;
  assign n176 = ~n170 & n175;
  assign n177 = n168 & n176;
  assign n178 = n162 & n177;
  assign n179 = n159 & n178;
  assign n180 = n153 & n164;
  assign n181 = n99 & n146;
  assign n182 = n90 & n110;
  assign n183 = n128 & n182;
  assign n184 = ~n181 & ~n183;
  assign n185 = n83 & n92;
  assign n186 = n146 & n185;
  assign n187 = n164 & n182;
  assign n188 = n130 & n182;
  assign n189 = ~n187 & ~n188;
  assign n190 = ~n186 & n189;
  assign n191 = n184 & n190;
  assign n192 = ~n180 & n191;
  assign n193 = n84 & n97;
  assign n194 = n111 & n133;
  assign n195 = n97 & n121;
  assign n196 = ~n194 & ~n195;
  assign n197 = n74 & n105;
  assign n198 = n105 & n182;
  assign n199 = ~n197 & ~n198;
  assign n200 = n196 & n199;
  assign n201 = ~n193 & n200;
  assign n202 = n192 & n201;
  assign n203 = n127 & n169;
  assign n204 = n103 & n133;
  assign n205 = ~n203 & ~n204;
  assign n206 = n87 & n103;
  assign n207 = n127 & n164;
  assign n208 = n103 & n164;
  assign n209 = ~n207 & ~n208;
  assign n210 = ~n206 & n209;
  assign n211 = n205 & n210;
  assign n212 = n202 & n211;
  assign n213 = n91 & n130;
  assign n214 = n146 & n164;
  assign n215 = ~n213 & ~n214;
  assign n216 = n99 & n111;
  assign n217 = n74 & n185;
  assign n218 = n80 & n91;
  assign n219 = n91 & n121;
  assign n220 = n77 & n91;
  assign n221 = ~n219 & ~n220;
  assign n222 = ~n218 & n221;
  assign n223 = ~n217 & n222;
  assign n224 = ~n216 & n223;
  assign n225 = n215 & n224;
  assign n226 = n212 & n225;
  assign n227 = n86 & n92;
  assign n228 = n103 & n227;
  assign n229 = n103 & n128;
  assign n230 = ~n228 & ~n229;
  assign n231 = n103 & n169;
  assign n232 = n103 & n185;
  assign n233 = ~n231 & ~n232;
  assign n234 = n230 & n233;
  assign n235 = n80 & n146;
  assign n236 = n146 & n227;
  assign n237 = ~n235 & ~n236;
  assign n238 = n121 & n182;
  assign n239 = n133 & n182;
  assign n240 = ~n238 & ~n239;
  assign n241 = n237 & n240;
  assign n242 = n87 & n97;
  assign n243 = n80 & n182;
  assign n244 = ~n242 & ~n243;
  assign n245 = n84 & n91;
  assign n246 = n80 & n97;
  assign n247 = n105 & n111;
  assign n248 = ~n246 & ~n247;
  assign n249 = ~n245 & n248;
  assign n250 = n244 & n249;
  assign n251 = n99 & n151;
  assign n252 = n130 & n146;
  assign n253 = ~n251 & ~n252;
  assign n254 = n182 & n185;
  assign n255 = n111 & n185;
  assign n256 = n111 & n227;
  assign n257 = ~n255 & ~n256;
  assign n258 = ~n254 & n257;
  assign n259 = n74 & n121;
  assign n260 = n84 & n146;
  assign n261 = n99 & n182;
  assign n262 = n113 & n182;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~n260 & n263;
  assign n265 = ~n259 & n264;
  assign n266 = n258 & n265;
  assign n267 = n253 & n266;
  assign n268 = n250 & n267;
  assign n269 = n241 & n268;
  assign n270 = n234 & n269;
  assign n271 = n226 & n270;
  assign n272 = n97 & n130;
  assign n273 = n74 & n227;
  assign n274 = n96 & n102;
  assign n275 = n99 & n274;
  assign n276 = ~n273 & ~n275;
  assign n277 = n121 & n274;
  assign n278 = n74 & n128;
  assign n279 = n74 & n169;
  assign n280 = n74 & n164;
  assign n281 = n130 & n274;
  assign n282 = ~n280 & ~n281;
  assign n283 = ~n279 & n282;
  assign n284 = ~n278 & n283;
  assign n285 = ~n277 & n284;
  assign n286 = n276 & n285;
  assign n287 = ~n272 & n286;
  assign n288 = n77 & n127;
  assign n289 = n127 & n185;
  assign n290 = n93 & n127;
  assign n291 = ~n289 & ~n290;
  assign n292 = n102 & n145;
  assign n293 = n169 & n292;
  assign n294 = n99 & n127;
  assign n295 = ~n293 & ~n294;
  assign n296 = n291 & n295;
  assign n297 = n133 & n292;
  assign n298 = n121 & n127;
  assign n299 = n80 & n127;
  assign n300 = ~n298 & ~n299;
  assign n301 = ~n297 & n300;
  assign n302 = n296 & n301;
  assign n303 = ~n288 & n302;
  assign n304 = n164 & n292;
  assign n305 = n127 & n227;
  assign n306 = ~n304 & ~n305;
  assign n307 = n128 & n292;
  assign n308 = n113 & n127;
  assign n309 = n87 & n127;
  assign n310 = n84 & n127;
  assign n311 = ~n309 & ~n310;
  assign n312 = ~n308 & n311;
  assign n313 = ~n307 & n312;
  assign n314 = n127 & n130;
  assign n315 = n105 & n127;
  assign n316 = ~n314 & ~n315;
  assign n317 = n313 & n316;
  assign n318 = n306 & n317;
  assign n319 = n303 & n318;
  assign n320 = n74 & n133;
  assign n321 = n77 & n274;
  assign n322 = ~n320 & ~n321;
  assign n323 = n99 & n292;
  assign n324 = n97 & n99;
  assign n325 = n93 & n97;
  assign n326 = n97 & n105;
  assign n327 = ~n325 & ~n326;
  assign n328 = ~n324 & n327;
  assign n329 = ~n323 & n328;
  assign n330 = n227 & n274;
  assign n331 = n80 & n292;
  assign n332 = n227 & n292;
  assign n333 = ~n331 & ~n332;
  assign n334 = n121 & n292;
  assign n335 = n333 & ~n334;
  assign n336 = n128 & n274;
  assign n337 = n185 & n274;
  assign n338 = ~n336 & ~n337;
  assign n339 = n335 & n338;
  assign n340 = ~n330 & n339;
  assign n341 = n164 & n274;
  assign n342 = n93 & n292;
  assign n343 = ~n341 & ~n342;
  assign n344 = n130 & n292;
  assign n345 = n87 & n292;
  assign n346 = ~n344 & ~n345;
  assign n347 = n343 & n346;
  assign n348 = n340 & n347;
  assign n349 = n97 & n113;
  assign n350 = n87 & n274;
  assign n351 = ~n349 & ~n350;
  assign n352 = n348 & n351;
  assign n353 = n77 & n292;
  assign n354 = n133 & n274;
  assign n355 = ~n353 & ~n354;
  assign n356 = n84 & n274;
  assign n357 = n185 & n292;
  assign n358 = ~n356 & ~n357;
  assign n359 = n355 & n358;
  assign n360 = n84 & n292;
  assign n361 = n169 & n274;
  assign n362 = n105 & n292;
  assign n363 = n113 & n292;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~n361 & n364;
  assign n366 = ~n360 & n365;
  assign n367 = n359 & n366;
  assign n368 = n352 & n367;
  assign n369 = n329 & n368;
  assign n370 = n322 & n369;
  assign n371 = n319 & n370;
  assign n372 = n105 & n274;
  assign n373 = n93 & n274;
  assign n374 = n113 & n274;
  assign n375 = n80 & n274;
  assign n376 = ~n374 & ~n375;
  assign n377 = ~n373 & n376;
  assign n378 = ~n372 & n377;
  assign n379 = n371 & n378;
  assign n380 = n287 & n379;
  assign n381 = n182 & n227;
  assign n382 = n146 & n169;
  assign n383 = n87 & n182;
  assign n384 = n77 & n146;
  assign n385 = n121 & n146;
  assign n386 = ~n384 & ~n385;
  assign n387 = ~n383 & n386;
  assign n388 = ~n382 & n387;
  assign n389 = ~n381 & n388;
  assign n390 = n84 & n182;
  assign n391 = n169 & n182;
  assign n392 = ~n390 & ~n391;
  assign n393 = n77 & n182;
  assign n394 = n93 & n146;
  assign n395 = n93 & n182;
  assign n396 = ~n394 & ~n395;
  assign n397 = ~n393 & n396;
  assign n398 = n105 & n146;
  assign n399 = n133 & n146;
  assign n400 = n87 & n146;
  assign n401 = n91 & n113;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~n399 & n402;
  assign n404 = ~n398 & n403;
  assign n405 = n397 & n404;
  assign n406 = n392 & n405;
  assign n407 = n389 & n406;
  assign n408 = n380 & n407;
  assign n409 = n271 & n408;
  assign n410 = n179 & n409;
  assign n411 = n148 & n410;
  assign n412 = n143 & n411;
  assign n413 = n87 & n151;
  assign n414 = n133 & n151;
  assign n415 = ~n242 & ~n324;
  assign n416 = ~n100 & ~n106;
  assign n417 = ~n349 & n416;
  assign n418 = ~n94 & n417;
  assign n419 = n415 & n418;
  assign n420 = ~n414 & n419;
  assign n421 = ~n413 & n420;
  assign n422 = n80 & n151;
  assign n423 = n121 & n151;
  assign n424 = n84 & n151;
  assign n425 = ~n423 & ~n424;
  assign n426 = ~n422 & n425;
  assign n427 = n77 & n151;
  assign n428 = n151 & n227;
  assign n429 = n151 & n185;
  assign n430 = n151 & n169;
  assign n431 = ~n429 & ~n430;
  assign n432 = ~n428 & n431;
  assign n433 = ~n427 & n432;
  assign n434 = n426 & n433;
  assign n435 = n130 & n151;
  assign n436 = n105 & n151;
  assign n437 = ~n435 & ~n436;
  assign n438 = n90 & n96;
  assign n439 = n164 & n438;
  assign n440 = n407 & ~n439;
  assign n441 = n185 & n438;
  assign n442 = n113 & n146;
  assign n443 = ~n147 & n241;
  assign n444 = ~n260 & n443;
  assign n445 = ~n198 & ~n254;
  assign n446 = ~n214 & n445;
  assign n447 = ~n252 & n446;
  assign n448 = ~n243 & n263;
  assign n449 = n191 & n448;
  assign n450 = n447 & n449;
  assign n451 = n444 & n450;
  assign n452 = ~n442 & n451;
  assign n453 = ~n441 & n452;
  assign n454 = n227 & n438;
  assign n455 = n169 & n438;
  assign n456 = ~n454 & ~n455;
  assign n457 = n84 & n438;
  assign n458 = n130 & n438;
  assign n459 = ~n457 & ~n458;
  assign n460 = n456 & n459;
  assign n461 = n93 & n438;
  assign n462 = n80 & n438;
  assign n463 = n133 & n438;
  assign n464 = n121 & n438;
  assign n465 = n128 & n438;
  assign n466 = n77 & n438;
  assign n467 = ~n465 & ~n466;
  assign n468 = n87 & n438;
  assign n469 = n128 & n151;
  assign n470 = ~n468 & ~n469;
  assign n471 = n467 & n470;
  assign n472 = ~n464 & n471;
  assign n473 = n105 & n438;
  assign n474 = n99 & n438;
  assign n475 = n151 & n164;
  assign n476 = ~n474 & ~n475;
  assign n477 = n113 & n438;
  assign n478 = n476 & ~n477;
  assign n479 = ~n473 & n478;
  assign n480 = n472 & n479;
  assign n481 = ~n463 & n480;
  assign n482 = ~n462 & n481;
  assign n483 = ~n461 & n482;
  assign n484 = n460 & n483;
  assign n485 = n453 & n484;
  assign n486 = n440 & n485;
  assign n487 = n437 & n486;
  assign n488 = ~n213 & ~n245;
  assign n489 = n222 & n488;
  assign n490 = ~n272 & n489;
  assign n491 = ~n193 & n327;
  assign n492 = ~n195 & ~n246;
  assign n493 = n491 & n492;
  assign n494 = n490 & n493;
  assign n495 = ~n98 & n494;
  assign n496 = n487 & n495;
  assign n497 = n434 & n496;
  assign n498 = n421 & n497;
  assign n499 = n412 & ~n498;
  assign n500 = n121 & n153;
  assign n501 = n80 & n153;
  assign n502 = n153 & n185;
  assign n503 = ~n501 & ~n502;
  assign n504 = n84 & n153;
  assign n505 = n77 & n153;
  assign n506 = n87 & n153;
  assign n507 = ~n505 & ~n506;
  assign n508 = ~n504 & n507;
  assign n509 = n503 & n508;
  assign n510 = ~n500 & n509;
  assign n511 = ~n216 & ~n247;
  assign n512 = n437 & n511;
  assign n513 = ~n251 & n512;
  assign n514 = ~n112 & n513;
  assign n515 = ~n180 & ~n413;
  assign n516 = n257 & n515;
  assign n517 = n153 & n169;
  assign n518 = n153 & n227;
  assign n519 = ~n517 & ~n518;
  assign n520 = n434 & n519;
  assign n521 = ~n194 & n520;
  assign n522 = n516 & n521;
  assign n523 = n179 & n522;
  assign n524 = n514 & n523;
  assign n525 = ~n414 & n524;
  assign n526 = n510 & n525;
  assign n527 = n97 & n164;
  assign n528 = ~n272 & ~n527;
  assign n529 = n415 & n528;
  assign n530 = ~n349 & n492;
  assign n531 = n529 & n530;
  assign n532 = ~n98 & n531;
  assign n533 = n97 & n133;
  assign n534 = n97 & n185;
  assign n535 = n97 & n169;
  assign n536 = n93 & n153;
  assign n537 = n97 & n227;
  assign n538 = n105 & n153;
  assign n539 = ~n537 & ~n538;
  assign n540 = ~n536 & n539;
  assign n541 = ~n535 & n540;
  assign n542 = ~n534 & n541;
  assign n543 = ~n533 & n542;
  assign n544 = n130 & n153;
  assign n545 = n97 & n128;
  assign n546 = ~n544 & ~n545;
  assign n547 = n113 & n153;
  assign n548 = n99 & n153;
  assign n549 = ~n547 & ~n548;
  assign n550 = n546 & n549;
  assign n551 = n543 & n550;
  assign n552 = n491 & n551;
  assign n553 = n532 & n552;
  assign n554 = n526 & n553;
  assign n555 = ~n73 & ~n90;
  assign n556 = pi31  & ~n555;
  assign n557 = ~n166 & n484;
  assign n558 = ~n149 & ~n441;
  assign n559 = n174 & n558;
  assign n560 = n557 & n559;
  assign n561 = ~n247 & n560;
  assign n562 = ~n160 & ~n181;
  assign n563 = ~n442 & n562;
  assign n564 = ~n398 & ~n439;
  assign n565 = n563 & n564;
  assign n566 = ~n216 & n565;
  assign n567 = n156 & ~n252;
  assign n568 = ~n180 & n567;
  assign n569 = ~n394 & n568;
  assign n570 = n566 & n569;
  assign n571 = n519 & n570;
  assign n572 = n561 & n571;
  assign n573 = ~n112 & n572;
  assign n574 = ~n104 & n380;
  assign n575 = n73 & n145;
  assign n576 = n93 & n575;
  assign n577 = n73 & n110;
  assign n578 = n130 & n577;
  assign n579 = n99 & n577;
  assign n580 = n164 & n575;
  assign n581 = n227 & n575;
  assign n582 = n80 & n575;
  assign n583 = n121 & n575;
  assign n584 = ~n582 & ~n583;
  assign n585 = ~n581 & n584;
  assign n586 = ~n580 & n585;
  assign n587 = ~n579 & n586;
  assign n588 = n169 & n575;
  assign n589 = n84 & n575;
  assign n590 = n128 & n575;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n588 & n591;
  assign n593 = n87 & n575;
  assign n594 = n77 & n575;
  assign n595 = n113 & n577;
  assign n596 = ~n594 & ~n595;
  assign n597 = ~n593 & n596;
  assign n598 = n185 & n575;
  assign n599 = n105 & n575;
  assign n600 = n133 & n575;
  assign n601 = n130 & n575;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~n599 & n602;
  assign n604 = ~n598 & n603;
  assign n605 = n597 & n604;
  assign n606 = n592 & n605;
  assign n607 = n587 & n606;
  assign n608 = ~n578 & n607;
  assign n609 = ~n576 & n608;
  assign n610 = n77 & n577;
  assign n611 = n105 & n577;
  assign n612 = n74 & n113;
  assign n613 = n99 & n575;
  assign n614 = n87 & n577;
  assign n615 = ~n613 & ~n614;
  assign n616 = ~n612 & n615;
  assign n617 = ~n611 & n616;
  assign n618 = ~n144 & n617;
  assign n619 = ~n610 & n618;
  assign n620 = n609 & n619;
  assign n621 = n74 & n93;
  assign n622 = n89 & ~n259;
  assign n623 = ~n81 & n622;
  assign n624 = ~n197 & n623;
  assign n625 = ~n621 & n624;
  assign n626 = n93 & n577;
  assign n627 = n169 & n577;
  assign n628 = n128 & n577;
  assign n629 = n185 & n577;
  assign n630 = ~n628 & ~n629;
  assign n631 = n84 & n577;
  assign n632 = n80 & n577;
  assign n633 = n227 & n577;
  assign n634 = ~n632 & ~n633;
  assign n635 = ~n631 & n634;
  assign n636 = n74 & n99;
  assign n637 = n164 & n577;
  assign n638 = n121 & n577;
  assign n639 = n133 & n577;
  assign n640 = ~n638 & ~n639;
  assign n641 = ~n637 & n640;
  assign n642 = ~n636 & n641;
  assign n643 = n635 & n642;
  assign n644 = n630 & n643;
  assign n645 = ~n627 & n644;
  assign n646 = ~n217 & n645;
  assign n647 = ~n78 & n646;
  assign n648 = ~n626 & n647;
  assign n649 = n625 & n648;
  assign n650 = n620 & n649;
  assign n651 = ~n98 & n650;
  assign n652 = n138 & n651;
  assign n653 = n574 & n652;
  assign n654 = ~n207 & n237;
  assign n655 = ~n399 & n654;
  assign n656 = ~n260 & ~n382;
  assign n657 = n655 & n656;
  assign n658 = ~n203 & n657;
  assign n659 = ~n186 & n492;
  assign n660 = ~n400 & n659;
  assign n661 = n658 & n660;
  assign n662 = n386 & n661;
  assign n663 = n653 & n662;
  assign n664 = n509 & n663;
  assign n665 = n573 & n664;
  assign n666 = n113 & n575;
  assign n667 = n91 & n227;
  assign n668 = n87 & n91;
  assign n669 = n91 & n133;
  assign n670 = n91 & n185;
  assign n671 = n91 & n169;
  assign n672 = n91 & n164;
  assign n673 = ~n671 & ~n672;
  assign n674 = ~n670 & n673;
  assign n675 = ~n669 & n674;
  assign n676 = ~n668 & n675;
  assign n677 = n73 & n96;
  assign n678 = n105 & n677;
  assign n679 = n130 & n677;
  assign n680 = ~n678 & ~n679;
  assign n681 = n113 & n677;
  assign n682 = n80 & n677;
  assign n683 = n99 & n677;
  assign n684 = ~n682 & ~n683;
  assign n685 = n121 & n677;
  assign n686 = n684 & ~n685;
  assign n687 = ~n681 & n686;
  assign n688 = n680 & n687;
  assign n689 = n164 & n677;
  assign n690 = n84 & n677;
  assign n691 = ~n689 & ~n690;
  assign n692 = n133 & n677;
  assign n693 = n91 & n128;
  assign n694 = ~n692 & ~n693;
  assign n695 = n185 & n677;
  assign n696 = n694 & ~n695;
  assign n697 = n227 & n677;
  assign n698 = n128 & n677;
  assign n699 = ~n697 & ~n698;
  assign n700 = n93 & n677;
  assign n701 = n77 & n677;
  assign n702 = ~n700 & ~n701;
  assign n703 = n699 & n702;
  assign n704 = n87 & n677;
  assign n705 = n169 & n677;
  assign n706 = ~n704 & ~n705;
  assign n707 = n703 & n706;
  assign n708 = n696 & n707;
  assign n709 = n691 & n708;
  assign n710 = n688 & n709;
  assign n711 = n676 & n710;
  assign n712 = ~n667 & n711;
  assign n713 = n488 & n712;
  assign n714 = ~n94 & n713;
  assign n715 = n222 & n416;
  assign n716 = n714 & n715;
  assign n717 = n486 & n716;
  assign n718 = ~n666 & n717;
  assign n719 = n553 & n718;
  assign n720 = ~n500 & n719;
  assign n721 = ~n665 & ~n720;
  assign n722 = ~n469 & ~n533;
  assign n723 = ~n537 & n722;
  assign n724 = ~n477 & n723;
  assign n725 = ~n183 & ~n534;
  assign n726 = ~n242 & ~n535;
  assign n727 = ~n401 & n623;
  assign n728 = n726 & n727;
  assign n729 = n725 & n728;
  assign n730 = n724 & n729;
  assign n731 = n476 & n730;
  assign n732 = ~n527 & n731;
  assign n733 = n519 & n607;
  assign n734 = ~n324 & n733;
  assign n735 = ~n214 & n734;
  assign n736 = n732 & n735;
  assign n737 = ~n197 & n736;
  assign n738 = ~n170 & ~n505;
  assign n739 = ~n457 & ~n610;
  assign n740 = ~n163 & n739;
  assign n741 = n738 & n740;
  assign n742 = ~n256 & n741;
  assign n743 = ~n461 & n742;
  assign n744 = ~n464 & ~n466;
  assign n745 = ~n502 & n744;
  assign n746 = ~n251 & ~n462;
  assign n747 = ~n611 & n746;
  assign n748 = n745 & n747;
  assign n749 = n645 & n748;
  assign n750 = ~n506 & n749;
  assign n751 = ~n254 & n750;
  assign n752 = n743 & n751;
  assign n753 = ~n504 & ~n578;
  assign n754 = ~n441 & ~n455;
  assign n755 = n753 & n754;
  assign n756 = ~n255 & n755;
  assign n757 = ~n468 & n756;
  assign n758 = ~n165 & ~n626;
  assign n759 = ~n381 & ~n458;
  assign n760 = n758 & n759;
  assign n761 = ~n612 & n760;
  assign n762 = ~n239 & n761;
  assign n763 = ~n501 & n762;
  assign n764 = n757 & n763;
  assign n765 = ~n393 & ~n454;
  assign n766 = ~n208 & n765;
  assign n767 = ~n198 & n766;
  assign n768 = ~n171 & ~n390;
  assign n769 = ~n161 & n768;
  assign n770 = ~n243 & n769;
  assign n771 = ~n621 & n770;
  assign n772 = n767 & n771;
  assign n773 = n764 & n772;
  assign n774 = n234 & n773;
  assign n775 = ~n391 & n774;
  assign n776 = ~n194 & n775;
  assign n777 = ~n150 & ~n206;
  assign n778 = ~n238 & n777;
  assign n779 = ~n383 & n778;
  assign n780 = n189 & n779;
  assign n781 = ~n614 & n780;
  assign n782 = ~n204 & n781;
  assign n783 = ~n473 & n782;
  assign n784 = n776 & n783;
  assign n785 = n752 & n784;
  assign n786 = n263 & n785;
  assign n787 = ~n78 & ~n395;
  assign n788 = ~n576 & ~n613;
  assign n789 = n418 & n788;
  assign n790 = n787 & n789;
  assign n791 = n786 & n790;
  assign n792 = ~n166 & n791;
  assign n793 = ~n193 & n792;
  assign n794 = n148 & n793;
  assign n795 = n737 & n794;
  assign n796 = ~n665 & ~n795;
  assign n797 = ~n463 & ~n547;
  assign n798 = n570 & n788;
  assign n799 = n797 & n798;
  assign n800 = ~n217 & n799;
  assign n801 = ~n232 & ~n534;
  assign n802 = ~n231 & ~n261;
  assign n803 = ~n461 & n802;
  assign n804 = n801 & n803;
  assign n805 = ~n354 & n804;
  assign n806 = ~n458 & n805;
  assign n807 = n276 & ~n580;
  assign n808 = ~n262 & ~n582;
  assign n809 = ~n361 & n808;
  assign n810 = ~n208 & n809;
  assign n811 = n807 & n810;
  assign n812 = ~n579 & n811;
  assign n813 = n806 & n812;
  assign n814 = ~n501 & ~n589;
  assign n815 = ~n350 & n814;
  assign n816 = ~n320 & ~n469;
  assign n817 = ~n395 & n816;
  assign n818 = ~n323 & n817;
  assign n819 = n815 & n818;
  assign n820 = ~n590 & n819;
  assign n821 = ~n170 & n820;
  assign n822 = n488 & ~n581;
  assign n823 = ~n342 & n822;
  assign n824 = ~n277 & n823;
  assign n825 = ~n163 & ~n372;
  assign n826 = n673 & n825;
  assign n827 = n824 & n826;
  assign n828 = ~n477 & n827;
  assign n829 = ~n218 & n828;
  assign n830 = n821 & n829;
  assign n831 = n813 & n830;
  assign n832 = n437 & n831;
  assign n833 = ~n465 & n832;
  assign n834 = n800 & n833;
  assign n835 = ~n595 & ~n681;
  assign n836 = ~n336 & n835;
  assign n837 = ~n147 & n836;
  assign n838 = ~n193 & ~n374;
  assign n839 = ~n279 & n838;
  assign n840 = ~n278 & n839;
  assign n841 = n837 & n840;
  assign n842 = n221 & n841;
  assign n843 = n476 & n842;
  assign n844 = ~n375 & n843;
  assign n845 = ~n242 & ~n280;
  assign n846 = ~n204 & n603;
  assign n847 = ~n337 & n846;
  assign n848 = n845 & n847;
  assign n849 = n257 & n848;
  assign n850 = ~n506 & n849;
  assign n851 = n844 & n850;
  assign n852 = ~n363 & ~n583;
  assign n853 = ~n341 & ~n667;
  assign n854 = n852 & n853;
  assign n855 = n777 & n854;
  assign n856 = ~n593 & n855;
  assign n857 = ~n214 & ~n668;
  assign n858 = ~n228 & ~n505;
  assign n859 = ~n588 & n858;
  assign n860 = ~n229 & ~n281;
  assign n861 = ~n504 & n860;
  assign n862 = ~n330 & ~n373;
  assign n863 = n861 & n862;
  assign n864 = ~n670 & n863;
  assign n865 = ~n598 & ~n693;
  assign n866 = ~n321 & n865;
  assign n867 = ~n473 & n866;
  assign n868 = n864 & n867;
  assign n869 = ~n669 & n868;
  assign n870 = ~n626 & n869;
  assign n871 = n859 & n870;
  assign n872 = n857 & n871;
  assign n873 = ~n594 & n872;
  assign n874 = ~n356 & n873;
  assign n875 = n856 & n874;
  assign n876 = n851 & n875;
  assign n877 = ~n152 & ~n427;
  assign n878 = ~n545 & n877;
  assign n879 = n876 & n878;
  assign n880 = ~n393 & n879;
  assign n881 = ~n272 & ~n548;
  assign n882 = ~n238 & ~n423;
  assign n883 = ~n243 & n882;
  assign n884 = ~n362 & ~n422;
  assign n885 = ~n188 & n884;
  assign n886 = ~n390 & ~n683;
  assign n887 = n885 & n886;
  assign n888 = ~n198 & n887;
  assign n889 = n883 & n888;
  assign n890 = n881 & n889;
  assign n891 = n327 & n890;
  assign n892 = ~n344 & n891;
  assign n893 = n880 & n892;
  assign n894 = n834 & n893;
  assign n895 = ~n795 & ~n894;
  assign n896 = ~n245 & ~n690;
  assign n897 = ~n435 & ~n594;
  assign n898 = n285 & n897;
  assign n899 = n896 & n898;
  assign n900 = ~n374 & n899;
  assign n901 = ~n599 & ~n610;
  assign n902 = n777 & n901;
  assign n903 = n156 & n902;
  assign n904 = ~n345 & n903;
  assign n905 = ~n357 & n904;
  assign n906 = n900 & n905;
  assign n907 = ~n601 & ~n701;
  assign n908 = ~n633 & n907;
  assign n909 = ~n195 & ~n639;
  assign n910 = ~n246 & ~n275;
  assign n911 = ~n260 & n910;
  assign n912 = n909 & n911;
  assign n913 = ~n293 & n912;
  assign n914 = ~n545 & n584;
  assign n915 = ~n627 & n914;
  assign n916 = n913 & n915;
  assign n917 = n908 & n916;
  assign n918 = n476 & n917;
  assign n919 = ~n232 & n918;
  assign n920 = ~n152 & ~n700;
  assign n921 = ~n360 & ~n682;
  assign n922 = ~n219 & n386;
  assign n923 = ~n477 & n922;
  assign n924 = n921 & n923;
  assign n925 = n920 & n924;
  assign n926 = ~n334 & n925;
  assign n927 = ~n501 & n926;
  assign n928 = n919 & n927;
  assign n929 = n906 & n928;
  assign n930 = ~n231 & ~n254;
  assign n931 = ~n578 & n930;
  assign n932 = ~n242 & n931;
  assign n933 = ~n314 & n932;
  assign n934 = ~n298 & ~n638;
  assign n935 = ~n261 & n934;
  assign n936 = ~n611 & n935;
  assign n937 = ~n165 & ~n424;
  assign n938 = n936 & n937;
  assign n939 = ~n294 & ~n307;
  assign n940 = ~n326 & n939;
  assign n941 = n938 & n940;
  assign n942 = n933 & n941;
  assign n943 = n929 & n942;
  assign n944 = n230 & n943;
  assign n945 = ~n395 & n944;
  assign n946 = ~n518 & ~n535;
  assign n947 = ~n290 & ~n325;
  assign n948 = ~n172 & n947;
  assign n949 = n857 & n948;
  assign n950 = n946 & n949;
  assign n951 = ~n217 & n950;
  assign n952 = ~n262 & n951;
  assign n953 = n945 & n952;
  assign n954 = ~n315 & ~n502;
  assign n955 = ~n147 & ~n308;
  assign n956 = ~n235 & ~n632;
  assign n957 = ~n304 & n956;
  assign n958 = ~n593 & n957;
  assign n959 = ~n218 & ~n332;
  assign n960 = ~n193 & n959;
  assign n961 = ~n180 & n960;
  assign n962 = ~n436 & n961;
  assign n963 = n958 & n962;
  assign n964 = n825 & n963;
  assign n965 = ~n220 & n964;
  assign n966 = ~n297 & ~n457;
  assign n967 = ~n505 & ~n679;
  assign n968 = ~n589 & n967;
  assign n969 = n797 & n968;
  assign n970 = n966 & n969;
  assign n971 = ~n614 & n970;
  assign n972 = ~n400 & n971;
  assign n973 = n965 & n972;
  assign n974 = ~n353 & ~n685;
  assign n975 = ~n631 & n816;
  assign n976 = ~n373 & n975;
  assign n977 = ~n273 & n976;
  assign n978 = n974 & n977;
  assign n979 = ~n678 & n978;
  assign n980 = ~n349 & ~n629;
  assign n981 = ~n383 & n980;
  assign n982 = ~n331 & n981;
  assign n983 = ~n213 & n982;
  assign n984 = n979 & n983;
  assign n985 = n973 & n984;
  assign n986 = ~n194 & ~n670;
  assign n987 = n467 & n986;
  assign n988 = ~n464 & n987;
  assign n989 = ~n239 & ~n413;
  assign n990 = ~n247 & n989;
  assign n991 = ~n381 & n990;
  assign n992 = n988 & n991;
  assign n993 = n985 & n992;
  assign n994 = n955 & n993;
  assign n995 = n954 & n994;
  assign n996 = ~n208 & n995;
  assign n997 = ~n204 & ~n462;
  assign n998 = ~n429 & ~n439;
  assign n999 = n540 & n998;
  assign n1000 = n788 & n999;
  assign n1001 = n997 & n1000;
  assign n1002 = ~n391 & n1001;
  assign n1003 = ~n442 & n1002;
  assign n1004 = n996 & n1003;
  assign n1005 = n953 & n1004;
  assign n1006 = ~n894 & ~n1005;
  assign n1007 = ~n228 & ~n638;
  assign n1008 = ~n463 & n1007;
  assign n1009 = n753 & n1008;
  assign n1010 = ~n299 & n1009;
  assign n1011 = ~n254 & ~n695;
  assign n1012 = ~n325 & ~n501;
  assign n1013 = ~n278 & ~n331;
  assign n1014 = ~n247 & n1013;
  assign n1015 = n1012 & n1014;
  assign n1016 = n1011 & n1015;
  assign n1017 = ~n147 & n1016;
  assign n1018 = n1010 & n1017;
  assign n1019 = n322 & n1018;
  assign n1020 = ~n163 & ~n533;
  assign n1021 = ~n461 & n1020;
  assign n1022 = ~n383 & ~n700;
  assign n1023 = n1021 & n1022;
  assign n1024 = ~n310 & ~n354;
  assign n1025 = ~n334 & ~n381;
  assign n1026 = n1024 & n1025;
  assign n1027 = ~n705 & n1026;
  assign n1028 = n1023 & n1027;
  assign n1029 = n1019 & n1028;
  assign n1030 = ~n580 & ~n697;
  assign n1031 = ~n413 & n1030;
  assign n1032 = ~n279 & n1031;
  assign n1033 = n1029 & n1032;
  assign n1034 = ~n436 & n1033;
  assign n1035 = ~n401 & n1034;
  assign n1036 = ~n598 & ~n704;
  assign n1037 = ~n360 & ~n385;
  assign n1038 = n1036 & n1037;
  assign n1039 = n226 & n1038;
  assign n1040 = ~n601 & n1039;
  assign n1041 = ~n309 & n1040;
  assign n1042 = ~n439 & n1041;
  assign n1043 = n1035 & n1042;
  assign n1044 = ~n134 & ~n375;
  assign n1045 = ~n171 & n1044;
  assign n1046 = ~n475 & n1045;
  assign n1047 = ~n238 & ~n517;
  assign n1048 = n1046 & n1047;
  assign n1049 = ~n581 & n1048;
  assign n1050 = ~n255 & ~n613;
  assign n1051 = ~n430 & n1050;
  assign n1052 = ~n161 & n1051;
  assign n1053 = ~n280 & n1052;
  assign n1054 = n1049 & n1053;
  assign n1055 = ~n337 & n1054;
  assign n1056 = ~n424 & n1055;
  assign n1057 = ~n273 & ~n361;
  assign n1058 = ~n232 & ~n423;
  assign n1059 = n1057 & n1058;
  assign n1060 = ~n576 & n1059;
  assign n1061 = ~n152 & n1060;
  assign n1062 = n1056 & n1061;
  assign n1063 = n237 & ~n305;
  assign n1064 = n558 & n1063;
  assign n1065 = ~n332 & n1064;
  assign n1066 = ~n537 & n1065;
  assign n1067 = n546 & ~n611;
  assign n1068 = ~n621 & ~n671;
  assign n1069 = ~n600 & n1068;
  assign n1070 = n1067 & n1069;
  assign n1071 = ~n679 & n1070;
  assign n1072 = ~n588 & n1071;
  assign n1073 = ~n356 & n1072;
  assign n1074 = n1066 & n1073;
  assign n1075 = n1062 & n1074;
  assign n1076 = ~n469 & ~n669;
  assign n1077 = ~n468 & n1076;
  assign n1078 = ~n464 & n1077;
  assign n1079 = ~n473 & ~n612;
  assign n1080 = ~n636 & n1079;
  assign n1081 = n1078 & n1080;
  assign n1082 = n1075 & n1081;
  assign n1083 = ~n637 & n1082;
  assign n1084 = ~n262 & n1083;
  assign n1085 = ~n678 & n1084;
  assign n1086 = ~n231 & ~n632;
  assign n1087 = ~n350 & n1086;
  assign n1088 = ~n628 & n1087;
  assign n1089 = ~n293 & ~n357;
  assign n1090 = ~n394 & ~n428;
  assign n1091 = ~n667 & n1090;
  assign n1092 = ~n330 & ~n353;
  assign n1093 = n1091 & n1092;
  assign n1094 = n1089 & n1093;
  assign n1095 = n1088 & n1094;
  assign n1096 = ~n288 & ~n534;
  assign n1097 = ~n631 & n901;
  assign n1098 = ~n229 & ~n502;
  assign n1099 = n1097 & n1098;
  assign n1100 = ~n536 & n1099;
  assign n1101 = n1096 & n1100;
  assign n1102 = n1095 & n1101;
  assign n1103 = ~n345 & n1102;
  assign n1104 = ~n462 & n1103;
  assign n1105 = ~n289 & n1104;
  assign n1106 = n1085 & n1105;
  assign n1107 = n1043 & n1106;
  assign n1108 = ~n1005 & ~n1107;
  assign n1109 = ~n461 & ~n536;
  assign n1110 = ~n375 & ~n637;
  assign n1111 = ~n243 & ~n350;
  assign n1112 = ~n116 & ~n310;
  assign n1113 = n1111 & n1112;
  assign n1114 = n1110 & n1113;
  assign n1115 = n1109 & n1114;
  assign n1116 = ~n219 & ~n595;
  assign n1117 = ~n166 & ~n183;
  assign n1118 = n1116 & n1117;
  assign n1119 = ~n147 & n1118;
  assign n1120 = ~n533 & ~n581;
  assign n1121 = ~n500 & n1120;
  assign n1122 = ~n289 & n1121;
  assign n1123 = n1119 & n1122;
  assign n1124 = ~n132 & ~n382;
  assign n1125 = ~n273 & ~n279;
  assign n1126 = ~n180 & n1125;
  assign n1127 = n1124 & n1126;
  assign n1128 = n1123 & n1127;
  assign n1129 = ~n475 & n1128;
  assign n1130 = n1115 & n1129;
  assign n1131 = ~n129 & ~n576;
  assign n1132 = ~n373 & ~n628;
  assign n1133 = ~n638 & n1132;
  assign n1134 = ~n188 & n1133;
  assign n1135 = n1131 & n1134;
  assign n1136 = n519 & n1135;
  assign n1137 = ~n231 & n1136;
  assign n1138 = ~n428 & ~n537;
  assign n1139 = ~n309 & ~n700;
  assign n1140 = ~n272 & n1139;
  assign n1141 = ~n154 & n1140;
  assign n1142 = n853 & n1141;
  assign n1143 = n1138 & n1142;
  assign n1144 = ~n259 & n1143;
  assign n1145 = n1137 & n1144;
  assign n1146 = n1130 & n1145;
  assign n1147 = ~n228 & ~n398;
  assign n1148 = ~n114 & ~n505;
  assign n1149 = ~n423 & n1148;
  assign n1150 = ~n672 & n1149;
  assign n1151 = n1147 & n1150;
  assign n1152 = n1146 & n1151;
  assign n1153 = ~n383 & ~n548;
  assign n1154 = ~n217 & ~n304;
  assign n1155 = ~n331 & n1154;
  assign n1156 = ~n324 & n1155;
  assign n1157 = n1153 & n1156;
  assign n1158 = n921 & n1157;
  assign n1159 = n1152 & n1158;
  assign n1160 = ~n299 & n1159;
  assign n1161 = ~n187 & n1160;
  assign n1162 = ~n204 & ~n611;
  assign n1163 = ~n463 & ~n477;
  assign n1164 = ~n504 & n1163;
  assign n1165 = ~n582 & n1164;
  assign n1166 = ~n260 & ~n261;
  assign n1167 = ~n193 & n1166;
  assign n1168 = n1165 & n1167;
  assign n1169 = ~n464 & ~n578;
  assign n1170 = n1050 & n1169;
  assign n1171 = ~n612 & n1170;
  assign n1172 = ~n195 & n1171;
  assign n1173 = ~n307 & ~n598;
  assign n1174 = ~n123 & n1173;
  assign n1175 = ~n356 & ~n391;
  assign n1176 = n101 & n1175;
  assign n1177 = n1012 & n1176;
  assign n1178 = n974 & n1177;
  assign n1179 = ~n614 & n1178;
  assign n1180 = ~n149 & ~n308;
  assign n1181 = ~n161 & ~n538;
  assign n1182 = ~n256 & ~n288;
  assign n1183 = n1181 & n1182;
  assign n1184 = n1180 & n1183;
  assign n1185 = n1179 & n1184;
  assign n1186 = ~n94 & ~n629;
  assign n1187 = n174 & ~n297;
  assign n1188 = ~n590 & n1187;
  assign n1189 = ~n198 & ~n385;
  assign n1190 = n1188 & n1189;
  assign n1191 = ~n414 & n1190;
  assign n1192 = ~n206 & ~n468;
  assign n1193 = ~n275 & n1192;
  assign n1194 = ~n422 & n1193;
  assign n1195 = ~n165 & n1194;
  assign n1196 = ~n181 & n1195;
  assign n1197 = n1191 & n1196;
  assign n1198 = n1186 & n1197;
  assign n1199 = ~n384 & n1198;
  assign n1200 = ~n208 & n467;
  assign n1201 = ~n186 & n852;
  assign n1202 = n1200 & n1201;
  assign n1203 = ~n232 & n1202;
  assign n1204 = ~n144 & ~n334;
  assign n1205 = ~n695 & n1204;
  assign n1206 = ~n704 & n1205;
  assign n1207 = n1203 & n1206;
  assign n1208 = ~n321 & n1207;
  assign n1209 = ~n689 & n1208;
  assign n1210 = n1199 & n1209;
  assign n1211 = n1185 & n1210;
  assign n1212 = ~n535 & n1211;
  assign n1213 = n1174 & n1212;
  assign n1214 = ~n294 & ~n506;
  assign n1215 = n488 & n1214;
  assign n1216 = n1213 & n1215;
  assign n1217 = n1172 & n1216;
  assign n1218 = n1168 & n1217;
  assign n1219 = n1162 & n1218;
  assign n1220 = ~n152 & ~n502;
  assign n1221 = ~n594 & n1220;
  assign n1222 = ~n336 & ~n454;
  assign n1223 = ~n214 & ~n424;
  assign n1224 = ~n374 & n1223;
  assign n1225 = n1222 & n1224;
  assign n1226 = n1221 & n1225;
  assign n1227 = ~n544 & n1226;
  assign n1228 = n1219 & n1227;
  assign n1229 = n694 & n1228;
  assign n1230 = n1161 & n1229;
  assign n1231 = ~n1107 & ~n1230;
  assign n1232 = ~n357 & ~n590;
  assign n1233 = ~n78 & ~n668;
  assign n1234 = ~n469 & n1233;
  assign n1235 = n343 & n1234;
  assign n1236 = n1232 & n1235;
  assign n1237 = ~n100 & n1236;
  assign n1238 = ~n315 & ~n578;
  assign n1239 = ~n217 & n1238;
  assign n1240 = ~n166 & n1239;
  assign n1241 = n244 & n1240;
  assign n1242 = n445 & n1241;
  assign n1243 = ~n466 & n1242;
  assign n1244 = ~n385 & n1243;
  assign n1245 = n1237 & n1244;
  assign n1246 = ~n614 & ~n692;
  assign n1247 = ~n331 & ~n637;
  assign n1248 = n703 & n1247;
  assign n1249 = n1181 & n1248;
  assign n1250 = n1246 & n1249;
  assign n1251 = ~n330 & n1250;
  assign n1252 = ~n122 & ~n548;
  assign n1253 = ~n114 & ~n475;
  assign n1254 = n1252 & n1253;
  assign n1255 = ~n462 & n1254;
  assign n1256 = ~n382 & n1255;
  assign n1257 = n1251 & n1256;
  assign n1258 = n1245 & n1257;
  assign n1259 = ~n290 & ~n320;
  assign n1260 = ~n214 & n1259;
  assign n1261 = ~n321 & n1260;
  assign n1262 = n1258 & n1261;
  assign n1263 = n306 & n1262;
  assign n1264 = ~n187 & n1263;
  assign n1265 = ~n81 & ~n422;
  assign n1266 = ~n464 & n528;
  assign n1267 = ~n180 & n1266;
  assign n1268 = ~n299 & ~n372;
  assign n1269 = ~n394 & n1268;
  assign n1270 = n1267 & n1269;
  assign n1271 = ~n399 & ~n588;
  assign n1272 = ~n435 & ~n667;
  assign n1273 = ~n252 & n1272;
  assign n1274 = ~n685 & n1273;
  assign n1275 = n1271 & n1274;
  assign n1276 = n1270 & n1275;
  assign n1277 = n1265 & n1276;
  assign n1278 = ~n206 & n1277;
  assign n1279 = ~n633 & n1278;
  assign n1280 = n1264 & n1279;
  assign n1281 = ~n173 & ~n427;
  assign n1282 = ~n104 & ~n611;
  assign n1283 = ~n203 & n1282;
  assign n1284 = ~n281 & ~n681;
  assign n1285 = ~n537 & ~n589;
  assign n1286 = ~n239 & n1285;
  assign n1287 = ~n401 & n1286;
  assign n1288 = n1284 & n1287;
  assign n1289 = ~n150 & n1288;
  assign n1290 = ~n194 & ~n232;
  assign n1291 = ~n129 & n1290;
  assign n1292 = ~n106 & n1291;
  assign n1293 = ~n627 & n1292;
  assign n1294 = ~n598 & n1293;
  assign n1295 = ~n213 & n1294;
  assign n1296 = n1289 & n1295;
  assign n1297 = n1283 & n1296;
  assign n1298 = n1281 & n1297;
  assign n1299 = ~n428 & n1298;
  assign n1300 = ~n458 & n1299;
  assign n1301 = ~n123 & ~n297;
  assign n1302 = ~n247 & ~n384;
  assign n1303 = ~n337 & n1302;
  assign n1304 = ~n98 & n1303;
  assign n1305 = ~n536 & n1304;
  assign n1306 = n1301 & n1305;
  assign n1307 = ~n704 & n1306;
  assign n1308 = ~n429 & n1307;
  assign n1309 = ~n632 & n1308;
  assign n1310 = n1300 & n1309;
  assign n1311 = ~n579 & ~n678;
  assign n1312 = ~n393 & n1311;
  assign n1313 = ~n583 & n1147;
  assign n1314 = ~n251 & n1313;
  assign n1315 = n1312 & n1314;
  assign n1316 = n1310 & n1315;
  assign n1317 = ~n261 & ~n349;
  assign n1318 = ~n324 & n1317;
  assign n1319 = ~n256 & ~n323;
  assign n1320 = ~n218 & n1319;
  assign n1321 = ~n457 & n1320;
  assign n1322 = ~n345 & n1321;
  assign n1323 = ~n154 & n1322;
  assign n1324 = ~n131 & n1323;
  assign n1325 = ~n395 & n1324;
  assign n1326 = ~n613 & n1325;
  assign n1327 = n1318 & n1326;
  assign n1328 = n1316 & n1327;
  assign n1329 = ~n229 & n1328;
  assign n1330 = ~n160 & n1329;
  assign n1331 = n376 & ~n636;
  assign n1332 = ~n599 & n1331;
  assign n1333 = n1204 & n1332;
  assign n1334 = n673 & n1333;
  assign n1335 = ~n235 & n1334;
  assign n1336 = ~n288 & n1335;
  assign n1337 = n1330 & n1336;
  assign n1338 = n1280 & n1337;
  assign n1339 = ~n1230 & ~n1338;
  assign n1340 = ~n98 & ~n464;
  assign n1341 = ~n85 & ~n132;
  assign n1342 = ~n336 & n1341;
  assign n1343 = ~n334 & ~n442;
  assign n1344 = ~n582 & ~n692;
  assign n1345 = n946 & n1344;
  assign n1346 = n1343 & n1345;
  assign n1347 = ~n186 & ~n637;
  assign n1348 = ~n341 & ~n429;
  assign n1349 = n1347 & n1348;
  assign n1350 = ~n672 & n1349;
  assign n1351 = n1346 & n1350;
  assign n1352 = ~n310 & ~n697;
  assign n1353 = ~n669 & n1352;
  assign n1354 = n1265 & n1353;
  assign n1355 = ~n100 & ~n307;
  assign n1356 = ~n399 & ~n474;
  assign n1357 = n1355 & n1356;
  assign n1358 = n1354 & n1357;
  assign n1359 = ~n689 & n1358;
  assign n1360 = n1351 & n1359;
  assign n1361 = n1342 & n1360;
  assign n1362 = ~n154 & ~n383;
  assign n1363 = ~n666 & n1362;
  assign n1364 = ~n259 & n1363;
  assign n1365 = ~n229 & n1364;
  assign n1366 = ~n299 & ~n583;
  assign n1367 = ~n129 & ~n690;
  assign n1368 = ~n198 & ~n314;
  assign n1369 = n215 & n1368;
  assign n1370 = ~n458 & n1369;
  assign n1371 = n1367 & n1370;
  assign n1372 = n1366 & n1371;
  assign n1373 = n1365 & n1372;
  assign n1374 = n1361 & n1373;
  assign n1375 = n1340 & n1374;
  assign n1376 = ~n374 & n511;
  assign n1377 = ~n633 & ~n678;
  assign n1378 = ~n626 & n1377;
  assign n1379 = n456 & n1378;
  assign n1380 = n1376 & n1379;
  assign n1381 = ~n682 & n706;
  assign n1382 = ~n290 & n1381;
  assign n1383 = n1192 & n1382;
  assign n1384 = n1380 & n1383;
  assign n1385 = n901 & n1384;
  assign n1386 = ~n245 & n1385;
  assign n1387 = n1375 & n1386;
  assign n1388 = ~n277 & ~n463;
  assign n1389 = ~n115 & ~n163;
  assign n1390 = ~n219 & ~n628;
  assign n1391 = n1389 & n1390;
  assign n1392 = n1388 & n1391;
  assign n1393 = ~n114 & n1392;
  assign n1394 = ~n131 & ~n297;
  assign n1395 = ~n393 & ~n698;
  assign n1396 = ~n150 & ~n262;
  assign n1397 = ~n345 & n1396;
  assign n1398 = n974 & n1397;
  assign n1399 = n1395 & n1398;
  assign n1400 = ~n668 & n1399;
  assign n1401 = ~n324 & ~n695;
  assign n1402 = ~n391 & ~n500;
  assign n1403 = n1401 & n1402;
  assign n1404 = ~n251 & n1403;
  assign n1405 = ~n181 & n1404;
  assign n1406 = n1400 & n1405;
  assign n1407 = ~n256 & n907;
  assign n1408 = ~n477 & n1407;
  assign n1409 = ~n323 & ~n465;
  assign n1410 = n910 & n1409;
  assign n1411 = n1086 & n1252;
  assign n1412 = n1410 & n1411;
  assign n1413 = ~n372 & n1412;
  assign n1414 = ~n579 & n1413;
  assign n1415 = n1408 & n1414;
  assign n1416 = n1406 & n1415;
  assign n1417 = ~n187 & ~n349;
  assign n1418 = ~n326 & ~n384;
  assign n1419 = ~n362 & n1418;
  assign n1420 = n1417 & n1419;
  assign n1421 = n1416 & n1420;
  assign n1422 = n1075 & n1421;
  assign n1423 = n1394 & n1422;
  assign n1424 = ~n439 & n1423;
  assign n1425 = n1393 & n1424;
  assign n1426 = n1387 & n1425;
  assign n1427 = ~n1338 & ~n1426;
  assign n1428 = ~n344 & ~n357;
  assign n1429 = ~n163 & n1428;
  assign n1430 = ~n275 & n1429;
  assign n1431 = ~n639 & n1430;
  assign n1432 = ~n116 & n1431;
  assign n1433 = ~n375 & n852;
  assign n1434 = ~n360 & n1433;
  assign n1435 = ~n129 & ~n636;
  assign n1436 = ~n458 & n1435;
  assign n1437 = ~n610 & n1436;
  assign n1438 = n1434 & n1437;
  assign n1439 = ~n465 & n1438;
  assign n1440 = n1432 & n1439;
  assign n1441 = ~n180 & ~n390;
  assign n1442 = ~n693 & n1441;
  assign n1443 = n1440 & n1442;
  assign n1444 = ~n100 & n1443;
  assign n1445 = ~n308 & n1109;
  assign n1446 = ~n242 & n1445;
  assign n1447 = ~n207 & ~n504;
  assign n1448 = ~n353 & ~n669;
  assign n1449 = n1447 & n1448;
  assign n1450 = ~n81 & n1449;
  assign n1451 = ~n173 & ~n517;
  assign n1452 = ~n600 & n1451;
  assign n1453 = ~n501 & n1452;
  assign n1454 = n1450 & n1453;
  assign n1455 = n1446 & n1454;
  assign n1456 = n997 & n1455;
  assign n1457 = ~n679 & n1456;
  assign n1458 = ~n231 & n1457;
  assign n1459 = n1444 & n1458;
  assign n1460 = ~n334 & n835;
  assign n1461 = ~n393 & n1460;
  assign n1462 = n546 & n1461;
  assign n1463 = ~n165 & n1462;
  assign n1464 = ~n307 & ~n593;
  assign n1465 = ~n468 & n491;
  assign n1466 = ~n246 & n1465;
  assign n1467 = n1222 & n1466;
  assign n1468 = n1464 & n1467;
  assign n1469 = n1268 & n1468;
  assign n1470 = ~n280 & n1469;
  assign n1471 = ~n309 & n779;
  assign n1472 = ~n293 & n1471;
  assign n1473 = ~n251 & n787;
  assign n1474 = n1472 & n1473;
  assign n1475 = n1394 & n1474;
  assign n1476 = ~n505 & n1475;
  assign n1477 = n1470 & n1476;
  assign n1478 = ~n245 & ~n288;
  assign n1479 = n184 & n447;
  assign n1480 = n1478 & n1479;
  assign n1481 = ~n535 & n1480;
  assign n1482 = ~n144 & ~n678;
  assign n1483 = ~n345 & ~n599;
  assign n1484 = ~n342 & n1483;
  assign n1485 = n1482 & n1484;
  assign n1486 = ~n469 & n1485;
  assign n1487 = ~n356 & n1486;
  assign n1488 = n1481 & n1487;
  assign n1489 = n1477 & n1488;
  assign n1490 = ~n310 & ~n427;
  assign n1491 = ~n601 & n1111;
  assign n1492 = ~n598 & n1491;
  assign n1493 = ~n506 & n1492;
  assign n1494 = ~n187 & ~n547;
  assign n1495 = ~n236 & n1220;
  assign n1496 = ~n218 & n1495;
  assign n1497 = ~n670 & n1496;
  assign n1498 = ~n629 & n1497;
  assign n1499 = ~n611 & n1498;
  assign n1500 = ~n362 & ~n435;
  assign n1501 = n1499 & n1500;
  assign n1502 = n1494 & n1501;
  assign n1503 = n1493 & n1502;
  assign n1504 = n1490 & n1503;
  assign n1505 = ~n188 & ~n671;
  assign n1506 = n386 & ~n638;
  assign n1507 = ~n194 & n1506;
  assign n1508 = n1505 & n1507;
  assign n1509 = n558 & n1508;
  assign n1510 = n1504 & n1509;
  assign n1511 = ~n117 & n1510;
  assign n1512 = ~n582 & n1511;
  assign n1513 = ~n94 & ~n477;
  assign n1514 = n1156 & n1513;
  assign n1515 = n1132 & n1514;
  assign n1516 = ~n332 & ~n534;
  assign n1517 = ~n323 & ~n442;
  assign n1518 = ~n527 & n1517;
  assign n1519 = ~n685 & n881;
  assign n1520 = ~n400 & n1519;
  assign n1521 = n1518 & n1520;
  assign n1522 = n1516 & n1521;
  assign n1523 = ~n213 & n1522;
  assign n1524 = n1515 & n1523;
  assign n1525 = n322 & n1524;
  assign n1526 = n1512 & n1525;
  assign n1527 = n1489 & n1526;
  assign n1528 = ~n422 & n1527;
  assign n1529 = ~n170 & n1528;
  assign n1530 = n1463 & n1529;
  assign n1531 = n1459 & n1530;
  assign n1532 = ~n1426 & ~n1531;
  assign n1533 = ~n194 & ~n320;
  assign n1534 = ~n193 & n1533;
  assign n1535 = n1362 & n1534;
  assign n1536 = n1131 & n1535;
  assign n1537 = n673 & n1536;
  assign n1538 = ~n170 & n1124;
  assign n1539 = ~n330 & ~n423;
  assign n1540 = ~n463 & n1539;
  assign n1541 = ~n375 & n1540;
  assign n1542 = ~n633 & n1541;
  assign n1543 = n1538 & n1542;
  assign n1544 = ~n85 & n1389;
  assign n1545 = ~n152 & ~n536;
  assign n1546 = n1513 & n1545;
  assign n1547 = ~n693 & n1546;
  assign n1548 = ~n106 & ~n598;
  assign n1549 = ~n682 & n1548;
  assign n1550 = ~n298 & n1549;
  assign n1551 = ~n398 & ~n527;
  assign n1552 = ~n629 & n1551;
  assign n1553 = ~n323 & n1552;
  assign n1554 = n1550 & n1553;
  assign n1555 = ~n304 & n1554;
  assign n1556 = ~n534 & n1555;
  assign n1557 = n1547 & n1556;
  assign n1558 = ~n502 & ~n701;
  assign n1559 = ~n466 & n1558;
  assign n1560 = ~n278 & ~n395;
  assign n1561 = n1559 & n1560;
  assign n1562 = n989 & n1561;
  assign n1563 = ~n342 & n1562;
  assign n1564 = ~n321 & n1563;
  assign n1565 = ~n455 & ~n626;
  assign n1566 = n415 & n1565;
  assign n1567 = ~n255 & n1566;
  assign n1568 = ~n259 & n1567;
  assign n1569 = n1564 & n1568;
  assign n1570 = n1557 & n1569;
  assign n1571 = n1544 & n1570;
  assign n1572 = n1543 & n1571;
  assign n1573 = ~n112 & n1572;
  assign n1574 = n1537 & n1573;
  assign n1575 = ~n314 & ~n690;
  assign n1576 = ~n436 & ~n621;
  assign n1577 = ~n203 & ~n683;
  assign n1578 = n814 & n1577;
  assign n1579 = ~n336 & n1578;
  assign n1580 = ~n337 & n1579;
  assign n1581 = ~n281 & ~n308;
  assign n1582 = ~n273 & ~n363;
  assign n1583 = n1272 & n1582;
  assign n1584 = n858 & n1583;
  assign n1585 = n1581 & n1584;
  assign n1586 = n615 & n1585;
  assign n1587 = ~n134 & ~n183;
  assign n1588 = ~n81 & ~n131;
  assign n1589 = n1587 & n1588;
  assign n1590 = ~n636 & n1589;
  assign n1591 = n1586 & n1590;
  assign n1592 = ~n147 & ~n254;
  assign n1593 = ~n583 & n1592;
  assign n1594 = ~n307 & n680;
  assign n1595 = ~n588 & n1594;
  assign n1596 = ~n475 & n1595;
  assign n1597 = ~n439 & n1596;
  assign n1598 = n1593 & n1597;
  assign n1599 = n1591 & n1598;
  assign n1600 = n1580 & n1599;
  assign n1601 = n1576 & n1600;
  assign n1602 = n1575 & n1601;
  assign n1603 = n1162 & n1602;
  assign n1604 = ~n229 & n1603;
  assign n1605 = ~n424 & ~n582;
  assign n1606 = n1197 & n1605;
  assign n1607 = n237 & n1606;
  assign n1608 = ~n309 & n1607;
  assign n1609 = n1604 & n1608;
  assign n1610 = n1574 & n1609;
  assign n1611 = ~n1531 & ~n1610;
  assign n1612 = ~n600 & n1565;
  assign n1613 = n1388 & n1612;
  assign n1614 = n402 & n1613;
  assign n1615 = ~n700 & n1614;
  assign n1616 = ~n537 & n1615;
  assign n1617 = ~n207 & ~n309;
  assign n1618 = ~n337 & ~n373;
  assign n1619 = n954 & n1618;
  assign n1620 = ~n132 & n1619;
  assign n1621 = ~n384 & n1620;
  assign n1622 = ~n588 & ~n695;
  assign n1623 = ~n422 & n1622;
  assign n1624 = ~n280 & ~n683;
  assign n1625 = ~n239 & n1624;
  assign n1626 = ~n693 & n1625;
  assign n1627 = n1623 & n1626;
  assign n1628 = ~n147 & ~n589;
  assign n1629 = ~n466 & n1628;
  assign n1630 = n1627 & n1629;
  assign n1631 = n1621 & n1630;
  assign n1632 = n1617 & n1631;
  assign n1633 = ~n681 & n1632;
  assign n1634 = ~n104 & ~n374;
  assign n1635 = ~n320 & ~n518;
  assign n1636 = n392 & n1635;
  assign n1637 = n1634 & n1636;
  assign n1638 = ~n594 & n1637;
  assign n1639 = ~n254 & n1638;
  assign n1640 = n1633 & n1639;
  assign n1641 = ~n229 & ~n593;
  assign n1642 = n1490 & n1641;
  assign n1643 = ~n144 & n1642;
  assign n1644 = ~n500 & ~n534;
  assign n1645 = ~n501 & n1644;
  assign n1646 = ~n163 & n1645;
  assign n1647 = n1234 & n1646;
  assign n1648 = ~n601 & n1647;
  assign n1649 = ~n582 & n1648;
  assign n1650 = n1643 & n1649;
  assign n1651 = n1640 & n1650;
  assign n1652 = ~n344 & ~n468;
  assign n1653 = ~n206 & n1652;
  assign n1654 = ~n349 & n1653;
  assign n1655 = ~n353 & n1654;
  assign n1656 = ~n208 & ~n213;
  assign n1657 = ~n666 & ~n698;
  assign n1658 = ~n117 & n1657;
  assign n1659 = ~n429 & ~n621;
  assign n1660 = n630 & n1659;
  assign n1661 = ~n477 & n1660;
  assign n1662 = n1658 & n1661;
  assign n1663 = n1656 & n1662;
  assign n1664 = n1655 & n1663;
  assign n1665 = n1651 & n1664;
  assign n1666 = ~n576 & n1665;
  assign n1667 = ~n228 & n1666;
  assign n1668 = ~n260 & n1667;
  assign n1669 = n1616 & n1668;
  assign n1670 = ~n331 & ~n356;
  assign n1671 = ~n332 & n1670;
  assign n1672 = ~n242 & ~n704;
  assign n1673 = n1671 & n1672;
  assign n1674 = ~n165 & n1673;
  assign n1675 = ~n361 & ~n638;
  assign n1676 = ~n115 & n1675;
  assign n1677 = ~n548 & n1676;
  assign n1678 = ~n214 & n1677;
  assign n1679 = n1674 & n1678;
  assign n1680 = n1126 & n1679;
  assign n1681 = n476 & n1680;
  assign n1682 = ~n430 & n1681;
  assign n1683 = n233 & ~n506;
  assign n1684 = ~n98 & ~n382;
  assign n1685 = ~n578 & n1684;
  assign n1686 = n1683 & n1685;
  assign n1687 = n1343 & n1686;
  assign n1688 = ~n428 & n1687;
  assign n1689 = n1682 & n1688;
  assign n1690 = ~n217 & n1377;
  assign n1691 = ~n538 & n1690;
  assign n1692 = ~n362 & n1691;
  assign n1693 = ~n171 & ~n395;
  assign n1694 = ~n441 & n1693;
  assign n1695 = ~n685 & n1694;
  assign n1696 = ~n307 & n1695;
  assign n1697 = ~n170 & n1696;
  assign n1698 = n189 & ~n345;
  assign n1699 = ~n272 & n1698;
  assign n1700 = ~n193 & ~n298;
  assign n1701 = ~n464 & n1700;
  assign n1702 = ~n81 & n1701;
  assign n1703 = n1699 & n1702;
  assign n1704 = ~n219 & n1703;
  assign n1705 = n1697 & n1704;
  assign n1706 = n1692 & n1705;
  assign n1707 = ~n305 & n1706;
  assign n1708 = ~n308 & ~n424;
  assign n1709 = ~n204 & n546;
  assign n1710 = ~n186 & n1709;
  assign n1711 = ~n262 & n1710;
  assign n1712 = n1708 & n1711;
  assign n1713 = ~n123 & n1712;
  assign n1714 = ~n670 & n1713;
  assign n1715 = n1707 & n1714;
  assign n1716 = n1689 & n1715;
  assign n1717 = ~n393 & n1587;
  assign n1718 = ~n360 & n1717;
  assign n1719 = ~n94 & n1718;
  assign n1720 = ~n278 & ~n385;
  assign n1721 = ~n375 & n1089;
  assign n1722 = n1720 & n1721;
  assign n1723 = ~n173 & ~n439;
  assign n1724 = ~n238 & ~n535;
  assign n1725 = n1723 & n1724;
  assign n1726 = n1722 & n1725;
  assign n1727 = n1120 & n1726;
  assign n1728 = n1719 & n1727;
  assign n1729 = n1716 & n1728;
  assign n1730 = ~n275 & n1729;
  assign n1731 = ~n194 & n1730;
  assign n1732 = ~n336 & ~n612;
  assign n1733 = ~n595 & n1732;
  assign n1734 = ~n682 & n1733;
  assign n1735 = ~n614 & n1734;
  assign n1736 = ~n504 & n1735;
  assign n1737 = ~n462 & n1736;
  assign n1738 = ~n671 & n1737;
  assign n1739 = n1731 & n1738;
  assign n1740 = n1669 & n1739;
  assign n1741 = ~n1610 & ~n1740;
  assign n1742 = ~n123 & ~n259;
  assign n1743 = ~n458 & n1742;
  assign n1744 = ~n293 & ~n632;
  assign n1745 = ~n423 & ~n590;
  assign n1746 = n1744 & n1745;
  assign n1747 = ~n220 & n1746;
  assign n1748 = n1743 & n1747;
  assign n1749 = ~n112 & ~n247;
  assign n1750 = ~n667 & n1749;
  assign n1751 = ~n611 & n1750;
  assign n1752 = ~n666 & n1751;
  assign n1753 = ~n474 & n1752;
  assign n1754 = ~n692 & n1753;
  assign n1755 = ~n304 & ~n600;
  assign n1756 = ~n81 & ~n583;
  assign n1757 = ~n401 & n1756;
  assign n1758 = ~n424 & n1757;
  assign n1759 = ~n315 & n1045;
  assign n1760 = ~n116 & n1759;
  assign n1761 = n1758 & n1760;
  assign n1762 = n1755 & n1761;
  assign n1763 = n1754 & n1762;
  assign n1764 = n1748 & n1763;
  assign n1765 = n1516 & n1764;
  assign n1766 = ~n441 & n1765;
  assign n1767 = ~n155 & ~n243;
  assign n1768 = n528 & n1767;
  assign n1769 = ~n537 & n1768;
  assign n1770 = n1353 & n1769;
  assign n1771 = n810 & n1770;
  assign n1772 = ~n578 & n1771;
  assign n1773 = ~n704 & n1772;
  assign n1774 = n1766 & n1773;
  assign n1775 = ~n422 & ~n689;
  assign n1776 = ~n701 & n797;
  assign n1777 = ~n290 & n1776;
  assign n1778 = ~n147 & n1777;
  assign n1779 = n1175 & n1778;
  assign n1780 = n1505 & n1779;
  assign n1781 = n1775 & n1780;
  assign n1782 = ~n115 & n1781;
  assign n1783 = ~n181 & ~n637;
  assign n1784 = ~n462 & ~n506;
  assign n1785 = ~n214 & ~n629;
  assign n1786 = n456 & n1785;
  assign n1787 = n1784 & n1786;
  assign n1788 = n1435 & n1787;
  assign n1789 = ~n354 & n1788;
  assign n1790 = ~n457 & n1789;
  assign n1791 = ~n439 & ~n500;
  assign n1792 = n1735 & n1791;
  assign n1793 = ~n154 & n1792;
  assign n1794 = ~n85 & n1793;
  assign n1795 = n1790 & n1794;
  assign n1796 = ~n705 & n1692;
  assign n1797 = ~n165 & n1796;
  assign n1798 = n491 & n1797;
  assign n1799 = n1445 & n1798;
  assign n1800 = ~n104 & n1799;
  assign n1801 = n868 & n1478;
  assign n1802 = ~n203 & n1801;
  assign n1803 = ~n218 & n1802;
  assign n1804 = n1800 & n1803;
  assign n1805 = n1795 & n1804;
  assign n1806 = n1783 & n1805;
  assign n1807 = n920 & n1806;
  assign n1808 = ~n363 & n1807;
  assign n1809 = ~n501 & n1808;
  assign n1810 = n1782 & n1809;
  assign n1811 = n1774 & n1810;
  assign n1812 = ~n1740 & ~n1811;
  assign n1813 = ~n170 & ~n670;
  assign n1814 = ~n621 & ~n689;
  assign n1815 = ~n310 & n1814;
  assign n1816 = ~n100 & n1815;
  assign n1817 = ~n204 & n1816;
  assign n1818 = n1271 & n1817;
  assign n1819 = ~n474 & n1818;
  assign n1820 = ~n537 & n1429;
  assign n1821 = ~n626 & n1820;
  assign n1822 = n1819 & n1821;
  assign n1823 = ~n256 & ~n273;
  assign n1824 = n233 & n1823;
  assign n1825 = ~n534 & n1824;
  assign n1826 = ~n247 & ~n390;
  assign n1827 = ~n197 & ~n350;
  assign n1828 = n1826 & n1827;
  assign n1829 = ~n147 & n1828;
  assign n1830 = ~n239 & ~n363;
  assign n1831 = ~n629 & n1830;
  assign n1832 = ~n155 & n1831;
  assign n1833 = ~n261 & n1832;
  assign n1834 = n1829 & n1833;
  assign n1835 = n1221 & n1834;
  assign n1836 = n1265 & n1835;
  assign n1837 = ~n117 & n1836;
  assign n1838 = ~n598 & n1837;
  assign n1839 = n1825 & n1838;
  assign n1840 = n1822 & n1839;
  assign n1841 = n1813 & n1840;
  assign n1842 = n1587 & n1841;
  assign n1843 = ~n590 & n1842;
  assign n1844 = ~n384 & ~n548;
  assign n1845 = ~n305 & n1844;
  assign n1846 = ~n166 & ~n171;
  assign n1847 = n1845 & n1846;
  assign n1848 = ~n277 & n1847;
  assign n1849 = ~n544 & n777;
  assign n1850 = ~n314 & n1849;
  assign n1851 = n1848 & n1850;
  assign n1852 = n1343 & n1851;
  assign n1853 = ~n455 & n1852;
  assign n1854 = n1281 & n1409;
  assign n1855 = n230 & n1854;
  assign n1856 = ~n375 & n1855;
  assign n1857 = ~n475 & n1856;
  assign n1858 = n1853 & n1857;
  assign n1859 = ~n112 & ~n243;
  assign n1860 = n1482 & n1859;
  assign n1861 = n1132 & n1860;
  assign n1862 = ~n436 & n1861;
  assign n1863 = ~n104 & ~n614;
  assign n1864 = ~n337 & n1863;
  assign n1865 = n1347 & n1864;
  assign n1866 = n684 & n1865;
  assign n1867 = ~n578 & n1866;
  assign n1868 = ~n214 & n1867;
  assign n1869 = n1862 & n1868;
  assign n1870 = n1858 & n1869;
  assign n1871 = ~n131 & n909;
  assign n1872 = ~n582 & ~n610;
  assign n1873 = ~n354 & ~n429;
  assign n1874 = n1872 & n1873;
  assign n1875 = ~n290 & n1874;
  assign n1876 = n1871 & n1875;
  assign n1877 = n1870 & n1876;
  assign n1878 = ~n149 & n1877;
  assign n1879 = n1843 & n1878;
  assign n1880 = ~n161 & n519;
  assign n1881 = ~n252 & ~n533;
  assign n1882 = ~n293 & ~n579;
  assign n1883 = n1881 & n1882;
  assign n1884 = ~n462 & n1883;
  assign n1885 = ~n430 & n488;
  assign n1886 = ~n275 & n1885;
  assign n1887 = ~n457 & n1886;
  assign n1888 = n1884 & n1887;
  assign n1889 = n1880 & n1888;
  assign n1890 = ~n506 & n1889;
  assign n1891 = ~n679 & n1109;
  assign n1892 = ~n262 & ~n681;
  assign n1893 = ~n613 & n1892;
  assign n1894 = ~n612 & n1893;
  assign n1895 = n1891 & n1894;
  assign n1896 = n908 & n1895;
  assign n1897 = n1791 & n1896;
  assign n1898 = ~n288 & n1897;
  assign n1899 = n1890 & n1898;
  assign n1900 = n1879 & n1899;
  assign n1901 = ~n1811 & ~n1900;
  assign n1902 = ~n194 & ~n545;
  assign n1903 = ~n701 & n1902;
  assign n1904 = ~n428 & n1903;
  assign n1905 = n1657 & n1904;
  assign n1906 = n415 & n1905;
  assign n1907 = ~n207 & n1906;
  assign n1908 = ~n427 & ~n580;
  assign n1909 = ~n217 & n1908;
  assign n1910 = ~n289 & n1909;
  assign n1911 = ~n279 & ~n613;
  assign n1912 = ~n260 & n1911;
  assign n1913 = ~n612 & n1912;
  assign n1914 = ~n116 & n1913;
  assign n1915 = n1910 & n1914;
  assign n1916 = ~n454 & n1915;
  assign n1917 = ~n172 & n396;
  assign n1918 = ~n401 & n1917;
  assign n1919 = ~n633 & ~n639;
  assign n1920 = ~n350 & n1919;
  assign n1921 = n1918 & n1920;
  assign n1922 = n1916 & n1921;
  assign n1923 = ~n381 & ~n457;
  assign n1924 = ~n323 & ~n423;
  assign n1925 = ~n390 & n1924;
  assign n1926 = n1770 & n1925;
  assign n1927 = ~n281 & n1926;
  assign n1928 = n1923 & n1927;
  assign n1929 = ~n275 & ~n598;
  assign n1930 = ~n413 & n1929;
  assign n1931 = ~n170 & n1930;
  assign n1932 = n897 & n1931;
  assign n1933 = n1565 & n1932;
  assign n1934 = ~n218 & ~n638;
  assign n1935 = ~n288 & ~n681;
  assign n1936 = ~n576 & n1935;
  assign n1937 = ~n466 & ~n579;
  assign n1938 = ~n374 & n1937;
  assign n1939 = ~n204 & n1938;
  assign n1940 = n1936 & n1939;
  assign n1941 = n1934 & n1940;
  assign n1942 = ~n362 & n1941;
  assign n1943 = n1933 & n1942;
  assign n1944 = ~n161 & n857;
  assign n1945 = ~n372 & n1944;
  assign n1946 = n1943 & n1945;
  assign n1947 = n1928 & n1946;
  assign n1948 = n1922 & n1947;
  assign n1949 = n797 & n1948;
  assign n1950 = ~n331 & n1949;
  assign n1951 = n1907 & n1950;
  assign n1952 = ~n693 & n1951;
  assign n1953 = ~n341 & ~n518;
  assign n1954 = ~n256 & n1953;
  assign n1955 = ~n236 & ~n538;
  assign n1956 = n1954 & n1955;
  assign n1957 = ~n383 & n1956;
  assign n1958 = ~n152 & ~n344;
  assign n1959 = n1957 & n1958;
  assign n1960 = ~n216 & n684;
  assign n1961 = ~n106 & n1960;
  assign n1962 = n1659 & n1961;
  assign n1963 = n1959 & n1962;
  assign n1964 = ~n117 & ~n375;
  assign n1965 = n253 & n1964;
  assign n1966 = ~n294 & n1965;
  assign n1967 = ~n477 & n1966;
  assign n1968 = ~n325 & ~n600;
  assign n1969 = ~n400 & n1968;
  assign n1970 = n1644 & n1969;
  assign n1971 = n1344 & n1970;
  assign n1972 = n558 & n1971;
  assign n1973 = ~n112 & n1972;
  assign n1974 = ~n599 & n1973;
  assign n1975 = n1967 & n1974;
  assign n1976 = ~n144 & ~n399;
  assign n1977 = ~n337 & n1976;
  assign n1978 = ~n186 & ~n430;
  assign n1979 = ~n171 & n1978;
  assign n1980 = n1977 & n1979;
  assign n1981 = ~n589 & n1980;
  assign n1982 = ~n361 & ~n627;
  assign n1983 = ~n297 & n1982;
  assign n1984 = ~n632 & n1983;
  assign n1985 = n1981 & n1984;
  assign n1986 = ~n246 & n1985;
  assign n1987 = ~n198 & n1986;
  assign n1988 = ~n220 & ~n636;
  assign n1989 = ~n363 & n1988;
  assign n1990 = ~n213 & ~n321;
  assign n1991 = ~n197 & n1990;
  assign n1992 = ~n517 & n1991;
  assign n1993 = n1989 & n1992;
  assign n1994 = n1109 & n1993;
  assign n1995 = ~n384 & n1994;
  assign n1996 = ~n187 & n1995;
  assign n1997 = n1987 & n1996;
  assign n1998 = n1975 & n1997;
  assign n1999 = ~n98 & ~n345;
  assign n2000 = ~n465 & n1999;
  assign n2001 = n263 & n2000;
  assign n2002 = n1998 & n2001;
  assign n2003 = n1963 & n2002;
  assign n2004 = ~n614 & n2003;
  assign n2005 = n1784 & n2004;
  assign n2006 = n1952 & n2005;
  assign n2007 = ~n1900 & ~n2006;
  assign n2008 = n1728 & n1947;
  assign n2009 = ~n611 & n797;
  assign n2010 = n1347 & n2009;
  assign n2011 = n896 & n2010;
  assign n2012 = ~n171 & n2011;
  assign n2013 = ~n106 & n2012;
  assign n2014 = n263 & n1545;
  assign n2015 = ~n689 & n2014;
  assign n2016 = ~n193 & n2015;
  assign n2017 = ~n610 & n2016;
  assign n2018 = n2013 & n2017;
  assign n2019 = n634 & n1686;
  assign n2020 = ~n475 & n2019;
  assign n2021 = ~n321 & ~n350;
  assign n2022 = n1664 & n2021;
  assign n2023 = ~n354 & n2022;
  assign n2024 = ~n172 & n2023;
  assign n2025 = ~n705 & n2024;
  assign n2026 = n2020 & n2025;
  assign n2027 = n2018 & n2026;
  assign n2028 = ~n298 & ~n534;
  assign n2029 = ~n672 & n2028;
  assign n2030 = n2027 & n2029;
  assign n2031 = n2008 & n2030;
  assign n2032 = ~n166 & ~n461;
  assign n2033 = ~n129 & ~n458;
  assign n2034 = n2032 & n2033;
  assign n2035 = ~n160 & n2034;
  assign n2036 = ~n198 & ~n342;
  assign n2037 = ~n220 & n2036;
  assign n2038 = ~n132 & n2037;
  assign n2039 = n2035 & n2038;
  assign n2040 = n2031 & n2039;
  assign n2041 = ~n78 & n2040;
  assign n2042 = ~n112 & ~n154;
  assign n2043 = ~n131 & n2042;
  assign n2044 = ~n582 & n1582;
  assign n2045 = n2043 & n2044;
  assign n2046 = ~n150 & ~n180;
  assign n2047 = ~n517 & n2046;
  assign n2048 = ~n474 & n2047;
  assign n2049 = n2045 & n2048;
  assign n2050 = n967 & n2049;
  assign n2051 = n1845 & n2050;
  assign n2052 = ~n235 & n2051;
  assign n2053 = ~n414 & n2052;
  assign n2054 = n2041 & n2053;
  assign n2055 = ~n391 & n2054;
  assign n2056 = ~n398 & ~n678;
  assign n2057 = ~n115 & n2056;
  assign n2058 = n2055 & n2057;
  assign n2059 = ~n2006 & ~n2058;
  assign n2060 = ~n639 & ~n689;
  assign n2061 = ~n666 & n2060;
  assign n2062 = ~n281 & n2061;
  assign n2063 = ~n384 & n2062;
  assign n2064 = ~n251 & ~n638;
  assign n2065 = ~n273 & ~n309;
  assign n2066 = ~n187 & ~n469;
  assign n2067 = ~n195 & n2066;
  assign n2068 = ~n242 & n2067;
  assign n2069 = n101 & n2068;
  assign n2070 = ~n326 & ~n401;
  assign n2071 = n1629 & n2070;
  assign n2072 = ~n500 & n694;
  assign n2073 = ~n207 & n2072;
  assign n2074 = n2071 & n2073;
  assign n2075 = n1694 & n2074;
  assign n2076 = n2069 & n2075;
  assign n2077 = n1908 & n2076;
  assign n2078 = n2065 & n2077;
  assign n2079 = n2064 & n2078;
  assign n2080 = ~n461 & n2079;
  assign n2081 = ~n354 & ~n690;
  assign n2082 = n1186 & n2081;
  assign n2083 = n1353 & n2082;
  assign n2084 = n1401 & n2083;
  assign n2085 = ~n122 & n2084;
  assign n2086 = ~n600 & n2085;
  assign n2087 = n2080 & n2086;
  assign n2088 = ~n474 & ~n544;
  assign n2089 = ~n413 & n1086;
  assign n2090 = n2088 & n2089;
  assign n2091 = ~n325 & ~n439;
  assign n2092 = ~n255 & n1265;
  assign n2093 = ~n166 & n2092;
  assign n2094 = n2091 & n2093;
  assign n2095 = n2090 & n2094;
  assign n2096 = ~n331 & n2095;
  assign n2097 = ~n88 & n2096;
  assign n2098 = n445 & ~n636;
  assign n2099 = ~n614 & n2098;
  assign n2100 = n291 & n2099;
  assign n2101 = ~n155 & n2100;
  assign n2102 = ~n598 & n2101;
  assign n2103 = n2097 & n2102;
  assign n2104 = n2087 & n2103;
  assign n2105 = ~n277 & ~n705;
  assign n2106 = n364 & n2105;
  assign n2107 = n797 & n2106;
  assign n2108 = n2104 & n2107;
  assign n2109 = ~n611 & n2108;
  assign n2110 = ~n134 & n2109;
  assign n2111 = ~n314 & ~n501;
  assign n2112 = ~n259 & n2111;
  assign n2113 = ~n262 & n2112;
  assign n2114 = ~n170 & ~n360;
  assign n2115 = ~n400 & n2114;
  assign n2116 = ~n428 & n2115;
  assign n2117 = ~n213 & ~n332;
  assign n2118 = n2116 & n2117;
  assign n2119 = n1924 & n2118;
  assign n2120 = n2113 & n2119;
  assign n2121 = n1708 & n2120;
  assign n2122 = ~n334 & n2121;
  assign n2123 = ~n78 & ~n536;
  assign n2124 = ~n385 & n2123;
  assign n2125 = ~n218 & ~n398;
  assign n2126 = ~n149 & n2125;
  assign n2127 = n2124 & n2126;
  assign n2128 = ~n701 & n2127;
  assign n2129 = ~n583 & n2128;
  assign n2130 = n2122 & n2129;
  assign n2131 = ~n337 & ~n590;
  assign n2132 = ~n235 & ~n238;
  assign n2133 = ~n275 & n2132;
  assign n2134 = n2131 & n2133;
  assign n2135 = ~n599 & n2134;
  assign n2136 = ~n186 & n1079;
  assign n2137 = ~n203 & ~n668;
  assign n2138 = ~n154 & n2137;
  assign n2139 = ~n116 & ~n436;
  assign n2140 = ~n272 & n2139;
  assign n2141 = ~n631 & n2140;
  assign n2142 = ~n353 & n2141;
  assign n2143 = n2138 & n2142;
  assign n2144 = n2136 & n2143;
  assign n2145 = ~n578 & n2144;
  assign n2146 = ~n341 & n2145;
  assign n2147 = n2135 & n2146;
  assign n2148 = n2130 & n2147;
  assign n2149 = ~n393 & ~n504;
  assign n2150 = n673 & n2149;
  assign n2151 = ~n435 & n2150;
  assign n2152 = ~n115 & ~n345;
  assign n2153 = ~n373 & n2152;
  assign n2154 = ~n588 & n2153;
  assign n2155 = ~n344 & n2154;
  assign n2156 = n2151 & n2155;
  assign n2157 = n596 & n2156;
  assign n2158 = ~n545 & n1192;
  assign n2159 = ~n304 & n2158;
  assign n2160 = ~n455 & n1700;
  assign n2161 = ~n667 & n2160;
  assign n2162 = n2159 & n2161;
  assign n2163 = ~n144 & ~n414;
  assign n2164 = ~n245 & n2163;
  assign n2165 = ~n163 & ~n228;
  assign n2166 = ~n256 & n2165;
  assign n2167 = ~n243 & n2166;
  assign n2168 = ~n621 & n2167;
  assign n2169 = n2164 & n2168;
  assign n2170 = n2162 & n2169;
  assign n2171 = n1637 & n2170;
  assign n2172 = n2157 & n2171;
  assign n2173 = n2148 & n2172;
  assign n2174 = ~n252 & n2173;
  assign n2175 = ~n534 & n2174;
  assign n2176 = n2110 & n2175;
  assign n2177 = ~n194 & n2176;
  assign n2178 = n2063 & n2177;
  assign n2179 = ~n2058 & ~n2178;
  assign n2180 = ~n414 & ~n442;
  assign n2181 = ~n464 & n2060;
  assign n2182 = n1924 & n1991;
  assign n2183 = ~n104 & ~n308;
  assign n2184 = ~n116 & n2183;
  assign n2185 = n174 & n2184;
  assign n2186 = n1784 & n2185;
  assign n2187 = n2182 & n2186;
  assign n2188 = ~n612 & n2187;
  assign n2189 = n392 & n592;
  assign n2190 = ~n171 & n2189;
  assign n2191 = ~n294 & ~n685;
  assign n2192 = ~n207 & ~n430;
  assign n2193 = ~n342 & n2192;
  assign n2194 = ~n131 & n2193;
  assign n2195 = ~n203 & ~n401;
  assign n2196 = n1964 & n2195;
  assign n2197 = ~n669 & n2048;
  assign n2198 = n2196 & n2197;
  assign n2199 = ~n382 & ~n579;
  assign n2200 = ~n670 & n2199;
  assign n2201 = ~n436 & n2200;
  assign n2202 = n2198 & n2201;
  assign n2203 = n2194 & n2202;
  assign n2204 = n2191 & n2203;
  assign n2205 = ~n373 & n2204;
  assign n2206 = ~n132 & n2205;
  assign n2207 = n2190 & n2206;
  assign n2208 = n2188 & n2207;
  assign n2209 = n2181 & n2208;
  assign n2210 = n528 & n2209;
  assign n2211 = ~n228 & n2210;
  assign n2212 = n2180 & n2211;
  assign n2213 = ~n144 & n2212;
  assign n2214 = ~n357 & ~n580;
  assign n2215 = ~n235 & n2214;
  assign n2216 = n1613 & n2215;
  assign n2217 = ~n697 & n2216;
  assign n2218 = ~n188 & ~n690;
  assign n2219 = ~n500 & n2218;
  assign n2220 = ~n112 & n2219;
  assign n2221 = ~n85 & ~n705;
  assign n2222 = n2220 & n2221;
  assign n2223 = n156 & n2222;
  assign n2224 = n1923 & n2223;
  assign n2225 = ~n147 & n2224;
  assign n2226 = n2217 & n2225;
  assign n2227 = ~n336 & n2226;
  assign n2228 = n306 & ~n683;
  assign n2229 = ~n395 & n2228;
  assign n2230 = n825 & n2229;
  assign n2231 = ~n252 & ~n631;
  assign n2232 = ~n259 & ~n594;
  assign n2233 = ~n533 & n2232;
  assign n2234 = ~n349 & n2233;
  assign n2235 = n2231 & n2234;
  assign n2236 = n2230 & n2235;
  assign n2237 = ~n217 & n2236;
  assign n2238 = n2056 & n2237;
  assign n2239 = n2227 & n2238;
  assign n2240 = ~n413 & ~n504;
  assign n2241 = ~n439 & n2240;
  assign n2242 = ~n362 & n2241;
  assign n2243 = n2239 & n2242;
  assign n2244 = ~n595 & n2243;
  assign n2245 = ~n344 & n2244;
  assign n2246 = n2213 & n2245;
  assign n2247 = ~n242 & ~n679;
  assign n2248 = ~n238 & n2247;
  assign n2249 = n1253 & n2248;
  assign n2250 = n1186 & n2249;
  assign n2251 = ~n208 & n2250;
  assign n2252 = n257 & ~n354;
  assign n2253 = ~n356 & n2252;
  assign n2254 = ~n288 & ~n518;
  assign n2255 = ~n260 & n2254;
  assign n2256 = ~n345 & n2255;
  assign n2257 = ~n231 & ~n610;
  assign n2258 = n2256 & n2257;
  assign n2259 = ~n181 & ~n545;
  assign n2260 = ~n290 & n2259;
  assign n2261 = n2258 & n2260;
  assign n2262 = n2253 & n2261;
  assign n2263 = ~n698 & n1720;
  assign n2264 = ~n239 & n2263;
  assign n2265 = ~n229 & ~n279;
  assign n2266 = ~n98 & n2265;
  assign n2267 = n2264 & n2266;
  assign n2268 = ~n477 & n2267;
  assign n2269 = ~n195 & ~n667;
  assign n2270 = ~n204 & n1301;
  assign n2271 = ~n424 & n2270;
  assign n2272 = n2269 & n2271;
  assign n2273 = n2268 & n2272;
  assign n2274 = n2262 & n2273;
  assign n2275 = ~n337 & n2274;
  assign n2276 = ~n216 & n2275;
  assign n2277 = n2251 & n2276;
  assign n2278 = n2246 & n2277;
  assign n2279 = ~n2178 & ~n2278;
  assign n2280 = ~n383 & ~n697;
  assign n2281 = ~n251 & ~n595;
  assign n2282 = ~n166 & ~n393;
  assign n2283 = n2281 & n2282;
  assign n2284 = ~n272 & n2283;
  assign n2285 = n237 & n907;
  assign n2286 = n2284 & n2285;
  assign n2287 = n1302 & n2286;
  assign n2288 = n2280 & n2287;
  assign n2289 = ~n670 & n2288;
  assign n2290 = ~n279 & ~n293;
  assign n2291 = ~n506 & n2290;
  assign n2292 = n753 & n2291;
  assign n2293 = ~n590 & n2292;
  assign n2294 = ~n315 & ~n361;
  assign n2295 = n416 & n2294;
  assign n2296 = ~n299 & n2295;
  assign n2297 = ~n668 & n2296;
  assign n2298 = n2293 & n2297;
  assign n2299 = ~n154 & ~n354;
  assign n2300 = ~n197 & ~n297;
  assign n2301 = ~n255 & n2300;
  assign n2302 = ~n391 & n2301;
  assign n2303 = n2299 & n2302;
  assign n2304 = ~n454 & n2303;
  assign n2305 = ~n149 & ~n350;
  assign n2306 = n2304 & n2305;
  assign n2307 = ~n171 & n2306;
  assign n2308 = ~n461 & n2307;
  assign n2309 = ~n385 & ~n695;
  assign n2310 = ~n441 & n2222;
  assign n2311 = n2309 & n2310;
  assign n2312 = ~n216 & n2311;
  assign n2313 = ~n123 & n1356;
  assign n2314 = ~n170 & n2313;
  assign n2315 = ~n261 & n2314;
  assign n2316 = n2312 & n2315;
  assign n2317 = n119 & n2316;
  assign n2318 = ~n398 & n2317;
  assign n2319 = n2308 & n2318;
  assign n2320 = n2298 & n2319;
  assign n2321 = ~n217 & ~n477;
  assign n2322 = n2320 & n2321;
  assign n2323 = n2231 & n2322;
  assign n2324 = ~n325 & n2323;
  assign n2325 = n2289 & n2324;
  assign n2326 = ~n229 & n921;
  assign n2327 = ~n94 & n2326;
  assign n2328 = n396 & n2327;
  assign n2329 = n2136 & n2328;
  assign n2330 = n673 & n2329;
  assign n2331 = ~n183 & n2330;
  assign n2332 = ~n207 & ~n332;
  assign n2333 = ~n172 & n2332;
  assign n2334 = ~n517 & n2333;
  assign n2335 = ~n462 & n2334;
  assign n2336 = n2199 & n2335;
  assign n2337 = ~n314 & n2336;
  assign n2338 = ~n505 & n2337;
  assign n2339 = n2331 & n2338;
  assign n2340 = ~n336 & ~n693;
  assign n2341 = n467 & n1934;
  assign n2342 = ~n538 & n2341;
  assign n2343 = n1494 & n2342;
  assign n2344 = n2340 & n2343;
  assign n2345 = ~n246 & ~n337;
  assign n2346 = n1670 & n2170;
  assign n2347 = n2345 & n2346;
  assign n2348 = n1396 & n2347;
  assign n2349 = n2344 & n2348;
  assign n2350 = n2339 & n2349;
  assign n2351 = ~n104 & ~n372;
  assign n2352 = ~n401 & n2351;
  assign n2353 = ~n700 & n2352;
  assign n2354 = ~n375 & n1872;
  assign n2355 = ~n429 & n2354;
  assign n2356 = ~n129 & ~n626;
  assign n2357 = ~n181 & n2356;
  assign n2358 = n2355 & n2357;
  assign n2359 = ~n628 & n2358;
  assign n2360 = n2353 & n2359;
  assign n2361 = n2350 & n2360;
  assign n2362 = n1252 & n2361;
  assign n2363 = ~n435 & n2362;
  assign n2364 = ~n536 & ~n629;
  assign n2365 = ~n324 & n2364;
  assign n2366 = n1598 & n2365;
  assign n2367 = n882 & n2366;
  assign n2368 = n2363 & n2367;
  assign n2369 = n2325 & n2368;
  assign n2370 = ~n2278 & ~n2369;
  assign n2371 = ~n115 & ~n203;
  assign n2372 = ~n698 & n2371;
  assign n2373 = ~n435 & ~n631;
  assign n2374 = ~n474 & n2373;
  assign n2375 = n2372 & n2374;
  assign n2376 = n1705 & n2375;
  assign n2377 = n1192 & n2376;
  assign n2378 = ~n477 & n2377;
  assign n2379 = ~n251 & ~n469;
  assign n2380 = ~n236 & n2379;
  assign n2381 = n1147 & n2380;
  assign n2382 = n1388 & n2381;
  assign n2383 = ~n122 & n2382;
  assign n2384 = n416 & n1708;
  assign n2385 = ~n589 & n2384;
  assign n2386 = n2383 & n2385;
  assign n2387 = n1138 & n2201;
  assign n2388 = ~n582 & n2387;
  assign n2389 = ~n372 & n920;
  assign n2390 = ~n439 & n2389;
  assign n2391 = n967 & n2390;
  assign n2392 = n402 & ~n527;
  assign n2393 = ~n614 & n2392;
  assign n2394 = n1353 & n2393;
  assign n2395 = n562 & n2394;
  assign n2396 = n2391 & n2395;
  assign n2397 = n1057 & n2396;
  assign n2398 = ~n613 & n2397;
  assign n2399 = n2388 & n2398;
  assign n2400 = n2386 & n2399;
  assign n2401 = ~n314 & ~n629;
  assign n2402 = ~n260 & n2401;
  assign n2403 = ~n256 & n2402;
  assign n2404 = n2400 & n2403;
  assign n2405 = n291 & n2404;
  assign n2406 = ~n229 & n2405;
  assign n2407 = ~n242 & n2406;
  assign n2408 = n2378 & n2407;
  assign n2409 = ~n255 & ~n666;
  assign n2410 = ~n336 & n694;
  assign n2411 = ~n154 & n2410;
  assign n2412 = n2409 & n2411;
  assign n2413 = n1011 & n2412;
  assign n2414 = ~n548 & n2413;
  assign n2415 = ~n536 & n2414;
  assign n2416 = ~n576 & n1516;
  assign n2417 = ~n132 & ~n208;
  assign n2418 = ~n238 & ~n705;
  assign n2419 = ~n595 & n2418;
  assign n2420 = ~n326 & n2419;
  assign n2421 = ~n462 & n2420;
  assign n2422 = ~n304 & n2421;
  assign n2423 = ~n414 & ~n610;
  assign n2424 = ~n239 & n2423;
  assign n2425 = ~n504 & n1409;
  assign n2426 = ~n518 & n2425;
  assign n2427 = ~n601 & ~n621;
  assign n2428 = ~n172 & ~n197;
  assign n2429 = ~n131 & ~n363;
  assign n2430 = n2428 & n2429;
  assign n2431 = n2427 & n2430;
  assign n2432 = n2426 & n2431;
  assign n2433 = n2424 & n2432;
  assign n2434 = ~n194 & n2433;
  assign n2435 = ~n114 & n2434;
  assign n2436 = ~n261 & ~n501;
  assign n2437 = ~n281 & n2436;
  assign n2438 = ~n88 & ~n547;
  assign n2439 = ~n129 & n2438;
  assign n2440 = n2437 & n2439;
  assign n2441 = ~n213 & ~n690;
  assign n2442 = ~n94 & n2441;
  assign n2443 = ~n166 & ~n683;
  assign n2444 = n2442 & n2443;
  assign n2445 = n2440 & n2444;
  assign n2446 = ~n117 & n2445;
  assign n2447 = ~n393 & n2446;
  assign n2448 = ~n632 & n2447;
  assign n2449 = n2435 & n2448;
  assign n2450 = ~n147 & n2449;
  assign n2451 = n2422 & n2450;
  assign n2452 = n2417 & n2451;
  assign n2453 = n1110 & n2452;
  assign n2454 = n2416 & n2453;
  assign n2455 = ~n394 & n2454;
  assign n2456 = n2415 & n2455;
  assign n2457 = n2408 & n2456;
  assign n2458 = ~n2369 & ~n2457;
  assign n2459 = ~n279 & ~n310;
  assign n2460 = ~n239 & n2459;
  assign n2461 = ~n106 & n2460;
  assign n2462 = ~n152 & ~n533;
  assign n2463 = n2461 & n2462;
  assign n2464 = n1652 & n2463;
  assign n2465 = n673 & n2464;
  assign n2466 = ~n475 & n2465;
  assign n2467 = ~n207 & ~n463;
  assign n2468 = ~n474 & n2427;
  assign n2469 = ~n204 & n2468;
  assign n2470 = n966 & n2469;
  assign n2471 = n2467 & n2470;
  assign n2472 = n135 & n2471;
  assign n2473 = ~n242 & n2472;
  assign n2474 = ~n281 & ~n422;
  assign n2475 = n2256 & n2474;
  assign n2476 = ~n289 & n2475;
  assign n2477 = ~n598 & n2476;
  assign n2478 = n2473 & n2477;
  assign n2479 = n748 & n1343;
  assign n2480 = ~n613 & n2479;
  assign n2481 = ~n627 & ~n682;
  assign n2482 = ~n161 & ~n639;
  assign n2483 = ~n94 & n2482;
  assign n2484 = n2481 & n2483;
  assign n2485 = ~n375 & n2484;
  assign n2486 = ~n259 & n2485;
  assign n2487 = n2480 & n2486;
  assign n2488 = n2478 & n2487;
  assign n2489 = ~n123 & n1902;
  assign n2490 = ~n332 & n2489;
  assign n2491 = ~n78 & ~n670;
  assign n2492 = n1095 & n2491;
  assign n2493 = ~n581 & n2492;
  assign n2494 = ~n100 & ~n216;
  assign n2495 = ~n326 & ~n361;
  assign n2496 = ~n219 & n2495;
  assign n2497 = n1656 & n2496;
  assign n2498 = n2494 & n2497;
  assign n2499 = ~n349 & n2498;
  assign n2500 = n2493 & n2499;
  assign n2501 = ~n122 & n2500;
  assign n2502 = ~n275 & ~n633;
  assign n2503 = ~n188 & n2502;
  assign n2504 = ~n307 & n2503;
  assign n2505 = ~n114 & ~n217;
  assign n2506 = n1767 & n2505;
  assign n2507 = ~n506 & n2506;
  assign n2508 = ~n252 & n2365;
  assign n2509 = ~n112 & n2508;
  assign n2510 = n2507 & n2509;
  assign n2511 = ~n669 & n2510;
  assign n2512 = ~n218 & n1723;
  assign n2513 = ~n538 & n1733;
  assign n2514 = ~n610 & n2513;
  assign n2515 = n2512 & n2514;
  assign n2516 = n2511 & n2515;
  assign n2517 = ~n116 & ~n414;
  assign n2518 = ~n165 & n2517;
  assign n2519 = ~n280 & ~n600;
  assign n2520 = n2518 & n2519;
  assign n2521 = n2516 & n2520;
  assign n2522 = ~n198 & n2521;
  assign n2523 = n2504 & n2522;
  assign n2524 = n2501 & n2523;
  assign n2525 = ~n685 & n2524;
  assign n2526 = ~n535 & n2525;
  assign n2527 = n2490 & n2526;
  assign n2528 = ~n441 & n2527;
  assign n2529 = ~n193 & ~n427;
  assign n2530 = ~n679 & n2131;
  assign n2531 = ~n232 & n2530;
  assign n2532 = n2529 & n2531;
  assign n2533 = n2528 & n2532;
  assign n2534 = n2488 & n2533;
  assign n2535 = ~n180 & n2534;
  assign n2536 = ~n678 & n2535;
  assign n2537 = n2466 & n2536;
  assign n2538 = ~n235 & ~n527;
  assign n2539 = ~n395 & n2538;
  assign n2540 = ~n704 & n2539;
  assign n2541 = ~n88 & n2540;
  assign n2542 = ~n626 & n2166;
  assign n2543 = n2541 & n2542;
  assign n2544 = n1605 & n2543;
  assign n2545 = ~n363 & n2544;
  assign n2546 = ~n220 & n2545;
  assign n2547 = n437 & ~n638;
  assign n2548 = ~n689 & n2547;
  assign n2549 = n699 & n2548;
  assign n2550 = n896 & n2549;
  assign n2551 = ~n458 & n2550;
  assign n2552 = ~n469 & n2551;
  assign n2553 = n2546 & n2552;
  assign n2554 = n2537 & n2553;
  assign n2555 = ~n2457 & ~n2554;
  assign n2556 = ~n85 & ~n362;
  assign n2557 = ~n188 & n2556;
  assign n2558 = n1657 & n2557;
  assign n2559 = n445 & n2558;
  assign n2560 = n907 & n2559;
  assign n2561 = ~n679 & n2560;
  assign n2562 = ~n154 & n1784;
  assign n2563 = ~n436 & n2562;
  assign n2564 = n2459 & n2563;
  assign n2565 = n162 & ~n342;
  assign n2566 = ~n382 & ~n600;
  assign n2567 = ~n288 & n2566;
  assign n2568 = ~n331 & n2567;
  assign n2569 = n2565 & n2568;
  assign n2570 = n807 & n2569;
  assign n2571 = n2564 & n2570;
  assign n2572 = ~n220 & ~n589;
  assign n2573 = ~n477 & ~n638;
  assign n2574 = ~n345 & n2573;
  assign n2575 = ~n305 & n2574;
  assign n2576 = n2572 & n2575;
  assign n2577 = n2571 & n2576;
  assign n2578 = n467 & n2577;
  assign n2579 = n1435 & n2578;
  assign n2580 = ~n474 & n2579;
  assign n2581 = n2561 & n2580;
  assign n2582 = ~n294 & n1162;
  assign n2583 = ~n353 & n2582;
  assign n2584 = ~n187 & n2583;
  assign n2585 = ~n208 & ~n427;
  assign n2586 = ~n252 & n2585;
  assign n2587 = ~n461 & n2586;
  assign n2588 = ~n289 & ~n334;
  assign n2589 = n2494 & n2588;
  assign n2590 = ~n213 & n2589;
  assign n2591 = n2587 & n2590;
  assign n2592 = ~n505 & n2591;
  assign n2593 = n2584 & n2592;
  assign n2594 = n1076 & n2593;
  assign n2595 = n1232 & n2594;
  assign n2596 = ~n235 & n2595;
  assign n2597 = n787 & n1635;
  assign n2598 = ~n690 & n2597;
  assign n2599 = ~n308 & n2598;
  assign n2600 = n2596 & n2599;
  assign n2601 = n754 & n1138;
  assign n2602 = ~n207 & n2601;
  assign n2603 = ~n321 & n909;
  assign n2604 = ~n172 & n838;
  assign n2605 = ~n588 & n2604;
  assign n2606 = ~n704 & n2605;
  assign n2607 = n2603 & n2606;
  assign n2608 = ~n594 & n2607;
  assign n2609 = ~n612 & n2608;
  assign n2610 = n2602 & n2609;
  assign n2611 = n2600 & n2610;
  assign n2612 = ~n501 & n2611;
  assign n2613 = ~n228 & n2612;
  assign n2614 = n107 & n2613;
  assign n2615 = ~n122 & n2614;
  assign n2616 = ~n473 & ~n671;
  assign n2617 = n1301 & n1451;
  assign n2618 = ~n500 & n2617;
  assign n2619 = ~n349 & n2618;
  assign n2620 = ~n290 & ~n309;
  assign n2621 = ~n293 & n2620;
  assign n2622 = ~n336 & n2621;
  assign n2623 = ~n219 & n2622;
  assign n2624 = n777 & n2623;
  assign n2625 = ~n613 & n2624;
  assign n2626 = ~n251 & n2625;
  assign n2627 = n2619 & n2626;
  assign n2628 = ~n373 & n1834;
  assign n2629 = ~n203 & ~n547;
  assign n2630 = ~n583 & n2629;
  assign n2631 = n546 & n2630;
  assign n2632 = ~n633 & n2631;
  assign n2633 = n2628 & n2632;
  assign n2634 = n2627 & n2633;
  assign n2635 = n2616 & n2634;
  assign n2636 = n1270 & n2635;
  assign n2637 = n1892 & n2636;
  assign n2638 = ~n341 & n2637;
  assign n2639 = n2615 & n2638;
  assign n2640 = n2581 & n2639;
  assign n2641 = ~n2554 & ~n2640;
  assign n2642 = ~n278 & ~n601;
  assign n2643 = ~n356 & n2642;
  assign n2644 = n615 & n2643;
  assign n2645 = n1840 & n2644;
  assign n2646 = n2496 & n2645;
  assign n2647 = ~n321 & n2646;
  assign n2648 = ~n430 & ~n527;
  assign n2649 = ~n636 & n2648;
  assign n2650 = ~n260 & n2064;
  assign n2651 = n2191 & n2650;
  assign n2652 = ~n98 & n2651;
  assign n2653 = n2649 & n2652;
  assign n2654 = ~n236 & ~n633;
  assign n2655 = ~n122 & n2654;
  assign n2656 = ~n246 & n2655;
  assign n2657 = n2653 & n2656;
  assign n2658 = ~n382 & n2657;
  assign n2659 = n2647 & n2658;
  assign n2660 = ~n315 & ~n354;
  assign n2661 = ~n535 & n2660;
  assign n2662 = ~n698 & n2661;
  assign n2663 = ~n324 & n2662;
  assign n2664 = ~n208 & n2663;
  assign n2665 = ~n454 & n2664;
  assign n2666 = ~n441 & ~n465;
  assign n2667 = ~n593 & n2666;
  assign n2668 = n2665 & n2667;
  assign n2669 = ~n330 & n2668;
  assign n2670 = n2039 & n2148;
  assign n2671 = n1110 & n2670;
  assign n2672 = n2280 & n2671;
  assign n2673 = ~n123 & n2672;
  assign n2674 = ~n580 & n2673;
  assign n2675 = n2669 & n2674;
  assign n2676 = n2659 & n2675;
  assign n2677 = ~n2640 & ~n2676;
  assign n2678 = ~n500 & n777;
  assign n2679 = ~n668 & n2678;
  assign n2680 = ~n173 & ~n374;
  assign n2681 = n1075 & n2680;
  assign n2682 = n955 & n2681;
  assign n2683 = ~n252 & ~n689;
  assign n2684 = ~n275 & ~n394;
  assign n2685 = ~n247 & n2684;
  assign n2686 = n1813 & n2685;
  assign n2687 = ~n429 & n2686;
  assign n2688 = ~n672 & n2687;
  assign n2689 = n1032 & n1859;
  assign n2690 = ~n277 & n2689;
  assign n2691 = ~n533 & n2690;
  assign n2692 = n2688 & n2691;
  assign n2693 = ~n354 & ~n632;
  assign n2694 = ~n115 & n2693;
  assign n2695 = ~n324 & n2694;
  assign n2696 = ~n245 & n2695;
  assign n2697 = ~n393 & n2199;
  assign n2698 = ~n314 & n2697;
  assign n2699 = ~n589 & n2698;
  assign n2700 = ~n304 & ~n598;
  assign n2701 = ~n349 & n2700;
  assign n2702 = n1265 & n2701;
  assign n2703 = ~n458 & n2702;
  assign n2704 = ~n256 & n1783;
  assign n2705 = ~n309 & n2704;
  assign n2706 = n2703 & n2705;
  assign n2707 = n2321 & n2706;
  assign n2708 = n2699 & n2707;
  assign n2709 = n327 & n2708;
  assign n2710 = ~n160 & n2709;
  assign n2711 = ~n261 & n2710;
  assign n2712 = n2696 & n2711;
  assign n2713 = n2692 & n2712;
  assign n2714 = n2683 & n2713;
  assign n2715 = n2682 & n2714;
  assign n2716 = ~n595 & n2715;
  assign n2717 = ~n505 & n2716;
  assign n2718 = n2679 & n2717;
  assign n2719 = ~n690 & ~n700;
  assign n2720 = ~n315 & n2719;
  assign n2721 = ~n262 & ~n538;
  assign n2722 = n2720 & n2721;
  assign n2723 = ~n216 & n2722;
  assign n2724 = ~n399 & ~n627;
  assign n2725 = ~n231 & n2724;
  assign n2726 = n2723 & n2725;
  assign n2727 = ~n614 & n2021;
  assign n2728 = ~n116 & n2727;
  assign n2729 = ~n183 & n2728;
  assign n2730 = ~n362 & n402;
  assign n2731 = n1464 & n1784;
  assign n2732 = ~n468 & n2731;
  assign n2733 = n2730 & n2732;
  assign n2734 = n1008 & n2733;
  assign n2735 = n2729 & n2734;
  assign n2736 = n2726 & n2735;
  assign n2737 = n291 & ~n464;
  assign n2738 = n1132 & n2737;
  assign n2739 = n1551 & n2738;
  assign n2740 = n1742 & n2739;
  assign n2741 = n343 & n2740;
  assign n2742 = n2736 & n2741;
  assign n2743 = ~n117 & n2742;
  assign n2744 = ~n435 & n2743;
  assign n2745 = ~n601 & n1011;
  assign n2746 = ~n465 & n2745;
  assign n2747 = n2744 & n2746;
  assign n2748 = n2718 & n2747;
  assign n2749 = ~n2676 & ~n2748;
  assign n2750 = n1181 & n1484;
  assign n2751 = n1079 & n2750;
  assign n2752 = ~n461 & n2751;
  assign n2753 = n1271 & n2520;
  assign n2754 = ~n203 & n2753;
  assign n2755 = n2752 & n2754;
  assign n2756 = ~n628 & n801;
  assign n2757 = ~n384 & n2756;
  assign n2758 = n2505 & n2757;
  assign n2759 = ~n544 & n2758;
  assign n2760 = ~n547 & ~n672;
  assign n2761 = n2131 & n2760;
  assign n2762 = n1169 & n2761;
  assign n2763 = ~n243 & n2762;
  assign n2764 = ~n194 & n2763;
  assign n2765 = n2759 & n2764;
  assign n2766 = n2755 & n2765;
  assign n2767 = ~n581 & ~n639;
  assign n2768 = ~n112 & n2767;
  assign n2769 = ~n423 & n1402;
  assign n2770 = n2768 & n2769;
  assign n2771 = ~n220 & ~n381;
  assign n2772 = ~n231 & ~n580;
  assign n2773 = ~n545 & n2772;
  assign n2774 = ~n462 & n2773;
  assign n2775 = n1724 & n2667;
  assign n2776 = ~n289 & n2775;
  assign n2777 = n2774 & n2776;
  assign n2778 = n2771 & n2777;
  assign n2779 = n2770 & n2778;
  assign n2780 = n2766 & n2779;
  assign n2781 = ~n595 & n2780;
  assign n2782 = ~n131 & n2781;
  assign n2783 = n684 & n1366;
  assign n2784 = ~n349 & n2783;
  assign n2785 = n2021 & n2784;
  assign n2786 = n2620 & n2785;
  assign n2787 = ~n693 & n2786;
  assign n2788 = n2782 & n2787;
  assign n2789 = ~n305 & n476;
  assign n2790 = ~n353 & n2789;
  assign n2791 = ~n435 & n2790;
  assign n2792 = ~n144 & ~n704;
  assign n2793 = ~n356 & n2792;
  assign n2794 = ~n187 & n2793;
  assign n2795 = n2400 & n2794;
  assign n2796 = n199 & n396;
  assign n2797 = ~n272 & n2796;
  assign n2798 = n431 & n2797;
  assign n2799 = n1015 & n2798;
  assign n2800 = n2795 & n2799;
  assign n2801 = n2309 & n2800;
  assign n2802 = n2791 & n2801;
  assign n2803 = n2788 & n2802;
  assign n2804 = ~n2748 & ~n2803;
  assign n2805 = n807 & n897;
  assign n2806 = n1058 & n2805;
  assign n2807 = n253 & n2806;
  assign n2808 = ~n681 & n2807;
  assign n2809 = ~n246 & n1700;
  assign n2810 = ~n504 & n1162;
  assign n2811 = ~n667 & n2810;
  assign n2812 = n2809 & n2811;
  assign n2813 = ~n152 & n2812;
  assign n2814 = ~n621 & ~n679;
  assign n2815 = ~n697 & n2814;
  assign n2816 = ~n315 & n2815;
  assign n2817 = ~n213 & n2816;
  assign n2818 = n2813 & n2817;
  assign n2819 = n1757 & n2818;
  assign n2820 = ~n414 & n2819;
  assign n2821 = n2808 & n2820;
  assign n2822 = ~n685 & n2066;
  assign n2823 = n291 & ~n462;
  assign n2824 = ~n692 & n2823;
  assign n2825 = n2822 & n2824;
  assign n2826 = n1618 & n2825;
  assign n2827 = ~n321 & n2826;
  assign n2828 = n282 & ~n394;
  assign n2829 = ~n307 & n2828;
  assign n2830 = n777 & n2829;
  assign n2831 = ~n360 & n2830;
  assign n2832 = n2827 & n2831;
  assign n2833 = n2821 & n2832;
  assign n2834 = ~n475 & n1285;
  assign n2835 = ~n165 & n2834;
  assign n2836 = ~n288 & ~n517;
  assign n2837 = ~n588 & n2836;
  assign n2838 = n1116 & n2837;
  assign n2839 = ~n183 & n2838;
  assign n2840 = n2835 & n2839;
  assign n2841 = ~n349 & n2840;
  assign n2842 = ~n98 & ~n336;
  assign n2843 = ~n628 & n1934;
  assign n2844 = n2081 & n2843;
  assign n2845 = n2842 & n2844;
  assign n2846 = n2841 & n2845;
  assign n2847 = n2833 & n2846;
  assign n2848 = ~n229 & n2847;
  assign n2849 = ~n106 & n2848;
  assign n2850 = ~n255 & ~n278;
  assign n2851 = ~n299 & ~n590;
  assign n2852 = n2850 & n2851;
  assign n2853 = ~n599 & n2852;
  assign n2854 = ~n85 & ~n518;
  assign n2855 = ~n598 & n2854;
  assign n2856 = n2853 & n2855;
  assign n2857 = n1204 & n2856;
  assign n2858 = n1964 & n2857;
  assign n2859 = ~n122 & n2858;
  assign n2860 = n1830 & n2648;
  assign n2861 = ~n627 & n1923;
  assign n2862 = ~n332 & n2861;
  assign n2863 = n1181 & n2862;
  assign n2864 = n2860 & n2863;
  assign n2865 = n2403 & n2864;
  assign n2866 = ~n330 & n2865;
  assign n2867 = n2859 & n2866;
  assign n2868 = ~n305 & n2867;
  assign n2869 = n1139 & n1394;
  assign n2870 = n2868 & n2869;
  assign n2871 = ~n576 & n2870;
  assign n2872 = ~n247 & n2871;
  assign n2873 = ~n350 & n2872;
  assign n2874 = n2849 & n2873;
  assign n2875 = n295 & n2090;
  assign n2876 = n706 & n2875;
  assign n2877 = ~n326 & n2876;
  assign n2878 = ~n78 & n2877;
  assign n2879 = ~n147 & ~n214;
  assign n2880 = ~n342 & n2879;
  assign n2881 = ~n535 & ~n639;
  assign n2882 = ~n242 & n2881;
  assign n2883 = n2880 & n2882;
  assign n2884 = n199 & n2883;
  assign n2885 = n1505 & n2884;
  assign n2886 = n1388 & n2885;
  assign n2887 = ~n304 & n2886;
  assign n2888 = ~n461 & n2887;
  assign n2889 = ~n361 & n2888;
  assign n2890 = n2878 & n2889;
  assign n2891 = n2874 & n2890;
  assign n2892 = ~n2803 & ~n2891;
  assign n2893 = n1711 & n2211;
  assign n2894 = n2064 & n2893;
  assign n2895 = n857 & n1659;
  assign n2896 = n233 & n2895;
  assign n2897 = n1561 & n2896;
  assign n2898 = n2505 & n2897;
  assign n2899 = n1516 & n2898;
  assign n2900 = ~n422 & n2899;
  assign n2901 = n2894 & n2900;
  assign n2902 = n1368 & n2127;
  assign n2903 = ~n477 & n2902;
  assign n2904 = ~n277 & ~n627;
  assign n2905 = n1923 & n2904;
  assign n2906 = ~n206 & n2905;
  assign n2907 = ~n594 & n2906;
  assign n2908 = n2903 & n2907;
  assign n2909 = ~n611 & n2665;
  assign n2910 = ~n350 & n2909;
  assign n2911 = n282 & n2231;
  assign n2912 = ~n88 & n2911;
  assign n2913 = ~n537 & n2912;
  assign n2914 = n2910 & n2913;
  assign n2915 = n2908 & n2914;
  assign n2916 = n1057 & n2656;
  assign n2917 = ~n134 & n2916;
  assign n2918 = n2915 & n2917;
  assign n2919 = n1268 & n2918;
  assign n2920 = ~n309 & ~n501;
  assign n2921 = ~n183 & n2920;
  assign n2922 = n167 & ~n331;
  assign n2923 = n706 & n2922;
  assign n2924 = n2921 & n2923;
  assign n2925 = ~n700 & n2924;
  assign n2926 = n2919 & n2925;
  assign n2927 = n2901 & n2926;
  assign n2928 = ~n2891 & ~n2927;
  assign n2929 = ~n414 & ~n504;
  assign n2930 = ~n206 & n2929;
  assign n2931 = ~n679 & n2930;
  assign n2932 = n1238 & n2931;
  assign n2933 = n1390 & n2932;
  assign n2934 = n1482 & n2933;
  assign n2935 = n1283 & n1646;
  assign n2936 = ~n589 & n2935;
  assign n2937 = ~n242 & n2936;
  assign n2938 = ~n505 & n1259;
  assign n2939 = ~n161 & n2938;
  assign n2940 = ~n180 & ~n297;
  assign n2941 = ~n272 & n511;
  assign n2942 = ~n600 & n2941;
  assign n2943 = ~n279 & n1247;
  assign n2944 = ~n170 & ~n373;
  assign n2945 = n2943 & n2944;
  assign n2946 = n2694 & n2945;
  assign n2947 = n2942 & n2946;
  assign n2948 = n2940 & n2947;
  assign n2949 = n2939 & n2948;
  assign n2950 = n901 & n2949;
  assign n2951 = ~n307 & n2950;
  assign n2952 = ~n633 & n2951;
  assign n2953 = n2937 & n2952;
  assign n2954 = ~n362 & n1182;
  assign n2955 = ~n705 & n2954;
  assign n2956 = ~n548 & n2955;
  assign n2957 = ~n332 & n1993;
  assign n2958 = ~n594 & n1539;
  assign n2959 = ~n535 & n2958;
  assign n2960 = n2957 & n2959;
  assign n2961 = n2842 & n2960;
  assign n2962 = n2956 & n2961;
  assign n2963 = n2772 & n2962;
  assign n2964 = ~n700 & n2963;
  assign n2965 = ~n360 & n2964;
  assign n2966 = n306 & n2548;
  assign n2967 = ~n353 & n2966;
  assign n2968 = ~n323 & n2967;
  assign n2969 = n2965 & n2968;
  assign n2970 = n2953 & n2969;
  assign n2971 = n480 & n2970;
  assign n2972 = ~n704 & n2971;
  assign n2973 = n2934 & n2972;
  assign n2974 = ~n681 & n865;
  assign n2975 = ~n195 & ~n428;
  assign n2976 = ~n538 & n2975;
  assign n2977 = n2974 & n2976;
  assign n2978 = ~n308 & n2977;
  assign n2979 = ~n356 & ~n544;
  assign n2980 = ~n701 & n2979;
  assign n2981 = ~n132 & n2980;
  assign n2982 = n2978 & n2981;
  assign n2983 = ~n670 & n2585;
  assign n2984 = ~n293 & n615;
  assign n2985 = ~n341 & n2984;
  assign n2986 = n2983 & n2985;
  assign n2987 = n2982 & n2986;
  assign n2988 = ~n692 & n2987;
  assign n2989 = n2281 & n2904;
  assign n2990 = ~n372 & n2989;
  assign n2991 = ~n149 & ~n579;
  assign n2992 = n1232 & n2991;
  assign n2993 = ~n698 & n2992;
  assign n2994 = ~n621 & n2993;
  assign n2995 = n2990 & n2994;
  assign n2996 = ~n374 & n2995;
  assign n2997 = ~n152 & ~n289;
  assign n2998 = ~n171 & n282;
  assign n2999 = n2997 & n2998;
  assign n3000 = n2996 & n2999;
  assign n3001 = n453 & n2094;
  assign n3002 = n3000 & n3001;
  assign n3003 = ~n683 & n3002;
  assign n3004 = n2988 & n3003;
  assign n3005 = n2973 & n3004;
  assign n3006 = ~n2927 & ~n3005;
  assign n3007 = ~n132 & ~n325;
  assign n3008 = ~n385 & n3007;
  assign n3009 = n884 & n3008;
  assign n3010 = n1625 & n3009;
  assign n3011 = ~n122 & n3010;
  assign n3012 = n1058 & n2342;
  assign n3013 = n1116 & n3012;
  assign n3014 = n1232 & n3013;
  assign n3015 = ~n85 & n3014;
  assign n3016 = n3011 & n3015;
  assign n3017 = n333 & ~n588;
  assign n3018 = ~n353 & n392;
  assign n3019 = ~n612 & n3018;
  assign n3020 = n3017 & n3019;
  assign n3021 = n2921 & n3020;
  assign n3022 = ~n208 & n3021;
  assign n3023 = n1936 & n2280;
  assign n3024 = ~n578 & n3023;
  assign n3025 = n1823 & n3024;
  assign n3026 = ~n172 & n3025;
  assign n3027 = ~n394 & n3026;
  assign n3028 = n3022 & n3027;
  assign n3029 = n3016 & n3028;
  assign n3030 = ~n88 & ~n112;
  assign n3031 = n196 & n3030;
  assign n3032 = ~n160 & n3031;
  assign n3033 = ~n580 & n1348;
  assign n3034 = ~n330 & n3033;
  assign n3035 = ~n129 & n3034;
  assign n3036 = n3032 & n3035;
  assign n3037 = n966 & n3036;
  assign n3038 = ~n134 & n515;
  assign n3039 = ~n502 & n3038;
  assign n3040 = ~n188 & n3039;
  assign n3041 = n2373 & n3040;
  assign n3042 = n3037 & n3041;
  assign n3043 = n3029 & n3042;
  assign n3044 = n797 & n3043;
  assign n3045 = ~n461 & ~n666;
  assign n3046 = n838 & n3045;
  assign n3047 = n1397 & n3046;
  assign n3048 = n1724 & n3047;
  assign n3049 = ~n682 & n1784;
  assign n3050 = ~n154 & ~n517;
  assign n3051 = ~n399 & n3050;
  assign n3052 = n1588 & n3051;
  assign n3053 = n865 & n3052;
  assign n3054 = ~n320 & n3053;
  assign n3055 = ~n213 & ~n414;
  assign n3056 = ~n278 & n3055;
  assign n3057 = ~n206 & n1111;
  assign n3058 = ~n398 & ~n632;
  assign n3059 = ~n314 & n3058;
  assign n3060 = ~n671 & n3059;
  assign n3061 = n3057 & n3060;
  assign n3062 = n1347 & n3061;
  assign n3063 = n3056 & n3062;
  assign n3064 = ~n117 & ~n705;
  assign n3065 = ~n372 & n3064;
  assign n3066 = ~n544 & ~n601;
  assign n3067 = n3065 & n3066;
  assign n3068 = ~n613 & n3067;
  assign n3069 = ~n323 & ~n475;
  assign n3070 = ~n242 & n3069;
  assign n3071 = n3068 & n3070;
  assign n3072 = n3063 & n3071;
  assign n3073 = ~n381 & n3072;
  assign n3074 = n3054 & n3073;
  assign n3075 = ~n361 & n3074;
  assign n3076 = n3049 & n3075;
  assign n3077 = n2494 & n3076;
  assign n3078 = n3048 & n3077;
  assign n3079 = ~n356 & ~n533;
  assign n3080 = ~n220 & n3079;
  assign n3081 = ~n173 & n930;
  assign n3082 = ~n468 & ~n701;
  assign n3083 = n3081 & n3082;
  assign n3084 = ~n78 & ~n114;
  assign n3085 = ~n537 & n3084;
  assign n3086 = n3083 & n3085;
  assign n3087 = n3080 & n3086;
  assign n3088 = n3078 & n3087;
  assign n3089 = ~n217 & n3088;
  assign n3090 = n3044 & n3089;
  assign n3091 = ~n123 & n3090;
  assign n3092 = ~n458 & n2066;
  assign n3093 = ~n473 & n3092;
  assign n3094 = n3091 & n3093;
  assign n3095 = ~n669 & n3094;
  assign n3096 = ~n149 & n1814;
  assign n3097 = n3095 & n3096;
  assign n3098 = ~n3005 & ~n3097;
  assign n3099 = n1321 & n2494;
  assign n3100 = n1435 & n3099;
  assign n3101 = ~n310 & n3100;
  assign n3102 = ~n149 & n3101;
  assign n3103 = ~n160 & ~n382;
  assign n3104 = ~n385 & ~n580;
  assign n3105 = ~n423 & n3104;
  assign n3106 = ~n281 & n3105;
  assign n3107 = n3103 & n3106;
  assign n3108 = n2064 & n3107;
  assign n3109 = ~n695 & n3108;
  assign n3110 = n940 & n1936;
  assign n3111 = ~n94 & n3110;
  assign n3112 = n3109 & n3111;
  assign n3113 = ~n321 & ~n336;
  assign n3114 = ~n155 & n1057;
  assign n3115 = n3113 & n3114;
  assign n3116 = ~n637 & n3115;
  assign n3117 = ~n463 & ~n537;
  assign n3118 = ~n104 & ~n228;
  assign n3119 = ~n429 & n2123;
  assign n3120 = n3118 & n3119;
  assign n3121 = ~n112 & n3120;
  assign n3122 = ~n356 & ~n477;
  assign n3123 = ~n424 & n3122;
  assign n3124 = ~n349 & n3123;
  assign n3125 = n3121 & n3124;
  assign n3126 = n3117 & n3125;
  assign n3127 = ~n247 & n3126;
  assign n3128 = ~n81 & n3127;
  assign n3129 = n3116 & n3128;
  assign n3130 = n3112 & n3129;
  assign n3131 = ~n670 & n3130;
  assign n3132 = n1252 & n3131;
  assign n3133 = n1089 & n3132;
  assign n3134 = n415 & n3133;
  assign n3135 = n2818 & n3134;
  assign n3136 = n2879 & n3135;
  assign n3137 = n3102 & n3136;
  assign n3138 = ~n98 & ~n400;
  assign n3139 = n174 & n2766;
  assign n3140 = n3138 & n3139;
  assign n3141 = ~n700 & n3140;
  assign n3142 = ~n466 & n3141;
  assign n3143 = n2218 & n2648;
  assign n3144 = ~n373 & n3143;
  assign n3145 = ~n208 & n3144;
  assign n3146 = n768 & n1911;
  assign n3147 = ~n235 & n3146;
  assign n3148 = ~n381 & n3147;
  assign n3149 = n3145 & n3148;
  assign n3150 = n437 & ~n593;
  assign n3151 = ~n325 & n3150;
  assign n3152 = ~n626 & n3151;
  assign n3153 = ~n353 & n1383;
  assign n3154 = ~n277 & n3153;
  assign n3155 = ~n181 & n3154;
  assign n3156 = n3152 & n3155;
  assign n3157 = n3149 & n3156;
  assign n3158 = ~n260 & ~n632;
  assign n3159 = ~n533 & n3158;
  assign n3160 = ~n506 & n3159;
  assign n3161 = ~n398 & n3160;
  assign n3162 = n3157 & n3161;
  assign n3163 = ~n254 & n3162;
  assign n3164 = ~n304 & n3163;
  assign n3165 = n3142 & n3164;
  assign n3166 = n3137 & n3165;
  assign n3167 = ~n3097 & ~n3166;
  assign n3168 = ~n115 & ~n204;
  assign n3169 = ~n309 & n3168;
  assign n3170 = ~n172 & n3169;
  assign n3171 = n910 & n3170;
  assign n3172 = n1784 & n3171;
  assign n3173 = ~n401 & n3172;
  assign n3174 = n1390 & n1577;
  assign n3175 = ~n610 & n3174;
  assign n3176 = ~n627 & n3175;
  assign n3177 = n3173 & n3176;
  assign n3178 = n1791 & n2032;
  assign n3179 = ~n374 & n3178;
  assign n3180 = ~n315 & n2683;
  assign n3181 = ~n261 & n3180;
  assign n3182 = n3179 & n3181;
  assign n3183 = n3177 & n3182;
  assign n3184 = n819 & n3183;
  assign n3185 = ~n373 & n3184;
  assign n3186 = ~n465 & n3185;
  assign n3187 = ~n345 & ~n400;
  assign n3188 = n546 & n3187;
  assign n3189 = ~n106 & n3188;
  assign n3190 = ~n353 & n655;
  assign n3191 = ~n183 & n3190;
  assign n3192 = n3189 & n3191;
  assign n3193 = n1246 & n1281;
  assign n3194 = ~n324 & n3193;
  assign n3195 = ~n384 & ~n436;
  assign n3196 = n1797 & n3195;
  assign n3197 = n196 & n3196;
  assign n3198 = ~n441 & n3197;
  assign n3199 = ~n360 & n3198;
  assign n3200 = n3194 & n3199;
  assign n3201 = n3192 & n3200;
  assign n3202 = ~n88 & ~n161;
  assign n3203 = n1373 & n3202;
  assign n3204 = n3130 & n3203;
  assign n3205 = n3201 & n3204;
  assign n3206 = ~n341 & n3205;
  assign n3207 = ~n533 & n3206;
  assign n3208 = n3186 & n3207;
  assign n3209 = ~n697 & n907;
  assign n3210 = ~n700 & n3209;
  assign n3211 = ~n669 & n3210;
  assign n3212 = n476 & n3211;
  assign n3213 = ~n180 & n3212;
  assign n3214 = ~n547 & n3213;
  assign n3215 = ~n502 & ~n517;
  assign n3216 = n240 & ~n331;
  assign n3217 = ~n232 & ~n330;
  assign n3218 = ~n422 & n3217;
  assign n3219 = ~n398 & n3218;
  assign n3220 = n3216 & n3219;
  assign n3221 = n3215 & n3220;
  assign n3222 = ~n334 & n3221;
  assign n3223 = ~n391 & n3222;
  assign n3224 = ~n600 & n3223;
  assign n3225 = n3214 & n3224;
  assign n3226 = n3208 & n3225;
  assign n3227 = ~n3166 & ~n3226;
  assign n3228 = ~n114 & ~n256;
  assign n3229 = ~n129 & n3228;
  assign n3230 = ~n307 & n3229;
  assign n3231 = ~n195 & ~n464;
  assign n3232 = n3230 & n3231;
  assign n3233 = ~n399 & n3232;
  assign n3234 = ~n247 & n680;
  assign n3235 = ~n442 & n3234;
  assign n3236 = n3233 & n3235;
  assign n3237 = n2231 & n3236;
  assign n3238 = ~n279 & n3237;
  assign n3239 = ~n122 & n167;
  assign n3240 = ~n150 & n3239;
  assign n3241 = ~n187 & n3240;
  assign n3242 = ~n330 & ~n636;
  assign n3243 = ~n669 & n3242;
  assign n3244 = ~n692 & n3114;
  assign n3245 = ~n203 & n3244;
  assign n3246 = n3243 & n3245;
  assign n3247 = ~n149 & ~n505;
  assign n3248 = ~n81 & n3247;
  assign n3249 = n3246 & n3248;
  assign n3250 = n3241 & n3249;
  assign n3251 = ~n297 & n3250;
  assign n3252 = ~n461 & n3251;
  assign n3253 = n3238 & n3252;
  assign n3254 = n1581 & n2648;
  assign n3255 = n853 & n3254;
  assign n3256 = n1651 & n3255;
  assign n3257 = n306 & n3256;
  assign n3258 = ~n538 & n3257;
  assign n3259 = n1859 & n2027;
  assign n3260 = ~n299 & n3259;
  assign n3261 = ~n639 & n3260;
  assign n3262 = n3258 & n3261;
  assign n3263 = n3253 & n3262;
  assign n3264 = ~n3226 & ~n3263;
  assign n3265 = ~n683 & n2481;
  assign n3266 = n907 & n1148;
  assign n3267 = ~n342 & n3266;
  assign n3268 = n3265 & n3267;
  assign n3269 = ~n669 & n3268;
  assign n3270 = ~n132 & ~n545;
  assign n3271 = ~n462 & n3270;
  assign n3272 = ~n324 & n3271;
  assign n3273 = ~n582 & ~n629;
  assign n3274 = ~n594 & n3273;
  assign n3275 = ~n614 & n3274;
  assign n3276 = ~n384 & n3275;
  assign n3277 = n3272 & n3276;
  assign n3278 = n2392 & n2474;
  assign n3279 = n1767 & n3278;
  assign n3280 = ~n693 & n3279;
  assign n3281 = ~n236 & ~n399;
  assign n3282 = ~n375 & n3281;
  assign n3283 = ~n468 & n3282;
  assign n3284 = ~n232 & n3283;
  assign n3285 = n1622 & n3284;
  assign n3286 = n758 & n3285;
  assign n3287 = ~n131 & n3286;
  assign n3288 = ~n639 & n3287;
  assign n3289 = n3280 & n3288;
  assign n3290 = ~n106 & n3289;
  assign n3291 = n2588 & n3215;
  assign n3292 = ~n186 & n3291;
  assign n3293 = n2273 & n3292;
  assign n3294 = n3290 & n3293;
  assign n3295 = n3277 & n3294;
  assign n3296 = n558 & n3295;
  assign n3297 = ~n393 & n3296;
  assign n3298 = ~n187 & n3297;
  assign n3299 = n3269 & n3298;
  assign n3300 = ~n183 & ~n325;
  assign n3301 = ~n280 & n3300;
  assign n3302 = n1089 & n3301;
  assign n3303 = n148 & n3302;
  assign n3304 = ~n290 & n3303;
  assign n3305 = ~n304 & ~n469;
  assign n3306 = ~n198 & n1285;
  assign n3307 = n1732 & n3306;
  assign n3308 = ~n536 & n3307;
  assign n3309 = ~n194 & ~n636;
  assign n3310 = ~n134 & n3309;
  assign n3311 = ~n381 & n3310;
  assign n3312 = n3308 & n3311;
  assign n3313 = n3305 & n3312;
  assign n3314 = ~n628 & n3313;
  assign n3315 = ~n435 & n3314;
  assign n3316 = n3304 & n3315;
  assign n3317 = n1813 & n3030;
  assign n3318 = ~n442 & n3317;
  assign n3319 = ~n160 & ~n535;
  assign n3320 = ~n429 & n3319;
  assign n3321 = ~n309 & n3320;
  assign n3322 = ~n245 & n3321;
  assign n3323 = n3318 & n3322;
  assign n3324 = ~n350 & n3323;
  assign n3325 = ~n464 & n2056;
  assign n3326 = n920 & n3325;
  assign n3327 = ~n599 & n838;
  assign n3328 = ~n254 & n3327;
  assign n3329 = n3326 & n3328;
  assign n3330 = n3324 & n3329;
  assign n3331 = n1539 & n3330;
  assign n3332 = n221 & n3331;
  assign n3333 = ~n277 & n3332;
  assign n3334 = n2418 & n2630;
  assign n3335 = ~n581 & n3334;
  assign n3336 = ~n413 & n3335;
  assign n3337 = n3333 & n3336;
  assign n3338 = n3316 & n3337;
  assign n3339 = ~n173 & ~n590;
  assign n3340 = ~n171 & n3339;
  assign n3341 = ~n320 & n3340;
  assign n3342 = n3338 & n3341;
  assign n3343 = n476 & n3342;
  assign n3344 = ~n390 & n3343;
  assign n3345 = ~n671 & n3344;
  assign n3346 = ~n593 & n1544;
  assign n3347 = ~n247 & n3346;
  assign n3348 = ~n81 & n3045;
  assign n3349 = n3347 & n3348;
  assign n3350 = ~n206 & n3349;
  assign n3351 = ~n595 & ~n611;
  assign n3352 = ~n428 & n3351;
  assign n3353 = ~n260 & n3352;
  assign n3354 = n3350 & n3353;
  assign n3355 = n459 & n3354;
  assign n3356 = ~n166 & n3355;
  assign n3357 = ~n78 & n3356;
  assign n3358 = ~n638 & n3357;
  assign n3359 = n3345 & n3358;
  assign n3360 = n3299 & n3359;
  assign n3361 = ~n3263 & ~n3360;
  assign n3362 = n3263 & n3360;
  assign n3363 = ~n3361 & ~n3362;
  assign n3364 = ~n428 & n2060;
  assign n3365 = n1063 & n1588;
  assign n3366 = ~n501 & n1132;
  assign n3367 = ~n535 & n3366;
  assign n3368 = n777 & n3367;
  assign n3369 = n3365 & n3368;
  assign n3370 = ~n462 & n3369;
  assign n3371 = ~n104 & ~n187;
  assign n3372 = ~n239 & ~n578;
  assign n3373 = n346 & n3372;
  assign n3374 = ~n197 & n3373;
  assign n3375 = n3371 & n3374;
  assign n3376 = ~n362 & n744;
  assign n3377 = ~n424 & n1442;
  assign n3378 = ~n598 & n3377;
  assign n3379 = n3376 & n3378;
  assign n3380 = n2772 & n3379;
  assign n3381 = n3375 & n3380;
  assign n3382 = ~n117 & n1272;
  assign n3383 = ~n165 & n3382;
  assign n3384 = n3381 & n3383;
  assign n3385 = n3370 & n3384;
  assign n3386 = n3364 & n3385;
  assign n3387 = n282 & ~n475;
  assign n3388 = ~n393 & n3387;
  assign n3389 = n3386 & n3388;
  assign n3390 = n955 & n3389;
  assign n3391 = ~n154 & n3390;
  assign n3392 = ~n216 & ~n458;
  assign n3393 = n2588 & n3392;
  assign n3394 = n2529 & n3393;
  assign n3395 = n2929 & n3394;
  assign n3396 = ~n251 & n3395;
  assign n3397 = n3391 & n3396;
  assign n3398 = ~n332 & n3397;
  assign n3399 = ~n666 & n1148;
  assign n3400 = ~n252 & n3399;
  assign n3401 = ~n547 & n1923;
  assign n3402 = ~n336 & n3401;
  assign n3403 = ~n678 & n3402;
  assign n3404 = ~n123 & n300;
  assign n3405 = ~n315 & n788;
  assign n3406 = ~n399 & n3405;
  assign n3407 = n3404 & n3406;
  assign n3408 = ~n704 & n1641;
  assign n3409 = ~n220 & n3408;
  assign n3410 = n3407 & n3409;
  assign n3411 = n3403 & n3410;
  assign n3412 = ~n614 & ~n679;
  assign n3413 = ~n277 & n3412;
  assign n3414 = n2114 & n3413;
  assign n3415 = n3411 & n3414;
  assign n3416 = ~n536 & n3415;
  assign n3417 = n3400 & n3416;
  assign n3418 = n3161 & n3242;
  assign n3419 = n89 & n3418;
  assign n3420 = n1478 & n3419;
  assign n3421 = ~n422 & n3420;
  assign n3422 = ~n363 & n787;
  assign n3423 = n244 & n3422;
  assign n3424 = n1451 & n3423;
  assign n3425 = n2070 & n3424;
  assign n3426 = ~n275 & n3425;
  assign n3427 = ~n582 & n3426;
  assign n3428 = n3421 & n3427;
  assign n3429 = n3417 & n3428;
  assign n3430 = ~n627 & n2418;
  assign n3431 = ~n454 & n3430;
  assign n3432 = ~n247 & n2199;
  assign n3433 = ~n144 & n3432;
  assign n3434 = n3431 & n3433;
  assign n3435 = ~n106 & n3434;
  assign n3436 = ~n183 & n1565;
  assign n3437 = ~n356 & n3436;
  assign n3438 = n1823 & n3437;
  assign n3439 = n3435 & n3438;
  assign n3440 = n3429 & n3439;
  assign n3441 = n562 & n3440;
  assign n3442 = ~n473 & ~n611;
  assign n3443 = ~n349 & ~n465;
  assign n3444 = n3442 & n3443;
  assign n3445 = n1720 & n3444;
  assign n3446 = n445 & n3445;
  assign n3447 = n3441 & n3446;
  assign n3448 = ~n695 & n3447;
  assign n3449 = n322 & n3448;
  assign n3450 = n3398 & n3449;
  assign n3451 = n3360 & n3450;
  assign n3452 = ~n363 & n2373;
  assign n3453 = ~n170 & n3452;
  assign n3454 = ~n134 & ~n391;
  assign n3455 = ~n207 & n3454;
  assign n3456 = ~n668 & n3455;
  assign n3457 = n3453 & n3456;
  assign n3458 = ~n208 & n3202;
  assign n3459 = ~n277 & n3458;
  assign n3460 = ~n220 & ~n414;
  assign n3461 = ~n197 & n3460;
  assign n3462 = ~n473 & n3461;
  assign n3463 = n3459 & n3462;
  assign n3464 = n3457 & n3463;
  assign n3465 = n725 & n3464;
  assign n3466 = n2021 & n3465;
  assign n3467 = ~n203 & n3466;
  assign n3468 = ~n262 & ~n429;
  assign n3469 = ~n704 & n3468;
  assign n3470 = ~n469 & n3469;
  assign n3471 = ~n150 & ~n272;
  assign n3472 = n2566 & n3471;
  assign n3473 = ~n100 & n3472;
  assign n3474 = n3470 & n3473;
  assign n3475 = ~n228 & n3474;
  assign n3476 = n3467 & n3475;
  assign n3477 = n295 & n768;
  assign n3478 = ~n122 & ~n672;
  assign n3479 = ~n599 & n3478;
  assign n3480 = n2234 & n3479;
  assign n3481 = n896 & n3480;
  assign n3482 = n3477 & n3481;
  assign n3483 = n3071 & n3482;
  assign n3484 = ~n360 & n3483;
  assign n3485 = ~n172 & n456;
  assign n3486 = ~n252 & n1954;
  assign n3487 = ~n160 & n3486;
  assign n3488 = n3485 & n3487;
  assign n3489 = n684 & n3488;
  assign n3490 = ~n280 & n3489;
  assign n3491 = ~n457 & n3490;
  assign n3492 = n3484 & n3491;
  assign n3493 = ~n464 & n3492;
  assign n3494 = n148 & ~n394;
  assign n3495 = n3493 & n3494;
  assign n3496 = n317 & n3495;
  assign n3497 = ~n235 & n3496;
  assign n3498 = ~n180 & ~n439;
  assign n3499 = ~n692 & n3498;
  assign n3500 = n1247 & n3499;
  assign n3501 = n3024 & n3500;
  assign n3502 = n3294 & n3501;
  assign n3503 = n797 & n3502;
  assign n3504 = ~n261 & n3503;
  assign n3505 = n3497 & n3504;
  assign n3506 = n3476 & n3505;
  assign n3507 = ~n3451 & ~n3506;
  assign n3508 = n3363 & n3507;
  assign n3509 = ~n3361 & ~n3508;
  assign n3510 = n3226 & n3263;
  assign n3511 = ~n3264 & ~n3510;
  assign n3512 = ~n3509 & n3511;
  assign n3513 = ~n3264 & ~n3512;
  assign n3514 = n3166 & n3226;
  assign n3515 = ~n3227 & ~n3514;
  assign n3516 = ~n3513 & n3515;
  assign n3517 = ~n3227 & ~n3516;
  assign n3518 = n3097 & n3166;
  assign n3519 = ~n3167 & ~n3518;
  assign n3520 = ~n3517 & n3519;
  assign n3521 = ~n3167 & ~n3520;
  assign n3522 = n3005 & n3097;
  assign n3523 = ~n3098 & ~n3522;
  assign n3524 = ~n3521 & n3523;
  assign n3525 = ~n3098 & ~n3524;
  assign n3526 = n2927 & n3005;
  assign n3527 = ~n3006 & ~n3526;
  assign n3528 = ~n3525 & n3527;
  assign n3529 = ~n3006 & ~n3528;
  assign n3530 = n2891 & n2927;
  assign n3531 = ~n2928 & ~n3530;
  assign n3532 = ~n3529 & n3531;
  assign n3533 = ~n2928 & ~n3532;
  assign n3534 = n2803 & n2891;
  assign n3535 = ~n2892 & ~n3534;
  assign n3536 = ~n3533 & n3535;
  assign n3537 = ~n2892 & ~n3536;
  assign n3538 = n2748 & n2803;
  assign n3539 = ~n2804 & ~n3538;
  assign n3540 = ~n3537 & n3539;
  assign n3541 = ~n2804 & ~n3540;
  assign n3542 = n2676 & n2748;
  assign n3543 = ~n2749 & ~n3542;
  assign n3544 = ~n3541 & n3543;
  assign n3545 = ~n2749 & ~n3544;
  assign n3546 = n2640 & n2676;
  assign n3547 = ~n2677 & ~n3546;
  assign n3548 = ~n3545 & n3547;
  assign n3549 = ~n2677 & ~n3548;
  assign n3550 = n2554 & n2640;
  assign n3551 = ~n2641 & ~n3550;
  assign n3552 = ~n3549 & n3551;
  assign n3553 = ~n2641 & ~n3552;
  assign n3554 = n2457 & n2554;
  assign n3555 = ~n2555 & ~n3554;
  assign n3556 = ~n3553 & n3555;
  assign n3557 = ~n2555 & ~n3556;
  assign n3558 = n2369 & n2457;
  assign n3559 = ~n2458 & ~n3558;
  assign n3560 = ~n3557 & n3559;
  assign n3561 = ~n2458 & ~n3560;
  assign n3562 = n2278 & n2369;
  assign n3563 = ~n2370 & ~n3562;
  assign n3564 = ~n3561 & n3563;
  assign n3565 = ~n2370 & ~n3564;
  assign n3566 = n2178 & n2278;
  assign n3567 = ~n2279 & ~n3566;
  assign n3568 = ~n3565 & n3567;
  assign n3569 = ~n2279 & ~n3568;
  assign n3570 = n2058 & n2178;
  assign n3571 = ~n2179 & ~n3570;
  assign n3572 = ~n3569 & n3571;
  assign n3573 = ~n2179 & ~n3572;
  assign n3574 = n2006 & n2058;
  assign n3575 = ~n2059 & ~n3574;
  assign n3576 = ~n3573 & n3575;
  assign n3577 = ~n2059 & ~n3576;
  assign n3578 = n1900 & n2006;
  assign n3579 = ~n2007 & ~n3578;
  assign n3580 = ~n3577 & n3579;
  assign n3581 = ~n2007 & ~n3580;
  assign n3582 = n1811 & n1900;
  assign n3583 = ~n1901 & ~n3582;
  assign n3584 = ~n3581 & n3583;
  assign n3585 = ~n1901 & ~n3584;
  assign n3586 = n1740 & n1811;
  assign n3587 = ~n1812 & ~n3586;
  assign n3588 = ~n3585 & n3587;
  assign n3589 = ~n1812 & ~n3588;
  assign n3590 = n1610 & n1740;
  assign n3591 = ~n1741 & ~n3590;
  assign n3592 = ~n3589 & n3591;
  assign n3593 = ~n1741 & ~n3592;
  assign n3594 = n1531 & n1610;
  assign n3595 = ~n1611 & ~n3594;
  assign n3596 = ~n3593 & n3595;
  assign n3597 = ~n1611 & ~n3596;
  assign n3598 = n1426 & n1531;
  assign n3599 = ~n1532 & ~n3598;
  assign n3600 = ~n3597 & n3599;
  assign n3601 = ~n1532 & ~n3600;
  assign n3602 = n1338 & n1426;
  assign n3603 = ~n1427 & ~n3602;
  assign n3604 = ~n3601 & n3603;
  assign n3605 = ~n1427 & ~n3604;
  assign n3606 = n1230 & n1338;
  assign n3607 = ~n1339 & ~n3606;
  assign n3608 = ~n3605 & n3607;
  assign n3609 = ~n1339 & ~n3608;
  assign n3610 = n1107 & n1230;
  assign n3611 = ~n1231 & ~n3610;
  assign n3612 = ~n3609 & n3611;
  assign n3613 = ~n1231 & ~n3612;
  assign n3614 = n1005 & n1107;
  assign n3615 = ~n1108 & ~n3614;
  assign n3616 = ~n3613 & n3615;
  assign n3617 = ~n1108 & ~n3616;
  assign n3618 = n894 & n1005;
  assign n3619 = ~n1006 & ~n3618;
  assign n3620 = ~n3617 & n3619;
  assign n3621 = ~n1006 & ~n3620;
  assign n3622 = n795 & n894;
  assign n3623 = ~n895 & ~n3622;
  assign n3624 = ~n3621 & n3623;
  assign n3625 = ~n895 & ~n3624;
  assign n3626 = n665 & n795;
  assign n3627 = ~n796 & ~n3626;
  assign n3628 = ~n3625 & n3627;
  assign n3629 = ~n796 & ~n3628;
  assign n3630 = n665 & n720;
  assign n3631 = ~n721 & ~n3630;
  assign n3632 = ~n3629 & n3631;
  assign n3633 = ~n721 & ~n3632;
  assign n3634 = ~n554 & ~n720;
  assign n3635 = n526 & n720;
  assign n3636 = ~n3634 & ~n3635;
  assign n3637 = ~n3633 & n3636;
  assign n3638 = n720 & ~n3637;
  assign n3639 = n556 & ~n3638;
  assign n3640 = pi30  & n555;
  assign n3641 = pi31  & n3640;
  assign n3642 = ~n3639 & ~n3641;
  assign n3643 = ~n554 & ~n3642;
  assign n3644 = ~n412 & n498;
  assign n3645 = ~n499 & ~n3644;
  assign n3646 = n3643 & n3645;
  assign n3647 = ~n499 & ~n3646;
  assign n3648 = n492 & ~n666;
  assign n3649 = ~n193 & n3648;
  assign n3650 = n211 & n234;
  assign n3651 = ~n242 & n3650;
  assign n3652 = n712 & n3651;
  assign n3653 = n653 & n3652;
  assign n3654 = n3649 & n3653;
  assign n3655 = n412 & n3654;
  assign n3656 = ~n412 & ~n3654;
  assign n3657 = ~n3655 & ~n3656;
  assign n3658 = ~n3647 & ~n3657;
  assign n3659 = ~n3647 & n3657;
  assign n3660 = n3647 & ~n3657;
  assign n3661 = ~n3659 & ~n3660;
  assign n3662 = ~n3643 & ~n3645;
  assign n3663 = ~n3646 & ~n3662;
  assign n3664 = ~n334 & n788;
  assign n3665 = ~n401 & n3664;
  assign n3666 = n222 & ~n504;
  assign n3667 = ~n149 & n3666;
  assign n3668 = n3665 & n3667;
  assign n3669 = ~n147 & n3668;
  assign n3670 = ~n697 & n1222;
  assign n3671 = ~n685 & n3670;
  assign n3672 = ~n337 & n3671;
  assign n3673 = ~n204 & n3672;
  assign n3674 = ~n439 & n3673;
  assign n3675 = n3669 & n3674;
  assign n3676 = ~n430 & n3675;
  assign n3677 = ~n517 & n3676;
  assign n3678 = ~n441 & n3677;
  assign n3679 = n2027 & n3678;
  assign n3680 = n3242 & n3679;
  assign n3681 = n1904 & n3680;
  assign n3682 = n2180 & n3681;
  assign n3683 = ~n362 & n3682;
  assign n3684 = ~n239 & n3683;
  assign n3685 = n2484 & n3282;
  assign n3686 = n1246 & n3685;
  assign n3687 = ~n626 & n3686;
  assign n3688 = ~n251 & n3687;
  assign n3689 = n3684 & n3688;
  assign n3690 = n343 & ~n518;
  assign n3691 = ~n357 & n3690;
  assign n3692 = ~n455 & n3691;
  assign n3693 = ~n160 & ~n363;
  assign n3694 = ~n395 & n3693;
  assign n3695 = ~n360 & ~n502;
  assign n3696 = ~n345 & n3695;
  assign n3697 = ~n465 & n3696;
  assign n3698 = n3694 & n3697;
  assign n3699 = ~n100 & ~n631;
  assign n3700 = ~n324 & n3699;
  assign n3701 = n3698 & n3700;
  assign n3702 = n3692 & n3701;
  assign n3703 = ~n104 & n248;
  assign n3704 = ~n173 & n3703;
  assign n3705 = n1679 & n3704;
  assign n3706 = n2066 & n3705;
  assign n3707 = n3702 & n3706;
  assign n3708 = ~n612 & n3707;
  assign n3709 = n230 & ~n695;
  assign n3710 = ~n183 & n3709;
  assign n3711 = ~n323 & n3710;
  assign n3712 = n3708 & n3711;
  assign n3713 = n3689 & n3712;
  assign n3714 = ~n152 & n1791;
  assign n3715 = ~n442 & ~n538;
  assign n3716 = n785 & n3715;
  assign n3717 = n3714 & n3716;
  assign n3718 = n2088 & n3717;
  assign n3719 = n2195 & n3718;
  assign n3720 = n2467 & n3719;
  assign n3721 = n319 & n607;
  assign n3722 = n3720 & n3721;
  assign n3723 = n494 & n3722;
  assign n3724 = ~n242 & ~n465;
  assign n3725 = n140 & n519;
  assign n3726 = ~n183 & n3725;
  assign n3727 = n3724 & n3726;
  assign n3728 = n3723 & n3727;
  assign n3729 = ~n3713 & ~n3728;
  assign n3730 = n3713 & n3728;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = ~pi29  & n3731;
  assign n3733 = ~n3729 & ~n3732;
  assign n3734 = n412 & ~n3733;
  assign n3735 = ~n412 & n3733;
  assign n3736 = ~n720 & n3641;
  assign n3737 = pi30  & ~pi31 ;
  assign n3738 = ~pi30  & pi31 ;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = n555 & ~n3739;
  assign n3741 = ~n554 & n3740;
  assign n3742 = ~n554 & n3638;
  assign n3743 = n554 & n3637;
  assign n3744 = ~n3742 & ~n3743;
  assign n3745 = n556 & ~n3744;
  assign n3746 = ~n3741 & ~n3745;
  assign n3747 = ~n3736 & n3746;
  assign n3748 = ~n3735 & ~n3747;
  assign n3749 = ~n3734 & ~n3748;
  assign n3750 = n3663 & ~n3749;
  assign n3751 = ~n3663 & n3749;
  assign n3752 = ~n3750 & ~n3751;
  assign n3753 = ~n116 & ~n527;
  assign n3754 = ~n462 & n3753;
  assign n3755 = n135 & ~n279;
  assign n3756 = ~n505 & n3755;
  assign n3757 = n3754 & n3756;
  assign n3758 = n630 & n1252;
  assign n3759 = n386 & n3758;
  assign n3760 = ~n427 & n3759;
  assign n3761 = ~n705 & n3760;
  assign n3762 = n1892 & n1931;
  assign n3763 = ~n383 & n3762;
  assign n3764 = ~n344 & n3763;
  assign n3765 = n3761 & n3764;
  assign n3766 = n3231 & n3765;
  assign n3767 = n3757 & n3766;
  assign n3768 = n467 & n3767;
  assign n3769 = ~n255 & n3768;
  assign n3770 = ~n424 & ~n475;
  assign n3771 = ~n193 & n3770;
  assign n3772 = ~n666 & n1577;
  assign n3773 = ~n106 & n3772;
  assign n3774 = ~n362 & n1635;
  assign n3775 = ~n216 & n3774;
  assign n3776 = n3773 & n3775;
  assign n3777 = ~n576 & n1163;
  assign n3778 = ~n235 & n3777;
  assign n3779 = ~n373 & ~n700;
  assign n3780 = ~n114 & n3779;
  assign n3781 = n3778 & n3780;
  assign n3782 = n3776 & n3781;
  assign n3783 = n3771 & n3782;
  assign n3784 = ~n469 & n3783;
  assign n3785 = ~n689 & n3784;
  assign n3786 = n3769 & n3785;
  assign n3787 = n1327 & n1451;
  assign n3788 = n680 & n3787;
  assign n3789 = n822 & n3788;
  assign n3790 = ~n305 & ~n533;
  assign n3791 = ~n254 & n3790;
  assign n3792 = n1617 & n3791;
  assign n3793 = ~n580 & n3792;
  assign n3794 = n1791 & n3020;
  assign n3795 = ~n260 & n3794;
  assign n3796 = n3793 & n3795;
  assign n3797 = ~n637 & n2771;
  assign n3798 = n2883 & n3797;
  assign n3799 = n1343 & n3798;
  assign n3800 = ~n278 & n3799;
  assign n3801 = n3000 & n3695;
  assign n3802 = n1435 & n3801;
  assign n3803 = ~n600 & n3802;
  assign n3804 = ~n633 & n3803;
  assign n3805 = n3800 & n3804;
  assign n3806 = n3796 & n3805;
  assign n3807 = ~n155 & ~n400;
  assign n3808 = ~n219 & n3807;
  assign n3809 = n3806 & n3808;
  assign n3810 = n3789 & n3809;
  assign n3811 = ~n123 & n3810;
  assign n3812 = ~n272 & n3811;
  assign n3813 = ~n536 & n694;
  assign n3814 = ~n501 & n3813;
  assign n3815 = n3812 & n3814;
  assign n3816 = n3786 & n3815;
  assign n3817 = n3713 & ~n3816;
  assign n3818 = ~n3713 & n3816;
  assign n3819 = ~n3817 & ~n3818;
  assign n3820 = ~n362 & ~n583;
  assign n3821 = ~n422 & n2436;
  assign n3822 = ~n363 & ~n373;
  assign n3823 = n1214 & n3822;
  assign n3824 = ~n117 & n1490;
  assign n3825 = ~n428 & n3824;
  assign n3826 = ~n180 & ~n320;
  assign n3827 = ~n544 & n3826;
  assign n3828 = n3825 & n3827;
  assign n3829 = n3823 & n3828;
  assign n3830 = n3821 & n3829;
  assign n3831 = n930 & n3830;
  assign n3832 = n2648 & n3831;
  assign n3833 = n3820 & n3832;
  assign n3834 = ~n273 & n3833;
  assign n3835 = ~n165 & ~n697;
  assign n3836 = ~n236 & n3835;
  assign n3837 = n3202 & n3836;
  assign n3838 = n562 & n3837;
  assign n3839 = n459 & n3838;
  assign n3840 = n901 & n3839;
  assign n3841 = ~n131 & n3840;
  assign n3842 = n3834 & n3841;
  assign n3843 = ~n170 & ~n238;
  assign n3844 = ~n398 & n3843;
  assign n3845 = ~n289 & ~n594;
  assign n3846 = ~n611 & n3845;
  assign n3847 = ~n321 & n3846;
  assign n3848 = ~n280 & n3847;
  assign n3849 = n3844 & n3848;
  assign n3850 = n1388 & n3849;
  assign n3851 = n706 & n3850;
  assign n3852 = ~n123 & n3851;
  assign n3853 = ~n195 & ~n354;
  assign n3854 = ~n666 & ~n701;
  assign n3855 = ~n305 & n3854;
  assign n3856 = ~n441 & n3855;
  assign n3857 = n3853 & n3856;
  assign n3858 = ~n81 & n3857;
  assign n3859 = ~n502 & ~n628;
  assign n3860 = ~n454 & n3859;
  assign n3861 = ~n122 & n3860;
  assign n3862 = ~n581 & n3861;
  assign n3863 = ~n439 & n3862;
  assign n3864 = n3858 & n3863;
  assign n3865 = n3412 & n3864;
  assign n3866 = ~n381 & n3865;
  assign n3867 = ~n132 & ~n633;
  assign n3868 = ~n372 & n3808;
  assign n3869 = ~n593 & n3868;
  assign n3870 = n3867 & n3869;
  assign n3871 = n2060 & n3870;
  assign n3872 = ~n152 & n3871;
  assign n3873 = ~n288 & n3872;
  assign n3874 = n3866 & n3873;
  assign n3875 = ~n576 & ~n600;
  assign n3876 = ~n590 & n3875;
  assign n3877 = ~n342 & n3876;
  assign n3878 = ~n683 & n3877;
  assign n3879 = n1340 & n1343;
  assign n3880 = n2680 & n3879;
  assign n3881 = n3878 & n3880;
  assign n3882 = n3874 & n3881;
  assign n3883 = n2350 & n3882;
  assign n3884 = ~n393 & n3883;
  assign n3885 = ~n668 & n3884;
  assign n3886 = n3852 & n3885;
  assign n3887 = n3842 & n3886;
  assign n3888 = ~n455 & n673;
  assign n3889 = ~n218 & n3888;
  assign n3890 = ~n384 & n3889;
  assign n3891 = n2321 & n3890;
  assign n3892 = n3429 & n3891;
  assign n3893 = n1079 & n3892;
  assign n3894 = n3138 & n3893;
  assign n3895 = ~n430 & n3894;
  assign n3896 = ~n161 & ~n216;
  assign n3897 = ~n131 & ~n465;
  assign n3898 = ~n610 & n3897;
  assign n3899 = ~n172 & n3898;
  assign n3900 = n3896 & n3899;
  assign n3901 = n1057 & n3900;
  assign n3902 = ~n697 & n3901;
  assign n3903 = n3895 & n3902;
  assign n3904 = ~n353 & n515;
  assign n3905 = ~n150 & n3904;
  assign n3906 = ~n527 & n3905;
  assign n3907 = ~n458 & n3906;
  assign n3908 = ~n290 & n3907;
  assign n3909 = ~n94 & n1076;
  assign n3910 = ~n372 & ~n423;
  assign n3911 = ~n195 & n3910;
  assign n3912 = ~n100 & n3911;
  assign n3913 = ~n152 & n3912;
  assign n3914 = n3909 & n3913;
  assign n3915 = n1132 & n3914;
  assign n3916 = n3908 & n3915;
  assign n3917 = n1285 & n3916;
  assign n3918 = ~n424 & n3917;
  assign n3919 = ~n116 & ~n391;
  assign n3920 = n596 & n3919;
  assign n3921 = ~n345 & n2199;
  assign n3922 = ~n261 & ~n341;
  assign n3923 = n3921 & n3922;
  assign n3924 = ~n281 & n3923;
  assign n3925 = ~n247 & n2417;
  assign n3926 = ~n621 & n3925;
  assign n3927 = n3924 & n3926;
  assign n3928 = n1401 & n3927;
  assign n3929 = n3920 & n3928;
  assign n3930 = ~n631 & n3929;
  assign n3931 = ~n466 & n3930;
  assign n3932 = ~n122 & n1232;
  assign n3933 = ~n544 & n3932;
  assign n3934 = n3931 & n3933;
  assign n3935 = ~n332 & ~n700;
  assign n3936 = ~n454 & n3935;
  assign n3937 = n1024 & n3936;
  assign n3938 = ~n204 & n3937;
  assign n3939 = ~n637 & n3938;
  assign n3940 = n1575 & n2180;
  assign n3941 = ~n518 & n3940;
  assign n3942 = ~n580 & n3941;
  assign n3943 = n3939 & n3942;
  assign n3944 = n3934 & n3943;
  assign n3945 = n1395 & n3944;
  assign n3946 = ~n129 & n3945;
  assign n3947 = n3918 & n3946;
  assign n3948 = n3903 & n3947;
  assign n3949 = ~n3887 & ~n3948;
  assign n3950 = n3887 & n3948;
  assign n3951 = ~n3949 & ~n3950;
  assign n3952 = ~pi26  & n3951;
  assign n3953 = ~n3949 & ~n3952;
  assign n3954 = n3816 & ~n3953;
  assign n3955 = ~n3816 & n3953;
  assign n3956 = ~n894 & n3641;
  assign n3957 = ~n795 & n3740;
  assign n3958 = n3625 & ~n3627;
  assign n3959 = ~n3628 & ~n3958;
  assign n3960 = n556 & n3959;
  assign n3961 = ~pi31  & ~n555;
  assign n3962 = ~n665 & n3961;
  assign n3963 = ~n3960 & ~n3962;
  assign n3964 = ~n3957 & n3963;
  assign n3965 = ~n3956 & n3964;
  assign n3966 = ~n3955 & ~n3965;
  assign n3967 = ~n3954 & ~n3966;
  assign n3968 = n3819 & ~n3967;
  assign n3969 = ~n3817 & ~n3968;
  assign n3970 = ~pi29  & ~n3732;
  assign n3971 = ~n3730 & n3733;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = ~n3969 & ~n3972;
  assign n3974 = n3969 & n3972;
  assign n3975 = ~n3973 & ~n3974;
  assign n3976 = ~n665 & n3641;
  assign n3977 = ~n720 & n3740;
  assign n3978 = n3633 & ~n3636;
  assign n3979 = ~n3637 & ~n3978;
  assign n3980 = n556 & n3979;
  assign n3981 = ~n554 & n3961;
  assign n3982 = ~n3980 & ~n3981;
  assign n3983 = ~n3977 & n3982;
  assign n3984 = ~n3976 & n3983;
  assign n3985 = n3975 & ~n3984;
  assign n3986 = ~n3973 & ~n3985;
  assign n3987 = ~n3734 & ~n3735;
  assign n3988 = ~n3747 & n3987;
  assign n3989 = n3747 & ~n3987;
  assign n3990 = ~n3988 & ~n3989;
  assign n3991 = ~n3986 & n3990;
  assign n3992 = n3986 & ~n3990;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = ~n3975 & n3984;
  assign n3995 = ~n3985 & ~n3994;
  assign n3996 = pi26  & ~pi27 ;
  assign n3997 = ~pi26  & pi27 ;
  assign n3998 = ~n3996 & ~n3997;
  assign n3999 = pi28  & ~pi29 ;
  assign n4000 = ~pi28  & pi29 ;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = ~n3998 & ~n4001;
  assign n4003 = ~n3638 & n4002;
  assign n4004 = ~n72 & ~n96;
  assign n4005 = n3998 & ~n4004;
  assign n4006 = ~n4001 & n4005;
  assign n4007 = ~n4003 & ~n4006;
  assign n4008 = ~n554 & ~n4007;
  assign n4009 = ~pi29  & n4008;
  assign n4010 = pi29  & ~n4008;
  assign n4011 = ~n4009 & ~n4010;
  assign n4012 = ~n795 & n3641;
  assign n4013 = ~n665 & n3740;
  assign n4014 = n3629 & ~n3631;
  assign n4015 = ~n3632 & ~n4014;
  assign n4016 = n556 & n4015;
  assign n4017 = ~n720 & n3961;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = ~n4013 & n4018;
  assign n4020 = ~n4012 & n4019;
  assign n4021 = n4011 & n4020;
  assign n4022 = ~n4011 & ~n4020;
  assign n4023 = ~n3819 & n3967;
  assign n4024 = ~n3968 & ~n4023;
  assign n4025 = ~n4022 & ~n4024;
  assign n4026 = ~n4021 & ~n4025;
  assign n4027 = n3995 & n4026;
  assign n4028 = ~n3954 & ~n3955;
  assign n4029 = ~n3965 & n4028;
  assign n4030 = n3965 & ~n4028;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = n549 & n3919;
  assign n4033 = n753 & n4032;
  assign n4034 = n558 & n4033;
  assign n4035 = ~n527 & n4034;
  assign n4036 = ~n299 & ~n350;
  assign n4037 = ~n399 & n4036;
  assign n4038 = n1109 & n4037;
  assign n4039 = ~n545 & n4038;
  assign n4040 = n4035 & n4039;
  assign n4041 = ~n695 & n4040;
  assign n4042 = ~n256 & n459;
  assign n4043 = ~n579 & n4042;
  assign n4044 = ~n331 & n1600;
  assign n4045 = ~n260 & n4044;
  assign n4046 = n4043 & n4045;
  assign n4047 = ~n669 & n4046;
  assign n4048 = ~n345 & ~n689;
  assign n4049 = ~n428 & n4048;
  assign n4050 = ~n155 & n221;
  assign n4051 = ~n442 & n4050;
  assign n4052 = n4049 & n4051;
  assign n4053 = n4047 & n4052;
  assign n4054 = n488 & n1461;
  assign n4055 = ~n252 & n4054;
  assign n4056 = n2064 & n2280;
  assign n4057 = ~n394 & n4056;
  assign n4058 = n4055 & n4057;
  assign n4059 = ~n232 & n4058;
  assign n4060 = ~n94 & ~n259;
  assign n4061 = ~n672 & n4060;
  assign n4062 = n167 & n907;
  assign n4063 = ~n413 & n4062;
  assign n4064 = n4061 & n4063;
  assign n4065 = n4059 & n4064;
  assign n4066 = n237 & n4065;
  assign n4067 = ~n231 & n4066;
  assign n4068 = ~n670 & n4067;
  assign n4069 = ~n400 & ~n576;
  assign n4070 = ~n294 & n4069;
  assign n4071 = ~n278 & ~n455;
  assign n4072 = ~n217 & n4071;
  assign n4073 = n4070 & n4072;
  assign n4074 = ~n341 & n4073;
  assign n4075 = ~n395 & n4074;
  assign n4076 = ~n344 & n4075;
  assign n4077 = n4068 & n4076;
  assign n4078 = ~n288 & ~n414;
  assign n4079 = ~n357 & n4078;
  assign n4080 = ~n692 & n4079;
  assign n4081 = ~n422 & n4080;
  assign n4082 = ~n374 & n4081;
  assign n4083 = ~n262 & ~n593;
  assign n4084 = ~n163 & n4083;
  assign n4085 = ~n600 & ~n639;
  assign n4086 = n4084 & n4085;
  assign n4087 = ~n310 & n4086;
  assign n4088 = ~n631 & n2904;
  assign n4089 = ~n238 & n4088;
  assign n4090 = n4087 & n4089;
  assign n4091 = n2335 & n4090;
  assign n4092 = ~n122 & n4091;
  assign n4093 = ~n477 & n4092;
  assign n4094 = ~n621 & n4093;
  assign n4095 = n4082 & n4094;
  assign n4096 = n4077 & n4095;
  assign n4097 = n2494 & n4096;
  assign n4098 = ~n188 & n4097;
  assign n4099 = n4053 & n4098;
  assign n4100 = n4041 & n4099;
  assign n4101 = n3887 & ~n4100;
  assign n4102 = ~n3887 & n4100;
  assign n4103 = ~n1107 & n3641;
  assign n4104 = ~n1005 & n3740;
  assign n4105 = n3617 & ~n3619;
  assign n4106 = ~n3620 & ~n4105;
  assign n4107 = n556 & n4106;
  assign n4108 = ~n894 & n3961;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = ~n4104 & n4109;
  assign n4111 = ~n4103 & n4110;
  assign n4112 = ~n4102 & ~n4111;
  assign n4113 = ~n4101 & ~n4112;
  assign n4114 = ~pi26  & ~n3952;
  assign n4115 = ~n3950 & n3953;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = ~n4113 & ~n4116;
  assign n4118 = n4113 & n4116;
  assign n4119 = ~n1005 & n3641;
  assign n4120 = ~n894 & n3740;
  assign n4121 = n3621 & ~n3623;
  assign n4122 = ~n3624 & ~n4121;
  assign n4123 = n556 & n4122;
  assign n4124 = ~n795 & n3961;
  assign n4125 = ~n4123 & ~n4124;
  assign n4126 = ~n4120 & n4125;
  assign n4127 = ~n4119 & n4126;
  assign n4128 = ~n4118 & ~n4127;
  assign n4129 = ~n4117 & ~n4128;
  assign n4130 = n4031 & ~n4129;
  assign n4131 = ~n4031 & n4129;
  assign n4132 = ~n3744 & n4002;
  assign n4133 = n3998 & n4004;
  assign n4134 = ~n554 & n4133;
  assign n4135 = ~n720 & n4006;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = ~n4132 & n4136;
  assign n4138 = pi29  & n4137;
  assign n4139 = ~pi29  & ~n4137;
  assign n4140 = ~n4138 & ~n4139;
  assign n4141 = ~n4131 & ~n4140;
  assign n4142 = ~n4130 & ~n4141;
  assign n4143 = ~n4021 & ~n4022;
  assign n4144 = ~n4024 & n4143;
  assign n4145 = n4024 & ~n4143;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = ~n4142 & ~n4146;
  assign n4148 = ~n4101 & ~n4102;
  assign n4149 = ~n4111 & n4148;
  assign n4150 = n4111 & ~n4148;
  assign n4151 = ~n4149 & ~n4150;
  assign n4152 = ~n181 & ~n469;
  assign n4153 = ~n672 & n4152;
  assign n4154 = ~n150 & ~n589;
  assign n4155 = n4153 & n4154;
  assign n4156 = n519 & n4155;
  assign n4157 = ~n527 & n4156;
  assign n4158 = ~n304 & n2724;
  assign n4159 = ~n372 & n4158;
  assign n4160 = ~n85 & ~n117;
  assign n4161 = ~n160 & n4160;
  assign n4162 = n4159 & n4161;
  assign n4163 = n2683 & n4162;
  assign n4164 = ~n280 & n4163;
  assign n4165 = ~n612 & n4164;
  assign n4166 = n4157 & n4165;
  assign n4167 = ~n261 & n2218;
  assign n4168 = ~n173 & n4167;
  assign n4169 = n1670 & n4168;
  assign n4170 = n3114 & n4169;
  assign n4171 = n2180 & n4170;
  assign n4172 = ~n576 & n4171;
  assign n4173 = ~n506 & n3277;
  assign n4174 = ~n106 & n4173;
  assign n4175 = ~n171 & ~n334;
  assign n4176 = ~n206 & n4175;
  assign n4177 = ~n613 & n4176;
  assign n4178 = ~n326 & n2248;
  assign n4179 = ~n667 & n4178;
  assign n4180 = n4177 & n4179;
  assign n4181 = ~n275 & n1141;
  assign n4182 = ~n636 & n4181;
  assign n4183 = ~n697 & n1301;
  assign n4184 = ~n464 & n4183;
  assign n4185 = ~n115 & n4184;
  assign n4186 = n4182 & n4185;
  assign n4187 = n4180 & n4186;
  assign n4188 = n1348 & n4187;
  assign n4189 = ~n633 & n4188;
  assign n4190 = ~n251 & n4189;
  assign n4191 = n4174 & n4190;
  assign n4192 = ~n203 & n467;
  assign n4193 = ~n294 & n1112;
  assign n4194 = ~n362 & ~n535;
  assign n4195 = n4193 & n4194;
  assign n4196 = ~n337 & n4195;
  assign n4197 = ~n144 & ~n298;
  assign n4198 = ~n593 & n4197;
  assign n4199 = ~n245 & n4198;
  assign n4200 = n4196 & n4199;
  assign n4201 = n4192 & n4200;
  assign n4202 = ~n534 & n4201;
  assign n4203 = ~n461 & ~n682;
  assign n4204 = n3896 & n4203;
  assign n4205 = ~n681 & n4204;
  assign n4206 = n237 & ~n422;
  assign n4207 = ~n134 & n4206;
  assign n4208 = n4205 & n4207;
  assign n4209 = ~n427 & n4208;
  assign n4210 = ~n214 & n4209;
  assign n4211 = n4202 & n4210;
  assign n4212 = n4191 & n4211;
  assign n4213 = n2120 & n4212;
  assign n4214 = ~n232 & n4213;
  assign n4215 = ~n277 & n4214;
  assign n4216 = n4172 & n4215;
  assign n4217 = n4166 & n4216;
  assign n4218 = n2306 & n2417;
  assign n4219 = n1791 & n4218;
  assign n4220 = ~n245 & n4219;
  assign n4221 = n1622 & n3906;
  assign n4222 = n1652 & n4221;
  assign n4223 = ~n435 & n4222;
  assign n4224 = ~n704 & n4223;
  assign n4225 = n4220 & n4224;
  assign n4226 = ~n305 & n445;
  assign n4227 = ~n611 & n4226;
  assign n4228 = n358 & n1978;
  assign n4229 = n4227 & n4228;
  assign n4230 = n1241 & n2070;
  assign n4231 = n4229 & n4230;
  assign n4232 = ~n114 & n4231;
  assign n4233 = ~n612 & n2772;
  assign n4234 = ~n579 & n4233;
  assign n4235 = ~n400 & n4234;
  assign n4236 = n4232 & n4235;
  assign n4237 = n4225 & n4236;
  assign n4238 = ~n172 & ~n534;
  assign n4239 = n89 & n1657;
  assign n4240 = n920 & n4239;
  assign n4241 = ~n170 & n4240;
  assign n4242 = ~n134 & ~n272;
  assign n4243 = ~n94 & n4242;
  assign n4244 = n1490 & n4243;
  assign n4245 = n282 & n4244;
  assign n4246 = ~n457 & n4245;
  assign n4247 = n4241 & n4246;
  assign n4248 = n1015 & n3876;
  assign n4249 = ~n238 & ~n252;
  assign n4250 = ~n262 & n4249;
  assign n4251 = ~n672 & n4250;
  assign n4252 = n754 & n4251;
  assign n4253 = ~n538 & n4252;
  assign n4254 = n4248 & n4253;
  assign n4255 = n4247 & n4254;
  assign n4256 = n4238 & n4255;
  assign n4257 = n4237 & n4256;
  assign n4258 = ~n697 & n4257;
  assign n4259 = ~n463 & n4258;
  assign n4260 = ~n506 & ~n581;
  assign n4261 = ~n685 & n2281;
  assign n4262 = ~n155 & ~n477;
  assign n4263 = n4261 & n4262;
  assign n4264 = ~n610 & n4263;
  assign n4265 = ~n385 & n3693;
  assign n4266 = ~n598 & n4265;
  assign n4267 = n4264 & n4266;
  assign n4268 = n4260 & n4267;
  assign n4269 = ~n206 & n4268;
  assign n4270 = ~n187 & n4269;
  assign n4271 = n4259 & n4270;
  assign n4272 = ~n362 & n1268;
  assign n4273 = ~n423 & n4272;
  assign n4274 = ~n207 & n4273;
  assign n4275 = ~n669 & n1252;
  assign n4276 = ~n626 & n4275;
  assign n4277 = n2929 & n4276;
  assign n4278 = n4274 & n4277;
  assign n4279 = ~n161 & ~n613;
  assign n4280 = n221 & n4279;
  assign n4281 = ~n374 & n3309;
  assign n4282 = n4280 & n4281;
  assign n4283 = n4278 & n4282;
  assign n4284 = n1962 & n4283;
  assign n4285 = ~n298 & n4284;
  assign n4286 = ~n308 & n4285;
  assign n4287 = ~n390 & ~n667;
  assign n4288 = ~n632 & n4287;
  assign n4289 = ~n537 & n4288;
  assign n4290 = n1356 & n4289;
  assign n4291 = n1676 & n4290;
  assign n4292 = ~n631 & n4291;
  assign n4293 = ~n461 & n4292;
  assign n4294 = ~n670 & n4293;
  assign n4295 = n4286 & n4294;
  assign n4296 = n4271 & n4295;
  assign n4297 = ~n4217 & ~n4296;
  assign n4298 = n4217 & n4296;
  assign n4299 = ~n4297 & ~n4298;
  assign n4300 = ~pi23  & n4299;
  assign n4301 = ~n4297 & ~n4300;
  assign n4302 = ~n3887 & n4301;
  assign n4303 = n3887 & ~n4301;
  assign n4304 = ~n1230 & n3641;
  assign n4305 = ~n1107 & n3740;
  assign n4306 = n3613 & ~n3615;
  assign n4307 = ~n3616 & ~n4306;
  assign n4308 = n556 & n4307;
  assign n4309 = ~n1005 & n3961;
  assign n4310 = ~n4308 & ~n4309;
  assign n4311 = ~n4305 & n4310;
  assign n4312 = ~n4304 & n4311;
  assign n4313 = ~n4303 & n4312;
  assign n4314 = ~n4302 & ~n4313;
  assign n4315 = n4151 & n4314;
  assign n4316 = ~n4151 & ~n4314;
  assign n4317 = ~n4315 & ~n4316;
  assign n4318 = ~pi23  & ~n4300;
  assign n4319 = ~n4298 & n4301;
  assign n4320 = ~n4318 & ~n4319;
  assign n4321 = ~n1338 & n3641;
  assign n4322 = n3609 & ~n3611;
  assign n4323 = ~n3612 & ~n4322;
  assign n4324 = n556 & n4323;
  assign n4325 = ~n1107 & n3961;
  assign n4326 = ~n1230 & n3740;
  assign n4327 = ~n4325 & ~n4326;
  assign n4328 = ~n4324 & n4327;
  assign n4329 = ~n4321 & n4328;
  assign n4330 = ~n4320 & ~n4329;
  assign n4331 = n4320 & n4329;
  assign n4332 = ~n4330 & ~n4331;
  assign n4333 = ~n279 & ~n589;
  assign n4334 = ~n281 & n4333;
  assign n4335 = n2132 & n4334;
  assign n4336 = ~n579 & n4335;
  assign n4337 = ~n204 & ~n261;
  assign n4338 = ~n639 & n4337;
  assign n4339 = n4336 & n4338;
  assign n4340 = n2191 & n4339;
  assign n4341 = ~n580 & n4340;
  assign n4342 = n1451 & n1763;
  assign n4343 = n1446 & n4342;
  assign n4344 = n1641 & n4343;
  assign n4345 = ~n682 & n4344;
  assign n4346 = n4341 & n4345;
  assign n4347 = ~n180 & n857;
  assign n4348 = n107 & n759;
  assign n4349 = ~n363 & ~n700;
  assign n4350 = ~n545 & n4349;
  assign n4351 = n1401 & n4350;
  assign n4352 = n4348 & n4351;
  assign n4353 = ~n298 & ~n671;
  assign n4354 = ~n342 & ~n621;
  assign n4355 = n4353 & n4354;
  assign n4356 = ~n144 & n4355;
  assign n4357 = ~n206 & n3414;
  assign n4358 = ~n147 & n4357;
  assign n4359 = ~n323 & ~n535;
  assign n4360 = ~n372 & n4359;
  assign n4361 = n746 & n4360;
  assign n4362 = n4358 & n4361;
  assign n4363 = n881 & n4362;
  assign n4364 = n445 & n4363;
  assign n4365 = ~n278 & n4364;
  assign n4366 = n4356 & n4365;
  assign n4367 = n4352 & n4366;
  assign n4368 = n4347 & n4367;
  assign n4369 = n3029 & n4368;
  assign n4370 = ~n629 & n4369;
  assign n4371 = ~n88 & ~n678;
  assign n4372 = n758 & n4371;
  assign n4373 = ~n693 & n4372;
  assign n4374 = n1417 & n4373;
  assign n4375 = n1148 & n4374;
  assign n4376 = ~n305 & n4375;
  assign n4377 = ~n429 & n4376;
  assign n4378 = n4370 & n4377;
  assign n4379 = n4346 & n4378;
  assign n4380 = ~n4217 & n4379;
  assign n4381 = n4217 & ~n4379;
  assign n4382 = ~n217 & n2991;
  assign n4383 = ~n171 & n702;
  assign n4384 = ~n160 & n4383;
  assign n4385 = n4382 & n4384;
  assign n4386 = n955 & n4385;
  assign n4387 = n291 & n4386;
  assign n4388 = n107 & n2133;
  assign n4389 = ~n454 & n4388;
  assign n4390 = n4387 & n4389;
  assign n4391 = ~n372 & n3038;
  assign n4392 = n822 & n4391;
  assign n4393 = ~n545 & n4392;
  assign n4394 = n897 & n3470;
  assign n4395 = n2180 & n4394;
  assign n4396 = ~n81 & n4395;
  assign n4397 = n4393 & n4396;
  assign n4398 = n4390 & n4397;
  assign n4399 = n2316 & n4398;
  assign n4400 = ~n477 & n4399;
  assign n4401 = n3791 & n4371;
  assign n4402 = ~n195 & ~n537;
  assign n4403 = ~n353 & n1131;
  assign n4404 = ~n666 & n1670;
  assign n4405 = ~n468 & n4404;
  assign n4406 = n4403 & n4405;
  assign n4407 = n4402 & n4406;
  assign n4408 = n4401 & n4407;
  assign n4409 = n459 & n1447;
  assign n4410 = n4408 & n4409;
  assign n4411 = ~n466 & n4410;
  assign n4412 = ~n375 & n2585;
  assign n4413 = ~n277 & n4412;
  assign n4414 = ~n505 & n4413;
  assign n4415 = n4411 & n4414;
  assign n4416 = ~n122 & n4334;
  assign n4417 = ~n633 & n4416;
  assign n4418 = n725 & n2653;
  assign n4419 = ~n255 & n4418;
  assign n4420 = ~n132 & n4419;
  assign n4421 = n4417 & n4420;
  assign n4422 = n4415 & n4421;
  assign n4423 = n1494 & n1785;
  assign n4424 = n1116 & n4423;
  assign n4425 = n4422 & n4424;
  assign n4426 = n2772 & n4425;
  assign n4427 = n615 & n1576;
  assign n4428 = ~n612 & n4427;
  assign n4429 = n1959 & n4428;
  assign n4430 = n2060 & n4429;
  assign n4431 = n4426 & n4430;
  assign n4432 = n1464 & n4431;
  assign n4433 = ~n631 & n4432;
  assign n4434 = ~n357 & n4433;
  assign n4435 = n4400 & n4434;
  assign n4436 = ~n304 & n4435;
  assign n4437 = ~n161 & n1368;
  assign n4438 = ~n501 & n4437;
  assign n4439 = n4436 & n4438;
  assign n4440 = n1112 & n3056;
  assign n4441 = n233 & n1166;
  assign n4442 = n1641 & n4441;
  assign n4443 = ~n373 & n4442;
  assign n4444 = ~n458 & ~n594;
  assign n4445 = n1924 & n4444;
  assign n4446 = n954 & n4445;
  assign n4447 = ~n692 & n4446;
  assign n4448 = n4443 & n4447;
  assign n4449 = ~n331 & n1744;
  assign n4450 = ~n246 & n3442;
  assign n4451 = ~n344 & n4450;
  assign n4452 = n4449 & n4451;
  assign n4453 = n1964 & n4452;
  assign n4454 = ~n298 & n4453;
  assign n4455 = ~n672 & n4260;
  assign n4456 = ~n188 & n4455;
  assign n4457 = n3030 & n4456;
  assign n4458 = n758 & n4457;
  assign n4459 = n415 & n4458;
  assign n4460 = n1368 & n4459;
  assign n4461 = ~n633 & n4460;
  assign n4462 = n4454 & n4461;
  assign n4463 = n4448 & n4462;
  assign n4464 = n992 & n4463;
  assign n4465 = n4440 & n4464;
  assign n4466 = ~n441 & n4465;
  assign n4467 = ~n700 & n4466;
  assign n4468 = ~n259 & ~n579;
  assign n4469 = ~n679 & n4468;
  assign n4470 = n1253 & n4469;
  assign n4471 = ~n129 & n4470;
  assign n4472 = ~n197 & n1478;
  assign n4473 = n1708 & n4472;
  assign n4474 = ~n98 & n4473;
  assign n4475 = n4471 & n4474;
  assign n4476 = ~n326 & n546;
  assign n4477 = ~n668 & n4476;
  assign n4478 = ~n256 & n852;
  assign n4479 = ~n610 & n4478;
  assign n4480 = n4477 & n4479;
  assign n4481 = ~n305 & n1482;
  assign n4482 = ~n391 & n4481;
  assign n4483 = ~n161 & ~n186;
  assign n4484 = ~n442 & n4483;
  assign n4485 = n4482 & n4484;
  assign n4486 = n4480 & n4485;
  assign n4487 = n1232 & n4486;
  assign n4488 = ~n309 & n4487;
  assign n4489 = n2066 & n2286;
  assign n4490 = ~n537 & n4489;
  assign n4491 = n4488 & n4490;
  assign n4492 = n4475 & n4491;
  assign n4493 = ~n395 & n456;
  assign n4494 = ~n505 & n3187;
  assign n4495 = n4493 & n4494;
  assign n4496 = ~n474 & n4495;
  assign n4497 = ~n217 & ~n299;
  assign n4498 = ~n252 & n4497;
  assign n4499 = ~n427 & n4498;
  assign n4500 = ~n219 & n4499;
  assign n4501 = n4496 & n4500;
  assign n4502 = n4492 & n4501;
  assign n4503 = n1388 & n4502;
  assign n4504 = ~n100 & n4503;
  assign n4505 = ~n131 & ~n637;
  assign n4506 = ~n614 & n4505;
  assign n4507 = ~n320 & n4506;
  assign n4508 = ~n289 & n4507;
  assign n4509 = ~n517 & n4508;
  assign n4510 = ~n279 & n691;
  assign n4511 = ~n307 & n4510;
  assign n4512 = ~n214 & n4511;
  assign n4513 = ~n104 & ~n533;
  assign n4514 = ~n382 & n4513;
  assign n4515 = n4512 & n4514;
  assign n4516 = ~n671 & n4515;
  assign n4517 = n4509 & n4516;
  assign n4518 = n1577 & n4517;
  assign n4519 = ~n468 & n4518;
  assign n4520 = n4504 & n4519;
  assign n4521 = n1011 & n4520;
  assign n4522 = n4467 & n4521;
  assign n4523 = ~n4439 & ~n4522;
  assign n4524 = n4439 & n4522;
  assign n4525 = ~n4523 & ~n4524;
  assign n4526 = ~pi20  & n4525;
  assign n4527 = ~n4523 & ~n4526;
  assign n4528 = ~n4379 & n4527;
  assign n4529 = n4379 & ~n4527;
  assign n4530 = ~n1531 & n3641;
  assign n4531 = ~n1426 & n3740;
  assign n4532 = n3601 & ~n3603;
  assign n4533 = ~n3604 & ~n4532;
  assign n4534 = n556 & n4533;
  assign n4535 = ~n1338 & n3961;
  assign n4536 = ~n4534 & ~n4535;
  assign n4537 = ~n4531 & n4536;
  assign n4538 = ~n4530 & n4537;
  assign n4539 = ~n4529 & n4538;
  assign n4540 = ~n4528 & ~n4539;
  assign n4541 = ~n4381 & ~n4540;
  assign n4542 = ~n4380 & ~n4541;
  assign n4543 = n4332 & n4542;
  assign n4544 = ~n4330 & ~n4543;
  assign n4545 = ~n4302 & ~n4303;
  assign n4546 = ~n4312 & n4545;
  assign n4547 = n4312 & ~n4545;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = ~n4544 & n4548;
  assign n4550 = n4544 & ~n4548;
  assign n4551 = ~n4549 & ~n4550;
  assign n4552 = ~n894 & n4006;
  assign n4553 = ~n795 & n4133;
  assign n4554 = n3959 & n4002;
  assign n4555 = ~n3998 & n4001;
  assign n4556 = ~n665 & n4555;
  assign n4557 = ~n4554 & ~n4556;
  assign n4558 = ~n4553 & n4557;
  assign n4559 = ~n4552 & n4558;
  assign n4560 = pi29  & n4559;
  assign n4561 = ~pi29  & ~n4559;
  assign n4562 = ~n4560 & ~n4561;
  assign n4563 = n4551 & ~n4562;
  assign n4564 = ~n4549 & ~n4563;
  assign n4565 = n4317 & ~n4564;
  assign n4566 = ~n4315 & ~n4565;
  assign n4567 = ~n4117 & ~n4118;
  assign n4568 = ~n4127 & n4567;
  assign n4569 = n4127 & ~n4567;
  assign n4570 = ~n4568 & ~n4569;
  assign n4571 = ~n4566 & n4570;
  assign n4572 = ~n665 & n4006;
  assign n4573 = ~n720 & n4133;
  assign n4574 = n3979 & n4002;
  assign n4575 = ~n554 & n4555;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = ~n4573 & n4576;
  assign n4578 = ~n4572 & n4577;
  assign n4579 = pi29  & n4578;
  assign n4580 = ~pi29  & ~n4578;
  assign n4581 = ~n4579 & ~n4580;
  assign n4582 = n4566 & ~n4570;
  assign n4583 = ~n4571 & ~n4582;
  assign n4584 = ~n4581 & n4583;
  assign n4585 = ~n4571 & ~n4584;
  assign n4586 = ~n4130 & ~n4131;
  assign n4587 = ~n4140 & n4586;
  assign n4588 = n4140 & ~n4586;
  assign n4589 = ~n4587 & ~n4588;
  assign n4590 = ~n4585 & n4589;
  assign n4591 = n4585 & ~n4589;
  assign n4592 = ~n4590 & ~n4591;
  assign n4593 = pi25  & ~pi26 ;
  assign n4594 = ~pi25  & pi26 ;
  assign n4595 = ~n4593 & ~n4594;
  assign n4596 = pi23  & ~pi24 ;
  assign n4597 = ~pi23  & pi24 ;
  assign n4598 = ~n4596 & ~n4597;
  assign n4599 = ~n76 & ~n82;
  assign n4600 = n4598 & ~n4599;
  assign n4601 = ~n4595 & n4600;
  assign n4602 = ~n4595 & ~n4598;
  assign n4603 = ~n3638 & n4602;
  assign n4604 = ~n4601 & ~n4603;
  assign n4605 = ~n554 & ~n4604;
  assign n4606 = ~pi26  & n4605;
  assign n4607 = pi26  & ~n4605;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = ~n795 & n4006;
  assign n4610 = ~n665 & n4133;
  assign n4611 = n4002 & n4015;
  assign n4612 = ~n720 & n4555;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 = ~n4610 & n4613;
  assign n4615 = ~n4609 & n4614;
  assign n4616 = pi29  & n4615;
  assign n4617 = ~pi29  & ~n4615;
  assign n4618 = ~n4616 & ~n4617;
  assign n4619 = ~n4608 & ~n4618;
  assign n4620 = ~n4317 & n4564;
  assign n4621 = ~n4565 & ~n4620;
  assign n4622 = n4608 & n4618;
  assign n4623 = ~n4619 & ~n4622;
  assign n4624 = n4621 & n4623;
  assign n4625 = ~n4619 & ~n4624;
  assign n4626 = n4581 & ~n4583;
  assign n4627 = ~n4584 & ~n4626;
  assign n4628 = ~n4625 & n4627;
  assign n4629 = ~n4551 & n4562;
  assign n4630 = ~n4563 & ~n4629;
  assign n4631 = ~n4528 & ~n4529;
  assign n4632 = ~n4538 & n4631;
  assign n4633 = n4538 & ~n4631;
  assign n4634 = ~n4632 & ~n4633;
  assign n4635 = ~n350 & ~n639;
  assign n4636 = ~n547 & n4635;
  assign n4637 = n1978 & n4636;
  assign n4638 = n1474 & n4637;
  assign n4639 = n810 & n4638;
  assign n4640 = ~n310 & n4639;
  assign n4641 = n2702 & n2947;
  assign n4642 = n1641 & n4641;
  assign n4643 = ~n330 & n4642;
  assign n4644 = n4640 & n4643;
  assign n4645 = n1109 & n4644;
  assign n4646 = ~n88 & ~n342;
  assign n4647 = ~n299 & n4646;
  assign n4648 = ~n594 & ~n668;
  assign n4649 = n4647 & n4648;
  assign n4650 = ~n681 & n4649;
  assign n4651 = ~n228 & ~n275;
  assign n4652 = ~n183 & n4651;
  assign n4653 = n4650 & n4652;
  assign n4654 = n1708 & n4653;
  assign n4655 = ~n400 & n4654;
  assign n4656 = ~n165 & n4655;
  assign n4657 = n1150 & n1478;
  assign n4658 = ~n252 & n4402;
  assign n4659 = ~n601 & n4658;
  assign n4660 = ~n123 & n476;
  assign n4661 = ~n155 & n4660;
  assign n4662 = n4659 & n4661;
  assign n4663 = n2345 & n4662;
  assign n4664 = n753 & n4663;
  assign n4665 = n456 & n4664;
  assign n4666 = n1516 & n4665;
  assign n4667 = ~n669 & n4666;
  assign n4668 = n4657 & n4667;
  assign n4669 = n3754 & n4668;
  assign n4670 = n4656 & n4669;
  assign n4671 = ~n692 & n2215;
  assign n4672 = ~n256 & n4671;
  assign n4673 = n923 & n4672;
  assign n4674 = ~n682 & n4673;
  assign n4675 = ~n689 & ~n705;
  assign n4676 = ~n466 & n4675;
  assign n4677 = n491 & n4676;
  assign n4678 = n1659 & n4677;
  assign n4679 = ~n180 & n4678;
  assign n4680 = ~n667 & n4679;
  assign n4681 = n4674 & n4680;
  assign n4682 = ~n442 & n1923;
  assign n4683 = n1964 & n4682;
  assign n4684 = n1830 & n4683;
  assign n4685 = n974 & n4684;
  assign n4686 = ~n290 & n4685;
  assign n4687 = ~n636 & ~n701;
  assign n4688 = ~n273 & ~n544;
  assign n4689 = n4687 & n4688;
  assign n4690 = ~n281 & n4689;
  assign n4691 = ~n298 & n3454;
  assign n4692 = ~n533 & n4691;
  assign n4693 = n4690 & n4692;
  assign n4694 = n1292 & n4693;
  assign n4695 = ~n589 & n4694;
  assign n4696 = ~n671 & n4695;
  assign n4697 = n4686 & n4696;
  assign n4698 = n4681 & n4697;
  assign n4699 = n4175 & n4698;
  assign n4700 = ~n441 & n4699;
  assign n4701 = n4670 & n4700;
  assign n4702 = n4645 & n4701;
  assign n4703 = n4439 & ~n4702;
  assign n4704 = ~n4439 & n4702;
  assign n4705 = ~n1740 & n3641;
  assign n4706 = ~n1610 & n3740;
  assign n4707 = n3593 & ~n3595;
  assign n4708 = ~n3596 & ~n4707;
  assign n4709 = n556 & n4708;
  assign n4710 = ~n1531 & n3961;
  assign n4711 = ~n4709 & ~n4710;
  assign n4712 = ~n4706 & n4711;
  assign n4713 = ~n4705 & n4712;
  assign n4714 = ~n4704 & ~n4713;
  assign n4715 = ~n4703 & ~n4714;
  assign n4716 = ~pi20  & ~n4526;
  assign n4717 = ~n4524 & n4527;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = ~n4715 & ~n4718;
  assign n4720 = n4715 & n4718;
  assign n4721 = ~n1610 & n3641;
  assign n4722 = ~n1531 & n3740;
  assign n4723 = n3597 & ~n3599;
  assign n4724 = ~n3600 & ~n4723;
  assign n4725 = n556 & n4724;
  assign n4726 = ~n1426 & n3961;
  assign n4727 = ~n4725 & ~n4726;
  assign n4728 = ~n4722 & n4727;
  assign n4729 = ~n4721 & n4728;
  assign n4730 = ~n4720 & ~n4729;
  assign n4731 = ~n4719 & ~n4730;
  assign n4732 = n4634 & ~n4731;
  assign n4733 = ~n4634 & n4731;
  assign n4734 = ~n4732 & ~n4733;
  assign n4735 = ~n1230 & n4006;
  assign n4736 = ~n1107 & n4133;
  assign n4737 = n4002 & n4307;
  assign n4738 = ~n1005 & n4555;
  assign n4739 = ~n4737 & ~n4738;
  assign n4740 = ~n4736 & n4739;
  assign n4741 = ~n4735 & n4740;
  assign n4742 = pi29  & n4741;
  assign n4743 = ~pi29  & ~n4741;
  assign n4744 = ~n4742 & ~n4743;
  assign n4745 = n4734 & ~n4744;
  assign n4746 = ~n4732 & ~n4745;
  assign n4747 = ~n4380 & ~n4381;
  assign n4748 = ~n4540 & n4747;
  assign n4749 = n4540 & ~n4747;
  assign n4750 = ~n4748 & ~n4749;
  assign n4751 = ~n1426 & n3641;
  assign n4752 = n3605 & ~n3607;
  assign n4753 = ~n3608 & ~n4752;
  assign n4754 = n556 & n4753;
  assign n4755 = ~n1230 & n3961;
  assign n4756 = ~n1338 & n3740;
  assign n4757 = ~n4755 & ~n4756;
  assign n4758 = ~n4754 & n4757;
  assign n4759 = ~n4751 & n4758;
  assign n4760 = ~n4750 & ~n4759;
  assign n4761 = n4750 & n4759;
  assign n4762 = ~n4760 & ~n4761;
  assign n4763 = ~n4746 & n4762;
  assign n4764 = ~n4760 & ~n4763;
  assign n4765 = ~n4332 & ~n4542;
  assign n4766 = ~n4543 & ~n4765;
  assign n4767 = n4764 & ~n4766;
  assign n4768 = ~n4764 & n4766;
  assign n4769 = ~n1005 & n4006;
  assign n4770 = ~n894 & n4133;
  assign n4771 = n4002 & n4122;
  assign n4772 = ~n795 & n4555;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = ~n4770 & n4773;
  assign n4775 = ~n4769 & n4774;
  assign n4776 = pi29  & n4775;
  assign n4777 = ~pi29  & ~n4775;
  assign n4778 = ~n4776 & ~n4777;
  assign n4779 = ~n4768 & n4778;
  assign n4780 = ~n4767 & ~n4779;
  assign n4781 = n4630 & n4780;
  assign n4782 = ~n3744 & n4602;
  assign n4783 = n4598 & n4599;
  assign n4784 = ~n554 & n4783;
  assign n4785 = ~n720 & n4601;
  assign n4786 = ~n4784 & ~n4785;
  assign n4787 = ~n4782 & n4786;
  assign n4788 = ~pi26  & ~n4787;
  assign n4789 = pi26  & n4787;
  assign n4790 = ~n4788 & ~n4789;
  assign n4791 = ~n4630 & ~n4780;
  assign n4792 = ~n4781 & ~n4791;
  assign n4793 = ~n4790 & n4792;
  assign n4794 = ~n4781 & ~n4793;
  assign n4795 = ~n4621 & ~n4623;
  assign n4796 = ~n4624 & ~n4795;
  assign n4797 = ~n4794 & n4796;
  assign n4798 = ~n665 & n4601;
  assign n4799 = ~n720 & n4783;
  assign n4800 = n3979 & n4602;
  assign n4801 = n4595 & ~n4598;
  assign n4802 = ~n554 & n4801;
  assign n4803 = ~n4800 & ~n4802;
  assign n4804 = ~n4799 & n4803;
  assign n4805 = ~n4798 & n4804;
  assign n4806 = pi26  & n4805;
  assign n4807 = ~pi26  & ~n4805;
  assign n4808 = ~n4806 & ~n4807;
  assign n4809 = ~n1107 & n4006;
  assign n4810 = ~n1005 & n4133;
  assign n4811 = n4002 & n4106;
  assign n4812 = ~n894 & n4555;
  assign n4813 = ~n4811 & ~n4812;
  assign n4814 = ~n4810 & n4813;
  assign n4815 = ~n4809 & n4814;
  assign n4816 = pi29  & n4815;
  assign n4817 = ~pi29  & ~n4815;
  assign n4818 = ~n4816 & ~n4817;
  assign n4819 = n4746 & ~n4762;
  assign n4820 = ~n4763 & ~n4819;
  assign n4821 = n4818 & ~n4820;
  assign n4822 = ~n4818 & n4820;
  assign n4823 = ~n795 & n4601;
  assign n4824 = ~n665 & n4783;
  assign n4825 = n4015 & n4602;
  assign n4826 = ~n720 & n4801;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = ~n4824 & n4827;
  assign n4829 = ~n4823 & n4828;
  assign n4830 = pi26  & n4829;
  assign n4831 = ~pi26  & ~n4829;
  assign n4832 = ~n4830 & ~n4831;
  assign n4833 = ~n4822 & n4832;
  assign n4834 = ~n4821 & ~n4833;
  assign n4835 = n4808 & n4834;
  assign n4836 = ~n4808 & ~n4834;
  assign n4837 = ~n4835 & ~n4836;
  assign n4838 = ~n4767 & ~n4768;
  assign n4839 = ~n4778 & n4838;
  assign n4840 = n4778 & ~n4838;
  assign n4841 = ~n4839 & ~n4840;
  assign n4842 = ~n4837 & n4841;
  assign n4843 = ~n4808 & n4834;
  assign n4844 = ~n4842 & ~n4843;
  assign n4845 = n4790 & ~n4792;
  assign n4846 = ~n4793 & ~n4845;
  assign n4847 = ~n4844 & n4846;
  assign n4848 = n4837 & ~n4841;
  assign n4849 = ~n4842 & ~n4848;
  assign n4850 = ~n1338 & n4006;
  assign n4851 = ~n1230 & n4133;
  assign n4852 = n4002 & n4323;
  assign n4853 = ~n1107 & n4555;
  assign n4854 = ~n4852 & ~n4853;
  assign n4855 = ~n4851 & n4854;
  assign n4856 = ~n4850 & n4855;
  assign n4857 = ~pi29  & ~n4856;
  assign n4858 = pi29  & n4856;
  assign n4859 = ~n4857 & ~n4858;
  assign n4860 = ~n4719 & ~n4720;
  assign n4861 = ~n4729 & n4860;
  assign n4862 = n4729 & ~n4860;
  assign n4863 = ~n4861 & ~n4862;
  assign n4864 = ~n4859 & n4863;
  assign n4865 = ~n4859 & ~n4863;
  assign n4866 = n4859 & n4863;
  assign n4867 = ~n4865 & ~n4866;
  assign n4868 = ~n4703 & ~n4704;
  assign n4869 = ~n4713 & n4868;
  assign n4870 = n4713 & ~n4868;
  assign n4871 = ~n4869 & ~n4870;
  assign n4872 = ~n375 & ~n705;
  assign n4873 = ~n197 & n4872;
  assign n4874 = ~n362 & n4873;
  assign n4875 = n1742 & n4874;
  assign n4876 = n3183 & n4875;
  assign n4877 = n2021 & n4876;
  assign n4878 = ~n129 & n4877;
  assign n4879 = n1305 & n2982;
  assign n4880 = n985 & n4879;
  assign n4881 = n1478 & n4880;
  assign n4882 = ~n394 & n4881;
  assign n4883 = n4878 & n4882;
  assign n4884 = n1120 & n2997;
  assign n4885 = n699 & n4884;
  assign n4886 = n1355 & n4885;
  assign n4887 = ~n548 & n4886;
  assign n4888 = ~n116 & ~n330;
  assign n4889 = n773 & n4888;
  assign n4890 = ~n323 & n4889;
  assign n4891 = n4887 & n4890;
  assign n4892 = n4883 & n4891;
  assign n4893 = ~n581 & n2616;
  assign n4894 = ~n160 & n4893;
  assign n4895 = n528 & n4894;
  assign n4896 = n2332 & n4895;
  assign n4897 = ~n344 & n967;
  assign n4898 = ~n117 & n4897;
  assign n4899 = n908 & n4898;
  assign n4900 = n1618 & n4899;
  assign n4901 = ~n299 & n4900;
  assign n4902 = ~n330 & n4901;
  assign n4903 = n2090 & n2491;
  assign n4904 = ~n436 & n4903;
  assign n4905 = ~n394 & n4904;
  assign n4906 = n4902 & n4905;
  assign n4907 = ~n155 & ~n163;
  assign n4908 = n1982 & n4907;
  assign n4909 = ~n166 & n4908;
  assign n4910 = ~n116 & ~n430;
  assign n4911 = ~n439 & n4910;
  assign n4912 = n4909 & n4911;
  assign n4913 = n997 & n4912;
  assign n4914 = ~n342 & n4913;
  assign n4915 = ~n289 & n4914;
  assign n4916 = ~n693 & n1924;
  assign n4917 = ~n81 & n4916;
  assign n4918 = n107 & n4917;
  assign n4919 = n857 & n4918;
  assign n4920 = ~n235 & n4919;
  assign n4921 = ~n626 & n4920;
  assign n4922 = n4915 & n4921;
  assign n4923 = n4906 & n4922;
  assign n4924 = n1353 & n4923;
  assign n4925 = ~n639 & n4924;
  assign n4926 = ~n236 & n4925;
  assign n4927 = n4896 & n4926;
  assign n4928 = n285 & n1217;
  assign n4929 = n1659 & n4928;
  assign n4930 = ~n705 & n4929;
  assign n4931 = ~n129 & n4930;
  assign n4932 = ~n229 & n4931;
  assign n4933 = ~n170 & n1395;
  assign n4934 = ~n112 & n4933;
  assign n4935 = n3045 & n4934;
  assign n4936 = n1892 & n4935;
  assign n4937 = n2214 & n4936;
  assign n4938 = ~n547 & n4937;
  assign n4939 = n4932 & n4938;
  assign n4940 = n4927 & n4939;
  assign n4941 = ~n4892 & ~n4940;
  assign n4942 = n4892 & n4940;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~pi17  & n4943;
  assign n4945 = ~n4941 & ~n4944;
  assign n4946 = n4439 & ~n4945;
  assign n4947 = ~n4439 & n4945;
  assign n4948 = ~n1811 & n3641;
  assign n4949 = ~n1740 & n3740;
  assign n4950 = n3589 & ~n3591;
  assign n4951 = ~n3592 & ~n4950;
  assign n4952 = n556 & n4951;
  assign n4953 = ~n1610 & n3961;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = ~n4949 & n4954;
  assign n4956 = ~n4948 & n4955;
  assign n4957 = ~n4947 & ~n4956;
  assign n4958 = ~n4946 & ~n4957;
  assign n4959 = n4871 & ~n4958;
  assign n4960 = ~n4871 & n4958;
  assign n4961 = ~n4959 & ~n4960;
  assign n4962 = ~pi17  & ~n4944;
  assign n4963 = ~n4942 & n4945;
  assign n4964 = ~n4962 & ~n4963;
  assign n4965 = ~n1900 & n3641;
  assign n4966 = n3585 & ~n3587;
  assign n4967 = ~n3588 & ~n4966;
  assign n4968 = n556 & n4967;
  assign n4969 = ~n1740 & n3961;
  assign n4970 = ~n1811 & n3740;
  assign n4971 = ~n4969 & ~n4970;
  assign n4972 = ~n4968 & n4971;
  assign n4973 = ~n4965 & n4972;
  assign n4974 = ~n4964 & ~n4973;
  assign n4975 = ~n629 & n3488;
  assign n4976 = ~n428 & n4975;
  assign n4977 = ~n401 & n4976;
  assign n4978 = ~n457 & ~n504;
  assign n4979 = n3195 & n4978;
  assign n4980 = ~n310 & n4979;
  assign n4981 = ~n599 & n4980;
  assign n4982 = n788 & n1656;
  assign n4983 = ~n506 & n4982;
  assign n4984 = ~n682 & n4983;
  assign n4985 = n4981 & n4984;
  assign n4986 = ~n626 & n2798;
  assign n4987 = ~n228 & n4986;
  assign n4988 = n549 & n1057;
  assign n4989 = ~n98 & n4988;
  assign n4990 = ~n150 & n4989;
  assign n4991 = n4987 & n4990;
  assign n4992 = n4985 & n4991;
  assign n4993 = n3806 & n4992;
  assign n4994 = ~n466 & n4993;
  assign n4995 = ~n229 & n4994;
  assign n4996 = n4977 & n4995;
  assign n4997 = n2940 & n3061;
  assign n4998 = n3202 & n4997;
  assign n4999 = n1466 & n4998;
  assign n5000 = n107 & n4999;
  assign n5001 = ~n262 & n5000;
  assign n5002 = ~n473 & n5001;
  assign n5003 = ~n219 & n3211;
  assign n5004 = n1813 & n5003;
  assign n5005 = ~n94 & n1285;
  assign n5006 = ~n464 & n5005;
  assign n5007 = n196 & n5006;
  assign n5008 = n5004 & n5007;
  assign n5009 = n3282 & n5008;
  assign n5010 = ~n304 & n5009;
  assign n5011 = ~n116 & n5010;
  assign n5012 = ~n132 & n5011;
  assign n5013 = n5002 & n5012;
  assign n5014 = n4996 & n5013;
  assign n5015 = n4892 & ~n5014;
  assign n5016 = ~n4892 & n5014;
  assign n5017 = ~n5015 & ~n5016;
  assign n5018 = ~n500 & n942;
  assign n5019 = ~n629 & n5018;
  assign n5020 = ~n236 & n4979;
  assign n5021 = ~n100 & n5020;
  assign n5022 = n5019 & n5021;
  assign n5023 = n199 & n4934;
  assign n5024 = ~n280 & n5023;
  assign n5025 = n1744 & n2979;
  assign n5026 = ~n621 & n5025;
  assign n5027 = n5024 & n5026;
  assign n5028 = ~n350 & n5027;
  assign n5029 = n3392 & n3897;
  assign n5030 = n5028 & n5029;
  assign n5031 = n1494 & n5030;
  assign n5032 = ~n332 & n5031;
  assign n5033 = ~n320 & n5032;
  assign n5034 = n2065 & n2281;
  assign n5035 = ~n477 & n5034;
  assign n5036 = ~n166 & n5035;
  assign n5037 = n5033 & n5036;
  assign n5038 = n5022 & n5037;
  assign n5039 = n902 & n5038;
  assign n5040 = n162 & n5039;
  assign n5041 = n1652 & n5040;
  assign n5042 = ~n462 & n5041;
  assign n5043 = ~n88 & ~n219;
  assign n5044 = ~n693 & n5043;
  assign n5045 = ~n685 & n2512;
  assign n5046 = ~n304 & n5045;
  assign n5047 = n5044 & n5046;
  assign n5048 = n431 & n5047;
  assign n5049 = n1401 & n5048;
  assign n5050 = ~n639 & n5049;
  assign n5051 = n5042 & n5050;
  assign n5052 = ~n305 & n1892;
  assign n5053 = ~n341 & n5052;
  assign n5054 = ~n692 & n5053;
  assign n5055 = ~n315 & n1939;
  assign n5056 = ~n413 & ~n631;
  assign n5057 = ~n697 & n5056;
  assign n5058 = ~n349 & n5057;
  assign n5059 = n5055 & n5058;
  assign n5060 = n3051 & n5059;
  assign n5061 = n5054 & n5060;
  assign n5062 = n2105 & n5061;
  assign n5063 = n725 & n5062;
  assign n5064 = ~n637 & n5063;
  assign n5065 = n230 & n3009;
  assign n5066 = ~n281 & n5065;
  assign n5067 = ~n278 & n5066;
  assign n5068 = n1131 & n1724;
  assign n5069 = ~n593 & n5068;
  assign n5070 = ~n704 & n5069;
  assign n5071 = ~n414 & n5070;
  assign n5072 = n5067 & n5071;
  assign n5073 = n392 & n673;
  assign n5074 = ~n297 & n5073;
  assign n5075 = ~n330 & n5074;
  assign n5076 = n1079 & n4662;
  assign n5077 = ~n679 & n5076;
  assign n5078 = ~n172 & n5077;
  assign n5079 = ~n214 & n5078;
  assign n5080 = n5075 & n5079;
  assign n5081 = n5072 & n5080;
  assign n5082 = n1864 & n5081;
  assign n5083 = ~n180 & n5082;
  assign n5084 = ~n583 & n5083;
  assign n5085 = n5064 & n5084;
  assign n5086 = n5051 & n5085;
  assign n5087 = ~n123 & ~n310;
  assign n5088 = n788 & n2921;
  assign n5089 = n5087 & n5088;
  assign n5090 = ~n144 & ~n544;
  assign n5091 = ~n198 & n5090;
  assign n5092 = n1168 & n3797;
  assign n5093 = n3284 & n5092;
  assign n5094 = ~n390 & n5093;
  assign n5095 = ~n259 & ~n385;
  assign n5096 = ~n98 & n5095;
  assign n5097 = ~n149 & n5096;
  assign n5098 = n1880 & n5097;
  assign n5099 = n89 & n5098;
  assign n5100 = ~n337 & n5099;
  assign n5101 = ~n626 & n5100;
  assign n5102 = n5094 & n5101;
  assign n5103 = ~n256 & n5102;
  assign n5104 = ~n115 & ~n314;
  assign n5105 = ~n214 & n5104;
  assign n5106 = ~n342 & n5105;
  assign n5107 = ~n595 & n5106;
  assign n5108 = ~n469 & n5107;
  assign n5109 = n5103 & n5108;
  assign n5110 = n5091 & n5109;
  assign n5111 = n5089 & n5110;
  assign n5112 = ~n393 & n5111;
  assign n5113 = ~n671 & n5112;
  assign n5114 = ~n439 & n5113;
  assign n5115 = ~n598 & ~n667;
  assign n5116 = ~n251 & n5115;
  assign n5117 = ~n298 & n5116;
  assign n5118 = n282 & ~n593;
  assign n5119 = n3045 & n5118;
  assign n5120 = ~n398 & n5119;
  assign n5121 = n5117 & n5120;
  assign n5122 = n4391 & n5121;
  assign n5123 = n997 & n5122;
  assign n5124 = ~n436 & n5123;
  assign n5125 = ~n208 & n1175;
  assign n5126 = ~n330 & n5125;
  assign n5127 = ~n527 & ~n678;
  assign n5128 = ~n324 & n5127;
  assign n5129 = ~n506 & n5128;
  assign n5130 = ~n533 & n5129;
  assign n5131 = n5126 & n5130;
  assign n5132 = ~n203 & ~n374;
  assign n5133 = ~n229 & n5132;
  assign n5134 = ~n273 & n2418;
  assign n5135 = ~n246 & n5134;
  assign n5136 = ~n360 & n5135;
  assign n5137 = n5133 & n5136;
  assign n5138 = n5131 & n5137;
  assign n5139 = ~n435 & ~n457;
  assign n5140 = ~n255 & ~n579;
  assign n5141 = ~n321 & n5140;
  assign n5142 = ~n357 & n5141;
  assign n5143 = n5139 & n5142;
  assign n5144 = n3479 & n5143;
  assign n5145 = n955 & n2685;
  assign n5146 = n5144 & n5145;
  assign n5147 = n5008 & n5146;
  assign n5148 = ~n155 & n5147;
  assign n5149 = ~n344 & n1355;
  assign n5150 = ~n361 & ~n588;
  assign n5151 = ~n279 & ~n502;
  assign n5152 = n5150 & n5151;
  assign n5153 = ~n218 & n5152;
  assign n5154 = n5149 & n5153;
  assign n5155 = n1659 & n5154;
  assign n5156 = ~n698 & n5155;
  assign n5157 = ~n332 & n5156;
  assign n5158 = n5148 & n5157;
  assign n5159 = ~n131 & n5158;
  assign n5160 = ~n345 & n2060;
  assign n5161 = ~n235 & n5160;
  assign n5162 = ~n187 & n5161;
  assign n5163 = n5159 & n5162;
  assign n5164 = n5138 & n5163;
  assign n5165 = ~n239 & n5164;
  assign n5166 = ~n277 & n5165;
  assign n5167 = n5124 & n5166;
  assign n5168 = n896 & n5167;
  assign n5169 = n5114 & n5168;
  assign n5170 = ~n5086 & ~n5169;
  assign n5171 = n5086 & n5169;
  assign n5172 = ~n5170 & ~n5171;
  assign n5173 = ~pi14  & n5172;
  assign n5174 = ~n5170 & ~n5173;
  assign n5175 = n5014 & ~n5174;
  assign n5176 = ~n5014 & n5174;
  assign n5177 = ~n2058 & n3641;
  assign n5178 = ~n2006 & n3740;
  assign n5179 = n3577 & ~n3579;
  assign n5180 = ~n3580 & ~n5179;
  assign n5181 = n556 & n5180;
  assign n5182 = ~n1900 & n3961;
  assign n5183 = ~n5181 & ~n5182;
  assign n5184 = ~n5178 & n5183;
  assign n5185 = ~n5177 & n5184;
  assign n5186 = ~n5176 & ~n5185;
  assign n5187 = ~n5175 & ~n5186;
  assign n5188 = n5017 & ~n5187;
  assign n5189 = ~n5015 & ~n5188;
  assign n5190 = n4964 & n4973;
  assign n5191 = ~n4974 & ~n5190;
  assign n5192 = ~n5189 & n5191;
  assign n5193 = ~n4974 & ~n5192;
  assign n5194 = ~n4946 & ~n4947;
  assign n5195 = ~n4956 & n5194;
  assign n5196 = n4956 & ~n5194;
  assign n5197 = ~n5195 & ~n5196;
  assign n5198 = ~n5193 & n5197;
  assign n5199 = n5193 & ~n5197;
  assign n5200 = ~n5198 & ~n5199;
  assign n5201 = ~n1531 & n4006;
  assign n5202 = ~n1426 & n4133;
  assign n5203 = n4002 & n4533;
  assign n5204 = ~n1338 & n4555;
  assign n5205 = ~n5203 & ~n5204;
  assign n5206 = ~n5202 & n5205;
  assign n5207 = ~n5201 & n5206;
  assign n5208 = pi29  & n5207;
  assign n5209 = ~pi29  & ~n5207;
  assign n5210 = ~n5208 & ~n5209;
  assign n5211 = n5200 & ~n5210;
  assign n5212 = ~n5198 & ~n5211;
  assign n5213 = n4961 & ~n5212;
  assign n5214 = ~n4959 & ~n5213;
  assign n5215 = ~n4867 & ~n5214;
  assign n5216 = ~n4864 & ~n5215;
  assign n5217 = ~n4734 & n4744;
  assign n5218 = ~n4745 & ~n5217;
  assign n5219 = ~n5216 & n5218;
  assign n5220 = ~n894 & n4601;
  assign n5221 = ~n795 & n4783;
  assign n5222 = n3959 & n4602;
  assign n5223 = ~n665 & n4801;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = ~n5221 & n5224;
  assign n5226 = ~n5220 & n5225;
  assign n5227 = ~pi26  & ~n5226;
  assign n5228 = pi26  & n5226;
  assign n5229 = ~n5227 & ~n5228;
  assign n5230 = n5216 & ~n5218;
  assign n5231 = ~n5219 & ~n5230;
  assign n5232 = ~n5229 & n5231;
  assign n5233 = ~n5219 & ~n5232;
  assign n5234 = ~pi22  & pi23 ;
  assign n5235 = pi22  & ~pi23 ;
  assign n5236 = ~n5234 & ~n5235;
  assign n5237 = n67 & n70;
  assign n5238 = ~n5236 & n5237;
  assign n5239 = ~n70 & ~n5236;
  assign n5240 = ~n3638 & n5239;
  assign n5241 = ~n5238 & ~n5240;
  assign n5242 = ~n554 & ~n5241;
  assign n5243 = pi23  & ~n5242;
  assign n5244 = ~pi23  & n5242;
  assign n5245 = ~n5243 & ~n5244;
  assign n5246 = n5233 & n5245;
  assign n5247 = ~n5233 & ~n5245;
  assign n5248 = ~n4821 & ~n4822;
  assign n5249 = ~n4832 & n5248;
  assign n5250 = n4832 & ~n5248;
  assign n5251 = ~n5249 & ~n5250;
  assign n5252 = ~n5247 & ~n5251;
  assign n5253 = ~n5246 & ~n5252;
  assign n5254 = n4849 & n5253;
  assign n5255 = n4867 & n5214;
  assign n5256 = ~n5215 & ~n5255;
  assign n5257 = ~n1005 & n4601;
  assign n5258 = ~n894 & n4783;
  assign n5259 = n4122 & n4602;
  assign n5260 = ~n795 & n4801;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = ~n5258 & n5261;
  assign n5263 = ~n5257 & n5262;
  assign n5264 = pi26  & n5263;
  assign n5265 = ~pi26  & ~n5263;
  assign n5266 = ~n5264 & ~n5265;
  assign n5267 = n5256 & ~n5266;
  assign n5268 = n5256 & n5266;
  assign n5269 = ~n5256 & ~n5266;
  assign n5270 = ~n5268 & ~n5269;
  assign n5271 = ~n4961 & n5212;
  assign n5272 = ~n5213 & ~n5271;
  assign n5273 = ~n1426 & n4006;
  assign n5274 = ~n1338 & n4133;
  assign n5275 = n4002 & n4753;
  assign n5276 = ~n1230 & n4555;
  assign n5277 = ~n5275 & ~n5276;
  assign n5278 = ~n5274 & n5277;
  assign n5279 = ~n5273 & n5278;
  assign n5280 = pi29  & n5279;
  assign n5281 = ~pi29  & ~n5279;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = n5272 & ~n5282;
  assign n5284 = ~n1107 & n4601;
  assign n5285 = ~n1005 & n4783;
  assign n5286 = n4106 & n4602;
  assign n5287 = ~n894 & n4801;
  assign n5288 = ~n5286 & ~n5287;
  assign n5289 = ~n5285 & n5288;
  assign n5290 = ~n5284 & n5289;
  assign n5291 = pi26  & n5290;
  assign n5292 = ~pi26  & ~n5290;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~n5272 & n5282;
  assign n5295 = ~n5293 & ~n5294;
  assign n5296 = ~n5283 & ~n5295;
  assign n5297 = ~n5270 & ~n5296;
  assign n5298 = ~n5267 & ~n5297;
  assign n5299 = n5229 & ~n5231;
  assign n5300 = ~n5232 & ~n5299;
  assign n5301 = ~n5298 & n5300;
  assign n5302 = ~n3744 & n5239;
  assign n5303 = n71 & ~n554;
  assign n5304 = ~n720 & n5238;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = ~n5302 & n5305;
  assign n5307 = ~pi23  & ~n5306;
  assign n5308 = pi23  & n5306;
  assign n5309 = ~n5307 & ~n5308;
  assign n5310 = n5298 & ~n5300;
  assign n5311 = ~n5301 & ~n5310;
  assign n5312 = ~n5309 & n5311;
  assign n5313 = ~n5301 & ~n5312;
  assign n5314 = ~n5246 & ~n5247;
  assign n5315 = n5251 & n5314;
  assign n5316 = ~n5251 & ~n5314;
  assign n5317 = ~n5315 & ~n5316;
  assign n5318 = ~n5313 & n5317;
  assign n5319 = n5313 & ~n5317;
  assign n5320 = ~n5318 & ~n5319;
  assign n5321 = n5309 & ~n5311;
  assign n5322 = ~n5312 & ~n5321;
  assign n5323 = ~n665 & n5238;
  assign n5324 = n71 & ~n720;
  assign n5325 = n3979 & n5239;
  assign n5326 = ~n70 & n5236;
  assign n5327 = ~n554 & n5326;
  assign n5328 = ~n5325 & ~n5327;
  assign n5329 = ~n5324 & n5328;
  assign n5330 = ~n5323 & n5329;
  assign n5331 = pi23  & n5330;
  assign n5332 = ~pi23  & ~n5330;
  assign n5333 = ~n5331 & ~n5332;
  assign n5334 = ~n5283 & ~n5294;
  assign n5335 = n5293 & ~n5334;
  assign n5336 = ~n5293 & n5334;
  assign n5337 = ~n5335 & ~n5336;
  assign n5338 = ~n5200 & n5210;
  assign n5339 = ~n5211 & ~n5338;
  assign n5340 = ~n5017 & n5187;
  assign n5341 = ~n5188 & ~n5340;
  assign n5342 = ~n2006 & n3641;
  assign n5343 = n3581 & ~n3583;
  assign n5344 = ~n3584 & ~n5343;
  assign n5345 = n556 & n5344;
  assign n5346 = ~n1811 & n3961;
  assign n5347 = ~n1900 & n3740;
  assign n5348 = ~n5346 & ~n5347;
  assign n5349 = ~n5345 & n5348;
  assign n5350 = ~n5342 & n5349;
  assign n5351 = n5341 & ~n5350;
  assign n5352 = ~n1740 & n4006;
  assign n5353 = ~n1610 & n4133;
  assign n5354 = n4002 & n4708;
  assign n5355 = ~n1531 & n4555;
  assign n5356 = ~n5354 & ~n5355;
  assign n5357 = ~n5353 & n5356;
  assign n5358 = ~n5352 & n5357;
  assign n5359 = ~pi29  & ~n5358;
  assign n5360 = pi29  & n5358;
  assign n5361 = ~n5359 & ~n5360;
  assign n5362 = n5341 & n5350;
  assign n5363 = ~n5341 & ~n5350;
  assign n5364 = ~n5362 & ~n5363;
  assign n5365 = ~n5361 & ~n5364;
  assign n5366 = ~n5351 & ~n5365;
  assign n5367 = n5189 & ~n5191;
  assign n5368 = ~n5192 & ~n5367;
  assign n5369 = ~n5366 & n5368;
  assign n5370 = ~n1610 & n4006;
  assign n5371 = ~n1531 & n4133;
  assign n5372 = n4002 & n4724;
  assign n5373 = ~n1426 & n4555;
  assign n5374 = ~n5372 & ~n5373;
  assign n5375 = ~n5371 & n5374;
  assign n5376 = ~n5370 & n5375;
  assign n5377 = pi29  & n5376;
  assign n5378 = ~pi29  & ~n5376;
  assign n5379 = ~n5377 & ~n5378;
  assign n5380 = n5366 & ~n5368;
  assign n5381 = ~n5379 & ~n5380;
  assign n5382 = ~n5369 & ~n5381;
  assign n5383 = n5339 & ~n5382;
  assign n5384 = ~n5339 & n5382;
  assign n5385 = ~n1230 & n4601;
  assign n5386 = ~n1107 & n4783;
  assign n5387 = n4307 & n4602;
  assign n5388 = ~n1005 & n4801;
  assign n5389 = ~n5387 & ~n5388;
  assign n5390 = ~n5386 & n5389;
  assign n5391 = ~n5385 & n5390;
  assign n5392 = pi26  & n5391;
  assign n5393 = ~pi26  & ~n5391;
  assign n5394 = ~n5392 & ~n5393;
  assign n5395 = ~n5384 & ~n5394;
  assign n5396 = ~n5383 & ~n5395;
  assign n5397 = n5337 & ~n5396;
  assign n5398 = ~n5337 & n5396;
  assign n5399 = ~n795 & n5238;
  assign n5400 = n71 & ~n665;
  assign n5401 = n4015 & n5239;
  assign n5402 = ~n720 & n5326;
  assign n5403 = ~n5401 & ~n5402;
  assign n5404 = ~n5400 & n5403;
  assign n5405 = ~n5399 & n5404;
  assign n5406 = pi23  & n5405;
  assign n5407 = ~pi23  & ~n5405;
  assign n5408 = ~n5406 & ~n5407;
  assign n5409 = ~n5398 & ~n5408;
  assign n5410 = ~n5397 & ~n5409;
  assign n5411 = ~n5333 & ~n5410;
  assign n5412 = n5333 & n5410;
  assign n5413 = n5270 & ~n5296;
  assign n5414 = ~n5270 & n5296;
  assign n5415 = ~n5413 & ~n5414;
  assign n5416 = ~n5412 & ~n5415;
  assign n5417 = ~n5411 & ~n5416;
  assign n5418 = n5322 & ~n5417;
  assign n5419 = ~n5411 & ~n5412;
  assign n5420 = ~n5415 & n5419;
  assign n5421 = n5415 & ~n5419;
  assign n5422 = ~n5420 & ~n5421;
  assign n5423 = pi17  & ~pi18 ;
  assign n5424 = ~pi17  & pi18 ;
  assign n5425 = ~n5423 & ~n5424;
  assign n5426 = pi19  & ~pi20 ;
  assign n5427 = ~pi19  & pi20 ;
  assign n5428 = ~n5426 & ~n5427;
  assign n5429 = ~n5425 & ~n5428;
  assign n5430 = ~n3638 & n5429;
  assign n5431 = ~pi18  & pi19 ;
  assign n5432 = pi18  & ~pi19 ;
  assign n5433 = ~n5431 & ~n5432;
  assign n5434 = n5425 & n5433;
  assign n5435 = ~n5428 & n5434;
  assign n5436 = ~n5430 & ~n5435;
  assign n5437 = ~n554 & ~n5436;
  assign n5438 = pi20  & ~n5437;
  assign n5439 = ~pi20  & n5437;
  assign n5440 = ~n5438 & ~n5439;
  assign n5441 = ~n1338 & n4601;
  assign n5442 = ~n1230 & n4783;
  assign n5443 = n4323 & n4602;
  assign n5444 = ~n1107 & n4801;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = ~n5442 & n5445;
  assign n5447 = ~n5441 & n5446;
  assign n5448 = pi26  & n5447;
  assign n5449 = ~pi26  & ~n5447;
  assign n5450 = ~n5448 & ~n5449;
  assign n5451 = ~n5369 & ~n5380;
  assign n5452 = n5379 & ~n5451;
  assign n5453 = ~n5379 & n5451;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = ~n5450 & n5454;
  assign n5456 = n5450 & ~n5454;
  assign n5457 = ~n5455 & ~n5456;
  assign n5458 = ~n5175 & ~n5176;
  assign n5459 = ~n5185 & n5458;
  assign n5460 = n5185 & ~n5458;
  assign n5461 = ~n5459 & ~n5460;
  assign n5462 = n1032 & n2738;
  assign n5463 = n3187 & n5462;
  assign n5464 = ~n477 & n5463;
  assign n5465 = n1283 & n4090;
  assign n5466 = ~n590 & n5465;
  assign n5467 = ~n579 & n3912;
  assign n5468 = ~n117 & n5467;
  assign n5469 = ~n533 & n5468;
  assign n5470 = n5466 & n5469;
  assign n5471 = n1767 & n3820;
  assign n5472 = ~n588 & n5471;
  assign n5473 = ~n545 & n5472;
  assign n5474 = ~n123 & n3897;
  assign n5475 = n437 & n5474;
  assign n5476 = n1402 & n5475;
  assign n5477 = n1494 & n5476;
  assign n5478 = n1368 & n5477;
  assign n5479 = ~n681 & n5478;
  assign n5480 = ~n638 & n5479;
  assign n5481 = n5473 & n5480;
  assign n5482 = n5470 & n5481;
  assign n5483 = ~n466 & ~n589;
  assign n5484 = ~n614 & n5483;
  assign n5485 = ~n273 & n5484;
  assign n5486 = ~n666 & n4354;
  assign n5487 = ~n170 & n5486;
  assign n5488 = n5485 & n5487;
  assign n5489 = n5482 & n5488;
  assign n5490 = ~n324 & n5489;
  assign n5491 = ~n422 & n5490;
  assign n5492 = n5464 & n5491;
  assign n5493 = ~n354 & ~n504;
  assign n5494 = n148 & ~n548;
  assign n5495 = n488 & n1783;
  assign n5496 = ~n94 & n306;
  assign n5497 = n1362 & n5496;
  assign n5498 = n930 & n5497;
  assign n5499 = n967 & n5498;
  assign n5500 = n2585 & n5499;
  assign n5501 = n5495 & n5500;
  assign n5502 = ~n399 & n5501;
  assign n5503 = n1380 & n4175;
  assign n5504 = ~n112 & n5503;
  assign n5505 = ~n390 & ~n473;
  assign n5506 = n1180 & n5505;
  assign n5507 = n4888 & n5506;
  assign n5508 = ~n280 & n5507;
  assign n5509 = n5504 & n5508;
  assign n5510 = n5502 & n5509;
  assign n5511 = n5494 & n5510;
  assign n5512 = n5493 & n5511;
  assign n5513 = n1138 & n5512;
  assign n5514 = ~n193 & n5513;
  assign n5515 = ~n278 & n5514;
  assign n5516 = ~n518 & n3309;
  assign n5517 = ~n197 & n5516;
  assign n5518 = n1109 & n5517;
  assign n5519 = n135 & ~n353;
  assign n5520 = ~n165 & n3499;
  assign n5521 = n5519 & n5520;
  assign n5522 = ~n239 & ~n325;
  assign n5523 = ~n235 & ~n475;
  assign n5524 = ~n595 & n5523;
  assign n5525 = n5522 & n5524;
  assign n5526 = n5521 & n5525;
  assign n5527 = n5518 & n5526;
  assign n5528 = n1516 & n5527;
  assign n5529 = ~n186 & n5528;
  assign n5530 = ~n114 & n5529;
  assign n5531 = n5515 & n5530;
  assign n5532 = n5492 & n5531;
  assign n5533 = n5169 & ~n5532;
  assign n5534 = ~n5169 & n5532;
  assign n5535 = ~n2278 & n3641;
  assign n5536 = ~n2178 & n3740;
  assign n5537 = n3569 & ~n3571;
  assign n5538 = ~n3572 & ~n5537;
  assign n5539 = n556 & n5538;
  assign n5540 = ~n2058 & n3961;
  assign n5541 = ~n5539 & ~n5540;
  assign n5542 = ~n5536 & n5541;
  assign n5543 = ~n5535 & n5542;
  assign n5544 = ~n5534 & ~n5543;
  assign n5545 = ~n5533 & ~n5544;
  assign n5546 = ~pi14  & ~n5173;
  assign n5547 = ~n5171 & n5174;
  assign n5548 = ~n5546 & ~n5547;
  assign n5549 = ~n5545 & ~n5548;
  assign n5550 = n5545 & n5548;
  assign n5551 = ~n2178 & n3641;
  assign n5552 = ~n2058 & n3740;
  assign n5553 = n3573 & ~n3575;
  assign n5554 = ~n3576 & ~n5553;
  assign n5555 = n556 & n5554;
  assign n5556 = ~n2006 & n3961;
  assign n5557 = ~n5555 & ~n5556;
  assign n5558 = ~n5552 & n5557;
  assign n5559 = ~n5551 & n5558;
  assign n5560 = ~n5550 & ~n5559;
  assign n5561 = ~n5549 & ~n5560;
  assign n5562 = n5461 & ~n5561;
  assign n5563 = ~n5461 & n5561;
  assign n5564 = ~n5562 & ~n5563;
  assign n5565 = ~n1811 & n4006;
  assign n5566 = ~n1740 & n4133;
  assign n5567 = n4002 & n4951;
  assign n5568 = ~n1610 & n4555;
  assign n5569 = ~n5567 & ~n5568;
  assign n5570 = ~n5566 & n5569;
  assign n5571 = ~n5565 & n5570;
  assign n5572 = pi29  & n5571;
  assign n5573 = ~pi29  & ~n5571;
  assign n5574 = ~n5572 & ~n5573;
  assign n5575 = n5564 & ~n5574;
  assign n5576 = ~n5562 & ~n5575;
  assign n5577 = n5361 & n5364;
  assign n5578 = ~n5365 & ~n5577;
  assign n5579 = ~n5576 & n5578;
  assign n5580 = n5576 & ~n5578;
  assign n5581 = ~n1426 & n4601;
  assign n5582 = ~n1338 & n4783;
  assign n5583 = n4602 & n4753;
  assign n5584 = ~n1230 & n4801;
  assign n5585 = ~n5583 & ~n5584;
  assign n5586 = ~n5582 & n5585;
  assign n5587 = ~n5581 & n5586;
  assign n5588 = pi26  & n5587;
  assign n5589 = ~pi26  & ~n5587;
  assign n5590 = ~n5588 & ~n5589;
  assign n5591 = ~n5580 & ~n5590;
  assign n5592 = ~n5579 & ~n5591;
  assign n5593 = n5457 & ~n5592;
  assign n5594 = ~n5455 & ~n5593;
  assign n5595 = ~n5383 & ~n5384;
  assign n5596 = ~n5394 & n5595;
  assign n5597 = n5394 & ~n5595;
  assign n5598 = ~n5596 & ~n5597;
  assign n5599 = ~n5594 & n5598;
  assign n5600 = n5594 & ~n5598;
  assign n5601 = ~n894 & n5238;
  assign n5602 = n71 & ~n795;
  assign n5603 = n3959 & n5239;
  assign n5604 = ~n665 & n5326;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = ~n5602 & n5605;
  assign n5607 = ~n5601 & n5606;
  assign n5608 = pi23  & n5607;
  assign n5609 = ~pi23  & ~n5607;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = ~n5600 & ~n5610;
  assign n5612 = ~n5599 & ~n5611;
  assign n5613 = ~n5440 & ~n5612;
  assign n5614 = n5440 & n5612;
  assign n5615 = ~n5397 & ~n5398;
  assign n5616 = ~n5408 & n5615;
  assign n5617 = n5408 & ~n5615;
  assign n5618 = ~n5616 & ~n5617;
  assign n5619 = ~n5614 & n5618;
  assign n5620 = ~n5613 & ~n5619;
  assign n5621 = n5422 & ~n5620;
  assign n5622 = ~n5422 & n5620;
  assign n5623 = ~n5621 & ~n5622;
  assign n5624 = ~n5613 & ~n5614;
  assign n5625 = n5618 & n5624;
  assign n5626 = ~n5618 & ~n5624;
  assign n5627 = ~n5625 & ~n5626;
  assign n5628 = ~n1005 & n5238;
  assign n5629 = n71 & ~n894;
  assign n5630 = n4122 & n5239;
  assign n5631 = ~n795 & n5326;
  assign n5632 = ~n5630 & ~n5631;
  assign n5633 = ~n5629 & n5632;
  assign n5634 = ~n5628 & n5633;
  assign n5635 = ~pi23  & ~n5634;
  assign n5636 = pi23  & n5634;
  assign n5637 = ~n5635 & ~n5636;
  assign n5638 = ~n5457 & n5592;
  assign n5639 = ~n5593 & ~n5638;
  assign n5640 = ~n5637 & n5639;
  assign n5641 = ~n5637 & ~n5639;
  assign n5642 = n5637 & n5639;
  assign n5643 = ~n5641 & ~n5642;
  assign n5644 = ~n5579 & ~n5580;
  assign n5645 = ~n5590 & n5644;
  assign n5646 = n5590 & ~n5644;
  assign n5647 = ~n5645 & ~n5646;
  assign n5648 = ~n1900 & n4006;
  assign n5649 = ~n1811 & n4133;
  assign n5650 = n4002 & n4967;
  assign n5651 = ~n1740 & n4555;
  assign n5652 = ~n5650 & ~n5651;
  assign n5653 = ~n5649 & n5652;
  assign n5654 = ~n5648 & n5653;
  assign n5655 = ~pi29  & ~n5654;
  assign n5656 = pi29  & n5654;
  assign n5657 = ~n5655 & ~n5656;
  assign n5658 = ~n5549 & ~n5550;
  assign n5659 = ~n5559 & n5658;
  assign n5660 = n5559 & ~n5658;
  assign n5661 = ~n5659 & ~n5660;
  assign n5662 = ~n5657 & n5661;
  assign n5663 = ~n5657 & ~n5661;
  assign n5664 = n5657 & n5661;
  assign n5665 = ~n5663 & ~n5664;
  assign n5666 = ~n5533 & ~n5534;
  assign n5667 = ~n5543 & n5666;
  assign n5668 = n5543 & ~n5666;
  assign n5669 = ~n5667 & ~n5668;
  assign n5670 = n3138 & n3265;
  assign n5671 = ~n262 & ~n293;
  assign n5672 = ~n474 & n5671;
  assign n5673 = n5670 & n5672;
  assign n5674 = ~n279 & n5673;
  assign n5675 = ~n273 & n2557;
  assign n5676 = ~n669 & n5675;
  assign n5677 = ~n441 & ~n534;
  assign n5678 = ~n628 & n5677;
  assign n5679 = ~n247 & n5678;
  assign n5680 = ~n458 & n2529;
  assign n5681 = ~n374 & n5680;
  assign n5682 = n5679 & n5681;
  assign n5683 = ~n678 & n5682;
  assign n5684 = ~n344 & n5683;
  assign n5685 = n5676 & n5684;
  assign n5686 = ~n104 & ~n255;
  assign n5687 = ~n395 & n5686;
  assign n5688 = n1622 & n5687;
  assign n5689 = ~n353 & n5688;
  assign n5690 = ~n115 & n5689;
  assign n5691 = n2136 & n4260;
  assign n5692 = ~n436 & n5691;
  assign n5693 = ~n580 & n5692;
  assign n5694 = n5690 & n5693;
  assign n5695 = n5685 & n5694;
  assign n5696 = n3695 & n5695;
  assign n5697 = ~n693 & n5696;
  assign n5698 = n5674 & n5697;
  assign n5699 = n2432 & n5121;
  assign n5700 = n1258 & n5699;
  assign n5701 = ~n236 & n5700;
  assign n5702 = n322 & n5056;
  assign n5703 = ~n231 & n5702;
  assign n5704 = ~n170 & ~n294;
  assign n5705 = n998 & n5704;
  assign n5706 = ~n112 & n5705;
  assign n5707 = ~n457 & n5706;
  assign n5708 = n5703 & n5707;
  assign n5709 = ~n194 & n5708;
  assign n5710 = n765 & n5160;
  assign n5711 = n3248 & n5710;
  assign n5712 = n5709 & n5711;
  assign n5713 = ~n314 & ~n636;
  assign n5714 = ~n324 & n5713;
  assign n5715 = n1618 & n5714;
  assign n5716 = n5712 & n5715;
  assign n5717 = ~n289 & n5716;
  assign n5718 = n5701 & n5717;
  assign n5719 = n5698 & n5718;
  assign n5720 = n4187 & n5712;
  assign n5721 = ~n330 & n5720;
  assign n5722 = ~n670 & n5721;
  assign n5723 = n1720 & n3704;
  assign n5724 = n167 & n5723;
  assign n5725 = n1132 & n5724;
  assign n5726 = ~n198 & n5725;
  assign n5727 = ~n288 & n5726;
  assign n5728 = n5722 & n5727;
  assign n5729 = ~n698 & n901;
  assign n5730 = ~n548 & n5729;
  assign n5731 = ~n435 & n5730;
  assign n5732 = n1554 & n2494;
  assign n5733 = ~n614 & n5732;
  assign n5734 = ~n441 & n5733;
  assign n5735 = ~n117 & n1577;
  assign n5736 = ~n152 & n5735;
  assign n5737 = n1784 & n3305;
  assign n5738 = ~n324 & ~n693;
  assign n5739 = ~n578 & n5738;
  assign n5740 = ~n593 & n5739;
  assign n5741 = ~n357 & n5740;
  assign n5742 = n5737 & n5741;
  assign n5743 = n4354 & n5742;
  assign n5744 = n5736 & n5743;
  assign n5745 = n706 & n5744;
  assign n5746 = ~n583 & n5745;
  assign n5747 = ~n280 & n5746;
  assign n5748 = n5734 & n5747;
  assign n5749 = n2505 & n3715;
  assign n5750 = ~n594 & n5749;
  assign n5751 = ~n690 & n5750;
  assign n5752 = ~n344 & ~n601;
  assign n5753 = ~n612 & n5752;
  assign n5754 = n2088 & n5753;
  assign n5755 = n1892 & n5754;
  assign n5756 = ~n163 & n5755;
  assign n5757 = ~n160 & n5756;
  assign n5758 = n5751 & n5757;
  assign n5759 = n5748 & n5758;
  assign n5760 = n1918 & n5759;
  assign n5761 = n1622 & n4408;
  assign n5762 = n1830 & n5761;
  assign n5763 = n1268 & n5762;
  assign n5764 = n5760 & n5763;
  assign n5765 = ~n155 & n5764;
  assign n5766 = ~n213 & n5765;
  assign n5767 = n5731 & n5766;
  assign n5768 = n5728 & n5767;
  assign n5769 = ~n5719 & ~n5768;
  assign n5770 = n5719 & n5768;
  assign n5771 = ~n5769 & ~n5770;
  assign n5772 = ~pi11  & n5771;
  assign n5773 = ~n5769 & ~n5772;
  assign n5774 = n5169 & ~n5773;
  assign n5775 = ~n5169 & n5773;
  assign n5776 = ~n2369 & n3641;
  assign n5777 = ~n2278 & n3740;
  assign n5778 = n3565 & ~n3567;
  assign n5779 = ~n3568 & ~n5778;
  assign n5780 = n556 & n5779;
  assign n5781 = ~n2178 & n3961;
  assign n5782 = ~n5780 & ~n5781;
  assign n5783 = ~n5777 & n5782;
  assign n5784 = ~n5776 & n5783;
  assign n5785 = ~n5775 & ~n5784;
  assign n5786 = ~n5774 & ~n5785;
  assign n5787 = n5669 & ~n5786;
  assign n5788 = ~n5669 & n5786;
  assign n5789 = ~n5787 & ~n5788;
  assign n5790 = ~pi11  & ~n5772;
  assign n5791 = ~n5770 & n5773;
  assign n5792 = ~n5790 & ~n5791;
  assign n5793 = ~n2457 & n3641;
  assign n5794 = n3561 & ~n3563;
  assign n5795 = ~n3564 & ~n5794;
  assign n5796 = n556 & n5795;
  assign n5797 = ~n2278 & n3961;
  assign n5798 = ~n2369 & n3740;
  assign n5799 = ~n5797 & ~n5798;
  assign n5800 = ~n5796 & n5799;
  assign n5801 = ~n5793 & n5800;
  assign n5802 = ~n5792 & ~n5801;
  assign n5803 = ~n581 & n1079;
  assign n5804 = ~n399 & n5803;
  assign n5805 = n1716 & n5804;
  assign n5806 = ~n458 & n5805;
  assign n5807 = n1751 & n4208;
  assign n5808 = ~n353 & n5807;
  assign n5809 = ~n309 & n5808;
  assign n5810 = n5806 & n5809;
  assign n5811 = ~n218 & n2345;
  assign n5812 = ~n668 & n5811;
  assign n5813 = n2396 & n5812;
  assign n5814 = n2683 & n5813;
  assign n5815 = ~n104 & n5814;
  assign n5816 = ~n413 & n5815;
  assign n5817 = ~n390 & n2021;
  assign n5818 = ~n423 & ~n599;
  assign n5819 = ~n297 & n5818;
  assign n5820 = n5817 & n5819;
  assign n5821 = n2451 & n5820;
  assign n5822 = n3215 & n5821;
  assign n5823 = ~n325 & n5822;
  assign n5824 = ~n627 & n5823;
  assign n5825 = n5816 & n5824;
  assign n5826 = n5810 & n5825;
  assign n5827 = n5719 & ~n5826;
  assign n5828 = ~n5719 & n5826;
  assign n5829 = ~n5827 & ~n5828;
  assign n5830 = ~n373 & n1817;
  assign n5831 = ~n461 & n5830;
  assign n5832 = ~n413 & ~n473;
  assign n5833 = ~n172 & n5832;
  assign n5834 = ~n229 & n2939;
  assign n5835 = ~n195 & n5834;
  assign n5836 = ~n384 & n5835;
  assign n5837 = n5833 & n5836;
  assign n5838 = n1936 & n5837;
  assign n5839 = ~n171 & n5838;
  assign n5840 = ~n147 & n5839;
  assign n5841 = n5831 & n5840;
  assign n5842 = ~n85 & ~n422;
  assign n5843 = ~n106 & ~n637;
  assign n5844 = n5842 & n5843;
  assign n5845 = ~n547 & n5844;
  assign n5846 = ~n578 & n4243;
  assign n5847 = ~n588 & n5846;
  assign n5848 = ~n349 & n5847;
  assign n5849 = n5845 & n5848;
  assign n5850 = n1124 & n5849;
  assign n5851 = ~n517 & n5850;
  assign n5852 = ~n683 & n5851;
  assign n5853 = n333 & n5128;
  assign n5854 = ~n610 & n5853;
  assign n5855 = ~n188 & n5854;
  assign n5856 = ~n394 & n5855;
  assign n5857 = n5852 & n5856;
  assign n5858 = n5841 & n5857;
  assign n5859 = n268 & n5858;
  assign n5860 = ~n590 & n5859;
  assign n5861 = ~n424 & n5860;
  assign n5862 = n1565 & n1785;
  assign n5863 = ~n308 & n5862;
  assign n5864 = ~n391 & n5863;
  assign n5865 = ~n122 & n1923;
  assign n5866 = ~n666 & n5865;
  assign n5867 = n706 & n5866;
  assign n5868 = ~n235 & n5867;
  assign n5869 = ~n228 & n5868;
  assign n5870 = n5864 & n5869;
  assign n5871 = n1464 & n5047;
  assign n5872 = ~n334 & n5871;
  assign n5873 = ~n360 & n5872;
  assign n5874 = n2931 & n4260;
  assign n5875 = ~n166 & n5874;
  assign n5876 = ~n181 & n5875;
  assign n5877 = n5873 & n5876;
  assign n5878 = n5870 & n5877;
  assign n5879 = n5753 & n5878;
  assign n5880 = ~n466 & n5879;
  assign n5881 = ~n670 & n5880;
  assign n5882 = n5861 & n5881;
  assign n5883 = ~n289 & ~n700;
  assign n5884 = ~n275 & ~n441;
  assign n5885 = n295 & n5884;
  assign n5886 = ~n697 & n5885;
  assign n5887 = ~n342 & n2481;
  assign n5888 = ~n692 & n5887;
  assign n5889 = n5886 & n5888;
  assign n5890 = n1583 & n5889;
  assign n5891 = n5883 & n5890;
  assign n5892 = ~n314 & n5891;
  assign n5893 = ~n217 & ~n280;
  assign n5894 = ~n548 & n5893;
  assign n5895 = ~n197 & n3117;
  assign n5896 = ~n129 & n5895;
  assign n5897 = n5894 & n5896;
  assign n5898 = n2576 & n5897;
  assign n5899 = ~n236 & n5898;
  assign n5900 = ~n213 & n5899;
  assign n5901 = n5892 & n5900;
  assign n5902 = n5882 & n5901;
  assign n5903 = ~n429 & n797;
  assign n5904 = ~n100 & ~n372;
  assign n5905 = n1272 & n5904;
  assign n5906 = ~n671 & n5905;
  assign n5907 = n5903 & n5906;
  assign n5908 = n920 & n5907;
  assign n5909 = ~n679 & n1181;
  assign n5910 = ~n628 & n5909;
  assign n5911 = ~n354 & n3113;
  assign n5912 = ~n394 & n5911;
  assign n5913 = n5910 & n5912;
  assign n5914 = ~n94 & n5913;
  assign n5915 = ~n599 & ~n704;
  assign n5916 = ~n545 & n5915;
  assign n5917 = n881 & n5916;
  assign n5918 = n5914 & n5917;
  assign n5919 = n515 & n5918;
  assign n5920 = n5908 & n5919;
  assign n5921 = n4683 & n5920;
  assign n5922 = ~n395 & n5921;
  assign n5923 = ~n218 & n237;
  assign n5924 = ~n293 & n5923;
  assign n5925 = n1124 & n5924;
  assign n5926 = n2409 & n5925;
  assign n5927 = n810 & n5926;
  assign n5928 = ~n631 & n5927;
  assign n5929 = ~n506 & n5928;
  assign n5930 = n5922 & n5929;
  assign n5931 = ~n149 & n5930;
  assign n5932 = ~n695 & n1577;
  assign n5933 = ~n150 & n5932;
  assign n5934 = n5931 & n5933;
  assign n5935 = n291 & ~n698;
  assign n5936 = ~n112 & ~n468;
  assign n5937 = n5935 & n5936;
  assign n5938 = ~n214 & n5937;
  assign n5939 = ~n260 & ~n273;
  assign n5940 = ~n278 & n5939;
  assign n5941 = ~n390 & n5940;
  assign n5942 = n5938 & n5941;
  assign n5943 = n5934 & n5942;
  assign n5944 = ~n583 & n5943;
  assign n5945 = n562 & n3352;
  assign n5946 = n946 & n5945;
  assign n5947 = ~n500 & n5946;
  assign n5948 = ~n670 & n5947;
  assign n5949 = n5944 & n5948;
  assign n5950 = ~n297 & n1908;
  assign n5951 = ~n122 & n5950;
  assign n5952 = ~n163 & n2428;
  assign n5953 = ~n626 & n5952;
  assign n5954 = n5951 & n5953;
  assign n5955 = ~n393 & n5954;
  assign n5956 = ~n345 & n816;
  assign n5957 = ~n204 & n5956;
  assign n5958 = n415 & n5957;
  assign n5959 = n5955 & n5958;
  assign n5960 = n694 & n5959;
  assign n5961 = n1340 & n5960;
  assign n5962 = ~n104 & n5961;
  assign n5963 = n4670 & n4677;
  assign n5964 = n1131 & n5963;
  assign n5965 = ~n544 & n5964;
  assign n5966 = ~n344 & n5965;
  assign n5967 = n5962 & n5966;
  assign n5968 = n5949 & n5967;
  assign n5969 = ~n5902 & ~n5968;
  assign n5970 = n5902 & n5968;
  assign n5971 = ~n5969 & ~n5970;
  assign n5972 = ~pi8  & n5971;
  assign n5973 = ~n5969 & ~n5972;
  assign n5974 = n5719 & ~n5973;
  assign n5975 = ~n5719 & n5973;
  assign n5976 = ~n2640 & n3641;
  assign n5977 = ~n2554 & n3740;
  assign n5978 = n3553 & ~n3555;
  assign n5979 = ~n3556 & ~n5978;
  assign n5980 = n556 & n5979;
  assign n5981 = ~n2457 & n3961;
  assign n5982 = ~n5980 & ~n5981;
  assign n5983 = ~n5977 & n5982;
  assign n5984 = ~n5976 & n5983;
  assign n5985 = ~n5975 & ~n5984;
  assign n5986 = ~n5974 & ~n5985;
  assign n5987 = n5829 & ~n5986;
  assign n5988 = ~n5827 & ~n5987;
  assign n5989 = n5792 & n5801;
  assign n5990 = ~n5802 & ~n5989;
  assign n5991 = ~n5988 & n5990;
  assign n5992 = ~n5802 & ~n5991;
  assign n5993 = ~n5774 & ~n5775;
  assign n5994 = ~n5784 & n5993;
  assign n5995 = n5784 & ~n5993;
  assign n5996 = ~n5994 & ~n5995;
  assign n5997 = ~n5992 & n5996;
  assign n5998 = n5992 & ~n5996;
  assign n5999 = ~n5997 & ~n5998;
  assign n6000 = ~n2058 & n4006;
  assign n6001 = ~n2006 & n4133;
  assign n6002 = n4002 & n5180;
  assign n6003 = ~n1900 & n4555;
  assign n6004 = ~n6002 & ~n6003;
  assign n6005 = ~n6001 & n6004;
  assign n6006 = ~n6000 & n6005;
  assign n6007 = pi29  & n6006;
  assign n6008 = ~pi29  & ~n6006;
  assign n6009 = ~n6007 & ~n6008;
  assign n6010 = n5999 & ~n6009;
  assign n6011 = ~n5997 & ~n6010;
  assign n6012 = n5789 & ~n6011;
  assign n6013 = ~n5787 & ~n6012;
  assign n6014 = ~n5665 & ~n6013;
  assign n6015 = ~n5662 & ~n6014;
  assign n6016 = ~n5564 & n5574;
  assign n6017 = ~n5575 & ~n6016;
  assign n6018 = ~n6015 & n6017;
  assign n6019 = n6015 & ~n6017;
  assign n6020 = ~n1531 & n4601;
  assign n6021 = ~n1426 & n4783;
  assign n6022 = n4533 & n4602;
  assign n6023 = ~n1338 & n4801;
  assign n6024 = ~n6022 & ~n6023;
  assign n6025 = ~n6021 & n6024;
  assign n6026 = ~n6020 & n6025;
  assign n6027 = pi26  & n6026;
  assign n6028 = ~pi26  & ~n6026;
  assign n6029 = ~n6027 & ~n6028;
  assign n6030 = ~n6019 & ~n6029;
  assign n6031 = ~n6018 & ~n6030;
  assign n6032 = n5647 & ~n6031;
  assign n6033 = ~n5647 & n6031;
  assign n6034 = ~n1107 & n5238;
  assign n6035 = n71 & ~n1005;
  assign n6036 = n4106 & n5239;
  assign n6037 = ~n894 & n5326;
  assign n6038 = ~n6036 & ~n6037;
  assign n6039 = ~n6035 & n6038;
  assign n6040 = ~n6034 & n6039;
  assign n6041 = pi23  & n6040;
  assign n6042 = ~pi23  & ~n6040;
  assign n6043 = ~n6041 & ~n6042;
  assign n6044 = ~n6033 & ~n6043;
  assign n6045 = ~n6032 & ~n6044;
  assign n6046 = ~n5643 & ~n6045;
  assign n6047 = ~n5640 & ~n6046;
  assign n6048 = ~n5599 & ~n5600;
  assign n6049 = ~n5610 & n6048;
  assign n6050 = n5610 & ~n6048;
  assign n6051 = ~n6049 & ~n6050;
  assign n6052 = ~n6047 & n6051;
  assign n6053 = n6047 & ~n6051;
  assign n6054 = ~n3744 & n5429;
  assign n6055 = n5425 & ~n5433;
  assign n6056 = ~n554 & n6055;
  assign n6057 = ~n720 & n5435;
  assign n6058 = ~n6056 & ~n6057;
  assign n6059 = ~n6054 & n6058;
  assign n6060 = pi20  & n6059;
  assign n6061 = ~pi20  & ~n6059;
  assign n6062 = ~n6060 & ~n6061;
  assign n6063 = ~n6053 & ~n6062;
  assign n6064 = ~n6052 & ~n6063;
  assign n6065 = n5627 & ~n6064;
  assign n6066 = ~n5627 & n6064;
  assign n6067 = ~n6065 & ~n6066;
  assign n6068 = ~n665 & n5435;
  assign n6069 = ~n720 & n6055;
  assign n6070 = n3979 & n5429;
  assign n6071 = ~n5425 & n5428;
  assign n6072 = ~n554 & n6071;
  assign n6073 = ~n6070 & ~n6072;
  assign n6074 = ~n6069 & n6073;
  assign n6075 = ~n6068 & n6074;
  assign n6076 = pi20  & n6075;
  assign n6077 = ~pi20  & ~n6075;
  assign n6078 = ~n6076 & ~n6077;
  assign n6079 = ~n6032 & ~n6033;
  assign n6080 = ~n6043 & n6079;
  assign n6081 = n6043 & ~n6079;
  assign n6082 = ~n6080 & ~n6081;
  assign n6083 = n5665 & n6013;
  assign n6084 = ~n6014 & ~n6083;
  assign n6085 = ~n1610 & n4601;
  assign n6086 = ~n1531 & n4783;
  assign n6087 = n4602 & n4724;
  assign n6088 = ~n1426 & n4801;
  assign n6089 = ~n6087 & ~n6088;
  assign n6090 = ~n6086 & n6089;
  assign n6091 = ~n6085 & n6090;
  assign n6092 = pi26  & n6091;
  assign n6093 = ~pi26  & ~n6091;
  assign n6094 = ~n6092 & ~n6093;
  assign n6095 = n6084 & ~n6094;
  assign n6096 = ~n6084 & n6094;
  assign n6097 = ~n6095 & ~n6096;
  assign n6098 = ~n5789 & n6011;
  assign n6099 = ~n6012 & ~n6098;
  assign n6100 = ~n2006 & n4006;
  assign n6101 = ~n1900 & n4133;
  assign n6102 = n4002 & n5344;
  assign n6103 = ~n1811 & n4555;
  assign n6104 = ~n6102 & ~n6103;
  assign n6105 = ~n6101 & n6104;
  assign n6106 = ~n6100 & n6105;
  assign n6107 = pi29  & n6106;
  assign n6108 = ~pi29  & ~n6106;
  assign n6109 = ~n6107 & ~n6108;
  assign n6110 = n6099 & ~n6109;
  assign n6111 = ~n1740 & n4601;
  assign n6112 = ~n1610 & n4783;
  assign n6113 = n4602 & n4708;
  assign n6114 = ~n1531 & n4801;
  assign n6115 = ~n6113 & ~n6114;
  assign n6116 = ~n6112 & n6115;
  assign n6117 = ~n6111 & n6116;
  assign n6118 = pi26  & n6117;
  assign n6119 = ~pi26  & ~n6117;
  assign n6120 = ~n6118 & ~n6119;
  assign n6121 = ~n6099 & n6109;
  assign n6122 = ~n6120 & ~n6121;
  assign n6123 = ~n6110 & ~n6122;
  assign n6124 = n6097 & ~n6123;
  assign n6125 = ~n6095 & ~n6124;
  assign n6126 = ~n6018 & ~n6019;
  assign n6127 = ~n6029 & n6126;
  assign n6128 = n6029 & ~n6126;
  assign n6129 = ~n6127 & ~n6128;
  assign n6130 = ~n6125 & n6129;
  assign n6131 = n6125 & ~n6129;
  assign n6132 = ~n1230 & n5238;
  assign n6133 = n71 & ~n1107;
  assign n6134 = n4307 & n5239;
  assign n6135 = ~n1005 & n5326;
  assign n6136 = ~n6134 & ~n6135;
  assign n6137 = ~n6133 & n6136;
  assign n6138 = ~n6132 & n6137;
  assign n6139 = pi23  & n6138;
  assign n6140 = ~pi23  & ~n6138;
  assign n6141 = ~n6139 & ~n6140;
  assign n6142 = ~n6131 & ~n6141;
  assign n6143 = ~n6130 & ~n6142;
  assign n6144 = n6082 & ~n6143;
  assign n6145 = ~n6082 & n6143;
  assign n6146 = ~n795 & n5435;
  assign n6147 = ~n665 & n6055;
  assign n6148 = n4015 & n5429;
  assign n6149 = ~n720 & n6071;
  assign n6150 = ~n6148 & ~n6149;
  assign n6151 = ~n6147 & n6150;
  assign n6152 = ~n6146 & n6151;
  assign n6153 = pi20  & n6152;
  assign n6154 = ~pi20  & ~n6152;
  assign n6155 = ~n6153 & ~n6154;
  assign n6156 = ~n6145 & ~n6155;
  assign n6157 = ~n6144 & ~n6156;
  assign n6158 = ~n6078 & ~n6157;
  assign n6159 = n5643 & n6045;
  assign n6160 = ~n6046 & ~n6159;
  assign n6161 = n6078 & n6157;
  assign n6162 = ~n6158 & ~n6161;
  assign n6163 = n6160 & n6162;
  assign n6164 = ~n6158 & ~n6163;
  assign n6165 = ~n6052 & ~n6053;
  assign n6166 = ~n6062 & n6165;
  assign n6167 = n6062 & ~n6165;
  assign n6168 = ~n6166 & ~n6167;
  assign n6169 = ~n6164 & n6168;
  assign n6170 = n6164 & ~n6168;
  assign n6171 = ~n6169 & ~n6170;
  assign n6172 = ~n6160 & ~n6162;
  assign n6173 = ~n6163 & ~n6172;
  assign n6174 = pi16  & ~pi17 ;
  assign n6175 = ~pi16  & pi17 ;
  assign n6176 = ~n6174 & ~n6175;
  assign n6177 = ~pi15  & pi16 ;
  assign n6178 = pi15  & ~pi16 ;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = pi14  & ~pi15 ;
  assign n6181 = ~pi14  & pi15 ;
  assign n6182 = ~n6180 & ~n6181;
  assign n6183 = n6179 & n6182;
  assign n6184 = ~n6176 & n6183;
  assign n6185 = ~n6176 & ~n6182;
  assign n6186 = ~n3638 & n6185;
  assign n6187 = ~n6184 & ~n6186;
  assign n6188 = ~n554 & ~n6187;
  assign n6189 = pi17  & ~n6188;
  assign n6190 = ~pi17  & n6188;
  assign n6191 = ~n6189 & ~n6190;
  assign n6192 = ~n1338 & n5238;
  assign n6193 = n71 & ~n1230;
  assign n6194 = n4323 & n5239;
  assign n6195 = ~n1107 & n5326;
  assign n6196 = ~n6194 & ~n6195;
  assign n6197 = ~n6193 & n6196;
  assign n6198 = ~n6192 & n6197;
  assign n6199 = ~pi23  & ~n6198;
  assign n6200 = pi23  & n6198;
  assign n6201 = ~n6199 & ~n6200;
  assign n6202 = ~n6097 & n6123;
  assign n6203 = ~n6124 & ~n6202;
  assign n6204 = ~n6201 & n6203;
  assign n6205 = ~n6201 & ~n6203;
  assign n6206 = n6201 & n6203;
  assign n6207 = ~n6205 & ~n6206;
  assign n6208 = ~n6110 & ~n6121;
  assign n6209 = n6120 & ~n6208;
  assign n6210 = ~n6120 & n6208;
  assign n6211 = ~n6209 & ~n6210;
  assign n6212 = ~n5999 & n6009;
  assign n6213 = ~n6010 & ~n6212;
  assign n6214 = ~n5829 & n5986;
  assign n6215 = ~n5987 & ~n6214;
  assign n6216 = ~n2554 & n3641;
  assign n6217 = n3557 & ~n3559;
  assign n6218 = ~n3560 & ~n6217;
  assign n6219 = n556 & n6218;
  assign n6220 = ~n2369 & n3961;
  assign n6221 = ~n2457 & n3740;
  assign n6222 = ~n6220 & ~n6221;
  assign n6223 = ~n6219 & n6222;
  assign n6224 = ~n6216 & n6223;
  assign n6225 = n6215 & ~n6224;
  assign n6226 = ~n2278 & n4006;
  assign n6227 = ~n2178 & n4133;
  assign n6228 = n4002 & n5538;
  assign n6229 = ~n2058 & n4555;
  assign n6230 = ~n6228 & ~n6229;
  assign n6231 = ~n6227 & n6230;
  assign n6232 = ~n6226 & n6231;
  assign n6233 = ~pi29  & ~n6232;
  assign n6234 = pi29  & n6232;
  assign n6235 = ~n6233 & ~n6234;
  assign n6236 = n6215 & n6224;
  assign n6237 = ~n6215 & ~n6224;
  assign n6238 = ~n6236 & ~n6237;
  assign n6239 = ~n6235 & ~n6238;
  assign n6240 = ~n6225 & ~n6239;
  assign n6241 = n5988 & ~n5990;
  assign n6242 = ~n5991 & ~n6241;
  assign n6243 = ~n6240 & n6242;
  assign n6244 = ~n2178 & n4006;
  assign n6245 = ~n2058 & n4133;
  assign n6246 = n4002 & n5554;
  assign n6247 = ~n2006 & n4555;
  assign n6248 = ~n6246 & ~n6247;
  assign n6249 = ~n6245 & n6248;
  assign n6250 = ~n6244 & n6249;
  assign n6251 = pi29  & n6250;
  assign n6252 = ~pi29  & ~n6250;
  assign n6253 = ~n6251 & ~n6252;
  assign n6254 = n6240 & ~n6242;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n6243 & ~n6255;
  assign n6257 = n6213 & ~n6256;
  assign n6258 = ~n6213 & n6256;
  assign n6259 = ~n1811 & n4601;
  assign n6260 = ~n1740 & n4783;
  assign n6261 = n4602 & n4951;
  assign n6262 = ~n1610 & n4801;
  assign n6263 = ~n6261 & ~n6262;
  assign n6264 = ~n6260 & n6263;
  assign n6265 = ~n6259 & n6264;
  assign n6266 = pi26  & n6265;
  assign n6267 = ~pi26  & ~n6265;
  assign n6268 = ~n6266 & ~n6267;
  assign n6269 = ~n6258 & ~n6268;
  assign n6270 = ~n6257 & ~n6269;
  assign n6271 = n6211 & ~n6270;
  assign n6272 = ~n6211 & n6270;
  assign n6273 = ~n1426 & n5238;
  assign n6274 = n71 & ~n1338;
  assign n6275 = n4753 & n5239;
  assign n6276 = ~n1230 & n5326;
  assign n6277 = ~n6275 & ~n6276;
  assign n6278 = ~n6274 & n6277;
  assign n6279 = ~n6273 & n6278;
  assign n6280 = pi23  & n6279;
  assign n6281 = ~pi23  & ~n6279;
  assign n6282 = ~n6280 & ~n6281;
  assign n6283 = ~n6272 & ~n6282;
  assign n6284 = ~n6271 & ~n6283;
  assign n6285 = ~n6207 & ~n6284;
  assign n6286 = ~n6204 & ~n6285;
  assign n6287 = ~n6130 & ~n6131;
  assign n6288 = ~n6141 & n6287;
  assign n6289 = n6141 & ~n6287;
  assign n6290 = ~n6288 & ~n6289;
  assign n6291 = ~n6286 & n6290;
  assign n6292 = n6286 & ~n6290;
  assign n6293 = ~n894 & n5435;
  assign n6294 = ~n795 & n6055;
  assign n6295 = n3959 & n5429;
  assign n6296 = ~n665 & n6071;
  assign n6297 = ~n6295 & ~n6296;
  assign n6298 = ~n6294 & n6297;
  assign n6299 = ~n6293 & n6298;
  assign n6300 = pi20  & n6299;
  assign n6301 = ~pi20  & ~n6299;
  assign n6302 = ~n6300 & ~n6301;
  assign n6303 = ~n6292 & ~n6302;
  assign n6304 = ~n6291 & ~n6303;
  assign n6305 = ~n6191 & ~n6304;
  assign n6306 = n6191 & n6304;
  assign n6307 = ~n6144 & ~n6145;
  assign n6308 = ~n6155 & n6307;
  assign n6309 = n6155 & ~n6307;
  assign n6310 = ~n6308 & ~n6309;
  assign n6311 = ~n6306 & n6310;
  assign n6312 = ~n6305 & ~n6311;
  assign n6313 = n6173 & ~n6312;
  assign n6314 = ~n6305 & ~n6306;
  assign n6315 = n6310 & n6314;
  assign n6316 = ~n6310 & ~n6314;
  assign n6317 = ~n6315 & ~n6316;
  assign n6318 = n6207 & n6284;
  assign n6319 = ~n6285 & ~n6318;
  assign n6320 = ~n1005 & n5435;
  assign n6321 = ~n894 & n6055;
  assign n6322 = n4122 & n5429;
  assign n6323 = ~n795 & n6071;
  assign n6324 = ~n6322 & ~n6323;
  assign n6325 = ~n6321 & n6324;
  assign n6326 = ~n6320 & n6325;
  assign n6327 = pi20  & n6326;
  assign n6328 = ~pi20  & ~n6326;
  assign n6329 = ~n6327 & ~n6328;
  assign n6330 = n6319 & ~n6329;
  assign n6331 = ~n6319 & n6329;
  assign n6332 = ~n6330 & ~n6331;
  assign n6333 = ~n6271 & ~n6272;
  assign n6334 = ~n6282 & n6333;
  assign n6335 = n6282 & ~n6333;
  assign n6336 = ~n6334 & ~n6335;
  assign n6337 = ~n1900 & n4601;
  assign n6338 = ~n1811 & n4783;
  assign n6339 = n4602 & n4967;
  assign n6340 = ~n1740 & n4801;
  assign n6341 = ~n6339 & ~n6340;
  assign n6342 = ~n6338 & n6341;
  assign n6343 = ~n6337 & n6342;
  assign n6344 = pi26  & n6343;
  assign n6345 = ~pi26  & ~n6343;
  assign n6346 = ~n6344 & ~n6345;
  assign n6347 = ~n6243 & ~n6254;
  assign n6348 = n6253 & ~n6347;
  assign n6349 = ~n6253 & n6347;
  assign n6350 = ~n6348 & ~n6349;
  assign n6351 = ~n6346 & n6350;
  assign n6352 = n6346 & ~n6350;
  assign n6353 = ~n6351 & ~n6352;
  assign n6354 = ~n5974 & ~n5975;
  assign n6355 = ~n5984 & n6354;
  assign n6356 = n5984 & ~n6354;
  assign n6357 = ~n6355 & ~n6356;
  assign n6358 = ~n354 & n1813;
  assign n6359 = ~n106 & n6358;
  assign n6360 = ~n500 & n1162;
  assign n6361 = n445 & n6360;
  assign n6362 = n4444 & n6361;
  assign n6363 = ~n160 & n6362;
  assign n6364 = n6359 & n6363;
  assign n6365 = n2192 & n2409;
  assign n6366 = ~n325 & n6365;
  assign n6367 = n1038 & n4168;
  assign n6368 = ~n94 & n6367;
  assign n6369 = ~n638 & n6368;
  assign n6370 = n6366 & n6369;
  assign n6371 = n6364 & n6370;
  assign n6372 = n1631 & n6371;
  assign n6373 = n758 & n6372;
  assign n6374 = ~n206 & n6373;
  assign n6375 = ~n324 & n6374;
  assign n6376 = ~n628 & ~n685;
  assign n6377 = ~n122 & n6376;
  assign n6378 = n1551 & n6377;
  assign n6379 = n1394 & n6378;
  assign n6380 = ~n180 & n6379;
  assign n6381 = ~n599 & n6380;
  assign n6382 = n6375 & n6381;
  assign n6383 = n4492 & n5889;
  assign n6384 = n1109 & n6383;
  assign n6385 = ~n171 & n6384;
  assign n6386 = n4872 & n5907;
  assign n6387 = ~n414 & n6386;
  assign n6388 = n6385 & n6387;
  assign n6389 = n6382 & n6388;
  assign n6390 = n5902 & ~n6389;
  assign n6391 = ~n5902 & n6389;
  assign n6392 = ~n6390 & ~n6391;
  assign n6393 = ~n466 & ~n469;
  assign n6394 = n1153 & n6393;
  assign n6395 = ~n423 & n6394;
  assign n6396 = ~n637 & n2294;
  assign n6397 = ~n325 & n6396;
  assign n6398 = n6395 & n6397;
  assign n6399 = n1275 & n6398;
  assign n6400 = n1148 & n6399;
  assign n6401 = ~n154 & n6400;
  assign n6402 = ~n669 & n6401;
  assign n6403 = n787 & n4061;
  assign n6404 = ~n612 & n6403;
  assign n6405 = ~n613 & n6404;
  assign n6406 = n6402 & n6405;
  assign n6407 = n3882 & n5038;
  assign n6408 = ~n518 & n6407;
  assign n6409 = ~n700 & n6408;
  assign n6410 = n1296 & n1544;
  assign n6411 = ~n331 & n6410;
  assign n6412 = ~n245 & n6411;
  assign n6413 = ~n147 & n6412;
  assign n6414 = n6409 & n6413;
  assign n6415 = n6406 & n6414;
  assign n6416 = ~pi2  & ~n6415;
  assign n6417 = pi2  & ~n6415;
  assign n6418 = ~pi2  & n6415;
  assign n6419 = ~n6417 & ~n6418;
  assign n6420 = ~pi5  & ~n6419;
  assign n6421 = ~n6416 & ~n6420;
  assign n6422 = n5902 & ~n6421;
  assign n6423 = ~n5902 & n6421;
  assign n6424 = ~n2803 & n3641;
  assign n6425 = ~n2748 & n3740;
  assign n6426 = n3541 & ~n3543;
  assign n6427 = ~n3544 & ~n6426;
  assign n6428 = n556 & n6427;
  assign n6429 = ~n2676 & n3961;
  assign n6430 = ~n6428 & ~n6429;
  assign n6431 = ~n6425 & n6430;
  assign n6432 = ~n6424 & n6431;
  assign n6433 = ~n6423 & ~n6432;
  assign n6434 = ~n6422 & ~n6433;
  assign n6435 = n6392 & ~n6434;
  assign n6436 = ~n6390 & ~n6435;
  assign n6437 = ~pi8  & ~n5972;
  assign n6438 = ~n5970 & n5973;
  assign n6439 = ~n6437 & ~n6438;
  assign n6440 = ~n6436 & ~n6439;
  assign n6441 = n6436 & n6439;
  assign n6442 = ~n2676 & n3641;
  assign n6443 = ~n2640 & n3740;
  assign n6444 = n3549 & ~n3551;
  assign n6445 = ~n3552 & ~n6444;
  assign n6446 = n556 & n6445;
  assign n6447 = ~n2554 & n3961;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = ~n6443 & n6448;
  assign n6450 = ~n6442 & n6449;
  assign n6451 = ~n6441 & ~n6450;
  assign n6452 = ~n6440 & ~n6451;
  assign n6453 = n6357 & ~n6452;
  assign n6454 = ~n6357 & n6452;
  assign n6455 = ~n6453 & ~n6454;
  assign n6456 = ~n2369 & n4006;
  assign n6457 = ~n2278 & n4133;
  assign n6458 = n4002 & n5779;
  assign n6459 = ~n2178 & n4555;
  assign n6460 = ~n6458 & ~n6459;
  assign n6461 = ~n6457 & n6460;
  assign n6462 = ~n6456 & n6461;
  assign n6463 = pi29  & n6462;
  assign n6464 = ~pi29  & ~n6462;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = n6455 & ~n6465;
  assign n6467 = ~n6453 & ~n6466;
  assign n6468 = n6235 & n6238;
  assign n6469 = ~n6239 & ~n6468;
  assign n6470 = ~n6467 & n6469;
  assign n6471 = n6467 & ~n6469;
  assign n6472 = ~n2006 & n4601;
  assign n6473 = ~n1900 & n4783;
  assign n6474 = n4602 & n5344;
  assign n6475 = ~n1811 & n4801;
  assign n6476 = ~n6474 & ~n6475;
  assign n6477 = ~n6473 & n6476;
  assign n6478 = ~n6472 & n6477;
  assign n6479 = pi26  & n6478;
  assign n6480 = ~pi26  & ~n6478;
  assign n6481 = ~n6479 & ~n6480;
  assign n6482 = ~n6471 & ~n6481;
  assign n6483 = ~n6470 & ~n6482;
  assign n6484 = n6353 & ~n6483;
  assign n6485 = ~n6351 & ~n6484;
  assign n6486 = ~n6257 & ~n6258;
  assign n6487 = ~n6268 & n6486;
  assign n6488 = n6268 & ~n6486;
  assign n6489 = ~n6487 & ~n6488;
  assign n6490 = ~n6485 & n6489;
  assign n6491 = n6485 & ~n6489;
  assign n6492 = ~n1531 & n5238;
  assign n6493 = n71 & ~n1426;
  assign n6494 = n4533 & n5239;
  assign n6495 = ~n1338 & n5326;
  assign n6496 = ~n6494 & ~n6495;
  assign n6497 = ~n6493 & n6496;
  assign n6498 = ~n6492 & n6497;
  assign n6499 = pi23  & n6498;
  assign n6500 = ~pi23  & ~n6498;
  assign n6501 = ~n6499 & ~n6500;
  assign n6502 = ~n6491 & ~n6501;
  assign n6503 = ~n6490 & ~n6502;
  assign n6504 = n6336 & ~n6503;
  assign n6505 = ~n6336 & n6503;
  assign n6506 = ~n1107 & n5435;
  assign n6507 = ~n1005 & n6055;
  assign n6508 = n4106 & n5429;
  assign n6509 = ~n894 & n6071;
  assign n6510 = ~n6508 & ~n6509;
  assign n6511 = ~n6507 & n6510;
  assign n6512 = ~n6506 & n6511;
  assign n6513 = pi20  & n6512;
  assign n6514 = ~pi20  & ~n6512;
  assign n6515 = ~n6513 & ~n6514;
  assign n6516 = ~n6505 & ~n6515;
  assign n6517 = ~n6504 & ~n6516;
  assign n6518 = n6332 & ~n6517;
  assign n6519 = ~n6330 & ~n6518;
  assign n6520 = ~n6291 & ~n6292;
  assign n6521 = ~n6302 & n6520;
  assign n6522 = n6302 & ~n6520;
  assign n6523 = ~n6521 & ~n6522;
  assign n6524 = ~n6519 & n6523;
  assign n6525 = n6519 & ~n6523;
  assign n6526 = ~n3744 & n6185;
  assign n6527 = ~n6179 & n6182;
  assign n6528 = ~n554 & n6527;
  assign n6529 = ~n720 & n6184;
  assign n6530 = ~n6528 & ~n6529;
  assign n6531 = ~n6526 & n6530;
  assign n6532 = pi17  & n6531;
  assign n6533 = ~pi17  & ~n6531;
  assign n6534 = ~n6532 & ~n6533;
  assign n6535 = ~n6525 & ~n6534;
  assign n6536 = ~n6524 & ~n6535;
  assign n6537 = n6317 & ~n6536;
  assign n6538 = ~n6317 & n6536;
  assign n6539 = ~n6537 & ~n6538;
  assign n6540 = ~n665 & n6184;
  assign n6541 = ~n720 & n6527;
  assign n6542 = n3979 & n6185;
  assign n6543 = n6176 & ~n6182;
  assign n6544 = ~n554 & n6543;
  assign n6545 = ~n6542 & ~n6544;
  assign n6546 = ~n6541 & n6545;
  assign n6547 = ~n6540 & n6546;
  assign n6548 = pi17  & n6547;
  assign n6549 = ~pi17  & ~n6547;
  assign n6550 = ~n6548 & ~n6549;
  assign n6551 = ~n6504 & ~n6505;
  assign n6552 = ~n6515 & n6551;
  assign n6553 = n6515 & ~n6551;
  assign n6554 = ~n6552 & ~n6553;
  assign n6555 = ~n1610 & n5238;
  assign n6556 = n71 & ~n1531;
  assign n6557 = n4724 & n5239;
  assign n6558 = ~n1426 & n5326;
  assign n6559 = ~n6557 & ~n6558;
  assign n6560 = ~n6556 & n6559;
  assign n6561 = ~n6555 & n6560;
  assign n6562 = ~pi23  & ~n6561;
  assign n6563 = pi23  & n6561;
  assign n6564 = ~n6562 & ~n6563;
  assign n6565 = ~n6353 & n6483;
  assign n6566 = ~n6484 & ~n6565;
  assign n6567 = ~n6564 & n6566;
  assign n6568 = ~n6564 & ~n6566;
  assign n6569 = n6564 & n6566;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = ~n6470 & ~n6471;
  assign n6572 = ~n6481 & n6571;
  assign n6573 = n6481 & ~n6571;
  assign n6574 = ~n6572 & ~n6573;
  assign n6575 = ~n2457 & n4006;
  assign n6576 = ~n2369 & n4133;
  assign n6577 = n4002 & n5795;
  assign n6578 = ~n2278 & n4555;
  assign n6579 = ~n6577 & ~n6578;
  assign n6580 = ~n6576 & n6579;
  assign n6581 = ~n6575 & n6580;
  assign n6582 = ~pi29  & ~n6581;
  assign n6583 = pi29  & n6581;
  assign n6584 = ~n6582 & ~n6583;
  assign n6585 = ~n6440 & ~n6441;
  assign n6586 = ~n6450 & n6585;
  assign n6587 = n6450 & ~n6585;
  assign n6588 = ~n6586 & ~n6587;
  assign n6589 = ~n6584 & n6588;
  assign n6590 = ~n6584 & ~n6588;
  assign n6591 = n6584 & n6588;
  assign n6592 = ~n6590 & ~n6591;
  assign n6593 = ~n6392 & n6434;
  assign n6594 = ~n6435 & ~n6593;
  assign n6595 = ~n2748 & n3641;
  assign n6596 = n3545 & ~n3547;
  assign n6597 = ~n3548 & ~n6596;
  assign n6598 = n556 & n6597;
  assign n6599 = ~n2640 & n3961;
  assign n6600 = ~n2676 & n3740;
  assign n6601 = ~n6599 & ~n6600;
  assign n6602 = ~n6598 & n6601;
  assign n6603 = ~n6595 & n6602;
  assign n6604 = n6594 & ~n6603;
  assign n6605 = ~n6422 & ~n6423;
  assign n6606 = ~n6432 & n6605;
  assign n6607 = n6432 & ~n6605;
  assign n6608 = ~n6606 & ~n6607;
  assign n6609 = n853 & n1090;
  assign n6610 = n744 & n6609;
  assign n6611 = ~n668 & n6610;
  assign n6612 = ~n427 & n3454;
  assign n6613 = ~n259 & n6612;
  assign n6614 = n6611 & n6613;
  assign n6615 = n3130 & n6614;
  assign n6616 = ~n395 & n6615;
  assign n6617 = n3820 & n5740;
  assign n6618 = ~n454 & n6617;
  assign n6619 = n6616 & n6618;
  assign n6620 = ~n170 & ~n290;
  assign n6621 = ~n172 & n6620;
  assign n6622 = ~n685 & n2814;
  assign n6623 = ~n683 & n6622;
  assign n6624 = n6621 & n6623;
  assign n6625 = n5087 & n5804;
  assign n6626 = n6624 & n6625;
  assign n6627 = n1221 & n6626;
  assign n6628 = ~n422 & n6627;
  assign n6629 = n1970 & n2870;
  assign n6630 = n226 & n6629;
  assign n6631 = n615 & n6630;
  assign n6632 = ~n245 & n6631;
  assign n6633 = n6628 & n6632;
  assign n6634 = n6619 & n6633;
  assign n6635 = pi2  & ~n6634;
  assign n6636 = n1063 & n5154;
  assign n6637 = n1708 & n6636;
  assign n6638 = ~n94 & n6637;
  assign n6639 = n4175 & n4427;
  assign n6640 = n5493 & n6639;
  assign n6641 = n528 & n6640;
  assign n6642 = n1516 & n6641;
  assign n6643 = ~n337 & n6642;
  assign n6644 = ~n382 & n6643;
  assign n6645 = n6638 & n6644;
  assign n6646 = n3338 & n3830;
  assign n6647 = n2231 & n6646;
  assign n6648 = ~n533 & n6647;
  assign n6649 = n1241 & n1416;
  assign n6650 = n174 & n6649;
  assign n6651 = ~n518 & n6650;
  assign n6652 = ~n473 & n6651;
  assign n6653 = n6648 & n6652;
  assign n6654 = n6645 & n6653;
  assign n6655 = pi2  & ~n6654;
  assign n6656 = ~pi2  & n6654;
  assign n6657 = ~n6655 & ~n6656;
  assign n6658 = ~n672 & n1505;
  assign n6659 = ~n232 & n6658;
  assign n6660 = ~n428 & ~n627;
  assign n6661 = ~n436 & n6660;
  assign n6662 = n6659 & n6661;
  assign n6663 = n2191 & n3919;
  assign n6664 = n1110 & n6663;
  assign n6665 = n528 & n6664;
  assign n6666 = ~n334 & n6665;
  assign n6667 = n1221 & n3320;
  assign n6668 = n5897 & n6667;
  assign n6669 = n5812 & n6668;
  assign n6670 = ~n689 & n6669;
  assign n6671 = n6666 & n6670;
  assign n6672 = ~n279 & n6671;
  assign n6673 = ~n372 & n684;
  assign n6674 = ~n400 & n6673;
  assign n6675 = n6672 & n6674;
  assign n6676 = n2104 & n6675;
  assign n6677 = n6662 & n6676;
  assign n6678 = n2940 & n3899;
  assign n6679 = n3392 & n6678;
  assign n6680 = n5150 & n6679;
  assign n6681 = n3820 & n6680;
  assign n6682 = n3411 & n3927;
  assign n6683 = n1362 & n6682;
  assign n6684 = ~n462 & n6683;
  assign n6685 = n6681 & n6684;
  assign n6686 = ~n236 & n6685;
  assign n6687 = n5505 & n6686;
  assign n6688 = n6677 & n6687;
  assign n6689 = pi2  & ~n6688;
  assign n6690 = ~pi2  & n6688;
  assign n6691 = ~n3097 & n3641;
  assign n6692 = ~n3005 & n3740;
  assign n6693 = n3525 & ~n3527;
  assign n6694 = ~n3528 & ~n6693;
  assign n6695 = n556 & n6694;
  assign n6696 = ~n2927 & n3961;
  assign n6697 = ~n6695 & ~n6696;
  assign n6698 = ~n6692 & n6697;
  assign n6699 = ~n6691 & n6698;
  assign n6700 = ~n6690 & ~n6699;
  assign n6701 = ~n6689 & ~n6700;
  assign n6702 = n6657 & ~n6701;
  assign n6703 = ~n6655 & ~n6702;
  assign n6704 = ~pi2  & n6634;
  assign n6705 = ~n6635 & ~n6704;
  assign n6706 = ~n6703 & n6705;
  assign n6707 = ~n6635 & ~n6706;
  assign n6708 = pi5  & n6419;
  assign n6709 = ~n6420 & ~n6708;
  assign n6710 = ~n6707 & n6709;
  assign n6711 = n6707 & ~n6709;
  assign n6712 = ~n2891 & n3641;
  assign n6713 = ~n2803 & n3740;
  assign n6714 = n3537 & ~n3539;
  assign n6715 = ~n3540 & ~n6714;
  assign n6716 = n556 & n6715;
  assign n6717 = ~n2748 & n3961;
  assign n6718 = ~n6716 & ~n6717;
  assign n6719 = ~n6713 & n6718;
  assign n6720 = ~n6712 & n6719;
  assign n6721 = ~n6711 & ~n6720;
  assign n6722 = ~n6710 & ~n6721;
  assign n6723 = n6608 & ~n6722;
  assign n6724 = ~n6608 & n6722;
  assign n6725 = ~n6723 & ~n6724;
  assign n6726 = ~n2640 & n4006;
  assign n6727 = ~n2554 & n4133;
  assign n6728 = n4002 & n5979;
  assign n6729 = ~n2457 & n4555;
  assign n6730 = ~n6728 & ~n6729;
  assign n6731 = ~n6727 & n6730;
  assign n6732 = ~n6726 & n6731;
  assign n6733 = pi29  & n6732;
  assign n6734 = ~pi29  & ~n6732;
  assign n6735 = ~n6733 & ~n6734;
  assign n6736 = n6725 & ~n6735;
  assign n6737 = ~n6723 & ~n6736;
  assign n6738 = n6594 & n6603;
  assign n6739 = ~n6594 & ~n6603;
  assign n6740 = ~n6738 & ~n6739;
  assign n6741 = ~n6737 & ~n6740;
  assign n6742 = ~n6604 & ~n6741;
  assign n6743 = ~n6592 & ~n6742;
  assign n6744 = ~n6589 & ~n6743;
  assign n6745 = ~n6455 & n6465;
  assign n6746 = ~n6466 & ~n6745;
  assign n6747 = ~n6744 & n6746;
  assign n6748 = n6744 & ~n6746;
  assign n6749 = ~n2058 & n4601;
  assign n6750 = ~n2006 & n4783;
  assign n6751 = n4602 & n5180;
  assign n6752 = ~n1900 & n4801;
  assign n6753 = ~n6751 & ~n6752;
  assign n6754 = ~n6750 & n6753;
  assign n6755 = ~n6749 & n6754;
  assign n6756 = pi26  & n6755;
  assign n6757 = ~pi26  & ~n6755;
  assign n6758 = ~n6756 & ~n6757;
  assign n6759 = ~n6748 & ~n6758;
  assign n6760 = ~n6747 & ~n6759;
  assign n6761 = n6574 & ~n6760;
  assign n6762 = ~n6574 & n6760;
  assign n6763 = ~n1740 & n5238;
  assign n6764 = n71 & ~n1610;
  assign n6765 = n4708 & n5239;
  assign n6766 = ~n1531 & n5326;
  assign n6767 = ~n6765 & ~n6766;
  assign n6768 = ~n6764 & n6767;
  assign n6769 = ~n6763 & n6768;
  assign n6770 = pi23  & n6769;
  assign n6771 = ~pi23  & ~n6769;
  assign n6772 = ~n6770 & ~n6771;
  assign n6773 = ~n6762 & ~n6772;
  assign n6774 = ~n6761 & ~n6773;
  assign n6775 = ~n6570 & ~n6774;
  assign n6776 = ~n6567 & ~n6775;
  assign n6777 = ~n6490 & ~n6491;
  assign n6778 = ~n6501 & n6777;
  assign n6779 = n6501 & ~n6777;
  assign n6780 = ~n6778 & ~n6779;
  assign n6781 = ~n6776 & n6780;
  assign n6782 = n6776 & ~n6780;
  assign n6783 = ~n1230 & n5435;
  assign n6784 = ~n1107 & n6055;
  assign n6785 = n4307 & n5429;
  assign n6786 = ~n1005 & n6071;
  assign n6787 = ~n6785 & ~n6786;
  assign n6788 = ~n6784 & n6787;
  assign n6789 = ~n6783 & n6788;
  assign n6790 = pi20  & n6789;
  assign n6791 = ~pi20  & ~n6789;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = ~n6782 & ~n6792;
  assign n6794 = ~n6781 & ~n6793;
  assign n6795 = n6554 & ~n6794;
  assign n6796 = ~n6554 & n6794;
  assign n6797 = ~n795 & n6184;
  assign n6798 = ~n665 & n6527;
  assign n6799 = n4015 & n6185;
  assign n6800 = ~n720 & n6543;
  assign n6801 = ~n6799 & ~n6800;
  assign n6802 = ~n6798 & n6801;
  assign n6803 = ~n6797 & n6802;
  assign n6804 = pi17  & n6803;
  assign n6805 = ~pi17  & ~n6803;
  assign n6806 = ~n6804 & ~n6805;
  assign n6807 = ~n6796 & ~n6806;
  assign n6808 = ~n6795 & ~n6807;
  assign n6809 = ~n6550 & ~n6808;
  assign n6810 = n6550 & n6808;
  assign n6811 = ~n6809 & ~n6810;
  assign n6812 = ~n6332 & n6517;
  assign n6813 = ~n6518 & ~n6812;
  assign n6814 = n6811 & n6813;
  assign n6815 = ~n6809 & ~n6814;
  assign n6816 = ~n6524 & ~n6525;
  assign n6817 = ~n6534 & n6816;
  assign n6818 = n6534 & ~n6816;
  assign n6819 = ~n6817 & ~n6818;
  assign n6820 = ~n6815 & n6819;
  assign n6821 = n6815 & ~n6819;
  assign n6822 = ~n6820 & ~n6821;
  assign n6823 = ~n6811 & ~n6813;
  assign n6824 = ~n6814 & ~n6823;
  assign n6825 = pi13  & ~pi14 ;
  assign n6826 = ~pi13  & pi14 ;
  assign n6827 = ~n6825 & ~n6826;
  assign n6828 = ~pi12  & pi13 ;
  assign n6829 = pi12  & ~pi13 ;
  assign n6830 = ~n6828 & ~n6829;
  assign n6831 = pi11  & ~pi12 ;
  assign n6832 = ~pi11  & pi12 ;
  assign n6833 = ~n6831 & ~n6832;
  assign n6834 = n6830 & n6833;
  assign n6835 = ~n6827 & n6834;
  assign n6836 = ~n6827 & ~n6833;
  assign n6837 = ~n3638 & n6836;
  assign n6838 = ~n6835 & ~n6837;
  assign n6839 = ~n554 & ~n6838;
  assign n6840 = pi14  & ~n6839;
  assign n6841 = ~pi14  & n6839;
  assign n6842 = ~n6840 & ~n6841;
  assign n6843 = n6570 & n6774;
  assign n6844 = ~n6775 & ~n6843;
  assign n6845 = ~n1338 & n5435;
  assign n6846 = ~n1230 & n6055;
  assign n6847 = n4323 & n5429;
  assign n6848 = ~n1107 & n6071;
  assign n6849 = ~n6847 & ~n6848;
  assign n6850 = ~n6846 & n6849;
  assign n6851 = ~n6845 & n6850;
  assign n6852 = pi20  & n6851;
  assign n6853 = ~pi20  & ~n6851;
  assign n6854 = ~n6852 & ~n6853;
  assign n6855 = n6844 & ~n6854;
  assign n6856 = ~n6844 & n6854;
  assign n6857 = ~n6855 & ~n6856;
  assign n6858 = ~n6761 & ~n6762;
  assign n6859 = ~n6772 & n6858;
  assign n6860 = n6772 & ~n6858;
  assign n6861 = ~n6859 & ~n6860;
  assign n6862 = n6592 & n6742;
  assign n6863 = ~n6743 & ~n6862;
  assign n6864 = ~n2178 & n4601;
  assign n6865 = ~n2058 & n4783;
  assign n6866 = n4602 & n5554;
  assign n6867 = ~n2006 & n4801;
  assign n6868 = ~n6866 & ~n6867;
  assign n6869 = ~n6865 & n6868;
  assign n6870 = ~n6864 & n6869;
  assign n6871 = pi26  & n6870;
  assign n6872 = ~pi26  & ~n6870;
  assign n6873 = ~n6871 & ~n6872;
  assign n6874 = n6863 & ~n6873;
  assign n6875 = ~n6863 & n6873;
  assign n6876 = ~n6874 & ~n6875;
  assign n6877 = ~n2554 & n4006;
  assign n6878 = ~n2457 & n4133;
  assign n6879 = n4002 & n6218;
  assign n6880 = ~n2369 & n4555;
  assign n6881 = ~n6879 & ~n6880;
  assign n6882 = ~n6878 & n6881;
  assign n6883 = ~n6877 & n6882;
  assign n6884 = pi29  & n6883;
  assign n6885 = ~pi29  & ~n6883;
  assign n6886 = ~n6884 & ~n6885;
  assign n6887 = n6737 & n6740;
  assign n6888 = ~n6741 & ~n6887;
  assign n6889 = ~n6886 & n6888;
  assign n6890 = n6886 & ~n6888;
  assign n6891 = ~n2278 & n4601;
  assign n6892 = ~n2178 & n4783;
  assign n6893 = n4602 & n5538;
  assign n6894 = ~n2058 & n4801;
  assign n6895 = ~n6893 & ~n6894;
  assign n6896 = ~n6892 & n6895;
  assign n6897 = ~n6891 & n6896;
  assign n6898 = pi26  & n6897;
  assign n6899 = ~pi26  & ~n6897;
  assign n6900 = ~n6898 & ~n6899;
  assign n6901 = ~n6890 & ~n6900;
  assign n6902 = ~n6889 & ~n6901;
  assign n6903 = n6876 & ~n6902;
  assign n6904 = ~n6874 & ~n6903;
  assign n6905 = ~n6747 & ~n6748;
  assign n6906 = ~n6758 & n6905;
  assign n6907 = n6758 & ~n6905;
  assign n6908 = ~n6906 & ~n6907;
  assign n6909 = ~n6904 & n6908;
  assign n6910 = n6904 & ~n6908;
  assign n6911 = ~n1811 & n5238;
  assign n6912 = n71 & ~n1740;
  assign n6913 = n4951 & n5239;
  assign n6914 = ~n1610 & n5326;
  assign n6915 = ~n6913 & ~n6914;
  assign n6916 = ~n6912 & n6915;
  assign n6917 = ~n6911 & n6916;
  assign n6918 = pi23  & n6917;
  assign n6919 = ~pi23  & ~n6917;
  assign n6920 = ~n6918 & ~n6919;
  assign n6921 = ~n6910 & ~n6920;
  assign n6922 = ~n6909 & ~n6921;
  assign n6923 = n6861 & ~n6922;
  assign n6924 = ~n6861 & n6922;
  assign n6925 = ~n1426 & n5435;
  assign n6926 = ~n1338 & n6055;
  assign n6927 = n4753 & n5429;
  assign n6928 = ~n1230 & n6071;
  assign n6929 = ~n6927 & ~n6928;
  assign n6930 = ~n6926 & n6929;
  assign n6931 = ~n6925 & n6930;
  assign n6932 = pi20  & n6931;
  assign n6933 = ~pi20  & ~n6931;
  assign n6934 = ~n6932 & ~n6933;
  assign n6935 = ~n6924 & ~n6934;
  assign n6936 = ~n6923 & ~n6935;
  assign n6937 = n6857 & ~n6936;
  assign n6938 = ~n6855 & ~n6937;
  assign n6939 = ~n6781 & ~n6782;
  assign n6940 = ~n6792 & n6939;
  assign n6941 = n6792 & ~n6939;
  assign n6942 = ~n6940 & ~n6941;
  assign n6943 = ~n6938 & n6942;
  assign n6944 = n6938 & ~n6942;
  assign n6945 = ~n894 & n6184;
  assign n6946 = ~n795 & n6527;
  assign n6947 = n3959 & n6185;
  assign n6948 = ~n665 & n6543;
  assign n6949 = ~n6947 & ~n6948;
  assign n6950 = ~n6946 & n6949;
  assign n6951 = ~n6945 & n6950;
  assign n6952 = pi17  & n6951;
  assign n6953 = ~pi17  & ~n6951;
  assign n6954 = ~n6952 & ~n6953;
  assign n6955 = ~n6944 & ~n6954;
  assign n6956 = ~n6943 & ~n6955;
  assign n6957 = ~n6842 & ~n6956;
  assign n6958 = n6842 & n6956;
  assign n6959 = ~n6795 & ~n6796;
  assign n6960 = ~n6806 & n6959;
  assign n6961 = n6806 & ~n6959;
  assign n6962 = ~n6960 & ~n6961;
  assign n6963 = ~n6958 & n6962;
  assign n6964 = ~n6957 & ~n6963;
  assign n6965 = n6824 & ~n6964;
  assign n6966 = ~n6824 & n6964;
  assign n6967 = ~n6965 & ~n6966;
  assign n6968 = ~n1005 & n6184;
  assign n6969 = ~n894 & n6527;
  assign n6970 = n4122 & n6185;
  assign n6971 = ~n795 & n6543;
  assign n6972 = ~n6970 & ~n6971;
  assign n6973 = ~n6969 & n6972;
  assign n6974 = ~n6968 & n6973;
  assign n6975 = ~pi17  & ~n6974;
  assign n6976 = pi17  & n6974;
  assign n6977 = ~n6975 & ~n6976;
  assign n6978 = ~n6857 & n6936;
  assign n6979 = ~n6937 & ~n6978;
  assign n6980 = ~n6977 & n6979;
  assign n6981 = ~n6977 & ~n6979;
  assign n6982 = n6977 & n6979;
  assign n6983 = ~n6981 & ~n6982;
  assign n6984 = ~n6923 & ~n6924;
  assign n6985 = ~n6934 & n6984;
  assign n6986 = n6934 & ~n6984;
  assign n6987 = ~n6985 & ~n6986;
  assign n6988 = ~n1900 & n5238;
  assign n6989 = n71 & ~n1811;
  assign n6990 = n4967 & n5239;
  assign n6991 = ~n1740 & n5326;
  assign n6992 = ~n6990 & ~n6991;
  assign n6993 = ~n6989 & n6992;
  assign n6994 = ~n6988 & n6993;
  assign n6995 = ~pi23  & ~n6994;
  assign n6996 = pi23  & n6994;
  assign n6997 = ~n6995 & ~n6996;
  assign n6998 = ~n6876 & n6902;
  assign n6999 = ~n6903 & ~n6998;
  assign n7000 = ~n6997 & n6999;
  assign n7001 = ~n6997 & ~n6999;
  assign n7002 = n6997 & n6999;
  assign n7003 = ~n7001 & ~n7002;
  assign n7004 = ~n6889 & ~n6890;
  assign n7005 = ~n6900 & n7004;
  assign n7006 = n6900 & ~n7004;
  assign n7007 = ~n7005 & ~n7006;
  assign n7008 = ~n6725 & n6735;
  assign n7009 = ~n6736 & ~n7008;
  assign n7010 = n6703 & ~n6705;
  assign n7011 = ~n6706 & ~n7010;
  assign n7012 = ~n2927 & n3641;
  assign n7013 = n3533 & ~n3535;
  assign n7014 = ~n3536 & ~n7013;
  assign n7015 = n556 & n7014;
  assign n7016 = ~n2803 & n3961;
  assign n7017 = ~n2891 & n3740;
  assign n7018 = ~n7016 & ~n7017;
  assign n7019 = ~n7015 & n7018;
  assign n7020 = ~n7012 & n7019;
  assign n7021 = n7011 & ~n7020;
  assign n7022 = ~n6657 & n6701;
  assign n7023 = ~n6702 & ~n7022;
  assign n7024 = ~n3005 & n3641;
  assign n7025 = n3529 & ~n3531;
  assign n7026 = ~n3532 & ~n7025;
  assign n7027 = n556 & n7026;
  assign n7028 = ~n2891 & n3961;
  assign n7029 = ~n2927 & n3740;
  assign n7030 = ~n7028 & ~n7029;
  assign n7031 = ~n7027 & n7030;
  assign n7032 = ~n7024 & n7031;
  assign n7033 = n7023 & ~n7032;
  assign n7034 = n1153 & n3860;
  assign n7035 = n1575 & n7034;
  assign n7036 = n5081 & n7035;
  assign n7037 = ~n243 & n7036;
  assign n7038 = n119 & n5030;
  assign n7039 = ~n246 & n7038;
  assign n7040 = n7037 & n7039;
  assign n7041 = ~n232 & n5883;
  assign n7042 = ~n134 & n7041;
  assign n7043 = ~n106 & n7042;
  assign n7044 = n2529 & n7043;
  assign n7045 = n1708 & n7044;
  assign n7046 = ~n307 & n7045;
  assign n7047 = n3305 & n5143;
  assign n7048 = n1924 & n7047;
  assign n7049 = ~n315 & n7048;
  assign n7050 = n596 & n5056;
  assign n7051 = n1783 & n7050;
  assign n7052 = n901 & n7051;
  assign n7053 = ~n533 & n7052;
  assign n7054 = n7049 & n7053;
  assign n7055 = n376 & n5493;
  assign n7056 = ~n614 & n7055;
  assign n7057 = ~n326 & n2571;
  assign n7058 = ~n582 & n7057;
  assign n7059 = n7056 & n7058;
  assign n7060 = n7054 & n7059;
  assign n7061 = ~n149 & n1233;
  assign n7062 = ~n626 & n7061;
  assign n7063 = n7060 & n7062;
  assign n7064 = n528 & n7063;
  assign n7065 = ~n256 & n7064;
  assign n7066 = ~n633 & n7065;
  assign n7067 = n7046 & n7066;
  assign n7068 = n7040 & n7067;
  assign n7069 = ~n3166 & n3641;
  assign n7070 = n3521 & ~n3523;
  assign n7071 = ~n3524 & ~n7070;
  assign n7072 = n556 & n7071;
  assign n7073 = ~n3005 & n3961;
  assign n7074 = ~n3097 & n3740;
  assign n7075 = ~n7073 & ~n7074;
  assign n7076 = ~n7072 & n7075;
  assign n7077 = ~n7069 & n7076;
  assign n7078 = ~n7068 & ~n7077;
  assign n7079 = n902 & n1361;
  assign n7080 = n1182 & n7079;
  assign n7081 = n2491 & n7080;
  assign n7082 = n1513 & n7081;
  assign n7083 = ~n235 & n7082;
  assign n7084 = n3897 & n5744;
  assign n7085 = ~n611 & n7084;
  assign n7086 = ~n576 & n7085;
  assign n7087 = n7083 & n7086;
  assign n7088 = ~n294 & n1516;
  assign n7089 = ~n183 & ~n246;
  assign n7090 = ~n354 & n7089;
  assign n7091 = n7088 & n7090;
  assign n7092 = n2467 & n7091;
  assign n7093 = n1742 & n7092;
  assign n7094 = n2529 & n7093;
  assign n7095 = n437 & n7094;
  assign n7096 = ~n372 & n7095;
  assign n7097 = ~n208 & ~n245;
  assign n7098 = n1147 & n5687;
  assign n7099 = n162 & n1340;
  assign n7100 = ~n600 & n7099;
  assign n7101 = n7098 & n7100;
  assign n7102 = ~n360 & ~n698;
  assign n7103 = ~n254 & n7102;
  assign n7104 = n4912 & n7103;
  assign n7105 = ~n278 & n7104;
  assign n7106 = n148 & ~n589;
  assign n7107 = ~n297 & n7106;
  assign n7108 = ~n390 & n7107;
  assign n7109 = n7105 & n7108;
  assign n7110 = n7101 & n7109;
  assign n7111 = n7097 & n7110;
  assign n7112 = ~n331 & n1923;
  assign n7113 = ~n695 & n7112;
  assign n7114 = n7111 & n7113;
  assign n7115 = ~n173 & n7114;
  assign n7116 = ~n171 & n7115;
  assign n7117 = n7096 & n7116;
  assign n7118 = n7087 & n7117;
  assign n7119 = ~n3226 & n3641;
  assign n7120 = n3517 & ~n3519;
  assign n7121 = ~n3520 & ~n7120;
  assign n7122 = n556 & n7121;
  assign n7123 = ~n3097 & n3961;
  assign n7124 = ~n3166 & n3740;
  assign n7125 = ~n7123 & ~n7124;
  assign n7126 = ~n7122 & n7125;
  assign n7127 = ~n7119 & n7126;
  assign n7128 = ~n7118 & ~n7127;
  assign n7129 = n2192 & n2380;
  assign n7130 = ~n326 & n7129;
  assign n7131 = ~n705 & n7130;
  assign n7132 = ~n279 & n754;
  assign n7133 = ~n538 & n7132;
  assign n7134 = ~n462 & n7133;
  assign n7135 = n476 & n7134;
  assign n7136 = ~n679 & n7135;
  assign n7137 = ~n208 & n7136;
  assign n7138 = ~n181 & n7137;
  assign n7139 = n7131 & n7138;
  assign n7140 = n3382 & n7139;
  assign n7141 = ~n666 & n777;
  assign n7142 = ~n360 & n7141;
  assign n7143 = ~n194 & n7142;
  assign n7144 = ~n636 & n7143;
  assign n7145 = ~n155 & n7144;
  assign n7146 = ~n260 & n7145;
  assign n7147 = n5820 & n7146;
  assign n7148 = n7140 & n7147;
  assign n7149 = n2294 & n7148;
  assign n7150 = ~n243 & n7149;
  assign n7151 = ~n595 & n2921;
  assign n7152 = ~n129 & n7151;
  assign n7153 = ~n314 & n7152;
  assign n7154 = n1050 & n7153;
  assign n7155 = ~n362 & n7154;
  assign n7156 = ~n545 & n7155;
  assign n7157 = n7150 & n7156;
  assign n7158 = n827 & n3087;
  assign n7159 = ~n442 & n7158;
  assign n7160 = ~n427 & n1757;
  assign n7161 = ~n518 & n7160;
  assign n7162 = n1395 & n7161;
  assign n7163 = ~n594 & ~n685;
  assign n7164 = ~n239 & n1340;
  assign n7165 = n7163 & n7164;
  assign n7166 = n2991 & n7165;
  assign n7167 = n7162 & n7166;
  assign n7168 = n5858 & n7167;
  assign n7169 = ~n104 & n7168;
  assign n7170 = ~n682 & n7169;
  assign n7171 = n7159 & n7170;
  assign n7172 = n7157 & n7171;
  assign n7173 = ~n3263 & n3641;
  assign n7174 = n3513 & ~n3515;
  assign n7175 = ~n3516 & ~n7174;
  assign n7176 = n556 & n7175;
  assign n7177 = ~n3166 & n3961;
  assign n7178 = ~n3226 & n3740;
  assign n7179 = ~n7177 & ~n7178;
  assign n7180 = ~n7176 & n7179;
  assign n7181 = ~n7173 & n7180;
  assign n7182 = ~n7172 & ~n7181;
  assign n7183 = ~n78 & ~n218;
  assign n7184 = ~n468 & n7183;
  assign n7185 = n392 & ~n441;
  assign n7186 = ~n150 & n7185;
  assign n7187 = n7184 & n7186;
  assign n7188 = n459 & n7187;
  assign n7189 = n2970 & n4251;
  assign n7190 = n857 & n7189;
  assign n7191 = n7188 & n7190;
  assign n7192 = ~n204 & n7191;
  assign n7193 = ~n147 & n7192;
  assign n7194 = ~n475 & n7193;
  assign n7195 = n230 & ~n536;
  assign n7196 = n174 & ~n383;
  assign n7197 = ~n601 & n7196;
  assign n7198 = n2392 & n7197;
  assign n7199 = n1617 & n7198;
  assign n7200 = n584 & n2345;
  assign n7201 = ~n198 & n7200;
  assign n7202 = ~n690 & n1025;
  assign n7203 = ~n626 & n7202;
  assign n7204 = n7201 & n7203;
  assign n7205 = n396 & ~n666;
  assign n7206 = ~n502 & n7205;
  assign n7207 = ~n629 & n4636;
  assign n7208 = ~n344 & n7207;
  assign n7209 = n7206 & n7208;
  assign n7210 = n7204 & n7209;
  assign n7211 = n5150 & n7210;
  assign n7212 = n467 & n7211;
  assign n7213 = n7199 & n7212;
  assign n7214 = ~n275 & n7213;
  assign n7215 = ~n682 & n7214;
  assign n7216 = n7195 & n7215;
  assign n7217 = n1902 & n7216;
  assign n7218 = n7194 & n7217;
  assign n7219 = ~n3360 & n3641;
  assign n7220 = n3509 & ~n3511;
  assign n7221 = ~n3512 & ~n7220;
  assign n7222 = n556 & n7221;
  assign n7223 = ~n3226 & n3961;
  assign n7224 = ~n3263 & n3740;
  assign n7225 = ~n7223 & ~n7224;
  assign n7226 = ~n7222 & n7225;
  assign n7227 = ~n7219 & n7226;
  assign n7228 = ~n7218 & ~n7227;
  assign n7229 = ~n7218 & n7227;
  assign n7230 = n7218 & ~n7227;
  assign n7231 = ~n7229 & ~n7230;
  assign n7232 = ~n180 & n910;
  assign n7233 = ~n187 & ~n610;
  assign n7234 = n7232 & n7233;
  assign n7235 = ~n154 & n7234;
  assign n7236 = ~n631 & n3460;
  assign n7237 = ~n115 & n7236;
  assign n7238 = n7235 & n7237;
  assign n7239 = n1482 & n7238;
  assign n7240 = ~n685 & n7239;
  assign n7241 = ~n362 & n7240;
  assign n7242 = n1246 & n4256;
  assign n7243 = ~n593 & n7242;
  assign n7244 = ~n518 & n7243;
  assign n7245 = n7241 & n7244;
  assign n7246 = n2846 & n4923;
  assign n7247 = n1775 & n7246;
  assign n7248 = ~n305 & n7247;
  assign n7249 = ~n637 & n7248;
  assign n7250 = ~n667 & n4192;
  assign n7251 = ~n381 & n7250;
  assign n7252 = n1147 & n7251;
  assign n7253 = n1700 & n7252;
  assign n7254 = n2505 & n7253;
  assign n7255 = n1252 & n7254;
  assign n7256 = n954 & n7255;
  assign n7257 = ~n208 & n7256;
  assign n7258 = ~n582 & n7257;
  assign n7259 = n7249 & n7258;
  assign n7260 = n7245 & n7259;
  assign n7261 = ~n3450 & n3641;
  assign n7262 = n3450 & ~n3506;
  assign n7263 = n3360 & ~n7262;
  assign n7264 = ~n3360 & n7262;
  assign n7265 = ~n7263 & ~n7264;
  assign n7266 = n556 & n7265;
  assign n7267 = ~n3360 & n3961;
  assign n7268 = ~n3506 & n3740;
  assign n7269 = ~n7267 & ~n7268;
  assign n7270 = ~n7266 & n7269;
  assign n7271 = ~n7261 & n7270;
  assign n7272 = ~n7260 & ~n7271;
  assign n7273 = n2209 & n2440;
  assign n7274 = n1181 & n7273;
  assign n7275 = ~n106 & n7274;
  assign n7276 = n3354 & n3771;
  assign n7277 = ~n154 & n7276;
  assign n7278 = ~n181 & n7277;
  assign n7279 = n7275 & n7278;
  assign n7280 = ~n122 & n910;
  assign n7281 = ~n229 & ~n632;
  assign n7282 = ~n580 & n7281;
  assign n7283 = ~n305 & n7282;
  assign n7284 = n7280 & n7283;
  assign n7285 = n2029 & n7284;
  assign n7286 = ~n400 & n7285;
  assign n7287 = ~n681 & n2843;
  assign n7288 = n3117 & n7287;
  assign n7289 = ~n254 & n7288;
  assign n7290 = ~n384 & n921;
  assign n7291 = ~n667 & n7290;
  assign n7292 = ~n123 & n2424;
  assign n7293 = ~n349 & n758;
  assign n7294 = n7292 & n7293;
  assign n7295 = n765 & n7294;
  assign n7296 = n7291 & n7295;
  assign n7297 = n1635 & n7296;
  assign n7298 = ~n155 & n7297;
  assign n7299 = ~n78 & n7298;
  assign n7300 = n7289 & n7299;
  assign n7301 = n1785 & n2280;
  assign n7302 = n1343 & n7301;
  assign n7303 = ~n544 & n7302;
  assign n7304 = ~n216 & n1036;
  assign n7305 = ~n236 & n7304;
  assign n7306 = n415 & n7305;
  assign n7307 = n467 & n7306;
  assign n7308 = ~n188 & n7307;
  assign n7309 = ~n289 & n7308;
  assign n7310 = n7303 & n7309;
  assign n7311 = n7300 & n7310;
  assign n7312 = ~n310 & n3714;
  assign n7313 = n7311 & n7312;
  assign n7314 = ~n693 & n7313;
  assign n7315 = ~n394 & n7314;
  assign n7316 = n7286 & n7315;
  assign n7317 = n7279 & n7316;
  assign n7318 = n7272 & ~n7317;
  assign n7319 = ~n7272 & n7317;
  assign n7320 = ~n3506 & n3641;
  assign n7321 = ~n3360 & n3740;
  assign n7322 = ~n3363 & ~n3507;
  assign n7323 = ~n3508 & ~n7322;
  assign n7324 = n556 & n7323;
  assign n7325 = ~n3263 & n3961;
  assign n7326 = ~n7324 & ~n7325;
  assign n7327 = ~n7321 & n7326;
  assign n7328 = ~n7320 & n7327;
  assign n7329 = ~n7319 & ~n7328;
  assign n7330 = ~n7318 & ~n7329;
  assign n7331 = ~n7231 & ~n7330;
  assign n7332 = ~n7228 & ~n7331;
  assign n7333 = ~n7172 & n7181;
  assign n7334 = n7172 & ~n7181;
  assign n7335 = ~n7333 & ~n7334;
  assign n7336 = ~n7332 & ~n7335;
  assign n7337 = ~n7182 & ~n7336;
  assign n7338 = ~n7118 & n7127;
  assign n7339 = n7118 & ~n7127;
  assign n7340 = ~n7338 & ~n7339;
  assign n7341 = ~n7337 & ~n7340;
  assign n7342 = ~n7128 & ~n7341;
  assign n7343 = ~n7068 & n7077;
  assign n7344 = n7068 & ~n7077;
  assign n7345 = ~n7343 & ~n7344;
  assign n7346 = ~n7342 & ~n7345;
  assign n7347 = ~n7078 & ~n7346;
  assign n7348 = ~n6689 & ~n6690;
  assign n7349 = ~n6699 & n7348;
  assign n7350 = n6699 & ~n7348;
  assign n7351 = ~n7349 & ~n7350;
  assign n7352 = ~n7347 & n7351;
  assign n7353 = n7347 & ~n7351;
  assign n7354 = ~n7352 & ~n7353;
  assign n7355 = ~n2891 & n4006;
  assign n7356 = ~n2803 & n4133;
  assign n7357 = n4002 & n6715;
  assign n7358 = ~n2748 & n4555;
  assign n7359 = ~n7357 & ~n7358;
  assign n7360 = ~n7356 & n7359;
  assign n7361 = ~n7355 & n7360;
  assign n7362 = pi29  & n7361;
  assign n7363 = ~pi29  & ~n7361;
  assign n7364 = ~n7362 & ~n7363;
  assign n7365 = n7354 & ~n7364;
  assign n7366 = ~n7352 & ~n7365;
  assign n7367 = n7023 & n7032;
  assign n7368 = ~n7023 & ~n7032;
  assign n7369 = ~n7367 & ~n7368;
  assign n7370 = ~n7366 & ~n7369;
  assign n7371 = ~n7033 & ~n7370;
  assign n7372 = n7011 & n7020;
  assign n7373 = ~n7011 & ~n7020;
  assign n7374 = ~n7372 & ~n7373;
  assign n7375 = ~n7371 & ~n7374;
  assign n7376 = ~n7021 & ~n7375;
  assign n7377 = ~n6710 & ~n6711;
  assign n7378 = ~n6720 & n7377;
  assign n7379 = n6720 & ~n7377;
  assign n7380 = ~n7378 & ~n7379;
  assign n7381 = ~n7376 & n7380;
  assign n7382 = n7376 & ~n7380;
  assign n7383 = ~n2676 & n4006;
  assign n7384 = ~n2640 & n4133;
  assign n7385 = n4002 & n6445;
  assign n7386 = ~n2554 & n4555;
  assign n7387 = ~n7385 & ~n7386;
  assign n7388 = ~n7384 & n7387;
  assign n7389 = ~n7383 & n7388;
  assign n7390 = pi29  & n7389;
  assign n7391 = ~pi29  & ~n7389;
  assign n7392 = ~n7390 & ~n7391;
  assign n7393 = ~n7382 & ~n7392;
  assign n7394 = ~n7381 & ~n7393;
  assign n7395 = n7009 & ~n7394;
  assign n7396 = ~n7009 & n7394;
  assign n7397 = ~n2369 & n4601;
  assign n7398 = ~n2278 & n4783;
  assign n7399 = n4602 & n5779;
  assign n7400 = ~n2178 & n4801;
  assign n7401 = ~n7399 & ~n7400;
  assign n7402 = ~n7398 & n7401;
  assign n7403 = ~n7397 & n7402;
  assign n7404 = pi26  & n7403;
  assign n7405 = ~pi26  & ~n7403;
  assign n7406 = ~n7404 & ~n7405;
  assign n7407 = ~n7396 & ~n7406;
  assign n7408 = ~n7395 & ~n7407;
  assign n7409 = n7007 & ~n7408;
  assign n7410 = ~n7007 & n7408;
  assign n7411 = ~n2006 & n5238;
  assign n7412 = n71 & ~n1900;
  assign n7413 = n5239 & n5344;
  assign n7414 = ~n1811 & n5326;
  assign n7415 = ~n7413 & ~n7414;
  assign n7416 = ~n7412 & n7415;
  assign n7417 = ~n7411 & n7416;
  assign n7418 = pi23  & n7417;
  assign n7419 = ~pi23  & ~n7417;
  assign n7420 = ~n7418 & ~n7419;
  assign n7421 = ~n7410 & ~n7420;
  assign n7422 = ~n7409 & ~n7421;
  assign n7423 = ~n7003 & ~n7422;
  assign n7424 = ~n7000 & ~n7423;
  assign n7425 = ~n6909 & ~n6910;
  assign n7426 = ~n6920 & n7425;
  assign n7427 = n6920 & ~n7425;
  assign n7428 = ~n7426 & ~n7427;
  assign n7429 = ~n7424 & n7428;
  assign n7430 = n7424 & ~n7428;
  assign n7431 = ~n1531 & n5435;
  assign n7432 = ~n1426 & n6055;
  assign n7433 = n4533 & n5429;
  assign n7434 = ~n1338 & n6071;
  assign n7435 = ~n7433 & ~n7434;
  assign n7436 = ~n7432 & n7435;
  assign n7437 = ~n7431 & n7436;
  assign n7438 = pi20  & n7437;
  assign n7439 = ~pi20  & ~n7437;
  assign n7440 = ~n7438 & ~n7439;
  assign n7441 = ~n7430 & ~n7440;
  assign n7442 = ~n7429 & ~n7441;
  assign n7443 = n6987 & ~n7442;
  assign n7444 = ~n6987 & n7442;
  assign n7445 = ~n1107 & n6184;
  assign n7446 = ~n1005 & n6527;
  assign n7447 = n4106 & n6185;
  assign n7448 = ~n894 & n6543;
  assign n7449 = ~n7447 & ~n7448;
  assign n7450 = ~n7446 & n7449;
  assign n7451 = ~n7445 & n7450;
  assign n7452 = pi17  & n7451;
  assign n7453 = ~pi17  & ~n7451;
  assign n7454 = ~n7452 & ~n7453;
  assign n7455 = ~n7444 & ~n7454;
  assign n7456 = ~n7443 & ~n7455;
  assign n7457 = ~n6983 & ~n7456;
  assign n7458 = ~n6980 & ~n7457;
  assign n7459 = ~n3744 & n6836;
  assign n7460 = ~n6830 & n6833;
  assign n7461 = ~n554 & n7460;
  assign n7462 = ~n720 & n6835;
  assign n7463 = ~n7461 & ~n7462;
  assign n7464 = ~n7459 & n7463;
  assign n7465 = pi14  & n7464;
  assign n7466 = ~pi14  & ~n7464;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = ~n7458 & ~n7467;
  assign n7469 = n7458 & n7467;
  assign n7470 = ~n7468 & ~n7469;
  assign n7471 = ~n6943 & ~n6944;
  assign n7472 = ~n6954 & n7471;
  assign n7473 = n6954 & ~n7471;
  assign n7474 = ~n7472 & ~n7473;
  assign n7475 = n7470 & n7474;
  assign n7476 = ~n7468 & ~n7475;
  assign n7477 = ~n6957 & ~n6958;
  assign n7478 = n6962 & n7477;
  assign n7479 = ~n6962 & ~n7477;
  assign n7480 = ~n7478 & ~n7479;
  assign n7481 = ~n7476 & n7480;
  assign n7482 = n7476 & ~n7480;
  assign n7483 = ~n7481 & ~n7482;
  assign n7484 = ~n665 & n6835;
  assign n7485 = ~n720 & n7460;
  assign n7486 = n3979 & n6836;
  assign n7487 = n6827 & ~n6833;
  assign n7488 = ~n554 & n7487;
  assign n7489 = ~n7486 & ~n7488;
  assign n7490 = ~n7485 & n7489;
  assign n7491 = ~n7484 & n7490;
  assign n7492 = pi14  & n7491;
  assign n7493 = ~pi14  & ~n7491;
  assign n7494 = ~n7492 & ~n7493;
  assign n7495 = ~n7443 & ~n7444;
  assign n7496 = ~n7454 & n7495;
  assign n7497 = n7454 & ~n7495;
  assign n7498 = ~n7496 & ~n7497;
  assign n7499 = n7003 & n7422;
  assign n7500 = ~n7423 & ~n7499;
  assign n7501 = ~n1610 & n5435;
  assign n7502 = ~n1531 & n6055;
  assign n7503 = n4724 & n5429;
  assign n7504 = ~n1426 & n6071;
  assign n7505 = ~n7503 & ~n7504;
  assign n7506 = ~n7502 & n7505;
  assign n7507 = ~n7501 & n7506;
  assign n7508 = pi20  & n7507;
  assign n7509 = ~pi20  & ~n7507;
  assign n7510 = ~n7508 & ~n7509;
  assign n7511 = n7500 & ~n7510;
  assign n7512 = ~n7500 & n7510;
  assign n7513 = ~n7511 & ~n7512;
  assign n7514 = ~n7409 & ~n7410;
  assign n7515 = ~n7420 & n7514;
  assign n7516 = n7420 & ~n7514;
  assign n7517 = ~n7515 & ~n7516;
  assign n7518 = ~n2457 & n4601;
  assign n7519 = ~n2369 & n4783;
  assign n7520 = n4602 & n5795;
  assign n7521 = ~n2278 & n4801;
  assign n7522 = ~n7520 & ~n7521;
  assign n7523 = ~n7519 & n7522;
  assign n7524 = ~n7518 & n7523;
  assign n7525 = pi26  & n7524;
  assign n7526 = ~pi26  & ~n7524;
  assign n7527 = ~n7525 & ~n7526;
  assign n7528 = ~n7381 & ~n7382;
  assign n7529 = ~n7392 & n7528;
  assign n7530 = n7392 & ~n7528;
  assign n7531 = ~n7529 & ~n7530;
  assign n7532 = ~n7527 & n7531;
  assign n7533 = n7527 & ~n7531;
  assign n7534 = ~n7532 & ~n7533;
  assign n7535 = ~n2748 & n4006;
  assign n7536 = ~n2676 & n4133;
  assign n7537 = n4002 & n6597;
  assign n7538 = ~n2640 & n4555;
  assign n7539 = ~n7537 & ~n7538;
  assign n7540 = ~n7536 & n7539;
  assign n7541 = ~n7535 & n7540;
  assign n7542 = pi29  & n7541;
  assign n7543 = ~pi29  & ~n7541;
  assign n7544 = ~n7542 & ~n7543;
  assign n7545 = n7371 & n7374;
  assign n7546 = ~n7375 & ~n7545;
  assign n7547 = ~n7544 & n7546;
  assign n7548 = n7544 & ~n7546;
  assign n7549 = ~n2554 & n4601;
  assign n7550 = ~n2457 & n4783;
  assign n7551 = n4602 & n6218;
  assign n7552 = ~n2369 & n4801;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = ~n7550 & n7553;
  assign n7555 = ~n7549 & n7554;
  assign n7556 = pi26  & n7555;
  assign n7557 = ~pi26  & ~n7555;
  assign n7558 = ~n7556 & ~n7557;
  assign n7559 = ~n7548 & ~n7558;
  assign n7560 = ~n7547 & ~n7559;
  assign n7561 = n7534 & ~n7560;
  assign n7562 = ~n7532 & ~n7561;
  assign n7563 = ~n7395 & ~n7396;
  assign n7564 = ~n7406 & n7563;
  assign n7565 = n7406 & ~n7563;
  assign n7566 = ~n7564 & ~n7565;
  assign n7567 = ~n7562 & n7566;
  assign n7568 = n7562 & ~n7566;
  assign n7569 = ~n2058 & n5238;
  assign n7570 = n71 & ~n2006;
  assign n7571 = n5180 & n5239;
  assign n7572 = ~n1900 & n5326;
  assign n7573 = ~n7571 & ~n7572;
  assign n7574 = ~n7570 & n7573;
  assign n7575 = ~n7569 & n7574;
  assign n7576 = pi23  & n7575;
  assign n7577 = ~pi23  & ~n7575;
  assign n7578 = ~n7576 & ~n7577;
  assign n7579 = ~n7568 & ~n7578;
  assign n7580 = ~n7567 & ~n7579;
  assign n7581 = n7517 & ~n7580;
  assign n7582 = ~n7517 & n7580;
  assign n7583 = ~n1740 & n5435;
  assign n7584 = ~n1610 & n6055;
  assign n7585 = n4708 & n5429;
  assign n7586 = ~n1531 & n6071;
  assign n7587 = ~n7585 & ~n7586;
  assign n7588 = ~n7584 & n7587;
  assign n7589 = ~n7583 & n7588;
  assign n7590 = pi20  & n7589;
  assign n7591 = ~pi20  & ~n7589;
  assign n7592 = ~n7590 & ~n7591;
  assign n7593 = ~n7582 & ~n7592;
  assign n7594 = ~n7581 & ~n7593;
  assign n7595 = n7513 & ~n7594;
  assign n7596 = ~n7511 & ~n7595;
  assign n7597 = ~n7429 & ~n7430;
  assign n7598 = ~n7440 & n7597;
  assign n7599 = n7440 & ~n7597;
  assign n7600 = ~n7598 & ~n7599;
  assign n7601 = ~n7596 & n7600;
  assign n7602 = n7596 & ~n7600;
  assign n7603 = ~n1230 & n6184;
  assign n7604 = ~n1107 & n6527;
  assign n7605 = n4307 & n6185;
  assign n7606 = ~n1005 & n6543;
  assign n7607 = ~n7605 & ~n7606;
  assign n7608 = ~n7604 & n7607;
  assign n7609 = ~n7603 & n7608;
  assign n7610 = pi17  & n7609;
  assign n7611 = ~pi17  & ~n7609;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = ~n7602 & ~n7612;
  assign n7614 = ~n7601 & ~n7613;
  assign n7615 = n7498 & ~n7614;
  assign n7616 = ~n7498 & n7614;
  assign n7617 = ~n795 & n6835;
  assign n7618 = ~n665 & n7460;
  assign n7619 = n4015 & n6836;
  assign n7620 = ~n720 & n7487;
  assign n7621 = ~n7619 & ~n7620;
  assign n7622 = ~n7618 & n7621;
  assign n7623 = ~n7617 & n7622;
  assign n7624 = pi14  & n7623;
  assign n7625 = ~pi14  & ~n7623;
  assign n7626 = ~n7624 & ~n7625;
  assign n7627 = ~n7616 & ~n7626;
  assign n7628 = ~n7615 & ~n7627;
  assign n7629 = ~n7494 & ~n7628;
  assign n7630 = n6983 & n7456;
  assign n7631 = ~n7457 & ~n7630;
  assign n7632 = n7494 & ~n7628;
  assign n7633 = ~n7494 & n7628;
  assign n7634 = ~n7632 & ~n7633;
  assign n7635 = n7631 & ~n7634;
  assign n7636 = ~n7629 & ~n7635;
  assign n7637 = ~n7470 & ~n7474;
  assign n7638 = ~n7475 & ~n7637;
  assign n7639 = ~n7636 & n7638;
  assign n7640 = ~n7631 & n7634;
  assign n7641 = ~n7635 & ~n7640;
  assign n7642 = pi8  & ~pi9 ;
  assign n7643 = ~pi8  & pi9 ;
  assign n7644 = ~n7642 & ~n7643;
  assign n7645 = pi10  & ~pi11 ;
  assign n7646 = ~pi10  & pi11 ;
  assign n7647 = ~n7645 & ~n7646;
  assign n7648 = ~n7644 & ~n7647;
  assign n7649 = ~n3638 & n7648;
  assign n7650 = ~pi9  & pi10 ;
  assign n7651 = pi9  & ~pi10 ;
  assign n7652 = ~n7650 & ~n7651;
  assign n7653 = n7644 & n7652;
  assign n7654 = ~n7647 & n7653;
  assign n7655 = ~n7649 & ~n7654;
  assign n7656 = ~n554 & ~n7655;
  assign n7657 = pi11  & ~n7656;
  assign n7658 = ~pi11  & n7656;
  assign n7659 = ~n7657 & ~n7658;
  assign n7660 = ~n1338 & n6184;
  assign n7661 = ~n1230 & n6527;
  assign n7662 = n4323 & n6185;
  assign n7663 = ~n1107 & n6543;
  assign n7664 = ~n7662 & ~n7663;
  assign n7665 = ~n7661 & n7664;
  assign n7666 = ~n7660 & n7665;
  assign n7667 = ~pi17  & ~n7666;
  assign n7668 = pi17  & n7666;
  assign n7669 = ~n7667 & ~n7668;
  assign n7670 = ~n7513 & n7594;
  assign n7671 = ~n7595 & ~n7670;
  assign n7672 = ~n7669 & n7671;
  assign n7673 = ~n7669 & ~n7671;
  assign n7674 = n7669 & n7671;
  assign n7675 = ~n7673 & ~n7674;
  assign n7676 = ~n7581 & ~n7582;
  assign n7677 = ~n7592 & n7676;
  assign n7678 = n7592 & ~n7676;
  assign n7679 = ~n7677 & ~n7678;
  assign n7680 = ~n2178 & n5238;
  assign n7681 = n71 & ~n2058;
  assign n7682 = n5239 & n5554;
  assign n7683 = ~n2006 & n5326;
  assign n7684 = ~n7682 & ~n7683;
  assign n7685 = ~n7681 & n7684;
  assign n7686 = ~n7680 & n7685;
  assign n7687 = ~pi23  & ~n7686;
  assign n7688 = pi23  & n7686;
  assign n7689 = ~n7687 & ~n7688;
  assign n7690 = ~n7534 & n7560;
  assign n7691 = ~n7561 & ~n7690;
  assign n7692 = ~n7689 & n7691;
  assign n7693 = ~n7689 & ~n7691;
  assign n7694 = n7689 & n7691;
  assign n7695 = ~n7693 & ~n7694;
  assign n7696 = ~n7547 & ~n7548;
  assign n7697 = ~n7558 & n7696;
  assign n7698 = n7558 & ~n7696;
  assign n7699 = ~n7697 & ~n7698;
  assign n7700 = ~n2803 & n4006;
  assign n7701 = ~n2748 & n4133;
  assign n7702 = n4002 & n6427;
  assign n7703 = ~n2676 & n4555;
  assign n7704 = ~n7702 & ~n7703;
  assign n7705 = ~n7701 & n7704;
  assign n7706 = ~n7700 & n7705;
  assign n7707 = pi29  & n7706;
  assign n7708 = ~pi29  & ~n7706;
  assign n7709 = ~n7707 & ~n7708;
  assign n7710 = n7366 & n7369;
  assign n7711 = ~n7370 & ~n7710;
  assign n7712 = ~n7709 & n7711;
  assign n7713 = n7709 & ~n7711;
  assign n7714 = ~n2640 & n4601;
  assign n7715 = ~n2554 & n4783;
  assign n7716 = n4602 & n5979;
  assign n7717 = ~n2457 & n4801;
  assign n7718 = ~n7716 & ~n7717;
  assign n7719 = ~n7715 & n7718;
  assign n7720 = ~n7714 & n7719;
  assign n7721 = pi26  & n7720;
  assign n7722 = ~pi26  & ~n7720;
  assign n7723 = ~n7721 & ~n7722;
  assign n7724 = ~n7713 & ~n7723;
  assign n7725 = ~n7712 & ~n7724;
  assign n7726 = n7699 & ~n7725;
  assign n7727 = ~n7699 & n7725;
  assign n7728 = ~n2278 & n5238;
  assign n7729 = n71 & ~n2178;
  assign n7730 = n5239 & n5538;
  assign n7731 = ~n2058 & n5326;
  assign n7732 = ~n7730 & ~n7731;
  assign n7733 = ~n7729 & n7732;
  assign n7734 = ~n7728 & n7733;
  assign n7735 = pi23  & n7734;
  assign n7736 = ~pi23  & ~n7734;
  assign n7737 = ~n7735 & ~n7736;
  assign n7738 = ~n7727 & ~n7737;
  assign n7739 = ~n7726 & ~n7738;
  assign n7740 = ~n7695 & ~n7739;
  assign n7741 = ~n7692 & ~n7740;
  assign n7742 = ~n7567 & ~n7568;
  assign n7743 = ~n7578 & n7742;
  assign n7744 = n7578 & ~n7742;
  assign n7745 = ~n7743 & ~n7744;
  assign n7746 = ~n7741 & n7745;
  assign n7747 = n7741 & ~n7745;
  assign n7748 = ~n1811 & n5435;
  assign n7749 = ~n1740 & n6055;
  assign n7750 = n4951 & n5429;
  assign n7751 = ~n1610 & n6071;
  assign n7752 = ~n7750 & ~n7751;
  assign n7753 = ~n7749 & n7752;
  assign n7754 = ~n7748 & n7753;
  assign n7755 = pi20  & n7754;
  assign n7756 = ~pi20  & ~n7754;
  assign n7757 = ~n7755 & ~n7756;
  assign n7758 = ~n7747 & ~n7757;
  assign n7759 = ~n7746 & ~n7758;
  assign n7760 = n7679 & ~n7759;
  assign n7761 = ~n7679 & n7759;
  assign n7762 = ~n1426 & n6184;
  assign n7763 = ~n1338 & n6527;
  assign n7764 = n4753 & n6185;
  assign n7765 = ~n1230 & n6543;
  assign n7766 = ~n7764 & ~n7765;
  assign n7767 = ~n7763 & n7766;
  assign n7768 = ~n7762 & n7767;
  assign n7769 = pi17  & n7768;
  assign n7770 = ~pi17  & ~n7768;
  assign n7771 = ~n7769 & ~n7770;
  assign n7772 = ~n7761 & ~n7771;
  assign n7773 = ~n7760 & ~n7772;
  assign n7774 = ~n7675 & ~n7773;
  assign n7775 = ~n7672 & ~n7774;
  assign n7776 = ~n7601 & ~n7602;
  assign n7777 = ~n7612 & n7776;
  assign n7778 = n7612 & ~n7776;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = ~n7775 & n7779;
  assign n7781 = n7775 & ~n7779;
  assign n7782 = ~n894 & n6835;
  assign n7783 = ~n795 & n7460;
  assign n7784 = n3959 & n6836;
  assign n7785 = ~n665 & n7487;
  assign n7786 = ~n7784 & ~n7785;
  assign n7787 = ~n7783 & n7786;
  assign n7788 = ~n7782 & n7787;
  assign n7789 = pi14  & n7788;
  assign n7790 = ~pi14  & ~n7788;
  assign n7791 = ~n7789 & ~n7790;
  assign n7792 = ~n7781 & ~n7791;
  assign n7793 = ~n7780 & ~n7792;
  assign n7794 = ~n7659 & ~n7793;
  assign n7795 = n7659 & n7793;
  assign n7796 = ~n7615 & ~n7616;
  assign n7797 = ~n7626 & n7796;
  assign n7798 = n7626 & ~n7796;
  assign n7799 = ~n7797 & ~n7798;
  assign n7800 = ~n7795 & n7799;
  assign n7801 = ~n7794 & ~n7800;
  assign n7802 = n7641 & ~n7801;
  assign n7803 = n7675 & n7773;
  assign n7804 = ~n7774 & ~n7803;
  assign n7805 = ~n1005 & n6835;
  assign n7806 = ~n894 & n7460;
  assign n7807 = n4122 & n6836;
  assign n7808 = ~n795 & n7487;
  assign n7809 = ~n7807 & ~n7808;
  assign n7810 = ~n7806 & n7809;
  assign n7811 = ~n7805 & n7810;
  assign n7812 = pi14  & n7811;
  assign n7813 = ~pi14  & ~n7811;
  assign n7814 = ~n7812 & ~n7813;
  assign n7815 = n7804 & ~n7814;
  assign n7816 = n7804 & n7814;
  assign n7817 = ~n7804 & ~n7814;
  assign n7818 = ~n7816 & ~n7817;
  assign n7819 = ~n7760 & ~n7761;
  assign n7820 = ~n7771 & n7819;
  assign n7821 = n7771 & ~n7819;
  assign n7822 = ~n7820 & ~n7821;
  assign n7823 = n7695 & n7739;
  assign n7824 = ~n7740 & ~n7823;
  assign n7825 = ~n1900 & n5435;
  assign n7826 = ~n1811 & n6055;
  assign n7827 = n4967 & n5429;
  assign n7828 = ~n1740 & n6071;
  assign n7829 = ~n7827 & ~n7828;
  assign n7830 = ~n7826 & n7829;
  assign n7831 = ~n7825 & n7830;
  assign n7832 = pi20  & n7831;
  assign n7833 = ~pi20  & ~n7831;
  assign n7834 = ~n7832 & ~n7833;
  assign n7835 = n7824 & ~n7834;
  assign n7836 = ~n7824 & n7834;
  assign n7837 = ~n7835 & ~n7836;
  assign n7838 = ~n7726 & ~n7727;
  assign n7839 = ~n7737 & n7838;
  assign n7840 = n7737 & ~n7838;
  assign n7841 = ~n7839 & ~n7840;
  assign n7842 = ~n2927 & n4006;
  assign n7843 = ~n2891 & n4133;
  assign n7844 = n4002 & n7014;
  assign n7845 = ~n2803 & n4555;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = ~n7843 & n7846;
  assign n7848 = ~n7842 & n7847;
  assign n7849 = pi29  & n7848;
  assign n7850 = ~pi29  & ~n7848;
  assign n7851 = ~n7849 & ~n7850;
  assign n7852 = n7342 & n7345;
  assign n7853 = ~n7346 & ~n7852;
  assign n7854 = ~n7851 & n7853;
  assign n7855 = ~n3005 & n4006;
  assign n7856 = ~n2927 & n4133;
  assign n7857 = n4002 & n7026;
  assign n7858 = ~n2891 & n4555;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = ~n7856 & n7859;
  assign n7861 = ~n7855 & n7860;
  assign n7862 = pi29  & n7861;
  assign n7863 = ~pi29  & ~n7861;
  assign n7864 = ~n7862 & ~n7863;
  assign n7865 = n7337 & n7340;
  assign n7866 = ~n7341 & ~n7865;
  assign n7867 = ~n7864 & n7866;
  assign n7868 = ~n3097 & n4006;
  assign n7869 = ~n3005 & n4133;
  assign n7870 = n4002 & n6694;
  assign n7871 = ~n2927 & n4555;
  assign n7872 = ~n7870 & ~n7871;
  assign n7873 = ~n7869 & n7872;
  assign n7874 = ~n7868 & n7873;
  assign n7875 = ~pi29  & ~n7874;
  assign n7876 = pi29  & n7874;
  assign n7877 = ~n7875 & ~n7876;
  assign n7878 = n7332 & n7335;
  assign n7879 = ~n7336 & ~n7878;
  assign n7880 = ~n7877 & n7879;
  assign n7881 = ~n7877 & ~n7879;
  assign n7882 = n7877 & n7879;
  assign n7883 = ~n7881 & ~n7882;
  assign n7884 = ~n3166 & n4006;
  assign n7885 = ~n3097 & n4133;
  assign n7886 = n4002 & n7071;
  assign n7887 = ~n3005 & n4555;
  assign n7888 = ~n7886 & ~n7887;
  assign n7889 = ~n7885 & n7888;
  assign n7890 = ~n7884 & n7889;
  assign n7891 = ~pi29  & ~n7890;
  assign n7892 = pi29  & n7890;
  assign n7893 = ~n7891 & ~n7892;
  assign n7894 = n7231 & n7330;
  assign n7895 = ~n7331 & ~n7894;
  assign n7896 = ~n7893 & n7895;
  assign n7897 = ~n7893 & ~n7895;
  assign n7898 = n7893 & n7895;
  assign n7899 = ~n7897 & ~n7898;
  assign n7900 = ~n3226 & n4006;
  assign n7901 = ~n3166 & n4133;
  assign n7902 = n4002 & n7121;
  assign n7903 = ~n3097 & n4555;
  assign n7904 = ~n7902 & ~n7903;
  assign n7905 = ~n7901 & n7904;
  assign n7906 = ~n7900 & n7905;
  assign n7907 = ~pi29  & ~n7906;
  assign n7908 = pi29  & n7906;
  assign n7909 = ~n7907 & ~n7908;
  assign n7910 = ~n7318 & ~n7319;
  assign n7911 = ~n7328 & n7910;
  assign n7912 = n7328 & ~n7910;
  assign n7913 = ~n7911 & ~n7912;
  assign n7914 = ~n7909 & n7913;
  assign n7915 = ~n3263 & n4006;
  assign n7916 = ~n3226 & n4133;
  assign n7917 = n4002 & n7175;
  assign n7918 = ~n3166 & n4555;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = ~n7916 & n7919;
  assign n7921 = ~n7915 & n7920;
  assign n7922 = ~pi29  & ~n7921;
  assign n7923 = pi29  & n7921;
  assign n7924 = ~n7922 & ~n7923;
  assign n7925 = ~n7260 & n7271;
  assign n7926 = n7260 & ~n7271;
  assign n7927 = ~n7925 & ~n7926;
  assign n7928 = ~n7924 & ~n7927;
  assign n7929 = ~n3360 & n4006;
  assign n7930 = ~n3263 & n4133;
  assign n7931 = n4002 & n7221;
  assign n7932 = ~n3226 & n4555;
  assign n7933 = ~n7931 & ~n7932;
  assign n7934 = ~n7930 & n7933;
  assign n7935 = ~n7929 & n7934;
  assign n7936 = ~pi29  & ~n7935;
  assign n7937 = pi29  & n7935;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = ~n3450 & n3740;
  assign n7940 = ~n3506 & n3961;
  assign n7941 = ~n3450 & n3506;
  assign n7942 = ~n7262 & ~n7941;
  assign n7943 = n556 & ~n7942;
  assign n7944 = ~n7940 & ~n7943;
  assign n7945 = ~n7939 & n7944;
  assign n7946 = ~n7938 & ~n7945;
  assign n7947 = ~n7938 & n7945;
  assign n7948 = n7938 & ~n7945;
  assign n7949 = ~n7947 & ~n7948;
  assign n7950 = ~n555 & ~n3450;
  assign n7951 = n4002 & ~n7942;
  assign n7952 = ~n3506 & n4555;
  assign n7953 = ~n3450 & n4133;
  assign n7954 = ~n7952 & ~n7953;
  assign n7955 = ~n7951 & n7954;
  assign n7956 = ~n3450 & ~n3998;
  assign n7957 = pi29  & ~n7956;
  assign n7958 = n7955 & n7957;
  assign n7959 = ~n3450 & n4006;
  assign n7960 = ~n3506 & n4133;
  assign n7961 = n4002 & n7265;
  assign n7962 = ~n3360 & n4555;
  assign n7963 = ~n7961 & ~n7962;
  assign n7964 = ~n7960 & n7963;
  assign n7965 = ~n7959 & n7964;
  assign n7966 = n7958 & n7965;
  assign n7967 = n7950 & n7966;
  assign n7968 = ~n3506 & n4006;
  assign n7969 = ~n3360 & n4133;
  assign n7970 = n4002 & n7323;
  assign n7971 = ~n3263 & n4555;
  assign n7972 = ~n7970 & ~n7971;
  assign n7973 = ~n7969 & n7972;
  assign n7974 = ~n7968 & n7973;
  assign n7975 = ~pi29  & ~n7974;
  assign n7976 = pi29  & n7974;
  assign n7977 = ~n7975 & ~n7976;
  assign n7978 = ~n7950 & n7966;
  assign n7979 = n7950 & ~n7966;
  assign n7980 = ~n7978 & ~n7979;
  assign n7981 = ~n7977 & ~n7980;
  assign n7982 = ~n7967 & ~n7981;
  assign n7983 = ~n7949 & ~n7982;
  assign n7984 = ~n7946 & ~n7983;
  assign n7985 = n7924 & n7927;
  assign n7986 = ~n7928 & ~n7985;
  assign n7987 = ~n7984 & n7986;
  assign n7988 = ~n7928 & ~n7987;
  assign n7989 = n7909 & ~n7913;
  assign n7990 = ~n7914 & ~n7989;
  assign n7991 = ~n7988 & n7990;
  assign n7992 = ~n7914 & ~n7991;
  assign n7993 = ~n7899 & ~n7992;
  assign n7994 = ~n7896 & ~n7993;
  assign n7995 = ~n7883 & ~n7994;
  assign n7996 = ~n7880 & ~n7995;
  assign n7997 = n7864 & ~n7866;
  assign n7998 = ~n7867 & ~n7997;
  assign n7999 = ~n7996 & n7998;
  assign n8000 = ~n7867 & ~n7999;
  assign n8001 = n7851 & ~n7853;
  assign n8002 = ~n7854 & ~n8001;
  assign n8003 = ~n8000 & n8002;
  assign n8004 = ~n7854 & ~n8003;
  assign n8005 = ~n7354 & n7364;
  assign n8006 = ~n7365 & ~n8005;
  assign n8007 = ~n8004 & n8006;
  assign n8008 = ~n2676 & n4601;
  assign n8009 = ~n2640 & n4783;
  assign n8010 = n4602 & n6445;
  assign n8011 = ~n2554 & n4801;
  assign n8012 = ~n8010 & ~n8011;
  assign n8013 = ~n8009 & n8012;
  assign n8014 = ~n8008 & n8013;
  assign n8015 = ~pi26  & ~n8014;
  assign n8016 = pi26  & n8014;
  assign n8017 = ~n8015 & ~n8016;
  assign n8018 = n8004 & ~n8006;
  assign n8019 = ~n8007 & ~n8018;
  assign n8020 = ~n8017 & n8019;
  assign n8021 = ~n8007 & ~n8020;
  assign n8022 = ~n7712 & ~n7713;
  assign n8023 = ~n7723 & n8022;
  assign n8024 = n7723 & ~n8022;
  assign n8025 = ~n8023 & ~n8024;
  assign n8026 = ~n8021 & n8025;
  assign n8027 = n8021 & ~n8025;
  assign n8028 = ~n2369 & n5238;
  assign n8029 = n71 & ~n2278;
  assign n8030 = n5239 & n5779;
  assign n8031 = ~n2178 & n5326;
  assign n8032 = ~n8030 & ~n8031;
  assign n8033 = ~n8029 & n8032;
  assign n8034 = ~n8028 & n8033;
  assign n8035 = pi23  & n8034;
  assign n8036 = ~pi23  & ~n8034;
  assign n8037 = ~n8035 & ~n8036;
  assign n8038 = ~n8027 & ~n8037;
  assign n8039 = ~n8026 & ~n8038;
  assign n8040 = n7841 & ~n8039;
  assign n8041 = ~n7841 & n8039;
  assign n8042 = ~n2006 & n5435;
  assign n8043 = ~n1900 & n6055;
  assign n8044 = n5344 & n5429;
  assign n8045 = ~n1811 & n6071;
  assign n8046 = ~n8044 & ~n8045;
  assign n8047 = ~n8043 & n8046;
  assign n8048 = ~n8042 & n8047;
  assign n8049 = pi20  & n8048;
  assign n8050 = ~pi20  & ~n8048;
  assign n8051 = ~n8049 & ~n8050;
  assign n8052 = ~n8041 & ~n8051;
  assign n8053 = ~n8040 & ~n8052;
  assign n8054 = n7837 & ~n8053;
  assign n8055 = ~n7835 & ~n8054;
  assign n8056 = ~n7746 & ~n7747;
  assign n8057 = ~n7757 & n8056;
  assign n8058 = n7757 & ~n8056;
  assign n8059 = ~n8057 & ~n8058;
  assign n8060 = ~n8055 & n8059;
  assign n8061 = n8055 & ~n8059;
  assign n8062 = ~n1531 & n6184;
  assign n8063 = ~n1426 & n6527;
  assign n8064 = n4533 & n6185;
  assign n8065 = ~n1338 & n6543;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = ~n8063 & n8066;
  assign n8068 = ~n8062 & n8067;
  assign n8069 = pi17  & n8068;
  assign n8070 = ~pi17  & ~n8068;
  assign n8071 = ~n8069 & ~n8070;
  assign n8072 = ~n8061 & ~n8071;
  assign n8073 = ~n8060 & ~n8072;
  assign n8074 = n7822 & ~n8073;
  assign n8075 = ~n7822 & n8073;
  assign n8076 = ~n1107 & n6835;
  assign n8077 = ~n1005 & n7460;
  assign n8078 = n4106 & n6836;
  assign n8079 = ~n894 & n7487;
  assign n8080 = ~n8078 & ~n8079;
  assign n8081 = ~n8077 & n8080;
  assign n8082 = ~n8076 & n8081;
  assign n8083 = pi14  & n8082;
  assign n8084 = ~pi14  & ~n8082;
  assign n8085 = ~n8083 & ~n8084;
  assign n8086 = ~n8075 & ~n8085;
  assign n8087 = ~n8074 & ~n8086;
  assign n8088 = ~n7818 & ~n8087;
  assign n8089 = ~n7815 & ~n8088;
  assign n8090 = ~n3744 & n7648;
  assign n8091 = n7644 & ~n7652;
  assign n8092 = ~n554 & n8091;
  assign n8093 = ~n720 & n7654;
  assign n8094 = ~n8092 & ~n8093;
  assign n8095 = ~n8090 & n8094;
  assign n8096 = pi11  & n8095;
  assign n8097 = ~pi11  & ~n8095;
  assign n8098 = ~n8096 & ~n8097;
  assign n8099 = ~n8089 & ~n8098;
  assign n8100 = n8089 & n8098;
  assign n8101 = ~n8099 & ~n8100;
  assign n8102 = ~n7780 & ~n7781;
  assign n8103 = ~n7791 & n8102;
  assign n8104 = n7791 & ~n8102;
  assign n8105 = ~n8103 & ~n8104;
  assign n8106 = n8101 & n8105;
  assign n8107 = ~n8099 & ~n8106;
  assign n8108 = ~n7794 & ~n7795;
  assign n8109 = n7799 & n8108;
  assign n8110 = ~n7799 & ~n8108;
  assign n8111 = ~n8109 & ~n8110;
  assign n8112 = ~n8107 & n8111;
  assign n8113 = n8107 & ~n8111;
  assign n8114 = ~n8112 & ~n8113;
  assign n8115 = ~n8101 & ~n8105;
  assign n8116 = ~n8106 & ~n8115;
  assign n8117 = ~n665 & n7654;
  assign n8118 = ~n720 & n8091;
  assign n8119 = n3979 & n7648;
  assign n8120 = ~n7644 & n7647;
  assign n8121 = ~n554 & n8120;
  assign n8122 = ~n8119 & ~n8121;
  assign n8123 = ~n8118 & n8122;
  assign n8124 = ~n8117 & n8123;
  assign n8125 = pi11  & n8124;
  assign n8126 = ~pi11  & ~n8124;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = ~n8074 & ~n8075;
  assign n8129 = ~n8085 & n8128;
  assign n8130 = n8085 & ~n8128;
  assign n8131 = ~n8129 & ~n8130;
  assign n8132 = ~n1610 & n6184;
  assign n8133 = ~n1531 & n6527;
  assign n8134 = n4724 & n6185;
  assign n8135 = ~n1426 & n6543;
  assign n8136 = ~n8134 & ~n8135;
  assign n8137 = ~n8133 & n8136;
  assign n8138 = ~n8132 & n8137;
  assign n8139 = ~pi17  & ~n8138;
  assign n8140 = pi17  & n8138;
  assign n8141 = ~n8139 & ~n8140;
  assign n8142 = ~n7837 & n8053;
  assign n8143 = ~n8054 & ~n8142;
  assign n8144 = ~n8141 & n8143;
  assign n8145 = ~n8141 & ~n8143;
  assign n8146 = n8141 & n8143;
  assign n8147 = ~n8145 & ~n8146;
  assign n8148 = ~n8040 & ~n8041;
  assign n8149 = ~n8051 & n8148;
  assign n8150 = n8051 & ~n8148;
  assign n8151 = ~n8149 & ~n8150;
  assign n8152 = n8000 & ~n8002;
  assign n8153 = ~n8003 & ~n8152;
  assign n8154 = ~n2748 & n4601;
  assign n8155 = ~n2676 & n4783;
  assign n8156 = n4602 & n6597;
  assign n8157 = ~n2640 & n4801;
  assign n8158 = ~n8156 & ~n8157;
  assign n8159 = ~n8155 & n8158;
  assign n8160 = ~n8154 & n8159;
  assign n8161 = pi26  & n8160;
  assign n8162 = ~pi26  & ~n8160;
  assign n8163 = ~n8161 & ~n8162;
  assign n8164 = n8153 & ~n8163;
  assign n8165 = n7996 & ~n7998;
  assign n8166 = ~n7999 & ~n8165;
  assign n8167 = ~n2803 & n4601;
  assign n8168 = ~n2748 & n4783;
  assign n8169 = n4602 & n6427;
  assign n8170 = ~n2676 & n4801;
  assign n8171 = ~n8169 & ~n8170;
  assign n8172 = ~n8168 & n8171;
  assign n8173 = ~n8167 & n8172;
  assign n8174 = pi26  & n8173;
  assign n8175 = ~pi26  & ~n8173;
  assign n8176 = ~n8174 & ~n8175;
  assign n8177 = n8166 & ~n8176;
  assign n8178 = n7883 & n7994;
  assign n8179 = ~n7995 & ~n8178;
  assign n8180 = ~n2891 & n4601;
  assign n8181 = ~n2803 & n4783;
  assign n8182 = n4602 & n6715;
  assign n8183 = ~n2748 & n4801;
  assign n8184 = ~n8182 & ~n8183;
  assign n8185 = ~n8181 & n8184;
  assign n8186 = ~n8180 & n8185;
  assign n8187 = pi26  & n8186;
  assign n8188 = ~pi26  & ~n8186;
  assign n8189 = ~n8187 & ~n8188;
  assign n8190 = n8179 & ~n8189;
  assign n8191 = n7899 & n7992;
  assign n8192 = ~n7993 & ~n8191;
  assign n8193 = ~n2927 & n4601;
  assign n8194 = ~n2891 & n4783;
  assign n8195 = n4602 & n7014;
  assign n8196 = ~n2803 & n4801;
  assign n8197 = ~n8195 & ~n8196;
  assign n8198 = ~n8194 & n8197;
  assign n8199 = ~n8193 & n8198;
  assign n8200 = pi26  & n8199;
  assign n8201 = ~pi26  & ~n8199;
  assign n8202 = ~n8200 & ~n8201;
  assign n8203 = n8192 & ~n8202;
  assign n8204 = n7988 & ~n7990;
  assign n8205 = ~n7991 & ~n8204;
  assign n8206 = ~n3005 & n4601;
  assign n8207 = ~n2927 & n4783;
  assign n8208 = n4602 & n7026;
  assign n8209 = ~n2891 & n4801;
  assign n8210 = ~n8208 & ~n8209;
  assign n8211 = ~n8207 & n8210;
  assign n8212 = ~n8206 & n8211;
  assign n8213 = pi26  & n8212;
  assign n8214 = ~pi26  & ~n8212;
  assign n8215 = ~n8213 & ~n8214;
  assign n8216 = n8205 & ~n8215;
  assign n8217 = n7984 & ~n7986;
  assign n8218 = ~n7987 & ~n8217;
  assign n8219 = ~n3097 & n4601;
  assign n8220 = ~n3005 & n4783;
  assign n8221 = n4602 & n6694;
  assign n8222 = ~n2927 & n4801;
  assign n8223 = ~n8221 & ~n8222;
  assign n8224 = ~n8220 & n8223;
  assign n8225 = ~n8219 & n8224;
  assign n8226 = pi26  & n8225;
  assign n8227 = ~pi26  & ~n8225;
  assign n8228 = ~n8226 & ~n8227;
  assign n8229 = n8218 & ~n8228;
  assign n8230 = ~n3166 & n4601;
  assign n8231 = ~n3097 & n4783;
  assign n8232 = n4602 & n7071;
  assign n8233 = ~n3005 & n4801;
  assign n8234 = ~n8232 & ~n8233;
  assign n8235 = ~n8231 & n8234;
  assign n8236 = ~n8230 & n8235;
  assign n8237 = pi26  & n8236;
  assign n8238 = ~pi26  & ~n8236;
  assign n8239 = ~n8237 & ~n8238;
  assign n8240 = n7949 & n7982;
  assign n8241 = ~n7983 & ~n8240;
  assign n8242 = ~n8239 & n8241;
  assign n8243 = ~n3226 & n4601;
  assign n8244 = ~n3166 & n4783;
  assign n8245 = n4602 & n7121;
  assign n8246 = ~n3097 & n4801;
  assign n8247 = ~n8245 & ~n8246;
  assign n8248 = ~n8244 & n8247;
  assign n8249 = ~n8243 & n8248;
  assign n8250 = ~pi26  & ~n8249;
  assign n8251 = pi26  & n8249;
  assign n8252 = ~n8250 & ~n8251;
  assign n8253 = n7977 & n7980;
  assign n8254 = ~n7981 & ~n8253;
  assign n8255 = ~n8252 & n8254;
  assign n8256 = ~n8252 & ~n8254;
  assign n8257 = n8252 & n8254;
  assign n8258 = ~n8256 & ~n8257;
  assign n8259 = ~n3263 & n4601;
  assign n8260 = ~n3226 & n4783;
  assign n8261 = n4602 & n7175;
  assign n8262 = ~n3166 & n4801;
  assign n8263 = ~n8261 & ~n8262;
  assign n8264 = ~n8260 & n8263;
  assign n8265 = ~n8259 & n8264;
  assign n8266 = ~pi26  & ~n8265;
  assign n8267 = pi26  & n8265;
  assign n8268 = ~n8266 & ~n8267;
  assign n8269 = pi29  & ~n7958;
  assign n8270 = n7965 & ~n8269;
  assign n8271 = ~n7965 & n8269;
  assign n8272 = ~n8270 & ~n8271;
  assign n8273 = ~n8268 & n8272;
  assign n8274 = ~n8268 & ~n8272;
  assign n8275 = n8268 & n8272;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = ~n3360 & n4601;
  assign n8278 = ~n3263 & n4783;
  assign n8279 = n4602 & n7221;
  assign n8280 = ~n3226 & n4801;
  assign n8281 = ~n8279 & ~n8280;
  assign n8282 = ~n8278 & n8281;
  assign n8283 = ~n8277 & n8282;
  assign n8284 = pi26  & n8283;
  assign n8285 = ~pi26  & ~n8283;
  assign n8286 = ~n8284 & ~n8285;
  assign n8287 = pi29  & n7956;
  assign n8288 = ~n7955 & n8287;
  assign n8289 = n7955 & ~n8287;
  assign n8290 = ~n8288 & ~n8289;
  assign n8291 = ~n8286 & n8290;
  assign n8292 = n4602 & ~n7942;
  assign n8293 = ~n3506 & n4801;
  assign n8294 = ~n3450 & n4783;
  assign n8295 = ~n8293 & ~n8294;
  assign n8296 = ~n8292 & n8295;
  assign n8297 = ~n3450 & ~n4598;
  assign n8298 = pi26  & ~n8297;
  assign n8299 = n8296 & n8298;
  assign n8300 = ~n3450 & n4601;
  assign n8301 = ~n3506 & n4783;
  assign n8302 = n4602 & n7265;
  assign n8303 = ~n3360 & n4801;
  assign n8304 = ~n8302 & ~n8303;
  assign n8305 = ~n8301 & n8304;
  assign n8306 = ~n8300 & n8305;
  assign n8307 = n8299 & n8306;
  assign n8308 = n7956 & n8307;
  assign n8309 = ~n7956 & n8307;
  assign n8310 = n7956 & ~n8307;
  assign n8311 = ~n8309 & ~n8310;
  assign n8312 = ~n3506 & n4601;
  assign n8313 = ~n3360 & n4783;
  assign n8314 = n4602 & n7323;
  assign n8315 = ~n3263 & n4801;
  assign n8316 = ~n8314 & ~n8315;
  assign n8317 = ~n8313 & n8316;
  assign n8318 = ~n8312 & n8317;
  assign n8319 = pi26  & n8318;
  assign n8320 = ~pi26  & ~n8318;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = ~n8311 & ~n8321;
  assign n8323 = ~n8308 & ~n8322;
  assign n8324 = n8286 & ~n8290;
  assign n8325 = ~n8291 & ~n8324;
  assign n8326 = ~n8323 & n8325;
  assign n8327 = ~n8291 & ~n8326;
  assign n8328 = ~n8276 & ~n8327;
  assign n8329 = ~n8273 & ~n8328;
  assign n8330 = ~n8258 & ~n8329;
  assign n8331 = ~n8255 & ~n8330;
  assign n8332 = n8239 & n8241;
  assign n8333 = ~n8239 & ~n8241;
  assign n8334 = ~n8332 & ~n8333;
  assign n8335 = ~n8331 & ~n8334;
  assign n8336 = ~n8242 & ~n8335;
  assign n8337 = n8218 & n8228;
  assign n8338 = ~n8218 & ~n8228;
  assign n8339 = ~n8337 & ~n8338;
  assign n8340 = ~n8336 & ~n8339;
  assign n8341 = ~n8229 & ~n8340;
  assign n8342 = n8205 & n8215;
  assign n8343 = ~n8205 & ~n8215;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = ~n8341 & ~n8344;
  assign n8346 = ~n8216 & ~n8345;
  assign n8347 = n8192 & n8202;
  assign n8348 = ~n8192 & ~n8202;
  assign n8349 = ~n8347 & ~n8348;
  assign n8350 = ~n8346 & ~n8349;
  assign n8351 = ~n8203 & ~n8350;
  assign n8352 = n8179 & n8189;
  assign n8353 = ~n8179 & ~n8189;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = ~n8351 & ~n8354;
  assign n8356 = ~n8190 & ~n8355;
  assign n8357 = n8166 & n8176;
  assign n8358 = ~n8166 & ~n8176;
  assign n8359 = ~n8357 & ~n8358;
  assign n8360 = ~n8356 & ~n8359;
  assign n8361 = ~n8177 & ~n8360;
  assign n8362 = n8153 & n8163;
  assign n8363 = ~n8153 & ~n8163;
  assign n8364 = ~n8362 & ~n8363;
  assign n8365 = ~n8361 & ~n8364;
  assign n8366 = ~n8164 & ~n8365;
  assign n8367 = n8017 & ~n8019;
  assign n8368 = ~n8020 & ~n8367;
  assign n8369 = ~n8366 & n8368;
  assign n8370 = ~n2457 & n5238;
  assign n8371 = n71 & ~n2369;
  assign n8372 = n5239 & n5795;
  assign n8373 = ~n2278 & n5326;
  assign n8374 = ~n8372 & ~n8373;
  assign n8375 = ~n8371 & n8374;
  assign n8376 = ~n8370 & n8375;
  assign n8377 = ~pi23  & ~n8376;
  assign n8378 = pi23  & n8376;
  assign n8379 = ~n8377 & ~n8378;
  assign n8380 = n8366 & ~n8368;
  assign n8381 = ~n8369 & ~n8380;
  assign n8382 = ~n8379 & n8381;
  assign n8383 = ~n8369 & ~n8382;
  assign n8384 = ~n8026 & ~n8027;
  assign n8385 = ~n8037 & n8384;
  assign n8386 = n8037 & ~n8384;
  assign n8387 = ~n8385 & ~n8386;
  assign n8388 = ~n8383 & n8387;
  assign n8389 = n8383 & ~n8387;
  assign n8390 = ~n2058 & n5435;
  assign n8391 = ~n2006 & n6055;
  assign n8392 = n5180 & n5429;
  assign n8393 = ~n1900 & n6071;
  assign n8394 = ~n8392 & ~n8393;
  assign n8395 = ~n8391 & n8394;
  assign n8396 = ~n8390 & n8395;
  assign n8397 = pi20  & n8396;
  assign n8398 = ~pi20  & ~n8396;
  assign n8399 = ~n8397 & ~n8398;
  assign n8400 = ~n8389 & ~n8399;
  assign n8401 = ~n8388 & ~n8400;
  assign n8402 = n8151 & ~n8401;
  assign n8403 = ~n8151 & n8401;
  assign n8404 = ~n1740 & n6184;
  assign n8405 = ~n1610 & n6527;
  assign n8406 = n4708 & n6185;
  assign n8407 = ~n1531 & n6543;
  assign n8408 = ~n8406 & ~n8407;
  assign n8409 = ~n8405 & n8408;
  assign n8410 = ~n8404 & n8409;
  assign n8411 = pi17  & n8410;
  assign n8412 = ~pi17  & ~n8410;
  assign n8413 = ~n8411 & ~n8412;
  assign n8414 = ~n8403 & ~n8413;
  assign n8415 = ~n8402 & ~n8414;
  assign n8416 = ~n8147 & ~n8415;
  assign n8417 = ~n8144 & ~n8416;
  assign n8418 = ~n8060 & ~n8061;
  assign n8419 = ~n8071 & n8418;
  assign n8420 = n8071 & ~n8418;
  assign n8421 = ~n8419 & ~n8420;
  assign n8422 = ~n8417 & n8421;
  assign n8423 = n8417 & ~n8421;
  assign n8424 = ~n1230 & n6835;
  assign n8425 = ~n1107 & n7460;
  assign n8426 = n4307 & n6836;
  assign n8427 = ~n1005 & n7487;
  assign n8428 = ~n8426 & ~n8427;
  assign n8429 = ~n8425 & n8428;
  assign n8430 = ~n8424 & n8429;
  assign n8431 = pi14  & n8430;
  assign n8432 = ~pi14  & ~n8430;
  assign n8433 = ~n8431 & ~n8432;
  assign n8434 = ~n8423 & ~n8433;
  assign n8435 = ~n8422 & ~n8434;
  assign n8436 = n8131 & ~n8435;
  assign n8437 = ~n8131 & n8435;
  assign n8438 = ~n795 & n7654;
  assign n8439 = ~n665 & n8091;
  assign n8440 = n4015 & n7648;
  assign n8441 = ~n720 & n8120;
  assign n8442 = ~n8440 & ~n8441;
  assign n8443 = ~n8439 & n8442;
  assign n8444 = ~n8438 & n8443;
  assign n8445 = pi11  & n8444;
  assign n8446 = ~pi11  & ~n8444;
  assign n8447 = ~n8445 & ~n8446;
  assign n8448 = ~n8437 & ~n8447;
  assign n8449 = ~n8436 & ~n8448;
  assign n8450 = ~n8127 & ~n8449;
  assign n8451 = n8127 & n8449;
  assign n8452 = n7818 & ~n8087;
  assign n8453 = ~n7818 & n8087;
  assign n8454 = ~n8452 & ~n8453;
  assign n8455 = ~n8451 & ~n8454;
  assign n8456 = ~n8450 & ~n8455;
  assign n8457 = n8116 & ~n8456;
  assign n8458 = ~n8450 & ~n8451;
  assign n8459 = ~n8454 & n8458;
  assign n8460 = n8454 & ~n8458;
  assign n8461 = ~n8459 & ~n8460;
  assign n8462 = pi5  & ~pi6 ;
  assign n8463 = ~pi5  & pi6 ;
  assign n8464 = ~n8462 & ~n8463;
  assign n8465 = pi7  & ~pi8 ;
  assign n8466 = ~pi7  & pi8 ;
  assign n8467 = ~n8465 & ~n8466;
  assign n8468 = ~n8464 & ~n8467;
  assign n8469 = ~n3638 & n8468;
  assign n8470 = ~pi6  & pi7 ;
  assign n8471 = pi6  & ~pi7 ;
  assign n8472 = ~n8470 & ~n8471;
  assign n8473 = n8464 & n8472;
  assign n8474 = ~n8467 & n8473;
  assign n8475 = ~n8469 & ~n8474;
  assign n8476 = ~n554 & ~n8475;
  assign n8477 = pi8  & ~n8476;
  assign n8478 = ~pi8  & n8476;
  assign n8479 = ~n8477 & ~n8478;
  assign n8480 = n8147 & n8415;
  assign n8481 = ~n8416 & ~n8480;
  assign n8482 = ~n1338 & n6835;
  assign n8483 = ~n1230 & n7460;
  assign n8484 = n4323 & n6836;
  assign n8485 = ~n1107 & n7487;
  assign n8486 = ~n8484 & ~n8485;
  assign n8487 = ~n8483 & n8486;
  assign n8488 = ~n8482 & n8487;
  assign n8489 = pi14  & n8488;
  assign n8490 = ~pi14  & ~n8488;
  assign n8491 = ~n8489 & ~n8490;
  assign n8492 = n8481 & ~n8491;
  assign n8493 = ~n8481 & n8491;
  assign n8494 = ~n8492 & ~n8493;
  assign n8495 = ~n8402 & ~n8403;
  assign n8496 = ~n8413 & n8495;
  assign n8497 = n8413 & ~n8495;
  assign n8498 = ~n8496 & ~n8497;
  assign n8499 = ~n2554 & n5238;
  assign n8500 = n71 & ~n2457;
  assign n8501 = n5239 & n6218;
  assign n8502 = ~n2369 & n5326;
  assign n8503 = ~n8501 & ~n8502;
  assign n8504 = ~n8500 & n8503;
  assign n8505 = ~n8499 & n8504;
  assign n8506 = ~pi23  & ~n8505;
  assign n8507 = pi23  & n8505;
  assign n8508 = ~n8506 & ~n8507;
  assign n8509 = n8361 & n8364;
  assign n8510 = ~n8365 & ~n8509;
  assign n8511 = ~n8508 & n8510;
  assign n8512 = ~n8508 & ~n8510;
  assign n8513 = n8508 & n8510;
  assign n8514 = ~n8512 & ~n8513;
  assign n8515 = ~n2640 & n5238;
  assign n8516 = n71 & ~n2554;
  assign n8517 = n5239 & n5979;
  assign n8518 = ~n2457 & n5326;
  assign n8519 = ~n8517 & ~n8518;
  assign n8520 = ~n8516 & n8519;
  assign n8521 = ~n8515 & n8520;
  assign n8522 = ~pi23  & ~n8521;
  assign n8523 = pi23  & n8521;
  assign n8524 = ~n8522 & ~n8523;
  assign n8525 = n8356 & n8359;
  assign n8526 = ~n8360 & ~n8525;
  assign n8527 = ~n8524 & n8526;
  assign n8528 = ~n8524 & ~n8526;
  assign n8529 = n8524 & n8526;
  assign n8530 = ~n8528 & ~n8529;
  assign n8531 = ~n2676 & n5238;
  assign n8532 = n71 & ~n2640;
  assign n8533 = n5239 & n6445;
  assign n8534 = ~n2554 & n5326;
  assign n8535 = ~n8533 & ~n8534;
  assign n8536 = ~n8532 & n8535;
  assign n8537 = ~n8531 & n8536;
  assign n8538 = ~pi23  & ~n8537;
  assign n8539 = pi23  & n8537;
  assign n8540 = ~n8538 & ~n8539;
  assign n8541 = ~n8351 & n8354;
  assign n8542 = n8351 & ~n8354;
  assign n8543 = ~n8541 & ~n8542;
  assign n8544 = ~n8540 & ~n8543;
  assign n8545 = ~n2748 & n5238;
  assign n8546 = n71 & ~n2676;
  assign n8547 = n5239 & n6597;
  assign n8548 = ~n2640 & n5326;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = ~n8546 & n8549;
  assign n8551 = ~n8545 & n8550;
  assign n8552 = ~pi23  & ~n8551;
  assign n8553 = pi23  & n8551;
  assign n8554 = ~n8552 & ~n8553;
  assign n8555 = ~n8346 & n8349;
  assign n8556 = n8346 & ~n8349;
  assign n8557 = ~n8555 & ~n8556;
  assign n8558 = ~n8554 & ~n8557;
  assign n8559 = ~n2803 & n5238;
  assign n8560 = n71 & ~n2748;
  assign n8561 = n5239 & n6427;
  assign n8562 = ~n2676 & n5326;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = ~n8560 & n8563;
  assign n8565 = ~n8559 & n8564;
  assign n8566 = ~pi23  & ~n8565;
  assign n8567 = pi23  & n8565;
  assign n8568 = ~n8566 & ~n8567;
  assign n8569 = n8341 & n8344;
  assign n8570 = ~n8345 & ~n8569;
  assign n8571 = ~n8568 & n8570;
  assign n8572 = ~n8568 & ~n8570;
  assign n8573 = n8568 & n8570;
  assign n8574 = ~n8572 & ~n8573;
  assign n8575 = ~n2891 & n5238;
  assign n8576 = n71 & ~n2803;
  assign n8577 = n5239 & n6715;
  assign n8578 = ~n2748 & n5326;
  assign n8579 = ~n8577 & ~n8578;
  assign n8580 = ~n8576 & n8579;
  assign n8581 = ~n8575 & n8580;
  assign n8582 = ~pi23  & ~n8581;
  assign n8583 = pi23  & n8581;
  assign n8584 = ~n8582 & ~n8583;
  assign n8585 = n8336 & n8339;
  assign n8586 = ~n8340 & ~n8585;
  assign n8587 = ~n8584 & n8586;
  assign n8588 = ~n8584 & ~n8586;
  assign n8589 = n8584 & n8586;
  assign n8590 = ~n8588 & ~n8589;
  assign n8591 = ~n2927 & n5238;
  assign n8592 = n71 & ~n2891;
  assign n8593 = n5239 & n7014;
  assign n8594 = ~n2803 & n5326;
  assign n8595 = ~n8593 & ~n8594;
  assign n8596 = ~n8592 & n8595;
  assign n8597 = ~n8591 & n8596;
  assign n8598 = ~pi23  & ~n8597;
  assign n8599 = pi23  & n8597;
  assign n8600 = ~n8598 & ~n8599;
  assign n8601 = ~n8331 & n8334;
  assign n8602 = n8331 & ~n8334;
  assign n8603 = ~n8601 & ~n8602;
  assign n8604 = ~n8600 & ~n8603;
  assign n8605 = n8258 & n8329;
  assign n8606 = ~n8330 & ~n8605;
  assign n8607 = ~n3005 & n5238;
  assign n8608 = n71 & ~n2927;
  assign n8609 = n5239 & n7026;
  assign n8610 = ~n2891 & n5326;
  assign n8611 = ~n8609 & ~n8610;
  assign n8612 = ~n8608 & n8611;
  assign n8613 = ~n8607 & n8612;
  assign n8614 = pi23  & n8613;
  assign n8615 = ~pi23  & ~n8613;
  assign n8616 = ~n8614 & ~n8615;
  assign n8617 = n8606 & ~n8616;
  assign n8618 = n8276 & n8327;
  assign n8619 = ~n8328 & ~n8618;
  assign n8620 = ~n3097 & n5238;
  assign n8621 = n71 & ~n3005;
  assign n8622 = n5239 & n6694;
  assign n8623 = ~n2927 & n5326;
  assign n8624 = ~n8622 & ~n8623;
  assign n8625 = ~n8621 & n8624;
  assign n8626 = ~n8620 & n8625;
  assign n8627 = pi23  & n8626;
  assign n8628 = ~pi23  & ~n8626;
  assign n8629 = ~n8627 & ~n8628;
  assign n8630 = n8619 & ~n8629;
  assign n8631 = ~n3166 & n5238;
  assign n8632 = n71 & ~n3097;
  assign n8633 = n5239 & n7071;
  assign n8634 = ~n3005 & n5326;
  assign n8635 = ~n8633 & ~n8634;
  assign n8636 = ~n8632 & n8635;
  assign n8637 = ~n8631 & n8636;
  assign n8638 = ~pi23  & ~n8637;
  assign n8639 = pi23  & n8637;
  assign n8640 = ~n8638 & ~n8639;
  assign n8641 = n8323 & ~n8325;
  assign n8642 = ~n8326 & ~n8641;
  assign n8643 = ~n8640 & n8642;
  assign n8644 = ~n8640 & ~n8642;
  assign n8645 = n8640 & n8642;
  assign n8646 = ~n8644 & ~n8645;
  assign n8647 = ~n3226 & n5238;
  assign n8648 = n71 & ~n3166;
  assign n8649 = n5239 & n7121;
  assign n8650 = ~n3097 & n5326;
  assign n8651 = ~n8649 & ~n8650;
  assign n8652 = ~n8648 & n8651;
  assign n8653 = ~n8647 & n8652;
  assign n8654 = pi23  & n8653;
  assign n8655 = ~pi23  & ~n8653;
  assign n8656 = ~n8654 & ~n8655;
  assign n8657 = n8311 & n8321;
  assign n8658 = ~n8322 & ~n8657;
  assign n8659 = ~n8656 & n8658;
  assign n8660 = ~n3263 & n5238;
  assign n8661 = n71 & ~n3226;
  assign n8662 = n5239 & n7175;
  assign n8663 = ~n3166 & n5326;
  assign n8664 = ~n8662 & ~n8663;
  assign n8665 = ~n8661 & n8664;
  assign n8666 = ~n8660 & n8665;
  assign n8667 = ~pi23  & ~n8666;
  assign n8668 = pi23  & n8666;
  assign n8669 = ~n8667 & ~n8668;
  assign n8670 = pi26  & ~n8299;
  assign n8671 = n8306 & ~n8670;
  assign n8672 = ~n8306 & n8670;
  assign n8673 = ~n8671 & ~n8672;
  assign n8674 = ~n8669 & n8673;
  assign n8675 = ~n8669 & ~n8673;
  assign n8676 = n8669 & n8673;
  assign n8677 = ~n8675 & ~n8676;
  assign n8678 = ~n3360 & n5238;
  assign n8679 = n71 & ~n3263;
  assign n8680 = n5239 & n7221;
  assign n8681 = ~n3226 & n5326;
  assign n8682 = ~n8680 & ~n8681;
  assign n8683 = ~n8679 & n8682;
  assign n8684 = ~n8678 & n8683;
  assign n8685 = pi23  & n8684;
  assign n8686 = ~pi23  & ~n8684;
  assign n8687 = ~n8685 & ~n8686;
  assign n8688 = pi26  & n8297;
  assign n8689 = ~n8296 & n8688;
  assign n8690 = n8296 & ~n8688;
  assign n8691 = ~n8689 & ~n8690;
  assign n8692 = ~n8687 & n8691;
  assign n8693 = n5239 & ~n7942;
  assign n8694 = ~n3506 & n5326;
  assign n8695 = n71 & ~n3450;
  assign n8696 = ~n8694 & ~n8695;
  assign n8697 = ~n8693 & n8696;
  assign n8698 = ~n70 & ~n3450;
  assign n8699 = pi23  & ~n8698;
  assign n8700 = n8697 & n8699;
  assign n8701 = ~n3450 & n5238;
  assign n8702 = n71 & ~n3506;
  assign n8703 = n5239 & n7265;
  assign n8704 = ~n3360 & n5326;
  assign n8705 = ~n8703 & ~n8704;
  assign n8706 = ~n8702 & n8705;
  assign n8707 = ~n8701 & n8706;
  assign n8708 = n8700 & n8707;
  assign n8709 = n8297 & n8708;
  assign n8710 = ~n8297 & n8708;
  assign n8711 = n8297 & ~n8708;
  assign n8712 = ~n8710 & ~n8711;
  assign n8713 = ~n3506 & n5238;
  assign n8714 = n71 & ~n3360;
  assign n8715 = n5239 & n7323;
  assign n8716 = ~n3263 & n5326;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = ~n8714 & n8717;
  assign n8719 = ~n8713 & n8718;
  assign n8720 = pi23  & n8719;
  assign n8721 = ~pi23  & ~n8719;
  assign n8722 = ~n8720 & ~n8721;
  assign n8723 = ~n8712 & ~n8722;
  assign n8724 = ~n8709 & ~n8723;
  assign n8725 = n8687 & ~n8691;
  assign n8726 = ~n8692 & ~n8725;
  assign n8727 = ~n8724 & n8726;
  assign n8728 = ~n8692 & ~n8727;
  assign n8729 = ~n8677 & ~n8728;
  assign n8730 = ~n8674 & ~n8729;
  assign n8731 = n8656 & ~n8658;
  assign n8732 = ~n8659 & ~n8731;
  assign n8733 = ~n8730 & n8732;
  assign n8734 = ~n8659 & ~n8733;
  assign n8735 = ~n8646 & ~n8734;
  assign n8736 = ~n8643 & ~n8735;
  assign n8737 = n8619 & n8629;
  assign n8738 = ~n8619 & ~n8629;
  assign n8739 = ~n8737 & ~n8738;
  assign n8740 = ~n8736 & ~n8739;
  assign n8741 = ~n8630 & ~n8740;
  assign n8742 = ~n8606 & n8616;
  assign n8743 = ~n8617 & ~n8742;
  assign n8744 = ~n8741 & n8743;
  assign n8745 = ~n8617 & ~n8744;
  assign n8746 = n8600 & n8603;
  assign n8747 = ~n8604 & ~n8746;
  assign n8748 = ~n8745 & n8747;
  assign n8749 = ~n8604 & ~n8748;
  assign n8750 = ~n8590 & ~n8749;
  assign n8751 = ~n8587 & ~n8750;
  assign n8752 = ~n8574 & ~n8751;
  assign n8753 = ~n8571 & ~n8752;
  assign n8754 = n8554 & n8557;
  assign n8755 = ~n8558 & ~n8754;
  assign n8756 = ~n8753 & n8755;
  assign n8757 = ~n8558 & ~n8756;
  assign n8758 = n8540 & n8543;
  assign n8759 = ~n8544 & ~n8758;
  assign n8760 = ~n8757 & n8759;
  assign n8761 = ~n8544 & ~n8760;
  assign n8762 = ~n8530 & ~n8761;
  assign n8763 = ~n8527 & ~n8762;
  assign n8764 = ~n8514 & ~n8763;
  assign n8765 = ~n8511 & ~n8764;
  assign n8766 = n8379 & ~n8381;
  assign n8767 = ~n8382 & ~n8766;
  assign n8768 = ~n8765 & n8767;
  assign n8769 = ~n2178 & n5435;
  assign n8770 = ~n2058 & n6055;
  assign n8771 = n5429 & n5554;
  assign n8772 = ~n2006 & n6071;
  assign n8773 = ~n8771 & ~n8772;
  assign n8774 = ~n8770 & n8773;
  assign n8775 = ~n8769 & n8774;
  assign n8776 = ~pi20  & ~n8775;
  assign n8777 = pi20  & n8775;
  assign n8778 = ~n8776 & ~n8777;
  assign n8779 = n8765 & ~n8767;
  assign n8780 = ~n8768 & ~n8779;
  assign n8781 = ~n8778 & n8780;
  assign n8782 = ~n8768 & ~n8781;
  assign n8783 = ~n8388 & ~n8389;
  assign n8784 = ~n8399 & n8783;
  assign n8785 = n8399 & ~n8783;
  assign n8786 = ~n8784 & ~n8785;
  assign n8787 = ~n8782 & n8786;
  assign n8788 = n8782 & ~n8786;
  assign n8789 = ~n1811 & n6184;
  assign n8790 = ~n1740 & n6527;
  assign n8791 = n4951 & n6185;
  assign n8792 = ~n1610 & n6543;
  assign n8793 = ~n8791 & ~n8792;
  assign n8794 = ~n8790 & n8793;
  assign n8795 = ~n8789 & n8794;
  assign n8796 = pi17  & n8795;
  assign n8797 = ~pi17  & ~n8795;
  assign n8798 = ~n8796 & ~n8797;
  assign n8799 = ~n8788 & ~n8798;
  assign n8800 = ~n8787 & ~n8799;
  assign n8801 = n8498 & ~n8800;
  assign n8802 = ~n8498 & n8800;
  assign n8803 = ~n1426 & n6835;
  assign n8804 = ~n1338 & n7460;
  assign n8805 = n4753 & n6836;
  assign n8806 = ~n1230 & n7487;
  assign n8807 = ~n8805 & ~n8806;
  assign n8808 = ~n8804 & n8807;
  assign n8809 = ~n8803 & n8808;
  assign n8810 = pi14  & n8809;
  assign n8811 = ~pi14  & ~n8809;
  assign n8812 = ~n8810 & ~n8811;
  assign n8813 = ~n8802 & ~n8812;
  assign n8814 = ~n8801 & ~n8813;
  assign n8815 = n8494 & ~n8814;
  assign n8816 = ~n8492 & ~n8815;
  assign n8817 = ~n8422 & ~n8423;
  assign n8818 = ~n8433 & n8817;
  assign n8819 = n8433 & ~n8817;
  assign n8820 = ~n8818 & ~n8819;
  assign n8821 = ~n8816 & n8820;
  assign n8822 = n8816 & ~n8820;
  assign n8823 = ~n894 & n7654;
  assign n8824 = ~n795 & n8091;
  assign n8825 = n3959 & n7648;
  assign n8826 = ~n665 & n8120;
  assign n8827 = ~n8825 & ~n8826;
  assign n8828 = ~n8824 & n8827;
  assign n8829 = ~n8823 & n8828;
  assign n8830 = pi11  & n8829;
  assign n8831 = ~pi11  & ~n8829;
  assign n8832 = ~n8830 & ~n8831;
  assign n8833 = ~n8822 & ~n8832;
  assign n8834 = ~n8821 & ~n8833;
  assign n8835 = ~n8479 & ~n8834;
  assign n8836 = n8479 & n8834;
  assign n8837 = ~n8436 & ~n8437;
  assign n8838 = ~n8447 & n8837;
  assign n8839 = n8447 & ~n8837;
  assign n8840 = ~n8838 & ~n8839;
  assign n8841 = ~n8836 & n8840;
  assign n8842 = ~n8835 & ~n8841;
  assign n8843 = n8461 & ~n8842;
  assign n8844 = ~n8461 & n8842;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = ~n1005 & n7654;
  assign n8847 = ~n894 & n8091;
  assign n8848 = n4122 & n7648;
  assign n8849 = ~n795 & n8120;
  assign n8850 = ~n8848 & ~n8849;
  assign n8851 = ~n8847 & n8850;
  assign n8852 = ~n8846 & n8851;
  assign n8853 = pi11  & n8852;
  assign n8854 = ~pi11  & ~n8852;
  assign n8855 = ~n8853 & ~n8854;
  assign n8856 = ~n8801 & ~n8802;
  assign n8857 = ~n8812 & n8856;
  assign n8858 = n8812 & ~n8856;
  assign n8859 = ~n8857 & ~n8858;
  assign n8860 = n8514 & n8763;
  assign n8861 = ~n8764 & ~n8860;
  assign n8862 = ~n2278 & n5435;
  assign n8863 = ~n2178 & n6055;
  assign n8864 = n5429 & n5538;
  assign n8865 = ~n2058 & n6071;
  assign n8866 = ~n8864 & ~n8865;
  assign n8867 = ~n8863 & n8866;
  assign n8868 = ~n8862 & n8867;
  assign n8869 = pi20  & n8868;
  assign n8870 = ~pi20  & ~n8868;
  assign n8871 = ~n8869 & ~n8870;
  assign n8872 = n8861 & ~n8871;
  assign n8873 = n8530 & n8761;
  assign n8874 = ~n8762 & ~n8873;
  assign n8875 = ~n2369 & n5435;
  assign n8876 = ~n2278 & n6055;
  assign n8877 = n5429 & n5779;
  assign n8878 = ~n2178 & n6071;
  assign n8879 = ~n8877 & ~n8878;
  assign n8880 = ~n8876 & n8879;
  assign n8881 = ~n8875 & n8880;
  assign n8882 = pi20  & n8881;
  assign n8883 = ~pi20  & ~n8881;
  assign n8884 = ~n8882 & ~n8883;
  assign n8885 = n8874 & ~n8884;
  assign n8886 = n8757 & ~n8759;
  assign n8887 = ~n8760 & ~n8886;
  assign n8888 = ~n2457 & n5435;
  assign n8889 = ~n2369 & n6055;
  assign n8890 = n5429 & n5795;
  assign n8891 = ~n2278 & n6071;
  assign n8892 = ~n8890 & ~n8891;
  assign n8893 = ~n8889 & n8892;
  assign n8894 = ~n8888 & n8893;
  assign n8895 = pi20  & n8894;
  assign n8896 = ~pi20  & ~n8894;
  assign n8897 = ~n8895 & ~n8896;
  assign n8898 = n8887 & ~n8897;
  assign n8899 = n8753 & ~n8755;
  assign n8900 = ~n8756 & ~n8899;
  assign n8901 = ~n2554 & n5435;
  assign n8902 = ~n2457 & n6055;
  assign n8903 = n5429 & n6218;
  assign n8904 = ~n2369 & n6071;
  assign n8905 = ~n8903 & ~n8904;
  assign n8906 = ~n8902 & n8905;
  assign n8907 = ~n8901 & n8906;
  assign n8908 = pi20  & n8907;
  assign n8909 = ~pi20  & ~n8907;
  assign n8910 = ~n8908 & ~n8909;
  assign n8911 = n8900 & ~n8910;
  assign n8912 = n8574 & n8751;
  assign n8913 = ~n8752 & ~n8912;
  assign n8914 = ~n2640 & n5435;
  assign n8915 = ~n2554 & n6055;
  assign n8916 = n5429 & n5979;
  assign n8917 = ~n2457 & n6071;
  assign n8918 = ~n8916 & ~n8917;
  assign n8919 = ~n8915 & n8918;
  assign n8920 = ~n8914 & n8919;
  assign n8921 = pi20  & n8920;
  assign n8922 = ~pi20  & ~n8920;
  assign n8923 = ~n8921 & ~n8922;
  assign n8924 = n8913 & ~n8923;
  assign n8925 = n8590 & n8749;
  assign n8926 = ~n8750 & ~n8925;
  assign n8927 = ~n2676 & n5435;
  assign n8928 = ~n2640 & n6055;
  assign n8929 = n5429 & n6445;
  assign n8930 = ~n2554 & n6071;
  assign n8931 = ~n8929 & ~n8930;
  assign n8932 = ~n8928 & n8931;
  assign n8933 = ~n8927 & n8932;
  assign n8934 = pi20  & n8933;
  assign n8935 = ~pi20  & ~n8933;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = n8926 & ~n8936;
  assign n8938 = n8745 & ~n8747;
  assign n8939 = ~n8748 & ~n8938;
  assign n8940 = ~n2748 & n5435;
  assign n8941 = ~n2676 & n6055;
  assign n8942 = n5429 & n6597;
  assign n8943 = ~n2640 & n6071;
  assign n8944 = ~n8942 & ~n8943;
  assign n8945 = ~n8941 & n8944;
  assign n8946 = ~n8940 & n8945;
  assign n8947 = pi20  & n8946;
  assign n8948 = ~pi20  & ~n8946;
  assign n8949 = ~n8947 & ~n8948;
  assign n8950 = n8939 & ~n8949;
  assign n8951 = ~n2803 & n5435;
  assign n8952 = ~n2748 & n6055;
  assign n8953 = n5429 & n6427;
  assign n8954 = ~n2676 & n6071;
  assign n8955 = ~n8953 & ~n8954;
  assign n8956 = ~n8952 & n8955;
  assign n8957 = ~n8951 & n8956;
  assign n8958 = ~pi20  & ~n8957;
  assign n8959 = pi20  & n8957;
  assign n8960 = ~n8958 & ~n8959;
  assign n8961 = n8741 & ~n8743;
  assign n8962 = ~n8744 & ~n8961;
  assign n8963 = ~n8960 & n8962;
  assign n8964 = ~n8960 & ~n8962;
  assign n8965 = n8960 & n8962;
  assign n8966 = ~n8964 & ~n8965;
  assign n8967 = ~n2891 & n5435;
  assign n8968 = ~n2803 & n6055;
  assign n8969 = n5429 & n6715;
  assign n8970 = ~n2748 & n6071;
  assign n8971 = ~n8969 & ~n8970;
  assign n8972 = ~n8968 & n8971;
  assign n8973 = ~n8967 & n8972;
  assign n8974 = ~pi20  & ~n8973;
  assign n8975 = pi20  & n8973;
  assign n8976 = ~n8974 & ~n8975;
  assign n8977 = ~n8736 & n8739;
  assign n8978 = n8736 & ~n8739;
  assign n8979 = ~n8977 & ~n8978;
  assign n8980 = ~n8976 & ~n8979;
  assign n8981 = n8646 & n8734;
  assign n8982 = ~n8735 & ~n8981;
  assign n8983 = ~n2927 & n5435;
  assign n8984 = ~n2891 & n6055;
  assign n8985 = n5429 & n7014;
  assign n8986 = ~n2803 & n6071;
  assign n8987 = ~n8985 & ~n8986;
  assign n8988 = ~n8984 & n8987;
  assign n8989 = ~n8983 & n8988;
  assign n8990 = pi20  & n8989;
  assign n8991 = ~pi20  & ~n8989;
  assign n8992 = ~n8990 & ~n8991;
  assign n8993 = n8982 & ~n8992;
  assign n8994 = n8730 & ~n8732;
  assign n8995 = ~n8733 & ~n8994;
  assign n8996 = ~n3005 & n5435;
  assign n8997 = ~n2927 & n6055;
  assign n8998 = n5429 & n7026;
  assign n8999 = ~n2891 & n6071;
  assign n9000 = ~n8998 & ~n8999;
  assign n9001 = ~n8997 & n9000;
  assign n9002 = ~n8996 & n9001;
  assign n9003 = pi20  & n9002;
  assign n9004 = ~pi20  & ~n9002;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = n8995 & ~n9005;
  assign n9007 = n8677 & n8728;
  assign n9008 = ~n8729 & ~n9007;
  assign n9009 = ~n3097 & n5435;
  assign n9010 = ~n3005 & n6055;
  assign n9011 = n5429 & n6694;
  assign n9012 = ~n2927 & n6071;
  assign n9013 = ~n9011 & ~n9012;
  assign n9014 = ~n9010 & n9013;
  assign n9015 = ~n9009 & n9014;
  assign n9016 = pi20  & n9015;
  assign n9017 = ~pi20  & ~n9015;
  assign n9018 = ~n9016 & ~n9017;
  assign n9019 = n9008 & ~n9018;
  assign n9020 = ~n3166 & n5435;
  assign n9021 = ~n3097 & n6055;
  assign n9022 = n5429 & n7071;
  assign n9023 = ~n3005 & n6071;
  assign n9024 = ~n9022 & ~n9023;
  assign n9025 = ~n9021 & n9024;
  assign n9026 = ~n9020 & n9025;
  assign n9027 = ~pi20  & ~n9026;
  assign n9028 = pi20  & n9026;
  assign n9029 = ~n9027 & ~n9028;
  assign n9030 = n8724 & ~n8726;
  assign n9031 = ~n8727 & ~n9030;
  assign n9032 = ~n9029 & n9031;
  assign n9033 = ~n9029 & ~n9031;
  assign n9034 = n9029 & n9031;
  assign n9035 = ~n9033 & ~n9034;
  assign n9036 = ~n3226 & n5435;
  assign n9037 = ~n3166 & n6055;
  assign n9038 = n5429 & n7121;
  assign n9039 = ~n3097 & n6071;
  assign n9040 = ~n9038 & ~n9039;
  assign n9041 = ~n9037 & n9040;
  assign n9042 = ~n9036 & n9041;
  assign n9043 = pi20  & n9042;
  assign n9044 = ~pi20  & ~n9042;
  assign n9045 = ~n9043 & ~n9044;
  assign n9046 = n8712 & n8722;
  assign n9047 = ~n8723 & ~n9046;
  assign n9048 = ~n9045 & n9047;
  assign n9049 = ~n3263 & n5435;
  assign n9050 = ~n3226 & n6055;
  assign n9051 = n5429 & n7175;
  assign n9052 = ~n3166 & n6071;
  assign n9053 = ~n9051 & ~n9052;
  assign n9054 = ~n9050 & n9053;
  assign n9055 = ~n9049 & n9054;
  assign n9056 = ~pi20  & ~n9055;
  assign n9057 = pi20  & n9055;
  assign n9058 = ~n9056 & ~n9057;
  assign n9059 = pi23  & ~n8700;
  assign n9060 = n8707 & ~n9059;
  assign n9061 = ~n8707 & n9059;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = ~n9058 & n9062;
  assign n9064 = ~n9058 & ~n9062;
  assign n9065 = n9058 & n9062;
  assign n9066 = ~n9064 & ~n9065;
  assign n9067 = ~n3360 & n5435;
  assign n9068 = ~n3263 & n6055;
  assign n9069 = n5429 & n7221;
  assign n9070 = ~n3226 & n6071;
  assign n9071 = ~n9069 & ~n9070;
  assign n9072 = ~n9068 & n9071;
  assign n9073 = ~n9067 & n9072;
  assign n9074 = pi20  & n9073;
  assign n9075 = ~pi20  & ~n9073;
  assign n9076 = ~n9074 & ~n9075;
  assign n9077 = pi23  & n8698;
  assign n9078 = ~n8697 & n9077;
  assign n9079 = n8697 & ~n9077;
  assign n9080 = ~n9078 & ~n9079;
  assign n9081 = ~n9076 & n9080;
  assign n9082 = n5429 & ~n7942;
  assign n9083 = ~n3506 & n6071;
  assign n9084 = ~n3450 & n6055;
  assign n9085 = ~n9083 & ~n9084;
  assign n9086 = ~n9082 & n9085;
  assign n9087 = ~n3450 & ~n5425;
  assign n9088 = pi20  & ~n9087;
  assign n9089 = n9086 & n9088;
  assign n9090 = ~n3450 & n5435;
  assign n9091 = ~n3506 & n6055;
  assign n9092 = n5429 & n7265;
  assign n9093 = ~n3360 & n6071;
  assign n9094 = ~n9092 & ~n9093;
  assign n9095 = ~n9091 & n9094;
  assign n9096 = ~n9090 & n9095;
  assign n9097 = n9089 & n9096;
  assign n9098 = n8698 & n9097;
  assign n9099 = ~n8698 & n9097;
  assign n9100 = n8698 & ~n9097;
  assign n9101 = ~n9099 & ~n9100;
  assign n9102 = ~n3506 & n5435;
  assign n9103 = ~n3360 & n6055;
  assign n9104 = n5429 & n7323;
  assign n9105 = ~n3263 & n6071;
  assign n9106 = ~n9104 & ~n9105;
  assign n9107 = ~n9103 & n9106;
  assign n9108 = ~n9102 & n9107;
  assign n9109 = pi20  & n9108;
  assign n9110 = ~pi20  & ~n9108;
  assign n9111 = ~n9109 & ~n9110;
  assign n9112 = ~n9101 & ~n9111;
  assign n9113 = ~n9098 & ~n9112;
  assign n9114 = n9076 & ~n9080;
  assign n9115 = ~n9081 & ~n9114;
  assign n9116 = ~n9113 & n9115;
  assign n9117 = ~n9081 & ~n9116;
  assign n9118 = ~n9066 & ~n9117;
  assign n9119 = ~n9063 & ~n9118;
  assign n9120 = n9045 & ~n9047;
  assign n9121 = ~n9048 & ~n9120;
  assign n9122 = ~n9119 & n9121;
  assign n9123 = ~n9048 & ~n9122;
  assign n9124 = ~n9035 & ~n9123;
  assign n9125 = ~n9032 & ~n9124;
  assign n9126 = n9008 & n9018;
  assign n9127 = ~n9008 & ~n9018;
  assign n9128 = ~n9126 & ~n9127;
  assign n9129 = ~n9125 & ~n9128;
  assign n9130 = ~n9019 & ~n9129;
  assign n9131 = n8995 & n9005;
  assign n9132 = ~n8995 & ~n9005;
  assign n9133 = ~n9131 & ~n9132;
  assign n9134 = ~n9130 & ~n9133;
  assign n9135 = ~n9006 & ~n9134;
  assign n9136 = ~n8982 & n8992;
  assign n9137 = ~n8993 & ~n9136;
  assign n9138 = ~n9135 & n9137;
  assign n9139 = ~n8993 & ~n9138;
  assign n9140 = n8976 & n8979;
  assign n9141 = ~n8980 & ~n9140;
  assign n9142 = ~n9139 & n9141;
  assign n9143 = ~n8980 & ~n9142;
  assign n9144 = ~n8966 & ~n9143;
  assign n9145 = ~n8963 & ~n9144;
  assign n9146 = n8939 & n8949;
  assign n9147 = ~n8939 & ~n8949;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = ~n9145 & ~n9148;
  assign n9150 = ~n8950 & ~n9149;
  assign n9151 = n8926 & n8936;
  assign n9152 = ~n8926 & ~n8936;
  assign n9153 = ~n9151 & ~n9152;
  assign n9154 = ~n9150 & ~n9153;
  assign n9155 = ~n8937 & ~n9154;
  assign n9156 = n8913 & n8923;
  assign n9157 = ~n8913 & ~n8923;
  assign n9158 = ~n9156 & ~n9157;
  assign n9159 = ~n9155 & ~n9158;
  assign n9160 = ~n8924 & ~n9159;
  assign n9161 = n8900 & n8910;
  assign n9162 = ~n8900 & ~n8910;
  assign n9163 = ~n9161 & ~n9162;
  assign n9164 = ~n9160 & ~n9163;
  assign n9165 = ~n8911 & ~n9164;
  assign n9166 = n8887 & n8897;
  assign n9167 = ~n8887 & ~n8897;
  assign n9168 = ~n9166 & ~n9167;
  assign n9169 = ~n9165 & ~n9168;
  assign n9170 = ~n8898 & ~n9169;
  assign n9171 = n8874 & n8884;
  assign n9172 = ~n8874 & ~n8884;
  assign n9173 = ~n9171 & ~n9172;
  assign n9174 = ~n9170 & ~n9173;
  assign n9175 = ~n8885 & ~n9174;
  assign n9176 = n8861 & n8871;
  assign n9177 = ~n8861 & ~n8871;
  assign n9178 = ~n9176 & ~n9177;
  assign n9179 = ~n9175 & ~n9178;
  assign n9180 = ~n8872 & ~n9179;
  assign n9181 = n8778 & ~n8780;
  assign n9182 = ~n8781 & ~n9181;
  assign n9183 = ~n9180 & n9182;
  assign n9184 = ~n1900 & n6184;
  assign n9185 = ~n1811 & n6527;
  assign n9186 = n4967 & n6185;
  assign n9187 = ~n1740 & n6543;
  assign n9188 = ~n9186 & ~n9187;
  assign n9189 = ~n9185 & n9188;
  assign n9190 = ~n9184 & n9189;
  assign n9191 = ~pi17  & ~n9190;
  assign n9192 = pi17  & n9190;
  assign n9193 = ~n9191 & ~n9192;
  assign n9194 = n9180 & ~n9182;
  assign n9195 = ~n9183 & ~n9194;
  assign n9196 = ~n9193 & n9195;
  assign n9197 = ~n9183 & ~n9196;
  assign n9198 = ~n8787 & ~n8788;
  assign n9199 = ~n8798 & n9198;
  assign n9200 = n8798 & ~n9198;
  assign n9201 = ~n9199 & ~n9200;
  assign n9202 = ~n9197 & n9201;
  assign n9203 = n9197 & ~n9201;
  assign n9204 = ~n1531 & n6835;
  assign n9205 = ~n1426 & n7460;
  assign n9206 = n4533 & n6836;
  assign n9207 = ~n1338 & n7487;
  assign n9208 = ~n9206 & ~n9207;
  assign n9209 = ~n9205 & n9208;
  assign n9210 = ~n9204 & n9209;
  assign n9211 = pi14  & n9210;
  assign n9212 = ~pi14  & ~n9210;
  assign n9213 = ~n9211 & ~n9212;
  assign n9214 = ~n9203 & ~n9213;
  assign n9215 = ~n9202 & ~n9214;
  assign n9216 = n8859 & ~n9215;
  assign n9217 = ~n8859 & n9215;
  assign n9218 = ~n1107 & n7654;
  assign n9219 = ~n1005 & n8091;
  assign n9220 = n4106 & n7648;
  assign n9221 = ~n894 & n8120;
  assign n9222 = ~n9220 & ~n9221;
  assign n9223 = ~n9219 & n9222;
  assign n9224 = ~n9218 & n9223;
  assign n9225 = pi11  & n9224;
  assign n9226 = ~pi11  & ~n9224;
  assign n9227 = ~n9225 & ~n9226;
  assign n9228 = ~n9217 & ~n9227;
  assign n9229 = ~n9216 & ~n9228;
  assign n9230 = ~n8855 & ~n9229;
  assign n9231 = n8855 & n9229;
  assign n9232 = ~n9230 & ~n9231;
  assign n9233 = ~n8494 & n8814;
  assign n9234 = ~n8815 & ~n9233;
  assign n9235 = n9232 & n9234;
  assign n9236 = ~n9230 & ~n9235;
  assign n9237 = ~n3744 & n8468;
  assign n9238 = n8464 & ~n8472;
  assign n9239 = ~n554 & n9238;
  assign n9240 = ~n720 & n8474;
  assign n9241 = ~n9239 & ~n9240;
  assign n9242 = ~n9237 & n9241;
  assign n9243 = pi8  & n9242;
  assign n9244 = ~pi8  & ~n9242;
  assign n9245 = ~n9243 & ~n9244;
  assign n9246 = ~n9236 & ~n9245;
  assign n9247 = n9236 & n9245;
  assign n9248 = ~n9246 & ~n9247;
  assign n9249 = ~n8821 & ~n8822;
  assign n9250 = ~n8832 & n9249;
  assign n9251 = n8832 & ~n9249;
  assign n9252 = ~n9250 & ~n9251;
  assign n9253 = n9248 & n9252;
  assign n9254 = ~n9246 & ~n9253;
  assign n9255 = ~n8835 & ~n8836;
  assign n9256 = n8840 & n9255;
  assign n9257 = ~n8840 & ~n9255;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = ~n9254 & n9258;
  assign n9260 = n9254 & ~n9258;
  assign n9261 = ~n9259 & ~n9260;
  assign n9262 = ~n665 & n8474;
  assign n9263 = ~n720 & n9238;
  assign n9264 = n3979 & n8468;
  assign n9265 = ~n8464 & n8467;
  assign n9266 = ~n554 & n9265;
  assign n9267 = ~n9264 & ~n9266;
  assign n9268 = ~n9263 & n9267;
  assign n9269 = ~n9262 & n9268;
  assign n9270 = pi8  & n9269;
  assign n9271 = ~pi8  & ~n9269;
  assign n9272 = ~n9270 & ~n9271;
  assign n9273 = ~n9216 & ~n9217;
  assign n9274 = ~n9227 & n9273;
  assign n9275 = n9227 & ~n9273;
  assign n9276 = ~n9274 & ~n9275;
  assign n9277 = ~n2006 & n6184;
  assign n9278 = ~n1900 & n6527;
  assign n9279 = n5344 & n6185;
  assign n9280 = ~n1811 & n6543;
  assign n9281 = ~n9279 & ~n9280;
  assign n9282 = ~n9278 & n9281;
  assign n9283 = ~n9277 & n9282;
  assign n9284 = ~pi17  & ~n9283;
  assign n9285 = pi17  & n9283;
  assign n9286 = ~n9284 & ~n9285;
  assign n9287 = ~n9175 & n9178;
  assign n9288 = n9175 & ~n9178;
  assign n9289 = ~n9287 & ~n9288;
  assign n9290 = ~n9286 & ~n9289;
  assign n9291 = ~n2058 & n6184;
  assign n9292 = ~n2006 & n6527;
  assign n9293 = n5180 & n6185;
  assign n9294 = ~n1900 & n6543;
  assign n9295 = ~n9293 & ~n9294;
  assign n9296 = ~n9292 & n9295;
  assign n9297 = ~n9291 & n9296;
  assign n9298 = ~pi17  & ~n9297;
  assign n9299 = pi17  & n9297;
  assign n9300 = ~n9298 & ~n9299;
  assign n9301 = ~n9170 & n9173;
  assign n9302 = n9170 & ~n9173;
  assign n9303 = ~n9301 & ~n9302;
  assign n9304 = ~n9300 & ~n9303;
  assign n9305 = ~n2178 & n6184;
  assign n9306 = ~n2058 & n6527;
  assign n9307 = n5554 & n6185;
  assign n9308 = ~n2006 & n6543;
  assign n9309 = ~n9307 & ~n9308;
  assign n9310 = ~n9306 & n9309;
  assign n9311 = ~n9305 & n9310;
  assign n9312 = ~pi17  & ~n9311;
  assign n9313 = pi17  & n9311;
  assign n9314 = ~n9312 & ~n9313;
  assign n9315 = n9165 & n9168;
  assign n9316 = ~n9169 & ~n9315;
  assign n9317 = ~n9314 & n9316;
  assign n9318 = ~n9314 & ~n9316;
  assign n9319 = n9314 & n9316;
  assign n9320 = ~n9318 & ~n9319;
  assign n9321 = ~n2278 & n6184;
  assign n9322 = ~n2178 & n6527;
  assign n9323 = n5538 & n6185;
  assign n9324 = ~n2058 & n6543;
  assign n9325 = ~n9323 & ~n9324;
  assign n9326 = ~n9322 & n9325;
  assign n9327 = ~n9321 & n9326;
  assign n9328 = ~pi17  & ~n9327;
  assign n9329 = pi17  & n9327;
  assign n9330 = ~n9328 & ~n9329;
  assign n9331 = n9160 & n9163;
  assign n9332 = ~n9164 & ~n9331;
  assign n9333 = ~n9330 & n9332;
  assign n9334 = ~n9330 & ~n9332;
  assign n9335 = n9330 & n9332;
  assign n9336 = ~n9334 & ~n9335;
  assign n9337 = ~n2369 & n6184;
  assign n9338 = ~n2278 & n6527;
  assign n9339 = n5779 & n6185;
  assign n9340 = ~n2178 & n6543;
  assign n9341 = ~n9339 & ~n9340;
  assign n9342 = ~n9338 & n9341;
  assign n9343 = ~n9337 & n9342;
  assign n9344 = ~pi17  & ~n9343;
  assign n9345 = pi17  & n9343;
  assign n9346 = ~n9344 & ~n9345;
  assign n9347 = ~n9155 & n9158;
  assign n9348 = n9155 & ~n9158;
  assign n9349 = ~n9347 & ~n9348;
  assign n9350 = ~n9346 & ~n9349;
  assign n9351 = ~n2457 & n6184;
  assign n9352 = ~n2369 & n6527;
  assign n9353 = n5795 & n6185;
  assign n9354 = ~n2278 & n6543;
  assign n9355 = ~n9353 & ~n9354;
  assign n9356 = ~n9352 & n9355;
  assign n9357 = ~n9351 & n9356;
  assign n9358 = ~pi17  & ~n9357;
  assign n9359 = pi17  & n9357;
  assign n9360 = ~n9358 & ~n9359;
  assign n9361 = ~n9150 & n9153;
  assign n9362 = n9150 & ~n9153;
  assign n9363 = ~n9361 & ~n9362;
  assign n9364 = ~n9360 & ~n9363;
  assign n9365 = ~n2554 & n6184;
  assign n9366 = ~n2457 & n6527;
  assign n9367 = n6185 & n6218;
  assign n9368 = ~n2369 & n6543;
  assign n9369 = ~n9367 & ~n9368;
  assign n9370 = ~n9366 & n9369;
  assign n9371 = ~n9365 & n9370;
  assign n9372 = ~pi17  & ~n9371;
  assign n9373 = pi17  & n9371;
  assign n9374 = ~n9372 & ~n9373;
  assign n9375 = n9145 & n9148;
  assign n9376 = ~n9149 & ~n9375;
  assign n9377 = ~n9374 & n9376;
  assign n9378 = ~n9374 & ~n9376;
  assign n9379 = n9374 & n9376;
  assign n9380 = ~n9378 & ~n9379;
  assign n9381 = n8966 & n9143;
  assign n9382 = ~n9144 & ~n9381;
  assign n9383 = ~n2640 & n6184;
  assign n9384 = ~n2554 & n6527;
  assign n9385 = n5979 & n6185;
  assign n9386 = ~n2457 & n6543;
  assign n9387 = ~n9385 & ~n9386;
  assign n9388 = ~n9384 & n9387;
  assign n9389 = ~n9383 & n9388;
  assign n9390 = pi17  & n9389;
  assign n9391 = ~pi17  & ~n9389;
  assign n9392 = ~n9390 & ~n9391;
  assign n9393 = n9382 & ~n9392;
  assign n9394 = n9139 & ~n9141;
  assign n9395 = ~n9142 & ~n9394;
  assign n9396 = ~n2676 & n6184;
  assign n9397 = ~n2640 & n6527;
  assign n9398 = n6185 & n6445;
  assign n9399 = ~n2554 & n6543;
  assign n9400 = ~n9398 & ~n9399;
  assign n9401 = ~n9397 & n9400;
  assign n9402 = ~n9396 & n9401;
  assign n9403 = pi17  & n9402;
  assign n9404 = ~pi17  & ~n9402;
  assign n9405 = ~n9403 & ~n9404;
  assign n9406 = n9395 & ~n9405;
  assign n9407 = ~n2748 & n6184;
  assign n9408 = ~n2676 & n6527;
  assign n9409 = n6185 & n6597;
  assign n9410 = ~n2640 & n6543;
  assign n9411 = ~n9409 & ~n9410;
  assign n9412 = ~n9408 & n9411;
  assign n9413 = ~n9407 & n9412;
  assign n9414 = ~pi17  & ~n9413;
  assign n9415 = pi17  & n9413;
  assign n9416 = ~n9414 & ~n9415;
  assign n9417 = n9135 & ~n9137;
  assign n9418 = ~n9138 & ~n9417;
  assign n9419 = ~n9416 & n9418;
  assign n9420 = ~n9416 & ~n9418;
  assign n9421 = n9416 & n9418;
  assign n9422 = ~n9420 & ~n9421;
  assign n9423 = ~n2803 & n6184;
  assign n9424 = ~n2748 & n6527;
  assign n9425 = n6185 & n6427;
  assign n9426 = ~n2676 & n6543;
  assign n9427 = ~n9425 & ~n9426;
  assign n9428 = ~n9424 & n9427;
  assign n9429 = ~n9423 & n9428;
  assign n9430 = ~pi17  & ~n9429;
  assign n9431 = pi17  & n9429;
  assign n9432 = ~n9430 & ~n9431;
  assign n9433 = n9130 & n9133;
  assign n9434 = ~n9134 & ~n9433;
  assign n9435 = ~n9432 & n9434;
  assign n9436 = ~n9432 & ~n9434;
  assign n9437 = n9432 & n9434;
  assign n9438 = ~n9436 & ~n9437;
  assign n9439 = ~n2891 & n6184;
  assign n9440 = ~n2803 & n6527;
  assign n9441 = n6185 & n6715;
  assign n9442 = ~n2748 & n6543;
  assign n9443 = ~n9441 & ~n9442;
  assign n9444 = ~n9440 & n9443;
  assign n9445 = ~n9439 & n9444;
  assign n9446 = ~pi17  & ~n9445;
  assign n9447 = pi17  & n9445;
  assign n9448 = ~n9446 & ~n9447;
  assign n9449 = ~n9125 & n9128;
  assign n9450 = n9125 & ~n9128;
  assign n9451 = ~n9449 & ~n9450;
  assign n9452 = ~n9448 & ~n9451;
  assign n9453 = n9035 & n9123;
  assign n9454 = ~n9124 & ~n9453;
  assign n9455 = ~n2927 & n6184;
  assign n9456 = ~n2891 & n6527;
  assign n9457 = n6185 & n7014;
  assign n9458 = ~n2803 & n6543;
  assign n9459 = ~n9457 & ~n9458;
  assign n9460 = ~n9456 & n9459;
  assign n9461 = ~n9455 & n9460;
  assign n9462 = pi17  & n9461;
  assign n9463 = ~pi17  & ~n9461;
  assign n9464 = ~n9462 & ~n9463;
  assign n9465 = n9454 & ~n9464;
  assign n9466 = n9119 & ~n9121;
  assign n9467 = ~n9122 & ~n9466;
  assign n9468 = ~n3005 & n6184;
  assign n9469 = ~n2927 & n6527;
  assign n9470 = n6185 & n7026;
  assign n9471 = ~n2891 & n6543;
  assign n9472 = ~n9470 & ~n9471;
  assign n9473 = ~n9469 & n9472;
  assign n9474 = ~n9468 & n9473;
  assign n9475 = pi17  & n9474;
  assign n9476 = ~pi17  & ~n9474;
  assign n9477 = ~n9475 & ~n9476;
  assign n9478 = n9467 & ~n9477;
  assign n9479 = n9066 & n9117;
  assign n9480 = ~n9118 & ~n9479;
  assign n9481 = ~n3097 & n6184;
  assign n9482 = ~n3005 & n6527;
  assign n9483 = n6185 & n6694;
  assign n9484 = ~n2927 & n6543;
  assign n9485 = ~n9483 & ~n9484;
  assign n9486 = ~n9482 & n9485;
  assign n9487 = ~n9481 & n9486;
  assign n9488 = pi17  & n9487;
  assign n9489 = ~pi17  & ~n9487;
  assign n9490 = ~n9488 & ~n9489;
  assign n9491 = n9480 & ~n9490;
  assign n9492 = ~n3166 & n6184;
  assign n9493 = ~n3097 & n6527;
  assign n9494 = n6185 & n7071;
  assign n9495 = ~n3005 & n6543;
  assign n9496 = ~n9494 & ~n9495;
  assign n9497 = ~n9493 & n9496;
  assign n9498 = ~n9492 & n9497;
  assign n9499 = ~pi17  & ~n9498;
  assign n9500 = pi17  & n9498;
  assign n9501 = ~n9499 & ~n9500;
  assign n9502 = n9113 & ~n9115;
  assign n9503 = ~n9116 & ~n9502;
  assign n9504 = ~n9501 & n9503;
  assign n9505 = ~n9501 & ~n9503;
  assign n9506 = n9501 & n9503;
  assign n9507 = ~n9505 & ~n9506;
  assign n9508 = ~n3226 & n6184;
  assign n9509 = ~n3166 & n6527;
  assign n9510 = n6185 & n7121;
  assign n9511 = ~n3097 & n6543;
  assign n9512 = ~n9510 & ~n9511;
  assign n9513 = ~n9509 & n9512;
  assign n9514 = ~n9508 & n9513;
  assign n9515 = pi17  & n9514;
  assign n9516 = ~pi17  & ~n9514;
  assign n9517 = ~n9515 & ~n9516;
  assign n9518 = n9101 & n9111;
  assign n9519 = ~n9112 & ~n9518;
  assign n9520 = ~n9517 & n9519;
  assign n9521 = ~n3263 & n6184;
  assign n9522 = ~n3226 & n6527;
  assign n9523 = n6185 & n7175;
  assign n9524 = ~n3166 & n6543;
  assign n9525 = ~n9523 & ~n9524;
  assign n9526 = ~n9522 & n9525;
  assign n9527 = ~n9521 & n9526;
  assign n9528 = ~pi17  & ~n9527;
  assign n9529 = pi17  & n9527;
  assign n9530 = ~n9528 & ~n9529;
  assign n9531 = pi20  & ~n9089;
  assign n9532 = n9096 & ~n9531;
  assign n9533 = ~n9096 & n9531;
  assign n9534 = ~n9532 & ~n9533;
  assign n9535 = ~n9530 & n9534;
  assign n9536 = ~n9530 & ~n9534;
  assign n9537 = n9530 & n9534;
  assign n9538 = ~n9536 & ~n9537;
  assign n9539 = ~n3360 & n6184;
  assign n9540 = ~n3263 & n6527;
  assign n9541 = n6185 & n7221;
  assign n9542 = ~n3226 & n6543;
  assign n9543 = ~n9541 & ~n9542;
  assign n9544 = ~n9540 & n9543;
  assign n9545 = ~n9539 & n9544;
  assign n9546 = pi17  & n9545;
  assign n9547 = ~pi17  & ~n9545;
  assign n9548 = ~n9546 & ~n9547;
  assign n9549 = pi20  & n9087;
  assign n9550 = ~n9086 & n9549;
  assign n9551 = n9086 & ~n9549;
  assign n9552 = ~n9550 & ~n9551;
  assign n9553 = ~n9548 & n9552;
  assign n9554 = n6185 & ~n7942;
  assign n9555 = ~n3506 & n6543;
  assign n9556 = ~n3450 & n6527;
  assign n9557 = ~n9555 & ~n9556;
  assign n9558 = ~n9554 & n9557;
  assign n9559 = ~n3450 & ~n6182;
  assign n9560 = pi17  & ~n9559;
  assign n9561 = n9558 & n9560;
  assign n9562 = ~n3450 & n6184;
  assign n9563 = ~n3506 & n6527;
  assign n9564 = n6185 & n7265;
  assign n9565 = ~n3360 & n6543;
  assign n9566 = ~n9564 & ~n9565;
  assign n9567 = ~n9563 & n9566;
  assign n9568 = ~n9562 & n9567;
  assign n9569 = n9561 & n9568;
  assign n9570 = n9087 & n9569;
  assign n9571 = ~n9087 & n9569;
  assign n9572 = n9087 & ~n9569;
  assign n9573 = ~n9571 & ~n9572;
  assign n9574 = ~n3506 & n6184;
  assign n9575 = ~n3360 & n6527;
  assign n9576 = n6185 & n7323;
  assign n9577 = ~n3263 & n6543;
  assign n9578 = ~n9576 & ~n9577;
  assign n9579 = ~n9575 & n9578;
  assign n9580 = ~n9574 & n9579;
  assign n9581 = pi17  & n9580;
  assign n9582 = ~pi17  & ~n9580;
  assign n9583 = ~n9581 & ~n9582;
  assign n9584 = ~n9573 & ~n9583;
  assign n9585 = ~n9570 & ~n9584;
  assign n9586 = n9548 & ~n9552;
  assign n9587 = ~n9553 & ~n9586;
  assign n9588 = ~n9585 & n9587;
  assign n9589 = ~n9553 & ~n9588;
  assign n9590 = ~n9538 & ~n9589;
  assign n9591 = ~n9535 & ~n9590;
  assign n9592 = n9517 & ~n9519;
  assign n9593 = ~n9520 & ~n9592;
  assign n9594 = ~n9591 & n9593;
  assign n9595 = ~n9520 & ~n9594;
  assign n9596 = ~n9507 & ~n9595;
  assign n9597 = ~n9504 & ~n9596;
  assign n9598 = n9480 & n9490;
  assign n9599 = ~n9480 & ~n9490;
  assign n9600 = ~n9598 & ~n9599;
  assign n9601 = ~n9597 & ~n9600;
  assign n9602 = ~n9491 & ~n9601;
  assign n9603 = n9467 & n9477;
  assign n9604 = ~n9467 & ~n9477;
  assign n9605 = ~n9603 & ~n9604;
  assign n9606 = ~n9602 & ~n9605;
  assign n9607 = ~n9478 & ~n9606;
  assign n9608 = ~n9454 & n9464;
  assign n9609 = ~n9465 & ~n9608;
  assign n9610 = ~n9607 & n9609;
  assign n9611 = ~n9465 & ~n9610;
  assign n9612 = n9448 & n9451;
  assign n9613 = ~n9452 & ~n9612;
  assign n9614 = ~n9611 & n9613;
  assign n9615 = ~n9452 & ~n9614;
  assign n9616 = ~n9438 & ~n9615;
  assign n9617 = ~n9435 & ~n9616;
  assign n9618 = ~n9422 & ~n9617;
  assign n9619 = ~n9419 & ~n9618;
  assign n9620 = n9395 & n9405;
  assign n9621 = ~n9395 & ~n9405;
  assign n9622 = ~n9620 & ~n9621;
  assign n9623 = ~n9619 & ~n9622;
  assign n9624 = ~n9406 & ~n9623;
  assign n9625 = ~n9382 & n9392;
  assign n9626 = ~n9393 & ~n9625;
  assign n9627 = ~n9624 & n9626;
  assign n9628 = ~n9393 & ~n9627;
  assign n9629 = ~n9380 & ~n9628;
  assign n9630 = ~n9377 & ~n9629;
  assign n9631 = n9360 & n9363;
  assign n9632 = ~n9364 & ~n9631;
  assign n9633 = ~n9630 & n9632;
  assign n9634 = ~n9364 & ~n9633;
  assign n9635 = n9346 & n9349;
  assign n9636 = ~n9350 & ~n9635;
  assign n9637 = ~n9634 & n9636;
  assign n9638 = ~n9350 & ~n9637;
  assign n9639 = ~n9336 & ~n9638;
  assign n9640 = ~n9333 & ~n9639;
  assign n9641 = ~n9320 & ~n9640;
  assign n9642 = ~n9317 & ~n9641;
  assign n9643 = n9300 & n9303;
  assign n9644 = ~n9304 & ~n9643;
  assign n9645 = ~n9642 & n9644;
  assign n9646 = ~n9304 & ~n9645;
  assign n9647 = n9286 & n9289;
  assign n9648 = ~n9290 & ~n9647;
  assign n9649 = ~n9646 & n9648;
  assign n9650 = ~n9290 & ~n9649;
  assign n9651 = n9193 & ~n9195;
  assign n9652 = ~n9196 & ~n9651;
  assign n9653 = ~n9650 & n9652;
  assign n9654 = ~n1610 & n6835;
  assign n9655 = ~n1531 & n7460;
  assign n9656 = n4724 & n6836;
  assign n9657 = ~n1426 & n7487;
  assign n9658 = ~n9656 & ~n9657;
  assign n9659 = ~n9655 & n9658;
  assign n9660 = ~n9654 & n9659;
  assign n9661 = ~pi14  & ~n9660;
  assign n9662 = pi14  & n9660;
  assign n9663 = ~n9661 & ~n9662;
  assign n9664 = n9650 & ~n9652;
  assign n9665 = ~n9653 & ~n9664;
  assign n9666 = ~n9663 & n9665;
  assign n9667 = ~n9653 & ~n9666;
  assign n9668 = ~n9202 & ~n9203;
  assign n9669 = ~n9213 & n9668;
  assign n9670 = n9213 & ~n9668;
  assign n9671 = ~n9669 & ~n9670;
  assign n9672 = ~n9667 & n9671;
  assign n9673 = n9667 & ~n9671;
  assign n9674 = ~n1230 & n7654;
  assign n9675 = ~n1107 & n8091;
  assign n9676 = n4307 & n7648;
  assign n9677 = ~n1005 & n8120;
  assign n9678 = ~n9676 & ~n9677;
  assign n9679 = ~n9675 & n9678;
  assign n9680 = ~n9674 & n9679;
  assign n9681 = pi11  & n9680;
  assign n9682 = ~pi11  & ~n9680;
  assign n9683 = ~n9681 & ~n9682;
  assign n9684 = ~n9673 & ~n9683;
  assign n9685 = ~n9672 & ~n9684;
  assign n9686 = n9276 & ~n9685;
  assign n9687 = ~n9276 & n9685;
  assign n9688 = ~n795 & n8474;
  assign n9689 = ~n665 & n9238;
  assign n9690 = n4015 & n8468;
  assign n9691 = ~n720 & n9265;
  assign n9692 = ~n9690 & ~n9691;
  assign n9693 = ~n9689 & n9692;
  assign n9694 = ~n9688 & n9693;
  assign n9695 = pi8  & n9694;
  assign n9696 = ~pi8  & ~n9694;
  assign n9697 = ~n9695 & ~n9696;
  assign n9698 = ~n9687 & ~n9697;
  assign n9699 = ~n9686 & ~n9698;
  assign n9700 = ~n9272 & ~n9699;
  assign n9701 = n9272 & ~n9699;
  assign n9702 = ~n9272 & n9699;
  assign n9703 = ~n9701 & ~n9702;
  assign n9704 = ~n9232 & ~n9234;
  assign n9705 = ~n9235 & ~n9704;
  assign n9706 = ~n9703 & n9705;
  assign n9707 = ~n9700 & ~n9706;
  assign n9708 = ~n9248 & ~n9252;
  assign n9709 = ~n9253 & ~n9708;
  assign n9710 = ~n9707 & n9709;
  assign n9711 = n9703 & ~n9705;
  assign n9712 = ~n9706 & ~n9711;
  assign n9713 = pi2  & ~pi3 ;
  assign n9714 = ~pi2  & pi3 ;
  assign n9715 = ~n9713 & ~n9714;
  assign n9716 = pi4  & ~pi5 ;
  assign n9717 = ~pi4  & pi5 ;
  assign n9718 = ~n9716 & ~n9717;
  assign n9719 = ~n9715 & ~n9718;
  assign n9720 = ~n3638 & n9719;
  assign n9721 = ~pi3  & pi4 ;
  assign n9722 = pi3  & ~pi4 ;
  assign n9723 = ~n9721 & ~n9722;
  assign n9724 = n9715 & n9723;
  assign n9725 = ~n9718 & n9724;
  assign n9726 = ~n9720 & ~n9725;
  assign n9727 = ~n554 & ~n9726;
  assign n9728 = pi5  & ~n9727;
  assign n9729 = ~pi5  & n9727;
  assign n9730 = ~n9728 & ~n9729;
  assign n9731 = n9646 & ~n9648;
  assign n9732 = ~n9649 & ~n9731;
  assign n9733 = ~n1740 & n6835;
  assign n9734 = ~n1610 & n7460;
  assign n9735 = n4708 & n6836;
  assign n9736 = ~n1531 & n7487;
  assign n9737 = ~n9735 & ~n9736;
  assign n9738 = ~n9734 & n9737;
  assign n9739 = ~n9733 & n9738;
  assign n9740 = pi14  & n9739;
  assign n9741 = ~pi14  & ~n9739;
  assign n9742 = ~n9740 & ~n9741;
  assign n9743 = n9732 & ~n9742;
  assign n9744 = n9642 & ~n9644;
  assign n9745 = ~n9645 & ~n9744;
  assign n9746 = ~n1811 & n6835;
  assign n9747 = ~n1740 & n7460;
  assign n9748 = n4951 & n6836;
  assign n9749 = ~n1610 & n7487;
  assign n9750 = ~n9748 & ~n9749;
  assign n9751 = ~n9747 & n9750;
  assign n9752 = ~n9746 & n9751;
  assign n9753 = pi14  & n9752;
  assign n9754 = ~pi14  & ~n9752;
  assign n9755 = ~n9753 & ~n9754;
  assign n9756 = n9745 & ~n9755;
  assign n9757 = n9320 & n9640;
  assign n9758 = ~n9641 & ~n9757;
  assign n9759 = ~n1900 & n6835;
  assign n9760 = ~n1811 & n7460;
  assign n9761 = n4967 & n6836;
  assign n9762 = ~n1740 & n7487;
  assign n9763 = ~n9761 & ~n9762;
  assign n9764 = ~n9760 & n9763;
  assign n9765 = ~n9759 & n9764;
  assign n9766 = pi14  & n9765;
  assign n9767 = ~pi14  & ~n9765;
  assign n9768 = ~n9766 & ~n9767;
  assign n9769 = n9758 & ~n9768;
  assign n9770 = n9336 & n9638;
  assign n9771 = ~n9639 & ~n9770;
  assign n9772 = ~n2006 & n6835;
  assign n9773 = ~n1900 & n7460;
  assign n9774 = n5344 & n6836;
  assign n9775 = ~n1811 & n7487;
  assign n9776 = ~n9774 & ~n9775;
  assign n9777 = ~n9773 & n9776;
  assign n9778 = ~n9772 & n9777;
  assign n9779 = pi14  & n9778;
  assign n9780 = ~pi14  & ~n9778;
  assign n9781 = ~n9779 & ~n9780;
  assign n9782 = n9771 & ~n9781;
  assign n9783 = n9634 & ~n9636;
  assign n9784 = ~n9637 & ~n9783;
  assign n9785 = ~n2058 & n6835;
  assign n9786 = ~n2006 & n7460;
  assign n9787 = n5180 & n6836;
  assign n9788 = ~n1900 & n7487;
  assign n9789 = ~n9787 & ~n9788;
  assign n9790 = ~n9786 & n9789;
  assign n9791 = ~n9785 & n9790;
  assign n9792 = pi14  & n9791;
  assign n9793 = ~pi14  & ~n9791;
  assign n9794 = ~n9792 & ~n9793;
  assign n9795 = n9784 & ~n9794;
  assign n9796 = n9630 & ~n9632;
  assign n9797 = ~n9633 & ~n9796;
  assign n9798 = ~n2178 & n6835;
  assign n9799 = ~n2058 & n7460;
  assign n9800 = n5554 & n6836;
  assign n9801 = ~n2006 & n7487;
  assign n9802 = ~n9800 & ~n9801;
  assign n9803 = ~n9799 & n9802;
  assign n9804 = ~n9798 & n9803;
  assign n9805 = pi14  & n9804;
  assign n9806 = ~pi14  & ~n9804;
  assign n9807 = ~n9805 & ~n9806;
  assign n9808 = n9797 & ~n9807;
  assign n9809 = n9380 & n9628;
  assign n9810 = ~n9629 & ~n9809;
  assign n9811 = ~n2278 & n6835;
  assign n9812 = ~n2178 & n7460;
  assign n9813 = n5538 & n6836;
  assign n9814 = ~n2058 & n7487;
  assign n9815 = ~n9813 & ~n9814;
  assign n9816 = ~n9812 & n9815;
  assign n9817 = ~n9811 & n9816;
  assign n9818 = pi14  & n9817;
  assign n9819 = ~pi14  & ~n9817;
  assign n9820 = ~n9818 & ~n9819;
  assign n9821 = n9810 & ~n9820;
  assign n9822 = ~n2369 & n6835;
  assign n9823 = ~n2278 & n7460;
  assign n9824 = n5779 & n6836;
  assign n9825 = ~n2178 & n7487;
  assign n9826 = ~n9824 & ~n9825;
  assign n9827 = ~n9823 & n9826;
  assign n9828 = ~n9822 & n9827;
  assign n9829 = ~pi14  & ~n9828;
  assign n9830 = pi14  & n9828;
  assign n9831 = ~n9829 & ~n9830;
  assign n9832 = n9624 & ~n9626;
  assign n9833 = ~n9627 & ~n9832;
  assign n9834 = ~n9831 & n9833;
  assign n9835 = ~n9831 & ~n9833;
  assign n9836 = n9831 & n9833;
  assign n9837 = ~n9835 & ~n9836;
  assign n9838 = ~n2457 & n6835;
  assign n9839 = ~n2369 & n7460;
  assign n9840 = n5795 & n6836;
  assign n9841 = ~n2278 & n7487;
  assign n9842 = ~n9840 & ~n9841;
  assign n9843 = ~n9839 & n9842;
  assign n9844 = ~n9838 & n9843;
  assign n9845 = ~pi14  & ~n9844;
  assign n9846 = pi14  & n9844;
  assign n9847 = ~n9845 & ~n9846;
  assign n9848 = n9619 & n9622;
  assign n9849 = ~n9623 & ~n9848;
  assign n9850 = ~n9847 & n9849;
  assign n9851 = ~n9847 & ~n9849;
  assign n9852 = n9847 & n9849;
  assign n9853 = ~n9851 & ~n9852;
  assign n9854 = n9422 & n9617;
  assign n9855 = ~n9618 & ~n9854;
  assign n9856 = ~n2554 & n6835;
  assign n9857 = ~n2457 & n7460;
  assign n9858 = n6218 & n6836;
  assign n9859 = ~n2369 & n7487;
  assign n9860 = ~n9858 & ~n9859;
  assign n9861 = ~n9857 & n9860;
  assign n9862 = ~n9856 & n9861;
  assign n9863 = pi14  & n9862;
  assign n9864 = ~pi14  & ~n9862;
  assign n9865 = ~n9863 & ~n9864;
  assign n9866 = n9855 & ~n9865;
  assign n9867 = n9438 & n9615;
  assign n9868 = ~n9616 & ~n9867;
  assign n9869 = ~n2640 & n6835;
  assign n9870 = ~n2554 & n7460;
  assign n9871 = n5979 & n6836;
  assign n9872 = ~n2457 & n7487;
  assign n9873 = ~n9871 & ~n9872;
  assign n9874 = ~n9870 & n9873;
  assign n9875 = ~n9869 & n9874;
  assign n9876 = pi14  & n9875;
  assign n9877 = ~pi14  & ~n9875;
  assign n9878 = ~n9876 & ~n9877;
  assign n9879 = n9868 & ~n9878;
  assign n9880 = n9611 & ~n9613;
  assign n9881 = ~n9614 & ~n9880;
  assign n9882 = ~n2676 & n6835;
  assign n9883 = ~n2640 & n7460;
  assign n9884 = n6445 & n6836;
  assign n9885 = ~n2554 & n7487;
  assign n9886 = ~n9884 & ~n9885;
  assign n9887 = ~n9883 & n9886;
  assign n9888 = ~n9882 & n9887;
  assign n9889 = pi14  & n9888;
  assign n9890 = ~pi14  & ~n9888;
  assign n9891 = ~n9889 & ~n9890;
  assign n9892 = n9881 & ~n9891;
  assign n9893 = ~n2748 & n6835;
  assign n9894 = ~n2676 & n7460;
  assign n9895 = n6597 & n6836;
  assign n9896 = ~n2640 & n7487;
  assign n9897 = ~n9895 & ~n9896;
  assign n9898 = ~n9894 & n9897;
  assign n9899 = ~n9893 & n9898;
  assign n9900 = ~pi14  & ~n9899;
  assign n9901 = pi14  & n9899;
  assign n9902 = ~n9900 & ~n9901;
  assign n9903 = n9607 & ~n9609;
  assign n9904 = ~n9610 & ~n9903;
  assign n9905 = ~n9902 & n9904;
  assign n9906 = ~n9902 & ~n9904;
  assign n9907 = n9902 & n9904;
  assign n9908 = ~n9906 & ~n9907;
  assign n9909 = ~n2803 & n6835;
  assign n9910 = ~n2748 & n7460;
  assign n9911 = n6427 & n6836;
  assign n9912 = ~n2676 & n7487;
  assign n9913 = ~n9911 & ~n9912;
  assign n9914 = ~n9910 & n9913;
  assign n9915 = ~n9909 & n9914;
  assign n9916 = ~pi14  & ~n9915;
  assign n9917 = pi14  & n9915;
  assign n9918 = ~n9916 & ~n9917;
  assign n9919 = n9602 & n9605;
  assign n9920 = ~n9606 & ~n9919;
  assign n9921 = ~n9918 & n9920;
  assign n9922 = ~n9918 & ~n9920;
  assign n9923 = n9918 & n9920;
  assign n9924 = ~n9922 & ~n9923;
  assign n9925 = ~n2891 & n6835;
  assign n9926 = ~n2803 & n7460;
  assign n9927 = n6715 & n6836;
  assign n9928 = ~n2748 & n7487;
  assign n9929 = ~n9927 & ~n9928;
  assign n9930 = ~n9926 & n9929;
  assign n9931 = ~n9925 & n9930;
  assign n9932 = ~pi14  & ~n9931;
  assign n9933 = pi14  & n9931;
  assign n9934 = ~n9932 & ~n9933;
  assign n9935 = ~n9597 & n9600;
  assign n9936 = n9597 & ~n9600;
  assign n9937 = ~n9935 & ~n9936;
  assign n9938 = ~n9934 & ~n9937;
  assign n9939 = n9507 & n9595;
  assign n9940 = ~n9596 & ~n9939;
  assign n9941 = ~n2927 & n6835;
  assign n9942 = ~n2891 & n7460;
  assign n9943 = n6836 & n7014;
  assign n9944 = ~n2803 & n7487;
  assign n9945 = ~n9943 & ~n9944;
  assign n9946 = ~n9942 & n9945;
  assign n9947 = ~n9941 & n9946;
  assign n9948 = pi14  & n9947;
  assign n9949 = ~pi14  & ~n9947;
  assign n9950 = ~n9948 & ~n9949;
  assign n9951 = n9940 & ~n9950;
  assign n9952 = n9591 & ~n9593;
  assign n9953 = ~n9594 & ~n9952;
  assign n9954 = ~n3005 & n6835;
  assign n9955 = ~n2927 & n7460;
  assign n9956 = n6836 & n7026;
  assign n9957 = ~n2891 & n7487;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = ~n9955 & n9958;
  assign n9960 = ~n9954 & n9959;
  assign n9961 = pi14  & n9960;
  assign n9962 = ~pi14  & ~n9960;
  assign n9963 = ~n9961 & ~n9962;
  assign n9964 = n9953 & ~n9963;
  assign n9965 = n9538 & n9589;
  assign n9966 = ~n9590 & ~n9965;
  assign n9967 = ~n3097 & n6835;
  assign n9968 = ~n3005 & n7460;
  assign n9969 = n6694 & n6836;
  assign n9970 = ~n2927 & n7487;
  assign n9971 = ~n9969 & ~n9970;
  assign n9972 = ~n9968 & n9971;
  assign n9973 = ~n9967 & n9972;
  assign n9974 = pi14  & n9973;
  assign n9975 = ~pi14  & ~n9973;
  assign n9976 = ~n9974 & ~n9975;
  assign n9977 = n9966 & ~n9976;
  assign n9978 = ~n3166 & n6835;
  assign n9979 = ~n3097 & n7460;
  assign n9980 = n6836 & n7071;
  assign n9981 = ~n3005 & n7487;
  assign n9982 = ~n9980 & ~n9981;
  assign n9983 = ~n9979 & n9982;
  assign n9984 = ~n9978 & n9983;
  assign n9985 = ~pi14  & ~n9984;
  assign n9986 = pi14  & n9984;
  assign n9987 = ~n9985 & ~n9986;
  assign n9988 = n9585 & ~n9587;
  assign n9989 = ~n9588 & ~n9988;
  assign n9990 = ~n9987 & n9989;
  assign n9991 = ~n9987 & ~n9989;
  assign n9992 = n9987 & n9989;
  assign n9993 = ~n9991 & ~n9992;
  assign n9994 = ~n3226 & n6835;
  assign n9995 = ~n3166 & n7460;
  assign n9996 = n6836 & n7121;
  assign n9997 = ~n3097 & n7487;
  assign n9998 = ~n9996 & ~n9997;
  assign n9999 = ~n9995 & n9998;
  assign n10000 = ~n9994 & n9999;
  assign n10001 = pi14  & n10000;
  assign n10002 = ~pi14  & ~n10000;
  assign n10003 = ~n10001 & ~n10002;
  assign n10004 = n9573 & n9583;
  assign n10005 = ~n9584 & ~n10004;
  assign n10006 = ~n10003 & n10005;
  assign n10007 = ~n3263 & n6835;
  assign n10008 = ~n3226 & n7460;
  assign n10009 = n6836 & n7175;
  assign n10010 = ~n3166 & n7487;
  assign n10011 = ~n10009 & ~n10010;
  assign n10012 = ~n10008 & n10011;
  assign n10013 = ~n10007 & n10012;
  assign n10014 = ~pi14  & ~n10013;
  assign n10015 = pi14  & n10013;
  assign n10016 = ~n10014 & ~n10015;
  assign n10017 = pi17  & ~n9561;
  assign n10018 = n9568 & ~n10017;
  assign n10019 = ~n9568 & n10017;
  assign n10020 = ~n10018 & ~n10019;
  assign n10021 = ~n10016 & n10020;
  assign n10022 = ~n10016 & ~n10020;
  assign n10023 = n10016 & n10020;
  assign n10024 = ~n10022 & ~n10023;
  assign n10025 = ~n3360 & n6835;
  assign n10026 = ~n3263 & n7460;
  assign n10027 = n6836 & n7221;
  assign n10028 = ~n3226 & n7487;
  assign n10029 = ~n10027 & ~n10028;
  assign n10030 = ~n10026 & n10029;
  assign n10031 = ~n10025 & n10030;
  assign n10032 = pi14  & n10031;
  assign n10033 = ~pi14  & ~n10031;
  assign n10034 = ~n10032 & ~n10033;
  assign n10035 = pi17  & n9559;
  assign n10036 = ~n9558 & n10035;
  assign n10037 = n9558 & ~n10035;
  assign n10038 = ~n10036 & ~n10037;
  assign n10039 = ~n10034 & n10038;
  assign n10040 = n6836 & ~n7942;
  assign n10041 = ~n3506 & n7487;
  assign n10042 = ~n3450 & n7460;
  assign n10043 = ~n10041 & ~n10042;
  assign n10044 = ~n10040 & n10043;
  assign n10045 = ~n3450 & ~n6833;
  assign n10046 = pi14  & ~n10045;
  assign n10047 = n10044 & n10046;
  assign n10048 = ~n3450 & n6835;
  assign n10049 = ~n3506 & n7460;
  assign n10050 = n6836 & n7265;
  assign n10051 = ~n3360 & n7487;
  assign n10052 = ~n10050 & ~n10051;
  assign n10053 = ~n10049 & n10052;
  assign n10054 = ~n10048 & n10053;
  assign n10055 = n10047 & n10054;
  assign n10056 = n9559 & n10055;
  assign n10057 = ~n9559 & n10055;
  assign n10058 = n9559 & ~n10055;
  assign n10059 = ~n10057 & ~n10058;
  assign n10060 = ~n3506 & n6835;
  assign n10061 = ~n3360 & n7460;
  assign n10062 = n6836 & n7323;
  assign n10063 = ~n3263 & n7487;
  assign n10064 = ~n10062 & ~n10063;
  assign n10065 = ~n10061 & n10064;
  assign n10066 = ~n10060 & n10065;
  assign n10067 = pi14  & n10066;
  assign n10068 = ~pi14  & ~n10066;
  assign n10069 = ~n10067 & ~n10068;
  assign n10070 = ~n10059 & ~n10069;
  assign n10071 = ~n10056 & ~n10070;
  assign n10072 = n10034 & ~n10038;
  assign n10073 = ~n10039 & ~n10072;
  assign n10074 = ~n10071 & n10073;
  assign n10075 = ~n10039 & ~n10074;
  assign n10076 = ~n10024 & ~n10075;
  assign n10077 = ~n10021 & ~n10076;
  assign n10078 = n10003 & ~n10005;
  assign n10079 = ~n10006 & ~n10078;
  assign n10080 = ~n10077 & n10079;
  assign n10081 = ~n10006 & ~n10080;
  assign n10082 = ~n9993 & ~n10081;
  assign n10083 = ~n9990 & ~n10082;
  assign n10084 = n9966 & n9976;
  assign n10085 = ~n9966 & ~n9976;
  assign n10086 = ~n10084 & ~n10085;
  assign n10087 = ~n10083 & ~n10086;
  assign n10088 = ~n9977 & ~n10087;
  assign n10089 = n9953 & n9963;
  assign n10090 = ~n9953 & ~n9963;
  assign n10091 = ~n10089 & ~n10090;
  assign n10092 = ~n10088 & ~n10091;
  assign n10093 = ~n9964 & ~n10092;
  assign n10094 = ~n9940 & n9950;
  assign n10095 = ~n9951 & ~n10094;
  assign n10096 = ~n10093 & n10095;
  assign n10097 = ~n9951 & ~n10096;
  assign n10098 = n9934 & n9937;
  assign n10099 = ~n9938 & ~n10098;
  assign n10100 = ~n10097 & n10099;
  assign n10101 = ~n9938 & ~n10100;
  assign n10102 = ~n9924 & ~n10101;
  assign n10103 = ~n9921 & ~n10102;
  assign n10104 = ~n9908 & ~n10103;
  assign n10105 = ~n9905 & ~n10104;
  assign n10106 = n9881 & n9891;
  assign n10107 = ~n9881 & ~n9891;
  assign n10108 = ~n10106 & ~n10107;
  assign n10109 = ~n10105 & ~n10108;
  assign n10110 = ~n9892 & ~n10109;
  assign n10111 = n9868 & n9878;
  assign n10112 = ~n9868 & ~n9878;
  assign n10113 = ~n10111 & ~n10112;
  assign n10114 = ~n10110 & ~n10113;
  assign n10115 = ~n9879 & ~n10114;
  assign n10116 = ~n9855 & n9865;
  assign n10117 = ~n9866 & ~n10116;
  assign n10118 = ~n10115 & n10117;
  assign n10119 = ~n9866 & ~n10118;
  assign n10120 = ~n9853 & ~n10119;
  assign n10121 = ~n9850 & ~n10120;
  assign n10122 = ~n9837 & ~n10121;
  assign n10123 = ~n9834 & ~n10122;
  assign n10124 = n9810 & n9820;
  assign n10125 = ~n9810 & ~n9820;
  assign n10126 = ~n10124 & ~n10125;
  assign n10127 = ~n10123 & ~n10126;
  assign n10128 = ~n9821 & ~n10127;
  assign n10129 = n9797 & n9807;
  assign n10130 = ~n9797 & ~n9807;
  assign n10131 = ~n10129 & ~n10130;
  assign n10132 = ~n10128 & ~n10131;
  assign n10133 = ~n9808 & ~n10132;
  assign n10134 = n9784 & n9794;
  assign n10135 = ~n9784 & ~n9794;
  assign n10136 = ~n10134 & ~n10135;
  assign n10137 = ~n10133 & ~n10136;
  assign n10138 = ~n9795 & ~n10137;
  assign n10139 = n9771 & n9781;
  assign n10140 = ~n9771 & ~n9781;
  assign n10141 = ~n10139 & ~n10140;
  assign n10142 = ~n10138 & ~n10141;
  assign n10143 = ~n9782 & ~n10142;
  assign n10144 = n9758 & n9768;
  assign n10145 = ~n9758 & ~n9768;
  assign n10146 = ~n10144 & ~n10145;
  assign n10147 = ~n10143 & ~n10146;
  assign n10148 = ~n9769 & ~n10147;
  assign n10149 = n9745 & n9755;
  assign n10150 = ~n9745 & ~n9755;
  assign n10151 = ~n10149 & ~n10150;
  assign n10152 = ~n10148 & ~n10151;
  assign n10153 = ~n9756 & ~n10152;
  assign n10154 = n9732 & n9742;
  assign n10155 = ~n9732 & ~n9742;
  assign n10156 = ~n10154 & ~n10155;
  assign n10157 = ~n10153 & ~n10156;
  assign n10158 = ~n9743 & ~n10157;
  assign n10159 = n9663 & ~n9665;
  assign n10160 = ~n9666 & ~n10159;
  assign n10161 = ~n10158 & n10160;
  assign n10162 = ~n1338 & n7654;
  assign n10163 = ~n1230 & n8091;
  assign n10164 = n4323 & n7648;
  assign n10165 = ~n1107 & n8120;
  assign n10166 = ~n10164 & ~n10165;
  assign n10167 = ~n10163 & n10166;
  assign n10168 = ~n10162 & n10167;
  assign n10169 = ~pi11  & ~n10168;
  assign n10170 = pi11  & n10168;
  assign n10171 = ~n10169 & ~n10170;
  assign n10172 = n10158 & ~n10160;
  assign n10173 = ~n10161 & ~n10172;
  assign n10174 = ~n10171 & n10173;
  assign n10175 = ~n10161 & ~n10174;
  assign n10176 = ~n9672 & ~n9673;
  assign n10177 = ~n9683 & n10176;
  assign n10178 = n9683 & ~n10176;
  assign n10179 = ~n10177 & ~n10178;
  assign n10180 = ~n10175 & n10179;
  assign n10181 = n10175 & ~n10179;
  assign n10182 = ~n894 & n8474;
  assign n10183 = ~n795 & n9238;
  assign n10184 = n3959 & n8468;
  assign n10185 = ~n665 & n9265;
  assign n10186 = ~n10184 & ~n10185;
  assign n10187 = ~n10183 & n10186;
  assign n10188 = ~n10182 & n10187;
  assign n10189 = pi8  & n10188;
  assign n10190 = ~pi8  & ~n10188;
  assign n10191 = ~n10189 & ~n10190;
  assign n10192 = ~n10181 & ~n10191;
  assign n10193 = ~n10180 & ~n10192;
  assign n10194 = ~n9730 & ~n10193;
  assign n10195 = n9730 & n10193;
  assign n10196 = ~n9686 & ~n9687;
  assign n10197 = ~n9697 & n10196;
  assign n10198 = n9697 & ~n10196;
  assign n10199 = ~n10197 & ~n10198;
  assign n10200 = ~n10195 & n10199;
  assign n10201 = ~n10194 & ~n10200;
  assign n10202 = n9712 & ~n10201;
  assign n10203 = ~n1426 & n7654;
  assign n10204 = ~n1338 & n8091;
  assign n10205 = n4753 & n7648;
  assign n10206 = ~n1230 & n8120;
  assign n10207 = ~n10205 & ~n10206;
  assign n10208 = ~n10204 & n10207;
  assign n10209 = ~n10203 & n10208;
  assign n10210 = ~pi11  & ~n10209;
  assign n10211 = pi11  & n10209;
  assign n10212 = ~n10210 & ~n10211;
  assign n10213 = n10153 & n10156;
  assign n10214 = ~n10157 & ~n10213;
  assign n10215 = ~n10212 & n10214;
  assign n10216 = ~n10212 & ~n10214;
  assign n10217 = n10212 & n10214;
  assign n10218 = ~n10216 & ~n10217;
  assign n10219 = ~n1531 & n7654;
  assign n10220 = ~n1426 & n8091;
  assign n10221 = n4533 & n7648;
  assign n10222 = ~n1338 & n8120;
  assign n10223 = ~n10221 & ~n10222;
  assign n10224 = ~n10220 & n10223;
  assign n10225 = ~n10219 & n10224;
  assign n10226 = ~pi11  & ~n10225;
  assign n10227 = pi11  & n10225;
  assign n10228 = ~n10226 & ~n10227;
  assign n10229 = n10148 & n10151;
  assign n10230 = ~n10152 & ~n10229;
  assign n10231 = ~n10228 & n10230;
  assign n10232 = ~n10228 & ~n10230;
  assign n10233 = n10228 & n10230;
  assign n10234 = ~n10232 & ~n10233;
  assign n10235 = ~n1610 & n7654;
  assign n10236 = ~n1531 & n8091;
  assign n10237 = n4724 & n7648;
  assign n10238 = ~n1426 & n8120;
  assign n10239 = ~n10237 & ~n10238;
  assign n10240 = ~n10236 & n10239;
  assign n10241 = ~n10235 & n10240;
  assign n10242 = ~pi11  & ~n10241;
  assign n10243 = pi11  & n10241;
  assign n10244 = ~n10242 & ~n10243;
  assign n10245 = ~n10143 & n10146;
  assign n10246 = n10143 & ~n10146;
  assign n10247 = ~n10245 & ~n10246;
  assign n10248 = ~n10244 & ~n10247;
  assign n10249 = ~n1740 & n7654;
  assign n10250 = ~n1610 & n8091;
  assign n10251 = n4708 & n7648;
  assign n10252 = ~n1531 & n8120;
  assign n10253 = ~n10251 & ~n10252;
  assign n10254 = ~n10250 & n10253;
  assign n10255 = ~n10249 & n10254;
  assign n10256 = ~pi11  & ~n10255;
  assign n10257 = pi11  & n10255;
  assign n10258 = ~n10256 & ~n10257;
  assign n10259 = ~n10138 & n10141;
  assign n10260 = n10138 & ~n10141;
  assign n10261 = ~n10259 & ~n10260;
  assign n10262 = ~n10258 & ~n10261;
  assign n10263 = ~n1811 & n7654;
  assign n10264 = ~n1740 & n8091;
  assign n10265 = n4951 & n7648;
  assign n10266 = ~n1610 & n8120;
  assign n10267 = ~n10265 & ~n10266;
  assign n10268 = ~n10264 & n10267;
  assign n10269 = ~n10263 & n10268;
  assign n10270 = ~pi11  & ~n10269;
  assign n10271 = pi11  & n10269;
  assign n10272 = ~n10270 & ~n10271;
  assign n10273 = n10133 & n10136;
  assign n10274 = ~n10137 & ~n10273;
  assign n10275 = ~n10272 & n10274;
  assign n10276 = ~n10272 & ~n10274;
  assign n10277 = n10272 & n10274;
  assign n10278 = ~n10276 & ~n10277;
  assign n10279 = ~n1900 & n7654;
  assign n10280 = ~n1811 & n8091;
  assign n10281 = n4967 & n7648;
  assign n10282 = ~n1740 & n8120;
  assign n10283 = ~n10281 & ~n10282;
  assign n10284 = ~n10280 & n10283;
  assign n10285 = ~n10279 & n10284;
  assign n10286 = ~pi11  & ~n10285;
  assign n10287 = pi11  & n10285;
  assign n10288 = ~n10286 & ~n10287;
  assign n10289 = n10128 & n10131;
  assign n10290 = ~n10132 & ~n10289;
  assign n10291 = ~n10288 & n10290;
  assign n10292 = ~n10288 & ~n10290;
  assign n10293 = n10288 & n10290;
  assign n10294 = ~n10292 & ~n10293;
  assign n10295 = ~n2006 & n7654;
  assign n10296 = ~n1900 & n8091;
  assign n10297 = n5344 & n7648;
  assign n10298 = ~n1811 & n8120;
  assign n10299 = ~n10297 & ~n10298;
  assign n10300 = ~n10296 & n10299;
  assign n10301 = ~n10295 & n10300;
  assign n10302 = ~pi11  & ~n10301;
  assign n10303 = pi11  & n10301;
  assign n10304 = ~n10302 & ~n10303;
  assign n10305 = ~n10123 & n10126;
  assign n10306 = n10123 & ~n10126;
  assign n10307 = ~n10305 & ~n10306;
  assign n10308 = ~n10304 & ~n10307;
  assign n10309 = n9837 & n10121;
  assign n10310 = ~n10122 & ~n10309;
  assign n10311 = ~n2058 & n7654;
  assign n10312 = ~n2006 & n8091;
  assign n10313 = n5180 & n7648;
  assign n10314 = ~n1900 & n8120;
  assign n10315 = ~n10313 & ~n10314;
  assign n10316 = ~n10312 & n10315;
  assign n10317 = ~n10311 & n10316;
  assign n10318 = pi11  & n10317;
  assign n10319 = ~pi11  & ~n10317;
  assign n10320 = ~n10318 & ~n10319;
  assign n10321 = n10310 & ~n10320;
  assign n10322 = n9853 & n10119;
  assign n10323 = ~n10120 & ~n10322;
  assign n10324 = ~n2178 & n7654;
  assign n10325 = ~n2058 & n8091;
  assign n10326 = n5554 & n7648;
  assign n10327 = ~n2006 & n8120;
  assign n10328 = ~n10326 & ~n10327;
  assign n10329 = ~n10325 & n10328;
  assign n10330 = ~n10324 & n10329;
  assign n10331 = pi11  & n10330;
  assign n10332 = ~pi11  & ~n10330;
  assign n10333 = ~n10331 & ~n10332;
  assign n10334 = n10323 & ~n10333;
  assign n10335 = ~n2278 & n7654;
  assign n10336 = ~n2178 & n8091;
  assign n10337 = n5538 & n7648;
  assign n10338 = ~n2058 & n8120;
  assign n10339 = ~n10337 & ~n10338;
  assign n10340 = ~n10336 & n10339;
  assign n10341 = ~n10335 & n10340;
  assign n10342 = ~pi11  & ~n10341;
  assign n10343 = pi11  & n10341;
  assign n10344 = ~n10342 & ~n10343;
  assign n10345 = n10115 & ~n10117;
  assign n10346 = ~n10118 & ~n10345;
  assign n10347 = ~n10344 & n10346;
  assign n10348 = ~n10344 & ~n10346;
  assign n10349 = n10344 & n10346;
  assign n10350 = ~n10348 & ~n10349;
  assign n10351 = ~n2369 & n7654;
  assign n10352 = ~n2278 & n8091;
  assign n10353 = n5779 & n7648;
  assign n10354 = ~n2178 & n8120;
  assign n10355 = ~n10353 & ~n10354;
  assign n10356 = ~n10352 & n10355;
  assign n10357 = ~n10351 & n10356;
  assign n10358 = ~pi11  & ~n10357;
  assign n10359 = pi11  & n10357;
  assign n10360 = ~n10358 & ~n10359;
  assign n10361 = ~n10110 & n10113;
  assign n10362 = n10110 & ~n10113;
  assign n10363 = ~n10361 & ~n10362;
  assign n10364 = ~n10360 & ~n10363;
  assign n10365 = ~n2457 & n7654;
  assign n10366 = ~n2369 & n8091;
  assign n10367 = n5795 & n7648;
  assign n10368 = ~n2278 & n8120;
  assign n10369 = ~n10367 & ~n10368;
  assign n10370 = ~n10366 & n10369;
  assign n10371 = ~n10365 & n10370;
  assign n10372 = ~pi11  & ~n10371;
  assign n10373 = pi11  & n10371;
  assign n10374 = ~n10372 & ~n10373;
  assign n10375 = n10105 & n10108;
  assign n10376 = ~n10109 & ~n10375;
  assign n10377 = ~n10374 & n10376;
  assign n10378 = ~n10374 & ~n10376;
  assign n10379 = n10374 & n10376;
  assign n10380 = ~n10378 & ~n10379;
  assign n10381 = n9908 & n10103;
  assign n10382 = ~n10104 & ~n10381;
  assign n10383 = ~n2554 & n7654;
  assign n10384 = ~n2457 & n8091;
  assign n10385 = n6218 & n7648;
  assign n10386 = ~n2369 & n8120;
  assign n10387 = ~n10385 & ~n10386;
  assign n10388 = ~n10384 & n10387;
  assign n10389 = ~n10383 & n10388;
  assign n10390 = pi11  & n10389;
  assign n10391 = ~pi11  & ~n10389;
  assign n10392 = ~n10390 & ~n10391;
  assign n10393 = n10382 & ~n10392;
  assign n10394 = n9924 & n10101;
  assign n10395 = ~n10102 & ~n10394;
  assign n10396 = ~n2640 & n7654;
  assign n10397 = ~n2554 & n8091;
  assign n10398 = n5979 & n7648;
  assign n10399 = ~n2457 & n8120;
  assign n10400 = ~n10398 & ~n10399;
  assign n10401 = ~n10397 & n10400;
  assign n10402 = ~n10396 & n10401;
  assign n10403 = pi11  & n10402;
  assign n10404 = ~pi11  & ~n10402;
  assign n10405 = ~n10403 & ~n10404;
  assign n10406 = n10395 & ~n10405;
  assign n10407 = n10097 & ~n10099;
  assign n10408 = ~n10100 & ~n10407;
  assign n10409 = ~n2676 & n7654;
  assign n10410 = ~n2640 & n8091;
  assign n10411 = n6445 & n7648;
  assign n10412 = ~n2554 & n8120;
  assign n10413 = ~n10411 & ~n10412;
  assign n10414 = ~n10410 & n10413;
  assign n10415 = ~n10409 & n10414;
  assign n10416 = pi11  & n10415;
  assign n10417 = ~pi11  & ~n10415;
  assign n10418 = ~n10416 & ~n10417;
  assign n10419 = n10408 & ~n10418;
  assign n10420 = ~n2748 & n7654;
  assign n10421 = ~n2676 & n8091;
  assign n10422 = n6597 & n7648;
  assign n10423 = ~n2640 & n8120;
  assign n10424 = ~n10422 & ~n10423;
  assign n10425 = ~n10421 & n10424;
  assign n10426 = ~n10420 & n10425;
  assign n10427 = ~pi11  & ~n10426;
  assign n10428 = pi11  & n10426;
  assign n10429 = ~n10427 & ~n10428;
  assign n10430 = n10093 & ~n10095;
  assign n10431 = ~n10096 & ~n10430;
  assign n10432 = ~n10429 & n10431;
  assign n10433 = ~n10429 & ~n10431;
  assign n10434 = n10429 & n10431;
  assign n10435 = ~n10433 & ~n10434;
  assign n10436 = ~n2803 & n7654;
  assign n10437 = ~n2748 & n8091;
  assign n10438 = n6427 & n7648;
  assign n10439 = ~n2676 & n8120;
  assign n10440 = ~n10438 & ~n10439;
  assign n10441 = ~n10437 & n10440;
  assign n10442 = ~n10436 & n10441;
  assign n10443 = ~pi11  & ~n10442;
  assign n10444 = pi11  & n10442;
  assign n10445 = ~n10443 & ~n10444;
  assign n10446 = n10088 & n10091;
  assign n10447 = ~n10092 & ~n10446;
  assign n10448 = ~n10445 & n10447;
  assign n10449 = ~n10445 & ~n10447;
  assign n10450 = n10445 & n10447;
  assign n10451 = ~n10449 & ~n10450;
  assign n10452 = ~n2891 & n7654;
  assign n10453 = ~n2803 & n8091;
  assign n10454 = n6715 & n7648;
  assign n10455 = ~n2748 & n8120;
  assign n10456 = ~n10454 & ~n10455;
  assign n10457 = ~n10453 & n10456;
  assign n10458 = ~n10452 & n10457;
  assign n10459 = ~pi11  & ~n10458;
  assign n10460 = pi11  & n10458;
  assign n10461 = ~n10459 & ~n10460;
  assign n10462 = ~n10083 & n10086;
  assign n10463 = n10083 & ~n10086;
  assign n10464 = ~n10462 & ~n10463;
  assign n10465 = ~n10461 & ~n10464;
  assign n10466 = n9993 & n10081;
  assign n10467 = ~n10082 & ~n10466;
  assign n10468 = ~n2927 & n7654;
  assign n10469 = ~n2891 & n8091;
  assign n10470 = n7014 & n7648;
  assign n10471 = ~n2803 & n8120;
  assign n10472 = ~n10470 & ~n10471;
  assign n10473 = ~n10469 & n10472;
  assign n10474 = ~n10468 & n10473;
  assign n10475 = pi11  & n10474;
  assign n10476 = ~pi11  & ~n10474;
  assign n10477 = ~n10475 & ~n10476;
  assign n10478 = n10467 & ~n10477;
  assign n10479 = n10077 & ~n10079;
  assign n10480 = ~n10080 & ~n10479;
  assign n10481 = ~n3005 & n7654;
  assign n10482 = ~n2927 & n8091;
  assign n10483 = n7026 & n7648;
  assign n10484 = ~n2891 & n8120;
  assign n10485 = ~n10483 & ~n10484;
  assign n10486 = ~n10482 & n10485;
  assign n10487 = ~n10481 & n10486;
  assign n10488 = pi11  & n10487;
  assign n10489 = ~pi11  & ~n10487;
  assign n10490 = ~n10488 & ~n10489;
  assign n10491 = n10480 & ~n10490;
  assign n10492 = n10024 & n10075;
  assign n10493 = ~n10076 & ~n10492;
  assign n10494 = ~n3097 & n7654;
  assign n10495 = ~n3005 & n8091;
  assign n10496 = n6694 & n7648;
  assign n10497 = ~n2927 & n8120;
  assign n10498 = ~n10496 & ~n10497;
  assign n10499 = ~n10495 & n10498;
  assign n10500 = ~n10494 & n10499;
  assign n10501 = pi11  & n10500;
  assign n10502 = ~pi11  & ~n10500;
  assign n10503 = ~n10501 & ~n10502;
  assign n10504 = n10493 & ~n10503;
  assign n10505 = ~n3166 & n7654;
  assign n10506 = ~n3097 & n8091;
  assign n10507 = n7071 & n7648;
  assign n10508 = ~n3005 & n8120;
  assign n10509 = ~n10507 & ~n10508;
  assign n10510 = ~n10506 & n10509;
  assign n10511 = ~n10505 & n10510;
  assign n10512 = ~pi11  & ~n10511;
  assign n10513 = pi11  & n10511;
  assign n10514 = ~n10512 & ~n10513;
  assign n10515 = n10071 & ~n10073;
  assign n10516 = ~n10074 & ~n10515;
  assign n10517 = ~n10514 & n10516;
  assign n10518 = ~n10514 & ~n10516;
  assign n10519 = n10514 & n10516;
  assign n10520 = ~n10518 & ~n10519;
  assign n10521 = ~n3226 & n7654;
  assign n10522 = ~n3166 & n8091;
  assign n10523 = n7121 & n7648;
  assign n10524 = ~n3097 & n8120;
  assign n10525 = ~n10523 & ~n10524;
  assign n10526 = ~n10522 & n10525;
  assign n10527 = ~n10521 & n10526;
  assign n10528 = pi11  & n10527;
  assign n10529 = ~pi11  & ~n10527;
  assign n10530 = ~n10528 & ~n10529;
  assign n10531 = n10059 & n10069;
  assign n10532 = ~n10070 & ~n10531;
  assign n10533 = ~n10530 & n10532;
  assign n10534 = ~n3263 & n7654;
  assign n10535 = ~n3226 & n8091;
  assign n10536 = n7175 & n7648;
  assign n10537 = ~n3166 & n8120;
  assign n10538 = ~n10536 & ~n10537;
  assign n10539 = ~n10535 & n10538;
  assign n10540 = ~n10534 & n10539;
  assign n10541 = ~pi11  & ~n10540;
  assign n10542 = pi11  & n10540;
  assign n10543 = ~n10541 & ~n10542;
  assign n10544 = pi14  & ~n10047;
  assign n10545 = n10054 & ~n10544;
  assign n10546 = ~n10054 & n10544;
  assign n10547 = ~n10545 & ~n10546;
  assign n10548 = ~n10543 & n10547;
  assign n10549 = ~n10543 & ~n10547;
  assign n10550 = n10543 & n10547;
  assign n10551 = ~n10549 & ~n10550;
  assign n10552 = ~n3360 & n7654;
  assign n10553 = ~n3263 & n8091;
  assign n10554 = n7221 & n7648;
  assign n10555 = ~n3226 & n8120;
  assign n10556 = ~n10554 & ~n10555;
  assign n10557 = ~n10553 & n10556;
  assign n10558 = ~n10552 & n10557;
  assign n10559 = pi11  & n10558;
  assign n10560 = ~pi11  & ~n10558;
  assign n10561 = ~n10559 & ~n10560;
  assign n10562 = pi14  & n10045;
  assign n10563 = ~n10044 & n10562;
  assign n10564 = n10044 & ~n10562;
  assign n10565 = ~n10563 & ~n10564;
  assign n10566 = ~n10561 & n10565;
  assign n10567 = n7648 & ~n7942;
  assign n10568 = ~n3506 & n8120;
  assign n10569 = ~n3450 & n8091;
  assign n10570 = ~n10568 & ~n10569;
  assign n10571 = ~n10567 & n10570;
  assign n10572 = ~n3450 & ~n7644;
  assign n10573 = pi11  & ~n10572;
  assign n10574 = n10571 & n10573;
  assign n10575 = ~n3450 & n7654;
  assign n10576 = ~n3506 & n8091;
  assign n10577 = n7265 & n7648;
  assign n10578 = ~n3360 & n8120;
  assign n10579 = ~n10577 & ~n10578;
  assign n10580 = ~n10576 & n10579;
  assign n10581 = ~n10575 & n10580;
  assign n10582 = n10574 & n10581;
  assign n10583 = n10045 & n10582;
  assign n10584 = ~n10045 & n10582;
  assign n10585 = n10045 & ~n10582;
  assign n10586 = ~n10584 & ~n10585;
  assign n10587 = ~n3506 & n7654;
  assign n10588 = ~n3360 & n8091;
  assign n10589 = n7323 & n7648;
  assign n10590 = ~n3263 & n8120;
  assign n10591 = ~n10589 & ~n10590;
  assign n10592 = ~n10588 & n10591;
  assign n10593 = ~n10587 & n10592;
  assign n10594 = pi11  & n10593;
  assign n10595 = ~pi11  & ~n10593;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = ~n10586 & ~n10596;
  assign n10598 = ~n10583 & ~n10597;
  assign n10599 = n10561 & ~n10565;
  assign n10600 = ~n10566 & ~n10599;
  assign n10601 = ~n10598 & n10600;
  assign n10602 = ~n10566 & ~n10601;
  assign n10603 = ~n10551 & ~n10602;
  assign n10604 = ~n10548 & ~n10603;
  assign n10605 = n10530 & ~n10532;
  assign n10606 = ~n10533 & ~n10605;
  assign n10607 = ~n10604 & n10606;
  assign n10608 = ~n10533 & ~n10607;
  assign n10609 = ~n10520 & ~n10608;
  assign n10610 = ~n10517 & ~n10609;
  assign n10611 = n10493 & n10503;
  assign n10612 = ~n10493 & ~n10503;
  assign n10613 = ~n10611 & ~n10612;
  assign n10614 = ~n10610 & ~n10613;
  assign n10615 = ~n10504 & ~n10614;
  assign n10616 = n10480 & n10490;
  assign n10617 = ~n10480 & ~n10490;
  assign n10618 = ~n10616 & ~n10617;
  assign n10619 = ~n10615 & ~n10618;
  assign n10620 = ~n10491 & ~n10619;
  assign n10621 = ~n10467 & n10477;
  assign n10622 = ~n10478 & ~n10621;
  assign n10623 = ~n10620 & n10622;
  assign n10624 = ~n10478 & ~n10623;
  assign n10625 = n10461 & n10464;
  assign n10626 = ~n10465 & ~n10625;
  assign n10627 = ~n10624 & n10626;
  assign n10628 = ~n10465 & ~n10627;
  assign n10629 = ~n10451 & ~n10628;
  assign n10630 = ~n10448 & ~n10629;
  assign n10631 = ~n10435 & ~n10630;
  assign n10632 = ~n10432 & ~n10631;
  assign n10633 = n10408 & n10418;
  assign n10634 = ~n10408 & ~n10418;
  assign n10635 = ~n10633 & ~n10634;
  assign n10636 = ~n10632 & ~n10635;
  assign n10637 = ~n10419 & ~n10636;
  assign n10638 = n10395 & n10405;
  assign n10639 = ~n10395 & ~n10405;
  assign n10640 = ~n10638 & ~n10639;
  assign n10641 = ~n10637 & ~n10640;
  assign n10642 = ~n10406 & ~n10641;
  assign n10643 = ~n10382 & n10392;
  assign n10644 = ~n10393 & ~n10643;
  assign n10645 = ~n10642 & n10644;
  assign n10646 = ~n10393 & ~n10645;
  assign n10647 = ~n10380 & ~n10646;
  assign n10648 = ~n10377 & ~n10647;
  assign n10649 = n10360 & n10363;
  assign n10650 = ~n10364 & ~n10649;
  assign n10651 = ~n10648 & n10650;
  assign n10652 = ~n10364 & ~n10651;
  assign n10653 = ~n10350 & ~n10652;
  assign n10654 = ~n10347 & ~n10653;
  assign n10655 = n10323 & n10333;
  assign n10656 = ~n10323 & ~n10333;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = ~n10654 & ~n10657;
  assign n10659 = ~n10334 & ~n10658;
  assign n10660 = ~n10310 & n10320;
  assign n10661 = ~n10321 & ~n10660;
  assign n10662 = ~n10659 & n10661;
  assign n10663 = ~n10321 & ~n10662;
  assign n10664 = n10304 & n10307;
  assign n10665 = ~n10308 & ~n10664;
  assign n10666 = ~n10663 & n10665;
  assign n10667 = ~n10308 & ~n10666;
  assign n10668 = ~n10294 & ~n10667;
  assign n10669 = ~n10291 & ~n10668;
  assign n10670 = ~n10278 & ~n10669;
  assign n10671 = ~n10275 & ~n10670;
  assign n10672 = n10258 & n10261;
  assign n10673 = ~n10262 & ~n10672;
  assign n10674 = ~n10671 & n10673;
  assign n10675 = ~n10262 & ~n10674;
  assign n10676 = n10244 & n10247;
  assign n10677 = ~n10248 & ~n10676;
  assign n10678 = ~n10675 & n10677;
  assign n10679 = ~n10248 & ~n10678;
  assign n10680 = ~n10234 & ~n10679;
  assign n10681 = ~n10231 & ~n10680;
  assign n10682 = ~n10218 & ~n10681;
  assign n10683 = ~n10215 & ~n10682;
  assign n10684 = n10171 & ~n10173;
  assign n10685 = ~n10174 & ~n10684;
  assign n10686 = ~n10683 & n10685;
  assign n10687 = ~n1005 & n8474;
  assign n10688 = ~n894 & n9238;
  assign n10689 = n4122 & n8468;
  assign n10690 = ~n795 & n9265;
  assign n10691 = ~n10689 & ~n10690;
  assign n10692 = ~n10688 & n10691;
  assign n10693 = ~n10687 & n10692;
  assign n10694 = ~pi8  & ~n10693;
  assign n10695 = pi8  & n10693;
  assign n10696 = ~n10694 & ~n10695;
  assign n10697 = n10683 & ~n10685;
  assign n10698 = ~n10686 & ~n10697;
  assign n10699 = ~n10696 & n10698;
  assign n10700 = ~n10686 & ~n10699;
  assign n10701 = ~n3744 & n9719;
  assign n10702 = n9715 & ~n9723;
  assign n10703 = ~n554 & n10702;
  assign n10704 = ~n720 & n9725;
  assign n10705 = ~n10703 & ~n10704;
  assign n10706 = ~n10701 & n10705;
  assign n10707 = pi5  & n10706;
  assign n10708 = ~pi5  & ~n10706;
  assign n10709 = ~n10707 & ~n10708;
  assign n10710 = ~n10700 & ~n10709;
  assign n10711 = n10700 & n10709;
  assign n10712 = ~n10710 & ~n10711;
  assign n10713 = ~n10180 & ~n10181;
  assign n10714 = ~n10191 & n10713;
  assign n10715 = n10191 & ~n10713;
  assign n10716 = ~n10714 & ~n10715;
  assign n10717 = n10712 & n10716;
  assign n10718 = ~n10710 & ~n10717;
  assign n10719 = ~n10194 & ~n10195;
  assign n10720 = n10199 & n10719;
  assign n10721 = ~n10199 & ~n10719;
  assign n10722 = ~n10720 & ~n10721;
  assign n10723 = ~n10718 & n10722;
  assign n10724 = n10718 & ~n10722;
  assign n10725 = ~n10723 & ~n10724;
  assign n10726 = n10218 & n10681;
  assign n10727 = ~n10682 & ~n10726;
  assign n10728 = ~n1107 & n8474;
  assign n10729 = ~n1005 & n9238;
  assign n10730 = n4106 & n8468;
  assign n10731 = ~n894 & n9265;
  assign n10732 = ~n10730 & ~n10731;
  assign n10733 = ~n10729 & n10732;
  assign n10734 = ~n10728 & n10733;
  assign n10735 = pi8  & n10734;
  assign n10736 = ~pi8  & ~n10734;
  assign n10737 = ~n10735 & ~n10736;
  assign n10738 = n10727 & ~n10737;
  assign n10739 = n10234 & n10679;
  assign n10740 = ~n10680 & ~n10739;
  assign n10741 = ~n1230 & n8474;
  assign n10742 = ~n1107 & n9238;
  assign n10743 = n4307 & n8468;
  assign n10744 = ~n1005 & n9265;
  assign n10745 = ~n10743 & ~n10744;
  assign n10746 = ~n10742 & n10745;
  assign n10747 = ~n10741 & n10746;
  assign n10748 = pi8  & n10747;
  assign n10749 = ~pi8  & ~n10747;
  assign n10750 = ~n10748 & ~n10749;
  assign n10751 = n10740 & ~n10750;
  assign n10752 = n10675 & ~n10677;
  assign n10753 = ~n10678 & ~n10752;
  assign n10754 = ~n1338 & n8474;
  assign n10755 = ~n1230 & n9238;
  assign n10756 = n4323 & n8468;
  assign n10757 = ~n1107 & n9265;
  assign n10758 = ~n10756 & ~n10757;
  assign n10759 = ~n10755 & n10758;
  assign n10760 = ~n10754 & n10759;
  assign n10761 = pi8  & n10760;
  assign n10762 = ~pi8  & ~n10760;
  assign n10763 = ~n10761 & ~n10762;
  assign n10764 = n10753 & ~n10763;
  assign n10765 = n10671 & ~n10673;
  assign n10766 = ~n10674 & ~n10765;
  assign n10767 = ~n1426 & n8474;
  assign n10768 = ~n1338 & n9238;
  assign n10769 = n4753 & n8468;
  assign n10770 = ~n1230 & n9265;
  assign n10771 = ~n10769 & ~n10770;
  assign n10772 = ~n10768 & n10771;
  assign n10773 = ~n10767 & n10772;
  assign n10774 = pi8  & n10773;
  assign n10775 = ~pi8  & ~n10773;
  assign n10776 = ~n10774 & ~n10775;
  assign n10777 = n10766 & ~n10776;
  assign n10778 = n10278 & n10669;
  assign n10779 = ~n10670 & ~n10778;
  assign n10780 = ~n1531 & n8474;
  assign n10781 = ~n1426 & n9238;
  assign n10782 = n4533 & n8468;
  assign n10783 = ~n1338 & n9265;
  assign n10784 = ~n10782 & ~n10783;
  assign n10785 = ~n10781 & n10784;
  assign n10786 = ~n10780 & n10785;
  assign n10787 = pi8  & n10786;
  assign n10788 = ~pi8  & ~n10786;
  assign n10789 = ~n10787 & ~n10788;
  assign n10790 = n10779 & ~n10789;
  assign n10791 = n10294 & n10667;
  assign n10792 = ~n10668 & ~n10791;
  assign n10793 = ~n1610 & n8474;
  assign n10794 = ~n1531 & n9238;
  assign n10795 = n4724 & n8468;
  assign n10796 = ~n1426 & n9265;
  assign n10797 = ~n10795 & ~n10796;
  assign n10798 = ~n10794 & n10797;
  assign n10799 = ~n10793 & n10798;
  assign n10800 = pi8  & n10799;
  assign n10801 = ~pi8  & ~n10799;
  assign n10802 = ~n10800 & ~n10801;
  assign n10803 = n10792 & ~n10802;
  assign n10804 = n10663 & ~n10665;
  assign n10805 = ~n10666 & ~n10804;
  assign n10806 = ~n1740 & n8474;
  assign n10807 = ~n1610 & n9238;
  assign n10808 = n4708 & n8468;
  assign n10809 = ~n1531 & n9265;
  assign n10810 = ~n10808 & ~n10809;
  assign n10811 = ~n10807 & n10810;
  assign n10812 = ~n10806 & n10811;
  assign n10813 = pi8  & n10812;
  assign n10814 = ~pi8  & ~n10812;
  assign n10815 = ~n10813 & ~n10814;
  assign n10816 = n10805 & ~n10815;
  assign n10817 = ~n1811 & n8474;
  assign n10818 = ~n1740 & n9238;
  assign n10819 = n4951 & n8468;
  assign n10820 = ~n1610 & n9265;
  assign n10821 = ~n10819 & ~n10820;
  assign n10822 = ~n10818 & n10821;
  assign n10823 = ~n10817 & n10822;
  assign n10824 = ~pi8  & ~n10823;
  assign n10825 = pi8  & n10823;
  assign n10826 = ~n10824 & ~n10825;
  assign n10827 = n10659 & ~n10661;
  assign n10828 = ~n10662 & ~n10827;
  assign n10829 = ~n10826 & n10828;
  assign n10830 = ~n10826 & ~n10828;
  assign n10831 = n10826 & n10828;
  assign n10832 = ~n10830 & ~n10831;
  assign n10833 = ~n1900 & n8474;
  assign n10834 = ~n1811 & n9238;
  assign n10835 = n4967 & n8468;
  assign n10836 = ~n1740 & n9265;
  assign n10837 = ~n10835 & ~n10836;
  assign n10838 = ~n10834 & n10837;
  assign n10839 = ~n10833 & n10838;
  assign n10840 = ~pi8  & ~n10839;
  assign n10841 = pi8  & n10839;
  assign n10842 = ~n10840 & ~n10841;
  assign n10843 = ~n10654 & n10657;
  assign n10844 = n10654 & ~n10657;
  assign n10845 = ~n10843 & ~n10844;
  assign n10846 = ~n10842 & ~n10845;
  assign n10847 = n10350 & n10652;
  assign n10848 = ~n10653 & ~n10847;
  assign n10849 = ~n2006 & n8474;
  assign n10850 = ~n1900 & n9238;
  assign n10851 = n5344 & n8468;
  assign n10852 = ~n1811 & n9265;
  assign n10853 = ~n10851 & ~n10852;
  assign n10854 = ~n10850 & n10853;
  assign n10855 = ~n10849 & n10854;
  assign n10856 = pi8  & n10855;
  assign n10857 = ~pi8  & ~n10855;
  assign n10858 = ~n10856 & ~n10857;
  assign n10859 = n10848 & ~n10858;
  assign n10860 = n10648 & ~n10650;
  assign n10861 = ~n10651 & ~n10860;
  assign n10862 = ~n2058 & n8474;
  assign n10863 = ~n2006 & n9238;
  assign n10864 = n5180 & n8468;
  assign n10865 = ~n1900 & n9265;
  assign n10866 = ~n10864 & ~n10865;
  assign n10867 = ~n10863 & n10866;
  assign n10868 = ~n10862 & n10867;
  assign n10869 = pi8  & n10868;
  assign n10870 = ~pi8  & ~n10868;
  assign n10871 = ~n10869 & ~n10870;
  assign n10872 = n10861 & ~n10871;
  assign n10873 = n10380 & n10646;
  assign n10874 = ~n10647 & ~n10873;
  assign n10875 = ~n2178 & n8474;
  assign n10876 = ~n2058 & n9238;
  assign n10877 = n5554 & n8468;
  assign n10878 = ~n2006 & n9265;
  assign n10879 = ~n10877 & ~n10878;
  assign n10880 = ~n10876 & n10879;
  assign n10881 = ~n10875 & n10880;
  assign n10882 = pi8  & n10881;
  assign n10883 = ~pi8  & ~n10881;
  assign n10884 = ~n10882 & ~n10883;
  assign n10885 = n10874 & ~n10884;
  assign n10886 = ~n2278 & n8474;
  assign n10887 = ~n2178 & n9238;
  assign n10888 = n5538 & n8468;
  assign n10889 = ~n2058 & n9265;
  assign n10890 = ~n10888 & ~n10889;
  assign n10891 = ~n10887 & n10890;
  assign n10892 = ~n10886 & n10891;
  assign n10893 = ~pi8  & ~n10892;
  assign n10894 = pi8  & n10892;
  assign n10895 = ~n10893 & ~n10894;
  assign n10896 = n10642 & ~n10644;
  assign n10897 = ~n10645 & ~n10896;
  assign n10898 = ~n10895 & n10897;
  assign n10899 = ~n10895 & ~n10897;
  assign n10900 = n10895 & n10897;
  assign n10901 = ~n10899 & ~n10900;
  assign n10902 = ~n2369 & n8474;
  assign n10903 = ~n2278 & n9238;
  assign n10904 = n5779 & n8468;
  assign n10905 = ~n2178 & n9265;
  assign n10906 = ~n10904 & ~n10905;
  assign n10907 = ~n10903 & n10906;
  assign n10908 = ~n10902 & n10907;
  assign n10909 = ~pi8  & ~n10908;
  assign n10910 = pi8  & n10908;
  assign n10911 = ~n10909 & ~n10910;
  assign n10912 = ~n10637 & n10640;
  assign n10913 = n10637 & ~n10640;
  assign n10914 = ~n10912 & ~n10913;
  assign n10915 = ~n10911 & ~n10914;
  assign n10916 = ~n2457 & n8474;
  assign n10917 = ~n2369 & n9238;
  assign n10918 = n5795 & n8468;
  assign n10919 = ~n2278 & n9265;
  assign n10920 = ~n10918 & ~n10919;
  assign n10921 = ~n10917 & n10920;
  assign n10922 = ~n10916 & n10921;
  assign n10923 = ~pi8  & ~n10922;
  assign n10924 = pi8  & n10922;
  assign n10925 = ~n10923 & ~n10924;
  assign n10926 = n10632 & n10635;
  assign n10927 = ~n10636 & ~n10926;
  assign n10928 = ~n10925 & n10927;
  assign n10929 = ~n10925 & ~n10927;
  assign n10930 = n10925 & n10927;
  assign n10931 = ~n10929 & ~n10930;
  assign n10932 = n10435 & n10630;
  assign n10933 = ~n10631 & ~n10932;
  assign n10934 = ~n2554 & n8474;
  assign n10935 = ~n2457 & n9238;
  assign n10936 = n6218 & n8468;
  assign n10937 = ~n2369 & n9265;
  assign n10938 = ~n10936 & ~n10937;
  assign n10939 = ~n10935 & n10938;
  assign n10940 = ~n10934 & n10939;
  assign n10941 = pi8  & n10940;
  assign n10942 = ~pi8  & ~n10940;
  assign n10943 = ~n10941 & ~n10942;
  assign n10944 = n10933 & ~n10943;
  assign n10945 = n10451 & n10628;
  assign n10946 = ~n10629 & ~n10945;
  assign n10947 = ~n2640 & n8474;
  assign n10948 = ~n2554 & n9238;
  assign n10949 = n5979 & n8468;
  assign n10950 = ~n2457 & n9265;
  assign n10951 = ~n10949 & ~n10950;
  assign n10952 = ~n10948 & n10951;
  assign n10953 = ~n10947 & n10952;
  assign n10954 = pi8  & n10953;
  assign n10955 = ~pi8  & ~n10953;
  assign n10956 = ~n10954 & ~n10955;
  assign n10957 = n10946 & ~n10956;
  assign n10958 = n10624 & ~n10626;
  assign n10959 = ~n10627 & ~n10958;
  assign n10960 = ~n2676 & n8474;
  assign n10961 = ~n2640 & n9238;
  assign n10962 = n6445 & n8468;
  assign n10963 = ~n2554 & n9265;
  assign n10964 = ~n10962 & ~n10963;
  assign n10965 = ~n10961 & n10964;
  assign n10966 = ~n10960 & n10965;
  assign n10967 = pi8  & n10966;
  assign n10968 = ~pi8  & ~n10966;
  assign n10969 = ~n10967 & ~n10968;
  assign n10970 = n10959 & ~n10969;
  assign n10971 = ~n2748 & n8474;
  assign n10972 = ~n2676 & n9238;
  assign n10973 = n6597 & n8468;
  assign n10974 = ~n2640 & n9265;
  assign n10975 = ~n10973 & ~n10974;
  assign n10976 = ~n10972 & n10975;
  assign n10977 = ~n10971 & n10976;
  assign n10978 = ~pi8  & ~n10977;
  assign n10979 = pi8  & n10977;
  assign n10980 = ~n10978 & ~n10979;
  assign n10981 = n10620 & ~n10622;
  assign n10982 = ~n10623 & ~n10981;
  assign n10983 = ~n10980 & n10982;
  assign n10984 = ~n10980 & ~n10982;
  assign n10985 = n10980 & n10982;
  assign n10986 = ~n10984 & ~n10985;
  assign n10987 = ~n2803 & n8474;
  assign n10988 = ~n2748 & n9238;
  assign n10989 = n6427 & n8468;
  assign n10990 = ~n2676 & n9265;
  assign n10991 = ~n10989 & ~n10990;
  assign n10992 = ~n10988 & n10991;
  assign n10993 = ~n10987 & n10992;
  assign n10994 = ~pi8  & ~n10993;
  assign n10995 = pi8  & n10993;
  assign n10996 = ~n10994 & ~n10995;
  assign n10997 = n10615 & n10618;
  assign n10998 = ~n10619 & ~n10997;
  assign n10999 = ~n10996 & n10998;
  assign n11000 = ~n10996 & ~n10998;
  assign n11001 = n10996 & n10998;
  assign n11002 = ~n11000 & ~n11001;
  assign n11003 = ~n2891 & n8474;
  assign n11004 = ~n2803 & n9238;
  assign n11005 = n6715 & n8468;
  assign n11006 = ~n2748 & n9265;
  assign n11007 = ~n11005 & ~n11006;
  assign n11008 = ~n11004 & n11007;
  assign n11009 = ~n11003 & n11008;
  assign n11010 = ~pi8  & ~n11009;
  assign n11011 = pi8  & n11009;
  assign n11012 = ~n11010 & ~n11011;
  assign n11013 = ~n10610 & n10613;
  assign n11014 = n10610 & ~n10613;
  assign n11015 = ~n11013 & ~n11014;
  assign n11016 = ~n11012 & ~n11015;
  assign n11017 = n10520 & n10608;
  assign n11018 = ~n10609 & ~n11017;
  assign n11019 = ~n2927 & n8474;
  assign n11020 = ~n2891 & n9238;
  assign n11021 = n7014 & n8468;
  assign n11022 = ~n2803 & n9265;
  assign n11023 = ~n11021 & ~n11022;
  assign n11024 = ~n11020 & n11023;
  assign n11025 = ~n11019 & n11024;
  assign n11026 = pi8  & n11025;
  assign n11027 = ~pi8  & ~n11025;
  assign n11028 = ~n11026 & ~n11027;
  assign n11029 = n11018 & ~n11028;
  assign n11030 = n10604 & ~n10606;
  assign n11031 = ~n10607 & ~n11030;
  assign n11032 = ~n3005 & n8474;
  assign n11033 = ~n2927 & n9238;
  assign n11034 = n7026 & n8468;
  assign n11035 = ~n2891 & n9265;
  assign n11036 = ~n11034 & ~n11035;
  assign n11037 = ~n11033 & n11036;
  assign n11038 = ~n11032 & n11037;
  assign n11039 = pi8  & n11038;
  assign n11040 = ~pi8  & ~n11038;
  assign n11041 = ~n11039 & ~n11040;
  assign n11042 = n11031 & ~n11041;
  assign n11043 = n10551 & n10602;
  assign n11044 = ~n10603 & ~n11043;
  assign n11045 = ~n3097 & n8474;
  assign n11046 = ~n3005 & n9238;
  assign n11047 = n6694 & n8468;
  assign n11048 = ~n2927 & n9265;
  assign n11049 = ~n11047 & ~n11048;
  assign n11050 = ~n11046 & n11049;
  assign n11051 = ~n11045 & n11050;
  assign n11052 = pi8  & n11051;
  assign n11053 = ~pi8  & ~n11051;
  assign n11054 = ~n11052 & ~n11053;
  assign n11055 = n11044 & ~n11054;
  assign n11056 = ~n3166 & n8474;
  assign n11057 = ~n3097 & n9238;
  assign n11058 = n7071 & n8468;
  assign n11059 = ~n3005 & n9265;
  assign n11060 = ~n11058 & ~n11059;
  assign n11061 = ~n11057 & n11060;
  assign n11062 = ~n11056 & n11061;
  assign n11063 = ~pi8  & ~n11062;
  assign n11064 = pi8  & n11062;
  assign n11065 = ~n11063 & ~n11064;
  assign n11066 = n10598 & ~n10600;
  assign n11067 = ~n10601 & ~n11066;
  assign n11068 = ~n11065 & n11067;
  assign n11069 = ~n11065 & ~n11067;
  assign n11070 = n11065 & n11067;
  assign n11071 = ~n11069 & ~n11070;
  assign n11072 = ~n3226 & n8474;
  assign n11073 = ~n3166 & n9238;
  assign n11074 = n7121 & n8468;
  assign n11075 = ~n3097 & n9265;
  assign n11076 = ~n11074 & ~n11075;
  assign n11077 = ~n11073 & n11076;
  assign n11078 = ~n11072 & n11077;
  assign n11079 = pi8  & n11078;
  assign n11080 = ~pi8  & ~n11078;
  assign n11081 = ~n11079 & ~n11080;
  assign n11082 = n10586 & n10596;
  assign n11083 = ~n10597 & ~n11082;
  assign n11084 = ~n11081 & n11083;
  assign n11085 = ~n3263 & n8474;
  assign n11086 = ~n3226 & n9238;
  assign n11087 = n7175 & n8468;
  assign n11088 = ~n3166 & n9265;
  assign n11089 = ~n11087 & ~n11088;
  assign n11090 = ~n11086 & n11089;
  assign n11091 = ~n11085 & n11090;
  assign n11092 = ~pi8  & ~n11091;
  assign n11093 = pi8  & n11091;
  assign n11094 = ~n11092 & ~n11093;
  assign n11095 = pi11  & ~n10574;
  assign n11096 = n10581 & ~n11095;
  assign n11097 = ~n10581 & n11095;
  assign n11098 = ~n11096 & ~n11097;
  assign n11099 = ~n11094 & n11098;
  assign n11100 = ~n11094 & ~n11098;
  assign n11101 = n11094 & n11098;
  assign n11102 = ~n11100 & ~n11101;
  assign n11103 = ~n3360 & n8474;
  assign n11104 = ~n3263 & n9238;
  assign n11105 = n7221 & n8468;
  assign n11106 = ~n3226 & n9265;
  assign n11107 = ~n11105 & ~n11106;
  assign n11108 = ~n11104 & n11107;
  assign n11109 = ~n11103 & n11108;
  assign n11110 = pi8  & n11109;
  assign n11111 = ~pi8  & ~n11109;
  assign n11112 = ~n11110 & ~n11111;
  assign n11113 = pi11  & n10572;
  assign n11114 = ~n10571 & n11113;
  assign n11115 = n10571 & ~n11113;
  assign n11116 = ~n11114 & ~n11115;
  assign n11117 = ~n11112 & n11116;
  assign n11118 = ~n7942 & n8468;
  assign n11119 = ~n3506 & n9265;
  assign n11120 = ~n3450 & n9238;
  assign n11121 = ~n11119 & ~n11120;
  assign n11122 = ~n11118 & n11121;
  assign n11123 = ~n3450 & ~n8464;
  assign n11124 = pi8  & ~n11123;
  assign n11125 = n11122 & n11124;
  assign n11126 = ~n3450 & n8474;
  assign n11127 = ~n3506 & n9238;
  assign n11128 = n7265 & n8468;
  assign n11129 = ~n3360 & n9265;
  assign n11130 = ~n11128 & ~n11129;
  assign n11131 = ~n11127 & n11130;
  assign n11132 = ~n11126 & n11131;
  assign n11133 = n11125 & n11132;
  assign n11134 = n10572 & n11133;
  assign n11135 = ~n10572 & n11133;
  assign n11136 = n10572 & ~n11133;
  assign n11137 = ~n11135 & ~n11136;
  assign n11138 = ~n3506 & n8474;
  assign n11139 = ~n3360 & n9238;
  assign n11140 = n7323 & n8468;
  assign n11141 = ~n3263 & n9265;
  assign n11142 = ~n11140 & ~n11141;
  assign n11143 = ~n11139 & n11142;
  assign n11144 = ~n11138 & n11143;
  assign n11145 = pi8  & n11144;
  assign n11146 = ~pi8  & ~n11144;
  assign n11147 = ~n11145 & ~n11146;
  assign n11148 = ~n11137 & ~n11147;
  assign n11149 = ~n11134 & ~n11148;
  assign n11150 = n11112 & ~n11116;
  assign n11151 = ~n11117 & ~n11150;
  assign n11152 = ~n11149 & n11151;
  assign n11153 = ~n11117 & ~n11152;
  assign n11154 = ~n11102 & ~n11153;
  assign n11155 = ~n11099 & ~n11154;
  assign n11156 = n11081 & ~n11083;
  assign n11157 = ~n11084 & ~n11156;
  assign n11158 = ~n11155 & n11157;
  assign n11159 = ~n11084 & ~n11158;
  assign n11160 = ~n11071 & ~n11159;
  assign n11161 = ~n11068 & ~n11160;
  assign n11162 = n11044 & n11054;
  assign n11163 = ~n11044 & ~n11054;
  assign n11164 = ~n11162 & ~n11163;
  assign n11165 = ~n11161 & ~n11164;
  assign n11166 = ~n11055 & ~n11165;
  assign n11167 = n11031 & n11041;
  assign n11168 = ~n11031 & ~n11041;
  assign n11169 = ~n11167 & ~n11168;
  assign n11170 = ~n11166 & ~n11169;
  assign n11171 = ~n11042 & ~n11170;
  assign n11172 = ~n11018 & n11028;
  assign n11173 = ~n11029 & ~n11172;
  assign n11174 = ~n11171 & n11173;
  assign n11175 = ~n11029 & ~n11174;
  assign n11176 = n11012 & n11015;
  assign n11177 = ~n11016 & ~n11176;
  assign n11178 = ~n11175 & n11177;
  assign n11179 = ~n11016 & ~n11178;
  assign n11180 = ~n11002 & ~n11179;
  assign n11181 = ~n10999 & ~n11180;
  assign n11182 = ~n10986 & ~n11181;
  assign n11183 = ~n10983 & ~n11182;
  assign n11184 = n10959 & n10969;
  assign n11185 = ~n10959 & ~n10969;
  assign n11186 = ~n11184 & ~n11185;
  assign n11187 = ~n11183 & ~n11186;
  assign n11188 = ~n10970 & ~n11187;
  assign n11189 = n10946 & n10956;
  assign n11190 = ~n10946 & ~n10956;
  assign n11191 = ~n11189 & ~n11190;
  assign n11192 = ~n11188 & ~n11191;
  assign n11193 = ~n10957 & ~n11192;
  assign n11194 = ~n10933 & n10943;
  assign n11195 = ~n10944 & ~n11194;
  assign n11196 = ~n11193 & n11195;
  assign n11197 = ~n10944 & ~n11196;
  assign n11198 = ~n10931 & ~n11197;
  assign n11199 = ~n10928 & ~n11198;
  assign n11200 = n10911 & n10914;
  assign n11201 = ~n10915 & ~n11200;
  assign n11202 = ~n11199 & n11201;
  assign n11203 = ~n10915 & ~n11202;
  assign n11204 = ~n10901 & ~n11203;
  assign n11205 = ~n10898 & ~n11204;
  assign n11206 = n10874 & n10884;
  assign n11207 = ~n10874 & ~n10884;
  assign n11208 = ~n11206 & ~n11207;
  assign n11209 = ~n11205 & ~n11208;
  assign n11210 = ~n10885 & ~n11209;
  assign n11211 = n10861 & n10871;
  assign n11212 = ~n10861 & ~n10871;
  assign n11213 = ~n11211 & ~n11212;
  assign n11214 = ~n11210 & ~n11213;
  assign n11215 = ~n10872 & ~n11214;
  assign n11216 = ~n10848 & n10858;
  assign n11217 = ~n10859 & ~n11216;
  assign n11218 = ~n11215 & n11217;
  assign n11219 = ~n10859 & ~n11218;
  assign n11220 = n10842 & n10845;
  assign n11221 = ~n10846 & ~n11220;
  assign n11222 = ~n11219 & n11221;
  assign n11223 = ~n10846 & ~n11222;
  assign n11224 = ~n10832 & ~n11223;
  assign n11225 = ~n10829 & ~n11224;
  assign n11226 = n10805 & n10815;
  assign n11227 = ~n10805 & ~n10815;
  assign n11228 = ~n11226 & ~n11227;
  assign n11229 = ~n11225 & ~n11228;
  assign n11230 = ~n10816 & ~n11229;
  assign n11231 = n10792 & n10802;
  assign n11232 = ~n10792 & ~n10802;
  assign n11233 = ~n11231 & ~n11232;
  assign n11234 = ~n11230 & ~n11233;
  assign n11235 = ~n10803 & ~n11234;
  assign n11236 = n10779 & n10789;
  assign n11237 = ~n10779 & ~n10789;
  assign n11238 = ~n11236 & ~n11237;
  assign n11239 = ~n11235 & ~n11238;
  assign n11240 = ~n10790 & ~n11239;
  assign n11241 = n10766 & n10776;
  assign n11242 = ~n10766 & ~n10776;
  assign n11243 = ~n11241 & ~n11242;
  assign n11244 = ~n11240 & ~n11243;
  assign n11245 = ~n10777 & ~n11244;
  assign n11246 = n10753 & n10763;
  assign n11247 = ~n10753 & ~n10763;
  assign n11248 = ~n11246 & ~n11247;
  assign n11249 = ~n11245 & ~n11248;
  assign n11250 = ~n10764 & ~n11249;
  assign n11251 = n10740 & n10750;
  assign n11252 = ~n10740 & ~n10750;
  assign n11253 = ~n11251 & ~n11252;
  assign n11254 = ~n11250 & ~n11253;
  assign n11255 = ~n10751 & ~n11254;
  assign n11256 = n10727 & n10737;
  assign n11257 = ~n10727 & ~n10737;
  assign n11258 = ~n11256 & ~n11257;
  assign n11259 = ~n11255 & ~n11258;
  assign n11260 = ~n10738 & ~n11259;
  assign n11261 = n10696 & ~n10698;
  assign n11262 = ~n10699 & ~n11261;
  assign n11263 = ~n11260 & n11262;
  assign n11264 = ~n665 & n9725;
  assign n11265 = ~n720 & n10702;
  assign n11266 = n3979 & n9719;
  assign n11267 = ~n9715 & n9718;
  assign n11268 = ~n554 & n11267;
  assign n11269 = ~n11266 & ~n11268;
  assign n11270 = ~n11265 & n11269;
  assign n11271 = ~n11264 & n11270;
  assign n11272 = ~pi5  & ~n11271;
  assign n11273 = pi5  & n11271;
  assign n11274 = ~n11272 & ~n11273;
  assign n11275 = n11260 & ~n11262;
  assign n11276 = ~n11263 & ~n11275;
  assign n11277 = ~n11274 & n11276;
  assign n11278 = ~n11263 & ~n11277;
  assign n11279 = ~n10712 & ~n10716;
  assign n11280 = ~n10717 & ~n11279;
  assign n11281 = ~n11278 & n11280;
  assign n11282 = n11274 & ~n11276;
  assign n11283 = ~n11277 & ~n11282;
  assign n11284 = pi1  & ~pi2 ;
  assign n11285 = ~pi1  & pi2 ;
  assign n11286 = ~n11284 & ~n11285;
  assign n11287 = ~pi0  & ~pi1 ;
  assign n11288 = ~n11286 & n11287;
  assign n11289 = pi0  & ~n11286;
  assign n11290 = ~n3638 & n11289;
  assign n11291 = ~n11288 & ~n11290;
  assign n11292 = ~n554 & ~n11291;
  assign n11293 = ~pi2  & n11292;
  assign n11294 = pi2  & ~n11292;
  assign n11295 = ~n11293 & ~n11294;
  assign n11296 = ~n795 & n9725;
  assign n11297 = ~n665 & n10702;
  assign n11298 = n4015 & n9719;
  assign n11299 = ~n720 & n11267;
  assign n11300 = ~n11298 & ~n11299;
  assign n11301 = ~n11297 & n11300;
  assign n11302 = ~n11296 & n11301;
  assign n11303 = pi5  & n11302;
  assign n11304 = ~pi5  & ~n11302;
  assign n11305 = ~n11303 & ~n11304;
  assign n11306 = ~n11295 & ~n11305;
  assign n11307 = ~n11255 & n11258;
  assign n11308 = n11255 & ~n11258;
  assign n11309 = ~n11307 & ~n11308;
  assign n11310 = n11295 & n11305;
  assign n11311 = ~n11309 & ~n11310;
  assign n11312 = ~n11306 & ~n11311;
  assign n11313 = n11283 & ~n11312;
  assign n11314 = ~n894 & n9725;
  assign n11315 = ~n795 & n10702;
  assign n11316 = n3959 & n9719;
  assign n11317 = ~n665 & n11267;
  assign n11318 = ~n11316 & ~n11317;
  assign n11319 = ~n11315 & n11318;
  assign n11320 = ~n11314 & n11319;
  assign n11321 = ~pi5  & ~n11320;
  assign n11322 = pi5  & n11320;
  assign n11323 = ~n11321 & ~n11322;
  assign n11324 = ~n11250 & n11253;
  assign n11325 = n11250 & ~n11253;
  assign n11326 = ~n11324 & ~n11325;
  assign n11327 = ~n11323 & ~n11326;
  assign n11328 = ~n1005 & n9725;
  assign n11329 = ~n894 & n10702;
  assign n11330 = n4122 & n9719;
  assign n11331 = ~n795 & n11267;
  assign n11332 = ~n11330 & ~n11331;
  assign n11333 = ~n11329 & n11332;
  assign n11334 = ~n11328 & n11333;
  assign n11335 = ~pi5  & ~n11334;
  assign n11336 = pi5  & n11334;
  assign n11337 = ~n11335 & ~n11336;
  assign n11338 = n11245 & n11248;
  assign n11339 = ~n11249 & ~n11338;
  assign n11340 = ~n11337 & n11339;
  assign n11341 = ~n11337 & ~n11339;
  assign n11342 = n11337 & n11339;
  assign n11343 = ~n11341 & ~n11342;
  assign n11344 = ~n1107 & n9725;
  assign n11345 = ~n1005 & n10702;
  assign n11346 = n4106 & n9719;
  assign n11347 = ~n894 & n11267;
  assign n11348 = ~n11346 & ~n11347;
  assign n11349 = ~n11345 & n11348;
  assign n11350 = ~n11344 & n11349;
  assign n11351 = ~pi5  & ~n11350;
  assign n11352 = pi5  & n11350;
  assign n11353 = ~n11351 & ~n11352;
  assign n11354 = n11240 & n11243;
  assign n11355 = ~n11244 & ~n11354;
  assign n11356 = ~n11353 & n11355;
  assign n11357 = ~n11353 & ~n11355;
  assign n11358 = n11353 & n11355;
  assign n11359 = ~n11357 & ~n11358;
  assign n11360 = ~n1230 & n9725;
  assign n11361 = ~n1107 & n10702;
  assign n11362 = n4307 & n9719;
  assign n11363 = ~n1005 & n11267;
  assign n11364 = ~n11362 & ~n11363;
  assign n11365 = ~n11361 & n11364;
  assign n11366 = ~n11360 & n11365;
  assign n11367 = ~pi5  & ~n11366;
  assign n11368 = pi5  & n11366;
  assign n11369 = ~n11367 & ~n11368;
  assign n11370 = ~n11235 & n11238;
  assign n11371 = n11235 & ~n11238;
  assign n11372 = ~n11370 & ~n11371;
  assign n11373 = ~n11369 & ~n11372;
  assign n11374 = ~n1338 & n9725;
  assign n11375 = ~n1230 & n10702;
  assign n11376 = n4323 & n9719;
  assign n11377 = ~n1107 & n11267;
  assign n11378 = ~n11376 & ~n11377;
  assign n11379 = ~n11375 & n11378;
  assign n11380 = ~n11374 & n11379;
  assign n11381 = ~pi5  & ~n11380;
  assign n11382 = pi5  & n11380;
  assign n11383 = ~n11381 & ~n11382;
  assign n11384 = ~n11230 & n11233;
  assign n11385 = n11230 & ~n11233;
  assign n11386 = ~n11384 & ~n11385;
  assign n11387 = ~n11383 & ~n11386;
  assign n11388 = ~n1426 & n9725;
  assign n11389 = ~n1338 & n10702;
  assign n11390 = n4753 & n9719;
  assign n11391 = ~n1230 & n11267;
  assign n11392 = ~n11390 & ~n11391;
  assign n11393 = ~n11389 & n11392;
  assign n11394 = ~n11388 & n11393;
  assign n11395 = ~pi5  & ~n11394;
  assign n11396 = pi5  & n11394;
  assign n11397 = ~n11395 & ~n11396;
  assign n11398 = n11225 & n11228;
  assign n11399 = ~n11229 & ~n11398;
  assign n11400 = ~n11397 & n11399;
  assign n11401 = ~n11397 & ~n11399;
  assign n11402 = n11397 & n11399;
  assign n11403 = ~n11401 & ~n11402;
  assign n11404 = n10832 & n11223;
  assign n11405 = ~n11224 & ~n11404;
  assign n11406 = ~n1531 & n9725;
  assign n11407 = ~n1426 & n10702;
  assign n11408 = n4533 & n9719;
  assign n11409 = ~n1338 & n11267;
  assign n11410 = ~n11408 & ~n11409;
  assign n11411 = ~n11407 & n11410;
  assign n11412 = ~n11406 & n11411;
  assign n11413 = pi5  & n11412;
  assign n11414 = ~pi5  & ~n11412;
  assign n11415 = ~n11413 & ~n11414;
  assign n11416 = n11405 & ~n11415;
  assign n11417 = n11219 & ~n11221;
  assign n11418 = ~n11222 & ~n11417;
  assign n11419 = ~n1610 & n9725;
  assign n11420 = ~n1531 & n10702;
  assign n11421 = n4724 & n9719;
  assign n11422 = ~n1426 & n11267;
  assign n11423 = ~n11421 & ~n11422;
  assign n11424 = ~n11420 & n11423;
  assign n11425 = ~n11419 & n11424;
  assign n11426 = pi5  & n11425;
  assign n11427 = ~pi5  & ~n11425;
  assign n11428 = ~n11426 & ~n11427;
  assign n11429 = n11418 & ~n11428;
  assign n11430 = ~n1740 & n9725;
  assign n11431 = ~n1610 & n10702;
  assign n11432 = n4708 & n9719;
  assign n11433 = ~n1531 & n11267;
  assign n11434 = ~n11432 & ~n11433;
  assign n11435 = ~n11431 & n11434;
  assign n11436 = ~n11430 & n11435;
  assign n11437 = ~pi5  & ~n11436;
  assign n11438 = pi5  & n11436;
  assign n11439 = ~n11437 & ~n11438;
  assign n11440 = n11215 & ~n11217;
  assign n11441 = ~n11218 & ~n11440;
  assign n11442 = ~n11439 & n11441;
  assign n11443 = ~n11439 & ~n11441;
  assign n11444 = n11439 & n11441;
  assign n11445 = ~n11443 & ~n11444;
  assign n11446 = ~n1811 & n9725;
  assign n11447 = ~n1740 & n10702;
  assign n11448 = n4951 & n9719;
  assign n11449 = ~n1610 & n11267;
  assign n11450 = ~n11448 & ~n11449;
  assign n11451 = ~n11447 & n11450;
  assign n11452 = ~n11446 & n11451;
  assign n11453 = ~pi5  & ~n11452;
  assign n11454 = pi5  & n11452;
  assign n11455 = ~n11453 & ~n11454;
  assign n11456 = n11210 & n11213;
  assign n11457 = ~n11214 & ~n11456;
  assign n11458 = ~n11455 & n11457;
  assign n11459 = ~n11455 & ~n11457;
  assign n11460 = n11455 & n11457;
  assign n11461 = ~n11459 & ~n11460;
  assign n11462 = ~n1900 & n9725;
  assign n11463 = ~n1811 & n10702;
  assign n11464 = n4967 & n9719;
  assign n11465 = ~n1740 & n11267;
  assign n11466 = ~n11464 & ~n11465;
  assign n11467 = ~n11463 & n11466;
  assign n11468 = ~n11462 & n11467;
  assign n11469 = ~pi5  & ~n11468;
  assign n11470 = pi5  & n11468;
  assign n11471 = ~n11469 & ~n11470;
  assign n11472 = ~n11205 & n11208;
  assign n11473 = n11205 & ~n11208;
  assign n11474 = ~n11472 & ~n11473;
  assign n11475 = ~n11471 & ~n11474;
  assign n11476 = n10901 & n11203;
  assign n11477 = ~n11204 & ~n11476;
  assign n11478 = ~n2006 & n9725;
  assign n11479 = ~n1900 & n10702;
  assign n11480 = n5344 & n9719;
  assign n11481 = ~n1811 & n11267;
  assign n11482 = ~n11480 & ~n11481;
  assign n11483 = ~n11479 & n11482;
  assign n11484 = ~n11478 & n11483;
  assign n11485 = pi5  & n11484;
  assign n11486 = ~pi5  & ~n11484;
  assign n11487 = ~n11485 & ~n11486;
  assign n11488 = n11477 & ~n11487;
  assign n11489 = n11199 & ~n11201;
  assign n11490 = ~n11202 & ~n11489;
  assign n11491 = ~n2058 & n9725;
  assign n11492 = ~n2006 & n10702;
  assign n11493 = n5180 & n9719;
  assign n11494 = ~n1900 & n11267;
  assign n11495 = ~n11493 & ~n11494;
  assign n11496 = ~n11492 & n11495;
  assign n11497 = ~n11491 & n11496;
  assign n11498 = pi5  & n11497;
  assign n11499 = ~pi5  & ~n11497;
  assign n11500 = ~n11498 & ~n11499;
  assign n11501 = n11490 & ~n11500;
  assign n11502 = n10931 & n11197;
  assign n11503 = ~n11198 & ~n11502;
  assign n11504 = ~n2178 & n9725;
  assign n11505 = ~n2058 & n10702;
  assign n11506 = n5554 & n9719;
  assign n11507 = ~n2006 & n11267;
  assign n11508 = ~n11506 & ~n11507;
  assign n11509 = ~n11505 & n11508;
  assign n11510 = ~n11504 & n11509;
  assign n11511 = pi5  & n11510;
  assign n11512 = ~pi5  & ~n11510;
  assign n11513 = ~n11511 & ~n11512;
  assign n11514 = n11503 & ~n11513;
  assign n11515 = ~n2278 & n9725;
  assign n11516 = ~n2178 & n10702;
  assign n11517 = n5538 & n9719;
  assign n11518 = ~n2058 & n11267;
  assign n11519 = ~n11517 & ~n11518;
  assign n11520 = ~n11516 & n11519;
  assign n11521 = ~n11515 & n11520;
  assign n11522 = ~pi5  & ~n11521;
  assign n11523 = pi5  & n11521;
  assign n11524 = ~n11522 & ~n11523;
  assign n11525 = n11193 & ~n11195;
  assign n11526 = ~n11196 & ~n11525;
  assign n11527 = ~n11524 & n11526;
  assign n11528 = ~n11524 & ~n11526;
  assign n11529 = n11524 & n11526;
  assign n11530 = ~n11528 & ~n11529;
  assign n11531 = ~n2369 & n9725;
  assign n11532 = ~n2278 & n10702;
  assign n11533 = n5779 & n9719;
  assign n11534 = ~n2178 & n11267;
  assign n11535 = ~n11533 & ~n11534;
  assign n11536 = ~n11532 & n11535;
  assign n11537 = ~n11531 & n11536;
  assign n11538 = ~pi5  & ~n11537;
  assign n11539 = pi5  & n11537;
  assign n11540 = ~n11538 & ~n11539;
  assign n11541 = ~n11188 & n11191;
  assign n11542 = n11188 & ~n11191;
  assign n11543 = ~n11541 & ~n11542;
  assign n11544 = ~n11540 & ~n11543;
  assign n11545 = ~n2457 & n9725;
  assign n11546 = ~n2369 & n10702;
  assign n11547 = n5795 & n9719;
  assign n11548 = ~n2278 & n11267;
  assign n11549 = ~n11547 & ~n11548;
  assign n11550 = ~n11546 & n11549;
  assign n11551 = ~n11545 & n11550;
  assign n11552 = ~pi5  & ~n11551;
  assign n11553 = pi5  & n11551;
  assign n11554 = ~n11552 & ~n11553;
  assign n11555 = n11183 & n11186;
  assign n11556 = ~n11187 & ~n11555;
  assign n11557 = ~n11554 & n11556;
  assign n11558 = ~n11554 & ~n11556;
  assign n11559 = n11554 & n11556;
  assign n11560 = ~n11558 & ~n11559;
  assign n11561 = n10986 & n11181;
  assign n11562 = ~n11182 & ~n11561;
  assign n11563 = ~n2554 & n9725;
  assign n11564 = ~n2457 & n10702;
  assign n11565 = n6218 & n9719;
  assign n11566 = ~n2369 & n11267;
  assign n11567 = ~n11565 & ~n11566;
  assign n11568 = ~n11564 & n11567;
  assign n11569 = ~n11563 & n11568;
  assign n11570 = pi5  & n11569;
  assign n11571 = ~pi5  & ~n11569;
  assign n11572 = ~n11570 & ~n11571;
  assign n11573 = n11562 & ~n11572;
  assign n11574 = n11002 & n11179;
  assign n11575 = ~n11180 & ~n11574;
  assign n11576 = ~n2640 & n9725;
  assign n11577 = ~n2554 & n10702;
  assign n11578 = n5979 & n9719;
  assign n11579 = ~n2457 & n11267;
  assign n11580 = ~n11578 & ~n11579;
  assign n11581 = ~n11577 & n11580;
  assign n11582 = ~n11576 & n11581;
  assign n11583 = pi5  & n11582;
  assign n11584 = ~pi5  & ~n11582;
  assign n11585 = ~n11583 & ~n11584;
  assign n11586 = n11575 & ~n11585;
  assign n11587 = n11175 & ~n11177;
  assign n11588 = ~n11178 & ~n11587;
  assign n11589 = ~n2676 & n9725;
  assign n11590 = ~n2640 & n10702;
  assign n11591 = n6445 & n9719;
  assign n11592 = ~n2554 & n11267;
  assign n11593 = ~n11591 & ~n11592;
  assign n11594 = ~n11590 & n11593;
  assign n11595 = ~n11589 & n11594;
  assign n11596 = pi5  & n11595;
  assign n11597 = ~pi5  & ~n11595;
  assign n11598 = ~n11596 & ~n11597;
  assign n11599 = n11588 & ~n11598;
  assign n11600 = ~n2748 & n9725;
  assign n11601 = ~n2676 & n10702;
  assign n11602 = n6597 & n9719;
  assign n11603 = ~n2640 & n11267;
  assign n11604 = ~n11602 & ~n11603;
  assign n11605 = ~n11601 & n11604;
  assign n11606 = ~n11600 & n11605;
  assign n11607 = ~pi5  & ~n11606;
  assign n11608 = pi5  & n11606;
  assign n11609 = ~n11607 & ~n11608;
  assign n11610 = n11171 & ~n11173;
  assign n11611 = ~n11174 & ~n11610;
  assign n11612 = ~n11609 & n11611;
  assign n11613 = ~n11609 & ~n11611;
  assign n11614 = n11609 & n11611;
  assign n11615 = ~n11613 & ~n11614;
  assign n11616 = ~n2803 & n9725;
  assign n11617 = ~n2748 & n10702;
  assign n11618 = n6427 & n9719;
  assign n11619 = ~n2676 & n11267;
  assign n11620 = ~n11618 & ~n11619;
  assign n11621 = ~n11617 & n11620;
  assign n11622 = ~n11616 & n11621;
  assign n11623 = ~pi5  & ~n11622;
  assign n11624 = pi5  & n11622;
  assign n11625 = ~n11623 & ~n11624;
  assign n11626 = n11166 & n11169;
  assign n11627 = ~n11170 & ~n11626;
  assign n11628 = ~n11625 & n11627;
  assign n11629 = ~n11625 & ~n11627;
  assign n11630 = n11625 & n11627;
  assign n11631 = ~n11629 & ~n11630;
  assign n11632 = ~n2891 & n9725;
  assign n11633 = ~n2803 & n10702;
  assign n11634 = n6715 & n9719;
  assign n11635 = ~n2748 & n11267;
  assign n11636 = ~n11634 & ~n11635;
  assign n11637 = ~n11633 & n11636;
  assign n11638 = ~n11632 & n11637;
  assign n11639 = ~pi5  & ~n11638;
  assign n11640 = pi5  & n11638;
  assign n11641 = ~n11639 & ~n11640;
  assign n11642 = ~n11161 & n11164;
  assign n11643 = n11161 & ~n11164;
  assign n11644 = ~n11642 & ~n11643;
  assign n11645 = ~n11641 & ~n11644;
  assign n11646 = n11071 & n11159;
  assign n11647 = ~n11160 & ~n11646;
  assign n11648 = ~n2927 & n9725;
  assign n11649 = ~n2891 & n10702;
  assign n11650 = n7014 & n9719;
  assign n11651 = ~n2803 & n11267;
  assign n11652 = ~n11650 & ~n11651;
  assign n11653 = ~n11649 & n11652;
  assign n11654 = ~n11648 & n11653;
  assign n11655 = pi5  & n11654;
  assign n11656 = ~pi5  & ~n11654;
  assign n11657 = ~n11655 & ~n11656;
  assign n11658 = n11647 & ~n11657;
  assign n11659 = n11155 & ~n11157;
  assign n11660 = ~n11158 & ~n11659;
  assign n11661 = ~n3005 & n9725;
  assign n11662 = ~n2927 & n10702;
  assign n11663 = n7026 & n9719;
  assign n11664 = ~n2891 & n11267;
  assign n11665 = ~n11663 & ~n11664;
  assign n11666 = ~n11662 & n11665;
  assign n11667 = ~n11661 & n11666;
  assign n11668 = pi5  & n11667;
  assign n11669 = ~pi5  & ~n11667;
  assign n11670 = ~n11668 & ~n11669;
  assign n11671 = n11660 & ~n11670;
  assign n11672 = n11102 & n11153;
  assign n11673 = ~n11154 & ~n11672;
  assign n11674 = ~n3097 & n9725;
  assign n11675 = ~n3005 & n10702;
  assign n11676 = n6694 & n9719;
  assign n11677 = ~n2927 & n11267;
  assign n11678 = ~n11676 & ~n11677;
  assign n11679 = ~n11675 & n11678;
  assign n11680 = ~n11674 & n11679;
  assign n11681 = pi5  & n11680;
  assign n11682 = ~pi5  & ~n11680;
  assign n11683 = ~n11681 & ~n11682;
  assign n11684 = n11673 & ~n11683;
  assign n11685 = ~n3166 & n9725;
  assign n11686 = ~n3097 & n10702;
  assign n11687 = n7071 & n9719;
  assign n11688 = ~n3005 & n11267;
  assign n11689 = ~n11687 & ~n11688;
  assign n11690 = ~n11686 & n11689;
  assign n11691 = ~n11685 & n11690;
  assign n11692 = ~pi5  & ~n11691;
  assign n11693 = pi5  & n11691;
  assign n11694 = ~n11692 & ~n11693;
  assign n11695 = n11149 & ~n11151;
  assign n11696 = ~n11152 & ~n11695;
  assign n11697 = ~n11694 & n11696;
  assign n11698 = ~n11694 & ~n11696;
  assign n11699 = n11694 & n11696;
  assign n11700 = ~n11698 & ~n11699;
  assign n11701 = ~n3226 & n9725;
  assign n11702 = ~n3166 & n10702;
  assign n11703 = n7121 & n9719;
  assign n11704 = ~n3097 & n11267;
  assign n11705 = ~n11703 & ~n11704;
  assign n11706 = ~n11702 & n11705;
  assign n11707 = ~n11701 & n11706;
  assign n11708 = pi5  & n11707;
  assign n11709 = ~pi5  & ~n11707;
  assign n11710 = ~n11708 & ~n11709;
  assign n11711 = n11137 & n11147;
  assign n11712 = ~n11148 & ~n11711;
  assign n11713 = ~n11710 & n11712;
  assign n11714 = ~n3263 & n9725;
  assign n11715 = ~n3226 & n10702;
  assign n11716 = n7175 & n9719;
  assign n11717 = ~n3166 & n11267;
  assign n11718 = ~n11716 & ~n11717;
  assign n11719 = ~n11715 & n11718;
  assign n11720 = ~n11714 & n11719;
  assign n11721 = ~pi5  & ~n11720;
  assign n11722 = pi5  & n11720;
  assign n11723 = ~n11721 & ~n11722;
  assign n11724 = pi8  & ~n11125;
  assign n11725 = n11132 & ~n11724;
  assign n11726 = ~n11132 & n11724;
  assign n11727 = ~n11725 & ~n11726;
  assign n11728 = ~n11723 & n11727;
  assign n11729 = ~n11723 & ~n11727;
  assign n11730 = n11723 & n11727;
  assign n11731 = ~n11729 & ~n11730;
  assign n11732 = ~n3360 & n9725;
  assign n11733 = ~n3263 & n10702;
  assign n11734 = n7221 & n9719;
  assign n11735 = ~n3226 & n11267;
  assign n11736 = ~n11734 & ~n11735;
  assign n11737 = ~n11733 & n11736;
  assign n11738 = ~n11732 & n11737;
  assign n11739 = pi5  & n11738;
  assign n11740 = ~pi5  & ~n11738;
  assign n11741 = ~n11739 & ~n11740;
  assign n11742 = pi8  & n11123;
  assign n11743 = ~n11122 & n11742;
  assign n11744 = n11122 & ~n11742;
  assign n11745 = ~n11743 & ~n11744;
  assign n11746 = ~n11741 & n11745;
  assign n11747 = ~n7942 & n9719;
  assign n11748 = ~n3506 & n11267;
  assign n11749 = ~n3450 & n10702;
  assign n11750 = ~n11748 & ~n11749;
  assign n11751 = ~n11747 & n11750;
  assign n11752 = ~n3450 & ~n9715;
  assign n11753 = pi5  & ~n11752;
  assign n11754 = n11751 & n11753;
  assign n11755 = ~n3450 & n9725;
  assign n11756 = ~n3506 & n10702;
  assign n11757 = n7265 & n9719;
  assign n11758 = ~n3360 & n11267;
  assign n11759 = ~n11757 & ~n11758;
  assign n11760 = ~n11756 & n11759;
  assign n11761 = ~n11755 & n11760;
  assign n11762 = n11754 & n11761;
  assign n11763 = n11123 & n11762;
  assign n11764 = ~n11123 & n11762;
  assign n11765 = n11123 & ~n11762;
  assign n11766 = ~n11764 & ~n11765;
  assign n11767 = ~n3506 & n9725;
  assign n11768 = ~n3360 & n10702;
  assign n11769 = n7323 & n9719;
  assign n11770 = ~n3263 & n11267;
  assign n11771 = ~n11769 & ~n11770;
  assign n11772 = ~n11768 & n11771;
  assign n11773 = ~n11767 & n11772;
  assign n11774 = pi5  & n11773;
  assign n11775 = ~pi5  & ~n11773;
  assign n11776 = ~n11774 & ~n11775;
  assign n11777 = ~n11766 & ~n11776;
  assign n11778 = ~n11763 & ~n11777;
  assign n11779 = n11741 & ~n11745;
  assign n11780 = ~n11746 & ~n11779;
  assign n11781 = ~n11778 & n11780;
  assign n11782 = ~n11746 & ~n11781;
  assign n11783 = ~n11731 & ~n11782;
  assign n11784 = ~n11728 & ~n11783;
  assign n11785 = n11710 & ~n11712;
  assign n11786 = ~n11713 & ~n11785;
  assign n11787 = ~n11784 & n11786;
  assign n11788 = ~n11713 & ~n11787;
  assign n11789 = ~n11700 & ~n11788;
  assign n11790 = ~n11697 & ~n11789;
  assign n11791 = n11673 & n11683;
  assign n11792 = ~n11673 & ~n11683;
  assign n11793 = ~n11791 & ~n11792;
  assign n11794 = ~n11790 & ~n11793;
  assign n11795 = ~n11684 & ~n11794;
  assign n11796 = n11660 & n11670;
  assign n11797 = ~n11660 & ~n11670;
  assign n11798 = ~n11796 & ~n11797;
  assign n11799 = ~n11795 & ~n11798;
  assign n11800 = ~n11671 & ~n11799;
  assign n11801 = ~n11647 & n11657;
  assign n11802 = ~n11658 & ~n11801;
  assign n11803 = ~n11800 & n11802;
  assign n11804 = ~n11658 & ~n11803;
  assign n11805 = n11641 & n11644;
  assign n11806 = ~n11645 & ~n11805;
  assign n11807 = ~n11804 & n11806;
  assign n11808 = ~n11645 & ~n11807;
  assign n11809 = ~n11631 & ~n11808;
  assign n11810 = ~n11628 & ~n11809;
  assign n11811 = ~n11615 & ~n11810;
  assign n11812 = ~n11612 & ~n11811;
  assign n11813 = n11588 & n11598;
  assign n11814 = ~n11588 & ~n11598;
  assign n11815 = ~n11813 & ~n11814;
  assign n11816 = ~n11812 & ~n11815;
  assign n11817 = ~n11599 & ~n11816;
  assign n11818 = n11575 & n11585;
  assign n11819 = ~n11575 & ~n11585;
  assign n11820 = ~n11818 & ~n11819;
  assign n11821 = ~n11817 & ~n11820;
  assign n11822 = ~n11586 & ~n11821;
  assign n11823 = ~n11562 & n11572;
  assign n11824 = ~n11573 & ~n11823;
  assign n11825 = ~n11822 & n11824;
  assign n11826 = ~n11573 & ~n11825;
  assign n11827 = ~n11560 & ~n11826;
  assign n11828 = ~n11557 & ~n11827;
  assign n11829 = n11540 & n11543;
  assign n11830 = ~n11544 & ~n11829;
  assign n11831 = ~n11828 & n11830;
  assign n11832 = ~n11544 & ~n11831;
  assign n11833 = ~n11530 & ~n11832;
  assign n11834 = ~n11527 & ~n11833;
  assign n11835 = n11503 & n11513;
  assign n11836 = ~n11503 & ~n11513;
  assign n11837 = ~n11835 & ~n11836;
  assign n11838 = ~n11834 & ~n11837;
  assign n11839 = ~n11514 & ~n11838;
  assign n11840 = n11490 & n11500;
  assign n11841 = ~n11490 & ~n11500;
  assign n11842 = ~n11840 & ~n11841;
  assign n11843 = ~n11839 & ~n11842;
  assign n11844 = ~n11501 & ~n11843;
  assign n11845 = ~n11477 & n11487;
  assign n11846 = ~n11488 & ~n11845;
  assign n11847 = ~n11844 & n11846;
  assign n11848 = ~n11488 & ~n11847;
  assign n11849 = n11471 & n11474;
  assign n11850 = ~n11475 & ~n11849;
  assign n11851 = ~n11848 & n11850;
  assign n11852 = ~n11475 & ~n11851;
  assign n11853 = ~n11461 & ~n11852;
  assign n11854 = ~n11458 & ~n11853;
  assign n11855 = ~n11445 & ~n11854;
  assign n11856 = ~n11442 & ~n11855;
  assign n11857 = n11418 & n11428;
  assign n11858 = ~n11418 & ~n11428;
  assign n11859 = ~n11857 & ~n11858;
  assign n11860 = ~n11856 & ~n11859;
  assign n11861 = ~n11429 & ~n11860;
  assign n11862 = ~n11405 & n11415;
  assign n11863 = ~n11416 & ~n11862;
  assign n11864 = ~n11861 & n11863;
  assign n11865 = ~n11416 & ~n11864;
  assign n11866 = ~n11403 & ~n11865;
  assign n11867 = ~n11400 & ~n11866;
  assign n11868 = n11383 & n11386;
  assign n11869 = ~n11387 & ~n11868;
  assign n11870 = ~n11867 & n11869;
  assign n11871 = ~n11387 & ~n11870;
  assign n11872 = n11369 & n11372;
  assign n11873 = ~n11373 & ~n11872;
  assign n11874 = ~n11871 & n11873;
  assign n11875 = ~n11373 & ~n11874;
  assign n11876 = ~n11359 & ~n11875;
  assign n11877 = ~n11356 & ~n11876;
  assign n11878 = ~n11343 & ~n11877;
  assign n11879 = ~n11340 & ~n11878;
  assign n11880 = n11323 & n11326;
  assign n11881 = ~n11327 & ~n11880;
  assign n11882 = ~n11879 & n11881;
  assign n11883 = ~n11327 & ~n11882;
  assign n11884 = ~n11306 & ~n11310;
  assign n11885 = n11309 & ~n11884;
  assign n11886 = ~n11309 & n11884;
  assign n11887 = ~n11885 & ~n11886;
  assign n11888 = ~n11883 & n11887;
  assign n11889 = n11883 & ~n11887;
  assign n11890 = ~n11888 & ~n11889;
  assign n11891 = n11879 & ~n11881;
  assign n11892 = ~n11882 & ~n11891;
  assign n11893 = ~n3744 & n11289;
  assign n11894 = ~pi0  & pi1 ;
  assign n11895 = ~n554 & n11894;
  assign n11896 = ~n720 & n11288;
  assign n11897 = ~n11895 & ~n11896;
  assign n11898 = ~n11893 & n11897;
  assign n11899 = pi2  & n11898;
  assign n11900 = ~pi2  & ~n11898;
  assign n11901 = ~n11899 & ~n11900;
  assign n11902 = n11892 & ~n11901;
  assign n11903 = n11343 & n11877;
  assign n11904 = ~n11878 & ~n11903;
  assign n11905 = ~n665 & n11288;
  assign n11906 = ~n720 & n11894;
  assign n11907 = n3979 & n11289;
  assign n11908 = pi0  & n11286;
  assign n11909 = ~n554 & n11908;
  assign n11910 = ~n11907 & ~n11909;
  assign n11911 = ~n11906 & n11910;
  assign n11912 = ~n11905 & n11911;
  assign n11913 = pi2  & n11912;
  assign n11914 = ~pi2  & ~n11912;
  assign n11915 = ~n11913 & ~n11914;
  assign n11916 = n11904 & ~n11915;
  assign n11917 = n11359 & n11875;
  assign n11918 = ~n11876 & ~n11917;
  assign n11919 = ~n795 & n11288;
  assign n11920 = ~n665 & n11894;
  assign n11921 = n4015 & n11289;
  assign n11922 = ~n720 & n11908;
  assign n11923 = ~n11921 & ~n11922;
  assign n11924 = ~n11920 & n11923;
  assign n11925 = ~n11919 & n11924;
  assign n11926 = pi2  & n11925;
  assign n11927 = ~pi2  & ~n11925;
  assign n11928 = ~n11926 & ~n11927;
  assign n11929 = n11918 & ~n11928;
  assign n11930 = n11871 & ~n11873;
  assign n11931 = ~n11874 & ~n11930;
  assign n11932 = ~n894 & n11288;
  assign n11933 = ~n795 & n11894;
  assign n11934 = n3959 & n11289;
  assign n11935 = ~n665 & n11908;
  assign n11936 = ~n11934 & ~n11935;
  assign n11937 = ~n11933 & n11936;
  assign n11938 = ~n11932 & n11937;
  assign n11939 = pi2  & n11938;
  assign n11940 = ~pi2  & ~n11938;
  assign n11941 = ~n11939 & ~n11940;
  assign n11942 = n11931 & ~n11941;
  assign n11943 = n11867 & ~n11869;
  assign n11944 = ~n11870 & ~n11943;
  assign n11945 = ~n1005 & n11288;
  assign n11946 = ~n894 & n11894;
  assign n11947 = n4122 & n11289;
  assign n11948 = ~n795 & n11908;
  assign n11949 = ~n11947 & ~n11948;
  assign n11950 = ~n11946 & n11949;
  assign n11951 = ~n11945 & n11950;
  assign n11952 = pi2  & n11951;
  assign n11953 = ~pi2  & ~n11951;
  assign n11954 = ~n11952 & ~n11953;
  assign n11955 = n11944 & ~n11954;
  assign n11956 = n11944 & n11954;
  assign n11957 = ~n11944 & ~n11954;
  assign n11958 = ~n11956 & ~n11957;
  assign n11959 = ~n1107 & n11288;
  assign n11960 = ~n1005 & n11894;
  assign n11961 = n4106 & n11289;
  assign n11962 = ~n894 & n11908;
  assign n11963 = ~n11961 & ~n11962;
  assign n11964 = ~n11960 & n11963;
  assign n11965 = ~n11959 & n11964;
  assign n11966 = pi2  & n11965;
  assign n11967 = ~pi2  & ~n11965;
  assign n11968 = ~n11966 & ~n11967;
  assign n11969 = n11861 & ~n11863;
  assign n11970 = ~n11864 & ~n11969;
  assign n11971 = n11856 & n11859;
  assign n11972 = ~n11860 & ~n11971;
  assign n11973 = ~n1426 & n11288;
  assign n11974 = ~n1338 & n11894;
  assign n11975 = n4753 & n11289;
  assign n11976 = ~n1230 & n11908;
  assign n11977 = ~n11975 & ~n11976;
  assign n11978 = ~n11974 & n11977;
  assign n11979 = ~n11973 & n11978;
  assign n11980 = pi2  & n11979;
  assign n11981 = ~pi2  & ~n11979;
  assign n11982 = ~n11980 & ~n11981;
  assign n11983 = ~n1531 & n11288;
  assign n11984 = ~n1426 & n11894;
  assign n11985 = n4533 & n11289;
  assign n11986 = ~n1338 & n11908;
  assign n11987 = ~n11985 & ~n11986;
  assign n11988 = ~n11984 & n11987;
  assign n11989 = ~n11983 & n11988;
  assign n11990 = pi2  & n11989;
  assign n11991 = ~pi2  & ~n11989;
  assign n11992 = ~n11990 & ~n11991;
  assign n11993 = ~n1610 & n11288;
  assign n11994 = ~n1531 & n11894;
  assign n11995 = n4724 & n11289;
  assign n11996 = ~n1426 & n11908;
  assign n11997 = ~n11995 & ~n11996;
  assign n11998 = ~n11994 & n11997;
  assign n11999 = ~n11993 & n11998;
  assign n12000 = pi2  & n11999;
  assign n12001 = ~pi2  & ~n11999;
  assign n12002 = ~n12000 & ~n12001;
  assign n12003 = n11844 & ~n11846;
  assign n12004 = ~n11847 & ~n12003;
  assign n12005 = n11839 & n11842;
  assign n12006 = ~n11843 & ~n12005;
  assign n12007 = n11834 & n11837;
  assign n12008 = ~n11838 & ~n12007;
  assign n12009 = ~n2006 & n11288;
  assign n12010 = ~n1900 & n11894;
  assign n12011 = n5344 & n11289;
  assign n12012 = ~n1811 & n11908;
  assign n12013 = ~n12011 & ~n12012;
  assign n12014 = ~n12010 & n12013;
  assign n12015 = ~n12009 & n12014;
  assign n12016 = pi2  & n12015;
  assign n12017 = ~pi2  & ~n12015;
  assign n12018 = ~n12016 & ~n12017;
  assign n12019 = ~n2058 & n11288;
  assign n12020 = ~n2006 & n11894;
  assign n12021 = n5180 & n11289;
  assign n12022 = ~n1900 & n11908;
  assign n12023 = ~n12021 & ~n12022;
  assign n12024 = ~n12020 & n12023;
  assign n12025 = ~n12019 & n12024;
  assign n12026 = pi2  & n12025;
  assign n12027 = ~pi2  & ~n12025;
  assign n12028 = ~n12026 & ~n12027;
  assign n12029 = ~n2178 & n11288;
  assign n12030 = ~n2058 & n11894;
  assign n12031 = n5554 & n11289;
  assign n12032 = ~n2006 & n11908;
  assign n12033 = ~n12031 & ~n12032;
  assign n12034 = ~n12030 & n12033;
  assign n12035 = ~n12029 & n12034;
  assign n12036 = pi2  & n12035;
  assign n12037 = ~pi2  & ~n12035;
  assign n12038 = ~n12036 & ~n12037;
  assign n12039 = n11822 & ~n11824;
  assign n12040 = ~n11825 & ~n12039;
  assign n12041 = n11817 & n11820;
  assign n12042 = ~n11821 & ~n12041;
  assign n12043 = n11812 & n11815;
  assign n12044 = ~n11816 & ~n12043;
  assign n12045 = ~n2554 & n11288;
  assign n12046 = ~n2457 & n11894;
  assign n12047 = n6218 & n11289;
  assign n12048 = ~n2369 & n11908;
  assign n12049 = ~n12047 & ~n12048;
  assign n12050 = ~n12046 & n12049;
  assign n12051 = ~n12045 & n12050;
  assign n12052 = pi2  & n12051;
  assign n12053 = ~pi2  & ~n12051;
  assign n12054 = ~n12052 & ~n12053;
  assign n12055 = ~n2640 & n11288;
  assign n12056 = ~n2554 & n11894;
  assign n12057 = n5979 & n11289;
  assign n12058 = ~n2457 & n11908;
  assign n12059 = ~n12057 & ~n12058;
  assign n12060 = ~n12056 & n12059;
  assign n12061 = ~n12055 & n12060;
  assign n12062 = pi2  & n12061;
  assign n12063 = ~pi2  & ~n12061;
  assign n12064 = ~n12062 & ~n12063;
  assign n12065 = ~n2676 & n11288;
  assign n12066 = ~n2640 & n11894;
  assign n12067 = n6445 & n11289;
  assign n12068 = ~n2554 & n11908;
  assign n12069 = ~n12067 & ~n12068;
  assign n12070 = ~n12066 & n12069;
  assign n12071 = ~n12065 & n12070;
  assign n12072 = pi2  & n12071;
  assign n12073 = ~pi2  & ~n12071;
  assign n12074 = ~n12072 & ~n12073;
  assign n12075 = n11800 & ~n11802;
  assign n12076 = ~n11803 & ~n12075;
  assign n12077 = n11795 & n11798;
  assign n12078 = ~n11799 & ~n12077;
  assign n12079 = n11790 & n11793;
  assign n12080 = ~n11794 & ~n12079;
  assign n12081 = ~n2927 & n11288;
  assign n12082 = ~n2891 & n11894;
  assign n12083 = n7014 & n11289;
  assign n12084 = ~n2803 & n11908;
  assign n12085 = ~n12083 & ~n12084;
  assign n12086 = ~n12082 & n12085;
  assign n12087 = ~n12081 & n12086;
  assign n12088 = pi2  & n12087;
  assign n12089 = ~pi2  & ~n12087;
  assign n12090 = ~n12088 & ~n12089;
  assign n12091 = ~n3005 & n11288;
  assign n12092 = ~n2927 & n11894;
  assign n12093 = n7026 & n11289;
  assign n12094 = ~n2891 & n11908;
  assign n12095 = ~n12093 & ~n12094;
  assign n12096 = ~n12092 & n12095;
  assign n12097 = ~n12091 & n12096;
  assign n12098 = pi2  & n12097;
  assign n12099 = ~pi2  & ~n12097;
  assign n12100 = ~n12098 & ~n12099;
  assign n12101 = ~n3097 & n11288;
  assign n12102 = ~n3005 & n11894;
  assign n12103 = n6694 & n11289;
  assign n12104 = ~n2927 & n11908;
  assign n12105 = ~n12103 & ~n12104;
  assign n12106 = ~n12102 & n12105;
  assign n12107 = ~n12101 & n12106;
  assign n12108 = pi2  & n12107;
  assign n12109 = ~pi2  & ~n12107;
  assign n12110 = ~n12108 & ~n12109;
  assign n12111 = n11778 & ~n11780;
  assign n12112 = ~n11781 & ~n12111;
  assign n12113 = ~n3226 & n11288;
  assign n12114 = ~n3166 & n11894;
  assign n12115 = n7121 & n11289;
  assign n12116 = ~n3097 & n11908;
  assign n12117 = ~n12115 & ~n12116;
  assign n12118 = ~n12114 & n12117;
  assign n12119 = ~n12113 & n12118;
  assign n12120 = pi2  & n12119;
  assign n12121 = ~pi2  & ~n12119;
  assign n12122 = ~n12120 & ~n12121;
  assign n12123 = pi5  & ~n11754;
  assign n12124 = n11761 & ~n12123;
  assign n12125 = ~n11761 & n12123;
  assign n12126 = ~n12124 & ~n12125;
  assign n12127 = ~n3360 & n11288;
  assign n12128 = ~n3263 & n11894;
  assign n12129 = n7221 & n11289;
  assign n12130 = ~n3226 & n11908;
  assign n12131 = ~n12129 & ~n12130;
  assign n12132 = ~n12128 & n12131;
  assign n12133 = ~n12127 & n12132;
  assign n12134 = pi2  & n12133;
  assign n12135 = ~pi2  & ~n12133;
  assign n12136 = ~n12134 & ~n12135;
  assign n12137 = ~n3450 & ~n11287;
  assign n12138 = ~n3506 & n11908;
  assign n12139 = pi2  & n11289;
  assign n12140 = n7265 & n12139;
  assign n12141 = ~n3450 & n11288;
  assign n12142 = ~n3506 & n11894;
  assign n12143 = ~n3360 & n11908;
  assign n12144 = ~n12142 & ~n12143;
  assign n12145 = ~n12141 & n12144;
  assign n12146 = pi2  & ~n12145;
  assign n12147 = ~n7942 & n12139;
  assign n12148 = pi2  & ~n12147;
  assign n12149 = ~n12146 & n12148;
  assign n12150 = ~n12140 & n12149;
  assign n12151 = ~n12138 & n12150;
  assign n12152 = ~n12137 & n12151;
  assign n12153 = n11752 & n12152;
  assign n12154 = ~n11752 & ~n12152;
  assign n12155 = ~n3506 & n11288;
  assign n12156 = ~n3360 & n11894;
  assign n12157 = n7323 & n11289;
  assign n12158 = ~n3263 & n11908;
  assign n12159 = ~n12157 & ~n12158;
  assign n12160 = ~n12156 & n12159;
  assign n12161 = ~n12155 & n12160;
  assign n12162 = pi2  & ~n12161;
  assign n12163 = ~pi2  & n12161;
  assign n12164 = ~n12162 & ~n12163;
  assign n12165 = ~n12154 & n12164;
  assign n12166 = ~n12153 & ~n12165;
  assign n12167 = ~n12136 & ~n12166;
  assign n12168 = n12136 & n12166;
  assign n12169 = pi5  & n11752;
  assign n12170 = ~n11751 & n12169;
  assign n12171 = n11751 & ~n12169;
  assign n12172 = ~n12170 & ~n12171;
  assign n12173 = ~n12168 & n12172;
  assign n12174 = ~n12167 & ~n12173;
  assign n12175 = n12126 & ~n12174;
  assign n12176 = ~n12126 & n12174;
  assign n12177 = ~n3263 & n11288;
  assign n12178 = ~n3226 & n11894;
  assign n12179 = n7175 & n11289;
  assign n12180 = ~n3166 & n11908;
  assign n12181 = ~n12179 & ~n12180;
  assign n12182 = ~n12178 & n12181;
  assign n12183 = ~n12177 & n12182;
  assign n12184 = pi2  & ~n12183;
  assign n12185 = ~pi2  & n12183;
  assign n12186 = ~n12184 & ~n12185;
  assign n12187 = ~n12176 & n12186;
  assign n12188 = ~n12175 & ~n12187;
  assign n12189 = ~n12122 & ~n12188;
  assign n12190 = n12122 & n12188;
  assign n12191 = n11766 & n11776;
  assign n12192 = ~n11777 & ~n12191;
  assign n12193 = ~n12190 & n12192;
  assign n12194 = ~n12189 & ~n12193;
  assign n12195 = n12112 & ~n12194;
  assign n12196 = ~n12112 & n12194;
  assign n12197 = ~n3166 & n11288;
  assign n12198 = ~n3097 & n11894;
  assign n12199 = n7071 & n11289;
  assign n12200 = ~n3005 & n11908;
  assign n12201 = ~n12199 & ~n12200;
  assign n12202 = ~n12198 & n12201;
  assign n12203 = ~n12197 & n12202;
  assign n12204 = pi2  & ~n12203;
  assign n12205 = ~pi2  & n12203;
  assign n12206 = ~n12204 & ~n12205;
  assign n12207 = ~n12196 & n12206;
  assign n12208 = ~n12195 & ~n12207;
  assign n12209 = ~n12110 & ~n12208;
  assign n12210 = n12110 & n12208;
  assign n12211 = n11731 & n11782;
  assign n12212 = ~n11783 & ~n12211;
  assign n12213 = ~n12210 & n12212;
  assign n12214 = ~n12209 & ~n12213;
  assign n12215 = ~n12100 & ~n12214;
  assign n12216 = n12100 & n12214;
  assign n12217 = n11784 & ~n11786;
  assign n12218 = ~n11787 & ~n12217;
  assign n12219 = ~n12216 & n12218;
  assign n12220 = ~n12215 & ~n12219;
  assign n12221 = ~n12090 & ~n12220;
  assign n12222 = n12090 & n12220;
  assign n12223 = n11700 & n11788;
  assign n12224 = ~n11789 & ~n12223;
  assign n12225 = ~n12222 & n12224;
  assign n12226 = ~n12221 & ~n12225;
  assign n12227 = n12080 & ~n12226;
  assign n12228 = ~n12080 & n12226;
  assign n12229 = ~n2891 & n11288;
  assign n12230 = ~n2803 & n11894;
  assign n12231 = n6715 & n11289;
  assign n12232 = ~n2748 & n11908;
  assign n12233 = ~n12231 & ~n12232;
  assign n12234 = ~n12230 & n12233;
  assign n12235 = ~n12229 & n12234;
  assign n12236 = pi2  & ~n12235;
  assign n12237 = ~pi2  & n12235;
  assign n12238 = ~n12236 & ~n12237;
  assign n12239 = ~n12228 & n12238;
  assign n12240 = ~n12227 & ~n12239;
  assign n12241 = n12078 & ~n12240;
  assign n12242 = ~n12078 & n12240;
  assign n12243 = ~n2803 & n11288;
  assign n12244 = ~n2748 & n11894;
  assign n12245 = n6427 & n11289;
  assign n12246 = ~n2676 & n11908;
  assign n12247 = ~n12245 & ~n12246;
  assign n12248 = ~n12244 & n12247;
  assign n12249 = ~n12243 & n12248;
  assign n12250 = pi2  & ~n12249;
  assign n12251 = ~pi2  & n12249;
  assign n12252 = ~n12250 & ~n12251;
  assign n12253 = ~n12242 & n12252;
  assign n12254 = ~n12241 & ~n12253;
  assign n12255 = n12076 & ~n12254;
  assign n12256 = ~n12076 & n12254;
  assign n12257 = ~n2748 & n11288;
  assign n12258 = ~n2676 & n11894;
  assign n12259 = n6597 & n11289;
  assign n12260 = ~n2640 & n11908;
  assign n12261 = ~n12259 & ~n12260;
  assign n12262 = ~n12258 & n12261;
  assign n12263 = ~n12257 & n12262;
  assign n12264 = pi2  & ~n12263;
  assign n12265 = ~pi2  & n12263;
  assign n12266 = ~n12264 & ~n12265;
  assign n12267 = ~n12256 & n12266;
  assign n12268 = ~n12255 & ~n12267;
  assign n12269 = ~n12074 & ~n12268;
  assign n12270 = n12074 & n12268;
  assign n12271 = n11804 & ~n11806;
  assign n12272 = ~n11807 & ~n12271;
  assign n12273 = ~n12270 & n12272;
  assign n12274 = ~n12269 & ~n12273;
  assign n12275 = ~n12064 & ~n12274;
  assign n12276 = n12064 & n12274;
  assign n12277 = n11631 & n11808;
  assign n12278 = ~n11809 & ~n12277;
  assign n12279 = ~n12276 & n12278;
  assign n12280 = ~n12275 & ~n12279;
  assign n12281 = ~n12054 & ~n12280;
  assign n12282 = n12054 & n12280;
  assign n12283 = n11615 & n11810;
  assign n12284 = ~n11811 & ~n12283;
  assign n12285 = ~n12282 & n12284;
  assign n12286 = ~n12281 & ~n12285;
  assign n12287 = n12044 & ~n12286;
  assign n12288 = ~n12044 & n12286;
  assign n12289 = ~n2457 & n11288;
  assign n12290 = ~n2369 & n11894;
  assign n12291 = n5795 & n11289;
  assign n12292 = ~n2278 & n11908;
  assign n12293 = ~n12291 & ~n12292;
  assign n12294 = ~n12290 & n12293;
  assign n12295 = ~n12289 & n12294;
  assign n12296 = pi2  & ~n12295;
  assign n12297 = ~pi2  & n12295;
  assign n12298 = ~n12296 & ~n12297;
  assign n12299 = ~n12288 & n12298;
  assign n12300 = ~n12287 & ~n12299;
  assign n12301 = n12042 & ~n12300;
  assign n12302 = ~n12042 & n12300;
  assign n12303 = ~n2369 & n11288;
  assign n12304 = ~n2278 & n11894;
  assign n12305 = n5779 & n11289;
  assign n12306 = ~n2178 & n11908;
  assign n12307 = ~n12305 & ~n12306;
  assign n12308 = ~n12304 & n12307;
  assign n12309 = ~n12303 & n12308;
  assign n12310 = pi2  & ~n12309;
  assign n12311 = ~pi2  & n12309;
  assign n12312 = ~n12310 & ~n12311;
  assign n12313 = ~n12302 & n12312;
  assign n12314 = ~n12301 & ~n12313;
  assign n12315 = n12040 & ~n12314;
  assign n12316 = ~n12040 & n12314;
  assign n12317 = ~n2278 & n11288;
  assign n12318 = ~n2178 & n11894;
  assign n12319 = n5538 & n11289;
  assign n12320 = ~n2058 & n11908;
  assign n12321 = ~n12319 & ~n12320;
  assign n12322 = ~n12318 & n12321;
  assign n12323 = ~n12317 & n12322;
  assign n12324 = pi2  & ~n12323;
  assign n12325 = ~pi2  & n12323;
  assign n12326 = ~n12324 & ~n12325;
  assign n12327 = ~n12316 & n12326;
  assign n12328 = ~n12315 & ~n12327;
  assign n12329 = ~n12038 & ~n12328;
  assign n12330 = n12038 & n12328;
  assign n12331 = n11560 & n11826;
  assign n12332 = ~n11827 & ~n12331;
  assign n12333 = ~n12330 & n12332;
  assign n12334 = ~n12329 & ~n12333;
  assign n12335 = ~n12028 & ~n12334;
  assign n12336 = n12028 & n12334;
  assign n12337 = n11828 & ~n11830;
  assign n12338 = ~n11831 & ~n12337;
  assign n12339 = ~n12336 & n12338;
  assign n12340 = ~n12335 & ~n12339;
  assign n12341 = ~n12018 & ~n12340;
  assign n12342 = n12018 & n12340;
  assign n12343 = n11530 & n11832;
  assign n12344 = ~n11833 & ~n12343;
  assign n12345 = ~n12342 & n12344;
  assign n12346 = ~n12341 & ~n12345;
  assign n12347 = n12008 & ~n12346;
  assign n12348 = ~n12008 & n12346;
  assign n12349 = ~n1900 & n11288;
  assign n12350 = ~n1811 & n11894;
  assign n12351 = n4967 & n11289;
  assign n12352 = ~n1740 & n11908;
  assign n12353 = ~n12351 & ~n12352;
  assign n12354 = ~n12350 & n12353;
  assign n12355 = ~n12349 & n12354;
  assign n12356 = pi2  & ~n12355;
  assign n12357 = ~pi2  & n12355;
  assign n12358 = ~n12356 & ~n12357;
  assign n12359 = ~n12348 & n12358;
  assign n12360 = ~n12347 & ~n12359;
  assign n12361 = n12006 & ~n12360;
  assign n12362 = ~n12006 & n12360;
  assign n12363 = ~n1811 & n11288;
  assign n12364 = ~n1740 & n11894;
  assign n12365 = n4951 & n11289;
  assign n12366 = ~n1610 & n11908;
  assign n12367 = ~n12365 & ~n12366;
  assign n12368 = ~n12364 & n12367;
  assign n12369 = ~n12363 & n12368;
  assign n12370 = pi2  & ~n12369;
  assign n12371 = ~pi2  & n12369;
  assign n12372 = ~n12370 & ~n12371;
  assign n12373 = ~n12362 & n12372;
  assign n12374 = ~n12361 & ~n12373;
  assign n12375 = n12004 & ~n12374;
  assign n12376 = ~n12004 & n12374;
  assign n12377 = ~n1740 & n11288;
  assign n12378 = ~n1610 & n11894;
  assign n12379 = n4708 & n11289;
  assign n12380 = ~n1531 & n11908;
  assign n12381 = ~n12379 & ~n12380;
  assign n12382 = ~n12378 & n12381;
  assign n12383 = ~n12377 & n12382;
  assign n12384 = pi2  & ~n12383;
  assign n12385 = ~pi2  & n12383;
  assign n12386 = ~n12384 & ~n12385;
  assign n12387 = ~n12376 & n12386;
  assign n12388 = ~n12375 & ~n12387;
  assign n12389 = ~n12002 & ~n12388;
  assign n12390 = n12002 & n12388;
  assign n12391 = n11848 & ~n11850;
  assign n12392 = ~n11851 & ~n12391;
  assign n12393 = ~n12390 & n12392;
  assign n12394 = ~n12389 & ~n12393;
  assign n12395 = ~n11992 & ~n12394;
  assign n12396 = n11992 & n12394;
  assign n12397 = n11461 & n11852;
  assign n12398 = ~n11853 & ~n12397;
  assign n12399 = ~n12396 & n12398;
  assign n12400 = ~n12395 & ~n12399;
  assign n12401 = ~n11982 & ~n12400;
  assign n12402 = n11982 & n12400;
  assign n12403 = n11445 & n11854;
  assign n12404 = ~n11855 & ~n12403;
  assign n12405 = ~n12402 & n12404;
  assign n12406 = ~n12401 & ~n12405;
  assign n12407 = n11972 & ~n12406;
  assign n12408 = ~n11972 & n12406;
  assign n12409 = ~n1338 & n11288;
  assign n12410 = ~n1230 & n11894;
  assign n12411 = n4323 & n11289;
  assign n12412 = ~n1107 & n11908;
  assign n12413 = ~n12411 & ~n12412;
  assign n12414 = ~n12410 & n12413;
  assign n12415 = ~n12409 & n12414;
  assign n12416 = pi2  & ~n12415;
  assign n12417 = ~pi2  & n12415;
  assign n12418 = ~n12416 & ~n12417;
  assign n12419 = ~n12408 & n12418;
  assign n12420 = ~n12407 & ~n12419;
  assign n12421 = n11970 & ~n12420;
  assign n12422 = ~n11970 & n12420;
  assign n12423 = ~n1230 & n11288;
  assign n12424 = ~n1107 & n11894;
  assign n12425 = n4307 & n11289;
  assign n12426 = ~n1005 & n11908;
  assign n12427 = ~n12425 & ~n12426;
  assign n12428 = ~n12424 & n12427;
  assign n12429 = ~n12423 & n12428;
  assign n12430 = pi2  & ~n12429;
  assign n12431 = ~pi2  & n12429;
  assign n12432 = ~n12430 & ~n12431;
  assign n12433 = ~n12422 & n12432;
  assign n12434 = ~n12421 & ~n12433;
  assign n12435 = ~n11968 & ~n12434;
  assign n12436 = n11968 & n12434;
  assign n12437 = n11403 & n11865;
  assign n12438 = ~n11866 & ~n12437;
  assign n12439 = ~n12436 & n12438;
  assign n12440 = ~n12435 & ~n12439;
  assign n12441 = ~n11958 & ~n12440;
  assign n12442 = ~n11955 & ~n12441;
  assign n12443 = ~n11931 & n11941;
  assign n12444 = ~n11942 & ~n12443;
  assign n12445 = ~n12442 & n12444;
  assign n12446 = ~n11942 & ~n12445;
  assign n12447 = ~n11918 & n11928;
  assign n12448 = ~n11929 & ~n12447;
  assign n12449 = ~n12446 & n12448;
  assign n12450 = ~n11929 & ~n12449;
  assign n12451 = ~n11904 & n11915;
  assign n12452 = ~n11916 & ~n12451;
  assign n12453 = ~n12450 & n12452;
  assign n12454 = ~n11916 & ~n12453;
  assign n12455 = ~n11892 & n11901;
  assign n12456 = ~n11902 & ~n12455;
  assign n12457 = ~n12454 & n12456;
  assign n12458 = ~n11902 & ~n12457;
  assign n12459 = n11890 & ~n12458;
  assign n12460 = ~n11888 & ~n12459;
  assign n12461 = ~n11283 & n11312;
  assign n12462 = ~n11313 & ~n12461;
  assign n12463 = ~n12460 & n12462;
  assign n12464 = ~n11313 & ~n12463;
  assign n12465 = n11278 & ~n11280;
  assign n12466 = ~n11281 & ~n12465;
  assign n12467 = ~n12464 & n12466;
  assign n12468 = ~n11281 & ~n12467;
  assign n12469 = n10725 & ~n12468;
  assign n12470 = ~n10723 & ~n12469;
  assign n12471 = ~n9712 & n10201;
  assign n12472 = ~n10202 & ~n12471;
  assign n12473 = ~n12470 & n12472;
  assign n12474 = ~n10202 & ~n12473;
  assign n12475 = n9707 & ~n9709;
  assign n12476 = ~n9710 & ~n12475;
  assign n12477 = ~n12474 & n12476;
  assign n12478 = ~n9710 & ~n12477;
  assign n12479 = n9261 & ~n12478;
  assign n12480 = ~n9259 & ~n12479;
  assign n12481 = n8845 & ~n12480;
  assign n12482 = ~n8843 & ~n12481;
  assign n12483 = ~n8116 & n8456;
  assign n12484 = ~n8457 & ~n12483;
  assign n12485 = ~n12482 & n12484;
  assign n12486 = ~n8457 & ~n12485;
  assign n12487 = n8114 & ~n12486;
  assign n12488 = ~n8112 & ~n12487;
  assign n12489 = ~n7641 & n7801;
  assign n12490 = ~n7802 & ~n12489;
  assign n12491 = ~n12488 & n12490;
  assign n12492 = ~n7802 & ~n12491;
  assign n12493 = n7636 & ~n7638;
  assign n12494 = ~n7639 & ~n12493;
  assign n12495 = ~n12492 & n12494;
  assign n12496 = ~n7639 & ~n12495;
  assign n12497 = n7483 & ~n12496;
  assign n12498 = ~n7481 & ~n12497;
  assign n12499 = n6967 & ~n12498;
  assign n12500 = ~n6965 & ~n12499;
  assign n12501 = n6822 & ~n12500;
  assign n12502 = ~n6820 & ~n12501;
  assign n12503 = n6539 & ~n12502;
  assign n12504 = ~n6537 & ~n12503;
  assign n12505 = ~n6173 & n6312;
  assign n12506 = ~n6313 & ~n12505;
  assign n12507 = ~n12504 & n12506;
  assign n12508 = ~n6313 & ~n12507;
  assign n12509 = n6171 & ~n12508;
  assign n12510 = ~n6169 & ~n12509;
  assign n12511 = n6067 & ~n12510;
  assign n12512 = ~n6065 & ~n12511;
  assign n12513 = n5623 & ~n12512;
  assign n12514 = ~n5621 & ~n12513;
  assign n12515 = ~n5322 & n5417;
  assign n12516 = ~n5418 & ~n12515;
  assign n12517 = ~n12514 & n12516;
  assign n12518 = ~n5418 & ~n12517;
  assign n12519 = n5320 & ~n12518;
  assign n12520 = ~n5318 & ~n12519;
  assign n12521 = ~n4849 & ~n5253;
  assign n12522 = ~n5254 & ~n12521;
  assign n12523 = ~n12520 & n12522;
  assign n12524 = ~n5254 & ~n12523;
  assign n12525 = n4844 & ~n4846;
  assign n12526 = ~n4847 & ~n12525;
  assign n12527 = ~n12524 & n12526;
  assign n12528 = ~n4847 & ~n12527;
  assign n12529 = n4794 & ~n4796;
  assign n12530 = ~n4797 & ~n12529;
  assign n12531 = ~n12528 & n12530;
  assign n12532 = ~n4797 & ~n12531;
  assign n12533 = n4625 & ~n4627;
  assign n12534 = ~n4628 & ~n12533;
  assign n12535 = ~n12532 & n12534;
  assign n12536 = ~n4628 & ~n12535;
  assign n12537 = n4592 & ~n12536;
  assign n12538 = ~n4590 & ~n12537;
  assign n12539 = n4142 & n4146;
  assign n12540 = ~n4147 & ~n12539;
  assign n12541 = ~n12538 & n12540;
  assign n12542 = ~n4147 & ~n12541;
  assign n12543 = ~n3995 & ~n4026;
  assign n12544 = ~n4027 & ~n12543;
  assign n12545 = ~n12542 & n12544;
  assign n12546 = ~n4027 & ~n12545;
  assign n12547 = n3993 & ~n12546;
  assign n12548 = ~n3991 & ~n12547;
  assign n12549 = n3752 & ~n12548;
  assign n12550 = ~n3750 & ~n12549;
  assign n12551 = ~n3661 & ~n12550;
  assign n12552 = ~n3658 & ~n12551;
  assign n12553 = n2360 & n4096;
  assign n12554 = n306 & n12553;
  assign n12555 = ~n342 & n4894;
  assign n12556 = ~n239 & n12555;
  assign n12557 = n1302 & n1785;
  assign n12558 = ~n330 & n12557;
  assign n12559 = n12556 & n12558;
  assign n12560 = ~n430 & n12559;
  assign n12561 = ~n298 & ~n373;
  assign n12562 = ~n465 & n12561;
  assign n12563 = n1162 & n12562;
  assign n12564 = n12560 & n12563;
  assign n12565 = n1221 & n12564;
  assign n12566 = n974 & n12565;
  assign n12567 = ~n580 & n12566;
  assign n12568 = n12554 & n12567;
  assign n12569 = n1124 & n7184;
  assign n12570 = n2794 & n12569;
  assign n12571 = n1924 & n12570;
  assign n12572 = n1368 & n12571;
  assign n12573 = ~n321 & ~n436;
  assign n12574 = ~n173 & n12573;
  assign n12575 = n3202 & n12574;
  assign n12576 = ~n599 & n12575;
  assign n12577 = ~n114 & n12576;
  assign n12578 = n2502 & n4053;
  assign n12579 = n2320 & n12578;
  assign n12580 = n2585 & n12579;
  assign n12581 = ~n469 & n12580;
  assign n12582 = ~n632 & n12581;
  assign n12583 = n12577 & n12582;
  assign n12584 = n5935 & n12583;
  assign n12585 = ~n612 & ~n682;
  assign n12586 = ~n229 & n12585;
  assign n12587 = ~n280 & ~n309;
  assign n12588 = ~n463 & n12587;
  assign n12589 = n1347 & n12588;
  assign n12590 = n3379 & n12589;
  assign n12591 = ~n243 & n12590;
  assign n12592 = n12586 & n12591;
  assign n12593 = n12584 & n12592;
  assign n12594 = n7143 & n12593;
  assign n12595 = n1635 & n12594;
  assign n12596 = ~n381 & n12595;
  assign n12597 = n12572 & n12596;
  assign n12598 = n12568 & n12597;
  assign n12599 = n551 & n12598;
  assign n12600 = ~n527 & n12599;
  assign n12601 = n3655 & ~n12600;
  assign n12602 = ~n3655 & n12600;
  assign n12603 = ~n12601 & ~n12602;
  assign n12604 = ~n12552 & n12603;
  assign n12605 = n12552 & ~n12603;
  assign n12606 = ~n12604 & ~n12605;
  assign n12607 = n71 & n12606;
  assign n12608 = ~n12600 & n12604;
  assign n12609 = n5326 & ~n12608;
  assign n12610 = n3655 & ~n12604;
  assign n12611 = n12600 & n12610;
  assign n12612 = n12609 & ~n12611;
  assign n12613 = n3661 & n12550;
  assign n12614 = ~n12551 & ~n12613;
  assign n12615 = n5238 & n12614;
  assign n12616 = ~n12608 & ~n12611;
  assign n12617 = ~n12606 & ~n12616;
  assign n12618 = n12606 & ~n12611;
  assign n12619 = ~n12617 & ~n12618;
  assign n12620 = ~n12606 & ~n12614;
  assign n12621 = ~n3752 & n12548;
  assign n12622 = ~n12549 & ~n12621;
  assign n12623 = n12614 & n12622;
  assign n12624 = ~n3993 & n12546;
  assign n12625 = ~n12547 & ~n12624;
  assign n12626 = n12622 & n12625;
  assign n12627 = ~n12622 & ~n12625;
  assign n12628 = ~n12626 & ~n12627;
  assign n12629 = n12542 & ~n12544;
  assign n12630 = ~n12545 & ~n12629;
  assign n12631 = ~n12625 & ~n12630;
  assign n12632 = n12538 & ~n12540;
  assign n12633 = ~n12541 & ~n12632;
  assign n12634 = n12630 & n12633;
  assign n12635 = ~n4592 & n12536;
  assign n12636 = ~n12537 & ~n12635;
  assign n12637 = n12633 & n12636;
  assign n12638 = n12532 & ~n12534;
  assign n12639 = ~n12535 & ~n12638;
  assign n12640 = n12636 & n12639;
  assign n12641 = ~n12636 & ~n12639;
  assign n12642 = ~n12640 & ~n12641;
  assign n12643 = n12528 & ~n12530;
  assign n12644 = ~n12531 & ~n12643;
  assign n12645 = ~n12639 & ~n12644;
  assign n12646 = n12524 & ~n12526;
  assign n12647 = ~n12527 & ~n12646;
  assign n12648 = n12644 & n12647;
  assign n12649 = n12520 & ~n12522;
  assign n12650 = ~n12523 & ~n12649;
  assign n12651 = n12647 & n12650;
  assign n12652 = ~n5320 & n12518;
  assign n12653 = ~n12519 & ~n12652;
  assign n12654 = n12650 & n12653;
  assign n12655 = n12514 & ~n12516;
  assign n12656 = ~n12517 & ~n12655;
  assign n12657 = n12653 & n12656;
  assign n12658 = ~n5623 & n12512;
  assign n12659 = ~n12513 & ~n12658;
  assign n12660 = n12656 & n12659;
  assign n12661 = ~n6067 & n12510;
  assign n12662 = ~n12511 & ~n12661;
  assign n12663 = n12659 & n12662;
  assign n12664 = ~n6171 & n12508;
  assign n12665 = ~n12509 & ~n12664;
  assign n12666 = n12662 & n12665;
  assign n12667 = n12504 & ~n12506;
  assign n12668 = ~n12507 & ~n12667;
  assign n12669 = n12665 & n12668;
  assign n12670 = ~n6539 & n12502;
  assign n12671 = ~n12503 & ~n12670;
  assign n12672 = n12668 & n12671;
  assign n12673 = ~n6822 & n12500;
  assign n12674 = ~n12501 & ~n12673;
  assign n12675 = n12671 & n12674;
  assign n12676 = ~n6967 & n12498;
  assign n12677 = ~n12499 & ~n12676;
  assign n12678 = n12674 & n12677;
  assign n12679 = ~n7483 & n12496;
  assign n12680 = ~n12497 & ~n12679;
  assign n12681 = n12677 & n12680;
  assign n12682 = n12492 & ~n12494;
  assign n12683 = ~n12495 & ~n12682;
  assign n12684 = n12680 & n12683;
  assign n12685 = n12488 & ~n12490;
  assign n12686 = ~n12491 & ~n12685;
  assign n12687 = n12683 & n12686;
  assign n12688 = ~n8114 & n12486;
  assign n12689 = ~n12487 & ~n12688;
  assign n12690 = n12686 & n12689;
  assign n12691 = n12482 & ~n12484;
  assign n12692 = ~n12485 & ~n12691;
  assign n12693 = n12689 & n12692;
  assign n12694 = ~n8845 & n12480;
  assign n12695 = ~n12481 & ~n12694;
  assign n12696 = n12692 & n12695;
  assign n12697 = ~n9261 & n12478;
  assign n12698 = ~n12479 & ~n12697;
  assign n12699 = n12695 & n12698;
  assign n12700 = n12474 & ~n12476;
  assign n12701 = ~n12477 & ~n12700;
  assign n12702 = n12698 & n12701;
  assign n12703 = n12470 & ~n12472;
  assign n12704 = ~n12473 & ~n12703;
  assign n12705 = n12701 & n12704;
  assign n12706 = ~n10725 & n12468;
  assign n12707 = ~n12469 & ~n12706;
  assign n12708 = n12704 & n12707;
  assign n12709 = n12464 & ~n12466;
  assign n12710 = ~n12467 & ~n12709;
  assign n12711 = n12707 & n12710;
  assign n12712 = n12460 & ~n12462;
  assign n12713 = ~n12463 & ~n12712;
  assign n12714 = n12710 & n12713;
  assign n12715 = ~n11890 & n12458;
  assign n12716 = ~n12459 & ~n12715;
  assign n12717 = n12713 & n12716;
  assign n12718 = n12454 & ~n12456;
  assign n12719 = ~n12457 & ~n12718;
  assign n12720 = n12716 & n12719;
  assign n12721 = n12450 & ~n12452;
  assign n12722 = ~n12453 & ~n12721;
  assign n12723 = n12719 & n12722;
  assign n12724 = n12446 & ~n12448;
  assign n12725 = ~n12449 & ~n12724;
  assign n12726 = n12722 & n12725;
  assign n12727 = ~n12722 & ~n12725;
  assign n12728 = ~n12726 & ~n12727;
  assign n12729 = n12442 & ~n12444;
  assign n12730 = ~n12445 & ~n12729;
  assign n12731 = n11958 & n12440;
  assign n12732 = ~n12441 & ~n12731;
  assign n12733 = ~n12725 & ~n12732;
  assign n12734 = n12730 & ~n12733;
  assign n12735 = n12728 & n12734;
  assign n12736 = ~n12726 & ~n12735;
  assign n12737 = ~n12719 & ~n12722;
  assign n12738 = ~n12723 & ~n12737;
  assign n12739 = ~n12736 & n12738;
  assign n12740 = ~n12723 & ~n12739;
  assign n12741 = ~n12716 & ~n12719;
  assign n12742 = ~n12720 & ~n12741;
  assign n12743 = ~n12740 & n12742;
  assign n12744 = ~n12720 & ~n12743;
  assign n12745 = ~n12713 & ~n12716;
  assign n12746 = ~n12717 & ~n12745;
  assign n12747 = ~n12744 & n12746;
  assign n12748 = ~n12717 & ~n12747;
  assign n12749 = ~n12710 & ~n12713;
  assign n12750 = ~n12714 & ~n12749;
  assign n12751 = ~n12748 & n12750;
  assign n12752 = ~n12714 & ~n12751;
  assign n12753 = ~n12707 & ~n12710;
  assign n12754 = ~n12711 & ~n12753;
  assign n12755 = ~n12752 & n12754;
  assign n12756 = ~n12711 & ~n12755;
  assign n12757 = ~n12704 & ~n12707;
  assign n12758 = ~n12708 & ~n12757;
  assign n12759 = ~n12756 & n12758;
  assign n12760 = ~n12708 & ~n12759;
  assign n12761 = ~n12701 & ~n12704;
  assign n12762 = ~n12705 & ~n12761;
  assign n12763 = ~n12760 & n12762;
  assign n12764 = ~n12705 & ~n12763;
  assign n12765 = ~n12698 & ~n12701;
  assign n12766 = ~n12702 & ~n12765;
  assign n12767 = ~n12764 & n12766;
  assign n12768 = ~n12702 & ~n12767;
  assign n12769 = ~n12695 & ~n12698;
  assign n12770 = ~n12699 & ~n12769;
  assign n12771 = ~n12768 & n12770;
  assign n12772 = ~n12699 & ~n12771;
  assign n12773 = ~n12692 & ~n12695;
  assign n12774 = ~n12696 & ~n12773;
  assign n12775 = ~n12772 & n12774;
  assign n12776 = ~n12696 & ~n12775;
  assign n12777 = ~n12689 & ~n12692;
  assign n12778 = ~n12693 & ~n12777;
  assign n12779 = ~n12776 & n12778;
  assign n12780 = ~n12693 & ~n12779;
  assign n12781 = ~n12686 & ~n12689;
  assign n12782 = ~n12690 & ~n12781;
  assign n12783 = ~n12780 & n12782;
  assign n12784 = ~n12690 & ~n12783;
  assign n12785 = ~n12683 & ~n12686;
  assign n12786 = ~n12687 & ~n12785;
  assign n12787 = ~n12784 & n12786;
  assign n12788 = ~n12687 & ~n12787;
  assign n12789 = ~n12680 & ~n12683;
  assign n12790 = ~n12684 & ~n12789;
  assign n12791 = ~n12788 & n12790;
  assign n12792 = ~n12684 & ~n12791;
  assign n12793 = ~n12677 & ~n12680;
  assign n12794 = ~n12681 & ~n12793;
  assign n12795 = ~n12792 & n12794;
  assign n12796 = ~n12681 & ~n12795;
  assign n12797 = ~n12674 & ~n12677;
  assign n12798 = ~n12678 & ~n12797;
  assign n12799 = ~n12796 & n12798;
  assign n12800 = ~n12678 & ~n12799;
  assign n12801 = ~n12671 & ~n12674;
  assign n12802 = ~n12675 & ~n12801;
  assign n12803 = ~n12800 & n12802;
  assign n12804 = ~n12675 & ~n12803;
  assign n12805 = ~n12668 & ~n12671;
  assign n12806 = ~n12672 & ~n12805;
  assign n12807 = ~n12804 & n12806;
  assign n12808 = ~n12672 & ~n12807;
  assign n12809 = ~n12665 & ~n12668;
  assign n12810 = ~n12669 & ~n12809;
  assign n12811 = ~n12808 & n12810;
  assign n12812 = ~n12669 & ~n12811;
  assign n12813 = ~n12662 & ~n12665;
  assign n12814 = ~n12666 & ~n12813;
  assign n12815 = ~n12812 & n12814;
  assign n12816 = ~n12666 & ~n12815;
  assign n12817 = ~n12659 & ~n12662;
  assign n12818 = ~n12663 & ~n12817;
  assign n12819 = ~n12816 & n12818;
  assign n12820 = ~n12663 & ~n12819;
  assign n12821 = ~n12656 & ~n12659;
  assign n12822 = ~n12660 & ~n12821;
  assign n12823 = ~n12820 & n12822;
  assign n12824 = ~n12660 & ~n12823;
  assign n12825 = ~n12653 & ~n12656;
  assign n12826 = ~n12657 & ~n12825;
  assign n12827 = ~n12824 & n12826;
  assign n12828 = ~n12657 & ~n12827;
  assign n12829 = ~n12650 & ~n12653;
  assign n12830 = ~n12654 & ~n12829;
  assign n12831 = ~n12828 & n12830;
  assign n12832 = ~n12654 & ~n12831;
  assign n12833 = ~n12647 & ~n12650;
  assign n12834 = ~n12651 & ~n12833;
  assign n12835 = ~n12832 & n12834;
  assign n12836 = ~n12651 & ~n12835;
  assign n12837 = ~n12644 & ~n12647;
  assign n12838 = ~n12648 & ~n12837;
  assign n12839 = ~n12836 & n12838;
  assign n12840 = ~n12648 & ~n12839;
  assign n12841 = n12639 & n12644;
  assign n12842 = n12840 & ~n12841;
  assign n12843 = ~n12645 & ~n12842;
  assign n12844 = n12642 & n12843;
  assign n12845 = ~n12640 & ~n12844;
  assign n12846 = ~n12633 & ~n12636;
  assign n12847 = ~n12637 & ~n12846;
  assign n12848 = ~n12845 & n12847;
  assign n12849 = ~n12637 & ~n12848;
  assign n12850 = ~n12630 & ~n12633;
  assign n12851 = ~n12634 & ~n12850;
  assign n12852 = ~n12849 & n12851;
  assign n12853 = ~n12634 & ~n12852;
  assign n12854 = n12625 & n12630;
  assign n12855 = n12853 & ~n12854;
  assign n12856 = ~n12631 & ~n12855;
  assign n12857 = n12628 & n12856;
  assign n12858 = ~n12626 & ~n12857;
  assign n12859 = ~n12614 & ~n12622;
  assign n12860 = ~n12623 & ~n12859;
  assign n12861 = ~n12858 & n12860;
  assign n12862 = ~n12623 & ~n12861;
  assign n12863 = n12606 & n12614;
  assign n12864 = n12862 & ~n12863;
  assign n12865 = ~n12620 & ~n12864;
  assign n12866 = n12619 & n12865;
  assign n12867 = ~n12619 & ~n12865;
  assign n12868 = ~n12866 & ~n12867;
  assign n12869 = n5239 & n12868;
  assign n12870 = ~n12615 & ~n12869;
  assign n12871 = ~n12612 & n12870;
  assign n12872 = ~n12607 & n12871;
  assign n12873 = pi23  & n12872;
  assign n12874 = ~pi23  & ~n12872;
  assign n12875 = ~n12873 & ~n12874;
  assign n12876 = ~n394 & n2436;
  assign n12877 = ~n150 & ~n181;
  assign n12878 = n1341 & n12877;
  assign n12879 = ~n213 & n12878;
  assign n12880 = n12876 & n12879;
  assign n12881 = ~n457 & n12880;
  assign n12882 = ~n361 & n5116;
  assign n12883 = ~n344 & n12882;
  assign n12884 = ~n671 & n12883;
  assign n12885 = n12881 & n12884;
  assign n12886 = ~n104 & n3724;
  assign n12887 = ~n341 & n2836;
  assign n12888 = ~n414 & n12887;
  assign n12889 = n12886 & n12888;
  assign n12890 = ~n633 & n12889;
  assign n12891 = ~n468 & n12890;
  assign n12892 = n858 & n3159;
  assign n12893 = ~n473 & n5670;
  assign n12894 = n12892 & n12893;
  assign n12895 = ~n81 & n2566;
  assign n12896 = ~n439 & n12895;
  assign n12897 = ~n356 & n12896;
  assign n12898 = ~n610 & n7062;
  assign n12899 = ~n116 & ~n129;
  assign n12900 = n12898 & n12899;
  assign n12901 = n2772 & n12900;
  assign n12902 = n12897 & n12901;
  assign n12903 = n12894 & n12902;
  assign n12904 = n12891 & n12903;
  assign n12905 = n12885 & n12904;
  assign n12906 = ~n259 & n12905;
  assign n12907 = ~n197 & ~n613;
  assign n12908 = ~n704 & n12907;
  assign n12909 = n1417 & n2060;
  assign n12910 = ~n390 & n12909;
  assign n12911 = n12908 & n12910;
  assign n12912 = n1934 & n12911;
  assign n12913 = ~n323 & n12912;
  assign n12914 = n12906 & n12913;
  assign n12915 = ~n216 & ~n534;
  assign n12916 = ~n360 & n12915;
  assign n12917 = ~n278 & ~n621;
  assign n12918 = ~n579 & n12917;
  assign n12919 = ~n289 & n12918;
  assign n12920 = ~n272 & n12919;
  assign n12921 = n12916 & n12920;
  assign n12922 = n2088 & n3195;
  assign n12923 = n12921 & n12922;
  assign n12924 = ~n582 & n12923;
  assign n12925 = n1247 & n1581;
  assign n12926 = n3338 & n12925;
  assign n12927 = n5105 & n12926;
  assign n12928 = ~n114 & n12927;
  assign n12929 = n12924 & n12928;
  assign n12930 = n12914 & n12929;
  assign n12931 = n754 & n5918;
  assign n12932 = n148 & n12931;
  assign n12933 = ~n236 & n12932;
  assign n12934 = ~n259 & ~n290;
  assign n12935 = n2184 & n3170;
  assign n12936 = n1182 & n12935;
  assign n12937 = n12934 & n12936;
  assign n12938 = ~n439 & n12937;
  assign n12939 = n12933 & n12938;
  assign n12940 = n3076 & n3820;
  assign n12941 = ~n298 & n12940;
  assign n12942 = ~n600 & n12941;
  assign n12943 = ~n423 & ~n681;
  assign n12944 = n3443 & n12943;
  assign n12945 = ~n536 & n12944;
  assign n12946 = ~n373 & ~n627;
  assign n12947 = ~n612 & n12946;
  assign n12948 = n12945 & n12947;
  assign n12949 = n402 & n12948;
  assign n12950 = n4422 & n12949;
  assign n12951 = n1246 & n12950;
  assign n12952 = ~n385 & n12951;
  assign n12953 = ~n501 & n12952;
  assign n12954 = n12942 & n12953;
  assign n12955 = n12939 & n12954;
  assign n12956 = ~n228 & n322;
  assign n12957 = ~n382 & n12956;
  assign n12958 = n3422 & n12957;
  assign n12959 = n2409 & n12958;
  assign n12960 = n3138 & n12959;
  assign n12961 = ~n668 & n12960;
  assign n12962 = n5482 & n7197;
  assign n12963 = n237 & n12962;
  assign n12964 = ~n129 & n12963;
  assign n12965 = n12961 & n12964;
  assign n12966 = n3330 & n3678;
  assign n12967 = ~n165 & n12966;
  assign n12968 = ~n298 & ~n424;
  assign n12969 = ~n315 & n12968;
  assign n12970 = ~n462 & n12969;
  assign n12971 = n12885 & n12970;
  assign n12972 = n2218 & n12971;
  assign n12973 = ~n633 & n12972;
  assign n12974 = n12967 & n12973;
  assign n12975 = n12965 & n12974;
  assign n12976 = ~n12955 & ~n12975;
  assign n12977 = n6176 & n6183;
  assign n12978 = ~n12608 & ~n12977;
  assign n12979 = pi17  & ~n12978;
  assign n12980 = ~pi17  & n12978;
  assign n12981 = ~n12979 & ~n12980;
  assign n12982 = n12955 & n12975;
  assign n12983 = ~n12976 & ~n12982;
  assign n12984 = n12981 & n12983;
  assign n12985 = ~n12976 & ~n12984;
  assign n12986 = n12930 & ~n12985;
  assign n12987 = ~n12930 & n12985;
  assign n12988 = ~n12986 & ~n12987;
  assign n12989 = n3641 & n12656;
  assign n12990 = n12828 & ~n12830;
  assign n12991 = ~n12831 & ~n12990;
  assign n12992 = n556 & n12991;
  assign n12993 = n3961 & n12650;
  assign n12994 = n3740 & n12653;
  assign n12995 = ~n12993 & ~n12994;
  assign n12996 = ~n12992 & n12995;
  assign n12997 = ~n12989 & n12996;
  assign n12998 = n12988 & ~n12997;
  assign n12999 = ~n12986 & ~n12998;
  assign n13000 = n2045 & n2735;
  assign n13001 = n1232 & n13000;
  assign n13002 = ~n704 & n13001;
  assign n13003 = ~n390 & n13002;
  assign n13004 = ~n598 & ~n669;
  assign n13005 = ~n701 & n1755;
  assign n13006 = n13004 & n13005;
  assign n13007 = n2345 & n13006;
  assign n13008 = ~n518 & n13007;
  assign n13009 = ~n163 & n13008;
  assign n13010 = ~n81 & n13009;
  assign n13011 = n13003 & n13010;
  assign n13012 = ~n186 & n13011;
  assign n13013 = n355 & n5858;
  assign n13014 = n758 & n13013;
  assign n13015 = n1222 & n1720;
  assign n13016 = ~n281 & n13015;
  assign n13017 = ~n383 & n13016;
  assign n13018 = n2585 & n2726;
  assign n13019 = ~n203 & n13018;
  assign n13020 = ~n170 & n13019;
  assign n13021 = n13017 & n13020;
  assign n13022 = n694 & n3479;
  assign n13023 = ~n166 & n13022;
  assign n13024 = ~n612 & n13023;
  assign n13025 = n998 & n1902;
  assign n13026 = ~n442 & n13025;
  assign n13027 = ~n361 & n13026;
  assign n13028 = n13024 & n13027;
  assign n13029 = n13021 & n13028;
  assign n13030 = n5091 & n13029;
  assign n13031 = n2066 & n13030;
  assign n13032 = n13014 & n13031;
  assign n13033 = ~n207 & n13032;
  assign n13034 = n3770 & n13033;
  assign n13035 = n13012 & n13034;
  assign n13036 = n12930 & ~n13035;
  assign n13037 = ~n12930 & n13035;
  assign n13038 = ~n13036 & ~n13037;
  assign n13039 = n3641 & n12653;
  assign n13040 = n3740 & n12650;
  assign n13041 = n12832 & ~n12834;
  assign n13042 = ~n12835 & ~n13041;
  assign n13043 = n556 & n13042;
  assign n13044 = n3961 & n12647;
  assign n13045 = ~n13043 & ~n13044;
  assign n13046 = ~n13040 & n13045;
  assign n13047 = ~n13039 & n13046;
  assign n13048 = n13038 & ~n13047;
  assign n13049 = ~n13038 & n13047;
  assign n13050 = ~n13048 & ~n13049;
  assign n13051 = ~n12999 & n13050;
  assign n13052 = n12999 & ~n13050;
  assign n13053 = ~n13051 & ~n13052;
  assign n13054 = ~n12981 & ~n12983;
  assign n13055 = ~n12984 & ~n13054;
  assign n13056 = n3641 & n12659;
  assign n13057 = n3740 & n12656;
  assign n13058 = n12824 & ~n12826;
  assign n13059 = ~n12827 & ~n13058;
  assign n13060 = n556 & n13059;
  assign n13061 = n3961 & n12653;
  assign n13062 = ~n13060 & ~n13061;
  assign n13063 = ~n13057 & n13062;
  assign n13064 = ~n13056 & n13063;
  assign n13065 = n13055 & ~n13064;
  assign n13066 = n2694 & n3386;
  assign n13067 = n1902 & n13066;
  assign n13068 = ~n262 & n13067;
  assign n13069 = ~n278 & ~n473;
  assign n13070 = ~n697 & n5138;
  assign n13071 = ~n350 & n6624;
  assign n13072 = n13070 & n13071;
  assign n13073 = ~n152 & ~n247;
  assign n13074 = n4444 & n13073;
  assign n13075 = ~n307 & n13074;
  assign n13076 = ~n114 & n13075;
  assign n13077 = ~n254 & ~n590;
  assign n13078 = ~n631 & n13077;
  assign n13079 = ~n548 & ~n614;
  assign n13080 = ~n279 & n13079;
  assign n13081 = n13078 & n13080;
  assign n13082 = n2180 & n13081;
  assign n13083 = ~n207 & n13082;
  assign n13084 = ~n181 & n13083;
  assign n13085 = n13076 & n13084;
  assign n13086 = n13072 & n13085;
  assign n13087 = n13069 & n13086;
  assign n13088 = n3478 & n13087;
  assign n13089 = ~n581 & n13088;
  assign n13090 = n2140 & n13089;
  assign n13091 = n3215 & n13090;
  assign n13092 = ~n242 & n13091;
  assign n13093 = ~n682 & n13092;
  assign n13094 = n13068 & n13093;
  assign n13095 = n2409 & n3870;
  assign n13096 = ~n690 & n13095;
  assign n13097 = ~n260 & n13096;
  assign n13098 = ~n629 & n1347;
  assign n13099 = ~n601 & n13098;
  assign n13100 = ~n331 & n13099;
  assign n13101 = n1285 & n2070;
  assign n13102 = ~n398 & n13101;
  assign n13103 = n300 & ~n583;
  assign n13104 = ~n341 & n13103;
  assign n13105 = n13102 & n13104;
  assign n13106 = ~n439 & n13105;
  assign n13107 = n13100 & n13106;
  assign n13108 = n558 & n13107;
  assign n13109 = ~n228 & n13108;
  assign n13110 = ~n85 & n13109;
  assign n13111 = n13097 & n13110;
  assign n13112 = n13094 & n13111;
  assign n13113 = n12955 & ~n13112;
  assign n13114 = n2593 & n4373;
  assign n13115 = ~n454 & n13114;
  assign n13116 = ~n163 & n2180;
  assign n13117 = ~n672 & n2416;
  assign n13118 = ~n325 & n13117;
  assign n13119 = n13116 & n13118;
  assign n13120 = n2635 & n13119;
  assign n13121 = ~n246 & n13120;
  assign n13122 = ~n281 & n13121;
  assign n13123 = n13115 & n13122;
  assign n13124 = n2105 & n5097;
  assign n13125 = n7060 & n13124;
  assign n13126 = ~n697 & n13125;
  assign n13127 = ~n231 & n13126;
  assign n13128 = n921 & n1659;
  assign n13129 = n1497 & n13128;
  assign n13130 = n1652 & n13129;
  assign n13131 = ~n391 & n13130;
  assign n13132 = ~n132 & n13131;
  assign n13133 = n13127 & n13132;
  assign n13134 = n13123 & n13133;
  assign n13135 = ~n633 & n5759;
  assign n13136 = ~n354 & n13135;
  assign n13137 = n3464 & n13136;
  assign n13138 = ~n332 & n13137;
  assign n13139 = ~n413 & n13138;
  assign n13140 = n759 & n1985;
  assign n13141 = ~n390 & n13140;
  assign n13142 = ~n78 & n13141;
  assign n13143 = n13139 & n13142;
  assign n13144 = n860 & n13143;
  assign n13145 = n1146 & n3897;
  assign n13146 = ~n590 & n13145;
  assign n13147 = ~n455 & n13146;
  assign n13148 = n5924 & n13147;
  assign n13149 = n13144 & n13148;
  assign n13150 = ~n13134 & ~n13149;
  assign n13151 = n6827 & n6834;
  assign n13152 = ~n12608 & ~n13151;
  assign n13153 = pi14  & ~n13152;
  assign n13154 = ~pi14  & n13152;
  assign n13155 = ~n13153 & ~n13154;
  assign n13156 = n13134 & n13149;
  assign n13157 = ~n13150 & ~n13156;
  assign n13158 = n13155 & n13157;
  assign n13159 = ~n13150 & ~n13158;
  assign n13160 = n13112 & ~n13159;
  assign n13161 = ~n13112 & n13159;
  assign n13162 = ~n13160 & ~n13161;
  assign n13163 = n3641 & n12665;
  assign n13164 = n12816 & ~n12818;
  assign n13165 = ~n12819 & ~n13164;
  assign n13166 = n556 & n13165;
  assign n13167 = n3961 & n12659;
  assign n13168 = n3740 & n12662;
  assign n13169 = ~n13167 & ~n13168;
  assign n13170 = ~n13166 & n13169;
  assign n13171 = ~n13163 & n13170;
  assign n13172 = n13162 & ~n13171;
  assign n13173 = ~n13160 & ~n13172;
  assign n13174 = ~n12955 & n13112;
  assign n13175 = ~n13113 & ~n13174;
  assign n13176 = ~n13173 & n13175;
  assign n13177 = ~n13113 & ~n13176;
  assign n13178 = n13055 & n13064;
  assign n13179 = ~n13055 & ~n13064;
  assign n13180 = ~n13178 & ~n13179;
  assign n13181 = ~n13177 & ~n13180;
  assign n13182 = ~n13065 & ~n13181;
  assign n13183 = ~n12988 & n12997;
  assign n13184 = ~n12998 & ~n13183;
  assign n13185 = ~n13182 & n13184;
  assign n13186 = n13182 & ~n13184;
  assign n13187 = ~n13185 & ~n13186;
  assign n13188 = n4006 & n12647;
  assign n13189 = n4133 & n12644;
  assign n13190 = ~n12645 & ~n12841;
  assign n13191 = n12840 & n13190;
  assign n13192 = ~n12840 & ~n13190;
  assign n13193 = ~n13191 & ~n13192;
  assign n13194 = n4002 & ~n13193;
  assign n13195 = n4555 & n12639;
  assign n13196 = ~n13194 & ~n13195;
  assign n13197 = ~n13189 & n13196;
  assign n13198 = ~n13188 & n13197;
  assign n13199 = pi29  & n13198;
  assign n13200 = ~pi29  & ~n13198;
  assign n13201 = ~n13199 & ~n13200;
  assign n13202 = n13187 & ~n13201;
  assign n13203 = ~n13185 & ~n13202;
  assign n13204 = n13053 & ~n13203;
  assign n13205 = ~n13053 & n13203;
  assign n13206 = ~n13204 & ~n13205;
  assign n13207 = n4006 & n12644;
  assign n13208 = n4133 & n12639;
  assign n13209 = ~n12642 & ~n12843;
  assign n13210 = ~n12844 & ~n13209;
  assign n13211 = n4002 & n13210;
  assign n13212 = n4555 & n12636;
  assign n13213 = ~n13211 & ~n13212;
  assign n13214 = ~n13208 & n13213;
  assign n13215 = ~n13207 & n13214;
  assign n13216 = pi29  & n13215;
  assign n13217 = ~pi29  & ~n13215;
  assign n13218 = ~n13216 & ~n13217;
  assign n13219 = n13206 & n13218;
  assign n13220 = ~n13206 & ~n13218;
  assign n13221 = ~n13219 & ~n13220;
  assign n13222 = n4601 & n12633;
  assign n13223 = n4783 & n12630;
  assign n13224 = ~n12631 & ~n12854;
  assign n13225 = n12853 & n13224;
  assign n13226 = ~n12853 & ~n13224;
  assign n13227 = ~n13225 & ~n13226;
  assign n13228 = n4602 & ~n13227;
  assign n13229 = n4801 & n12625;
  assign n13230 = ~n13228 & ~n13229;
  assign n13231 = ~n13223 & n13230;
  assign n13232 = ~n13222 & n13231;
  assign n13233 = pi26  & n13232;
  assign n13234 = ~pi26  & ~n13232;
  assign n13235 = ~n13233 & ~n13234;
  assign n13236 = ~n13221 & ~n13235;
  assign n13237 = n13221 & n13235;
  assign n13238 = ~n13236 & ~n13237;
  assign n13239 = ~n13187 & n13201;
  assign n13240 = ~n13202 & ~n13239;
  assign n13241 = n13173 & ~n13175;
  assign n13242 = ~n13176 & ~n13241;
  assign n13243 = n3641 & n12662;
  assign n13244 = n3740 & n12659;
  assign n13245 = n12820 & ~n12822;
  assign n13246 = ~n12823 & ~n13245;
  assign n13247 = n556 & n13246;
  assign n13248 = n3961 & n12656;
  assign n13249 = ~n13247 & ~n13248;
  assign n13250 = ~n13244 & n13249;
  assign n13251 = ~n13243 & n13250;
  assign n13252 = n13242 & ~n13251;
  assign n13253 = n13242 & n13251;
  assign n13254 = ~n13242 & ~n13251;
  assign n13255 = ~n13253 & ~n13254;
  assign n13256 = n4006 & n12653;
  assign n13257 = n4133 & n12650;
  assign n13258 = n4002 & n13042;
  assign n13259 = n4555 & n12647;
  assign n13260 = ~n13258 & ~n13259;
  assign n13261 = ~n13257 & n13260;
  assign n13262 = ~n13256 & n13261;
  assign n13263 = pi29  & n13262;
  assign n13264 = ~pi29  & ~n13262;
  assign n13265 = ~n13263 & ~n13264;
  assign n13266 = ~n13255 & ~n13265;
  assign n13267 = ~n13252 & ~n13266;
  assign n13268 = n13177 & ~n13180;
  assign n13269 = ~n13177 & n13180;
  assign n13270 = ~n13268 & ~n13269;
  assign n13271 = ~n13267 & ~n13270;
  assign n13272 = n4006 & n12650;
  assign n13273 = n4133 & n12647;
  assign n13274 = n12836 & ~n12838;
  assign n13275 = ~n12839 & ~n13274;
  assign n13276 = n4002 & n13275;
  assign n13277 = n4555 & n12644;
  assign n13278 = ~n13276 & ~n13277;
  assign n13279 = ~n13273 & n13278;
  assign n13280 = ~n13272 & n13279;
  assign n13281 = pi29  & n13280;
  assign n13282 = ~pi29  & ~n13280;
  assign n13283 = ~n13281 & ~n13282;
  assign n13284 = n13267 & n13270;
  assign n13285 = ~n13283 & ~n13284;
  assign n13286 = ~n13271 & ~n13285;
  assign n13287 = n13240 & ~n13286;
  assign n13288 = ~n13240 & n13286;
  assign n13289 = n4601 & n12636;
  assign n13290 = n4783 & n12633;
  assign n13291 = n12849 & ~n12851;
  assign n13292 = ~n12852 & ~n13291;
  assign n13293 = n4602 & n13292;
  assign n13294 = n4801 & n12630;
  assign n13295 = ~n13293 & ~n13294;
  assign n13296 = ~n13290 & n13295;
  assign n13297 = ~n13289 & n13296;
  assign n13298 = pi26  & n13297;
  assign n13299 = ~pi26  & ~n13297;
  assign n13300 = ~n13298 & ~n13299;
  assign n13301 = ~n13288 & ~n13300;
  assign n13302 = ~n13287 & ~n13301;
  assign n13303 = n13238 & ~n13302;
  assign n13304 = ~n13238 & n13302;
  assign n13305 = n5238 & n12622;
  assign n13306 = n71 & n12614;
  assign n13307 = ~n12620 & ~n12863;
  assign n13308 = n12862 & n13307;
  assign n13309 = ~n12862 & ~n13307;
  assign n13310 = ~n13308 & ~n13309;
  assign n13311 = n5239 & ~n13310;
  assign n13312 = n5326 & n12606;
  assign n13313 = ~n13311 & ~n13312;
  assign n13314 = ~n13306 & n13313;
  assign n13315 = ~n13305 & n13314;
  assign n13316 = pi23  & n13315;
  assign n13317 = ~pi23  & ~n13315;
  assign n13318 = ~n13316 & ~n13317;
  assign n13319 = ~n13304 & ~n13318;
  assign n13320 = ~n13303 & ~n13319;
  assign n13321 = ~n12875 & ~n13320;
  assign n13322 = n4601 & n12630;
  assign n13323 = n4783 & n12625;
  assign n13324 = ~n12628 & ~n12856;
  assign n13325 = ~n12857 & ~n13324;
  assign n13326 = n4602 & n13325;
  assign n13327 = n4801 & n12622;
  assign n13328 = ~n13326 & ~n13327;
  assign n13329 = ~n13323 & n13328;
  assign n13330 = ~n13322 & n13329;
  assign n13331 = pi26  & n13330;
  assign n13332 = ~pi26  & ~n13330;
  assign n13333 = ~n13331 & ~n13332;
  assign n13334 = ~n13051 & ~n13204;
  assign n13335 = n5428 & n5434;
  assign n13336 = ~n12608 & ~n13335;
  assign n13337 = pi20  & ~n13336;
  assign n13338 = ~pi20  & n13336;
  assign n13339 = ~n13337 & ~n13338;
  assign n13340 = n1617 & n2524;
  assign n13341 = n1775 & n13340;
  assign n13342 = ~n399 & n13341;
  assign n13343 = n1851 & n4472;
  assign n13344 = ~n461 & n13343;
  assign n13345 = ~n220 & n13344;
  assign n13346 = n13342 & n13345;
  assign n13347 = n1605 & n3439;
  assign n13348 = ~n681 & n13347;
  assign n13349 = ~n692 & n13348;
  assign n13350 = ~n695 & n2066;
  assign n13351 = n1348 & n2156;
  assign n13352 = n949 & n1366;
  assign n13353 = n13351 & n13352;
  assign n13354 = ~n693 & n13353;
  assign n13355 = n1409 & n3326;
  assign n13356 = ~n260 & n13355;
  assign n13357 = n2642 & n5704;
  assign n13358 = ~n697 & n13357;
  assign n13359 = ~n85 & n13358;
  assign n13360 = n13356 & n13359;
  assign n13361 = n13354 & n13360;
  assign n13362 = n13350 & n13361;
  assign n13363 = n1577 & n13362;
  assign n13364 = n1513 & n13363;
  assign n13365 = ~n401 & n13364;
  assign n13366 = ~n457 & n13365;
  assign n13367 = n13349 & n13366;
  assign n13368 = n13346 & n13367;
  assign n13369 = n12930 & n13368;
  assign n13370 = ~n12930 & ~n13368;
  assign n13371 = ~n13369 & ~n13370;
  assign n13372 = n13339 & n13371;
  assign n13373 = ~n13339 & ~n13371;
  assign n13374 = ~n13372 & ~n13373;
  assign n13375 = ~n13037 & ~n13047;
  assign n13376 = ~n13036 & ~n13375;
  assign n13377 = n13374 & ~n13376;
  assign n13378 = ~n13374 & n13376;
  assign n13379 = ~n13377 & ~n13378;
  assign n13380 = n3641 & n12650;
  assign n13381 = n3740 & n12647;
  assign n13382 = n556 & n13275;
  assign n13383 = n3961 & n12644;
  assign n13384 = ~n13382 & ~n13383;
  assign n13385 = ~n13381 & n13384;
  assign n13386 = ~n13380 & n13385;
  assign n13387 = n13379 & ~n13386;
  assign n13388 = ~n13379 & n13386;
  assign n13389 = ~n13387 & ~n13388;
  assign n13390 = ~n13334 & n13389;
  assign n13391 = n13334 & ~n13389;
  assign n13392 = ~n13390 & ~n13391;
  assign n13393 = n4006 & n12639;
  assign n13394 = n4133 & n12636;
  assign n13395 = n12845 & ~n12847;
  assign n13396 = ~n12848 & ~n13395;
  assign n13397 = n4002 & n13396;
  assign n13398 = n4555 & n12633;
  assign n13399 = ~n13397 & ~n13398;
  assign n13400 = ~n13394 & n13399;
  assign n13401 = ~n13393 & n13400;
  assign n13402 = pi29  & n13401;
  assign n13403 = ~pi29  & ~n13401;
  assign n13404 = ~n13402 & ~n13403;
  assign n13405 = n13392 & ~n13404;
  assign n13406 = ~n13392 & n13404;
  assign n13407 = ~n13405 & ~n13406;
  assign n13408 = n13333 & n13407;
  assign n13409 = ~n13333 & ~n13407;
  assign n13410 = ~n13408 & ~n13409;
  assign n13411 = n13206 & ~n13218;
  assign n13412 = ~n13236 & ~n13411;
  assign n13413 = ~n13410 & ~n13412;
  assign n13414 = n13410 & n13412;
  assign n13415 = ~n13413 & ~n13414;
  assign n13416 = n12875 & ~n13320;
  assign n13417 = ~n12875 & n13320;
  assign n13418 = ~n13416 & ~n13417;
  assign n13419 = n13415 & ~n13418;
  assign n13420 = ~n13321 & ~n13419;
  assign n13421 = ~n13333 & n13407;
  assign n13422 = ~n13413 & ~n13421;
  assign n13423 = ~n13370 & ~n13372;
  assign n13424 = n12593 & ~n13423;
  assign n13425 = ~n12593 & n13423;
  assign n13426 = ~n13424 & ~n13425;
  assign n13427 = n3641 & n12647;
  assign n13428 = n556 & ~n13193;
  assign n13429 = n3961 & n12639;
  assign n13430 = n3740 & n12644;
  assign n13431 = ~n13429 & ~n13430;
  assign n13432 = ~n13428 & n13431;
  assign n13433 = ~n13427 & n13432;
  assign n13434 = n13426 & ~n13433;
  assign n13435 = ~n13426 & n13433;
  assign n13436 = ~n13434 & ~n13435;
  assign n13437 = ~n13378 & ~n13386;
  assign n13438 = ~n13377 & ~n13437;
  assign n13439 = n13436 & ~n13438;
  assign n13440 = ~n13436 & n13438;
  assign n13441 = ~n13439 & ~n13440;
  assign n13442 = n4006 & n12636;
  assign n13443 = n4133 & n12633;
  assign n13444 = n4002 & n13292;
  assign n13445 = n4555 & n12630;
  assign n13446 = ~n13444 & ~n13445;
  assign n13447 = ~n13443 & n13446;
  assign n13448 = ~n13442 & n13447;
  assign n13449 = pi29  & n13448;
  assign n13450 = ~pi29  & ~n13448;
  assign n13451 = ~n13449 & ~n13450;
  assign n13452 = n13441 & ~n13451;
  assign n13453 = ~n13441 & n13451;
  assign n13454 = ~n13452 & ~n13453;
  assign n13455 = ~n13391 & ~n13404;
  assign n13456 = ~n13390 & ~n13455;
  assign n13457 = n13454 & ~n13456;
  assign n13458 = ~n13454 & n13456;
  assign n13459 = ~n13457 & ~n13458;
  assign n13460 = n4601 & n12625;
  assign n13461 = n4783 & n12622;
  assign n13462 = n12858 & ~n12860;
  assign n13463 = ~n12861 & ~n13462;
  assign n13464 = n4602 & n13463;
  assign n13465 = n4801 & n12614;
  assign n13466 = ~n13464 & ~n13465;
  assign n13467 = ~n13461 & n13466;
  assign n13468 = ~n13460 & n13467;
  assign n13469 = pi26  & n13468;
  assign n13470 = ~pi26  & ~n13468;
  assign n13471 = ~n13469 & ~n13470;
  assign n13472 = n13459 & ~n13471;
  assign n13473 = ~n13459 & n13471;
  assign n13474 = ~n13472 & ~n13473;
  assign n13475 = ~n13422 & n13474;
  assign n13476 = n13422 & ~n13474;
  assign n13477 = ~n13475 & ~n13476;
  assign n13478 = n5238 & n12606;
  assign n13479 = n71 & n12616;
  assign n13480 = n12611 & n12866;
  assign n13481 = ~n12611 & ~n12866;
  assign n13482 = ~n13480 & ~n13481;
  assign n13483 = ~n12618 & ~n13482;
  assign n13484 = n5239 & ~n13483;
  assign n13485 = ~n12609 & ~n13484;
  assign n13486 = ~n13479 & n13485;
  assign n13487 = ~n13478 & n13486;
  assign n13488 = pi23  & n13487;
  assign n13489 = ~pi23  & ~n13487;
  assign n13490 = ~n13488 & ~n13489;
  assign n13491 = n13477 & ~n13490;
  assign n13492 = ~n13477 & n13490;
  assign n13493 = ~n13491 & ~n13492;
  assign n13494 = n13420 & n13493;
  assign n13495 = ~n13420 & ~n13493;
  assign n13496 = ~n13494 & ~n13495;
  assign n13497 = ~n13415 & n13418;
  assign n13498 = ~n13419 & ~n13497;
  assign n13499 = ~n12616 & ~n13480;
  assign n13500 = n5429 & ~n13499;
  assign n13501 = n5435 & ~n12611;
  assign n13502 = ~n5429 & ~n5434;
  assign n13503 = ~n13501 & ~n13502;
  assign n13504 = ~n12608 & ~n13503;
  assign n13505 = ~n13500 & ~n13504;
  assign n13506 = pi20  & n13505;
  assign n13507 = ~pi20  & ~n13505;
  assign n13508 = ~n13506 & ~n13507;
  assign n13509 = n4601 & n12639;
  assign n13510 = n4783 & n12636;
  assign n13511 = n4602 & n13396;
  assign n13512 = n4801 & n12633;
  assign n13513 = ~n13511 & ~n13512;
  assign n13514 = ~n13510 & n13513;
  assign n13515 = ~n13509 & n13514;
  assign n13516 = pi26  & n13515;
  assign n13517 = ~pi26  & ~n13515;
  assign n13518 = ~n13516 & ~n13517;
  assign n13519 = ~n13271 & ~n13284;
  assign n13520 = n13283 & ~n13519;
  assign n13521 = ~n13283 & n13519;
  assign n13522 = ~n13520 & ~n13521;
  assign n13523 = ~n13518 & n13522;
  assign n13524 = n13518 & n13522;
  assign n13525 = ~n13518 & ~n13522;
  assign n13526 = ~n13524 & ~n13525;
  assign n13527 = ~n13162 & n13171;
  assign n13528 = ~n13172 & ~n13527;
  assign n13529 = ~n13155 & ~n13157;
  assign n13530 = ~n13158 & ~n13529;
  assign n13531 = ~n612 & n2566;
  assign n13532 = n768 & n1859;
  assign n13533 = n814 & n4456;
  assign n13534 = ~n197 & n13533;
  assign n13535 = ~n154 & n13534;
  assign n13536 = n13532 & n13535;
  assign n13537 = ~n216 & n13536;
  assign n13538 = n13531 & n13537;
  assign n13539 = n1513 & n13538;
  assign n13540 = n797 & n13539;
  assign n13541 = ~n294 & n13540;
  assign n13542 = ~n544 & n13541;
  assign n13543 = n1484 & n3009;
  assign n13544 = n519 & n13543;
  assign n13545 = n4888 & n13544;
  assign n13546 = n2654 & n13545;
  assign n13547 = n13542 & n13546;
  assign n13548 = n2833 & n4162;
  assign n13549 = ~n502 & n13548;
  assign n13550 = ~n441 & n13549;
  assign n13551 = ~n238 & n706;
  assign n13552 = ~n247 & n4238;
  assign n13553 = ~n383 & n13552;
  assign n13554 = ~n288 & ~n537;
  assign n13555 = n13553 & n13554;
  assign n13556 = n1169 & n13555;
  assign n13557 = n1587 & n13556;
  assign n13558 = n1912 & n13557;
  assign n13559 = ~n631 & n13558;
  assign n13560 = n1224 & n1783;
  assign n13561 = n1652 & n3855;
  assign n13562 = n13560 & n13561;
  assign n13563 = n810 & n13562;
  assign n13564 = ~n106 & n13563;
  assign n13565 = n13559 & n13564;
  assign n13566 = ~n357 & n13565;
  assign n13567 = n13551 & n13566;
  assign n13568 = n2340 & n13567;
  assign n13569 = ~n398 & n13568;
  assign n13570 = ~n231 & n13569;
  assign n13571 = n13550 & n13570;
  assign n13572 = n13547 & n13571;
  assign n13573 = n13149 & ~n13572;
  assign n13574 = ~n13149 & n13572;
  assign n13575 = n3641 & n12671;
  assign n13576 = n3740 & n12668;
  assign n13577 = n12808 & ~n12810;
  assign n13578 = ~n12811 & ~n13577;
  assign n13579 = n556 & n13578;
  assign n13580 = n3961 & n12665;
  assign n13581 = ~n13579 & ~n13580;
  assign n13582 = ~n13576 & n13581;
  assign n13583 = ~n13575 & n13582;
  assign n13584 = ~n13574 & ~n13583;
  assign n13585 = ~n13573 & ~n13584;
  assign n13586 = n13530 & ~n13585;
  assign n13587 = ~n13530 & n13585;
  assign n13588 = n3641 & n12668;
  assign n13589 = n3740 & n12665;
  assign n13590 = n12812 & ~n12814;
  assign n13591 = ~n12815 & ~n13590;
  assign n13592 = n556 & n13591;
  assign n13593 = n3961 & n12662;
  assign n13594 = ~n13592 & ~n13593;
  assign n13595 = ~n13589 & n13594;
  assign n13596 = ~n13588 & n13595;
  assign n13597 = ~n13587 & ~n13596;
  assign n13598 = ~n13586 & ~n13597;
  assign n13599 = n13528 & ~n13598;
  assign n13600 = ~n13528 & n13598;
  assign n13601 = ~n13599 & ~n13600;
  assign n13602 = n4006 & n12656;
  assign n13603 = n4133 & n12653;
  assign n13604 = n4002 & n12991;
  assign n13605 = n4555 & n12650;
  assign n13606 = ~n13604 & ~n13605;
  assign n13607 = ~n13603 & n13606;
  assign n13608 = ~n13602 & n13607;
  assign n13609 = pi29  & n13608;
  assign n13610 = ~pi29  & ~n13608;
  assign n13611 = ~n13609 & ~n13610;
  assign n13612 = n13601 & ~n13611;
  assign n13613 = ~n13599 & ~n13612;
  assign n13614 = n13255 & n13265;
  assign n13615 = ~n13266 & ~n13614;
  assign n13616 = ~n13613 & n13615;
  assign n13617 = n13613 & ~n13615;
  assign n13618 = n4601 & n12644;
  assign n13619 = n4783 & n12639;
  assign n13620 = n4602 & n13210;
  assign n13621 = n4801 & n12636;
  assign n13622 = ~n13620 & ~n13621;
  assign n13623 = ~n13619 & n13622;
  assign n13624 = ~n13618 & n13623;
  assign n13625 = pi26  & n13624;
  assign n13626 = ~pi26  & ~n13624;
  assign n13627 = ~n13625 & ~n13626;
  assign n13628 = ~n13617 & ~n13627;
  assign n13629 = ~n13616 & ~n13628;
  assign n13630 = ~n13526 & ~n13629;
  assign n13631 = ~n13523 & ~n13630;
  assign n13632 = ~n13287 & ~n13288;
  assign n13633 = ~n13300 & n13632;
  assign n13634 = n13300 & ~n13632;
  assign n13635 = ~n13633 & ~n13634;
  assign n13636 = ~n13631 & n13635;
  assign n13637 = n13631 & ~n13635;
  assign n13638 = n5238 & n12625;
  assign n13639 = n71 & n12622;
  assign n13640 = n5239 & n13463;
  assign n13641 = n5326 & n12614;
  assign n13642 = ~n13640 & ~n13641;
  assign n13643 = ~n13639 & n13642;
  assign n13644 = ~n13638 & n13643;
  assign n13645 = pi23  & n13644;
  assign n13646 = ~pi23  & ~n13644;
  assign n13647 = ~n13645 & ~n13646;
  assign n13648 = ~n13637 & ~n13647;
  assign n13649 = ~n13636 & ~n13648;
  assign n13650 = ~n13508 & ~n13649;
  assign n13651 = n13508 & n13649;
  assign n13652 = ~n13303 & ~n13304;
  assign n13653 = ~n13318 & n13652;
  assign n13654 = n13318 & ~n13652;
  assign n13655 = ~n13653 & ~n13654;
  assign n13656 = ~n13651 & n13655;
  assign n13657 = ~n13650 & ~n13656;
  assign n13658 = n13498 & ~n13657;
  assign n13659 = ~n13650 & ~n13651;
  assign n13660 = n13655 & n13659;
  assign n13661 = ~n13655 & ~n13659;
  assign n13662 = ~n13660 & ~n13661;
  assign n13663 = n13526 & n13629;
  assign n13664 = ~n13630 & ~n13663;
  assign n13665 = n5238 & n12630;
  assign n13666 = n71 & n12625;
  assign n13667 = n5239 & n13325;
  assign n13668 = n5326 & n12622;
  assign n13669 = ~n13667 & ~n13668;
  assign n13670 = ~n13666 & n13669;
  assign n13671 = ~n13665 & n13670;
  assign n13672 = pi23  & n13671;
  assign n13673 = ~pi23  & ~n13671;
  assign n13674 = ~n13672 & ~n13673;
  assign n13675 = n13664 & ~n13674;
  assign n13676 = n13664 & n13674;
  assign n13677 = ~n13664 & ~n13674;
  assign n13678 = ~n13676 & ~n13677;
  assign n13679 = ~n13616 & ~n13617;
  assign n13680 = ~n13627 & n13679;
  assign n13681 = n13627 & ~n13679;
  assign n13682 = ~n13680 & ~n13681;
  assign n13683 = n4006 & n12659;
  assign n13684 = n4133 & n12656;
  assign n13685 = n4002 & n13059;
  assign n13686 = n4555 & n12653;
  assign n13687 = ~n13685 & ~n13686;
  assign n13688 = ~n13684 & n13687;
  assign n13689 = ~n13683 & n13688;
  assign n13690 = pi29  & n13689;
  assign n13691 = ~pi29  & ~n13689;
  assign n13692 = ~n13690 & ~n13691;
  assign n13693 = ~n13586 & ~n13587;
  assign n13694 = ~n13596 & n13693;
  assign n13695 = n13596 & ~n13693;
  assign n13696 = ~n13694 & ~n13695;
  assign n13697 = ~n13692 & n13696;
  assign n13698 = ~n320 & n5104;
  assign n13699 = ~n165 & n13698;
  assign n13700 = ~n626 & ~n681;
  assign n13701 = ~n545 & n13700;
  assign n13702 = ~n204 & n2418;
  assign n13703 = ~n293 & n13702;
  assign n13704 = n13701 & n13703;
  assign n13705 = ~n349 & n13704;
  assign n13706 = ~n308 & n2082;
  assign n13707 = ~n231 & n13706;
  assign n13708 = n725 & n13707;
  assign n13709 = n13705 & n13708;
  assign n13710 = n1169 & n13709;
  assign n13711 = n257 & n13710;
  assign n13712 = n2768 & n4918;
  assign n13713 = n148 & n13712;
  assign n13714 = ~n701 & n13713;
  assign n13715 = n13711 & n13714;
  assign n13716 = n6675 & n13715;
  assign n13717 = ~n239 & n13716;
  assign n13718 = ~n357 & ~n384;
  assign n13719 = ~n307 & n13718;
  assign n13720 = ~n698 & n3715;
  assign n13721 = ~n475 & n13720;
  assign n13722 = n13719 & n13721;
  assign n13723 = n3429 & n13722;
  assign n13724 = n306 & n13723;
  assign n13725 = n3700 & n13724;
  assign n13726 = ~n181 & n13725;
  assign n13727 = n13717 & n13726;
  assign n13728 = ~n187 & n13727;
  assign n13729 = n13699 & n13728;
  assign n13730 = ~n363 & n5105;
  assign n13731 = n1361 & n6371;
  assign n13732 = n985 & n13731;
  assign n13733 = n1767 & n13732;
  assign n13734 = n1141 & n13733;
  assign n13735 = ~n232 & n13734;
  assign n13736 = n861 & n3085;
  assign n13737 = n253 & n13736;
  assign n13738 = ~n203 & n1925;
  assign n13739 = ~n455 & n2979;
  assign n13740 = ~n149 & n13739;
  assign n13741 = n13738 & n13740;
  assign n13742 = n3242 & n13741;
  assign n13743 = n13737 & n13742;
  assign n13744 = n1922 & n13743;
  assign n13745 = ~n581 & n13744;
  assign n13746 = n13735 & n13745;
  assign n13747 = ~n424 & n13746;
  assign n13748 = n13730 & n13747;
  assign n13749 = ~n13729 & ~n13748;
  assign n13750 = n7647 & n7653;
  assign n13751 = ~n12608 & ~n13750;
  assign n13752 = pi11  & ~n13751;
  assign n13753 = ~pi11  & n13751;
  assign n13754 = ~n13752 & ~n13753;
  assign n13755 = n13729 & n13748;
  assign n13756 = ~n13749 & ~n13755;
  assign n13757 = n13754 & n13756;
  assign n13758 = ~n13749 & ~n13757;
  assign n13759 = n13149 & ~n13758;
  assign n13760 = ~n13149 & n13758;
  assign n13761 = ~n13759 & ~n13760;
  assign n13762 = n3641 & n12674;
  assign n13763 = n12804 & ~n12806;
  assign n13764 = ~n12807 & ~n13763;
  assign n13765 = n556 & n13764;
  assign n13766 = n3961 & n12668;
  assign n13767 = n3740 & n12671;
  assign n13768 = ~n13766 & ~n13767;
  assign n13769 = ~n13765 & n13768;
  assign n13770 = ~n13762 & n13769;
  assign n13771 = n13761 & ~n13770;
  assign n13772 = ~n13759 & ~n13771;
  assign n13773 = ~n13573 & ~n13574;
  assign n13774 = ~n13583 & n13773;
  assign n13775 = n13583 & ~n13773;
  assign n13776 = ~n13774 & ~n13775;
  assign n13777 = ~n13772 & n13776;
  assign n13778 = n13772 & ~n13776;
  assign n13779 = ~n13777 & ~n13778;
  assign n13780 = ~n13754 & ~n13756;
  assign n13781 = ~n13757 & ~n13780;
  assign n13782 = n3641 & n12677;
  assign n13783 = n3740 & n12674;
  assign n13784 = n12800 & ~n12802;
  assign n13785 = ~n12803 & ~n13784;
  assign n13786 = n556 & n13785;
  assign n13787 = n3961 & n12671;
  assign n13788 = ~n13786 & ~n13787;
  assign n13789 = ~n13783 & n13788;
  assign n13790 = ~n13782 & n13789;
  assign n13791 = n13781 & ~n13790;
  assign n13792 = n13781 & n13790;
  assign n13793 = ~n13781 & ~n13790;
  assign n13794 = ~n13792 & ~n13793;
  assign n13795 = n355 & n2411;
  assign n13796 = n989 & n13795;
  assign n13797 = n1058 & n13796;
  assign n13798 = n558 & n13797;
  assign n13799 = ~n463 & n13798;
  assign n13800 = n300 & n4992;
  assign n13801 = ~n117 & n13800;
  assign n13802 = ~n683 & n13801;
  assign n13803 = n13799 & n13802;
  assign n13804 = ~n455 & n1186;
  assign n13805 = n1070 & n2708;
  assign n13806 = n1079 & n13805;
  assign n13807 = ~n315 & n1482;
  assign n13808 = ~n435 & n13807;
  assign n13809 = ~n536 & n13808;
  assign n13810 = n1025 & n13809;
  assign n13811 = n2195 & n13810;
  assign n13812 = n392 & n13811;
  assign n13813 = n13806 & n13812;
  assign n13814 = ~n698 & n13813;
  assign n13815 = n2218 & n3267;
  assign n13816 = ~n88 & n13815;
  assign n13817 = ~n289 & ~n474;
  assign n13818 = ~n414 & n13817;
  assign n13819 = ~n668 & n13818;
  assign n13820 = n596 & n13819;
  assign n13821 = ~n464 & n13820;
  assign n13822 = ~n639 & n13821;
  assign n13823 = n13816 & n13822;
  assign n13824 = n13814 & n13823;
  assign n13825 = n13804 & n13824;
  assign n13826 = n706 & n13825;
  assign n13827 = ~n186 & n13826;
  assign n13828 = ~n280 & n3168;
  assign n13829 = n415 & n13828;
  assign n13830 = ~n278 & ~n344;
  assign n13831 = ~n614 & n2904;
  assign n13832 = ~n216 & n13831;
  assign n13833 = n13830 & n13832;
  assign n13834 = n2032 & n13833;
  assign n13835 = n13829 & n13834;
  assign n13836 = n1587 & n13835;
  assign n13837 = ~n307 & n13836;
  assign n13838 = ~n85 & n13837;
  assign n13839 = n13827 & n13838;
  assign n13840 = n13803 & n13839;
  assign n13841 = n13729 & ~n13840;
  assign n13842 = ~n455 & n2056;
  assign n13843 = n196 & ~n330;
  assign n13844 = ~n668 & n1138;
  assign n13845 = n13843 & n13844;
  assign n13846 = ~n216 & n13845;
  assign n13847 = ~n277 & n528;
  assign n13848 = ~n430 & n13847;
  assign n13849 = ~n308 & n13848;
  assign n13850 = ~n261 & n13849;
  assign n13851 = n13846 & n13850;
  assign n13852 = n4385 & n13851;
  assign n13853 = n1332 & n2760;
  assign n13854 = n3029 & n13853;
  assign n13855 = n1174 & n13854;
  assign n13856 = n476 & n13855;
  assign n13857 = n13852 & n13856;
  assign n13858 = ~n186 & n1343;
  assign n13859 = n2115 & n2997;
  assign n13860 = n1513 & n13859;
  assign n13861 = ~n350 & n13860;
  assign n13862 = n1447 & n4898;
  assign n13863 = ~n594 & n13862;
  assign n13864 = ~n150 & n13863;
  assign n13865 = n13861 & n13864;
  assign n13866 = ~n304 & n13865;
  assign n13867 = n13858 & n13866;
  assign n13868 = n13857 & n13867;
  assign n13869 = ~n154 & n584;
  assign n13870 = ~n413 & n13869;
  assign n13871 = ~n436 & n13870;
  assign n13872 = ~n188 & n12957;
  assign n13873 = ~n294 & n1976;
  assign n13874 = ~n315 & n13873;
  assign n13875 = n13872 & n13874;
  assign n13876 = n1369 & n13875;
  assign n13877 = n13871 & n13876;
  assign n13878 = n758 & n13877;
  assign n13879 = n3159 & n13878;
  assign n13880 = n706 & n13879;
  assign n13881 = ~n611 & n13880;
  assign n13882 = n13868 & n13881;
  assign n13883 = ~n299 & n13882;
  assign n13884 = n13842 & n13883;
  assign n13885 = n2491 & n5672;
  assign n13886 = n1998 & n13885;
  assign n13887 = n884 & n3944;
  assign n13888 = n1388 & n13887;
  assign n13889 = n13886 & n13888;
  assign n13890 = ~n330 & ~n538;
  assign n13891 = ~n154 & n13890;
  assign n13892 = ~n342 & n13891;
  assign n13893 = ~n236 & n13892;
  assign n13894 = ~n88 & ~n685;
  assign n13895 = n13893 & n13894;
  assign n13896 = n13889 & n13895;
  assign n13897 = ~n173 & n13896;
  assign n13898 = ~n504 & n2504;
  assign n13899 = ~n181 & n13898;
  assign n13900 = ~n548 & n2418;
  assign n13901 = ~n576 & n2784;
  assign n13902 = n13900 & n13901;
  assign n13903 = n954 & n13902;
  assign n13904 = n13899 & n13903;
  assign n13905 = n1534 & n13904;
  assign n13906 = n2644 & n13905;
  assign n13907 = ~n629 & n13906;
  assign n13908 = ~n639 & n13907;
  assign n13909 = n13897 & n13908;
  assign n13910 = ~n232 & n13909;
  assign n13911 = ~n255 & n1192;
  assign n13912 = ~n505 & n13911;
  assign n13913 = n13910 & n13912;
  assign n13914 = ~n13884 & ~n13913;
  assign n13915 = n8467 & n8473;
  assign n13916 = ~n12608 & ~n13915;
  assign n13917 = pi8  & ~n13916;
  assign n13918 = ~pi8  & n13916;
  assign n13919 = ~n13917 & ~n13918;
  assign n13920 = n13884 & n13913;
  assign n13921 = ~n13914 & ~n13920;
  assign n13922 = n13919 & n13921;
  assign n13923 = ~n13914 & ~n13922;
  assign n13924 = n13729 & ~n13923;
  assign n13925 = ~n13729 & n13923;
  assign n13926 = ~n13924 & ~n13925;
  assign n13927 = n3641 & n12683;
  assign n13928 = n12792 & ~n12794;
  assign n13929 = ~n12795 & ~n13928;
  assign n13930 = n556 & n13929;
  assign n13931 = n3961 & n12677;
  assign n13932 = n3740 & n12680;
  assign n13933 = ~n13931 & ~n13932;
  assign n13934 = ~n13930 & n13933;
  assign n13935 = ~n13927 & n13934;
  assign n13936 = n13926 & ~n13935;
  assign n13937 = ~n13924 & ~n13936;
  assign n13938 = ~n13729 & n13840;
  assign n13939 = ~n13841 & ~n13938;
  assign n13940 = ~n13937 & n13939;
  assign n13941 = ~n13841 & ~n13940;
  assign n13942 = ~n13794 & ~n13941;
  assign n13943 = ~n13791 & ~n13942;
  assign n13944 = ~n13761 & n13770;
  assign n13945 = ~n13771 & ~n13944;
  assign n13946 = ~n13943 & n13945;
  assign n13947 = n13943 & ~n13945;
  assign n13948 = ~n13946 & ~n13947;
  assign n13949 = n4006 & n12665;
  assign n13950 = n4133 & n12662;
  assign n13951 = n4002 & n13165;
  assign n13952 = n4555 & n12659;
  assign n13953 = ~n13951 & ~n13952;
  assign n13954 = ~n13950 & n13953;
  assign n13955 = ~n13949 & n13954;
  assign n13956 = pi29  & n13955;
  assign n13957 = ~pi29  & ~n13955;
  assign n13958 = ~n13956 & ~n13957;
  assign n13959 = n13948 & ~n13958;
  assign n13960 = ~n13946 & ~n13959;
  assign n13961 = n13779 & ~n13960;
  assign n13962 = ~n13777 & ~n13961;
  assign n13963 = n13692 & ~n13696;
  assign n13964 = ~n13697 & ~n13963;
  assign n13965 = ~n13962 & n13964;
  assign n13966 = ~n13697 & ~n13965;
  assign n13967 = ~n13601 & n13611;
  assign n13968 = ~n13612 & ~n13967;
  assign n13969 = ~n13966 & n13968;
  assign n13970 = n13966 & ~n13968;
  assign n13971 = n4601 & n12647;
  assign n13972 = n4783 & n12644;
  assign n13973 = n4602 & ~n13193;
  assign n13974 = n4801 & n12639;
  assign n13975 = ~n13973 & ~n13974;
  assign n13976 = ~n13972 & n13975;
  assign n13977 = ~n13971 & n13976;
  assign n13978 = pi26  & n13977;
  assign n13979 = ~pi26  & ~n13977;
  assign n13980 = ~n13978 & ~n13979;
  assign n13981 = ~n13970 & ~n13980;
  assign n13982 = ~n13969 & ~n13981;
  assign n13983 = n13682 & ~n13982;
  assign n13984 = ~n13682 & n13982;
  assign n13985 = n5238 & n12633;
  assign n13986 = n71 & n12630;
  assign n13987 = n5239 & ~n13227;
  assign n13988 = n5326 & n12625;
  assign n13989 = ~n13987 & ~n13988;
  assign n13990 = ~n13986 & n13989;
  assign n13991 = ~n13985 & n13990;
  assign n13992 = pi23  & n13991;
  assign n13993 = ~pi23  & ~n13991;
  assign n13994 = ~n13992 & ~n13993;
  assign n13995 = ~n13984 & ~n13994;
  assign n13996 = ~n13983 & ~n13995;
  assign n13997 = ~n13678 & ~n13996;
  assign n13998 = ~n13675 & ~n13997;
  assign n13999 = ~n13636 & ~n13637;
  assign n14000 = ~n13647 & n13999;
  assign n14001 = n13647 & ~n13999;
  assign n14002 = ~n14000 & ~n14001;
  assign n14003 = ~n13998 & n14002;
  assign n14004 = n13998 & ~n14002;
  assign n14005 = n5435 & n12606;
  assign n14006 = n6055 & n12616;
  assign n14007 = n5429 & ~n13483;
  assign n14008 = n6071 & ~n12608;
  assign n14009 = ~n14007 & ~n14008;
  assign n14010 = ~n14006 & n14009;
  assign n14011 = ~n14005 & n14010;
  assign n14012 = pi20  & n14011;
  assign n14013 = ~pi20  & ~n14011;
  assign n14014 = ~n14012 & ~n14013;
  assign n14015 = ~n14004 & ~n14014;
  assign n14016 = ~n14003 & ~n14015;
  assign n14017 = n13662 & ~n14016;
  assign n14018 = ~n13662 & n14016;
  assign n14019 = ~n14017 & ~n14018;
  assign n14020 = n6055 & n12606;
  assign n14021 = ~n12611 & n14008;
  assign n14022 = n5435 & n12614;
  assign n14023 = n5429 & n12868;
  assign n14024 = ~n14022 & ~n14023;
  assign n14025 = ~n14021 & n14024;
  assign n14026 = ~n14020 & n14025;
  assign n14027 = pi20  & n14026;
  assign n14028 = ~pi20  & ~n14026;
  assign n14029 = ~n14027 & ~n14028;
  assign n14030 = ~n13983 & ~n13984;
  assign n14031 = ~n13994 & n14030;
  assign n14032 = n13994 & ~n14030;
  assign n14033 = ~n14031 & ~n14032;
  assign n14034 = n13962 & ~n13964;
  assign n14035 = ~n13965 & ~n14034;
  assign n14036 = n4601 & n12650;
  assign n14037 = n4783 & n12647;
  assign n14038 = n4602 & n13275;
  assign n14039 = n4801 & n12644;
  assign n14040 = ~n14038 & ~n14039;
  assign n14041 = ~n14037 & n14040;
  assign n14042 = ~n14036 & n14041;
  assign n14043 = pi26  & n14042;
  assign n14044 = ~pi26  & ~n14042;
  assign n14045 = ~n14043 & ~n14044;
  assign n14046 = n14035 & ~n14045;
  assign n14047 = n14035 & n14045;
  assign n14048 = ~n14035 & ~n14045;
  assign n14049 = ~n14047 & ~n14048;
  assign n14050 = ~n13779 & n13960;
  assign n14051 = ~n13961 & ~n14050;
  assign n14052 = n4006 & n12662;
  assign n14053 = n4133 & n12659;
  assign n14054 = n4002 & n13246;
  assign n14055 = n4555 & n12656;
  assign n14056 = ~n14054 & ~n14055;
  assign n14057 = ~n14053 & n14056;
  assign n14058 = ~n14052 & n14057;
  assign n14059 = pi29  & n14058;
  assign n14060 = ~pi29  & ~n14058;
  assign n14061 = ~n14059 & ~n14060;
  assign n14062 = n14051 & ~n14061;
  assign n14063 = n14051 & n14061;
  assign n14064 = ~n14051 & ~n14061;
  assign n14065 = ~n14063 & ~n14064;
  assign n14066 = n4601 & n12653;
  assign n14067 = n4783 & n12650;
  assign n14068 = n4602 & n13042;
  assign n14069 = n4801 & n12647;
  assign n14070 = ~n14068 & ~n14069;
  assign n14071 = ~n14067 & n14070;
  assign n14072 = ~n14066 & n14071;
  assign n14073 = pi26  & n14072;
  assign n14074 = ~pi26  & ~n14072;
  assign n14075 = ~n14073 & ~n14074;
  assign n14076 = ~n14065 & ~n14075;
  assign n14077 = ~n14062 & ~n14076;
  assign n14078 = ~n14049 & ~n14077;
  assign n14079 = ~n14046 & ~n14078;
  assign n14080 = ~n13969 & ~n13970;
  assign n14081 = ~n13980 & n14080;
  assign n14082 = n13980 & ~n14080;
  assign n14083 = ~n14081 & ~n14082;
  assign n14084 = ~n14079 & n14083;
  assign n14085 = n14079 & ~n14083;
  assign n14086 = n5238 & n12636;
  assign n14087 = n71 & n12633;
  assign n14088 = n5239 & n13292;
  assign n14089 = n5326 & n12630;
  assign n14090 = ~n14088 & ~n14089;
  assign n14091 = ~n14087 & n14090;
  assign n14092 = ~n14086 & n14091;
  assign n14093 = pi23  & n14092;
  assign n14094 = ~pi23  & ~n14092;
  assign n14095 = ~n14093 & ~n14094;
  assign n14096 = ~n14085 & ~n14095;
  assign n14097 = ~n14084 & ~n14096;
  assign n14098 = n14033 & ~n14097;
  assign n14099 = ~n14033 & n14097;
  assign n14100 = n5435 & n12622;
  assign n14101 = n6055 & n12614;
  assign n14102 = n5429 & ~n13310;
  assign n14103 = n6071 & n12606;
  assign n14104 = ~n14102 & ~n14103;
  assign n14105 = ~n14101 & n14104;
  assign n14106 = ~n14100 & n14105;
  assign n14107 = pi20  & n14106;
  assign n14108 = ~pi20  & ~n14106;
  assign n14109 = ~n14107 & ~n14108;
  assign n14110 = ~n14099 & ~n14109;
  assign n14111 = ~n14098 & ~n14110;
  assign n14112 = ~n14029 & ~n14111;
  assign n14113 = n13678 & n13996;
  assign n14114 = ~n13997 & ~n14113;
  assign n14115 = n14029 & ~n14111;
  assign n14116 = ~n14029 & n14111;
  assign n14117 = ~n14115 & ~n14116;
  assign n14118 = n14114 & ~n14117;
  assign n14119 = ~n14112 & ~n14118;
  assign n14120 = ~n14003 & ~n14004;
  assign n14121 = ~n14014 & n14120;
  assign n14122 = n14014 & ~n14120;
  assign n14123 = ~n14121 & ~n14122;
  assign n14124 = ~n14119 & n14123;
  assign n14125 = n14119 & n14123;
  assign n14126 = ~n14119 & ~n14123;
  assign n14127 = ~n14125 & ~n14126;
  assign n14128 = ~n14114 & n14117;
  assign n14129 = ~n14118 & ~n14128;
  assign n14130 = n6185 & ~n13499;
  assign n14131 = n6184 & ~n12611;
  assign n14132 = ~n6527 & ~n6543;
  assign n14133 = ~n14131 & n14132;
  assign n14134 = ~n12608 & ~n14133;
  assign n14135 = ~n14130 & ~n14134;
  assign n14136 = pi17  & n14135;
  assign n14137 = ~pi17  & ~n14135;
  assign n14138 = ~n14136 & ~n14137;
  assign n14139 = n14049 & n14077;
  assign n14140 = ~n14078 & ~n14139;
  assign n14141 = n5238 & n12639;
  assign n14142 = n71 & n12636;
  assign n14143 = n5239 & n13396;
  assign n14144 = n5326 & n12633;
  assign n14145 = ~n14143 & ~n14144;
  assign n14146 = ~n14142 & n14145;
  assign n14147 = ~n14141 & n14146;
  assign n14148 = pi23  & n14147;
  assign n14149 = ~pi23  & ~n14147;
  assign n14150 = ~n14148 & ~n14149;
  assign n14151 = n14140 & ~n14150;
  assign n14152 = n14140 & n14150;
  assign n14153 = ~n14140 & ~n14150;
  assign n14154 = ~n14152 & ~n14153;
  assign n14155 = n14065 & n14075;
  assign n14156 = ~n14076 & ~n14155;
  assign n14157 = ~n13948 & n13958;
  assign n14158 = ~n13959 & ~n14157;
  assign n14159 = n13937 & ~n13939;
  assign n14160 = ~n13940 & ~n14159;
  assign n14161 = n3641 & n12680;
  assign n14162 = n3740 & n12677;
  assign n14163 = n12796 & ~n12798;
  assign n14164 = ~n12799 & ~n14163;
  assign n14165 = n556 & n14164;
  assign n14166 = n3961 & n12674;
  assign n14167 = ~n14165 & ~n14166;
  assign n14168 = ~n14162 & n14167;
  assign n14169 = ~n14161 & n14168;
  assign n14170 = n14160 & ~n14169;
  assign n14171 = n14160 & n14169;
  assign n14172 = ~n14160 & ~n14169;
  assign n14173 = ~n14171 & ~n14172;
  assign n14174 = n4006 & n12671;
  assign n14175 = n4133 & n12668;
  assign n14176 = n4002 & n13578;
  assign n14177 = n4555 & n12665;
  assign n14178 = ~n14176 & ~n14177;
  assign n14179 = ~n14175 & n14178;
  assign n14180 = ~n14174 & n14179;
  assign n14181 = pi29  & n14180;
  assign n14182 = ~pi29  & ~n14180;
  assign n14183 = ~n14181 & ~n14182;
  assign n14184 = ~n14173 & ~n14183;
  assign n14185 = ~n14170 & ~n14184;
  assign n14186 = ~n13794 & n13941;
  assign n14187 = n13794 & ~n13941;
  assign n14188 = ~n14186 & ~n14187;
  assign n14189 = ~n14185 & ~n14188;
  assign n14190 = n4006 & n12668;
  assign n14191 = n4133 & n12665;
  assign n14192 = n4002 & n13591;
  assign n14193 = n4555 & n12662;
  assign n14194 = ~n14192 & ~n14193;
  assign n14195 = ~n14191 & n14194;
  assign n14196 = ~n14190 & n14195;
  assign n14197 = pi29  & n14196;
  assign n14198 = ~pi29  & ~n14196;
  assign n14199 = ~n14197 & ~n14198;
  assign n14200 = n14185 & n14188;
  assign n14201 = ~n14199 & ~n14200;
  assign n14202 = ~n14189 & ~n14201;
  assign n14203 = n14158 & ~n14202;
  assign n14204 = ~n14158 & n14202;
  assign n14205 = n4601 & n12656;
  assign n14206 = n4783 & n12653;
  assign n14207 = n4602 & n12991;
  assign n14208 = n4801 & n12650;
  assign n14209 = ~n14207 & ~n14208;
  assign n14210 = ~n14206 & n14209;
  assign n14211 = ~n14205 & n14210;
  assign n14212 = pi26  & n14211;
  assign n14213 = ~pi26  & ~n14211;
  assign n14214 = ~n14212 & ~n14213;
  assign n14215 = ~n14204 & ~n14214;
  assign n14216 = ~n14203 & ~n14215;
  assign n14217 = n14156 & ~n14216;
  assign n14218 = ~n14156 & n14216;
  assign n14219 = n5238 & n12644;
  assign n14220 = n71 & n12639;
  assign n14221 = n5239 & n13210;
  assign n14222 = n5326 & n12636;
  assign n14223 = ~n14221 & ~n14222;
  assign n14224 = ~n14220 & n14223;
  assign n14225 = ~n14219 & n14224;
  assign n14226 = pi23  & n14225;
  assign n14227 = ~pi23  & ~n14225;
  assign n14228 = ~n14226 & ~n14227;
  assign n14229 = ~n14218 & ~n14228;
  assign n14230 = ~n14217 & ~n14229;
  assign n14231 = ~n14154 & ~n14230;
  assign n14232 = ~n14151 & ~n14231;
  assign n14233 = ~n14084 & ~n14085;
  assign n14234 = ~n14095 & n14233;
  assign n14235 = n14095 & ~n14233;
  assign n14236 = ~n14234 & ~n14235;
  assign n14237 = ~n14232 & n14236;
  assign n14238 = n14232 & ~n14236;
  assign n14239 = n5435 & n12625;
  assign n14240 = n6055 & n12622;
  assign n14241 = n5429 & n13463;
  assign n14242 = n6071 & n12614;
  assign n14243 = ~n14241 & ~n14242;
  assign n14244 = ~n14240 & n14243;
  assign n14245 = ~n14239 & n14244;
  assign n14246 = pi20  & n14245;
  assign n14247 = ~pi20  & ~n14245;
  assign n14248 = ~n14246 & ~n14247;
  assign n14249 = ~n14238 & ~n14248;
  assign n14250 = ~n14237 & ~n14249;
  assign n14251 = ~n14138 & ~n14250;
  assign n14252 = n14138 & n14250;
  assign n14253 = ~n14098 & ~n14099;
  assign n14254 = ~n14109 & n14253;
  assign n14255 = n14109 & ~n14253;
  assign n14256 = ~n14254 & ~n14255;
  assign n14257 = ~n14252 & n14256;
  assign n14258 = ~n14251 & ~n14257;
  assign n14259 = n14129 & ~n14258;
  assign n14260 = ~n14251 & ~n14252;
  assign n14261 = n14256 & n14260;
  assign n14262 = ~n14256 & ~n14260;
  assign n14263 = ~n14261 & ~n14262;
  assign n14264 = n14154 & n14230;
  assign n14265 = ~n14231 & ~n14264;
  assign n14266 = n5435 & n12630;
  assign n14267 = n6055 & n12625;
  assign n14268 = n5429 & n13325;
  assign n14269 = n6071 & n12622;
  assign n14270 = ~n14268 & ~n14269;
  assign n14271 = ~n14267 & n14270;
  assign n14272 = ~n14266 & n14271;
  assign n14273 = pi20  & n14272;
  assign n14274 = ~pi20  & ~n14272;
  assign n14275 = ~n14273 & ~n14274;
  assign n14276 = n14265 & ~n14275;
  assign n14277 = n14265 & n14275;
  assign n14278 = ~n14265 & ~n14275;
  assign n14279 = ~n14277 & ~n14278;
  assign n14280 = ~n14217 & ~n14218;
  assign n14281 = ~n14228 & n14280;
  assign n14282 = n14228 & ~n14280;
  assign n14283 = ~n14281 & ~n14282;
  assign n14284 = n4601 & n12659;
  assign n14285 = n4783 & n12656;
  assign n14286 = n4602 & n13059;
  assign n14287 = n4801 & n12653;
  assign n14288 = ~n14286 & ~n14287;
  assign n14289 = ~n14285 & n14288;
  assign n14290 = ~n14284 & n14289;
  assign n14291 = pi26  & n14290;
  assign n14292 = ~pi26  & ~n14290;
  assign n14293 = ~n14291 & ~n14292;
  assign n14294 = ~n14189 & ~n14200;
  assign n14295 = n14199 & ~n14294;
  assign n14296 = ~n14199 & n14294;
  assign n14297 = ~n14295 & ~n14296;
  assign n14298 = ~n14293 & n14297;
  assign n14299 = n14293 & n14297;
  assign n14300 = ~n14293 & ~n14297;
  assign n14301 = ~n14299 & ~n14300;
  assign n14302 = ~n13926 & n13935;
  assign n14303 = ~n13936 & ~n14302;
  assign n14304 = n1924 & n13069;
  assign n14305 = n1344 & n14304;
  assign n14306 = n2713 & n14305;
  assign n14307 = n2611 & n14306;
  assign n14308 = ~n681 & n14307;
  assign n14309 = n1054 & n2842;
  assign n14310 = ~n685 & n14309;
  assign n14311 = ~n186 & n14310;
  assign n14312 = n14308 & n14311;
  assign n14313 = ~n701 & n14312;
  assign n14314 = n89 & n1101;
  assign n14315 = n167 & n5866;
  assign n14316 = n14314 & n14315;
  assign n14317 = ~n629 & n14316;
  assign n14318 = ~n236 & n14317;
  assign n14319 = n386 & n14318;
  assign n14320 = n14313 & n14319;
  assign n14321 = n13884 & ~n14320;
  assign n14322 = n1268 & n1976;
  assign n14323 = ~n401 & n14322;
  assign n14324 = ~n195 & n1023;
  assign n14325 = ~n261 & n14324;
  assign n14326 = n14323 & n14325;
  assign n14327 = ~n255 & n3896;
  assign n14328 = ~n581 & n14327;
  assign n14329 = n1494 & n2474;
  assign n14330 = ~n462 & n14329;
  assign n14331 = ~n344 & n14330;
  assign n14332 = n14328 & n14331;
  assign n14333 = n14326 & n14332;
  assign n14334 = n4073 & n14333;
  assign n14335 = ~n373 & n14334;
  assign n14336 = n2940 & n4469;
  assign n14337 = n13128 & n14336;
  assign n14338 = n107 & n14337;
  assign n14339 = n1419 & n3312;
  assign n14340 = n1409 & n14339;
  assign n14341 = n306 & n14340;
  assign n14342 = n14338 & n14341;
  assign n14343 = ~n632 & n1148;
  assign n14344 = ~n85 & n14343;
  assign n14345 = n13819 & n14344;
  assign n14346 = n14342 & n14345;
  assign n14347 = n14335 & n14346;
  assign n14348 = n2345 & n14347;
  assign n14349 = ~n254 & n14348;
  assign n14350 = n946 & n13709;
  assign n14351 = ~n683 & n14350;
  assign n14352 = n14349 & n14351;
  assign n14353 = n4267 & n6662;
  assign n14354 = ~n277 & n14353;
  assign n14355 = n1377 & n7187;
  assign n14356 = n4472 & n14355;
  assign n14357 = n4175 & n14356;
  assign n14358 = ~n290 & n14357;
  assign n14359 = n14354 & n14358;
  assign n14360 = n14352 & n14359;
  assign n14361 = n11286 & n11287;
  assign n14362 = ~pi2  & ~n14361;
  assign n14363 = ~n12608 & n14362;
  assign n14364 = pi2  & n12608;
  assign n14365 = ~n14363 & ~n14364;
  assign n14366 = ~n14360 & n14365;
  assign n14367 = n14360 & n14365;
  assign n14368 = ~n14360 & ~n14365;
  assign n14369 = ~n14367 & ~n14368;
  assign n14370 = n9718 & n9724;
  assign n14371 = ~n12608 & ~n14370;
  assign n14372 = ~pi5  & n14371;
  assign n14373 = pi5  & ~n14371;
  assign n14374 = ~n14372 & ~n14373;
  assign n14375 = ~n14369 & n14374;
  assign n14376 = ~n14366 & ~n14375;
  assign n14377 = n13884 & ~n14376;
  assign n14378 = ~n13884 & n14376;
  assign n14379 = ~n14377 & ~n14378;
  assign n14380 = n3641 & n12692;
  assign n14381 = n12780 & ~n12782;
  assign n14382 = ~n12783 & ~n14381;
  assign n14383 = n556 & n14382;
  assign n14384 = n3961 & n12686;
  assign n14385 = n3740 & n12689;
  assign n14386 = ~n14384 & ~n14385;
  assign n14387 = ~n14383 & n14386;
  assign n14388 = ~n14380 & n14387;
  assign n14389 = n14379 & ~n14388;
  assign n14390 = ~n14377 & ~n14389;
  assign n14391 = ~n13884 & n14320;
  assign n14392 = ~n14321 & ~n14391;
  assign n14393 = ~n14390 & n14392;
  assign n14394 = ~n14321 & ~n14393;
  assign n14395 = ~n13919 & ~n13921;
  assign n14396 = ~n13922 & ~n14395;
  assign n14397 = ~n14394 & n14396;
  assign n14398 = n14394 & ~n14396;
  assign n14399 = n3641 & n12686;
  assign n14400 = n3740 & n12683;
  assign n14401 = n12788 & ~n12790;
  assign n14402 = ~n12791 & ~n14401;
  assign n14403 = n556 & n14402;
  assign n14404 = n3961 & n12680;
  assign n14405 = ~n14403 & ~n14404;
  assign n14406 = ~n14400 & n14405;
  assign n14407 = ~n14399 & n14406;
  assign n14408 = ~n14398 & ~n14407;
  assign n14409 = ~n14397 & ~n14408;
  assign n14410 = n14303 & ~n14409;
  assign n14411 = ~n14303 & n14409;
  assign n14412 = ~n14410 & ~n14411;
  assign n14413 = n4006 & n12674;
  assign n14414 = n4133 & n12671;
  assign n14415 = n4002 & n13764;
  assign n14416 = n4555 & n12668;
  assign n14417 = ~n14415 & ~n14416;
  assign n14418 = ~n14414 & n14417;
  assign n14419 = ~n14413 & n14418;
  assign n14420 = pi29  & n14419;
  assign n14421 = ~pi29  & ~n14419;
  assign n14422 = ~n14420 & ~n14421;
  assign n14423 = n14412 & ~n14422;
  assign n14424 = ~n14410 & ~n14423;
  assign n14425 = n14173 & n14183;
  assign n14426 = ~n14184 & ~n14425;
  assign n14427 = ~n14424 & n14426;
  assign n14428 = n14424 & ~n14426;
  assign n14429 = n4601 & n12662;
  assign n14430 = n4783 & n12659;
  assign n14431 = n4602 & n13246;
  assign n14432 = n4801 & n12656;
  assign n14433 = ~n14431 & ~n14432;
  assign n14434 = ~n14430 & n14433;
  assign n14435 = ~n14429 & n14434;
  assign n14436 = pi26  & n14435;
  assign n14437 = ~pi26  & ~n14435;
  assign n14438 = ~n14436 & ~n14437;
  assign n14439 = ~n14428 & ~n14438;
  assign n14440 = ~n14427 & ~n14439;
  assign n14441 = ~n14301 & ~n14440;
  assign n14442 = ~n14298 & ~n14441;
  assign n14443 = ~n14203 & ~n14204;
  assign n14444 = ~n14214 & n14443;
  assign n14445 = n14214 & ~n14443;
  assign n14446 = ~n14444 & ~n14445;
  assign n14447 = ~n14442 & n14446;
  assign n14448 = n14442 & ~n14446;
  assign n14449 = n5238 & n12647;
  assign n14450 = n71 & n12644;
  assign n14451 = n5239 & ~n13193;
  assign n14452 = n5326 & n12639;
  assign n14453 = ~n14451 & ~n14452;
  assign n14454 = ~n14450 & n14453;
  assign n14455 = ~n14449 & n14454;
  assign n14456 = pi23  & n14455;
  assign n14457 = ~pi23  & ~n14455;
  assign n14458 = ~n14456 & ~n14457;
  assign n14459 = ~n14448 & ~n14458;
  assign n14460 = ~n14447 & ~n14459;
  assign n14461 = n14283 & ~n14460;
  assign n14462 = ~n14283 & n14460;
  assign n14463 = n5435 & n12633;
  assign n14464 = n6055 & n12630;
  assign n14465 = n5429 & ~n13227;
  assign n14466 = n6071 & n12625;
  assign n14467 = ~n14465 & ~n14466;
  assign n14468 = ~n14464 & n14467;
  assign n14469 = ~n14463 & n14468;
  assign n14470 = pi20  & n14469;
  assign n14471 = ~pi20  & ~n14469;
  assign n14472 = ~n14470 & ~n14471;
  assign n14473 = ~n14462 & ~n14472;
  assign n14474 = ~n14461 & ~n14473;
  assign n14475 = ~n14279 & ~n14474;
  assign n14476 = ~n14276 & ~n14475;
  assign n14477 = ~n14237 & ~n14238;
  assign n14478 = ~n14248 & n14477;
  assign n14479 = n14248 & ~n14477;
  assign n14480 = ~n14478 & ~n14479;
  assign n14481 = ~n14476 & n14480;
  assign n14482 = n14476 & ~n14480;
  assign n14483 = n6184 & n12606;
  assign n14484 = n6527 & n12616;
  assign n14485 = n6185 & ~n13483;
  assign n14486 = n6543 & ~n12608;
  assign n14487 = ~n14485 & ~n14486;
  assign n14488 = ~n14484 & n14487;
  assign n14489 = ~n14483 & n14488;
  assign n14490 = pi17  & n14489;
  assign n14491 = ~pi17  & ~n14489;
  assign n14492 = ~n14490 & ~n14491;
  assign n14493 = ~n14482 & ~n14492;
  assign n14494 = ~n14481 & ~n14493;
  assign n14495 = n14263 & ~n14494;
  assign n14496 = ~n14263 & n14494;
  assign n14497 = ~n14495 & ~n14496;
  assign n14498 = n6527 & n12606;
  assign n14499 = ~n12611 & n14486;
  assign n14500 = n6184 & n12614;
  assign n14501 = n6185 & n12868;
  assign n14502 = ~n14500 & ~n14501;
  assign n14503 = ~n14499 & n14502;
  assign n14504 = ~n14498 & n14503;
  assign n14505 = pi17  & n14504;
  assign n14506 = ~pi17  & ~n14504;
  assign n14507 = ~n14505 & ~n14506;
  assign n14508 = ~n14461 & ~n14462;
  assign n14509 = ~n14472 & n14508;
  assign n14510 = n14472 & ~n14508;
  assign n14511 = ~n14509 & ~n14510;
  assign n14512 = n14301 & n14440;
  assign n14513 = ~n14441 & ~n14512;
  assign n14514 = n5238 & n12650;
  assign n14515 = n71 & n12647;
  assign n14516 = n5239 & n13275;
  assign n14517 = n5326 & n12644;
  assign n14518 = ~n14516 & ~n14517;
  assign n14519 = ~n14515 & n14518;
  assign n14520 = ~n14514 & n14519;
  assign n14521 = pi23  & n14520;
  assign n14522 = ~pi23  & ~n14520;
  assign n14523 = ~n14521 & ~n14522;
  assign n14524 = n14513 & ~n14523;
  assign n14525 = n14513 & n14523;
  assign n14526 = ~n14513 & ~n14523;
  assign n14527 = ~n14525 & ~n14526;
  assign n14528 = ~n14427 & ~n14428;
  assign n14529 = ~n14438 & n14528;
  assign n14530 = n14438 & ~n14528;
  assign n14531 = ~n14529 & ~n14530;
  assign n14532 = n4006 & n12677;
  assign n14533 = n4133 & n12674;
  assign n14534 = n4002 & n13785;
  assign n14535 = n4555 & n12671;
  assign n14536 = ~n14534 & ~n14535;
  assign n14537 = ~n14533 & n14536;
  assign n14538 = ~n14532 & n14537;
  assign n14539 = pi29  & n14538;
  assign n14540 = ~pi29  & ~n14538;
  assign n14541 = ~n14539 & ~n14540;
  assign n14542 = ~n14397 & ~n14398;
  assign n14543 = ~n14407 & n14542;
  assign n14544 = n14407 & ~n14542;
  assign n14545 = ~n14543 & ~n14544;
  assign n14546 = ~n14541 & n14545;
  assign n14547 = n14390 & ~n14392;
  assign n14548 = ~n14393 & ~n14547;
  assign n14549 = n3641 & n12689;
  assign n14550 = n3740 & n12686;
  assign n14551 = n12784 & ~n12786;
  assign n14552 = ~n12787 & ~n14551;
  assign n14553 = n556 & n14552;
  assign n14554 = n3961 & n12683;
  assign n14555 = ~n14553 & ~n14554;
  assign n14556 = ~n14550 & n14555;
  assign n14557 = ~n14549 & n14556;
  assign n14558 = n14548 & ~n14557;
  assign n14559 = n14548 & n14557;
  assign n14560 = ~n14548 & ~n14557;
  assign n14561 = ~n14559 & ~n14560;
  assign n14562 = n2010 & n3375;
  assign n14563 = ~n289 & n14562;
  assign n14564 = ~n183 & n14563;
  assign n14565 = n871 & n3030;
  assign n14566 = n2642 & n14565;
  assign n14567 = ~n246 & n14566;
  assign n14568 = ~n382 & n14567;
  assign n14569 = ~n149 & n14568;
  assign n14570 = n14564 & n14569;
  assign n14571 = n2056 & n4212;
  assign n14572 = ~n349 & n14571;
  assign n14573 = ~n394 & n14572;
  assign n14574 = ~n293 & n3864;
  assign n14575 = ~n391 & n14574;
  assign n14576 = ~n638 & n14575;
  assign n14577 = n14573 & n14576;
  assign n14578 = n14570 & n14577;
  assign n14579 = ~n14365 & ~n14578;
  assign n14580 = n1454 & n2529;
  assign n14581 = n1464 & n14580;
  assign n14582 = n4888 & n14581;
  assign n14583 = ~n457 & n14582;
  assign n14584 = n1272 & n13073;
  assign n14585 = ~n666 & n14584;
  assign n14586 = n1679 & n14585;
  assign n14587 = ~n544 & n14586;
  assign n14588 = ~n213 & n14587;
  assign n14589 = n14583 & n14588;
  assign n14590 = n276 & n14347;
  assign n14591 = ~n578 & n14590;
  assign n14592 = ~n272 & n14591;
  assign n14593 = n2683 & n12589;
  assign n14594 = n2021 & n14593;
  assign n14595 = n1401 & n14594;
  assign n14596 = n237 & n14595;
  assign n14597 = ~n341 & n14596;
  assign n14598 = ~n473 & n14597;
  assign n14599 = n14592 & n14598;
  assign n14600 = n14589 & n14599;
  assign n14601 = ~n14365 & ~n14600;
  assign n14602 = n14365 & n14600;
  assign n14603 = ~n14601 & ~n14602;
  assign n14604 = ~n372 & n3704;
  assign n14605 = ~n147 & n14604;
  assign n14606 = ~n547 & n14605;
  assign n14607 = n3195 & n4289;
  assign n14608 = n1390 & n14607;
  assign n14609 = n2131 & n14608;
  assign n14610 = ~n576 & n14609;
  assign n14611 = n515 & n2543;
  assign n14612 = ~n160 & n14611;
  assign n14613 = n14610 & n14612;
  assign n14614 = ~n320 & ~n461;
  assign n14615 = n2975 & n14614;
  assign n14616 = ~n112 & n14615;
  assign n14617 = ~n698 & n2321;
  assign n14618 = ~n350 & n14617;
  assign n14619 = n14616 & n14618;
  assign n14620 = n14613 & n14619;
  assign n14621 = n14606 & n14620;
  assign n14622 = ~n254 & ~n500;
  assign n14623 = n14621 & n14622;
  assign n14624 = ~n581 & n14623;
  assign n14625 = ~n705 & n2491;
  assign n14626 = ~n394 & n14625;
  assign n14627 = n14624 & n14626;
  assign n14628 = n1505 & n14627;
  assign n14629 = n2463 & n3443;
  assign n14630 = n14628 & n14629;
  assign n14631 = ~n308 & n14630;
  assign n14632 = ~n297 & n2060;
  assign n14633 = ~n382 & n14632;
  assign n14634 = n14631 & n14633;
  assign n14635 = ~n631 & ~n697;
  assign n14636 = ~n535 & n14635;
  assign n14637 = ~n305 & n14636;
  assign n14638 = ~n155 & ~n578;
  assign n14639 = ~n679 & n14638;
  assign n14640 = n960 & n14639;
  assign n14641 = n14637 & n14640;
  assign n14642 = n13029 & n14641;
  assign n14643 = ~n588 & n14642;
  assign n14644 = ~n277 & n14643;
  assign n14645 = n2327 & n13819;
  assign n14646 = ~n548 & n14645;
  assign n14647 = ~n610 & n14646;
  assign n14648 = n14644 & n14647;
  assign n14649 = n14634 & n14648;
  assign n14650 = ~n14365 & ~n14649;
  assign n14651 = n14365 & n14649;
  assign n14652 = n3641 & n12704;
  assign n14653 = n3740 & n12701;
  assign n14654 = n12764 & ~n12766;
  assign n14655 = ~n12767 & ~n14654;
  assign n14656 = n556 & n14655;
  assign n14657 = n3961 & n12698;
  assign n14658 = ~n14656 & ~n14657;
  assign n14659 = ~n14653 & n14658;
  assign n14660 = ~n14652 & n14659;
  assign n14661 = ~n14651 & ~n14660;
  assign n14662 = ~n14650 & ~n14661;
  assign n14663 = n14603 & ~n14662;
  assign n14664 = ~n14601 & ~n14663;
  assign n14665 = n14365 & n14578;
  assign n14666 = ~n14579 & ~n14665;
  assign n14667 = ~n14664 & n14666;
  assign n14668 = ~n14579 & ~n14667;
  assign n14669 = n14369 & ~n14374;
  assign n14670 = ~n14375 & ~n14669;
  assign n14671 = ~n14668 & n14670;
  assign n14672 = n14668 & ~n14670;
  assign n14673 = ~n14671 & ~n14672;
  assign n14674 = n3641 & n12695;
  assign n14675 = n3740 & n12692;
  assign n14676 = n12776 & ~n12778;
  assign n14677 = ~n12779 & ~n14676;
  assign n14678 = n556 & n14677;
  assign n14679 = n3961 & n12689;
  assign n14680 = ~n14678 & ~n14679;
  assign n14681 = ~n14675 & n14680;
  assign n14682 = ~n14674 & n14681;
  assign n14683 = n14673 & ~n14682;
  assign n14684 = ~n14671 & ~n14683;
  assign n14685 = ~n14379 & n14388;
  assign n14686 = ~n14389 & ~n14685;
  assign n14687 = ~n14684 & n14686;
  assign n14688 = n14684 & ~n14686;
  assign n14689 = ~n14687 & ~n14688;
  assign n14690 = n4006 & n12683;
  assign n14691 = n4133 & n12680;
  assign n14692 = n4002 & n13929;
  assign n14693 = n4555 & n12677;
  assign n14694 = ~n14692 & ~n14693;
  assign n14695 = ~n14691 & n14694;
  assign n14696 = ~n14690 & n14695;
  assign n14697 = pi29  & n14696;
  assign n14698 = ~pi29  & ~n14696;
  assign n14699 = ~n14697 & ~n14698;
  assign n14700 = n14689 & ~n14699;
  assign n14701 = ~n14687 & ~n14700;
  assign n14702 = ~n14561 & ~n14701;
  assign n14703 = ~n14558 & ~n14702;
  assign n14704 = n14541 & ~n14545;
  assign n14705 = ~n14546 & ~n14704;
  assign n14706 = ~n14703 & n14705;
  assign n14707 = ~n14546 & ~n14706;
  assign n14708 = ~n14412 & n14422;
  assign n14709 = ~n14423 & ~n14708;
  assign n14710 = ~n14707 & n14709;
  assign n14711 = n14707 & ~n14709;
  assign n14712 = n4601 & n12665;
  assign n14713 = n4783 & n12662;
  assign n14714 = n4602 & n13165;
  assign n14715 = n4801 & n12659;
  assign n14716 = ~n14714 & ~n14715;
  assign n14717 = ~n14713 & n14716;
  assign n14718 = ~n14712 & n14717;
  assign n14719 = pi26  & n14718;
  assign n14720 = ~pi26  & ~n14718;
  assign n14721 = ~n14719 & ~n14720;
  assign n14722 = ~n14711 & ~n14721;
  assign n14723 = ~n14710 & ~n14722;
  assign n14724 = n14531 & ~n14723;
  assign n14725 = ~n14531 & n14723;
  assign n14726 = n5238 & n12653;
  assign n14727 = n71 & n12650;
  assign n14728 = n5239 & n13042;
  assign n14729 = n5326 & n12647;
  assign n14730 = ~n14728 & ~n14729;
  assign n14731 = ~n14727 & n14730;
  assign n14732 = ~n14726 & n14731;
  assign n14733 = pi23  & n14732;
  assign n14734 = ~pi23  & ~n14732;
  assign n14735 = ~n14733 & ~n14734;
  assign n14736 = ~n14725 & ~n14735;
  assign n14737 = ~n14724 & ~n14736;
  assign n14738 = ~n14527 & ~n14737;
  assign n14739 = ~n14524 & ~n14738;
  assign n14740 = ~n14447 & ~n14448;
  assign n14741 = ~n14458 & n14740;
  assign n14742 = n14458 & ~n14740;
  assign n14743 = ~n14741 & ~n14742;
  assign n14744 = ~n14739 & n14743;
  assign n14745 = n14739 & ~n14743;
  assign n14746 = n5435 & n12636;
  assign n14747 = n6055 & n12633;
  assign n14748 = n5429 & n13292;
  assign n14749 = n6071 & n12630;
  assign n14750 = ~n14748 & ~n14749;
  assign n14751 = ~n14747 & n14750;
  assign n14752 = ~n14746 & n14751;
  assign n14753 = pi20  & n14752;
  assign n14754 = ~pi20  & ~n14752;
  assign n14755 = ~n14753 & ~n14754;
  assign n14756 = ~n14745 & ~n14755;
  assign n14757 = ~n14744 & ~n14756;
  assign n14758 = n14511 & ~n14757;
  assign n14759 = ~n14511 & n14757;
  assign n14760 = n6184 & n12622;
  assign n14761 = n6527 & n12614;
  assign n14762 = n6185 & ~n13310;
  assign n14763 = n6543 & n12606;
  assign n14764 = ~n14762 & ~n14763;
  assign n14765 = ~n14761 & n14764;
  assign n14766 = ~n14760 & n14765;
  assign n14767 = pi17  & n14766;
  assign n14768 = ~pi17  & ~n14766;
  assign n14769 = ~n14767 & ~n14768;
  assign n14770 = ~n14759 & ~n14769;
  assign n14771 = ~n14758 & ~n14770;
  assign n14772 = ~n14507 & ~n14771;
  assign n14773 = n14279 & n14474;
  assign n14774 = ~n14475 & ~n14773;
  assign n14775 = n14507 & ~n14771;
  assign n14776 = ~n14507 & n14771;
  assign n14777 = ~n14775 & ~n14776;
  assign n14778 = n14774 & ~n14777;
  assign n14779 = ~n14772 & ~n14778;
  assign n14780 = ~n14481 & ~n14482;
  assign n14781 = ~n14492 & n14780;
  assign n14782 = n14492 & ~n14780;
  assign n14783 = ~n14781 & ~n14782;
  assign n14784 = ~n14779 & n14783;
  assign n14785 = n14779 & n14783;
  assign n14786 = ~n14779 & ~n14783;
  assign n14787 = ~n14785 & ~n14786;
  assign n14788 = ~n14774 & n14777;
  assign n14789 = ~n14778 & ~n14788;
  assign n14790 = n6836 & ~n13499;
  assign n14791 = n6835 & ~n12611;
  assign n14792 = ~n7460 & ~n7487;
  assign n14793 = ~n14791 & n14792;
  assign n14794 = ~n12608 & ~n14793;
  assign n14795 = ~n14790 & ~n14794;
  assign n14796 = pi14  & n14795;
  assign n14797 = ~pi14  & ~n14795;
  assign n14798 = ~n14796 & ~n14797;
  assign n14799 = n14527 & n14737;
  assign n14800 = ~n14738 & ~n14799;
  assign n14801 = n5435 & n12639;
  assign n14802 = n6055 & n12636;
  assign n14803 = n5429 & n13396;
  assign n14804 = n6071 & n12633;
  assign n14805 = ~n14803 & ~n14804;
  assign n14806 = ~n14802 & n14805;
  assign n14807 = ~n14801 & n14806;
  assign n14808 = pi20  & n14807;
  assign n14809 = ~pi20  & ~n14807;
  assign n14810 = ~n14808 & ~n14809;
  assign n14811 = n14800 & ~n14810;
  assign n14812 = n14800 & n14810;
  assign n14813 = ~n14800 & ~n14810;
  assign n14814 = ~n14812 & ~n14813;
  assign n14815 = ~n14724 & ~n14725;
  assign n14816 = ~n14735 & n14815;
  assign n14817 = n14735 & ~n14815;
  assign n14818 = ~n14816 & ~n14817;
  assign n14819 = n14703 & ~n14705;
  assign n14820 = ~n14706 & ~n14819;
  assign n14821 = n4601 & n12668;
  assign n14822 = n4783 & n12665;
  assign n14823 = n4602 & n13591;
  assign n14824 = n4801 & n12662;
  assign n14825 = ~n14823 & ~n14824;
  assign n14826 = ~n14822 & n14825;
  assign n14827 = ~n14821 & n14826;
  assign n14828 = pi26  & n14827;
  assign n14829 = ~pi26  & ~n14827;
  assign n14830 = ~n14828 & ~n14829;
  assign n14831 = n14820 & ~n14830;
  assign n14832 = n14820 & n14830;
  assign n14833 = ~n14820 & ~n14830;
  assign n14834 = ~n14832 & ~n14833;
  assign n14835 = n14561 & n14701;
  assign n14836 = ~n14702 & ~n14835;
  assign n14837 = n4006 & n12680;
  assign n14838 = n4133 & n12677;
  assign n14839 = n4002 & n14164;
  assign n14840 = n4555 & n12674;
  assign n14841 = ~n14839 & ~n14840;
  assign n14842 = ~n14838 & n14841;
  assign n14843 = ~n14837 & n14842;
  assign n14844 = pi29  & n14843;
  assign n14845 = ~pi29  & ~n14843;
  assign n14846 = ~n14844 & ~n14845;
  assign n14847 = n14836 & ~n14846;
  assign n14848 = n14836 & n14846;
  assign n14849 = ~n14836 & ~n14846;
  assign n14850 = ~n14848 & ~n14849;
  assign n14851 = n4601 & n12671;
  assign n14852 = n4783 & n12668;
  assign n14853 = n4602 & n13578;
  assign n14854 = n4801 & n12665;
  assign n14855 = ~n14853 & ~n14854;
  assign n14856 = ~n14852 & n14855;
  assign n14857 = ~n14851 & n14856;
  assign n14858 = pi26  & n14857;
  assign n14859 = ~pi26  & ~n14857;
  assign n14860 = ~n14858 & ~n14859;
  assign n14861 = ~n14850 & ~n14860;
  assign n14862 = ~n14847 & ~n14861;
  assign n14863 = ~n14834 & ~n14862;
  assign n14864 = ~n14831 & ~n14863;
  assign n14865 = ~n14710 & ~n14711;
  assign n14866 = ~n14721 & n14865;
  assign n14867 = n14721 & ~n14865;
  assign n14868 = ~n14866 & ~n14867;
  assign n14869 = ~n14864 & n14868;
  assign n14870 = n14864 & ~n14868;
  assign n14871 = n5238 & n12656;
  assign n14872 = n71 & n12653;
  assign n14873 = n5239 & n12991;
  assign n14874 = n5326 & n12650;
  assign n14875 = ~n14873 & ~n14874;
  assign n14876 = ~n14872 & n14875;
  assign n14877 = ~n14871 & n14876;
  assign n14878 = pi23  & n14877;
  assign n14879 = ~pi23  & ~n14877;
  assign n14880 = ~n14878 & ~n14879;
  assign n14881 = ~n14870 & ~n14880;
  assign n14882 = ~n14869 & ~n14881;
  assign n14883 = n14818 & ~n14882;
  assign n14884 = ~n14818 & n14882;
  assign n14885 = n5435 & n12644;
  assign n14886 = n6055 & n12639;
  assign n14887 = n5429 & n13210;
  assign n14888 = n6071 & n12636;
  assign n14889 = ~n14887 & ~n14888;
  assign n14890 = ~n14886 & n14889;
  assign n14891 = ~n14885 & n14890;
  assign n14892 = pi20  & n14891;
  assign n14893 = ~pi20  & ~n14891;
  assign n14894 = ~n14892 & ~n14893;
  assign n14895 = ~n14884 & ~n14894;
  assign n14896 = ~n14883 & ~n14895;
  assign n14897 = ~n14814 & ~n14896;
  assign n14898 = ~n14811 & ~n14897;
  assign n14899 = ~n14744 & ~n14745;
  assign n14900 = ~n14755 & n14899;
  assign n14901 = n14755 & ~n14899;
  assign n14902 = ~n14900 & ~n14901;
  assign n14903 = ~n14898 & n14902;
  assign n14904 = n14898 & ~n14902;
  assign n14905 = n6184 & n12625;
  assign n14906 = n6527 & n12622;
  assign n14907 = n6185 & n13463;
  assign n14908 = n6543 & n12614;
  assign n14909 = ~n14907 & ~n14908;
  assign n14910 = ~n14906 & n14909;
  assign n14911 = ~n14905 & n14910;
  assign n14912 = pi17  & n14911;
  assign n14913 = ~pi17  & ~n14911;
  assign n14914 = ~n14912 & ~n14913;
  assign n14915 = ~n14904 & ~n14914;
  assign n14916 = ~n14903 & ~n14915;
  assign n14917 = ~n14798 & ~n14916;
  assign n14918 = n14798 & n14916;
  assign n14919 = ~n14758 & ~n14759;
  assign n14920 = ~n14769 & n14919;
  assign n14921 = n14769 & ~n14919;
  assign n14922 = ~n14920 & ~n14921;
  assign n14923 = ~n14918 & n14922;
  assign n14924 = ~n14917 & ~n14923;
  assign n14925 = n14789 & ~n14924;
  assign n14926 = ~n14917 & ~n14918;
  assign n14927 = n14922 & n14926;
  assign n14928 = ~n14922 & ~n14926;
  assign n14929 = ~n14927 & ~n14928;
  assign n14930 = n14814 & n14896;
  assign n14931 = ~n14897 & ~n14930;
  assign n14932 = n6184 & n12630;
  assign n14933 = n6527 & n12625;
  assign n14934 = n6185 & n13325;
  assign n14935 = n6543 & n12622;
  assign n14936 = ~n14934 & ~n14935;
  assign n14937 = ~n14933 & n14936;
  assign n14938 = ~n14932 & n14937;
  assign n14939 = pi17  & n14938;
  assign n14940 = ~pi17  & ~n14938;
  assign n14941 = ~n14939 & ~n14940;
  assign n14942 = n14931 & ~n14941;
  assign n14943 = n14931 & n14941;
  assign n14944 = ~n14931 & ~n14941;
  assign n14945 = ~n14943 & ~n14944;
  assign n14946 = ~n14883 & ~n14884;
  assign n14947 = ~n14894 & n14946;
  assign n14948 = n14894 & ~n14946;
  assign n14949 = ~n14947 & ~n14948;
  assign n14950 = n14834 & n14862;
  assign n14951 = ~n14863 & ~n14950;
  assign n14952 = n5238 & n12659;
  assign n14953 = n71 & n12656;
  assign n14954 = n5239 & n13059;
  assign n14955 = n5326 & n12653;
  assign n14956 = ~n14954 & ~n14955;
  assign n14957 = ~n14953 & n14956;
  assign n14958 = ~n14952 & n14957;
  assign n14959 = pi23  & n14958;
  assign n14960 = ~pi23  & ~n14958;
  assign n14961 = ~n14959 & ~n14960;
  assign n14962 = n14951 & ~n14961;
  assign n14963 = n14951 & n14961;
  assign n14964 = ~n14951 & ~n14961;
  assign n14965 = ~n14963 & ~n14964;
  assign n14966 = ~n14850 & n14860;
  assign n14967 = n14850 & ~n14860;
  assign n14968 = ~n14966 & ~n14967;
  assign n14969 = ~n14689 & n14699;
  assign n14970 = ~n14700 & ~n14969;
  assign n14971 = n14664 & ~n14666;
  assign n14972 = ~n14667 & ~n14971;
  assign n14973 = n3641 & n12698;
  assign n14974 = n3740 & n12695;
  assign n14975 = n12772 & ~n12774;
  assign n14976 = ~n12775 & ~n14975;
  assign n14977 = n556 & n14976;
  assign n14978 = n3961 & n12692;
  assign n14979 = ~n14977 & ~n14978;
  assign n14980 = ~n14974 & n14979;
  assign n14981 = ~n14973 & n14980;
  assign n14982 = n14972 & ~n14981;
  assign n14983 = n14972 & n14981;
  assign n14984 = ~n14972 & ~n14981;
  assign n14985 = ~n14983 & ~n14984;
  assign n14986 = ~n14603 & n14662;
  assign n14987 = ~n14663 & ~n14986;
  assign n14988 = n3641 & n12701;
  assign n14989 = n3740 & n12698;
  assign n14990 = n12768 & ~n12770;
  assign n14991 = ~n12771 & ~n14990;
  assign n14992 = n556 & n14991;
  assign n14993 = n3961 & n12695;
  assign n14994 = ~n14992 & ~n14993;
  assign n14995 = ~n14989 & n14994;
  assign n14996 = ~n14988 & n14995;
  assign n14997 = n14987 & ~n14996;
  assign n14998 = n14987 & n14996;
  assign n14999 = ~n14987 & ~n14996;
  assign n15000 = ~n14998 & ~n14999;
  assign n15001 = n3392 & n4441;
  assign n15002 = ~n186 & n15001;
  assign n15003 = ~n116 & ~n150;
  assign n15004 = ~n171 & n15003;
  assign n15005 = ~n685 & n4037;
  assign n15006 = ~n668 & n15005;
  assign n15007 = n15004 & n15006;
  assign n15008 = n1252 & n15007;
  assign n15009 = n901 & n15008;
  assign n15010 = ~n517 & n15009;
  assign n15011 = n15002 & n15010;
  assign n15012 = n1116 & n3367;
  assign n15013 = n1570 & n15012;
  assign n15014 = n5482 & n15013;
  assign n15015 = n706 & n15014;
  assign n15016 = ~n360 & n15015;
  assign n15017 = n2986 & n13722;
  assign n15018 = ~n337 & n15017;
  assign n15019 = ~n98 & n15018;
  assign n15020 = n15016 & n15019;
  assign n15021 = n15011 & n15020;
  assign n15022 = n3641 & n12707;
  assign n15023 = n12760 & ~n12762;
  assign n15024 = ~n12763 & ~n15023;
  assign n15025 = n556 & n15024;
  assign n15026 = n3961 & n12701;
  assign n15027 = n3740 & n12704;
  assign n15028 = ~n15026 & ~n15027;
  assign n15029 = ~n15025 & n15028;
  assign n15030 = ~n15022 & n15029;
  assign n15031 = ~n15021 & ~n15030;
  assign n15032 = ~n632 & n1341;
  assign n15033 = ~n670 & n15032;
  assign n15034 = n1489 & n3782;
  assign n15035 = n6614 & n15034;
  assign n15036 = ~n98 & n15035;
  assign n15037 = n15033 & n15036;
  assign n15038 = n3107 & n3460;
  assign n15039 = n528 & n15038;
  assign n15040 = ~n289 & n15039;
  assign n15041 = n1982 & n4353;
  assign n15042 = n3442 & n15041;
  assign n15043 = n1840 & n15042;
  assign n15044 = ~n538 & n15043;
  assign n15045 = ~n439 & n15044;
  assign n15046 = n15040 & n15045;
  assign n15047 = n15037 & n15046;
  assign n15048 = n3641 & n12710;
  assign n15049 = n12756 & ~n12758;
  assign n15050 = ~n12759 & ~n15049;
  assign n15051 = n556 & n15050;
  assign n15052 = n3961 & n12704;
  assign n15053 = n3740 & n12707;
  assign n15054 = ~n15052 & ~n15053;
  assign n15055 = ~n15051 & n15054;
  assign n15056 = ~n15048 & n15055;
  assign n15057 = ~n15047 & ~n15056;
  assign n15058 = n1783 & n14627;
  assign n15059 = ~n255 & n15058;
  assign n15060 = n1892 & n3250;
  assign n15061 = ~n401 & n15060;
  assign n15062 = n15059 & n15061;
  assign n15063 = ~n701 & n5105;
  assign n15064 = ~n398 & n15063;
  assign n15065 = n2428 & n3301;
  assign n15066 = n2488 & n15065;
  assign n15067 = n359 & n2365;
  assign n15068 = n15066 & n15067;
  assign n15069 = ~n589 & n15068;
  assign n15070 = n15064 & n15069;
  assign n15071 = n15062 & n15070;
  assign n15072 = n3641 & n12713;
  assign n15073 = n12752 & ~n12754;
  assign n15074 = ~n12755 & ~n15073;
  assign n15075 = n556 & n15074;
  assign n15076 = n3961 & n12707;
  assign n15077 = n3740 & n12710;
  assign n15078 = ~n15076 & ~n15077;
  assign n15079 = ~n15075 & n15078;
  assign n15080 = ~n15072 & n15079;
  assign n15081 = ~n15071 & ~n15080;
  assign n15082 = n916 & n2365;
  assign n15083 = ~n393 & n15082;
  assign n15084 = n467 & n4256;
  assign n15085 = ~n436 & n15084;
  assign n15086 = ~n144 & n15085;
  assign n15087 = n15083 & n15086;
  assign n15088 = ~n173 & n1742;
  assign n15089 = ~n442 & ~n628;
  assign n15090 = n237 & n15089;
  assign n15091 = ~n314 & n15090;
  assign n15092 = n15088 & n15091;
  assign n15093 = n1147 & n4517;
  assign n15094 = n2065 & n15093;
  assign n15095 = n15092 & n15094;
  assign n15096 = ~n290 & n15095;
  assign n15097 = n3771 & n4237;
  assign n15098 = n343 & n15097;
  assign n15099 = ~n304 & n15098;
  assign n15100 = ~n98 & n15099;
  assign n15101 = n15096 & n15100;
  assign n15102 = n15087 & n15101;
  assign n15103 = n3641 & n12716;
  assign n15104 = n12748 & ~n12750;
  assign n15105 = ~n12751 & ~n15104;
  assign n15106 = n556 & n15105;
  assign n15107 = n3961 & n12710;
  assign n15108 = n3740 & n12713;
  assign n15109 = ~n15107 & ~n15108;
  assign n15110 = ~n15106 & n15109;
  assign n15111 = ~n15103 & n15110;
  assign n15112 = ~n15102 & ~n15111;
  assign n15113 = n317 & n7043;
  assign n15114 = n237 & n15113;
  assign n15115 = ~n576 & n15114;
  assign n15116 = n2683 & n13538;
  assign n15117 = n1934 & n15116;
  assign n15118 = n148 & n15117;
  assign n15119 = ~n163 & n15118;
  assign n15120 = ~n187 & n15119;
  assign n15121 = n15115 & n15120;
  assign n15122 = ~n115 & ~n505;
  assign n15123 = ~n160 & n15122;
  assign n15124 = n1576 & n15123;
  assign n15125 = n2340 & n15124;
  assign n15126 = ~n100 & n15125;
  assign n15127 = n2229 & n4888;
  assign n15128 = ~n123 & n15127;
  assign n15129 = ~n341 & n15128;
  assign n15130 = n15126 & n15129;
  assign n15131 = ~n590 & n4452;
  assign n15132 = ~n214 & n15131;
  assign n15133 = ~n391 & n7167;
  assign n15134 = ~n517 & n15133;
  assign n15135 = n15132 & n15134;
  assign n15136 = n15130 & n15135;
  assign n15137 = n367 & n2975;
  assign n15138 = n797 & n15137;
  assign n15139 = ~n78 & n15138;
  assign n15140 = n546 & n13848;
  assign n15141 = ~n468 & n15140;
  assign n15142 = n15139 & n15141;
  assign n15143 = n459 & n5894;
  assign n15144 = ~n454 & n15143;
  assign n15145 = n378 & n3771;
  assign n15146 = n1109 & n15145;
  assign n15147 = ~n413 & n15146;
  assign n15148 = n15144 & n15147;
  assign n15149 = n15142 & n15148;
  assign n15150 = n3409 & n15149;
  assign n15151 = n15136 & n15150;
  assign n15152 = ~n682 & n15151;
  assign n15153 = n3835 & n7097;
  assign n15154 = n2099 & n15153;
  assign n15155 = ~n207 & n15154;
  assign n15156 = ~n394 & n15155;
  assign n15157 = n15152 & n15156;
  assign n15158 = n15121 & n15157;
  assign n15159 = n3641 & n12719;
  assign n15160 = n12744 & ~n12746;
  assign n15161 = ~n12747 & ~n15160;
  assign n15162 = n556 & n15161;
  assign n15163 = n3961 & n12713;
  assign n15164 = n3740 & n12716;
  assign n15165 = ~n15163 & ~n15164;
  assign n15166 = ~n15162 & n15165;
  assign n15167 = ~n15159 & n15166;
  assign n15168 = ~n15158 & ~n15167;
  assign n15169 = n3158 & n4065;
  assign n15170 = n230 & n15169;
  assign n15171 = ~n255 & n15170;
  assign n15172 = n1169 & n2623;
  assign n15173 = ~n590 & n15172;
  assign n15174 = ~n544 & n15173;
  assign n15175 = n15171 & n15174;
  assign n15176 = ~n363 & n12564;
  assign n15177 = ~n88 & n15176;
  assign n15178 = n1587 & n3936;
  assign n15179 = ~n436 & n15178;
  assign n15180 = n3187 & n4079;
  assign n15181 = ~n533 & n15180;
  assign n15182 = n15179 & n15181;
  assign n15183 = n107 & n13904;
  assign n15184 = ~n170 & n15183;
  assign n15185 = n946 & n2076;
  assign n15186 = n2021 & n15185;
  assign n15187 = n1964 & n15186;
  assign n15188 = n1272 & n15187;
  assign n15189 = ~n704 & n15188;
  assign n15190 = n15184 & n15189;
  assign n15191 = n15182 & n15190;
  assign n15192 = n1708 & n15191;
  assign n15193 = ~n637 & n15192;
  assign n15194 = ~n325 & n15193;
  assign n15195 = n15177 & n15194;
  assign n15196 = n15175 & n15195;
  assign n15197 = n3641 & n12722;
  assign n15198 = n12740 & ~n12742;
  assign n15199 = ~n12743 & ~n15198;
  assign n15200 = n556 & n15199;
  assign n15201 = n3961 & n12716;
  assign n15202 = n3740 & n12719;
  assign n15203 = ~n15201 & ~n15202;
  assign n15204 = ~n15200 & n15203;
  assign n15205 = ~n15197 & n15204;
  assign n15206 = ~n15196 & ~n15205;
  assign n15207 = n2070 & n3042;
  assign n15208 = ~n428 & n15207;
  assign n15209 = n1936 & n2350;
  assign n15210 = ~n373 & n15209;
  assign n15211 = n15208 & n15210;
  assign n15212 = ~n171 & n1634;
  assign n15213 = n12934 & n15212;
  assign n15214 = n1271 & n15213;
  assign n15215 = ~n281 & n15214;
  assign n15216 = ~n273 & n3159;
  assign n15217 = ~n427 & n15216;
  assign n15218 = ~n219 & n15217;
  assign n15219 = n15215 & n15218;
  assign n15220 = ~n197 & n4444;
  assign n15221 = ~n581 & n981;
  assign n15222 = ~n501 & n15221;
  assign n15223 = n15220 & n15222;
  assign n15224 = n386 & n15223;
  assign n15225 = ~n578 & n15224;
  assign n15226 = ~n231 & n15225;
  assign n15227 = n392 & n13835;
  assign n15228 = ~n147 & n15227;
  assign n15229 = ~n251 & n15228;
  assign n15230 = n15226 & n15229;
  assign n15231 = n15219 & n15230;
  assign n15232 = n1521 & n15231;
  assign n15233 = ~n678 & n15232;
  assign n15234 = n156 & n5525;
  assign n15235 = n2502 & n15234;
  assign n15236 = n2997 & n15235;
  assign n15237 = ~n504 & n15236;
  assign n15238 = ~n589 & n15237;
  assign n15239 = n15233 & n15238;
  assign n15240 = n15211 & n15239;
  assign n15241 = n3641 & n12725;
  assign n15242 = n12736 & ~n12738;
  assign n15243 = ~n12739 & ~n15242;
  assign n15244 = n556 & n15243;
  assign n15245 = n3961 & n12719;
  assign n15246 = n3740 & n12722;
  assign n15247 = ~n15245 & ~n15246;
  assign n15248 = ~n15244 & n15247;
  assign n15249 = ~n15241 & n15248;
  assign n15250 = ~n15240 & ~n15249;
  assign n15251 = n282 & n3675;
  assign n15252 = ~n194 & n15251;
  assign n15253 = ~n588 & n15252;
  assign n15254 = n3347 & n4498;
  assign n15255 = n4492 & n15254;
  assign n15256 = n643 & n15255;
  assign n15257 = ~n180 & n15256;
  assign n15258 = n1539 & n7091;
  assign n15259 = n5942 & n15258;
  assign n15260 = n343 & n15259;
  assign n15261 = ~n538 & n15260;
  assign n15262 = n15257 & n15261;
  assign n15263 = n3767 & n15262;
  assign n15264 = n15253 & n15263;
  assign n15265 = n3641 & n12730;
  assign n15266 = ~n12728 & ~n12734;
  assign n15267 = ~n12735 & ~n15266;
  assign n15268 = n556 & n15267;
  assign n15269 = n3961 & n12722;
  assign n15270 = n3740 & n12725;
  assign n15271 = ~n15269 & ~n15270;
  assign n15272 = ~n15268 & n15271;
  assign n15273 = ~n15265 & n15272;
  assign n15274 = ~n15264 & ~n15273;
  assign n15275 = ~n15264 & n15273;
  assign n15276 = n15264 & ~n15273;
  assign n15277 = ~n15275 & ~n15276;
  assign n15278 = n2269 & n3132;
  assign n15279 = n2417 & n15278;
  assign n15280 = ~n243 & n15279;
  assign n15281 = ~n332 & ~n341;
  assign n15282 = n2000 & n15281;
  assign n15283 = ~n527 & n15282;
  assign n15284 = ~n279 & n2991;
  assign n15285 = ~n238 & n15284;
  assign n15286 = n15283 & n15285;
  assign n15287 = n907 & n15286;
  assign n15288 = ~n297 & n15287;
  assign n15289 = n1012 & n3890;
  assign n15290 = ~n669 & n15289;
  assign n15291 = n15288 & n15290;
  assign n15292 = n616 & n741;
  assign n15293 = ~n229 & n15292;
  assign n15294 = n1089 & n15092;
  assign n15295 = n392 & n15294;
  assign n15296 = ~n245 & n15295;
  assign n15297 = n15293 & n15296;
  assign n15298 = n15291 & n15297;
  assign n15299 = n7210 & n15298;
  assign n15300 = ~n544 & n15299;
  assign n15301 = n15280 & n15300;
  assign n15302 = n804 & n2825;
  assign n15303 = n515 & n15302;
  assign n15304 = ~n171 & n15303;
  assign n15305 = n2856 & n2923;
  assign n15306 = ~n578 & n15305;
  assign n15307 = ~n323 & n15306;
  assign n15308 = n15304 & n15307;
  assign n15309 = n15301 & n15308;
  assign n15310 = n12730 & ~n12732;
  assign n15311 = ~n12730 & n12732;
  assign n15312 = ~n15310 & ~n15311;
  assign n15313 = n556 & ~n15312;
  assign n15314 = n3740 & n12732;
  assign n15315 = n3961 & n12730;
  assign n15316 = ~n15314 & ~n15315;
  assign n15317 = ~n15313 & n15316;
  assign n15318 = ~n15309 & ~n15317;
  assign n15319 = n3704 & n13825;
  assign n15320 = ~n593 & n15319;
  assign n15321 = ~n672 & n15320;
  assign n15322 = n584 & n4049;
  assign n15323 = n1551 & n15322;
  assign n15324 = n1261 & n15323;
  assign n15325 = n1132 & n15324;
  assign n15326 = ~n538 & n15325;
  assign n15327 = ~n293 & n15326;
  assign n15328 = n15321 & n15327;
  assign n15329 = n2064 & n14641;
  assign n15330 = ~n356 & n15329;
  assign n15331 = ~n116 & n15330;
  assign n15332 = n1908 & n2269;
  assign n15333 = ~n670 & n15332;
  assign n15334 = n416 & n1742;
  assign n15335 = ~n610 & n15334;
  assign n15336 = ~n129 & n15335;
  assign n15337 = n15333 & n15336;
  assign n15338 = ~n502 & n15337;
  assign n15339 = ~n588 & ~n700;
  assign n15340 = ~n112 & n15339;
  assign n15341 = n1646 & n1708;
  assign n15342 = ~n465 & n15341;
  assign n15343 = n15340 & n15342;
  assign n15344 = n15338 & n15343;
  assign n15345 = ~n666 & n15344;
  assign n15346 = ~n243 & n15345;
  assign n15347 = ~n323 & n15346;
  assign n15348 = n15331 & n15347;
  assign n15349 = n15328 & n15348;
  assign n15350 = n15318 & ~n15349;
  assign n15351 = ~n15318 & n15349;
  assign n15352 = n3641 & n12732;
  assign n15353 = n3740 & n12730;
  assign n15354 = n12725 & ~n15310;
  assign n15355 = ~n12725 & n15310;
  assign n15356 = ~n15354 & ~n15355;
  assign n15357 = n556 & ~n15356;
  assign n15358 = n3961 & n12725;
  assign n15359 = ~n15357 & ~n15358;
  assign n15360 = ~n15353 & n15359;
  assign n15361 = ~n15352 & n15360;
  assign n15362 = ~n15351 & ~n15361;
  assign n15363 = ~n15350 & ~n15362;
  assign n15364 = ~n15277 & ~n15363;
  assign n15365 = ~n15274 & ~n15364;
  assign n15366 = ~n15240 & n15249;
  assign n15367 = n15240 & ~n15249;
  assign n15368 = ~n15366 & ~n15367;
  assign n15369 = ~n15365 & ~n15368;
  assign n15370 = ~n15250 & ~n15369;
  assign n15371 = ~n15196 & n15205;
  assign n15372 = n15196 & ~n15205;
  assign n15373 = ~n15371 & ~n15372;
  assign n15374 = ~n15370 & ~n15373;
  assign n15375 = ~n15206 & ~n15374;
  assign n15376 = ~n15158 & n15167;
  assign n15377 = n15158 & ~n15167;
  assign n15378 = ~n15376 & ~n15377;
  assign n15379 = ~n15375 & ~n15378;
  assign n15380 = ~n15168 & ~n15379;
  assign n15381 = ~n15102 & n15111;
  assign n15382 = n15102 & ~n15111;
  assign n15383 = ~n15381 & ~n15382;
  assign n15384 = ~n15380 & ~n15383;
  assign n15385 = ~n15112 & ~n15384;
  assign n15386 = ~n15071 & n15080;
  assign n15387 = n15071 & ~n15080;
  assign n15388 = ~n15386 & ~n15387;
  assign n15389 = ~n15385 & ~n15388;
  assign n15390 = ~n15081 & ~n15389;
  assign n15391 = ~n15047 & n15056;
  assign n15392 = n15047 & ~n15056;
  assign n15393 = ~n15391 & ~n15392;
  assign n15394 = ~n15390 & ~n15393;
  assign n15395 = ~n15057 & ~n15394;
  assign n15396 = ~n15021 & n15030;
  assign n15397 = n15021 & ~n15030;
  assign n15398 = ~n15396 & ~n15397;
  assign n15399 = ~n15395 & ~n15398;
  assign n15400 = ~n15031 & ~n15399;
  assign n15401 = ~n14650 & ~n14651;
  assign n15402 = ~n14660 & n15401;
  assign n15403 = n14660 & ~n15401;
  assign n15404 = ~n15402 & ~n15403;
  assign n15405 = ~n15400 & n15404;
  assign n15406 = n15400 & ~n15404;
  assign n15407 = ~n15405 & ~n15406;
  assign n15408 = n4006 & n12695;
  assign n15409 = n4133 & n12692;
  assign n15410 = n4002 & n14677;
  assign n15411 = n4555 & n12689;
  assign n15412 = ~n15410 & ~n15411;
  assign n15413 = ~n15409 & n15412;
  assign n15414 = ~n15408 & n15413;
  assign n15415 = pi29  & n15414;
  assign n15416 = ~pi29  & ~n15414;
  assign n15417 = ~n15415 & ~n15416;
  assign n15418 = n15407 & ~n15417;
  assign n15419 = ~n15405 & ~n15418;
  assign n15420 = ~n15000 & ~n15419;
  assign n15421 = ~n14997 & ~n15420;
  assign n15422 = ~n14985 & ~n15421;
  assign n15423 = ~n14982 & ~n15422;
  assign n15424 = ~n14673 & n14682;
  assign n15425 = ~n14683 & ~n15424;
  assign n15426 = ~n15423 & n15425;
  assign n15427 = n15423 & ~n15425;
  assign n15428 = n4006 & n12686;
  assign n15429 = n4133 & n12683;
  assign n15430 = n4002 & n14402;
  assign n15431 = n4555 & n12680;
  assign n15432 = ~n15430 & ~n15431;
  assign n15433 = ~n15429 & n15432;
  assign n15434 = ~n15428 & n15433;
  assign n15435 = pi29  & n15434;
  assign n15436 = ~pi29  & ~n15434;
  assign n15437 = ~n15435 & ~n15436;
  assign n15438 = ~n15427 & ~n15437;
  assign n15439 = ~n15426 & ~n15438;
  assign n15440 = n14970 & ~n15439;
  assign n15441 = ~n14970 & n15439;
  assign n15442 = n4601 & n12674;
  assign n15443 = n4783 & n12671;
  assign n15444 = n4602 & n13764;
  assign n15445 = n4801 & n12668;
  assign n15446 = ~n15444 & ~n15445;
  assign n15447 = ~n15443 & n15446;
  assign n15448 = ~n15442 & n15447;
  assign n15449 = pi26  & n15448;
  assign n15450 = ~pi26  & ~n15448;
  assign n15451 = ~n15449 & ~n15450;
  assign n15452 = ~n15441 & ~n15451;
  assign n15453 = ~n15440 & ~n15452;
  assign n15454 = ~n14968 & ~n15453;
  assign n15455 = n14968 & n15453;
  assign n15456 = n5238 & n12662;
  assign n15457 = n71 & n12659;
  assign n15458 = n5239 & n13246;
  assign n15459 = n5326 & n12656;
  assign n15460 = ~n15458 & ~n15459;
  assign n15461 = ~n15457 & n15460;
  assign n15462 = ~n15456 & n15461;
  assign n15463 = pi23  & n15462;
  assign n15464 = ~pi23  & ~n15462;
  assign n15465 = ~n15463 & ~n15464;
  assign n15466 = ~n15455 & ~n15465;
  assign n15467 = ~n15454 & ~n15466;
  assign n15468 = ~n14965 & ~n15467;
  assign n15469 = ~n14962 & ~n15468;
  assign n15470 = ~n14869 & ~n14870;
  assign n15471 = ~n14880 & n15470;
  assign n15472 = n14880 & ~n15470;
  assign n15473 = ~n15471 & ~n15472;
  assign n15474 = ~n15469 & n15473;
  assign n15475 = n15469 & ~n15473;
  assign n15476 = n5435 & n12647;
  assign n15477 = n6055 & n12644;
  assign n15478 = n5429 & ~n13193;
  assign n15479 = n6071 & n12639;
  assign n15480 = ~n15478 & ~n15479;
  assign n15481 = ~n15477 & n15480;
  assign n15482 = ~n15476 & n15481;
  assign n15483 = pi20  & n15482;
  assign n15484 = ~pi20  & ~n15482;
  assign n15485 = ~n15483 & ~n15484;
  assign n15486 = ~n15475 & ~n15485;
  assign n15487 = ~n15474 & ~n15486;
  assign n15488 = n14949 & ~n15487;
  assign n15489 = ~n14949 & n15487;
  assign n15490 = n6184 & n12633;
  assign n15491 = n6527 & n12630;
  assign n15492 = n6185 & ~n13227;
  assign n15493 = n6543 & n12625;
  assign n15494 = ~n15492 & ~n15493;
  assign n15495 = ~n15491 & n15494;
  assign n15496 = ~n15490 & n15495;
  assign n15497 = pi17  & n15496;
  assign n15498 = ~pi17  & ~n15496;
  assign n15499 = ~n15497 & ~n15498;
  assign n15500 = ~n15489 & ~n15499;
  assign n15501 = ~n15488 & ~n15500;
  assign n15502 = ~n14945 & ~n15501;
  assign n15503 = ~n14942 & ~n15502;
  assign n15504 = ~n14903 & ~n14904;
  assign n15505 = ~n14914 & n15504;
  assign n15506 = n14914 & ~n15504;
  assign n15507 = ~n15505 & ~n15506;
  assign n15508 = ~n15503 & n15507;
  assign n15509 = n15503 & ~n15507;
  assign n15510 = n6835 & n12606;
  assign n15511 = n7460 & n12616;
  assign n15512 = n6836 & ~n13483;
  assign n15513 = n7487 & ~n12608;
  assign n15514 = ~n15512 & ~n15513;
  assign n15515 = ~n15511 & n15514;
  assign n15516 = ~n15510 & n15515;
  assign n15517 = pi14  & n15516;
  assign n15518 = ~pi14  & ~n15516;
  assign n15519 = ~n15517 & ~n15518;
  assign n15520 = ~n15509 & ~n15519;
  assign n15521 = ~n15508 & ~n15520;
  assign n15522 = n14929 & ~n15521;
  assign n15523 = ~n14929 & n15521;
  assign n15524 = ~n15522 & ~n15523;
  assign n15525 = n7460 & n12606;
  assign n15526 = ~n12611 & n15513;
  assign n15527 = n6835 & n12614;
  assign n15528 = n6836 & n12868;
  assign n15529 = ~n15527 & ~n15528;
  assign n15530 = ~n15526 & n15529;
  assign n15531 = ~n15525 & n15530;
  assign n15532 = pi14  & n15531;
  assign n15533 = ~pi14  & ~n15531;
  assign n15534 = ~n15532 & ~n15533;
  assign n15535 = ~n15488 & ~n15489;
  assign n15536 = ~n15499 & n15535;
  assign n15537 = n15499 & ~n15535;
  assign n15538 = ~n15536 & ~n15537;
  assign n15539 = n14965 & n15467;
  assign n15540 = ~n15468 & ~n15539;
  assign n15541 = n5435 & n12650;
  assign n15542 = n6055 & n12647;
  assign n15543 = n5429 & n13275;
  assign n15544 = n6071 & n12644;
  assign n15545 = ~n15543 & ~n15544;
  assign n15546 = ~n15542 & n15545;
  assign n15547 = ~n15541 & n15546;
  assign n15548 = pi20  & n15547;
  assign n15549 = ~pi20  & ~n15547;
  assign n15550 = ~n15548 & ~n15549;
  assign n15551 = n15540 & ~n15550;
  assign n15552 = n15540 & n15550;
  assign n15553 = ~n15540 & ~n15550;
  assign n15554 = ~n15552 & ~n15553;
  assign n15555 = ~n15454 & ~n15455;
  assign n15556 = ~n15465 & n15555;
  assign n15557 = n15465 & ~n15555;
  assign n15558 = ~n15556 & ~n15557;
  assign n15559 = n4601 & n12677;
  assign n15560 = n4783 & n12674;
  assign n15561 = n4602 & n13785;
  assign n15562 = n4801 & n12671;
  assign n15563 = ~n15561 & ~n15562;
  assign n15564 = ~n15560 & n15563;
  assign n15565 = ~n15559 & n15564;
  assign n15566 = pi26  & n15565;
  assign n15567 = ~pi26  & ~n15565;
  assign n15568 = ~n15566 & ~n15567;
  assign n15569 = ~n15426 & ~n15427;
  assign n15570 = ~n15437 & n15569;
  assign n15571 = n15437 & ~n15569;
  assign n15572 = ~n15570 & ~n15571;
  assign n15573 = ~n15568 & n15572;
  assign n15574 = n14985 & n15421;
  assign n15575 = ~n15422 & ~n15574;
  assign n15576 = n4006 & n12689;
  assign n15577 = n4133 & n12686;
  assign n15578 = n4002 & n14552;
  assign n15579 = n4555 & n12683;
  assign n15580 = ~n15578 & ~n15579;
  assign n15581 = ~n15577 & n15580;
  assign n15582 = ~n15576 & n15581;
  assign n15583 = pi29  & n15582;
  assign n15584 = ~pi29  & ~n15582;
  assign n15585 = ~n15583 & ~n15584;
  assign n15586 = n15575 & ~n15585;
  assign n15587 = n15575 & n15585;
  assign n15588 = ~n15575 & ~n15585;
  assign n15589 = ~n15587 & ~n15588;
  assign n15590 = n4783 & n12677;
  assign n15591 = n4801 & n12674;
  assign n15592 = n4602 & n14164;
  assign n15593 = n4601 & n12680;
  assign n15594 = ~n15592 & ~n15593;
  assign n15595 = ~n15591 & n15594;
  assign n15596 = ~n15590 & n15595;
  assign n15597 = pi26  & n15596;
  assign n15598 = ~pi26  & ~n15596;
  assign n15599 = ~n15597 & ~n15598;
  assign n15600 = ~n15589 & ~n15599;
  assign n15601 = ~n15586 & ~n15600;
  assign n15602 = n15568 & ~n15572;
  assign n15603 = ~n15573 & ~n15602;
  assign n15604 = ~n15601 & n15603;
  assign n15605 = ~n15573 & ~n15604;
  assign n15606 = ~n15440 & ~n15441;
  assign n15607 = ~n15451 & n15606;
  assign n15608 = n15451 & ~n15606;
  assign n15609 = ~n15607 & ~n15608;
  assign n15610 = ~n15605 & n15609;
  assign n15611 = n15605 & ~n15609;
  assign n15612 = n5238 & n12665;
  assign n15613 = n71 & n12662;
  assign n15614 = n5239 & n13165;
  assign n15615 = n5326 & n12659;
  assign n15616 = ~n15614 & ~n15615;
  assign n15617 = ~n15613 & n15616;
  assign n15618 = ~n15612 & n15617;
  assign n15619 = pi23  & n15618;
  assign n15620 = ~pi23  & ~n15618;
  assign n15621 = ~n15619 & ~n15620;
  assign n15622 = ~n15611 & ~n15621;
  assign n15623 = ~n15610 & ~n15622;
  assign n15624 = n15558 & ~n15623;
  assign n15625 = ~n15558 & n15623;
  assign n15626 = n5435 & n12653;
  assign n15627 = n6055 & n12650;
  assign n15628 = n5429 & n13042;
  assign n15629 = n6071 & n12647;
  assign n15630 = ~n15628 & ~n15629;
  assign n15631 = ~n15627 & n15630;
  assign n15632 = ~n15626 & n15631;
  assign n15633 = pi20  & n15632;
  assign n15634 = ~pi20  & ~n15632;
  assign n15635 = ~n15633 & ~n15634;
  assign n15636 = ~n15625 & ~n15635;
  assign n15637 = ~n15624 & ~n15636;
  assign n15638 = ~n15554 & ~n15637;
  assign n15639 = ~n15551 & ~n15638;
  assign n15640 = ~n15474 & ~n15475;
  assign n15641 = ~n15485 & n15640;
  assign n15642 = n15485 & ~n15640;
  assign n15643 = ~n15641 & ~n15642;
  assign n15644 = ~n15639 & n15643;
  assign n15645 = n15639 & ~n15643;
  assign n15646 = n6184 & n12636;
  assign n15647 = n6527 & n12633;
  assign n15648 = n6185 & n13292;
  assign n15649 = n6543 & n12630;
  assign n15650 = ~n15648 & ~n15649;
  assign n15651 = ~n15647 & n15650;
  assign n15652 = ~n15646 & n15651;
  assign n15653 = pi17  & n15652;
  assign n15654 = ~pi17  & ~n15652;
  assign n15655 = ~n15653 & ~n15654;
  assign n15656 = ~n15645 & ~n15655;
  assign n15657 = ~n15644 & ~n15656;
  assign n15658 = n15538 & ~n15657;
  assign n15659 = ~n15538 & n15657;
  assign n15660 = n6835 & n12622;
  assign n15661 = n7460 & n12614;
  assign n15662 = n6836 & ~n13310;
  assign n15663 = n7487 & n12606;
  assign n15664 = ~n15662 & ~n15663;
  assign n15665 = ~n15661 & n15664;
  assign n15666 = ~n15660 & n15665;
  assign n15667 = pi14  & n15666;
  assign n15668 = ~pi14  & ~n15666;
  assign n15669 = ~n15667 & ~n15668;
  assign n15670 = ~n15659 & ~n15669;
  assign n15671 = ~n15658 & ~n15670;
  assign n15672 = ~n15534 & ~n15671;
  assign n15673 = n14945 & n15501;
  assign n15674 = ~n15502 & ~n15673;
  assign n15675 = n15534 & ~n15671;
  assign n15676 = ~n15534 & n15671;
  assign n15677 = ~n15675 & ~n15676;
  assign n15678 = n15674 & ~n15677;
  assign n15679 = ~n15672 & ~n15678;
  assign n15680 = ~n15508 & ~n15509;
  assign n15681 = ~n15519 & n15680;
  assign n15682 = n15519 & ~n15680;
  assign n15683 = ~n15681 & ~n15682;
  assign n15684 = ~n15679 & n15683;
  assign n15685 = n15679 & n15683;
  assign n15686 = ~n15679 & ~n15683;
  assign n15687 = ~n15685 & ~n15686;
  assign n15688 = ~n15674 & n15677;
  assign n15689 = ~n15678 & ~n15688;
  assign n15690 = n7648 & ~n13499;
  assign n15691 = n7654 & ~n12611;
  assign n15692 = ~n7648 & ~n7653;
  assign n15693 = ~n15691 & ~n15692;
  assign n15694 = ~n12608 & ~n15693;
  assign n15695 = ~n15690 & ~n15694;
  assign n15696 = pi11  & n15695;
  assign n15697 = ~pi11  & ~n15695;
  assign n15698 = ~n15696 & ~n15697;
  assign n15699 = n15554 & n15637;
  assign n15700 = ~n15638 & ~n15699;
  assign n15701 = n6184 & n12639;
  assign n15702 = n6527 & n12636;
  assign n15703 = n6185 & n13396;
  assign n15704 = n6543 & n12633;
  assign n15705 = ~n15703 & ~n15704;
  assign n15706 = ~n15702 & n15705;
  assign n15707 = ~n15701 & n15706;
  assign n15708 = pi17  & n15707;
  assign n15709 = ~pi17  & ~n15707;
  assign n15710 = ~n15708 & ~n15709;
  assign n15711 = n15700 & ~n15710;
  assign n15712 = n15700 & n15710;
  assign n15713 = ~n15700 & ~n15710;
  assign n15714 = ~n15712 & ~n15713;
  assign n15715 = ~n15624 & ~n15625;
  assign n15716 = ~n15635 & n15715;
  assign n15717 = n15635 & ~n15715;
  assign n15718 = ~n15716 & ~n15717;
  assign n15719 = n15601 & ~n15603;
  assign n15720 = ~n15604 & ~n15719;
  assign n15721 = n5238 & n12668;
  assign n15722 = n71 & n12665;
  assign n15723 = n5239 & n13591;
  assign n15724 = n5326 & n12662;
  assign n15725 = ~n15723 & ~n15724;
  assign n15726 = ~n15722 & n15725;
  assign n15727 = ~n15721 & n15726;
  assign n15728 = pi23  & n15727;
  assign n15729 = ~pi23  & ~n15727;
  assign n15730 = ~n15728 & ~n15729;
  assign n15731 = n15720 & ~n15730;
  assign n15732 = n15720 & n15730;
  assign n15733 = ~n15720 & ~n15730;
  assign n15734 = ~n15732 & ~n15733;
  assign n15735 = ~n15589 & n15599;
  assign n15736 = n15589 & ~n15599;
  assign n15737 = ~n15735 & ~n15736;
  assign n15738 = n15000 & n15419;
  assign n15739 = ~n15420 & ~n15738;
  assign n15740 = n4006 & n12692;
  assign n15741 = n4133 & n12689;
  assign n15742 = n4002 & n14382;
  assign n15743 = n4555 & n12686;
  assign n15744 = ~n15742 & ~n15743;
  assign n15745 = ~n15741 & n15744;
  assign n15746 = ~n15740 & n15745;
  assign n15747 = pi29  & n15746;
  assign n15748 = ~pi29  & ~n15746;
  assign n15749 = ~n15747 & ~n15748;
  assign n15750 = n15739 & ~n15749;
  assign n15751 = n15739 & n15749;
  assign n15752 = ~n15739 & ~n15749;
  assign n15753 = ~n15751 & ~n15752;
  assign n15754 = n4801 & n12677;
  assign n15755 = n4601 & n12683;
  assign n15756 = n4602 & n13929;
  assign n15757 = n4783 & n12680;
  assign n15758 = ~n15756 & ~n15757;
  assign n15759 = ~n15755 & n15758;
  assign n15760 = ~n15754 & n15759;
  assign n15761 = pi26  & n15760;
  assign n15762 = ~pi26  & ~n15760;
  assign n15763 = ~n15761 & ~n15762;
  assign n15764 = ~n15753 & ~n15763;
  assign n15765 = ~n15750 & ~n15764;
  assign n15766 = ~n15737 & ~n15765;
  assign n15767 = n15737 & n15765;
  assign n15768 = n5238 & n12671;
  assign n15769 = n71 & n12668;
  assign n15770 = n5239 & n13578;
  assign n15771 = n5326 & n12665;
  assign n15772 = ~n15770 & ~n15771;
  assign n15773 = ~n15769 & n15772;
  assign n15774 = ~n15768 & n15773;
  assign n15775 = pi23  & n15774;
  assign n15776 = ~pi23  & ~n15774;
  assign n15777 = ~n15775 & ~n15776;
  assign n15778 = ~n15767 & ~n15777;
  assign n15779 = ~n15766 & ~n15778;
  assign n15780 = ~n15734 & ~n15779;
  assign n15781 = ~n15731 & ~n15780;
  assign n15782 = ~n15610 & ~n15611;
  assign n15783 = ~n15621 & n15782;
  assign n15784 = n15621 & ~n15782;
  assign n15785 = ~n15783 & ~n15784;
  assign n15786 = ~n15781 & n15785;
  assign n15787 = n15781 & ~n15785;
  assign n15788 = n5435 & n12656;
  assign n15789 = n6055 & n12653;
  assign n15790 = n5429 & n12991;
  assign n15791 = n6071 & n12650;
  assign n15792 = ~n15790 & ~n15791;
  assign n15793 = ~n15789 & n15792;
  assign n15794 = ~n15788 & n15793;
  assign n15795 = pi20  & n15794;
  assign n15796 = ~pi20  & ~n15794;
  assign n15797 = ~n15795 & ~n15796;
  assign n15798 = ~n15787 & ~n15797;
  assign n15799 = ~n15786 & ~n15798;
  assign n15800 = n15718 & ~n15799;
  assign n15801 = ~n15718 & n15799;
  assign n15802 = n6184 & n12644;
  assign n15803 = n6527 & n12639;
  assign n15804 = n6185 & n13210;
  assign n15805 = n6543 & n12636;
  assign n15806 = ~n15804 & ~n15805;
  assign n15807 = ~n15803 & n15806;
  assign n15808 = ~n15802 & n15807;
  assign n15809 = pi17  & n15808;
  assign n15810 = ~pi17  & ~n15808;
  assign n15811 = ~n15809 & ~n15810;
  assign n15812 = ~n15801 & ~n15811;
  assign n15813 = ~n15800 & ~n15812;
  assign n15814 = ~n15714 & ~n15813;
  assign n15815 = ~n15711 & ~n15814;
  assign n15816 = ~n15644 & ~n15645;
  assign n15817 = ~n15655 & n15816;
  assign n15818 = n15655 & ~n15816;
  assign n15819 = ~n15817 & ~n15818;
  assign n15820 = ~n15815 & n15819;
  assign n15821 = n15815 & ~n15819;
  assign n15822 = n6835 & n12625;
  assign n15823 = n7460 & n12622;
  assign n15824 = n6836 & n13463;
  assign n15825 = n7487 & n12614;
  assign n15826 = ~n15824 & ~n15825;
  assign n15827 = ~n15823 & n15826;
  assign n15828 = ~n15822 & n15827;
  assign n15829 = pi14  & n15828;
  assign n15830 = ~pi14  & ~n15828;
  assign n15831 = ~n15829 & ~n15830;
  assign n15832 = ~n15821 & ~n15831;
  assign n15833 = ~n15820 & ~n15832;
  assign n15834 = ~n15698 & ~n15833;
  assign n15835 = n15698 & n15833;
  assign n15836 = ~n15658 & ~n15659;
  assign n15837 = ~n15669 & n15836;
  assign n15838 = n15669 & ~n15836;
  assign n15839 = ~n15837 & ~n15838;
  assign n15840 = ~n15835 & n15839;
  assign n15841 = ~n15834 & ~n15840;
  assign n15842 = n15689 & ~n15841;
  assign n15843 = ~n15834 & ~n15835;
  assign n15844 = n15839 & n15843;
  assign n15845 = ~n15839 & ~n15843;
  assign n15846 = ~n15844 & ~n15845;
  assign n15847 = n15714 & n15813;
  assign n15848 = ~n15814 & ~n15847;
  assign n15849 = n6835 & n12630;
  assign n15850 = n7460 & n12625;
  assign n15851 = n6836 & n13325;
  assign n15852 = n7487 & n12622;
  assign n15853 = ~n15851 & ~n15852;
  assign n15854 = ~n15850 & n15853;
  assign n15855 = ~n15849 & n15854;
  assign n15856 = pi14  & n15855;
  assign n15857 = ~pi14  & ~n15855;
  assign n15858 = ~n15856 & ~n15857;
  assign n15859 = n15848 & ~n15858;
  assign n15860 = n15848 & n15858;
  assign n15861 = ~n15848 & ~n15858;
  assign n15862 = ~n15860 & ~n15861;
  assign n15863 = ~n15800 & ~n15801;
  assign n15864 = ~n15811 & n15863;
  assign n15865 = n15811 & ~n15863;
  assign n15866 = ~n15864 & ~n15865;
  assign n15867 = n15734 & n15779;
  assign n15868 = ~n15780 & ~n15867;
  assign n15869 = n5435 & n12659;
  assign n15870 = n6055 & n12656;
  assign n15871 = n5429 & n13059;
  assign n15872 = n6071 & n12653;
  assign n15873 = ~n15871 & ~n15872;
  assign n15874 = ~n15870 & n15873;
  assign n15875 = ~n15869 & n15874;
  assign n15876 = pi20  & n15875;
  assign n15877 = ~pi20  & ~n15875;
  assign n15878 = ~n15876 & ~n15877;
  assign n15879 = n15868 & ~n15878;
  assign n15880 = n15868 & n15878;
  assign n15881 = ~n15868 & ~n15878;
  assign n15882 = ~n15880 & ~n15881;
  assign n15883 = ~n15766 & ~n15767;
  assign n15884 = ~n15777 & n15883;
  assign n15885 = n15777 & ~n15883;
  assign n15886 = ~n15884 & ~n15885;
  assign n15887 = ~n15753 & n15763;
  assign n15888 = n15753 & ~n15763;
  assign n15889 = ~n15887 & ~n15888;
  assign n15890 = n4006 & n12698;
  assign n15891 = n4133 & n12695;
  assign n15892 = n4002 & n14976;
  assign n15893 = n4555 & n12692;
  assign n15894 = ~n15892 & ~n15893;
  assign n15895 = ~n15891 & n15894;
  assign n15896 = ~n15890 & n15895;
  assign n15897 = pi29  & n15896;
  assign n15898 = ~pi29  & ~n15896;
  assign n15899 = ~n15897 & ~n15898;
  assign n15900 = n15395 & n15398;
  assign n15901 = ~n15399 & ~n15900;
  assign n15902 = ~n15899 & n15901;
  assign n15903 = n4006 & n12701;
  assign n15904 = n4133 & n12698;
  assign n15905 = n4002 & n14991;
  assign n15906 = n4555 & n12695;
  assign n15907 = ~n15905 & ~n15906;
  assign n15908 = ~n15904 & n15907;
  assign n15909 = ~n15903 & n15908;
  assign n15910 = pi29  & n15909;
  assign n15911 = ~pi29  & ~n15909;
  assign n15912 = ~n15910 & ~n15911;
  assign n15913 = n15390 & n15393;
  assign n15914 = ~n15394 & ~n15913;
  assign n15915 = ~n15912 & n15914;
  assign n15916 = n4006 & n12704;
  assign n15917 = n4133 & n12701;
  assign n15918 = n4002 & n14655;
  assign n15919 = n4555 & n12698;
  assign n15920 = ~n15918 & ~n15919;
  assign n15921 = ~n15917 & n15920;
  assign n15922 = ~n15916 & n15921;
  assign n15923 = pi29  & n15922;
  assign n15924 = ~pi29  & ~n15922;
  assign n15925 = ~n15923 & ~n15924;
  assign n15926 = n15385 & n15388;
  assign n15927 = ~n15389 & ~n15926;
  assign n15928 = ~n15925 & n15927;
  assign n15929 = n4006 & n12707;
  assign n15930 = n4133 & n12704;
  assign n15931 = n4002 & n15024;
  assign n15932 = n4555 & n12701;
  assign n15933 = ~n15931 & ~n15932;
  assign n15934 = ~n15930 & n15933;
  assign n15935 = ~n15929 & n15934;
  assign n15936 = pi29  & n15935;
  assign n15937 = ~pi29  & ~n15935;
  assign n15938 = ~n15936 & ~n15937;
  assign n15939 = n15380 & n15383;
  assign n15940 = ~n15384 & ~n15939;
  assign n15941 = ~n15938 & n15940;
  assign n15942 = n4006 & n12710;
  assign n15943 = n4133 & n12707;
  assign n15944 = n4002 & n15050;
  assign n15945 = n4555 & n12704;
  assign n15946 = ~n15944 & ~n15945;
  assign n15947 = ~n15943 & n15946;
  assign n15948 = ~n15942 & n15947;
  assign n15949 = pi29  & n15948;
  assign n15950 = ~pi29  & ~n15948;
  assign n15951 = ~n15949 & ~n15950;
  assign n15952 = n15375 & n15378;
  assign n15953 = ~n15379 & ~n15952;
  assign n15954 = ~n15951 & n15953;
  assign n15955 = n4006 & n12713;
  assign n15956 = n4133 & n12710;
  assign n15957 = n4002 & n15074;
  assign n15958 = n4555 & n12707;
  assign n15959 = ~n15957 & ~n15958;
  assign n15960 = ~n15956 & n15959;
  assign n15961 = ~n15955 & n15960;
  assign n15962 = ~pi29  & ~n15961;
  assign n15963 = pi29  & n15961;
  assign n15964 = ~n15962 & ~n15963;
  assign n15965 = n15370 & n15373;
  assign n15966 = ~n15374 & ~n15965;
  assign n15967 = ~n15964 & n15966;
  assign n15968 = ~n15964 & ~n15966;
  assign n15969 = n15964 & n15966;
  assign n15970 = ~n15968 & ~n15969;
  assign n15971 = n4006 & n12716;
  assign n15972 = n4133 & n12713;
  assign n15973 = n4002 & n15105;
  assign n15974 = n4555 & n12710;
  assign n15975 = ~n15973 & ~n15974;
  assign n15976 = ~n15972 & n15975;
  assign n15977 = ~n15971 & n15976;
  assign n15978 = ~pi29  & ~n15977;
  assign n15979 = pi29  & n15977;
  assign n15980 = ~n15978 & ~n15979;
  assign n15981 = n15365 & n15368;
  assign n15982 = ~n15369 & ~n15981;
  assign n15983 = ~n15980 & n15982;
  assign n15984 = ~n15980 & ~n15982;
  assign n15985 = n15980 & n15982;
  assign n15986 = ~n15984 & ~n15985;
  assign n15987 = n4006 & n12719;
  assign n15988 = n4133 & n12716;
  assign n15989 = n4002 & n15161;
  assign n15990 = n4555 & n12713;
  assign n15991 = ~n15989 & ~n15990;
  assign n15992 = ~n15988 & n15991;
  assign n15993 = ~n15987 & n15992;
  assign n15994 = ~pi29  & ~n15993;
  assign n15995 = pi29  & n15993;
  assign n15996 = ~n15994 & ~n15995;
  assign n15997 = n15277 & n15363;
  assign n15998 = ~n15364 & ~n15997;
  assign n15999 = ~n15996 & n15998;
  assign n16000 = ~n15996 & ~n15998;
  assign n16001 = n15996 & n15998;
  assign n16002 = ~n16000 & ~n16001;
  assign n16003 = n4006 & n12722;
  assign n16004 = n4133 & n12719;
  assign n16005 = n4002 & n15199;
  assign n16006 = n4555 & n12716;
  assign n16007 = ~n16005 & ~n16006;
  assign n16008 = ~n16004 & n16007;
  assign n16009 = ~n16003 & n16008;
  assign n16010 = ~pi29  & ~n16009;
  assign n16011 = pi29  & n16009;
  assign n16012 = ~n16010 & ~n16011;
  assign n16013 = ~n15350 & ~n15351;
  assign n16014 = ~n15361 & n16013;
  assign n16015 = n15361 & ~n16013;
  assign n16016 = ~n16014 & ~n16015;
  assign n16017 = ~n16012 & n16016;
  assign n16018 = n4006 & n12725;
  assign n16019 = n4133 & n12722;
  assign n16020 = n4002 & n15243;
  assign n16021 = n4555 & n12719;
  assign n16022 = ~n16020 & ~n16021;
  assign n16023 = ~n16019 & n16022;
  assign n16024 = ~n16018 & n16023;
  assign n16025 = ~pi29  & ~n16024;
  assign n16026 = pi29  & n16024;
  assign n16027 = ~n16025 & ~n16026;
  assign n16028 = ~n15309 & n15317;
  assign n16029 = n15309 & ~n15317;
  assign n16030 = ~n16028 & ~n16029;
  assign n16031 = ~n16027 & ~n16030;
  assign n16032 = ~n555 & n12732;
  assign n16033 = n4002 & ~n15312;
  assign n16034 = n4555 & n12730;
  assign n16035 = n4133 & n12732;
  assign n16036 = ~n16034 & ~n16035;
  assign n16037 = ~n16033 & n16036;
  assign n16038 = ~n3998 & n12732;
  assign n16039 = pi29  & ~n16038;
  assign n16040 = n16037 & n16039;
  assign n16041 = n4006 & n12732;
  assign n16042 = n4133 & n12730;
  assign n16043 = n4002 & ~n15356;
  assign n16044 = n4555 & n12725;
  assign n16045 = ~n16043 & ~n16044;
  assign n16046 = ~n16042 & n16045;
  assign n16047 = ~n16041 & n16046;
  assign n16048 = n16040 & n16047;
  assign n16049 = n16032 & n16048;
  assign n16050 = n4006 & n12730;
  assign n16051 = n4133 & n12725;
  assign n16052 = n4002 & n15267;
  assign n16053 = n4555 & n12722;
  assign n16054 = ~n16052 & ~n16053;
  assign n16055 = ~n16051 & n16054;
  assign n16056 = ~n16050 & n16055;
  assign n16057 = ~pi29  & ~n16056;
  assign n16058 = pi29  & n16056;
  assign n16059 = ~n16057 & ~n16058;
  assign n16060 = ~n16032 & n16048;
  assign n16061 = n16032 & ~n16048;
  assign n16062 = ~n16060 & ~n16061;
  assign n16063 = ~n16059 & ~n16062;
  assign n16064 = ~n16049 & ~n16063;
  assign n16065 = n16027 & n16030;
  assign n16066 = ~n16031 & ~n16065;
  assign n16067 = ~n16064 & n16066;
  assign n16068 = ~n16031 & ~n16067;
  assign n16069 = n16012 & ~n16016;
  assign n16070 = ~n16017 & ~n16069;
  assign n16071 = ~n16068 & n16070;
  assign n16072 = ~n16017 & ~n16071;
  assign n16073 = ~n16002 & ~n16072;
  assign n16074 = ~n15999 & ~n16073;
  assign n16075 = ~n15986 & ~n16074;
  assign n16076 = ~n15983 & ~n16075;
  assign n16077 = ~n15970 & ~n16076;
  assign n16078 = ~n15967 & ~n16077;
  assign n16079 = n15951 & ~n15953;
  assign n16080 = ~n15954 & ~n16079;
  assign n16081 = ~n16078 & n16080;
  assign n16082 = ~n15954 & ~n16081;
  assign n16083 = n15938 & ~n15940;
  assign n16084 = ~n15941 & ~n16083;
  assign n16085 = ~n16082 & n16084;
  assign n16086 = ~n15941 & ~n16085;
  assign n16087 = n15925 & ~n15927;
  assign n16088 = ~n15928 & ~n16087;
  assign n16089 = ~n16086 & n16088;
  assign n16090 = ~n15928 & ~n16089;
  assign n16091 = n15912 & ~n15914;
  assign n16092 = ~n15915 & ~n16091;
  assign n16093 = ~n16090 & n16092;
  assign n16094 = ~n15915 & ~n16093;
  assign n16095 = n15899 & ~n15901;
  assign n16096 = ~n15902 & ~n16095;
  assign n16097 = ~n16094 & n16096;
  assign n16098 = ~n15902 & ~n16097;
  assign n16099 = ~n15407 & n15417;
  assign n16100 = ~n15418 & ~n16099;
  assign n16101 = ~n16098 & n16100;
  assign n16102 = n16098 & ~n16100;
  assign n16103 = n4601 & n12686;
  assign n16104 = n4783 & n12683;
  assign n16105 = n4602 & n14402;
  assign n16106 = n4801 & n12680;
  assign n16107 = ~n16105 & ~n16106;
  assign n16108 = ~n16104 & n16107;
  assign n16109 = ~n16103 & n16108;
  assign n16110 = pi26  & n16109;
  assign n16111 = ~pi26  & ~n16109;
  assign n16112 = ~n16110 & ~n16111;
  assign n16113 = ~n16102 & ~n16112;
  assign n16114 = ~n16101 & ~n16113;
  assign n16115 = ~n15889 & ~n16114;
  assign n16116 = n15889 & n16114;
  assign n16117 = n5238 & n12674;
  assign n16118 = n71 & n12671;
  assign n16119 = n5239 & n13764;
  assign n16120 = n5326 & n12668;
  assign n16121 = ~n16119 & ~n16120;
  assign n16122 = ~n16118 & n16121;
  assign n16123 = ~n16117 & n16122;
  assign n16124 = pi23  & n16123;
  assign n16125 = ~pi23  & ~n16123;
  assign n16126 = ~n16124 & ~n16125;
  assign n16127 = ~n16116 & ~n16126;
  assign n16128 = ~n16115 & ~n16127;
  assign n16129 = n15886 & ~n16128;
  assign n16130 = ~n15886 & n16128;
  assign n16131 = n5435 & n12662;
  assign n16132 = n6055 & n12659;
  assign n16133 = n5429 & n13246;
  assign n16134 = n6071 & n12656;
  assign n16135 = ~n16133 & ~n16134;
  assign n16136 = ~n16132 & n16135;
  assign n16137 = ~n16131 & n16136;
  assign n16138 = pi20  & n16137;
  assign n16139 = ~pi20  & ~n16137;
  assign n16140 = ~n16138 & ~n16139;
  assign n16141 = ~n16130 & ~n16140;
  assign n16142 = ~n16129 & ~n16141;
  assign n16143 = ~n15882 & ~n16142;
  assign n16144 = ~n15879 & ~n16143;
  assign n16145 = ~n15786 & ~n15787;
  assign n16146 = ~n15797 & n16145;
  assign n16147 = n15797 & ~n16145;
  assign n16148 = ~n16146 & ~n16147;
  assign n16149 = ~n16144 & n16148;
  assign n16150 = n16144 & ~n16148;
  assign n16151 = n6184 & n12647;
  assign n16152 = n6527 & n12644;
  assign n16153 = n6185 & ~n13193;
  assign n16154 = n6543 & n12639;
  assign n16155 = ~n16153 & ~n16154;
  assign n16156 = ~n16152 & n16155;
  assign n16157 = ~n16151 & n16156;
  assign n16158 = pi17  & n16157;
  assign n16159 = ~pi17  & ~n16157;
  assign n16160 = ~n16158 & ~n16159;
  assign n16161 = ~n16150 & ~n16160;
  assign n16162 = ~n16149 & ~n16161;
  assign n16163 = n15866 & ~n16162;
  assign n16164 = ~n15866 & n16162;
  assign n16165 = n6835 & n12633;
  assign n16166 = n7460 & n12630;
  assign n16167 = n6836 & ~n13227;
  assign n16168 = n7487 & n12625;
  assign n16169 = ~n16167 & ~n16168;
  assign n16170 = ~n16166 & n16169;
  assign n16171 = ~n16165 & n16170;
  assign n16172 = pi14  & n16171;
  assign n16173 = ~pi14  & ~n16171;
  assign n16174 = ~n16172 & ~n16173;
  assign n16175 = ~n16164 & ~n16174;
  assign n16176 = ~n16163 & ~n16175;
  assign n16177 = ~n15862 & ~n16176;
  assign n16178 = ~n15859 & ~n16177;
  assign n16179 = ~n15820 & ~n15821;
  assign n16180 = ~n15831 & n16179;
  assign n16181 = n15831 & ~n16179;
  assign n16182 = ~n16180 & ~n16181;
  assign n16183 = ~n16178 & n16182;
  assign n16184 = n16178 & ~n16182;
  assign n16185 = n7654 & n12606;
  assign n16186 = n8091 & n12616;
  assign n16187 = n7648 & ~n13483;
  assign n16188 = n8120 & ~n12608;
  assign n16189 = ~n16187 & ~n16188;
  assign n16190 = ~n16186 & n16189;
  assign n16191 = ~n16185 & n16190;
  assign n16192 = pi11  & n16191;
  assign n16193 = ~pi11  & ~n16191;
  assign n16194 = ~n16192 & ~n16193;
  assign n16195 = ~n16184 & ~n16194;
  assign n16196 = ~n16183 & ~n16195;
  assign n16197 = n15846 & ~n16196;
  assign n16198 = ~n15846 & n16196;
  assign n16199 = ~n16197 & ~n16198;
  assign n16200 = n8091 & n12606;
  assign n16201 = ~n12611 & n16188;
  assign n16202 = n7654 & n12614;
  assign n16203 = n7648 & n12868;
  assign n16204 = ~n16202 & ~n16203;
  assign n16205 = ~n16201 & n16204;
  assign n16206 = ~n16200 & n16205;
  assign n16207 = pi11  & n16206;
  assign n16208 = ~pi11  & ~n16206;
  assign n16209 = ~n16207 & ~n16208;
  assign n16210 = ~n16163 & ~n16164;
  assign n16211 = ~n16174 & n16210;
  assign n16212 = n16174 & ~n16210;
  assign n16213 = ~n16211 & ~n16212;
  assign n16214 = n15882 & n16142;
  assign n16215 = ~n16143 & ~n16214;
  assign n16216 = n6184 & n12650;
  assign n16217 = n6527 & n12647;
  assign n16218 = n6185 & n13275;
  assign n16219 = n6543 & n12644;
  assign n16220 = ~n16218 & ~n16219;
  assign n16221 = ~n16217 & n16220;
  assign n16222 = ~n16216 & n16221;
  assign n16223 = pi17  & n16222;
  assign n16224 = ~pi17  & ~n16222;
  assign n16225 = ~n16223 & ~n16224;
  assign n16226 = n16215 & ~n16225;
  assign n16227 = n16215 & n16225;
  assign n16228 = ~n16215 & ~n16225;
  assign n16229 = ~n16227 & ~n16228;
  assign n16230 = ~n16129 & ~n16130;
  assign n16231 = ~n16140 & n16230;
  assign n16232 = n16140 & ~n16230;
  assign n16233 = ~n16231 & ~n16232;
  assign n16234 = ~n16115 & ~n16116;
  assign n16235 = ~n16126 & n16234;
  assign n16236 = n16126 & ~n16234;
  assign n16237 = ~n16235 & ~n16236;
  assign n16238 = n16094 & ~n16096;
  assign n16239 = ~n16097 & ~n16238;
  assign n16240 = n4601 & n12689;
  assign n16241 = n4783 & n12686;
  assign n16242 = n4602 & n14552;
  assign n16243 = n4801 & n12683;
  assign n16244 = ~n16242 & ~n16243;
  assign n16245 = ~n16241 & n16244;
  assign n16246 = ~n16240 & n16245;
  assign n16247 = pi26  & n16246;
  assign n16248 = ~pi26  & ~n16246;
  assign n16249 = ~n16247 & ~n16248;
  assign n16250 = n16239 & ~n16249;
  assign n16251 = n16090 & ~n16092;
  assign n16252 = ~n16093 & ~n16251;
  assign n16253 = n4601 & n12692;
  assign n16254 = n4783 & n12689;
  assign n16255 = n4602 & n14382;
  assign n16256 = n4801 & n12686;
  assign n16257 = ~n16255 & ~n16256;
  assign n16258 = ~n16254 & n16257;
  assign n16259 = ~n16253 & n16258;
  assign n16260 = pi26  & n16259;
  assign n16261 = ~pi26  & ~n16259;
  assign n16262 = ~n16260 & ~n16261;
  assign n16263 = n16252 & ~n16262;
  assign n16264 = n16086 & ~n16088;
  assign n16265 = ~n16089 & ~n16264;
  assign n16266 = n4601 & n12695;
  assign n16267 = n4783 & n12692;
  assign n16268 = n4602 & n14677;
  assign n16269 = n4801 & n12689;
  assign n16270 = ~n16268 & ~n16269;
  assign n16271 = ~n16267 & n16270;
  assign n16272 = ~n16266 & n16271;
  assign n16273 = pi26  & n16272;
  assign n16274 = ~pi26  & ~n16272;
  assign n16275 = ~n16273 & ~n16274;
  assign n16276 = n16265 & ~n16275;
  assign n16277 = n16082 & ~n16084;
  assign n16278 = ~n16085 & ~n16277;
  assign n16279 = n4601 & n12698;
  assign n16280 = n4783 & n12695;
  assign n16281 = n4602 & n14976;
  assign n16282 = n4801 & n12692;
  assign n16283 = ~n16281 & ~n16282;
  assign n16284 = ~n16280 & n16283;
  assign n16285 = ~n16279 & n16284;
  assign n16286 = pi26  & n16285;
  assign n16287 = ~pi26  & ~n16285;
  assign n16288 = ~n16286 & ~n16287;
  assign n16289 = n16278 & ~n16288;
  assign n16290 = n16078 & ~n16080;
  assign n16291 = ~n16081 & ~n16290;
  assign n16292 = n4601 & n12701;
  assign n16293 = n4783 & n12698;
  assign n16294 = n4602 & n14991;
  assign n16295 = n4801 & n12695;
  assign n16296 = ~n16294 & ~n16295;
  assign n16297 = ~n16293 & n16296;
  assign n16298 = ~n16292 & n16297;
  assign n16299 = pi26  & n16298;
  assign n16300 = ~pi26  & ~n16298;
  assign n16301 = ~n16299 & ~n16300;
  assign n16302 = n16291 & ~n16301;
  assign n16303 = n15970 & n16076;
  assign n16304 = ~n16077 & ~n16303;
  assign n16305 = n4601 & n12704;
  assign n16306 = n4783 & n12701;
  assign n16307 = n4602 & n14655;
  assign n16308 = n4801 & n12698;
  assign n16309 = ~n16307 & ~n16308;
  assign n16310 = ~n16306 & n16309;
  assign n16311 = ~n16305 & n16310;
  assign n16312 = pi26  & n16311;
  assign n16313 = ~pi26  & ~n16311;
  assign n16314 = ~n16312 & ~n16313;
  assign n16315 = n16304 & ~n16314;
  assign n16316 = n15986 & n16074;
  assign n16317 = ~n16075 & ~n16316;
  assign n16318 = n4783 & n12704;
  assign n16319 = n4801 & n12701;
  assign n16320 = n4602 & n15024;
  assign n16321 = n4601 & n12707;
  assign n16322 = ~n16320 & ~n16321;
  assign n16323 = ~n16319 & n16322;
  assign n16324 = ~n16318 & n16323;
  assign n16325 = pi26  & n16324;
  assign n16326 = ~pi26  & ~n16324;
  assign n16327 = ~n16325 & ~n16326;
  assign n16328 = n16317 & ~n16327;
  assign n16329 = n16002 & n16072;
  assign n16330 = ~n16073 & ~n16329;
  assign n16331 = n4801 & n12704;
  assign n16332 = n4783 & n12707;
  assign n16333 = n4602 & n15050;
  assign n16334 = n4601 & n12710;
  assign n16335 = ~n16333 & ~n16334;
  assign n16336 = ~n16332 & n16335;
  assign n16337 = ~n16331 & n16336;
  assign n16338 = pi26  & n16337;
  assign n16339 = ~pi26  & ~n16337;
  assign n16340 = ~n16338 & ~n16339;
  assign n16341 = n16330 & ~n16340;
  assign n16342 = n16068 & ~n16070;
  assign n16343 = ~n16071 & ~n16342;
  assign n16344 = n4801 & n12707;
  assign n16345 = n4601 & n12713;
  assign n16346 = n4602 & n15074;
  assign n16347 = n4783 & n12710;
  assign n16348 = ~n16346 & ~n16347;
  assign n16349 = ~n16345 & n16348;
  assign n16350 = ~n16344 & n16349;
  assign n16351 = pi26  & n16350;
  assign n16352 = ~pi26  & ~n16350;
  assign n16353 = ~n16351 & ~n16352;
  assign n16354 = n16343 & ~n16353;
  assign n16355 = n4783 & n12713;
  assign n16356 = n4801 & n12710;
  assign n16357 = n4602 & n15105;
  assign n16358 = n4601 & n12716;
  assign n16359 = ~n16357 & ~n16358;
  assign n16360 = ~n16356 & n16359;
  assign n16361 = ~n16355 & n16360;
  assign n16362 = pi26  & n16361;
  assign n16363 = ~pi26  & ~n16361;
  assign n16364 = ~n16362 & ~n16363;
  assign n16365 = n16064 & ~n16066;
  assign n16366 = ~n16067 & ~n16365;
  assign n16367 = ~n16364 & n16366;
  assign n16368 = n4801 & n12713;
  assign n16369 = n4601 & n12719;
  assign n16370 = n4602 & n15161;
  assign n16371 = n4783 & n12716;
  assign n16372 = ~n16370 & ~n16371;
  assign n16373 = ~n16369 & n16372;
  assign n16374 = ~n16368 & n16373;
  assign n16375 = ~pi26  & ~n16374;
  assign n16376 = pi26  & n16374;
  assign n16377 = ~n16375 & ~n16376;
  assign n16378 = n16059 & n16062;
  assign n16379 = ~n16063 & ~n16378;
  assign n16380 = ~n16377 & n16379;
  assign n16381 = ~n16377 & ~n16379;
  assign n16382 = n16377 & n16379;
  assign n16383 = ~n16381 & ~n16382;
  assign n16384 = n4783 & n12719;
  assign n16385 = n4801 & n12716;
  assign n16386 = n4602 & n15199;
  assign n16387 = n4601 & n12722;
  assign n16388 = ~n16386 & ~n16387;
  assign n16389 = ~n16385 & n16388;
  assign n16390 = ~n16384 & n16389;
  assign n16391 = ~pi26  & ~n16390;
  assign n16392 = pi26  & n16390;
  assign n16393 = ~n16391 & ~n16392;
  assign n16394 = pi29  & ~n16040;
  assign n16395 = n16047 & ~n16394;
  assign n16396 = ~n16047 & n16394;
  assign n16397 = ~n16395 & ~n16396;
  assign n16398 = ~n16393 & n16397;
  assign n16399 = ~n16393 & ~n16397;
  assign n16400 = n16393 & n16397;
  assign n16401 = ~n16399 & ~n16400;
  assign n16402 = n4801 & n12719;
  assign n16403 = n4783 & n12722;
  assign n16404 = n4602 & n15243;
  assign n16405 = n4601 & n12725;
  assign n16406 = ~n16404 & ~n16405;
  assign n16407 = ~n16403 & n16406;
  assign n16408 = ~n16402 & n16407;
  assign n16409 = pi26  & n16408;
  assign n16410 = ~pi26  & ~n16408;
  assign n16411 = ~n16409 & ~n16410;
  assign n16412 = pi29  & n16038;
  assign n16413 = ~n16037 & n16412;
  assign n16414 = n16037 & ~n16412;
  assign n16415 = ~n16413 & ~n16414;
  assign n16416 = ~n16411 & n16415;
  assign n16417 = n4602 & ~n15312;
  assign n16418 = n4783 & n12732;
  assign n16419 = n4801 & n12730;
  assign n16420 = ~n16418 & ~n16419;
  assign n16421 = ~n16417 & n16420;
  assign n16422 = ~n4598 & n12732;
  assign n16423 = pi26  & ~n16422;
  assign n16424 = n16421 & n16423;
  assign n16425 = n4801 & n12725;
  assign n16426 = n4783 & n12730;
  assign n16427 = n4602 & ~n15356;
  assign n16428 = n4601 & n12732;
  assign n16429 = ~n16427 & ~n16428;
  assign n16430 = ~n16426 & n16429;
  assign n16431 = ~n16425 & n16430;
  assign n16432 = n16424 & n16431;
  assign n16433 = n16038 & n16432;
  assign n16434 = ~n16038 & n16432;
  assign n16435 = n16038 & ~n16432;
  assign n16436 = ~n16434 & ~n16435;
  assign n16437 = n4801 & n12722;
  assign n16438 = n4783 & n12725;
  assign n16439 = n4602 & n15267;
  assign n16440 = n4601 & n12730;
  assign n16441 = ~n16439 & ~n16440;
  assign n16442 = ~n16438 & n16441;
  assign n16443 = ~n16437 & n16442;
  assign n16444 = pi26  & n16443;
  assign n16445 = ~pi26  & ~n16443;
  assign n16446 = ~n16444 & ~n16445;
  assign n16447 = ~n16436 & ~n16446;
  assign n16448 = ~n16433 & ~n16447;
  assign n16449 = n16411 & ~n16415;
  assign n16450 = ~n16416 & ~n16449;
  assign n16451 = ~n16448 & n16450;
  assign n16452 = ~n16416 & ~n16451;
  assign n16453 = ~n16401 & ~n16452;
  assign n16454 = ~n16398 & ~n16453;
  assign n16455 = ~n16383 & ~n16454;
  assign n16456 = ~n16380 & ~n16455;
  assign n16457 = n16364 & n16366;
  assign n16458 = ~n16364 & ~n16366;
  assign n16459 = ~n16457 & ~n16458;
  assign n16460 = ~n16456 & ~n16459;
  assign n16461 = ~n16367 & ~n16460;
  assign n16462 = n16343 & n16353;
  assign n16463 = ~n16343 & ~n16353;
  assign n16464 = ~n16462 & ~n16463;
  assign n16465 = ~n16461 & ~n16464;
  assign n16466 = ~n16354 & ~n16465;
  assign n16467 = n16330 & n16340;
  assign n16468 = ~n16330 & ~n16340;
  assign n16469 = ~n16467 & ~n16468;
  assign n16470 = ~n16466 & ~n16469;
  assign n16471 = ~n16341 & ~n16470;
  assign n16472 = n16317 & n16327;
  assign n16473 = ~n16317 & ~n16327;
  assign n16474 = ~n16472 & ~n16473;
  assign n16475 = ~n16471 & ~n16474;
  assign n16476 = ~n16328 & ~n16475;
  assign n16477 = n16304 & n16314;
  assign n16478 = ~n16304 & ~n16314;
  assign n16479 = ~n16477 & ~n16478;
  assign n16480 = ~n16476 & ~n16479;
  assign n16481 = ~n16315 & ~n16480;
  assign n16482 = n16291 & n16301;
  assign n16483 = ~n16291 & ~n16301;
  assign n16484 = ~n16482 & ~n16483;
  assign n16485 = ~n16481 & ~n16484;
  assign n16486 = ~n16302 & ~n16485;
  assign n16487 = n16278 & n16288;
  assign n16488 = ~n16278 & ~n16288;
  assign n16489 = ~n16487 & ~n16488;
  assign n16490 = ~n16486 & ~n16489;
  assign n16491 = ~n16289 & ~n16490;
  assign n16492 = n16265 & n16275;
  assign n16493 = ~n16265 & ~n16275;
  assign n16494 = ~n16492 & ~n16493;
  assign n16495 = ~n16491 & ~n16494;
  assign n16496 = ~n16276 & ~n16495;
  assign n16497 = n16252 & n16262;
  assign n16498 = ~n16252 & ~n16262;
  assign n16499 = ~n16497 & ~n16498;
  assign n16500 = ~n16496 & ~n16499;
  assign n16501 = ~n16263 & ~n16500;
  assign n16502 = ~n16239 & n16249;
  assign n16503 = ~n16250 & ~n16502;
  assign n16504 = ~n16501 & n16503;
  assign n16505 = ~n16250 & ~n16504;
  assign n16506 = ~n16101 & ~n16102;
  assign n16507 = ~n16112 & n16506;
  assign n16508 = n16112 & ~n16506;
  assign n16509 = ~n16507 & ~n16508;
  assign n16510 = ~n16505 & n16509;
  assign n16511 = n16505 & ~n16509;
  assign n16512 = n5238 & n12677;
  assign n16513 = n71 & n12674;
  assign n16514 = n5239 & n13785;
  assign n16515 = n5326 & n12671;
  assign n16516 = ~n16514 & ~n16515;
  assign n16517 = ~n16513 & n16516;
  assign n16518 = ~n16512 & n16517;
  assign n16519 = pi23  & n16518;
  assign n16520 = ~pi23  & ~n16518;
  assign n16521 = ~n16519 & ~n16520;
  assign n16522 = ~n16511 & ~n16521;
  assign n16523 = ~n16510 & ~n16522;
  assign n16524 = n16237 & ~n16523;
  assign n16525 = ~n16237 & n16523;
  assign n16526 = n5435 & n12665;
  assign n16527 = n6055 & n12662;
  assign n16528 = n5429 & n13165;
  assign n16529 = n6071 & n12659;
  assign n16530 = ~n16528 & ~n16529;
  assign n16531 = ~n16527 & n16530;
  assign n16532 = ~n16526 & n16531;
  assign n16533 = pi20  & n16532;
  assign n16534 = ~pi20  & ~n16532;
  assign n16535 = ~n16533 & ~n16534;
  assign n16536 = ~n16525 & ~n16535;
  assign n16537 = ~n16524 & ~n16536;
  assign n16538 = n16233 & ~n16537;
  assign n16539 = ~n16233 & n16537;
  assign n16540 = n6184 & n12653;
  assign n16541 = n6527 & n12650;
  assign n16542 = n6185 & n13042;
  assign n16543 = n6543 & n12647;
  assign n16544 = ~n16542 & ~n16543;
  assign n16545 = ~n16541 & n16544;
  assign n16546 = ~n16540 & n16545;
  assign n16547 = pi17  & n16546;
  assign n16548 = ~pi17  & ~n16546;
  assign n16549 = ~n16547 & ~n16548;
  assign n16550 = ~n16539 & ~n16549;
  assign n16551 = ~n16538 & ~n16550;
  assign n16552 = ~n16229 & ~n16551;
  assign n16553 = ~n16226 & ~n16552;
  assign n16554 = ~n16149 & ~n16150;
  assign n16555 = ~n16160 & n16554;
  assign n16556 = n16160 & ~n16554;
  assign n16557 = ~n16555 & ~n16556;
  assign n16558 = ~n16553 & n16557;
  assign n16559 = n16553 & ~n16557;
  assign n16560 = n6835 & n12636;
  assign n16561 = n7460 & n12633;
  assign n16562 = n6836 & n13292;
  assign n16563 = n7487 & n12630;
  assign n16564 = ~n16562 & ~n16563;
  assign n16565 = ~n16561 & n16564;
  assign n16566 = ~n16560 & n16565;
  assign n16567 = pi14  & n16566;
  assign n16568 = ~pi14  & ~n16566;
  assign n16569 = ~n16567 & ~n16568;
  assign n16570 = ~n16559 & ~n16569;
  assign n16571 = ~n16558 & ~n16570;
  assign n16572 = n16213 & ~n16571;
  assign n16573 = ~n16213 & n16571;
  assign n16574 = n7654 & n12622;
  assign n16575 = n8091 & n12614;
  assign n16576 = n7648 & ~n13310;
  assign n16577 = n8120 & n12606;
  assign n16578 = ~n16576 & ~n16577;
  assign n16579 = ~n16575 & n16578;
  assign n16580 = ~n16574 & n16579;
  assign n16581 = pi11  & n16580;
  assign n16582 = ~pi11  & ~n16580;
  assign n16583 = ~n16581 & ~n16582;
  assign n16584 = ~n16573 & ~n16583;
  assign n16585 = ~n16572 & ~n16584;
  assign n16586 = ~n16209 & ~n16585;
  assign n16587 = n15862 & n16176;
  assign n16588 = ~n16177 & ~n16587;
  assign n16589 = n16209 & ~n16585;
  assign n16590 = ~n16209 & n16585;
  assign n16591 = ~n16589 & ~n16590;
  assign n16592 = n16588 & ~n16591;
  assign n16593 = ~n16586 & ~n16592;
  assign n16594 = ~n16183 & ~n16184;
  assign n16595 = ~n16194 & n16594;
  assign n16596 = n16194 & ~n16594;
  assign n16597 = ~n16595 & ~n16596;
  assign n16598 = ~n16593 & n16597;
  assign n16599 = n16593 & n16597;
  assign n16600 = ~n16593 & ~n16597;
  assign n16601 = ~n16599 & ~n16600;
  assign n16602 = ~n16588 & n16591;
  assign n16603 = ~n16592 & ~n16602;
  assign n16604 = n8468 & ~n13499;
  assign n16605 = n8474 & ~n12611;
  assign n16606 = ~n8468 & ~n8473;
  assign n16607 = ~n16605 & ~n16606;
  assign n16608 = ~n12608 & ~n16607;
  assign n16609 = ~n16604 & ~n16608;
  assign n16610 = pi8  & n16609;
  assign n16611 = ~pi8  & ~n16609;
  assign n16612 = ~n16610 & ~n16611;
  assign n16613 = n16229 & n16551;
  assign n16614 = ~n16552 & ~n16613;
  assign n16615 = n6835 & n12639;
  assign n16616 = n7460 & n12636;
  assign n16617 = n6836 & n13396;
  assign n16618 = n7487 & n12633;
  assign n16619 = ~n16617 & ~n16618;
  assign n16620 = ~n16616 & n16619;
  assign n16621 = ~n16615 & n16620;
  assign n16622 = pi14  & n16621;
  assign n16623 = ~pi14  & ~n16621;
  assign n16624 = ~n16622 & ~n16623;
  assign n16625 = n16614 & ~n16624;
  assign n16626 = n16614 & n16624;
  assign n16627 = ~n16614 & ~n16624;
  assign n16628 = ~n16626 & ~n16627;
  assign n16629 = ~n16538 & ~n16539;
  assign n16630 = ~n16549 & n16629;
  assign n16631 = n16549 & ~n16629;
  assign n16632 = ~n16630 & ~n16631;
  assign n16633 = ~n16524 & ~n16525;
  assign n16634 = ~n16535 & n16633;
  assign n16635 = n16535 & ~n16633;
  assign n16636 = ~n16634 & ~n16635;
  assign n16637 = n5238 & n12680;
  assign n16638 = n71 & n12677;
  assign n16639 = n5239 & n14164;
  assign n16640 = n5326 & n12674;
  assign n16641 = ~n16639 & ~n16640;
  assign n16642 = ~n16638 & n16641;
  assign n16643 = ~n16637 & n16642;
  assign n16644 = ~pi23  & ~n16643;
  assign n16645 = pi23  & n16643;
  assign n16646 = ~n16644 & ~n16645;
  assign n16647 = n16501 & ~n16503;
  assign n16648 = ~n16504 & ~n16647;
  assign n16649 = ~n16646 & n16648;
  assign n16650 = ~n16646 & ~n16648;
  assign n16651 = n16646 & n16648;
  assign n16652 = ~n16650 & ~n16651;
  assign n16653 = n5238 & n12683;
  assign n16654 = n71 & n12680;
  assign n16655 = n5239 & n13929;
  assign n16656 = n5326 & n12677;
  assign n16657 = ~n16655 & ~n16656;
  assign n16658 = ~n16654 & n16657;
  assign n16659 = ~n16653 & n16658;
  assign n16660 = ~pi23  & ~n16659;
  assign n16661 = pi23  & n16659;
  assign n16662 = ~n16660 & ~n16661;
  assign n16663 = n16496 & n16499;
  assign n16664 = ~n16500 & ~n16663;
  assign n16665 = ~n16662 & n16664;
  assign n16666 = ~n16662 & ~n16664;
  assign n16667 = n16662 & n16664;
  assign n16668 = ~n16666 & ~n16667;
  assign n16669 = n5238 & n12686;
  assign n16670 = n71 & n12683;
  assign n16671 = n5239 & n14402;
  assign n16672 = n5326 & n12680;
  assign n16673 = ~n16671 & ~n16672;
  assign n16674 = ~n16670 & n16673;
  assign n16675 = ~n16669 & n16674;
  assign n16676 = ~pi23  & ~n16675;
  assign n16677 = pi23  & n16675;
  assign n16678 = ~n16676 & ~n16677;
  assign n16679 = n16491 & n16494;
  assign n16680 = ~n16495 & ~n16679;
  assign n16681 = ~n16678 & n16680;
  assign n16682 = ~n16678 & ~n16680;
  assign n16683 = n16678 & n16680;
  assign n16684 = ~n16682 & ~n16683;
  assign n16685 = n5238 & n12689;
  assign n16686 = n71 & n12686;
  assign n16687 = n5239 & n14552;
  assign n16688 = n5326 & n12683;
  assign n16689 = ~n16687 & ~n16688;
  assign n16690 = ~n16686 & n16689;
  assign n16691 = ~n16685 & n16690;
  assign n16692 = ~pi23  & ~n16691;
  assign n16693 = pi23  & n16691;
  assign n16694 = ~n16692 & ~n16693;
  assign n16695 = n16486 & n16489;
  assign n16696 = ~n16490 & ~n16695;
  assign n16697 = ~n16694 & n16696;
  assign n16698 = ~n16694 & ~n16696;
  assign n16699 = n16694 & n16696;
  assign n16700 = ~n16698 & ~n16699;
  assign n16701 = n5238 & n12692;
  assign n16702 = n71 & n12689;
  assign n16703 = n5239 & n14382;
  assign n16704 = n5326 & n12686;
  assign n16705 = ~n16703 & ~n16704;
  assign n16706 = ~n16702 & n16705;
  assign n16707 = ~n16701 & n16706;
  assign n16708 = ~pi23  & ~n16707;
  assign n16709 = pi23  & n16707;
  assign n16710 = ~n16708 & ~n16709;
  assign n16711 = n16481 & n16484;
  assign n16712 = ~n16485 & ~n16711;
  assign n16713 = ~n16710 & n16712;
  assign n16714 = ~n16710 & ~n16712;
  assign n16715 = n16710 & n16712;
  assign n16716 = ~n16714 & ~n16715;
  assign n16717 = n5238 & n12695;
  assign n16718 = n71 & n12692;
  assign n16719 = n5239 & n14677;
  assign n16720 = n5326 & n12689;
  assign n16721 = ~n16719 & ~n16720;
  assign n16722 = ~n16718 & n16721;
  assign n16723 = ~n16717 & n16722;
  assign n16724 = ~pi23  & ~n16723;
  assign n16725 = pi23  & n16723;
  assign n16726 = ~n16724 & ~n16725;
  assign n16727 = ~n16476 & n16479;
  assign n16728 = n16476 & ~n16479;
  assign n16729 = ~n16727 & ~n16728;
  assign n16730 = ~n16726 & ~n16729;
  assign n16731 = n5238 & n12698;
  assign n16732 = n71 & n12695;
  assign n16733 = n5239 & n14976;
  assign n16734 = n5326 & n12692;
  assign n16735 = ~n16733 & ~n16734;
  assign n16736 = ~n16732 & n16735;
  assign n16737 = ~n16731 & n16736;
  assign n16738 = ~pi23  & ~n16737;
  assign n16739 = pi23  & n16737;
  assign n16740 = ~n16738 & ~n16739;
  assign n16741 = ~n16471 & n16474;
  assign n16742 = n16471 & ~n16474;
  assign n16743 = ~n16741 & ~n16742;
  assign n16744 = ~n16740 & ~n16743;
  assign n16745 = n5238 & n12701;
  assign n16746 = n71 & n12698;
  assign n16747 = n5239 & n14991;
  assign n16748 = n5326 & n12695;
  assign n16749 = ~n16747 & ~n16748;
  assign n16750 = ~n16746 & n16749;
  assign n16751 = ~n16745 & n16750;
  assign n16752 = ~pi23  & ~n16751;
  assign n16753 = pi23  & n16751;
  assign n16754 = ~n16752 & ~n16753;
  assign n16755 = ~n16466 & n16469;
  assign n16756 = n16466 & ~n16469;
  assign n16757 = ~n16755 & ~n16756;
  assign n16758 = ~n16754 & ~n16757;
  assign n16759 = n5238 & n12704;
  assign n16760 = n71 & n12701;
  assign n16761 = n5239 & n14655;
  assign n16762 = n5326 & n12698;
  assign n16763 = ~n16761 & ~n16762;
  assign n16764 = ~n16760 & n16763;
  assign n16765 = ~n16759 & n16764;
  assign n16766 = ~pi23  & ~n16765;
  assign n16767 = pi23  & n16765;
  assign n16768 = ~n16766 & ~n16767;
  assign n16769 = n16461 & n16464;
  assign n16770 = ~n16465 & ~n16769;
  assign n16771 = ~n16768 & n16770;
  assign n16772 = ~n16768 & ~n16770;
  assign n16773 = n16768 & n16770;
  assign n16774 = ~n16772 & ~n16773;
  assign n16775 = n5238 & n12707;
  assign n16776 = n71 & n12704;
  assign n16777 = n5239 & n15024;
  assign n16778 = n5326 & n12701;
  assign n16779 = ~n16777 & ~n16778;
  assign n16780 = ~n16776 & n16779;
  assign n16781 = ~n16775 & n16780;
  assign n16782 = ~pi23  & ~n16781;
  assign n16783 = pi23  & n16781;
  assign n16784 = ~n16782 & ~n16783;
  assign n16785 = n16456 & n16459;
  assign n16786 = ~n16460 & ~n16785;
  assign n16787 = ~n16784 & n16786;
  assign n16788 = ~n16784 & ~n16786;
  assign n16789 = n16784 & n16786;
  assign n16790 = ~n16788 & ~n16789;
  assign n16791 = n16383 & n16454;
  assign n16792 = ~n16455 & ~n16791;
  assign n16793 = n5238 & n12710;
  assign n16794 = n71 & n12707;
  assign n16795 = n5239 & n15050;
  assign n16796 = n5326 & n12704;
  assign n16797 = ~n16795 & ~n16796;
  assign n16798 = ~n16794 & n16797;
  assign n16799 = ~n16793 & n16798;
  assign n16800 = pi23  & n16799;
  assign n16801 = ~pi23  & ~n16799;
  assign n16802 = ~n16800 & ~n16801;
  assign n16803 = n16792 & ~n16802;
  assign n16804 = n16401 & n16452;
  assign n16805 = ~n16453 & ~n16804;
  assign n16806 = n5238 & n12713;
  assign n16807 = n71 & n12710;
  assign n16808 = n5239 & n15074;
  assign n16809 = n5326 & n12707;
  assign n16810 = ~n16808 & ~n16809;
  assign n16811 = ~n16807 & n16810;
  assign n16812 = ~n16806 & n16811;
  assign n16813 = pi23  & n16812;
  assign n16814 = ~pi23  & ~n16812;
  assign n16815 = ~n16813 & ~n16814;
  assign n16816 = n16805 & ~n16815;
  assign n16817 = n5238 & n12716;
  assign n16818 = n71 & n12713;
  assign n16819 = n5239 & n15105;
  assign n16820 = n5326 & n12710;
  assign n16821 = ~n16819 & ~n16820;
  assign n16822 = ~n16818 & n16821;
  assign n16823 = ~n16817 & n16822;
  assign n16824 = ~pi23  & ~n16823;
  assign n16825 = pi23  & n16823;
  assign n16826 = ~n16824 & ~n16825;
  assign n16827 = n16448 & ~n16450;
  assign n16828 = ~n16451 & ~n16827;
  assign n16829 = ~n16826 & n16828;
  assign n16830 = ~n16826 & ~n16828;
  assign n16831 = n16826 & n16828;
  assign n16832 = ~n16830 & ~n16831;
  assign n16833 = n5238 & n12719;
  assign n16834 = n71 & n12716;
  assign n16835 = n5239 & n15161;
  assign n16836 = n5326 & n12713;
  assign n16837 = ~n16835 & ~n16836;
  assign n16838 = ~n16834 & n16837;
  assign n16839 = ~n16833 & n16838;
  assign n16840 = pi23  & n16839;
  assign n16841 = ~pi23  & ~n16839;
  assign n16842 = ~n16840 & ~n16841;
  assign n16843 = n16436 & n16446;
  assign n16844 = ~n16447 & ~n16843;
  assign n16845 = ~n16842 & n16844;
  assign n16846 = n5238 & n12722;
  assign n16847 = n71 & n12719;
  assign n16848 = n5239 & n15199;
  assign n16849 = n5326 & n12716;
  assign n16850 = ~n16848 & ~n16849;
  assign n16851 = ~n16847 & n16850;
  assign n16852 = ~n16846 & n16851;
  assign n16853 = ~pi23  & ~n16852;
  assign n16854 = pi23  & n16852;
  assign n16855 = ~n16853 & ~n16854;
  assign n16856 = pi26  & ~n16424;
  assign n16857 = n16431 & ~n16856;
  assign n16858 = ~n16431 & n16856;
  assign n16859 = ~n16857 & ~n16858;
  assign n16860 = ~n16855 & n16859;
  assign n16861 = ~n16855 & ~n16859;
  assign n16862 = n16855 & n16859;
  assign n16863 = ~n16861 & ~n16862;
  assign n16864 = n5238 & n12725;
  assign n16865 = n71 & n12722;
  assign n16866 = n5239 & n15243;
  assign n16867 = n5326 & n12719;
  assign n16868 = ~n16866 & ~n16867;
  assign n16869 = ~n16865 & n16868;
  assign n16870 = ~n16864 & n16869;
  assign n16871 = pi23  & n16870;
  assign n16872 = ~pi23  & ~n16870;
  assign n16873 = ~n16871 & ~n16872;
  assign n16874 = pi26  & n16422;
  assign n16875 = ~n16421 & n16874;
  assign n16876 = n16421 & ~n16874;
  assign n16877 = ~n16875 & ~n16876;
  assign n16878 = ~n16873 & n16877;
  assign n16879 = n5239 & ~n15312;
  assign n16880 = n5326 & n12730;
  assign n16881 = n71 & n12732;
  assign n16882 = ~n16880 & ~n16881;
  assign n16883 = ~n16879 & n16882;
  assign n16884 = ~n70 & n12732;
  assign n16885 = pi23  & ~n16884;
  assign n16886 = n16883 & n16885;
  assign n16887 = n5238 & n12732;
  assign n16888 = n71 & n12730;
  assign n16889 = n5239 & ~n15356;
  assign n16890 = n5326 & n12725;
  assign n16891 = ~n16889 & ~n16890;
  assign n16892 = ~n16888 & n16891;
  assign n16893 = ~n16887 & n16892;
  assign n16894 = n16886 & n16893;
  assign n16895 = n16422 & n16894;
  assign n16896 = ~n16422 & n16894;
  assign n16897 = n16422 & ~n16894;
  assign n16898 = ~n16896 & ~n16897;
  assign n16899 = n5238 & n12730;
  assign n16900 = n71 & n12725;
  assign n16901 = n5239 & n15267;
  assign n16902 = n5326 & n12722;
  assign n16903 = ~n16901 & ~n16902;
  assign n16904 = ~n16900 & n16903;
  assign n16905 = ~n16899 & n16904;
  assign n16906 = pi23  & n16905;
  assign n16907 = ~pi23  & ~n16905;
  assign n16908 = ~n16906 & ~n16907;
  assign n16909 = ~n16898 & ~n16908;
  assign n16910 = ~n16895 & ~n16909;
  assign n16911 = n16873 & ~n16877;
  assign n16912 = ~n16878 & ~n16911;
  assign n16913 = ~n16910 & n16912;
  assign n16914 = ~n16878 & ~n16913;
  assign n16915 = ~n16863 & ~n16914;
  assign n16916 = ~n16860 & ~n16915;
  assign n16917 = n16842 & ~n16844;
  assign n16918 = ~n16845 & ~n16917;
  assign n16919 = ~n16916 & n16918;
  assign n16920 = ~n16845 & ~n16919;
  assign n16921 = ~n16832 & ~n16920;
  assign n16922 = ~n16829 & ~n16921;
  assign n16923 = n16805 & n16815;
  assign n16924 = ~n16805 & ~n16815;
  assign n16925 = ~n16923 & ~n16924;
  assign n16926 = ~n16922 & ~n16925;
  assign n16927 = ~n16816 & ~n16926;
  assign n16928 = ~n16792 & n16802;
  assign n16929 = ~n16803 & ~n16928;
  assign n16930 = ~n16927 & n16929;
  assign n16931 = ~n16803 & ~n16930;
  assign n16932 = ~n16790 & ~n16931;
  assign n16933 = ~n16787 & ~n16932;
  assign n16934 = ~n16774 & ~n16933;
  assign n16935 = ~n16771 & ~n16934;
  assign n16936 = n16754 & n16757;
  assign n16937 = ~n16758 & ~n16936;
  assign n16938 = ~n16935 & n16937;
  assign n16939 = ~n16758 & ~n16938;
  assign n16940 = n16740 & n16743;
  assign n16941 = ~n16744 & ~n16940;
  assign n16942 = ~n16939 & n16941;
  assign n16943 = ~n16744 & ~n16942;
  assign n16944 = n16726 & n16729;
  assign n16945 = ~n16730 & ~n16944;
  assign n16946 = ~n16943 & n16945;
  assign n16947 = ~n16730 & ~n16946;
  assign n16948 = ~n16716 & ~n16947;
  assign n16949 = ~n16713 & ~n16948;
  assign n16950 = ~n16700 & ~n16949;
  assign n16951 = ~n16697 & ~n16950;
  assign n16952 = ~n16684 & ~n16951;
  assign n16953 = ~n16681 & ~n16952;
  assign n16954 = ~n16668 & ~n16953;
  assign n16955 = ~n16665 & ~n16954;
  assign n16956 = ~n16652 & ~n16955;
  assign n16957 = ~n16649 & ~n16956;
  assign n16958 = ~n16510 & ~n16511;
  assign n16959 = ~n16521 & n16958;
  assign n16960 = n16521 & ~n16958;
  assign n16961 = ~n16959 & ~n16960;
  assign n16962 = ~n16957 & n16961;
  assign n16963 = n16957 & ~n16961;
  assign n16964 = n5435 & n12668;
  assign n16965 = n6055 & n12665;
  assign n16966 = n5429 & n13591;
  assign n16967 = n6071 & n12662;
  assign n16968 = ~n16966 & ~n16967;
  assign n16969 = ~n16965 & n16968;
  assign n16970 = ~n16964 & n16969;
  assign n16971 = pi20  & n16970;
  assign n16972 = ~pi20  & ~n16970;
  assign n16973 = ~n16971 & ~n16972;
  assign n16974 = ~n16963 & ~n16973;
  assign n16975 = ~n16962 & ~n16974;
  assign n16976 = n16636 & ~n16975;
  assign n16977 = ~n16636 & n16975;
  assign n16978 = n6184 & n12656;
  assign n16979 = n6527 & n12653;
  assign n16980 = n6185 & n12991;
  assign n16981 = n6543 & n12650;
  assign n16982 = ~n16980 & ~n16981;
  assign n16983 = ~n16979 & n16982;
  assign n16984 = ~n16978 & n16983;
  assign n16985 = pi17  & n16984;
  assign n16986 = ~pi17  & ~n16984;
  assign n16987 = ~n16985 & ~n16986;
  assign n16988 = ~n16977 & ~n16987;
  assign n16989 = ~n16976 & ~n16988;
  assign n16990 = n16632 & ~n16989;
  assign n16991 = ~n16632 & n16989;
  assign n16992 = n6835 & n12644;
  assign n16993 = n7460 & n12639;
  assign n16994 = n6836 & n13210;
  assign n16995 = n7487 & n12636;
  assign n16996 = ~n16994 & ~n16995;
  assign n16997 = ~n16993 & n16996;
  assign n16998 = ~n16992 & n16997;
  assign n16999 = pi14  & n16998;
  assign n17000 = ~pi14  & ~n16998;
  assign n17001 = ~n16999 & ~n17000;
  assign n17002 = ~n16991 & ~n17001;
  assign n17003 = ~n16990 & ~n17002;
  assign n17004 = ~n16628 & ~n17003;
  assign n17005 = ~n16625 & ~n17004;
  assign n17006 = ~n16558 & ~n16559;
  assign n17007 = ~n16569 & n17006;
  assign n17008 = n16569 & ~n17006;
  assign n17009 = ~n17007 & ~n17008;
  assign n17010 = ~n17005 & n17009;
  assign n17011 = n17005 & ~n17009;
  assign n17012 = n7654 & n12625;
  assign n17013 = n8091 & n12622;
  assign n17014 = n7648 & n13463;
  assign n17015 = n8120 & n12614;
  assign n17016 = ~n17014 & ~n17015;
  assign n17017 = ~n17013 & n17016;
  assign n17018 = ~n17012 & n17017;
  assign n17019 = pi11  & n17018;
  assign n17020 = ~pi11  & ~n17018;
  assign n17021 = ~n17019 & ~n17020;
  assign n17022 = ~n17011 & ~n17021;
  assign n17023 = ~n17010 & ~n17022;
  assign n17024 = ~n16612 & ~n17023;
  assign n17025 = n16612 & n17023;
  assign n17026 = ~n16572 & ~n16573;
  assign n17027 = ~n16583 & n17026;
  assign n17028 = n16583 & ~n17026;
  assign n17029 = ~n17027 & ~n17028;
  assign n17030 = ~n17025 & n17029;
  assign n17031 = ~n17024 & ~n17030;
  assign n17032 = n16603 & ~n17031;
  assign n17033 = ~n17024 & ~n17025;
  assign n17034 = n17029 & n17033;
  assign n17035 = ~n17029 & ~n17033;
  assign n17036 = ~n17034 & ~n17035;
  assign n17037 = n16628 & n17003;
  assign n17038 = ~n17004 & ~n17037;
  assign n17039 = n7654 & n12630;
  assign n17040 = n8091 & n12625;
  assign n17041 = n7648 & n13325;
  assign n17042 = n8120 & n12622;
  assign n17043 = ~n17041 & ~n17042;
  assign n17044 = ~n17040 & n17043;
  assign n17045 = ~n17039 & n17044;
  assign n17046 = pi11  & n17045;
  assign n17047 = ~pi11  & ~n17045;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = n17038 & ~n17048;
  assign n17050 = n17038 & n17048;
  assign n17051 = ~n17038 & ~n17048;
  assign n17052 = ~n17050 & ~n17051;
  assign n17053 = ~n16990 & ~n16991;
  assign n17054 = ~n17001 & n17053;
  assign n17055 = n17001 & ~n17053;
  assign n17056 = ~n17054 & ~n17055;
  assign n17057 = ~n16976 & ~n16977;
  assign n17058 = ~n16987 & n17057;
  assign n17059 = n16987 & ~n17057;
  assign n17060 = ~n17058 & ~n17059;
  assign n17061 = n16652 & n16955;
  assign n17062 = ~n16956 & ~n17061;
  assign n17063 = n5435 & n12671;
  assign n17064 = n6055 & n12668;
  assign n17065 = n5429 & n13578;
  assign n17066 = n6071 & n12665;
  assign n17067 = ~n17065 & ~n17066;
  assign n17068 = ~n17064 & n17067;
  assign n17069 = ~n17063 & n17068;
  assign n17070 = pi20  & n17069;
  assign n17071 = ~pi20  & ~n17069;
  assign n17072 = ~n17070 & ~n17071;
  assign n17073 = n17062 & ~n17072;
  assign n17074 = n16668 & n16953;
  assign n17075 = ~n16954 & ~n17074;
  assign n17076 = n5435 & n12674;
  assign n17077 = n6055 & n12671;
  assign n17078 = n5429 & n13764;
  assign n17079 = n6071 & n12668;
  assign n17080 = ~n17078 & ~n17079;
  assign n17081 = ~n17077 & n17080;
  assign n17082 = ~n17076 & n17081;
  assign n17083 = pi20  & n17082;
  assign n17084 = ~pi20  & ~n17082;
  assign n17085 = ~n17083 & ~n17084;
  assign n17086 = n17075 & ~n17085;
  assign n17087 = n16684 & n16951;
  assign n17088 = ~n16952 & ~n17087;
  assign n17089 = n5435 & n12677;
  assign n17090 = n6055 & n12674;
  assign n17091 = n5429 & n13785;
  assign n17092 = n6071 & n12671;
  assign n17093 = ~n17091 & ~n17092;
  assign n17094 = ~n17090 & n17093;
  assign n17095 = ~n17089 & n17094;
  assign n17096 = pi20  & n17095;
  assign n17097 = ~pi20  & ~n17095;
  assign n17098 = ~n17096 & ~n17097;
  assign n17099 = n17088 & ~n17098;
  assign n17100 = n16700 & n16949;
  assign n17101 = ~n16950 & ~n17100;
  assign n17102 = n5435 & n12680;
  assign n17103 = n6055 & n12677;
  assign n17104 = n5429 & n14164;
  assign n17105 = n6071 & n12674;
  assign n17106 = ~n17104 & ~n17105;
  assign n17107 = ~n17103 & n17106;
  assign n17108 = ~n17102 & n17107;
  assign n17109 = pi20  & n17108;
  assign n17110 = ~pi20  & ~n17108;
  assign n17111 = ~n17109 & ~n17110;
  assign n17112 = n17101 & ~n17111;
  assign n17113 = n16716 & n16947;
  assign n17114 = ~n16948 & ~n17113;
  assign n17115 = n5435 & n12683;
  assign n17116 = n6055 & n12680;
  assign n17117 = n5429 & n13929;
  assign n17118 = n6071 & n12677;
  assign n17119 = ~n17117 & ~n17118;
  assign n17120 = ~n17116 & n17119;
  assign n17121 = ~n17115 & n17120;
  assign n17122 = pi20  & n17121;
  assign n17123 = ~pi20  & ~n17121;
  assign n17124 = ~n17122 & ~n17123;
  assign n17125 = n17114 & ~n17124;
  assign n17126 = n16943 & ~n16945;
  assign n17127 = ~n16946 & ~n17126;
  assign n17128 = n5435 & n12686;
  assign n17129 = n6055 & n12683;
  assign n17130 = n5429 & n14402;
  assign n17131 = n6071 & n12680;
  assign n17132 = ~n17130 & ~n17131;
  assign n17133 = ~n17129 & n17132;
  assign n17134 = ~n17128 & n17133;
  assign n17135 = pi20  & n17134;
  assign n17136 = ~pi20  & ~n17134;
  assign n17137 = ~n17135 & ~n17136;
  assign n17138 = n17127 & ~n17137;
  assign n17139 = n16939 & ~n16941;
  assign n17140 = ~n16942 & ~n17139;
  assign n17141 = n5435 & n12689;
  assign n17142 = n6055 & n12686;
  assign n17143 = n5429 & n14552;
  assign n17144 = n6071 & n12683;
  assign n17145 = ~n17143 & ~n17144;
  assign n17146 = ~n17142 & n17145;
  assign n17147 = ~n17141 & n17146;
  assign n17148 = pi20  & n17147;
  assign n17149 = ~pi20  & ~n17147;
  assign n17150 = ~n17148 & ~n17149;
  assign n17151 = n17140 & ~n17150;
  assign n17152 = n16935 & ~n16937;
  assign n17153 = ~n16938 & ~n17152;
  assign n17154 = n5435 & n12692;
  assign n17155 = n6055 & n12689;
  assign n17156 = n5429 & n14382;
  assign n17157 = n6071 & n12686;
  assign n17158 = ~n17156 & ~n17157;
  assign n17159 = ~n17155 & n17158;
  assign n17160 = ~n17154 & n17159;
  assign n17161 = pi20  & n17160;
  assign n17162 = ~pi20  & ~n17160;
  assign n17163 = ~n17161 & ~n17162;
  assign n17164 = n17153 & ~n17163;
  assign n17165 = n16774 & n16933;
  assign n17166 = ~n16934 & ~n17165;
  assign n17167 = n5435 & n12695;
  assign n17168 = n6055 & n12692;
  assign n17169 = n5429 & n14677;
  assign n17170 = n6071 & n12689;
  assign n17171 = ~n17169 & ~n17170;
  assign n17172 = ~n17168 & n17171;
  assign n17173 = ~n17167 & n17172;
  assign n17174 = pi20  & n17173;
  assign n17175 = ~pi20  & ~n17173;
  assign n17176 = ~n17174 & ~n17175;
  assign n17177 = n17166 & ~n17176;
  assign n17178 = n16790 & n16931;
  assign n17179 = ~n16932 & ~n17178;
  assign n17180 = n5435 & n12698;
  assign n17181 = n6055 & n12695;
  assign n17182 = n5429 & n14976;
  assign n17183 = n6071 & n12692;
  assign n17184 = ~n17182 & ~n17183;
  assign n17185 = ~n17181 & n17184;
  assign n17186 = ~n17180 & n17185;
  assign n17187 = pi20  & n17186;
  assign n17188 = ~pi20  & ~n17186;
  assign n17189 = ~n17187 & ~n17188;
  assign n17190 = n17179 & ~n17189;
  assign n17191 = n5435 & n12701;
  assign n17192 = n6055 & n12698;
  assign n17193 = n5429 & n14991;
  assign n17194 = n6071 & n12695;
  assign n17195 = ~n17193 & ~n17194;
  assign n17196 = ~n17192 & n17195;
  assign n17197 = ~n17191 & n17196;
  assign n17198 = ~pi20  & ~n17197;
  assign n17199 = pi20  & n17197;
  assign n17200 = ~n17198 & ~n17199;
  assign n17201 = n16927 & ~n16929;
  assign n17202 = ~n16930 & ~n17201;
  assign n17203 = ~n17200 & n17202;
  assign n17204 = ~n17200 & ~n17202;
  assign n17205 = n17200 & n17202;
  assign n17206 = ~n17204 & ~n17205;
  assign n17207 = n5435 & n12704;
  assign n17208 = n6055 & n12701;
  assign n17209 = n5429 & n14655;
  assign n17210 = n6071 & n12698;
  assign n17211 = ~n17209 & ~n17210;
  assign n17212 = ~n17208 & n17211;
  assign n17213 = ~n17207 & n17212;
  assign n17214 = ~pi20  & ~n17213;
  assign n17215 = pi20  & n17213;
  assign n17216 = ~n17214 & ~n17215;
  assign n17217 = ~n16922 & n16925;
  assign n17218 = n16922 & ~n16925;
  assign n17219 = ~n17217 & ~n17218;
  assign n17220 = ~n17216 & ~n17219;
  assign n17221 = n16832 & n16920;
  assign n17222 = ~n16921 & ~n17221;
  assign n17223 = n5435 & n12707;
  assign n17224 = n6055 & n12704;
  assign n17225 = n5429 & n15024;
  assign n17226 = n6071 & n12701;
  assign n17227 = ~n17225 & ~n17226;
  assign n17228 = ~n17224 & n17227;
  assign n17229 = ~n17223 & n17228;
  assign n17230 = pi20  & n17229;
  assign n17231 = ~pi20  & ~n17229;
  assign n17232 = ~n17230 & ~n17231;
  assign n17233 = n17222 & ~n17232;
  assign n17234 = n16916 & ~n16918;
  assign n17235 = ~n16919 & ~n17234;
  assign n17236 = n5435 & n12710;
  assign n17237 = n6055 & n12707;
  assign n17238 = n5429 & n15050;
  assign n17239 = n6071 & n12704;
  assign n17240 = ~n17238 & ~n17239;
  assign n17241 = ~n17237 & n17240;
  assign n17242 = ~n17236 & n17241;
  assign n17243 = pi20  & n17242;
  assign n17244 = ~pi20  & ~n17242;
  assign n17245 = ~n17243 & ~n17244;
  assign n17246 = n17235 & ~n17245;
  assign n17247 = n16863 & n16914;
  assign n17248 = ~n16915 & ~n17247;
  assign n17249 = n5435 & n12713;
  assign n17250 = n6055 & n12710;
  assign n17251 = n5429 & n15074;
  assign n17252 = n6071 & n12707;
  assign n17253 = ~n17251 & ~n17252;
  assign n17254 = ~n17250 & n17253;
  assign n17255 = ~n17249 & n17254;
  assign n17256 = pi20  & n17255;
  assign n17257 = ~pi20  & ~n17255;
  assign n17258 = ~n17256 & ~n17257;
  assign n17259 = n17248 & ~n17258;
  assign n17260 = n5435 & n12716;
  assign n17261 = n6055 & n12713;
  assign n17262 = n5429 & n15105;
  assign n17263 = n6071 & n12710;
  assign n17264 = ~n17262 & ~n17263;
  assign n17265 = ~n17261 & n17264;
  assign n17266 = ~n17260 & n17265;
  assign n17267 = ~pi20  & ~n17266;
  assign n17268 = pi20  & n17266;
  assign n17269 = ~n17267 & ~n17268;
  assign n17270 = n16910 & ~n16912;
  assign n17271 = ~n16913 & ~n17270;
  assign n17272 = ~n17269 & n17271;
  assign n17273 = ~n17269 & ~n17271;
  assign n17274 = n17269 & n17271;
  assign n17275 = ~n17273 & ~n17274;
  assign n17276 = n5435 & n12719;
  assign n17277 = n6055 & n12716;
  assign n17278 = n5429 & n15161;
  assign n17279 = n6071 & n12713;
  assign n17280 = ~n17278 & ~n17279;
  assign n17281 = ~n17277 & n17280;
  assign n17282 = ~n17276 & n17281;
  assign n17283 = pi20  & n17282;
  assign n17284 = ~pi20  & ~n17282;
  assign n17285 = ~n17283 & ~n17284;
  assign n17286 = n16898 & n16908;
  assign n17287 = ~n16909 & ~n17286;
  assign n17288 = ~n17285 & n17287;
  assign n17289 = n5435 & n12722;
  assign n17290 = n6055 & n12719;
  assign n17291 = n5429 & n15199;
  assign n17292 = n6071 & n12716;
  assign n17293 = ~n17291 & ~n17292;
  assign n17294 = ~n17290 & n17293;
  assign n17295 = ~n17289 & n17294;
  assign n17296 = ~pi20  & ~n17295;
  assign n17297 = pi20  & n17295;
  assign n17298 = ~n17296 & ~n17297;
  assign n17299 = pi23  & ~n16886;
  assign n17300 = n16893 & ~n17299;
  assign n17301 = ~n16893 & n17299;
  assign n17302 = ~n17300 & ~n17301;
  assign n17303 = ~n17298 & n17302;
  assign n17304 = ~n17298 & ~n17302;
  assign n17305 = n17298 & n17302;
  assign n17306 = ~n17304 & ~n17305;
  assign n17307 = n5435 & n12725;
  assign n17308 = n6055 & n12722;
  assign n17309 = n5429 & n15243;
  assign n17310 = n6071 & n12719;
  assign n17311 = ~n17309 & ~n17310;
  assign n17312 = ~n17308 & n17311;
  assign n17313 = ~n17307 & n17312;
  assign n17314 = pi20  & n17313;
  assign n17315 = ~pi20  & ~n17313;
  assign n17316 = ~n17314 & ~n17315;
  assign n17317 = pi23  & n16884;
  assign n17318 = ~n16883 & n17317;
  assign n17319 = n16883 & ~n17317;
  assign n17320 = ~n17318 & ~n17319;
  assign n17321 = ~n17316 & n17320;
  assign n17322 = n5429 & ~n15312;
  assign n17323 = n6071 & n12730;
  assign n17324 = n6055 & n12732;
  assign n17325 = ~n17323 & ~n17324;
  assign n17326 = ~n17322 & n17325;
  assign n17327 = ~n5425 & n12732;
  assign n17328 = pi20  & ~n17327;
  assign n17329 = n17326 & n17328;
  assign n17330 = n5435 & n12732;
  assign n17331 = n6055 & n12730;
  assign n17332 = n5429 & ~n15356;
  assign n17333 = n6071 & n12725;
  assign n17334 = ~n17332 & ~n17333;
  assign n17335 = ~n17331 & n17334;
  assign n17336 = ~n17330 & n17335;
  assign n17337 = n17329 & n17336;
  assign n17338 = n16884 & n17337;
  assign n17339 = ~n16884 & n17337;
  assign n17340 = n16884 & ~n17337;
  assign n17341 = ~n17339 & ~n17340;
  assign n17342 = n5435 & n12730;
  assign n17343 = n6055 & n12725;
  assign n17344 = n5429 & n15267;
  assign n17345 = n6071 & n12722;
  assign n17346 = ~n17344 & ~n17345;
  assign n17347 = ~n17343 & n17346;
  assign n17348 = ~n17342 & n17347;
  assign n17349 = pi20  & n17348;
  assign n17350 = ~pi20  & ~n17348;
  assign n17351 = ~n17349 & ~n17350;
  assign n17352 = ~n17341 & ~n17351;
  assign n17353 = ~n17338 & ~n17352;
  assign n17354 = n17316 & ~n17320;
  assign n17355 = ~n17321 & ~n17354;
  assign n17356 = ~n17353 & n17355;
  assign n17357 = ~n17321 & ~n17356;
  assign n17358 = ~n17306 & ~n17357;
  assign n17359 = ~n17303 & ~n17358;
  assign n17360 = n17285 & ~n17287;
  assign n17361 = ~n17288 & ~n17360;
  assign n17362 = ~n17359 & n17361;
  assign n17363 = ~n17288 & ~n17362;
  assign n17364 = ~n17275 & ~n17363;
  assign n17365 = ~n17272 & ~n17364;
  assign n17366 = n17248 & n17258;
  assign n17367 = ~n17248 & ~n17258;
  assign n17368 = ~n17366 & ~n17367;
  assign n17369 = ~n17365 & ~n17368;
  assign n17370 = ~n17259 & ~n17369;
  assign n17371 = n17235 & n17245;
  assign n17372 = ~n17235 & ~n17245;
  assign n17373 = ~n17371 & ~n17372;
  assign n17374 = ~n17370 & ~n17373;
  assign n17375 = ~n17246 & ~n17374;
  assign n17376 = ~n17222 & n17232;
  assign n17377 = ~n17233 & ~n17376;
  assign n17378 = ~n17375 & n17377;
  assign n17379 = ~n17233 & ~n17378;
  assign n17380 = n17216 & n17219;
  assign n17381 = ~n17220 & ~n17380;
  assign n17382 = ~n17379 & n17381;
  assign n17383 = ~n17220 & ~n17382;
  assign n17384 = ~n17206 & ~n17383;
  assign n17385 = ~n17203 & ~n17384;
  assign n17386 = n17179 & n17189;
  assign n17387 = ~n17179 & ~n17189;
  assign n17388 = ~n17386 & ~n17387;
  assign n17389 = ~n17385 & ~n17388;
  assign n17390 = ~n17190 & ~n17389;
  assign n17391 = n17166 & n17176;
  assign n17392 = ~n17166 & ~n17176;
  assign n17393 = ~n17391 & ~n17392;
  assign n17394 = ~n17390 & ~n17393;
  assign n17395 = ~n17177 & ~n17394;
  assign n17396 = n17153 & n17163;
  assign n17397 = ~n17153 & ~n17163;
  assign n17398 = ~n17396 & ~n17397;
  assign n17399 = ~n17395 & ~n17398;
  assign n17400 = ~n17164 & ~n17399;
  assign n17401 = n17140 & n17150;
  assign n17402 = ~n17140 & ~n17150;
  assign n17403 = ~n17401 & ~n17402;
  assign n17404 = ~n17400 & ~n17403;
  assign n17405 = ~n17151 & ~n17404;
  assign n17406 = n17127 & n17137;
  assign n17407 = ~n17127 & ~n17137;
  assign n17408 = ~n17406 & ~n17407;
  assign n17409 = ~n17405 & ~n17408;
  assign n17410 = ~n17138 & ~n17409;
  assign n17411 = n17114 & n17124;
  assign n17412 = ~n17114 & ~n17124;
  assign n17413 = ~n17411 & ~n17412;
  assign n17414 = ~n17410 & ~n17413;
  assign n17415 = ~n17125 & ~n17414;
  assign n17416 = n17101 & n17111;
  assign n17417 = ~n17101 & ~n17111;
  assign n17418 = ~n17416 & ~n17417;
  assign n17419 = ~n17415 & ~n17418;
  assign n17420 = ~n17112 & ~n17419;
  assign n17421 = n17088 & n17098;
  assign n17422 = ~n17088 & ~n17098;
  assign n17423 = ~n17421 & ~n17422;
  assign n17424 = ~n17420 & ~n17423;
  assign n17425 = ~n17099 & ~n17424;
  assign n17426 = n17075 & n17085;
  assign n17427 = ~n17075 & ~n17085;
  assign n17428 = ~n17426 & ~n17427;
  assign n17429 = ~n17425 & ~n17428;
  assign n17430 = ~n17086 & ~n17429;
  assign n17431 = ~n17062 & n17072;
  assign n17432 = ~n17073 & ~n17431;
  assign n17433 = ~n17430 & n17432;
  assign n17434 = ~n17073 & ~n17433;
  assign n17435 = ~n16962 & ~n16963;
  assign n17436 = ~n16973 & n17435;
  assign n17437 = n16973 & ~n17435;
  assign n17438 = ~n17436 & ~n17437;
  assign n17439 = ~n17434 & n17438;
  assign n17440 = n17434 & ~n17438;
  assign n17441 = n6184 & n12659;
  assign n17442 = n6527 & n12656;
  assign n17443 = n6185 & n13059;
  assign n17444 = n6543 & n12653;
  assign n17445 = ~n17443 & ~n17444;
  assign n17446 = ~n17442 & n17445;
  assign n17447 = ~n17441 & n17446;
  assign n17448 = pi17  & n17447;
  assign n17449 = ~pi17  & ~n17447;
  assign n17450 = ~n17448 & ~n17449;
  assign n17451 = ~n17440 & ~n17450;
  assign n17452 = ~n17439 & ~n17451;
  assign n17453 = n17060 & ~n17452;
  assign n17454 = ~n17060 & n17452;
  assign n17455 = n6835 & n12647;
  assign n17456 = n7460 & n12644;
  assign n17457 = n6836 & ~n13193;
  assign n17458 = n7487 & n12639;
  assign n17459 = ~n17457 & ~n17458;
  assign n17460 = ~n17456 & n17459;
  assign n17461 = ~n17455 & n17460;
  assign n17462 = pi14  & n17461;
  assign n17463 = ~pi14  & ~n17461;
  assign n17464 = ~n17462 & ~n17463;
  assign n17465 = ~n17454 & ~n17464;
  assign n17466 = ~n17453 & ~n17465;
  assign n17467 = n17056 & ~n17466;
  assign n17468 = ~n17056 & n17466;
  assign n17469 = n7654 & n12633;
  assign n17470 = n8091 & n12630;
  assign n17471 = n7648 & ~n13227;
  assign n17472 = n8120 & n12625;
  assign n17473 = ~n17471 & ~n17472;
  assign n17474 = ~n17470 & n17473;
  assign n17475 = ~n17469 & n17474;
  assign n17476 = pi11  & n17475;
  assign n17477 = ~pi11  & ~n17475;
  assign n17478 = ~n17476 & ~n17477;
  assign n17479 = ~n17468 & ~n17478;
  assign n17480 = ~n17467 & ~n17479;
  assign n17481 = ~n17052 & ~n17480;
  assign n17482 = ~n17049 & ~n17481;
  assign n17483 = ~n17010 & ~n17011;
  assign n17484 = ~n17021 & n17483;
  assign n17485 = n17021 & ~n17483;
  assign n17486 = ~n17484 & ~n17485;
  assign n17487 = ~n17482 & n17486;
  assign n17488 = n17482 & ~n17486;
  assign n17489 = n8474 & n12606;
  assign n17490 = n9238 & n12616;
  assign n17491 = n8468 & ~n13483;
  assign n17492 = n9265 & ~n12608;
  assign n17493 = ~n17491 & ~n17492;
  assign n17494 = ~n17490 & n17493;
  assign n17495 = ~n17489 & n17494;
  assign n17496 = pi8  & n17495;
  assign n17497 = ~pi8  & ~n17495;
  assign n17498 = ~n17496 & ~n17497;
  assign n17499 = ~n17488 & ~n17498;
  assign n17500 = ~n17487 & ~n17499;
  assign n17501 = n17036 & ~n17500;
  assign n17502 = ~n17036 & n17500;
  assign n17503 = ~n17501 & ~n17502;
  assign n17504 = n9238 & n12606;
  assign n17505 = ~n12611 & n17492;
  assign n17506 = n8474 & n12614;
  assign n17507 = n8468 & n12868;
  assign n17508 = ~n17506 & ~n17507;
  assign n17509 = ~n17505 & n17508;
  assign n17510 = ~n17504 & n17509;
  assign n17511 = pi8  & n17510;
  assign n17512 = ~pi8  & ~n17510;
  assign n17513 = ~n17511 & ~n17512;
  assign n17514 = ~n17467 & ~n17468;
  assign n17515 = ~n17478 & n17514;
  assign n17516 = n17478 & ~n17514;
  assign n17517 = ~n17515 & ~n17516;
  assign n17518 = ~n17453 & ~n17454;
  assign n17519 = ~n17464 & n17518;
  assign n17520 = n17464 & ~n17518;
  assign n17521 = ~n17519 & ~n17520;
  assign n17522 = n6184 & n12662;
  assign n17523 = n6527 & n12659;
  assign n17524 = n6185 & n13246;
  assign n17525 = n6543 & n12656;
  assign n17526 = ~n17524 & ~n17525;
  assign n17527 = ~n17523 & n17526;
  assign n17528 = ~n17522 & n17527;
  assign n17529 = ~pi17  & ~n17528;
  assign n17530 = pi17  & n17528;
  assign n17531 = ~n17529 & ~n17530;
  assign n17532 = n17430 & ~n17432;
  assign n17533 = ~n17433 & ~n17532;
  assign n17534 = ~n17531 & n17533;
  assign n17535 = ~n17531 & ~n17533;
  assign n17536 = n17531 & n17533;
  assign n17537 = ~n17535 & ~n17536;
  assign n17538 = n6184 & n12665;
  assign n17539 = n6527 & n12662;
  assign n17540 = n6185 & n13165;
  assign n17541 = n6543 & n12659;
  assign n17542 = ~n17540 & ~n17541;
  assign n17543 = ~n17539 & n17542;
  assign n17544 = ~n17538 & n17543;
  assign n17545 = ~pi17  & ~n17544;
  assign n17546 = pi17  & n17544;
  assign n17547 = ~n17545 & ~n17546;
  assign n17548 = ~n17425 & n17428;
  assign n17549 = n17425 & ~n17428;
  assign n17550 = ~n17548 & ~n17549;
  assign n17551 = ~n17547 & ~n17550;
  assign n17552 = n6184 & n12668;
  assign n17553 = n6527 & n12665;
  assign n17554 = n6185 & n13591;
  assign n17555 = n6543 & n12662;
  assign n17556 = ~n17554 & ~n17555;
  assign n17557 = ~n17553 & n17556;
  assign n17558 = ~n17552 & n17557;
  assign n17559 = ~pi17  & ~n17558;
  assign n17560 = pi17  & n17558;
  assign n17561 = ~n17559 & ~n17560;
  assign n17562 = ~n17420 & n17423;
  assign n17563 = n17420 & ~n17423;
  assign n17564 = ~n17562 & ~n17563;
  assign n17565 = ~n17561 & ~n17564;
  assign n17566 = n6184 & n12671;
  assign n17567 = n6527 & n12668;
  assign n17568 = n6185 & n13578;
  assign n17569 = n6543 & n12665;
  assign n17570 = ~n17568 & ~n17569;
  assign n17571 = ~n17567 & n17570;
  assign n17572 = ~n17566 & n17571;
  assign n17573 = ~pi17  & ~n17572;
  assign n17574 = pi17  & n17572;
  assign n17575 = ~n17573 & ~n17574;
  assign n17576 = ~n17415 & n17418;
  assign n17577 = n17415 & ~n17418;
  assign n17578 = ~n17576 & ~n17577;
  assign n17579 = ~n17575 & ~n17578;
  assign n17580 = n6184 & n12674;
  assign n17581 = n6527 & n12671;
  assign n17582 = n6185 & n13764;
  assign n17583 = n6543 & n12668;
  assign n17584 = ~n17582 & ~n17583;
  assign n17585 = ~n17581 & n17584;
  assign n17586 = ~n17580 & n17585;
  assign n17587 = ~pi17  & ~n17586;
  assign n17588 = pi17  & n17586;
  assign n17589 = ~n17587 & ~n17588;
  assign n17590 = ~n17410 & n17413;
  assign n17591 = n17410 & ~n17413;
  assign n17592 = ~n17590 & ~n17591;
  assign n17593 = ~n17589 & ~n17592;
  assign n17594 = n6184 & n12677;
  assign n17595 = n6527 & n12674;
  assign n17596 = n6185 & n13785;
  assign n17597 = n6543 & n12671;
  assign n17598 = ~n17596 & ~n17597;
  assign n17599 = ~n17595 & n17598;
  assign n17600 = ~n17594 & n17599;
  assign n17601 = ~pi17  & ~n17600;
  assign n17602 = pi17  & n17600;
  assign n17603 = ~n17601 & ~n17602;
  assign n17604 = n17405 & n17408;
  assign n17605 = ~n17409 & ~n17604;
  assign n17606 = ~n17603 & n17605;
  assign n17607 = ~n17603 & ~n17605;
  assign n17608 = n17603 & n17605;
  assign n17609 = ~n17607 & ~n17608;
  assign n17610 = n6184 & n12680;
  assign n17611 = n6527 & n12677;
  assign n17612 = n6185 & n14164;
  assign n17613 = n6543 & n12674;
  assign n17614 = ~n17612 & ~n17613;
  assign n17615 = ~n17611 & n17614;
  assign n17616 = ~n17610 & n17615;
  assign n17617 = ~pi17  & ~n17616;
  assign n17618 = pi17  & n17616;
  assign n17619 = ~n17617 & ~n17618;
  assign n17620 = n17400 & n17403;
  assign n17621 = ~n17404 & ~n17620;
  assign n17622 = ~n17619 & n17621;
  assign n17623 = ~n17619 & ~n17621;
  assign n17624 = n17619 & n17621;
  assign n17625 = ~n17623 & ~n17624;
  assign n17626 = n6184 & n12683;
  assign n17627 = n6527 & n12680;
  assign n17628 = n6185 & n13929;
  assign n17629 = n6543 & n12677;
  assign n17630 = ~n17628 & ~n17629;
  assign n17631 = ~n17627 & n17630;
  assign n17632 = ~n17626 & n17631;
  assign n17633 = ~pi17  & ~n17632;
  assign n17634 = pi17  & n17632;
  assign n17635 = ~n17633 & ~n17634;
  assign n17636 = n17395 & n17398;
  assign n17637 = ~n17399 & ~n17636;
  assign n17638 = ~n17635 & n17637;
  assign n17639 = ~n17635 & ~n17637;
  assign n17640 = n17635 & n17637;
  assign n17641 = ~n17639 & ~n17640;
  assign n17642 = n6184 & n12686;
  assign n17643 = n6527 & n12683;
  assign n17644 = n6185 & n14402;
  assign n17645 = n6543 & n12680;
  assign n17646 = ~n17644 & ~n17645;
  assign n17647 = ~n17643 & n17646;
  assign n17648 = ~n17642 & n17647;
  assign n17649 = ~pi17  & ~n17648;
  assign n17650 = pi17  & n17648;
  assign n17651 = ~n17649 & ~n17650;
  assign n17652 = ~n17390 & n17393;
  assign n17653 = n17390 & ~n17393;
  assign n17654 = ~n17652 & ~n17653;
  assign n17655 = ~n17651 & ~n17654;
  assign n17656 = n6184 & n12689;
  assign n17657 = n6527 & n12686;
  assign n17658 = n6185 & n14552;
  assign n17659 = n6543 & n12683;
  assign n17660 = ~n17658 & ~n17659;
  assign n17661 = ~n17657 & n17660;
  assign n17662 = ~n17656 & n17661;
  assign n17663 = ~pi17  & ~n17662;
  assign n17664 = pi17  & n17662;
  assign n17665 = ~n17663 & ~n17664;
  assign n17666 = ~n17385 & n17388;
  assign n17667 = n17385 & ~n17388;
  assign n17668 = ~n17666 & ~n17667;
  assign n17669 = ~n17665 & ~n17668;
  assign n17670 = n17206 & n17383;
  assign n17671 = ~n17384 & ~n17670;
  assign n17672 = n6184 & n12692;
  assign n17673 = n6527 & n12689;
  assign n17674 = n6185 & n14382;
  assign n17675 = n6543 & n12686;
  assign n17676 = ~n17674 & ~n17675;
  assign n17677 = ~n17673 & n17676;
  assign n17678 = ~n17672 & n17677;
  assign n17679 = pi17  & n17678;
  assign n17680 = ~pi17  & ~n17678;
  assign n17681 = ~n17679 & ~n17680;
  assign n17682 = n17671 & ~n17681;
  assign n17683 = n17379 & ~n17381;
  assign n17684 = ~n17382 & ~n17683;
  assign n17685 = n6184 & n12695;
  assign n17686 = n6527 & n12692;
  assign n17687 = n6185 & n14677;
  assign n17688 = n6543 & n12689;
  assign n17689 = ~n17687 & ~n17688;
  assign n17690 = ~n17686 & n17689;
  assign n17691 = ~n17685 & n17690;
  assign n17692 = pi17  & n17691;
  assign n17693 = ~pi17  & ~n17691;
  assign n17694 = ~n17692 & ~n17693;
  assign n17695 = n17684 & ~n17694;
  assign n17696 = n6184 & n12698;
  assign n17697 = n6527 & n12695;
  assign n17698 = n6185 & n14976;
  assign n17699 = n6543 & n12692;
  assign n17700 = ~n17698 & ~n17699;
  assign n17701 = ~n17697 & n17700;
  assign n17702 = ~n17696 & n17701;
  assign n17703 = ~pi17  & ~n17702;
  assign n17704 = pi17  & n17702;
  assign n17705 = ~n17703 & ~n17704;
  assign n17706 = n17375 & ~n17377;
  assign n17707 = ~n17378 & ~n17706;
  assign n17708 = ~n17705 & n17707;
  assign n17709 = ~n17705 & ~n17707;
  assign n17710 = n17705 & n17707;
  assign n17711 = ~n17709 & ~n17710;
  assign n17712 = n6184 & n12701;
  assign n17713 = n6527 & n12698;
  assign n17714 = n6185 & n14991;
  assign n17715 = n6543 & n12695;
  assign n17716 = ~n17714 & ~n17715;
  assign n17717 = ~n17713 & n17716;
  assign n17718 = ~n17712 & n17717;
  assign n17719 = ~pi17  & ~n17718;
  assign n17720 = pi17  & n17718;
  assign n17721 = ~n17719 & ~n17720;
  assign n17722 = n17370 & n17373;
  assign n17723 = ~n17374 & ~n17722;
  assign n17724 = ~n17721 & n17723;
  assign n17725 = ~n17721 & ~n17723;
  assign n17726 = n17721 & n17723;
  assign n17727 = ~n17725 & ~n17726;
  assign n17728 = n6184 & n12704;
  assign n17729 = n6527 & n12701;
  assign n17730 = n6185 & n14655;
  assign n17731 = n6543 & n12698;
  assign n17732 = ~n17730 & ~n17731;
  assign n17733 = ~n17729 & n17732;
  assign n17734 = ~n17728 & n17733;
  assign n17735 = ~pi17  & ~n17734;
  assign n17736 = pi17  & n17734;
  assign n17737 = ~n17735 & ~n17736;
  assign n17738 = ~n17365 & n17368;
  assign n17739 = n17365 & ~n17368;
  assign n17740 = ~n17738 & ~n17739;
  assign n17741 = ~n17737 & ~n17740;
  assign n17742 = n17275 & n17363;
  assign n17743 = ~n17364 & ~n17742;
  assign n17744 = n6184 & n12707;
  assign n17745 = n6527 & n12704;
  assign n17746 = n6185 & n15024;
  assign n17747 = n6543 & n12701;
  assign n17748 = ~n17746 & ~n17747;
  assign n17749 = ~n17745 & n17748;
  assign n17750 = ~n17744 & n17749;
  assign n17751 = pi17  & n17750;
  assign n17752 = ~pi17  & ~n17750;
  assign n17753 = ~n17751 & ~n17752;
  assign n17754 = n17743 & ~n17753;
  assign n17755 = n17359 & ~n17361;
  assign n17756 = ~n17362 & ~n17755;
  assign n17757 = n6184 & n12710;
  assign n17758 = n6527 & n12707;
  assign n17759 = n6185 & n15050;
  assign n17760 = n6543 & n12704;
  assign n17761 = ~n17759 & ~n17760;
  assign n17762 = ~n17758 & n17761;
  assign n17763 = ~n17757 & n17762;
  assign n17764 = pi17  & n17763;
  assign n17765 = ~pi17  & ~n17763;
  assign n17766 = ~n17764 & ~n17765;
  assign n17767 = n17756 & ~n17766;
  assign n17768 = n17306 & n17357;
  assign n17769 = ~n17358 & ~n17768;
  assign n17770 = n6184 & n12713;
  assign n17771 = n6527 & n12710;
  assign n17772 = n6185 & n15074;
  assign n17773 = n6543 & n12707;
  assign n17774 = ~n17772 & ~n17773;
  assign n17775 = ~n17771 & n17774;
  assign n17776 = ~n17770 & n17775;
  assign n17777 = pi17  & n17776;
  assign n17778 = ~pi17  & ~n17776;
  assign n17779 = ~n17777 & ~n17778;
  assign n17780 = n17769 & ~n17779;
  assign n17781 = n6184 & n12716;
  assign n17782 = n6527 & n12713;
  assign n17783 = n6185 & n15105;
  assign n17784 = n6543 & n12710;
  assign n17785 = ~n17783 & ~n17784;
  assign n17786 = ~n17782 & n17785;
  assign n17787 = ~n17781 & n17786;
  assign n17788 = ~pi17  & ~n17787;
  assign n17789 = pi17  & n17787;
  assign n17790 = ~n17788 & ~n17789;
  assign n17791 = n17353 & ~n17355;
  assign n17792 = ~n17356 & ~n17791;
  assign n17793 = ~n17790 & n17792;
  assign n17794 = ~n17790 & ~n17792;
  assign n17795 = n17790 & n17792;
  assign n17796 = ~n17794 & ~n17795;
  assign n17797 = n6184 & n12719;
  assign n17798 = n6527 & n12716;
  assign n17799 = n6185 & n15161;
  assign n17800 = n6543 & n12713;
  assign n17801 = ~n17799 & ~n17800;
  assign n17802 = ~n17798 & n17801;
  assign n17803 = ~n17797 & n17802;
  assign n17804 = pi17  & n17803;
  assign n17805 = ~pi17  & ~n17803;
  assign n17806 = ~n17804 & ~n17805;
  assign n17807 = n17341 & n17351;
  assign n17808 = ~n17352 & ~n17807;
  assign n17809 = ~n17806 & n17808;
  assign n17810 = n6184 & n12722;
  assign n17811 = n6527 & n12719;
  assign n17812 = n6185 & n15199;
  assign n17813 = n6543 & n12716;
  assign n17814 = ~n17812 & ~n17813;
  assign n17815 = ~n17811 & n17814;
  assign n17816 = ~n17810 & n17815;
  assign n17817 = ~pi17  & ~n17816;
  assign n17818 = pi17  & n17816;
  assign n17819 = ~n17817 & ~n17818;
  assign n17820 = pi20  & ~n17329;
  assign n17821 = n17336 & ~n17820;
  assign n17822 = ~n17336 & n17820;
  assign n17823 = ~n17821 & ~n17822;
  assign n17824 = ~n17819 & n17823;
  assign n17825 = ~n17819 & ~n17823;
  assign n17826 = n17819 & n17823;
  assign n17827 = ~n17825 & ~n17826;
  assign n17828 = n6184 & n12725;
  assign n17829 = n6527 & n12722;
  assign n17830 = n6185 & n15243;
  assign n17831 = n6543 & n12719;
  assign n17832 = ~n17830 & ~n17831;
  assign n17833 = ~n17829 & n17832;
  assign n17834 = ~n17828 & n17833;
  assign n17835 = pi17  & n17834;
  assign n17836 = ~pi17  & ~n17834;
  assign n17837 = ~n17835 & ~n17836;
  assign n17838 = pi20  & n17327;
  assign n17839 = ~n17326 & n17838;
  assign n17840 = n17326 & ~n17838;
  assign n17841 = ~n17839 & ~n17840;
  assign n17842 = ~n17837 & n17841;
  assign n17843 = n6185 & ~n15312;
  assign n17844 = n6543 & n12730;
  assign n17845 = n6527 & n12732;
  assign n17846 = ~n17844 & ~n17845;
  assign n17847 = ~n17843 & n17846;
  assign n17848 = ~n6182 & n12732;
  assign n17849 = pi17  & ~n17848;
  assign n17850 = n17847 & n17849;
  assign n17851 = n6184 & n12732;
  assign n17852 = n6527 & n12730;
  assign n17853 = n6185 & ~n15356;
  assign n17854 = n6543 & n12725;
  assign n17855 = ~n17853 & ~n17854;
  assign n17856 = ~n17852 & n17855;
  assign n17857 = ~n17851 & n17856;
  assign n17858 = n17850 & n17857;
  assign n17859 = n17327 & n17858;
  assign n17860 = ~n17327 & n17858;
  assign n17861 = n17327 & ~n17858;
  assign n17862 = ~n17860 & ~n17861;
  assign n17863 = n6184 & n12730;
  assign n17864 = n6527 & n12725;
  assign n17865 = n6185 & n15267;
  assign n17866 = n6543 & n12722;
  assign n17867 = ~n17865 & ~n17866;
  assign n17868 = ~n17864 & n17867;
  assign n17869 = ~n17863 & n17868;
  assign n17870 = pi17  & n17869;
  assign n17871 = ~pi17  & ~n17869;
  assign n17872 = ~n17870 & ~n17871;
  assign n17873 = ~n17862 & ~n17872;
  assign n17874 = ~n17859 & ~n17873;
  assign n17875 = n17837 & ~n17841;
  assign n17876 = ~n17842 & ~n17875;
  assign n17877 = ~n17874 & n17876;
  assign n17878 = ~n17842 & ~n17877;
  assign n17879 = ~n17827 & ~n17878;
  assign n17880 = ~n17824 & ~n17879;
  assign n17881 = n17806 & ~n17808;
  assign n17882 = ~n17809 & ~n17881;
  assign n17883 = ~n17880 & n17882;
  assign n17884 = ~n17809 & ~n17883;
  assign n17885 = ~n17796 & ~n17884;
  assign n17886 = ~n17793 & ~n17885;
  assign n17887 = n17769 & n17779;
  assign n17888 = ~n17769 & ~n17779;
  assign n17889 = ~n17887 & ~n17888;
  assign n17890 = ~n17886 & ~n17889;
  assign n17891 = ~n17780 & ~n17890;
  assign n17892 = n17756 & n17766;
  assign n17893 = ~n17756 & ~n17766;
  assign n17894 = ~n17892 & ~n17893;
  assign n17895 = ~n17891 & ~n17894;
  assign n17896 = ~n17767 & ~n17895;
  assign n17897 = ~n17743 & n17753;
  assign n17898 = ~n17754 & ~n17897;
  assign n17899 = ~n17896 & n17898;
  assign n17900 = ~n17754 & ~n17899;
  assign n17901 = n17737 & n17740;
  assign n17902 = ~n17741 & ~n17901;
  assign n17903 = ~n17900 & n17902;
  assign n17904 = ~n17741 & ~n17903;
  assign n17905 = ~n17727 & ~n17904;
  assign n17906 = ~n17724 & ~n17905;
  assign n17907 = ~n17711 & ~n17906;
  assign n17908 = ~n17708 & ~n17907;
  assign n17909 = n17684 & n17694;
  assign n17910 = ~n17684 & ~n17694;
  assign n17911 = ~n17909 & ~n17910;
  assign n17912 = ~n17908 & ~n17911;
  assign n17913 = ~n17695 & ~n17912;
  assign n17914 = ~n17671 & n17681;
  assign n17915 = ~n17682 & ~n17914;
  assign n17916 = ~n17913 & n17915;
  assign n17917 = ~n17682 & ~n17916;
  assign n17918 = n17665 & n17668;
  assign n17919 = ~n17669 & ~n17918;
  assign n17920 = ~n17917 & n17919;
  assign n17921 = ~n17669 & ~n17920;
  assign n17922 = n17651 & n17654;
  assign n17923 = ~n17655 & ~n17922;
  assign n17924 = ~n17921 & n17923;
  assign n17925 = ~n17655 & ~n17924;
  assign n17926 = ~n17641 & ~n17925;
  assign n17927 = ~n17638 & ~n17926;
  assign n17928 = ~n17625 & ~n17927;
  assign n17929 = ~n17622 & ~n17928;
  assign n17930 = ~n17609 & ~n17929;
  assign n17931 = ~n17606 & ~n17930;
  assign n17932 = n17589 & n17592;
  assign n17933 = ~n17593 & ~n17932;
  assign n17934 = ~n17931 & n17933;
  assign n17935 = ~n17593 & ~n17934;
  assign n17936 = n17575 & n17578;
  assign n17937 = ~n17579 & ~n17936;
  assign n17938 = ~n17935 & n17937;
  assign n17939 = ~n17579 & ~n17938;
  assign n17940 = n17561 & n17564;
  assign n17941 = ~n17565 & ~n17940;
  assign n17942 = ~n17939 & n17941;
  assign n17943 = ~n17565 & ~n17942;
  assign n17944 = n17547 & n17550;
  assign n17945 = ~n17551 & ~n17944;
  assign n17946 = ~n17943 & n17945;
  assign n17947 = ~n17551 & ~n17946;
  assign n17948 = ~n17537 & ~n17947;
  assign n17949 = ~n17534 & ~n17948;
  assign n17950 = ~n17439 & ~n17440;
  assign n17951 = ~n17450 & n17950;
  assign n17952 = n17450 & ~n17950;
  assign n17953 = ~n17951 & ~n17952;
  assign n17954 = ~n17949 & n17953;
  assign n17955 = n17949 & ~n17953;
  assign n17956 = n6835 & n12650;
  assign n17957 = n7460 & n12647;
  assign n17958 = n6836 & n13275;
  assign n17959 = n7487 & n12644;
  assign n17960 = ~n17958 & ~n17959;
  assign n17961 = ~n17957 & n17960;
  assign n17962 = ~n17956 & n17961;
  assign n17963 = pi14  & n17962;
  assign n17964 = ~pi14  & ~n17962;
  assign n17965 = ~n17963 & ~n17964;
  assign n17966 = ~n17955 & ~n17965;
  assign n17967 = ~n17954 & ~n17966;
  assign n17968 = n17521 & ~n17967;
  assign n17969 = ~n17521 & n17967;
  assign n17970 = n7654 & n12636;
  assign n17971 = n8091 & n12633;
  assign n17972 = n7648 & n13292;
  assign n17973 = n8120 & n12630;
  assign n17974 = ~n17972 & ~n17973;
  assign n17975 = ~n17971 & n17974;
  assign n17976 = ~n17970 & n17975;
  assign n17977 = pi11  & n17976;
  assign n17978 = ~pi11  & ~n17976;
  assign n17979 = ~n17977 & ~n17978;
  assign n17980 = ~n17969 & ~n17979;
  assign n17981 = ~n17968 & ~n17980;
  assign n17982 = n17517 & ~n17981;
  assign n17983 = ~n17517 & n17981;
  assign n17984 = n8474 & n12622;
  assign n17985 = n9238 & n12614;
  assign n17986 = n8468 & ~n13310;
  assign n17987 = n9265 & n12606;
  assign n17988 = ~n17986 & ~n17987;
  assign n17989 = ~n17985 & n17988;
  assign n17990 = ~n17984 & n17989;
  assign n17991 = pi8  & n17990;
  assign n17992 = ~pi8  & ~n17990;
  assign n17993 = ~n17991 & ~n17992;
  assign n17994 = ~n17983 & ~n17993;
  assign n17995 = ~n17982 & ~n17994;
  assign n17996 = ~n17513 & ~n17995;
  assign n17997 = n17513 & ~n17995;
  assign n17998 = ~n17513 & n17995;
  assign n17999 = ~n17997 & ~n17998;
  assign n18000 = n17052 & n17480;
  assign n18001 = ~n17481 & ~n18000;
  assign n18002 = ~n17999 & n18001;
  assign n18003 = ~n17996 & ~n18002;
  assign n18004 = ~n17487 & ~n17488;
  assign n18005 = ~n17498 & n18004;
  assign n18006 = n17498 & ~n18004;
  assign n18007 = ~n18005 & ~n18006;
  assign n18008 = ~n18003 & n18007;
  assign n18009 = n18003 & n18007;
  assign n18010 = ~n18003 & ~n18007;
  assign n18011 = ~n18009 & ~n18010;
  assign n18012 = n17999 & ~n18001;
  assign n18013 = ~n18002 & ~n18012;
  assign n18014 = n9719 & ~n13499;
  assign n18015 = n9725 & ~n12611;
  assign n18016 = ~n9719 & ~n9724;
  assign n18017 = ~n18015 & ~n18016;
  assign n18018 = ~n12608 & ~n18017;
  assign n18019 = ~n18014 & ~n18018;
  assign n18020 = pi5  & n18019;
  assign n18021 = ~pi5  & ~n18019;
  assign n18022 = ~n18020 & ~n18021;
  assign n18023 = ~n17968 & ~n17969;
  assign n18024 = ~n17979 & n18023;
  assign n18025 = n17979 & ~n18023;
  assign n18026 = ~n18024 & ~n18025;
  assign n18027 = n17537 & n17947;
  assign n18028 = ~n17948 & ~n18027;
  assign n18029 = n6835 & n12653;
  assign n18030 = n7460 & n12650;
  assign n18031 = n6836 & n13042;
  assign n18032 = n7487 & n12647;
  assign n18033 = ~n18031 & ~n18032;
  assign n18034 = ~n18030 & n18033;
  assign n18035 = ~n18029 & n18034;
  assign n18036 = pi14  & n18035;
  assign n18037 = ~pi14  & ~n18035;
  assign n18038 = ~n18036 & ~n18037;
  assign n18039 = n18028 & ~n18038;
  assign n18040 = n17943 & ~n17945;
  assign n18041 = ~n17946 & ~n18040;
  assign n18042 = n6835 & n12656;
  assign n18043 = n7460 & n12653;
  assign n18044 = n6836 & n12991;
  assign n18045 = n7487 & n12650;
  assign n18046 = ~n18044 & ~n18045;
  assign n18047 = ~n18043 & n18046;
  assign n18048 = ~n18042 & n18047;
  assign n18049 = pi14  & n18048;
  assign n18050 = ~pi14  & ~n18048;
  assign n18051 = ~n18049 & ~n18050;
  assign n18052 = n18041 & ~n18051;
  assign n18053 = n17939 & ~n17941;
  assign n18054 = ~n17942 & ~n18053;
  assign n18055 = n6835 & n12659;
  assign n18056 = n7460 & n12656;
  assign n18057 = n6836 & n13059;
  assign n18058 = n7487 & n12653;
  assign n18059 = ~n18057 & ~n18058;
  assign n18060 = ~n18056 & n18059;
  assign n18061 = ~n18055 & n18060;
  assign n18062 = pi14  & n18061;
  assign n18063 = ~pi14  & ~n18061;
  assign n18064 = ~n18062 & ~n18063;
  assign n18065 = n18054 & ~n18064;
  assign n18066 = n17935 & ~n17937;
  assign n18067 = ~n17938 & ~n18066;
  assign n18068 = n6835 & n12662;
  assign n18069 = n7460 & n12659;
  assign n18070 = n6836 & n13246;
  assign n18071 = n7487 & n12656;
  assign n18072 = ~n18070 & ~n18071;
  assign n18073 = ~n18069 & n18072;
  assign n18074 = ~n18068 & n18073;
  assign n18075 = pi14  & n18074;
  assign n18076 = ~pi14  & ~n18074;
  assign n18077 = ~n18075 & ~n18076;
  assign n18078 = n18067 & ~n18077;
  assign n18079 = n17931 & ~n17933;
  assign n18080 = ~n17934 & ~n18079;
  assign n18081 = n6835 & n12665;
  assign n18082 = n7460 & n12662;
  assign n18083 = n6836 & n13165;
  assign n18084 = n7487 & n12659;
  assign n18085 = ~n18083 & ~n18084;
  assign n18086 = ~n18082 & n18085;
  assign n18087 = ~n18081 & n18086;
  assign n18088 = pi14  & n18087;
  assign n18089 = ~pi14  & ~n18087;
  assign n18090 = ~n18088 & ~n18089;
  assign n18091 = n18080 & ~n18090;
  assign n18092 = n17609 & n17929;
  assign n18093 = ~n17930 & ~n18092;
  assign n18094 = n6835 & n12668;
  assign n18095 = n7460 & n12665;
  assign n18096 = n6836 & n13591;
  assign n18097 = n7487 & n12662;
  assign n18098 = ~n18096 & ~n18097;
  assign n18099 = ~n18095 & n18098;
  assign n18100 = ~n18094 & n18099;
  assign n18101 = pi14  & n18100;
  assign n18102 = ~pi14  & ~n18100;
  assign n18103 = ~n18101 & ~n18102;
  assign n18104 = n18093 & ~n18103;
  assign n18105 = n17625 & n17927;
  assign n18106 = ~n17928 & ~n18105;
  assign n18107 = n6835 & n12671;
  assign n18108 = n7460 & n12668;
  assign n18109 = n6836 & n13578;
  assign n18110 = n7487 & n12665;
  assign n18111 = ~n18109 & ~n18110;
  assign n18112 = ~n18108 & n18111;
  assign n18113 = ~n18107 & n18112;
  assign n18114 = pi14  & n18113;
  assign n18115 = ~pi14  & ~n18113;
  assign n18116 = ~n18114 & ~n18115;
  assign n18117 = n18106 & ~n18116;
  assign n18118 = n17641 & n17925;
  assign n18119 = ~n17926 & ~n18118;
  assign n18120 = n6835 & n12674;
  assign n18121 = n7460 & n12671;
  assign n18122 = n6836 & n13764;
  assign n18123 = n7487 & n12668;
  assign n18124 = ~n18122 & ~n18123;
  assign n18125 = ~n18121 & n18124;
  assign n18126 = ~n18120 & n18125;
  assign n18127 = pi14  & n18126;
  assign n18128 = ~pi14  & ~n18126;
  assign n18129 = ~n18127 & ~n18128;
  assign n18130 = n18119 & ~n18129;
  assign n18131 = n17921 & ~n17923;
  assign n18132 = ~n17924 & ~n18131;
  assign n18133 = n6835 & n12677;
  assign n18134 = n7460 & n12674;
  assign n18135 = n6836 & n13785;
  assign n18136 = n7487 & n12671;
  assign n18137 = ~n18135 & ~n18136;
  assign n18138 = ~n18134 & n18137;
  assign n18139 = ~n18133 & n18138;
  assign n18140 = pi14  & n18139;
  assign n18141 = ~pi14  & ~n18139;
  assign n18142 = ~n18140 & ~n18141;
  assign n18143 = n18132 & ~n18142;
  assign n18144 = n17917 & ~n17919;
  assign n18145 = ~n17920 & ~n18144;
  assign n18146 = n6835 & n12680;
  assign n18147 = n7460 & n12677;
  assign n18148 = n6836 & n14164;
  assign n18149 = n7487 & n12674;
  assign n18150 = ~n18148 & ~n18149;
  assign n18151 = ~n18147 & n18150;
  assign n18152 = ~n18146 & n18151;
  assign n18153 = pi14  & n18152;
  assign n18154 = ~pi14  & ~n18152;
  assign n18155 = ~n18153 & ~n18154;
  assign n18156 = n18145 & ~n18155;
  assign n18157 = n6835 & n12683;
  assign n18158 = n7460 & n12680;
  assign n18159 = n6836 & n13929;
  assign n18160 = n7487 & n12677;
  assign n18161 = ~n18159 & ~n18160;
  assign n18162 = ~n18158 & n18161;
  assign n18163 = ~n18157 & n18162;
  assign n18164 = ~pi14  & ~n18163;
  assign n18165 = pi14  & n18163;
  assign n18166 = ~n18164 & ~n18165;
  assign n18167 = n17913 & ~n17915;
  assign n18168 = ~n17916 & ~n18167;
  assign n18169 = ~n18166 & n18168;
  assign n18170 = ~n18166 & ~n18168;
  assign n18171 = n18166 & n18168;
  assign n18172 = ~n18170 & ~n18171;
  assign n18173 = n6835 & n12686;
  assign n18174 = n7460 & n12683;
  assign n18175 = n6836 & n14402;
  assign n18176 = n7487 & n12680;
  assign n18177 = ~n18175 & ~n18176;
  assign n18178 = ~n18174 & n18177;
  assign n18179 = ~n18173 & n18178;
  assign n18180 = ~pi14  & ~n18179;
  assign n18181 = pi14  & n18179;
  assign n18182 = ~n18180 & ~n18181;
  assign n18183 = n17908 & n17911;
  assign n18184 = ~n17912 & ~n18183;
  assign n18185 = ~n18182 & n18184;
  assign n18186 = ~n18182 & ~n18184;
  assign n18187 = n18182 & n18184;
  assign n18188 = ~n18186 & ~n18187;
  assign n18189 = n17711 & n17906;
  assign n18190 = ~n17907 & ~n18189;
  assign n18191 = n6835 & n12689;
  assign n18192 = n7460 & n12686;
  assign n18193 = n6836 & n14552;
  assign n18194 = n7487 & n12683;
  assign n18195 = ~n18193 & ~n18194;
  assign n18196 = ~n18192 & n18195;
  assign n18197 = ~n18191 & n18196;
  assign n18198 = pi14  & n18197;
  assign n18199 = ~pi14  & ~n18197;
  assign n18200 = ~n18198 & ~n18199;
  assign n18201 = n18190 & ~n18200;
  assign n18202 = n17727 & n17904;
  assign n18203 = ~n17905 & ~n18202;
  assign n18204 = n6835 & n12692;
  assign n18205 = n7460 & n12689;
  assign n18206 = n6836 & n14382;
  assign n18207 = n7487 & n12686;
  assign n18208 = ~n18206 & ~n18207;
  assign n18209 = ~n18205 & n18208;
  assign n18210 = ~n18204 & n18209;
  assign n18211 = pi14  & n18210;
  assign n18212 = ~pi14  & ~n18210;
  assign n18213 = ~n18211 & ~n18212;
  assign n18214 = n18203 & ~n18213;
  assign n18215 = n17900 & ~n17902;
  assign n18216 = ~n17903 & ~n18215;
  assign n18217 = n6835 & n12695;
  assign n18218 = n7460 & n12692;
  assign n18219 = n6836 & n14677;
  assign n18220 = n7487 & n12689;
  assign n18221 = ~n18219 & ~n18220;
  assign n18222 = ~n18218 & n18221;
  assign n18223 = ~n18217 & n18222;
  assign n18224 = pi14  & n18223;
  assign n18225 = ~pi14  & ~n18223;
  assign n18226 = ~n18224 & ~n18225;
  assign n18227 = n18216 & ~n18226;
  assign n18228 = n6835 & n12698;
  assign n18229 = n7460 & n12695;
  assign n18230 = n6836 & n14976;
  assign n18231 = n7487 & n12692;
  assign n18232 = ~n18230 & ~n18231;
  assign n18233 = ~n18229 & n18232;
  assign n18234 = ~n18228 & n18233;
  assign n18235 = ~pi14  & ~n18234;
  assign n18236 = pi14  & n18234;
  assign n18237 = ~n18235 & ~n18236;
  assign n18238 = n17896 & ~n17898;
  assign n18239 = ~n17899 & ~n18238;
  assign n18240 = ~n18237 & n18239;
  assign n18241 = ~n18237 & ~n18239;
  assign n18242 = n18237 & n18239;
  assign n18243 = ~n18241 & ~n18242;
  assign n18244 = n6835 & n12701;
  assign n18245 = n7460 & n12698;
  assign n18246 = n6836 & n14991;
  assign n18247 = n7487 & n12695;
  assign n18248 = ~n18246 & ~n18247;
  assign n18249 = ~n18245 & n18248;
  assign n18250 = ~n18244 & n18249;
  assign n18251 = ~pi14  & ~n18250;
  assign n18252 = pi14  & n18250;
  assign n18253 = ~n18251 & ~n18252;
  assign n18254 = n17891 & n17894;
  assign n18255 = ~n17895 & ~n18254;
  assign n18256 = ~n18253 & n18255;
  assign n18257 = ~n18253 & ~n18255;
  assign n18258 = n18253 & n18255;
  assign n18259 = ~n18257 & ~n18258;
  assign n18260 = n6835 & n12704;
  assign n18261 = n7460 & n12701;
  assign n18262 = n6836 & n14655;
  assign n18263 = n7487 & n12698;
  assign n18264 = ~n18262 & ~n18263;
  assign n18265 = ~n18261 & n18264;
  assign n18266 = ~n18260 & n18265;
  assign n18267 = ~pi14  & ~n18266;
  assign n18268 = pi14  & n18266;
  assign n18269 = ~n18267 & ~n18268;
  assign n18270 = ~n17886 & n17889;
  assign n18271 = n17886 & ~n17889;
  assign n18272 = ~n18270 & ~n18271;
  assign n18273 = ~n18269 & ~n18272;
  assign n18274 = n17796 & n17884;
  assign n18275 = ~n17885 & ~n18274;
  assign n18276 = n6835 & n12707;
  assign n18277 = n7460 & n12704;
  assign n18278 = n6836 & n15024;
  assign n18279 = n7487 & n12701;
  assign n18280 = ~n18278 & ~n18279;
  assign n18281 = ~n18277 & n18280;
  assign n18282 = ~n18276 & n18281;
  assign n18283 = pi14  & n18282;
  assign n18284 = ~pi14  & ~n18282;
  assign n18285 = ~n18283 & ~n18284;
  assign n18286 = n18275 & ~n18285;
  assign n18287 = n17880 & ~n17882;
  assign n18288 = ~n17883 & ~n18287;
  assign n18289 = n6835 & n12710;
  assign n18290 = n7460 & n12707;
  assign n18291 = n6836 & n15050;
  assign n18292 = n7487 & n12704;
  assign n18293 = ~n18291 & ~n18292;
  assign n18294 = ~n18290 & n18293;
  assign n18295 = ~n18289 & n18294;
  assign n18296 = pi14  & n18295;
  assign n18297 = ~pi14  & ~n18295;
  assign n18298 = ~n18296 & ~n18297;
  assign n18299 = n18288 & ~n18298;
  assign n18300 = n17827 & n17878;
  assign n18301 = ~n17879 & ~n18300;
  assign n18302 = n6835 & n12713;
  assign n18303 = n7460 & n12710;
  assign n18304 = n6836 & n15074;
  assign n18305 = n7487 & n12707;
  assign n18306 = ~n18304 & ~n18305;
  assign n18307 = ~n18303 & n18306;
  assign n18308 = ~n18302 & n18307;
  assign n18309 = pi14  & n18308;
  assign n18310 = ~pi14  & ~n18308;
  assign n18311 = ~n18309 & ~n18310;
  assign n18312 = n18301 & ~n18311;
  assign n18313 = n6835 & n12716;
  assign n18314 = n7460 & n12713;
  assign n18315 = n6836 & n15105;
  assign n18316 = n7487 & n12710;
  assign n18317 = ~n18315 & ~n18316;
  assign n18318 = ~n18314 & n18317;
  assign n18319 = ~n18313 & n18318;
  assign n18320 = ~pi14  & ~n18319;
  assign n18321 = pi14  & n18319;
  assign n18322 = ~n18320 & ~n18321;
  assign n18323 = n17874 & ~n17876;
  assign n18324 = ~n17877 & ~n18323;
  assign n18325 = ~n18322 & n18324;
  assign n18326 = ~n18322 & ~n18324;
  assign n18327 = n18322 & n18324;
  assign n18328 = ~n18326 & ~n18327;
  assign n18329 = n6835 & n12719;
  assign n18330 = n7460 & n12716;
  assign n18331 = n6836 & n15161;
  assign n18332 = n7487 & n12713;
  assign n18333 = ~n18331 & ~n18332;
  assign n18334 = ~n18330 & n18333;
  assign n18335 = ~n18329 & n18334;
  assign n18336 = pi14  & n18335;
  assign n18337 = ~pi14  & ~n18335;
  assign n18338 = ~n18336 & ~n18337;
  assign n18339 = n17862 & n17872;
  assign n18340 = ~n17873 & ~n18339;
  assign n18341 = ~n18338 & n18340;
  assign n18342 = n6835 & n12722;
  assign n18343 = n7460 & n12719;
  assign n18344 = n6836 & n15199;
  assign n18345 = n7487 & n12716;
  assign n18346 = ~n18344 & ~n18345;
  assign n18347 = ~n18343 & n18346;
  assign n18348 = ~n18342 & n18347;
  assign n18349 = ~pi14  & ~n18348;
  assign n18350 = pi14  & n18348;
  assign n18351 = ~n18349 & ~n18350;
  assign n18352 = pi17  & ~n17850;
  assign n18353 = n17857 & ~n18352;
  assign n18354 = ~n17857 & n18352;
  assign n18355 = ~n18353 & ~n18354;
  assign n18356 = ~n18351 & n18355;
  assign n18357 = ~n18351 & ~n18355;
  assign n18358 = n18351 & n18355;
  assign n18359 = ~n18357 & ~n18358;
  assign n18360 = n6835 & n12725;
  assign n18361 = n7460 & n12722;
  assign n18362 = n6836 & n15243;
  assign n18363 = n7487 & n12719;
  assign n18364 = ~n18362 & ~n18363;
  assign n18365 = ~n18361 & n18364;
  assign n18366 = ~n18360 & n18365;
  assign n18367 = pi14  & n18366;
  assign n18368 = ~pi14  & ~n18366;
  assign n18369 = ~n18367 & ~n18368;
  assign n18370 = pi17  & n17848;
  assign n18371 = ~n17847 & n18370;
  assign n18372 = n17847 & ~n18370;
  assign n18373 = ~n18371 & ~n18372;
  assign n18374 = ~n18369 & n18373;
  assign n18375 = n6836 & ~n15312;
  assign n18376 = n7487 & n12730;
  assign n18377 = n7460 & n12732;
  assign n18378 = ~n18376 & ~n18377;
  assign n18379 = ~n18375 & n18378;
  assign n18380 = ~n6833 & n12732;
  assign n18381 = pi14  & ~n18380;
  assign n18382 = n18379 & n18381;
  assign n18383 = n6835 & n12732;
  assign n18384 = n7460 & n12730;
  assign n18385 = n6836 & ~n15356;
  assign n18386 = n7487 & n12725;
  assign n18387 = ~n18385 & ~n18386;
  assign n18388 = ~n18384 & n18387;
  assign n18389 = ~n18383 & n18388;
  assign n18390 = n18382 & n18389;
  assign n18391 = n17848 & n18390;
  assign n18392 = ~n17848 & n18390;
  assign n18393 = n17848 & ~n18390;
  assign n18394 = ~n18392 & ~n18393;
  assign n18395 = n6835 & n12730;
  assign n18396 = n7460 & n12725;
  assign n18397 = n6836 & n15267;
  assign n18398 = n7487 & n12722;
  assign n18399 = ~n18397 & ~n18398;
  assign n18400 = ~n18396 & n18399;
  assign n18401 = ~n18395 & n18400;
  assign n18402 = pi14  & n18401;
  assign n18403 = ~pi14  & ~n18401;
  assign n18404 = ~n18402 & ~n18403;
  assign n18405 = ~n18394 & ~n18404;
  assign n18406 = ~n18391 & ~n18405;
  assign n18407 = n18369 & ~n18373;
  assign n18408 = ~n18374 & ~n18407;
  assign n18409 = ~n18406 & n18408;
  assign n18410 = ~n18374 & ~n18409;
  assign n18411 = ~n18359 & ~n18410;
  assign n18412 = ~n18356 & ~n18411;
  assign n18413 = n18338 & ~n18340;
  assign n18414 = ~n18341 & ~n18413;
  assign n18415 = ~n18412 & n18414;
  assign n18416 = ~n18341 & ~n18415;
  assign n18417 = ~n18328 & ~n18416;
  assign n18418 = ~n18325 & ~n18417;
  assign n18419 = n18301 & n18311;
  assign n18420 = ~n18301 & ~n18311;
  assign n18421 = ~n18419 & ~n18420;
  assign n18422 = ~n18418 & ~n18421;
  assign n18423 = ~n18312 & ~n18422;
  assign n18424 = n18288 & n18298;
  assign n18425 = ~n18288 & ~n18298;
  assign n18426 = ~n18424 & ~n18425;
  assign n18427 = ~n18423 & ~n18426;
  assign n18428 = ~n18299 & ~n18427;
  assign n18429 = ~n18275 & n18285;
  assign n18430 = ~n18286 & ~n18429;
  assign n18431 = ~n18428 & n18430;
  assign n18432 = ~n18286 & ~n18431;
  assign n18433 = n18269 & n18272;
  assign n18434 = ~n18273 & ~n18433;
  assign n18435 = ~n18432 & n18434;
  assign n18436 = ~n18273 & ~n18435;
  assign n18437 = ~n18259 & ~n18436;
  assign n18438 = ~n18256 & ~n18437;
  assign n18439 = ~n18243 & ~n18438;
  assign n18440 = ~n18240 & ~n18439;
  assign n18441 = n18216 & n18226;
  assign n18442 = ~n18216 & ~n18226;
  assign n18443 = ~n18441 & ~n18442;
  assign n18444 = ~n18440 & ~n18443;
  assign n18445 = ~n18227 & ~n18444;
  assign n18446 = n18203 & n18213;
  assign n18447 = ~n18203 & ~n18213;
  assign n18448 = ~n18446 & ~n18447;
  assign n18449 = ~n18445 & ~n18448;
  assign n18450 = ~n18214 & ~n18449;
  assign n18451 = ~n18190 & n18200;
  assign n18452 = ~n18201 & ~n18451;
  assign n18453 = ~n18450 & n18452;
  assign n18454 = ~n18201 & ~n18453;
  assign n18455 = ~n18188 & ~n18454;
  assign n18456 = ~n18185 & ~n18455;
  assign n18457 = ~n18172 & ~n18456;
  assign n18458 = ~n18169 & ~n18457;
  assign n18459 = n18145 & n18155;
  assign n18460 = ~n18145 & ~n18155;
  assign n18461 = ~n18459 & ~n18460;
  assign n18462 = ~n18458 & ~n18461;
  assign n18463 = ~n18156 & ~n18462;
  assign n18464 = n18132 & n18142;
  assign n18465 = ~n18132 & ~n18142;
  assign n18466 = ~n18464 & ~n18465;
  assign n18467 = ~n18463 & ~n18466;
  assign n18468 = ~n18143 & ~n18467;
  assign n18469 = n18119 & n18129;
  assign n18470 = ~n18119 & ~n18129;
  assign n18471 = ~n18469 & ~n18470;
  assign n18472 = ~n18468 & ~n18471;
  assign n18473 = ~n18130 & ~n18472;
  assign n18474 = n18106 & n18116;
  assign n18475 = ~n18106 & ~n18116;
  assign n18476 = ~n18474 & ~n18475;
  assign n18477 = ~n18473 & ~n18476;
  assign n18478 = ~n18117 & ~n18477;
  assign n18479 = n18093 & n18103;
  assign n18480 = ~n18093 & ~n18103;
  assign n18481 = ~n18479 & ~n18480;
  assign n18482 = ~n18478 & ~n18481;
  assign n18483 = ~n18104 & ~n18482;
  assign n18484 = n18080 & n18090;
  assign n18485 = ~n18080 & ~n18090;
  assign n18486 = ~n18484 & ~n18485;
  assign n18487 = ~n18483 & ~n18486;
  assign n18488 = ~n18091 & ~n18487;
  assign n18489 = n18067 & n18077;
  assign n18490 = ~n18067 & ~n18077;
  assign n18491 = ~n18489 & ~n18490;
  assign n18492 = ~n18488 & ~n18491;
  assign n18493 = ~n18078 & ~n18492;
  assign n18494 = n18054 & n18064;
  assign n18495 = ~n18054 & ~n18064;
  assign n18496 = ~n18494 & ~n18495;
  assign n18497 = ~n18493 & ~n18496;
  assign n18498 = ~n18065 & ~n18497;
  assign n18499 = n18041 & n18051;
  assign n18500 = ~n18041 & ~n18051;
  assign n18501 = ~n18499 & ~n18500;
  assign n18502 = ~n18498 & ~n18501;
  assign n18503 = ~n18052 & ~n18502;
  assign n18504 = ~n18028 & n18038;
  assign n18505 = ~n18039 & ~n18504;
  assign n18506 = ~n18503 & n18505;
  assign n18507 = ~n18039 & ~n18506;
  assign n18508 = ~n17954 & ~n17955;
  assign n18509 = ~n17965 & n18508;
  assign n18510 = n17965 & ~n18508;
  assign n18511 = ~n18509 & ~n18510;
  assign n18512 = ~n18507 & n18511;
  assign n18513 = n18507 & ~n18511;
  assign n18514 = n7654 & n12639;
  assign n18515 = n8091 & n12636;
  assign n18516 = n7648 & n13396;
  assign n18517 = n8120 & n12633;
  assign n18518 = ~n18516 & ~n18517;
  assign n18519 = ~n18515 & n18518;
  assign n18520 = ~n18514 & n18519;
  assign n18521 = pi11  & n18520;
  assign n18522 = ~pi11  & ~n18520;
  assign n18523 = ~n18521 & ~n18522;
  assign n18524 = ~n18513 & ~n18523;
  assign n18525 = ~n18512 & ~n18524;
  assign n18526 = n18026 & ~n18525;
  assign n18527 = ~n18026 & n18525;
  assign n18528 = n8474 & n12625;
  assign n18529 = n9238 & n12622;
  assign n18530 = n8468 & n13463;
  assign n18531 = n9265 & n12614;
  assign n18532 = ~n18530 & ~n18531;
  assign n18533 = ~n18529 & n18532;
  assign n18534 = ~n18528 & n18533;
  assign n18535 = pi8  & n18534;
  assign n18536 = ~pi8  & ~n18534;
  assign n18537 = ~n18535 & ~n18536;
  assign n18538 = ~n18527 & ~n18537;
  assign n18539 = ~n18526 & ~n18538;
  assign n18540 = ~n18022 & ~n18539;
  assign n18541 = n18022 & n18539;
  assign n18542 = ~n17982 & ~n17983;
  assign n18543 = ~n17993 & n18542;
  assign n18544 = n17993 & ~n18542;
  assign n18545 = ~n18543 & ~n18544;
  assign n18546 = ~n18541 & n18545;
  assign n18547 = ~n18540 & ~n18546;
  assign n18548 = n18013 & ~n18547;
  assign n18549 = ~n18540 & ~n18541;
  assign n18550 = n18545 & n18549;
  assign n18551 = ~n18545 & ~n18549;
  assign n18552 = ~n18550 & ~n18551;
  assign n18553 = ~n18526 & ~n18527;
  assign n18554 = ~n18537 & n18553;
  assign n18555 = n18537 & ~n18553;
  assign n18556 = ~n18554 & ~n18555;
  assign n18557 = n7654 & n12644;
  assign n18558 = n8091 & n12639;
  assign n18559 = n7648 & n13210;
  assign n18560 = n8120 & n12636;
  assign n18561 = ~n18559 & ~n18560;
  assign n18562 = ~n18558 & n18561;
  assign n18563 = ~n18557 & n18562;
  assign n18564 = ~pi11  & ~n18563;
  assign n18565 = pi11  & n18563;
  assign n18566 = ~n18564 & ~n18565;
  assign n18567 = n18503 & ~n18505;
  assign n18568 = ~n18506 & ~n18567;
  assign n18569 = ~n18566 & n18568;
  assign n18570 = ~n18566 & ~n18568;
  assign n18571 = n18566 & n18568;
  assign n18572 = ~n18570 & ~n18571;
  assign n18573 = n7654 & n12647;
  assign n18574 = n8091 & n12644;
  assign n18575 = n7648 & ~n13193;
  assign n18576 = n8120 & n12639;
  assign n18577 = ~n18575 & ~n18576;
  assign n18578 = ~n18574 & n18577;
  assign n18579 = ~n18573 & n18578;
  assign n18580 = ~pi11  & ~n18579;
  assign n18581 = pi11  & n18579;
  assign n18582 = ~n18580 & ~n18581;
  assign n18583 = n18498 & n18501;
  assign n18584 = ~n18502 & ~n18583;
  assign n18585 = ~n18582 & n18584;
  assign n18586 = ~n18582 & ~n18584;
  assign n18587 = n18582 & n18584;
  assign n18588 = ~n18586 & ~n18587;
  assign n18589 = n7654 & n12650;
  assign n18590 = n8091 & n12647;
  assign n18591 = n7648 & n13275;
  assign n18592 = n8120 & n12644;
  assign n18593 = ~n18591 & ~n18592;
  assign n18594 = ~n18590 & n18593;
  assign n18595 = ~n18589 & n18594;
  assign n18596 = ~pi11  & ~n18595;
  assign n18597 = pi11  & n18595;
  assign n18598 = ~n18596 & ~n18597;
  assign n18599 = n18493 & n18496;
  assign n18600 = ~n18497 & ~n18599;
  assign n18601 = ~n18598 & n18600;
  assign n18602 = ~n18598 & ~n18600;
  assign n18603 = n18598 & n18600;
  assign n18604 = ~n18602 & ~n18603;
  assign n18605 = n7654 & n12653;
  assign n18606 = n8091 & n12650;
  assign n18607 = n7648 & n13042;
  assign n18608 = n8120 & n12647;
  assign n18609 = ~n18607 & ~n18608;
  assign n18610 = ~n18606 & n18609;
  assign n18611 = ~n18605 & n18610;
  assign n18612 = ~pi11  & ~n18611;
  assign n18613 = pi11  & n18611;
  assign n18614 = ~n18612 & ~n18613;
  assign n18615 = n18488 & n18491;
  assign n18616 = ~n18492 & ~n18615;
  assign n18617 = ~n18614 & n18616;
  assign n18618 = ~n18614 & ~n18616;
  assign n18619 = n18614 & n18616;
  assign n18620 = ~n18618 & ~n18619;
  assign n18621 = n7654 & n12656;
  assign n18622 = n8091 & n12653;
  assign n18623 = n7648 & n12991;
  assign n18624 = n8120 & n12650;
  assign n18625 = ~n18623 & ~n18624;
  assign n18626 = ~n18622 & n18625;
  assign n18627 = ~n18621 & n18626;
  assign n18628 = ~pi11  & ~n18627;
  assign n18629 = pi11  & n18627;
  assign n18630 = ~n18628 & ~n18629;
  assign n18631 = n18483 & n18486;
  assign n18632 = ~n18487 & ~n18631;
  assign n18633 = ~n18630 & n18632;
  assign n18634 = ~n18630 & ~n18632;
  assign n18635 = n18630 & n18632;
  assign n18636 = ~n18634 & ~n18635;
  assign n18637 = n7654 & n12659;
  assign n18638 = n8091 & n12656;
  assign n18639 = n7648 & n13059;
  assign n18640 = n8120 & n12653;
  assign n18641 = ~n18639 & ~n18640;
  assign n18642 = ~n18638 & n18641;
  assign n18643 = ~n18637 & n18642;
  assign n18644 = ~pi11  & ~n18643;
  assign n18645 = pi11  & n18643;
  assign n18646 = ~n18644 & ~n18645;
  assign n18647 = ~n18478 & n18481;
  assign n18648 = n18478 & ~n18481;
  assign n18649 = ~n18647 & ~n18648;
  assign n18650 = ~n18646 & ~n18649;
  assign n18651 = n7654 & n12662;
  assign n18652 = n8091 & n12659;
  assign n18653 = n7648 & n13246;
  assign n18654 = n8120 & n12656;
  assign n18655 = ~n18653 & ~n18654;
  assign n18656 = ~n18652 & n18655;
  assign n18657 = ~n18651 & n18656;
  assign n18658 = ~pi11  & ~n18657;
  assign n18659 = pi11  & n18657;
  assign n18660 = ~n18658 & ~n18659;
  assign n18661 = ~n18473 & n18476;
  assign n18662 = n18473 & ~n18476;
  assign n18663 = ~n18661 & ~n18662;
  assign n18664 = ~n18660 & ~n18663;
  assign n18665 = n7654 & n12665;
  assign n18666 = n8091 & n12662;
  assign n18667 = n7648 & n13165;
  assign n18668 = n8120 & n12659;
  assign n18669 = ~n18667 & ~n18668;
  assign n18670 = ~n18666 & n18669;
  assign n18671 = ~n18665 & n18670;
  assign n18672 = ~pi11  & ~n18671;
  assign n18673 = pi11  & n18671;
  assign n18674 = ~n18672 & ~n18673;
  assign n18675 = ~n18468 & n18471;
  assign n18676 = n18468 & ~n18471;
  assign n18677 = ~n18675 & ~n18676;
  assign n18678 = ~n18674 & ~n18677;
  assign n18679 = n7654 & n12668;
  assign n18680 = n8091 & n12665;
  assign n18681 = n7648 & n13591;
  assign n18682 = n8120 & n12662;
  assign n18683 = ~n18681 & ~n18682;
  assign n18684 = ~n18680 & n18683;
  assign n18685 = ~n18679 & n18684;
  assign n18686 = ~pi11  & ~n18685;
  assign n18687 = pi11  & n18685;
  assign n18688 = ~n18686 & ~n18687;
  assign n18689 = n18463 & n18466;
  assign n18690 = ~n18467 & ~n18689;
  assign n18691 = ~n18688 & n18690;
  assign n18692 = ~n18688 & ~n18690;
  assign n18693 = n18688 & n18690;
  assign n18694 = ~n18692 & ~n18693;
  assign n18695 = n7654 & n12671;
  assign n18696 = n8091 & n12668;
  assign n18697 = n7648 & n13578;
  assign n18698 = n8120 & n12665;
  assign n18699 = ~n18697 & ~n18698;
  assign n18700 = ~n18696 & n18699;
  assign n18701 = ~n18695 & n18700;
  assign n18702 = ~pi11  & ~n18701;
  assign n18703 = pi11  & n18701;
  assign n18704 = ~n18702 & ~n18703;
  assign n18705 = n18458 & n18461;
  assign n18706 = ~n18462 & ~n18705;
  assign n18707 = ~n18704 & n18706;
  assign n18708 = ~n18704 & ~n18706;
  assign n18709 = n18704 & n18706;
  assign n18710 = ~n18708 & ~n18709;
  assign n18711 = n18172 & n18456;
  assign n18712 = ~n18457 & ~n18711;
  assign n18713 = n7654 & n12674;
  assign n18714 = n8091 & n12671;
  assign n18715 = n7648 & n13764;
  assign n18716 = n8120 & n12668;
  assign n18717 = ~n18715 & ~n18716;
  assign n18718 = ~n18714 & n18717;
  assign n18719 = ~n18713 & n18718;
  assign n18720 = pi11  & n18719;
  assign n18721 = ~pi11  & ~n18719;
  assign n18722 = ~n18720 & ~n18721;
  assign n18723 = n18712 & ~n18722;
  assign n18724 = n18188 & n18454;
  assign n18725 = ~n18455 & ~n18724;
  assign n18726 = n7654 & n12677;
  assign n18727 = n8091 & n12674;
  assign n18728 = n7648 & n13785;
  assign n18729 = n8120 & n12671;
  assign n18730 = ~n18728 & ~n18729;
  assign n18731 = ~n18727 & n18730;
  assign n18732 = ~n18726 & n18731;
  assign n18733 = pi11  & n18732;
  assign n18734 = ~pi11  & ~n18732;
  assign n18735 = ~n18733 & ~n18734;
  assign n18736 = n18725 & ~n18735;
  assign n18737 = n7654 & n12680;
  assign n18738 = n8091 & n12677;
  assign n18739 = n7648 & n14164;
  assign n18740 = n8120 & n12674;
  assign n18741 = ~n18739 & ~n18740;
  assign n18742 = ~n18738 & n18741;
  assign n18743 = ~n18737 & n18742;
  assign n18744 = ~pi11  & ~n18743;
  assign n18745 = pi11  & n18743;
  assign n18746 = ~n18744 & ~n18745;
  assign n18747 = n18450 & ~n18452;
  assign n18748 = ~n18453 & ~n18747;
  assign n18749 = ~n18746 & n18748;
  assign n18750 = ~n18746 & ~n18748;
  assign n18751 = n18746 & n18748;
  assign n18752 = ~n18750 & ~n18751;
  assign n18753 = n7654 & n12683;
  assign n18754 = n8091 & n12680;
  assign n18755 = n7648 & n13929;
  assign n18756 = n8120 & n12677;
  assign n18757 = ~n18755 & ~n18756;
  assign n18758 = ~n18754 & n18757;
  assign n18759 = ~n18753 & n18758;
  assign n18760 = ~pi11  & ~n18759;
  assign n18761 = pi11  & n18759;
  assign n18762 = ~n18760 & ~n18761;
  assign n18763 = ~n18445 & n18448;
  assign n18764 = n18445 & ~n18448;
  assign n18765 = ~n18763 & ~n18764;
  assign n18766 = ~n18762 & ~n18765;
  assign n18767 = n7654 & n12686;
  assign n18768 = n8091 & n12683;
  assign n18769 = n7648 & n14402;
  assign n18770 = n8120 & n12680;
  assign n18771 = ~n18769 & ~n18770;
  assign n18772 = ~n18768 & n18771;
  assign n18773 = ~n18767 & n18772;
  assign n18774 = ~pi11  & ~n18773;
  assign n18775 = pi11  & n18773;
  assign n18776 = ~n18774 & ~n18775;
  assign n18777 = n18440 & n18443;
  assign n18778 = ~n18444 & ~n18777;
  assign n18779 = ~n18776 & n18778;
  assign n18780 = ~n18776 & ~n18778;
  assign n18781 = n18776 & n18778;
  assign n18782 = ~n18780 & ~n18781;
  assign n18783 = n18243 & n18438;
  assign n18784 = ~n18439 & ~n18783;
  assign n18785 = n7654 & n12689;
  assign n18786 = n8091 & n12686;
  assign n18787 = n7648 & n14552;
  assign n18788 = n8120 & n12683;
  assign n18789 = ~n18787 & ~n18788;
  assign n18790 = ~n18786 & n18789;
  assign n18791 = ~n18785 & n18790;
  assign n18792 = pi11  & n18791;
  assign n18793 = ~pi11  & ~n18791;
  assign n18794 = ~n18792 & ~n18793;
  assign n18795 = n18784 & ~n18794;
  assign n18796 = n18259 & n18436;
  assign n18797 = ~n18437 & ~n18796;
  assign n18798 = n7654 & n12692;
  assign n18799 = n8091 & n12689;
  assign n18800 = n7648 & n14382;
  assign n18801 = n8120 & n12686;
  assign n18802 = ~n18800 & ~n18801;
  assign n18803 = ~n18799 & n18802;
  assign n18804 = ~n18798 & n18803;
  assign n18805 = pi11  & n18804;
  assign n18806 = ~pi11  & ~n18804;
  assign n18807 = ~n18805 & ~n18806;
  assign n18808 = n18797 & ~n18807;
  assign n18809 = n18432 & ~n18434;
  assign n18810 = ~n18435 & ~n18809;
  assign n18811 = n7654 & n12695;
  assign n18812 = n8091 & n12692;
  assign n18813 = n7648 & n14677;
  assign n18814 = n8120 & n12689;
  assign n18815 = ~n18813 & ~n18814;
  assign n18816 = ~n18812 & n18815;
  assign n18817 = ~n18811 & n18816;
  assign n18818 = pi11  & n18817;
  assign n18819 = ~pi11  & ~n18817;
  assign n18820 = ~n18818 & ~n18819;
  assign n18821 = n18810 & ~n18820;
  assign n18822 = n7654 & n12698;
  assign n18823 = n8091 & n12695;
  assign n18824 = n7648 & n14976;
  assign n18825 = n8120 & n12692;
  assign n18826 = ~n18824 & ~n18825;
  assign n18827 = ~n18823 & n18826;
  assign n18828 = ~n18822 & n18827;
  assign n18829 = ~pi11  & ~n18828;
  assign n18830 = pi11  & n18828;
  assign n18831 = ~n18829 & ~n18830;
  assign n18832 = n18428 & ~n18430;
  assign n18833 = ~n18431 & ~n18832;
  assign n18834 = ~n18831 & n18833;
  assign n18835 = ~n18831 & ~n18833;
  assign n18836 = n18831 & n18833;
  assign n18837 = ~n18835 & ~n18836;
  assign n18838 = n7654 & n12701;
  assign n18839 = n8091 & n12698;
  assign n18840 = n7648 & n14991;
  assign n18841 = n8120 & n12695;
  assign n18842 = ~n18840 & ~n18841;
  assign n18843 = ~n18839 & n18842;
  assign n18844 = ~n18838 & n18843;
  assign n18845 = ~pi11  & ~n18844;
  assign n18846 = pi11  & n18844;
  assign n18847 = ~n18845 & ~n18846;
  assign n18848 = n18423 & n18426;
  assign n18849 = ~n18427 & ~n18848;
  assign n18850 = ~n18847 & n18849;
  assign n18851 = ~n18847 & ~n18849;
  assign n18852 = n18847 & n18849;
  assign n18853 = ~n18851 & ~n18852;
  assign n18854 = n7654 & n12704;
  assign n18855 = n8091 & n12701;
  assign n18856 = n7648 & n14655;
  assign n18857 = n8120 & n12698;
  assign n18858 = ~n18856 & ~n18857;
  assign n18859 = ~n18855 & n18858;
  assign n18860 = ~n18854 & n18859;
  assign n18861 = ~pi11  & ~n18860;
  assign n18862 = pi11  & n18860;
  assign n18863 = ~n18861 & ~n18862;
  assign n18864 = ~n18418 & n18421;
  assign n18865 = n18418 & ~n18421;
  assign n18866 = ~n18864 & ~n18865;
  assign n18867 = ~n18863 & ~n18866;
  assign n18868 = n18328 & n18416;
  assign n18869 = ~n18417 & ~n18868;
  assign n18870 = n7654 & n12707;
  assign n18871 = n8091 & n12704;
  assign n18872 = n7648 & n15024;
  assign n18873 = n8120 & n12701;
  assign n18874 = ~n18872 & ~n18873;
  assign n18875 = ~n18871 & n18874;
  assign n18876 = ~n18870 & n18875;
  assign n18877 = pi11  & n18876;
  assign n18878 = ~pi11  & ~n18876;
  assign n18879 = ~n18877 & ~n18878;
  assign n18880 = n18869 & ~n18879;
  assign n18881 = n18412 & ~n18414;
  assign n18882 = ~n18415 & ~n18881;
  assign n18883 = n7654 & n12710;
  assign n18884 = n8091 & n12707;
  assign n18885 = n7648 & n15050;
  assign n18886 = n8120 & n12704;
  assign n18887 = ~n18885 & ~n18886;
  assign n18888 = ~n18884 & n18887;
  assign n18889 = ~n18883 & n18888;
  assign n18890 = pi11  & n18889;
  assign n18891 = ~pi11  & ~n18889;
  assign n18892 = ~n18890 & ~n18891;
  assign n18893 = n18882 & ~n18892;
  assign n18894 = n18359 & n18410;
  assign n18895 = ~n18411 & ~n18894;
  assign n18896 = n7654 & n12713;
  assign n18897 = n8091 & n12710;
  assign n18898 = n7648 & n15074;
  assign n18899 = n8120 & n12707;
  assign n18900 = ~n18898 & ~n18899;
  assign n18901 = ~n18897 & n18900;
  assign n18902 = ~n18896 & n18901;
  assign n18903 = pi11  & n18902;
  assign n18904 = ~pi11  & ~n18902;
  assign n18905 = ~n18903 & ~n18904;
  assign n18906 = n18895 & ~n18905;
  assign n18907 = n7654 & n12716;
  assign n18908 = n8091 & n12713;
  assign n18909 = n7648 & n15105;
  assign n18910 = n8120 & n12710;
  assign n18911 = ~n18909 & ~n18910;
  assign n18912 = ~n18908 & n18911;
  assign n18913 = ~n18907 & n18912;
  assign n18914 = ~pi11  & ~n18913;
  assign n18915 = pi11  & n18913;
  assign n18916 = ~n18914 & ~n18915;
  assign n18917 = n18406 & ~n18408;
  assign n18918 = ~n18409 & ~n18917;
  assign n18919 = ~n18916 & n18918;
  assign n18920 = ~n18916 & ~n18918;
  assign n18921 = n18916 & n18918;
  assign n18922 = ~n18920 & ~n18921;
  assign n18923 = n7654 & n12719;
  assign n18924 = n8091 & n12716;
  assign n18925 = n7648 & n15161;
  assign n18926 = n8120 & n12713;
  assign n18927 = ~n18925 & ~n18926;
  assign n18928 = ~n18924 & n18927;
  assign n18929 = ~n18923 & n18928;
  assign n18930 = pi11  & n18929;
  assign n18931 = ~pi11  & ~n18929;
  assign n18932 = ~n18930 & ~n18931;
  assign n18933 = n18394 & n18404;
  assign n18934 = ~n18405 & ~n18933;
  assign n18935 = ~n18932 & n18934;
  assign n18936 = n7654 & n12722;
  assign n18937 = n8091 & n12719;
  assign n18938 = n7648 & n15199;
  assign n18939 = n8120 & n12716;
  assign n18940 = ~n18938 & ~n18939;
  assign n18941 = ~n18937 & n18940;
  assign n18942 = ~n18936 & n18941;
  assign n18943 = ~pi11  & ~n18942;
  assign n18944 = pi11  & n18942;
  assign n18945 = ~n18943 & ~n18944;
  assign n18946 = pi14  & ~n18382;
  assign n18947 = n18389 & ~n18946;
  assign n18948 = ~n18389 & n18946;
  assign n18949 = ~n18947 & ~n18948;
  assign n18950 = ~n18945 & n18949;
  assign n18951 = ~n18945 & ~n18949;
  assign n18952 = n18945 & n18949;
  assign n18953 = ~n18951 & ~n18952;
  assign n18954 = n7654 & n12725;
  assign n18955 = n8091 & n12722;
  assign n18956 = n7648 & n15243;
  assign n18957 = n8120 & n12719;
  assign n18958 = ~n18956 & ~n18957;
  assign n18959 = ~n18955 & n18958;
  assign n18960 = ~n18954 & n18959;
  assign n18961 = pi11  & n18960;
  assign n18962 = ~pi11  & ~n18960;
  assign n18963 = ~n18961 & ~n18962;
  assign n18964 = pi14  & n18380;
  assign n18965 = ~n18379 & n18964;
  assign n18966 = n18379 & ~n18964;
  assign n18967 = ~n18965 & ~n18966;
  assign n18968 = ~n18963 & n18967;
  assign n18969 = n7648 & ~n15312;
  assign n18970 = n8120 & n12730;
  assign n18971 = n8091 & n12732;
  assign n18972 = ~n18970 & ~n18971;
  assign n18973 = ~n18969 & n18972;
  assign n18974 = ~n7644 & n12732;
  assign n18975 = pi11  & ~n18974;
  assign n18976 = n18973 & n18975;
  assign n18977 = n7654 & n12732;
  assign n18978 = n8091 & n12730;
  assign n18979 = n7648 & ~n15356;
  assign n18980 = n8120 & n12725;
  assign n18981 = ~n18979 & ~n18980;
  assign n18982 = ~n18978 & n18981;
  assign n18983 = ~n18977 & n18982;
  assign n18984 = n18976 & n18983;
  assign n18985 = n18380 & n18984;
  assign n18986 = ~n18380 & n18984;
  assign n18987 = n18380 & ~n18984;
  assign n18988 = ~n18986 & ~n18987;
  assign n18989 = n7654 & n12730;
  assign n18990 = n8091 & n12725;
  assign n18991 = n7648 & n15267;
  assign n18992 = n8120 & n12722;
  assign n18993 = ~n18991 & ~n18992;
  assign n18994 = ~n18990 & n18993;
  assign n18995 = ~n18989 & n18994;
  assign n18996 = pi11  & n18995;
  assign n18997 = ~pi11  & ~n18995;
  assign n18998 = ~n18996 & ~n18997;
  assign n18999 = ~n18988 & ~n18998;
  assign n19000 = ~n18985 & ~n18999;
  assign n19001 = n18963 & ~n18967;
  assign n19002 = ~n18968 & ~n19001;
  assign n19003 = ~n19000 & n19002;
  assign n19004 = ~n18968 & ~n19003;
  assign n19005 = ~n18953 & ~n19004;
  assign n19006 = ~n18950 & ~n19005;
  assign n19007 = n18932 & ~n18934;
  assign n19008 = ~n18935 & ~n19007;
  assign n19009 = ~n19006 & n19008;
  assign n19010 = ~n18935 & ~n19009;
  assign n19011 = ~n18922 & ~n19010;
  assign n19012 = ~n18919 & ~n19011;
  assign n19013 = n18895 & n18905;
  assign n19014 = ~n18895 & ~n18905;
  assign n19015 = ~n19013 & ~n19014;
  assign n19016 = ~n19012 & ~n19015;
  assign n19017 = ~n18906 & ~n19016;
  assign n19018 = n18882 & n18892;
  assign n19019 = ~n18882 & ~n18892;
  assign n19020 = ~n19018 & ~n19019;
  assign n19021 = ~n19017 & ~n19020;
  assign n19022 = ~n18893 & ~n19021;
  assign n19023 = ~n18869 & n18879;
  assign n19024 = ~n18880 & ~n19023;
  assign n19025 = ~n19022 & n19024;
  assign n19026 = ~n18880 & ~n19025;
  assign n19027 = n18863 & n18866;
  assign n19028 = ~n18867 & ~n19027;
  assign n19029 = ~n19026 & n19028;
  assign n19030 = ~n18867 & ~n19029;
  assign n19031 = ~n18853 & ~n19030;
  assign n19032 = ~n18850 & ~n19031;
  assign n19033 = ~n18837 & ~n19032;
  assign n19034 = ~n18834 & ~n19033;
  assign n19035 = n18810 & n18820;
  assign n19036 = ~n18810 & ~n18820;
  assign n19037 = ~n19035 & ~n19036;
  assign n19038 = ~n19034 & ~n19037;
  assign n19039 = ~n18821 & ~n19038;
  assign n19040 = n18797 & n18807;
  assign n19041 = ~n18797 & ~n18807;
  assign n19042 = ~n19040 & ~n19041;
  assign n19043 = ~n19039 & ~n19042;
  assign n19044 = ~n18808 & ~n19043;
  assign n19045 = ~n18784 & n18794;
  assign n19046 = ~n18795 & ~n19045;
  assign n19047 = ~n19044 & n19046;
  assign n19048 = ~n18795 & ~n19047;
  assign n19049 = ~n18782 & ~n19048;
  assign n19050 = ~n18779 & ~n19049;
  assign n19051 = n18762 & n18765;
  assign n19052 = ~n18766 & ~n19051;
  assign n19053 = ~n19050 & n19052;
  assign n19054 = ~n18766 & ~n19053;
  assign n19055 = ~n18752 & ~n19054;
  assign n19056 = ~n18749 & ~n19055;
  assign n19057 = n18725 & n18735;
  assign n19058 = ~n18725 & ~n18735;
  assign n19059 = ~n19057 & ~n19058;
  assign n19060 = ~n19056 & ~n19059;
  assign n19061 = ~n18736 & ~n19060;
  assign n19062 = ~n18712 & n18722;
  assign n19063 = ~n18723 & ~n19062;
  assign n19064 = ~n19061 & n19063;
  assign n19065 = ~n18723 & ~n19064;
  assign n19066 = ~n18710 & ~n19065;
  assign n19067 = ~n18707 & ~n19066;
  assign n19068 = ~n18694 & ~n19067;
  assign n19069 = ~n18691 & ~n19068;
  assign n19070 = n18674 & n18677;
  assign n19071 = ~n18678 & ~n19070;
  assign n19072 = ~n19069 & n19071;
  assign n19073 = ~n18678 & ~n19072;
  assign n19074 = n18660 & n18663;
  assign n19075 = ~n18664 & ~n19074;
  assign n19076 = ~n19073 & n19075;
  assign n19077 = ~n18664 & ~n19076;
  assign n19078 = n18646 & n18649;
  assign n19079 = ~n18650 & ~n19078;
  assign n19080 = ~n19077 & n19079;
  assign n19081 = ~n18650 & ~n19080;
  assign n19082 = ~n18636 & ~n19081;
  assign n19083 = ~n18633 & ~n19082;
  assign n19084 = ~n18620 & ~n19083;
  assign n19085 = ~n18617 & ~n19084;
  assign n19086 = ~n18604 & ~n19085;
  assign n19087 = ~n18601 & ~n19086;
  assign n19088 = ~n18588 & ~n19087;
  assign n19089 = ~n18585 & ~n19088;
  assign n19090 = ~n18572 & ~n19089;
  assign n19091 = ~n18569 & ~n19090;
  assign n19092 = ~n18512 & ~n18513;
  assign n19093 = ~n18523 & n19092;
  assign n19094 = n18523 & ~n19092;
  assign n19095 = ~n19093 & ~n19094;
  assign n19096 = ~n19091 & n19095;
  assign n19097 = n19091 & ~n19095;
  assign n19098 = n8474 & n12630;
  assign n19099 = n9238 & n12625;
  assign n19100 = n8468 & n13325;
  assign n19101 = n9265 & n12622;
  assign n19102 = ~n19100 & ~n19101;
  assign n19103 = ~n19099 & n19102;
  assign n19104 = ~n19098 & n19103;
  assign n19105 = pi8  & n19104;
  assign n19106 = ~pi8  & ~n19104;
  assign n19107 = ~n19105 & ~n19106;
  assign n19108 = ~n19097 & ~n19107;
  assign n19109 = ~n19096 & ~n19108;
  assign n19110 = n18556 & ~n19109;
  assign n19111 = ~n18556 & n19109;
  assign n19112 = n9725 & n12606;
  assign n19113 = n10702 & n12616;
  assign n19114 = n9719 & ~n13483;
  assign n19115 = n11267 & ~n12608;
  assign n19116 = ~n19114 & ~n19115;
  assign n19117 = ~n19113 & n19116;
  assign n19118 = ~n19112 & n19117;
  assign n19119 = pi5  & n19118;
  assign n19120 = ~pi5  & ~n19118;
  assign n19121 = ~n19119 & ~n19120;
  assign n19122 = ~n19111 & ~n19121;
  assign n19123 = ~n19110 & ~n19122;
  assign n19124 = n18552 & ~n19123;
  assign n19125 = ~n18552 & n19123;
  assign n19126 = ~n19124 & ~n19125;
  assign n19127 = ~n19110 & ~n19111;
  assign n19128 = ~n19121 & n19127;
  assign n19129 = n19121 & ~n19127;
  assign n19130 = ~n19128 & ~n19129;
  assign n19131 = n18572 & n19089;
  assign n19132 = ~n19090 & ~n19131;
  assign n19133 = n8474 & n12633;
  assign n19134 = n9238 & n12630;
  assign n19135 = n8468 & ~n13227;
  assign n19136 = n9265 & n12625;
  assign n19137 = ~n19135 & ~n19136;
  assign n19138 = ~n19134 & n19137;
  assign n19139 = ~n19133 & n19138;
  assign n19140 = pi8  & n19139;
  assign n19141 = ~pi8  & ~n19139;
  assign n19142 = ~n19140 & ~n19141;
  assign n19143 = n19132 & ~n19142;
  assign n19144 = n18588 & n19087;
  assign n19145 = ~n19088 & ~n19144;
  assign n19146 = n8474 & n12636;
  assign n19147 = n9238 & n12633;
  assign n19148 = n8468 & n13292;
  assign n19149 = n9265 & n12630;
  assign n19150 = ~n19148 & ~n19149;
  assign n19151 = ~n19147 & n19150;
  assign n19152 = ~n19146 & n19151;
  assign n19153 = pi8  & n19152;
  assign n19154 = ~pi8  & ~n19152;
  assign n19155 = ~n19153 & ~n19154;
  assign n19156 = n19145 & ~n19155;
  assign n19157 = n18604 & n19085;
  assign n19158 = ~n19086 & ~n19157;
  assign n19159 = n8474 & n12639;
  assign n19160 = n9238 & n12636;
  assign n19161 = n8468 & n13396;
  assign n19162 = n9265 & n12633;
  assign n19163 = ~n19161 & ~n19162;
  assign n19164 = ~n19160 & n19163;
  assign n19165 = ~n19159 & n19164;
  assign n19166 = pi8  & n19165;
  assign n19167 = ~pi8  & ~n19165;
  assign n19168 = ~n19166 & ~n19167;
  assign n19169 = n19158 & ~n19168;
  assign n19170 = n18620 & n19083;
  assign n19171 = ~n19084 & ~n19170;
  assign n19172 = n8474 & n12644;
  assign n19173 = n9238 & n12639;
  assign n19174 = n8468 & n13210;
  assign n19175 = n9265 & n12636;
  assign n19176 = ~n19174 & ~n19175;
  assign n19177 = ~n19173 & n19176;
  assign n19178 = ~n19172 & n19177;
  assign n19179 = pi8  & n19178;
  assign n19180 = ~pi8  & ~n19178;
  assign n19181 = ~n19179 & ~n19180;
  assign n19182 = n19171 & ~n19181;
  assign n19183 = n18636 & n19081;
  assign n19184 = ~n19082 & ~n19183;
  assign n19185 = n8474 & n12647;
  assign n19186 = n9238 & n12644;
  assign n19187 = n8468 & ~n13193;
  assign n19188 = n9265 & n12639;
  assign n19189 = ~n19187 & ~n19188;
  assign n19190 = ~n19186 & n19189;
  assign n19191 = ~n19185 & n19190;
  assign n19192 = pi8  & n19191;
  assign n19193 = ~pi8  & ~n19191;
  assign n19194 = ~n19192 & ~n19193;
  assign n19195 = n19184 & ~n19194;
  assign n19196 = n19077 & ~n19079;
  assign n19197 = ~n19080 & ~n19196;
  assign n19198 = n8474 & n12650;
  assign n19199 = n9238 & n12647;
  assign n19200 = n8468 & n13275;
  assign n19201 = n9265 & n12644;
  assign n19202 = ~n19200 & ~n19201;
  assign n19203 = ~n19199 & n19202;
  assign n19204 = ~n19198 & n19203;
  assign n19205 = pi8  & n19204;
  assign n19206 = ~pi8  & ~n19204;
  assign n19207 = ~n19205 & ~n19206;
  assign n19208 = n19197 & ~n19207;
  assign n19209 = n19073 & ~n19075;
  assign n19210 = ~n19076 & ~n19209;
  assign n19211 = n8474 & n12653;
  assign n19212 = n9238 & n12650;
  assign n19213 = n8468 & n13042;
  assign n19214 = n9265 & n12647;
  assign n19215 = ~n19213 & ~n19214;
  assign n19216 = ~n19212 & n19215;
  assign n19217 = ~n19211 & n19216;
  assign n19218 = pi8  & n19217;
  assign n19219 = ~pi8  & ~n19217;
  assign n19220 = ~n19218 & ~n19219;
  assign n19221 = n19210 & ~n19220;
  assign n19222 = n19069 & ~n19071;
  assign n19223 = ~n19072 & ~n19222;
  assign n19224 = n8474 & n12656;
  assign n19225 = n9238 & n12653;
  assign n19226 = n8468 & n12991;
  assign n19227 = n9265 & n12650;
  assign n19228 = ~n19226 & ~n19227;
  assign n19229 = ~n19225 & n19228;
  assign n19230 = ~n19224 & n19229;
  assign n19231 = pi8  & n19230;
  assign n19232 = ~pi8  & ~n19230;
  assign n19233 = ~n19231 & ~n19232;
  assign n19234 = n19223 & ~n19233;
  assign n19235 = n18694 & n19067;
  assign n19236 = ~n19068 & ~n19235;
  assign n19237 = n8474 & n12659;
  assign n19238 = n9238 & n12656;
  assign n19239 = n8468 & n13059;
  assign n19240 = n9265 & n12653;
  assign n19241 = ~n19239 & ~n19240;
  assign n19242 = ~n19238 & n19241;
  assign n19243 = ~n19237 & n19242;
  assign n19244 = pi8  & n19243;
  assign n19245 = ~pi8  & ~n19243;
  assign n19246 = ~n19244 & ~n19245;
  assign n19247 = n19236 & ~n19246;
  assign n19248 = n18710 & n19065;
  assign n19249 = ~n19066 & ~n19248;
  assign n19250 = n8474 & n12662;
  assign n19251 = n9238 & n12659;
  assign n19252 = n8468 & n13246;
  assign n19253 = n9265 & n12656;
  assign n19254 = ~n19252 & ~n19253;
  assign n19255 = ~n19251 & n19254;
  assign n19256 = ~n19250 & n19255;
  assign n19257 = pi8  & n19256;
  assign n19258 = ~pi8  & ~n19256;
  assign n19259 = ~n19257 & ~n19258;
  assign n19260 = n19249 & ~n19259;
  assign n19261 = n8474 & n12665;
  assign n19262 = n9238 & n12662;
  assign n19263 = n8468 & n13165;
  assign n19264 = n9265 & n12659;
  assign n19265 = ~n19263 & ~n19264;
  assign n19266 = ~n19262 & n19265;
  assign n19267 = ~n19261 & n19266;
  assign n19268 = ~pi8  & ~n19267;
  assign n19269 = pi8  & n19267;
  assign n19270 = ~n19268 & ~n19269;
  assign n19271 = n19061 & ~n19063;
  assign n19272 = ~n19064 & ~n19271;
  assign n19273 = ~n19270 & n19272;
  assign n19274 = ~n19270 & ~n19272;
  assign n19275 = n19270 & n19272;
  assign n19276 = ~n19274 & ~n19275;
  assign n19277 = n8474 & n12668;
  assign n19278 = n9238 & n12665;
  assign n19279 = n8468 & n13591;
  assign n19280 = n9265 & n12662;
  assign n19281 = ~n19279 & ~n19280;
  assign n19282 = ~n19278 & n19281;
  assign n19283 = ~n19277 & n19282;
  assign n19284 = ~pi8  & ~n19283;
  assign n19285 = pi8  & n19283;
  assign n19286 = ~n19284 & ~n19285;
  assign n19287 = ~n19056 & n19059;
  assign n19288 = n19056 & ~n19059;
  assign n19289 = ~n19287 & ~n19288;
  assign n19290 = ~n19286 & ~n19289;
  assign n19291 = n18752 & n19054;
  assign n19292 = ~n19055 & ~n19291;
  assign n19293 = n8474 & n12671;
  assign n19294 = n9238 & n12668;
  assign n19295 = n8468 & n13578;
  assign n19296 = n9265 & n12665;
  assign n19297 = ~n19295 & ~n19296;
  assign n19298 = ~n19294 & n19297;
  assign n19299 = ~n19293 & n19298;
  assign n19300 = pi8  & n19299;
  assign n19301 = ~pi8  & ~n19299;
  assign n19302 = ~n19300 & ~n19301;
  assign n19303 = n19292 & ~n19302;
  assign n19304 = n19050 & ~n19052;
  assign n19305 = ~n19053 & ~n19304;
  assign n19306 = n8474 & n12674;
  assign n19307 = n9238 & n12671;
  assign n19308 = n8468 & n13764;
  assign n19309 = n9265 & n12668;
  assign n19310 = ~n19308 & ~n19309;
  assign n19311 = ~n19307 & n19310;
  assign n19312 = ~n19306 & n19311;
  assign n19313 = pi8  & n19312;
  assign n19314 = ~pi8  & ~n19312;
  assign n19315 = ~n19313 & ~n19314;
  assign n19316 = n19305 & ~n19315;
  assign n19317 = n18782 & n19048;
  assign n19318 = ~n19049 & ~n19317;
  assign n19319 = n8474 & n12677;
  assign n19320 = n9238 & n12674;
  assign n19321 = n8468 & n13785;
  assign n19322 = n9265 & n12671;
  assign n19323 = ~n19321 & ~n19322;
  assign n19324 = ~n19320 & n19323;
  assign n19325 = ~n19319 & n19324;
  assign n19326 = pi8  & n19325;
  assign n19327 = ~pi8  & ~n19325;
  assign n19328 = ~n19326 & ~n19327;
  assign n19329 = n19318 & ~n19328;
  assign n19330 = n8474 & n12680;
  assign n19331 = n9238 & n12677;
  assign n19332 = n8468 & n14164;
  assign n19333 = n9265 & n12674;
  assign n19334 = ~n19332 & ~n19333;
  assign n19335 = ~n19331 & n19334;
  assign n19336 = ~n19330 & n19335;
  assign n19337 = ~pi8  & ~n19336;
  assign n19338 = pi8  & n19336;
  assign n19339 = ~n19337 & ~n19338;
  assign n19340 = n19044 & ~n19046;
  assign n19341 = ~n19047 & ~n19340;
  assign n19342 = ~n19339 & n19341;
  assign n19343 = ~n19339 & ~n19341;
  assign n19344 = n19339 & n19341;
  assign n19345 = ~n19343 & ~n19344;
  assign n19346 = n8474 & n12683;
  assign n19347 = n9238 & n12680;
  assign n19348 = n8468 & n13929;
  assign n19349 = n9265 & n12677;
  assign n19350 = ~n19348 & ~n19349;
  assign n19351 = ~n19347 & n19350;
  assign n19352 = ~n19346 & n19351;
  assign n19353 = ~pi8  & ~n19352;
  assign n19354 = pi8  & n19352;
  assign n19355 = ~n19353 & ~n19354;
  assign n19356 = ~n19039 & n19042;
  assign n19357 = n19039 & ~n19042;
  assign n19358 = ~n19356 & ~n19357;
  assign n19359 = ~n19355 & ~n19358;
  assign n19360 = n8474 & n12686;
  assign n19361 = n9238 & n12683;
  assign n19362 = n8468 & n14402;
  assign n19363 = n9265 & n12680;
  assign n19364 = ~n19362 & ~n19363;
  assign n19365 = ~n19361 & n19364;
  assign n19366 = ~n19360 & n19365;
  assign n19367 = ~pi8  & ~n19366;
  assign n19368 = pi8  & n19366;
  assign n19369 = ~n19367 & ~n19368;
  assign n19370 = n19034 & n19037;
  assign n19371 = ~n19038 & ~n19370;
  assign n19372 = ~n19369 & n19371;
  assign n19373 = ~n19369 & ~n19371;
  assign n19374 = n19369 & n19371;
  assign n19375 = ~n19373 & ~n19374;
  assign n19376 = n18837 & n19032;
  assign n19377 = ~n19033 & ~n19376;
  assign n19378 = n8474 & n12689;
  assign n19379 = n9238 & n12686;
  assign n19380 = n8468 & n14552;
  assign n19381 = n9265 & n12683;
  assign n19382 = ~n19380 & ~n19381;
  assign n19383 = ~n19379 & n19382;
  assign n19384 = ~n19378 & n19383;
  assign n19385 = pi8  & n19384;
  assign n19386 = ~pi8  & ~n19384;
  assign n19387 = ~n19385 & ~n19386;
  assign n19388 = n19377 & ~n19387;
  assign n19389 = n18853 & n19030;
  assign n19390 = ~n19031 & ~n19389;
  assign n19391 = n8474 & n12692;
  assign n19392 = n9238 & n12689;
  assign n19393 = n8468 & n14382;
  assign n19394 = n9265 & n12686;
  assign n19395 = ~n19393 & ~n19394;
  assign n19396 = ~n19392 & n19395;
  assign n19397 = ~n19391 & n19396;
  assign n19398 = pi8  & n19397;
  assign n19399 = ~pi8  & ~n19397;
  assign n19400 = ~n19398 & ~n19399;
  assign n19401 = n19390 & ~n19400;
  assign n19402 = n19026 & ~n19028;
  assign n19403 = ~n19029 & ~n19402;
  assign n19404 = n8474 & n12695;
  assign n19405 = n9238 & n12692;
  assign n19406 = n8468 & n14677;
  assign n19407 = n9265 & n12689;
  assign n19408 = ~n19406 & ~n19407;
  assign n19409 = ~n19405 & n19408;
  assign n19410 = ~n19404 & n19409;
  assign n19411 = pi8  & n19410;
  assign n19412 = ~pi8  & ~n19410;
  assign n19413 = ~n19411 & ~n19412;
  assign n19414 = n19403 & ~n19413;
  assign n19415 = n8474 & n12698;
  assign n19416 = n9238 & n12695;
  assign n19417 = n8468 & n14976;
  assign n19418 = n9265 & n12692;
  assign n19419 = ~n19417 & ~n19418;
  assign n19420 = ~n19416 & n19419;
  assign n19421 = ~n19415 & n19420;
  assign n19422 = ~pi8  & ~n19421;
  assign n19423 = pi8  & n19421;
  assign n19424 = ~n19422 & ~n19423;
  assign n19425 = n19022 & ~n19024;
  assign n19426 = ~n19025 & ~n19425;
  assign n19427 = ~n19424 & n19426;
  assign n19428 = ~n19424 & ~n19426;
  assign n19429 = n19424 & n19426;
  assign n19430 = ~n19428 & ~n19429;
  assign n19431 = n8474 & n12701;
  assign n19432 = n9238 & n12698;
  assign n19433 = n8468 & n14991;
  assign n19434 = n9265 & n12695;
  assign n19435 = ~n19433 & ~n19434;
  assign n19436 = ~n19432 & n19435;
  assign n19437 = ~n19431 & n19436;
  assign n19438 = ~pi8  & ~n19437;
  assign n19439 = pi8  & n19437;
  assign n19440 = ~n19438 & ~n19439;
  assign n19441 = n19017 & n19020;
  assign n19442 = ~n19021 & ~n19441;
  assign n19443 = ~n19440 & n19442;
  assign n19444 = ~n19440 & ~n19442;
  assign n19445 = n19440 & n19442;
  assign n19446 = ~n19444 & ~n19445;
  assign n19447 = n8474 & n12704;
  assign n19448 = n9238 & n12701;
  assign n19449 = n8468 & n14655;
  assign n19450 = n9265 & n12698;
  assign n19451 = ~n19449 & ~n19450;
  assign n19452 = ~n19448 & n19451;
  assign n19453 = ~n19447 & n19452;
  assign n19454 = ~pi8  & ~n19453;
  assign n19455 = pi8  & n19453;
  assign n19456 = ~n19454 & ~n19455;
  assign n19457 = ~n19012 & n19015;
  assign n19458 = n19012 & ~n19015;
  assign n19459 = ~n19457 & ~n19458;
  assign n19460 = ~n19456 & ~n19459;
  assign n19461 = n18922 & n19010;
  assign n19462 = ~n19011 & ~n19461;
  assign n19463 = n8474 & n12707;
  assign n19464 = n9238 & n12704;
  assign n19465 = n8468 & n15024;
  assign n19466 = n9265 & n12701;
  assign n19467 = ~n19465 & ~n19466;
  assign n19468 = ~n19464 & n19467;
  assign n19469 = ~n19463 & n19468;
  assign n19470 = pi8  & n19469;
  assign n19471 = ~pi8  & ~n19469;
  assign n19472 = ~n19470 & ~n19471;
  assign n19473 = n19462 & ~n19472;
  assign n19474 = n19006 & ~n19008;
  assign n19475 = ~n19009 & ~n19474;
  assign n19476 = n8474 & n12710;
  assign n19477 = n9238 & n12707;
  assign n19478 = n8468 & n15050;
  assign n19479 = n9265 & n12704;
  assign n19480 = ~n19478 & ~n19479;
  assign n19481 = ~n19477 & n19480;
  assign n19482 = ~n19476 & n19481;
  assign n19483 = pi8  & n19482;
  assign n19484 = ~pi8  & ~n19482;
  assign n19485 = ~n19483 & ~n19484;
  assign n19486 = n19475 & ~n19485;
  assign n19487 = n18953 & n19004;
  assign n19488 = ~n19005 & ~n19487;
  assign n19489 = n8474 & n12713;
  assign n19490 = n9238 & n12710;
  assign n19491 = n8468 & n15074;
  assign n19492 = n9265 & n12707;
  assign n19493 = ~n19491 & ~n19492;
  assign n19494 = ~n19490 & n19493;
  assign n19495 = ~n19489 & n19494;
  assign n19496 = pi8  & n19495;
  assign n19497 = ~pi8  & ~n19495;
  assign n19498 = ~n19496 & ~n19497;
  assign n19499 = n19488 & ~n19498;
  assign n19500 = n8474 & n12716;
  assign n19501 = n9238 & n12713;
  assign n19502 = n8468 & n15105;
  assign n19503 = n9265 & n12710;
  assign n19504 = ~n19502 & ~n19503;
  assign n19505 = ~n19501 & n19504;
  assign n19506 = ~n19500 & n19505;
  assign n19507 = ~pi8  & ~n19506;
  assign n19508 = pi8  & n19506;
  assign n19509 = ~n19507 & ~n19508;
  assign n19510 = n19000 & ~n19002;
  assign n19511 = ~n19003 & ~n19510;
  assign n19512 = ~n19509 & n19511;
  assign n19513 = ~n19509 & ~n19511;
  assign n19514 = n19509 & n19511;
  assign n19515 = ~n19513 & ~n19514;
  assign n19516 = n8474 & n12719;
  assign n19517 = n9238 & n12716;
  assign n19518 = n8468 & n15161;
  assign n19519 = n9265 & n12713;
  assign n19520 = ~n19518 & ~n19519;
  assign n19521 = ~n19517 & n19520;
  assign n19522 = ~n19516 & n19521;
  assign n19523 = pi8  & n19522;
  assign n19524 = ~pi8  & ~n19522;
  assign n19525 = ~n19523 & ~n19524;
  assign n19526 = n18988 & n18998;
  assign n19527 = ~n18999 & ~n19526;
  assign n19528 = ~n19525 & n19527;
  assign n19529 = n8474 & n12722;
  assign n19530 = n9238 & n12719;
  assign n19531 = n8468 & n15199;
  assign n19532 = n9265 & n12716;
  assign n19533 = ~n19531 & ~n19532;
  assign n19534 = ~n19530 & n19533;
  assign n19535 = ~n19529 & n19534;
  assign n19536 = ~pi8  & ~n19535;
  assign n19537 = pi8  & n19535;
  assign n19538 = ~n19536 & ~n19537;
  assign n19539 = pi11  & ~n18976;
  assign n19540 = n18983 & ~n19539;
  assign n19541 = ~n18983 & n19539;
  assign n19542 = ~n19540 & ~n19541;
  assign n19543 = ~n19538 & n19542;
  assign n19544 = ~n19538 & ~n19542;
  assign n19545 = n19538 & n19542;
  assign n19546 = ~n19544 & ~n19545;
  assign n19547 = n8474 & n12725;
  assign n19548 = n9238 & n12722;
  assign n19549 = n8468 & n15243;
  assign n19550 = n9265 & n12719;
  assign n19551 = ~n19549 & ~n19550;
  assign n19552 = ~n19548 & n19551;
  assign n19553 = ~n19547 & n19552;
  assign n19554 = pi8  & n19553;
  assign n19555 = ~pi8  & ~n19553;
  assign n19556 = ~n19554 & ~n19555;
  assign n19557 = pi11  & n18974;
  assign n19558 = ~n18973 & n19557;
  assign n19559 = n18973 & ~n19557;
  assign n19560 = ~n19558 & ~n19559;
  assign n19561 = ~n19556 & n19560;
  assign n19562 = n8468 & ~n15312;
  assign n19563 = n9265 & n12730;
  assign n19564 = n9238 & n12732;
  assign n19565 = ~n19563 & ~n19564;
  assign n19566 = ~n19562 & n19565;
  assign n19567 = ~n8464 & n12732;
  assign n19568 = pi8  & ~n19567;
  assign n19569 = n19566 & n19568;
  assign n19570 = n8474 & n12732;
  assign n19571 = n9238 & n12730;
  assign n19572 = n8468 & ~n15356;
  assign n19573 = n9265 & n12725;
  assign n19574 = ~n19572 & ~n19573;
  assign n19575 = ~n19571 & n19574;
  assign n19576 = ~n19570 & n19575;
  assign n19577 = n19569 & n19576;
  assign n19578 = n18974 & n19577;
  assign n19579 = ~n18974 & n19577;
  assign n19580 = n18974 & ~n19577;
  assign n19581 = ~n19579 & ~n19580;
  assign n19582 = n8474 & n12730;
  assign n19583 = n9238 & n12725;
  assign n19584 = n8468 & n15267;
  assign n19585 = n9265 & n12722;
  assign n19586 = ~n19584 & ~n19585;
  assign n19587 = ~n19583 & n19586;
  assign n19588 = ~n19582 & n19587;
  assign n19589 = pi8  & n19588;
  assign n19590 = ~pi8  & ~n19588;
  assign n19591 = ~n19589 & ~n19590;
  assign n19592 = ~n19581 & ~n19591;
  assign n19593 = ~n19578 & ~n19592;
  assign n19594 = n19556 & ~n19560;
  assign n19595 = ~n19561 & ~n19594;
  assign n19596 = ~n19593 & n19595;
  assign n19597 = ~n19561 & ~n19596;
  assign n19598 = ~n19546 & ~n19597;
  assign n19599 = ~n19543 & ~n19598;
  assign n19600 = n19525 & ~n19527;
  assign n19601 = ~n19528 & ~n19600;
  assign n19602 = ~n19599 & n19601;
  assign n19603 = ~n19528 & ~n19602;
  assign n19604 = ~n19515 & ~n19603;
  assign n19605 = ~n19512 & ~n19604;
  assign n19606 = n19488 & n19498;
  assign n19607 = ~n19488 & ~n19498;
  assign n19608 = ~n19606 & ~n19607;
  assign n19609 = ~n19605 & ~n19608;
  assign n19610 = ~n19499 & ~n19609;
  assign n19611 = n19475 & n19485;
  assign n19612 = ~n19475 & ~n19485;
  assign n19613 = ~n19611 & ~n19612;
  assign n19614 = ~n19610 & ~n19613;
  assign n19615 = ~n19486 & ~n19614;
  assign n19616 = ~n19462 & n19472;
  assign n19617 = ~n19473 & ~n19616;
  assign n19618 = ~n19615 & n19617;
  assign n19619 = ~n19473 & ~n19618;
  assign n19620 = n19456 & n19459;
  assign n19621 = ~n19460 & ~n19620;
  assign n19622 = ~n19619 & n19621;
  assign n19623 = ~n19460 & ~n19622;
  assign n19624 = ~n19446 & ~n19623;
  assign n19625 = ~n19443 & ~n19624;
  assign n19626 = ~n19430 & ~n19625;
  assign n19627 = ~n19427 & ~n19626;
  assign n19628 = n19403 & n19413;
  assign n19629 = ~n19403 & ~n19413;
  assign n19630 = ~n19628 & ~n19629;
  assign n19631 = ~n19627 & ~n19630;
  assign n19632 = ~n19414 & ~n19631;
  assign n19633 = n19390 & n19400;
  assign n19634 = ~n19390 & ~n19400;
  assign n19635 = ~n19633 & ~n19634;
  assign n19636 = ~n19632 & ~n19635;
  assign n19637 = ~n19401 & ~n19636;
  assign n19638 = ~n19377 & n19387;
  assign n19639 = ~n19388 & ~n19638;
  assign n19640 = ~n19637 & n19639;
  assign n19641 = ~n19388 & ~n19640;
  assign n19642 = ~n19375 & ~n19641;
  assign n19643 = ~n19372 & ~n19642;
  assign n19644 = n19355 & n19358;
  assign n19645 = ~n19359 & ~n19644;
  assign n19646 = ~n19643 & n19645;
  assign n19647 = ~n19359 & ~n19646;
  assign n19648 = ~n19345 & ~n19647;
  assign n19649 = ~n19342 & ~n19648;
  assign n19650 = n19318 & n19328;
  assign n19651 = ~n19318 & ~n19328;
  assign n19652 = ~n19650 & ~n19651;
  assign n19653 = ~n19649 & ~n19652;
  assign n19654 = ~n19329 & ~n19653;
  assign n19655 = n19305 & n19315;
  assign n19656 = ~n19305 & ~n19315;
  assign n19657 = ~n19655 & ~n19656;
  assign n19658 = ~n19654 & ~n19657;
  assign n19659 = ~n19316 & ~n19658;
  assign n19660 = ~n19292 & n19302;
  assign n19661 = ~n19303 & ~n19660;
  assign n19662 = ~n19659 & n19661;
  assign n19663 = ~n19303 & ~n19662;
  assign n19664 = n19286 & n19289;
  assign n19665 = ~n19290 & ~n19664;
  assign n19666 = ~n19663 & n19665;
  assign n19667 = ~n19290 & ~n19666;
  assign n19668 = ~n19276 & ~n19667;
  assign n19669 = ~n19273 & ~n19668;
  assign n19670 = n19249 & n19259;
  assign n19671 = ~n19249 & ~n19259;
  assign n19672 = ~n19670 & ~n19671;
  assign n19673 = ~n19669 & ~n19672;
  assign n19674 = ~n19260 & ~n19673;
  assign n19675 = n19236 & n19246;
  assign n19676 = ~n19236 & ~n19246;
  assign n19677 = ~n19675 & ~n19676;
  assign n19678 = ~n19674 & ~n19677;
  assign n19679 = ~n19247 & ~n19678;
  assign n19680 = n19223 & n19233;
  assign n19681 = ~n19223 & ~n19233;
  assign n19682 = ~n19680 & ~n19681;
  assign n19683 = ~n19679 & ~n19682;
  assign n19684 = ~n19234 & ~n19683;
  assign n19685 = n19210 & n19220;
  assign n19686 = ~n19210 & ~n19220;
  assign n19687 = ~n19685 & ~n19686;
  assign n19688 = ~n19684 & ~n19687;
  assign n19689 = ~n19221 & ~n19688;
  assign n19690 = n19197 & n19207;
  assign n19691 = ~n19197 & ~n19207;
  assign n19692 = ~n19690 & ~n19691;
  assign n19693 = ~n19689 & ~n19692;
  assign n19694 = ~n19208 & ~n19693;
  assign n19695 = n19184 & n19194;
  assign n19696 = ~n19184 & ~n19194;
  assign n19697 = ~n19695 & ~n19696;
  assign n19698 = ~n19694 & ~n19697;
  assign n19699 = ~n19195 & ~n19698;
  assign n19700 = n19171 & n19181;
  assign n19701 = ~n19171 & ~n19181;
  assign n19702 = ~n19700 & ~n19701;
  assign n19703 = ~n19699 & ~n19702;
  assign n19704 = ~n19182 & ~n19703;
  assign n19705 = n19158 & n19168;
  assign n19706 = ~n19158 & ~n19168;
  assign n19707 = ~n19705 & ~n19706;
  assign n19708 = ~n19704 & ~n19707;
  assign n19709 = ~n19169 & ~n19708;
  assign n19710 = n19145 & n19155;
  assign n19711 = ~n19145 & ~n19155;
  assign n19712 = ~n19710 & ~n19711;
  assign n19713 = ~n19709 & ~n19712;
  assign n19714 = ~n19156 & ~n19713;
  assign n19715 = ~n19132 & n19142;
  assign n19716 = ~n19143 & ~n19715;
  assign n19717 = ~n19714 & n19716;
  assign n19718 = ~n19143 & ~n19717;
  assign n19719 = ~n19096 & ~n19097;
  assign n19720 = ~n19107 & n19719;
  assign n19721 = n19107 & ~n19719;
  assign n19722 = ~n19720 & ~n19721;
  assign n19723 = ~n19718 & n19722;
  assign n19724 = n19718 & ~n19722;
  assign n19725 = n10702 & n12606;
  assign n19726 = ~n12611 & n19115;
  assign n19727 = n9725 & n12614;
  assign n19728 = n9719 & n12868;
  assign n19729 = ~n19727 & ~n19728;
  assign n19730 = ~n19726 & n19729;
  assign n19731 = ~n19725 & n19730;
  assign n19732 = pi5  & n19731;
  assign n19733 = ~pi5  & ~n19731;
  assign n19734 = ~n19732 & ~n19733;
  assign n19735 = ~n19724 & ~n19734;
  assign n19736 = ~n19723 & ~n19735;
  assign n19737 = n19130 & ~n19736;
  assign n19738 = ~n19130 & n19736;
  assign n19739 = ~n19737 & ~n19738;
  assign n19740 = n9725 & n12622;
  assign n19741 = n10702 & n12614;
  assign n19742 = n9719 & ~n13310;
  assign n19743 = n11267 & n12606;
  assign n19744 = ~n19742 & ~n19743;
  assign n19745 = ~n19741 & n19744;
  assign n19746 = ~n19740 & n19745;
  assign n19747 = ~pi5  & ~n19746;
  assign n19748 = pi5  & n19746;
  assign n19749 = ~n19747 & ~n19748;
  assign n19750 = n19714 & ~n19716;
  assign n19751 = ~n19717 & ~n19750;
  assign n19752 = ~n19749 & n19751;
  assign n19753 = ~n19749 & ~n19751;
  assign n19754 = n19749 & n19751;
  assign n19755 = ~n19753 & ~n19754;
  assign n19756 = n11289 & ~n13499;
  assign n19757 = ~n11287 & ~n11289;
  assign n19758 = n11288 & ~n12611;
  assign n19759 = ~n19757 & ~n19758;
  assign n19760 = ~n12608 & ~n19759;
  assign n19761 = ~n19756 & ~n19760;
  assign n19762 = pi2  & n19761;
  assign n19763 = ~pi2  & ~n19761;
  assign n19764 = ~n19762 & ~n19763;
  assign n19765 = ~n19755 & ~n19764;
  assign n19766 = ~n19752 & ~n19765;
  assign n19767 = ~n19723 & ~n19724;
  assign n19768 = ~n19734 & n19767;
  assign n19769 = n19734 & ~n19767;
  assign n19770 = ~n19768 & ~n19769;
  assign n19771 = ~n19766 & n19770;
  assign n19772 = n19766 & ~n19770;
  assign n19773 = ~n19771 & ~n19772;
  assign n19774 = n9725 & n12625;
  assign n19775 = n10702 & n12622;
  assign n19776 = n9719 & n13463;
  assign n19777 = n11267 & n12614;
  assign n19778 = ~n19776 & ~n19777;
  assign n19779 = ~n19775 & n19778;
  assign n19780 = ~n19774 & n19779;
  assign n19781 = ~pi5  & ~n19780;
  assign n19782 = pi5  & n19780;
  assign n19783 = ~n19781 & ~n19782;
  assign n19784 = ~n19709 & n19712;
  assign n19785 = n19709 & ~n19712;
  assign n19786 = ~n19784 & ~n19785;
  assign n19787 = ~n19783 & ~n19786;
  assign n19788 = n9725 & n12630;
  assign n19789 = n10702 & n12625;
  assign n19790 = n9719 & n13325;
  assign n19791 = n11267 & n12622;
  assign n19792 = ~n19790 & ~n19791;
  assign n19793 = ~n19789 & n19792;
  assign n19794 = ~n19788 & n19793;
  assign n19795 = ~pi5  & ~n19794;
  assign n19796 = pi5  & n19794;
  assign n19797 = ~n19795 & ~n19796;
  assign n19798 = ~n19704 & n19707;
  assign n19799 = n19704 & ~n19707;
  assign n19800 = ~n19798 & ~n19799;
  assign n19801 = ~n19797 & ~n19800;
  assign n19802 = n9725 & n12633;
  assign n19803 = n10702 & n12630;
  assign n19804 = n9719 & ~n13227;
  assign n19805 = n11267 & n12625;
  assign n19806 = ~n19804 & ~n19805;
  assign n19807 = ~n19803 & n19806;
  assign n19808 = ~n19802 & n19807;
  assign n19809 = ~pi5  & ~n19808;
  assign n19810 = pi5  & n19808;
  assign n19811 = ~n19809 & ~n19810;
  assign n19812 = ~n19699 & n19702;
  assign n19813 = n19699 & ~n19702;
  assign n19814 = ~n19812 & ~n19813;
  assign n19815 = ~n19811 & ~n19814;
  assign n19816 = n9725 & n12636;
  assign n19817 = n10702 & n12633;
  assign n19818 = n9719 & n13292;
  assign n19819 = n11267 & n12630;
  assign n19820 = ~n19818 & ~n19819;
  assign n19821 = ~n19817 & n19820;
  assign n19822 = ~n19816 & n19821;
  assign n19823 = ~pi5  & ~n19822;
  assign n19824 = pi5  & n19822;
  assign n19825 = ~n19823 & ~n19824;
  assign n19826 = ~n19694 & n19697;
  assign n19827 = n19694 & ~n19697;
  assign n19828 = ~n19826 & ~n19827;
  assign n19829 = ~n19825 & ~n19828;
  assign n19830 = n9725 & n12639;
  assign n19831 = n10702 & n12636;
  assign n19832 = n9719 & n13396;
  assign n19833 = n11267 & n12633;
  assign n19834 = ~n19832 & ~n19833;
  assign n19835 = ~n19831 & n19834;
  assign n19836 = ~n19830 & n19835;
  assign n19837 = ~pi5  & ~n19836;
  assign n19838 = pi5  & n19836;
  assign n19839 = ~n19837 & ~n19838;
  assign n19840 = n19689 & n19692;
  assign n19841 = ~n19693 & ~n19840;
  assign n19842 = ~n19839 & n19841;
  assign n19843 = ~n19839 & ~n19841;
  assign n19844 = n19839 & n19841;
  assign n19845 = ~n19843 & ~n19844;
  assign n19846 = n9725 & n12644;
  assign n19847 = n10702 & n12639;
  assign n19848 = n9719 & n13210;
  assign n19849 = n11267 & n12636;
  assign n19850 = ~n19848 & ~n19849;
  assign n19851 = ~n19847 & n19850;
  assign n19852 = ~n19846 & n19851;
  assign n19853 = ~pi5  & ~n19852;
  assign n19854 = pi5  & n19852;
  assign n19855 = ~n19853 & ~n19854;
  assign n19856 = n19684 & n19687;
  assign n19857 = ~n19688 & ~n19856;
  assign n19858 = ~n19855 & n19857;
  assign n19859 = ~n19855 & ~n19857;
  assign n19860 = n19855 & n19857;
  assign n19861 = ~n19859 & ~n19860;
  assign n19862 = n9725 & n12647;
  assign n19863 = n10702 & n12644;
  assign n19864 = n9719 & ~n13193;
  assign n19865 = n11267 & n12639;
  assign n19866 = ~n19864 & ~n19865;
  assign n19867 = ~n19863 & n19866;
  assign n19868 = ~n19862 & n19867;
  assign n19869 = ~pi5  & ~n19868;
  assign n19870 = pi5  & n19868;
  assign n19871 = ~n19869 & ~n19870;
  assign n19872 = n19679 & n19682;
  assign n19873 = ~n19683 & ~n19872;
  assign n19874 = ~n19871 & n19873;
  assign n19875 = ~n19871 & ~n19873;
  assign n19876 = n19871 & n19873;
  assign n19877 = ~n19875 & ~n19876;
  assign n19878 = n9725 & n12650;
  assign n19879 = n10702 & n12647;
  assign n19880 = n9719 & n13275;
  assign n19881 = n11267 & n12644;
  assign n19882 = ~n19880 & ~n19881;
  assign n19883 = ~n19879 & n19882;
  assign n19884 = ~n19878 & n19883;
  assign n19885 = ~pi5  & ~n19884;
  assign n19886 = pi5  & n19884;
  assign n19887 = ~n19885 & ~n19886;
  assign n19888 = ~n19674 & n19677;
  assign n19889 = n19674 & ~n19677;
  assign n19890 = ~n19888 & ~n19889;
  assign n19891 = ~n19887 & ~n19890;
  assign n19892 = n9725 & n12653;
  assign n19893 = n10702 & n12650;
  assign n19894 = n9719 & n13042;
  assign n19895 = n11267 & n12647;
  assign n19896 = ~n19894 & ~n19895;
  assign n19897 = ~n19893 & n19896;
  assign n19898 = ~n19892 & n19897;
  assign n19899 = ~pi5  & ~n19898;
  assign n19900 = pi5  & n19898;
  assign n19901 = ~n19899 & ~n19900;
  assign n19902 = ~n19669 & n19672;
  assign n19903 = n19669 & ~n19672;
  assign n19904 = ~n19902 & ~n19903;
  assign n19905 = ~n19901 & ~n19904;
  assign n19906 = n19276 & n19667;
  assign n19907 = ~n19668 & ~n19906;
  assign n19908 = n9725 & n12656;
  assign n19909 = n10702 & n12653;
  assign n19910 = n9719 & n12991;
  assign n19911 = n11267 & n12650;
  assign n19912 = ~n19910 & ~n19911;
  assign n19913 = ~n19909 & n19912;
  assign n19914 = ~n19908 & n19913;
  assign n19915 = pi5  & n19914;
  assign n19916 = ~pi5  & ~n19914;
  assign n19917 = ~n19915 & ~n19916;
  assign n19918 = n19907 & ~n19917;
  assign n19919 = n19663 & ~n19665;
  assign n19920 = ~n19666 & ~n19919;
  assign n19921 = n9725 & n12659;
  assign n19922 = n10702 & n12656;
  assign n19923 = n9719 & n13059;
  assign n19924 = n11267 & n12653;
  assign n19925 = ~n19923 & ~n19924;
  assign n19926 = ~n19922 & n19925;
  assign n19927 = ~n19921 & n19926;
  assign n19928 = pi5  & n19927;
  assign n19929 = ~pi5  & ~n19927;
  assign n19930 = ~n19928 & ~n19929;
  assign n19931 = n19920 & ~n19930;
  assign n19932 = n9725 & n12662;
  assign n19933 = n10702 & n12659;
  assign n19934 = n9719 & n13246;
  assign n19935 = n11267 & n12656;
  assign n19936 = ~n19934 & ~n19935;
  assign n19937 = ~n19933 & n19936;
  assign n19938 = ~n19932 & n19937;
  assign n19939 = ~pi5  & ~n19938;
  assign n19940 = pi5  & n19938;
  assign n19941 = ~n19939 & ~n19940;
  assign n19942 = n19659 & ~n19661;
  assign n19943 = ~n19662 & ~n19942;
  assign n19944 = ~n19941 & n19943;
  assign n19945 = ~n19941 & ~n19943;
  assign n19946 = n19941 & n19943;
  assign n19947 = ~n19945 & ~n19946;
  assign n19948 = n9725 & n12665;
  assign n19949 = n10702 & n12662;
  assign n19950 = n9719 & n13165;
  assign n19951 = n11267 & n12659;
  assign n19952 = ~n19950 & ~n19951;
  assign n19953 = ~n19949 & n19952;
  assign n19954 = ~n19948 & n19953;
  assign n19955 = ~pi5  & ~n19954;
  assign n19956 = pi5  & n19954;
  assign n19957 = ~n19955 & ~n19956;
  assign n19958 = n19654 & n19657;
  assign n19959 = ~n19658 & ~n19958;
  assign n19960 = ~n19957 & n19959;
  assign n19961 = ~n19957 & ~n19959;
  assign n19962 = n19957 & n19959;
  assign n19963 = ~n19961 & ~n19962;
  assign n19964 = n9725 & n12668;
  assign n19965 = n10702 & n12665;
  assign n19966 = n9719 & n13591;
  assign n19967 = n11267 & n12662;
  assign n19968 = ~n19966 & ~n19967;
  assign n19969 = ~n19965 & n19968;
  assign n19970 = ~n19964 & n19969;
  assign n19971 = ~pi5  & ~n19970;
  assign n19972 = pi5  & n19970;
  assign n19973 = ~n19971 & ~n19972;
  assign n19974 = ~n19649 & n19652;
  assign n19975 = n19649 & ~n19652;
  assign n19976 = ~n19974 & ~n19975;
  assign n19977 = ~n19973 & ~n19976;
  assign n19978 = n19345 & n19647;
  assign n19979 = ~n19648 & ~n19978;
  assign n19980 = n9725 & n12671;
  assign n19981 = n10702 & n12668;
  assign n19982 = n9719 & n13578;
  assign n19983 = n11267 & n12665;
  assign n19984 = ~n19982 & ~n19983;
  assign n19985 = ~n19981 & n19984;
  assign n19986 = ~n19980 & n19985;
  assign n19987 = pi5  & n19986;
  assign n19988 = ~pi5  & ~n19986;
  assign n19989 = ~n19987 & ~n19988;
  assign n19990 = n19979 & ~n19989;
  assign n19991 = n19643 & ~n19645;
  assign n19992 = ~n19646 & ~n19991;
  assign n19993 = n9725 & n12674;
  assign n19994 = n10702 & n12671;
  assign n19995 = n9719 & n13764;
  assign n19996 = n11267 & n12668;
  assign n19997 = ~n19995 & ~n19996;
  assign n19998 = ~n19994 & n19997;
  assign n19999 = ~n19993 & n19998;
  assign n20000 = pi5  & n19999;
  assign n20001 = ~pi5  & ~n19999;
  assign n20002 = ~n20000 & ~n20001;
  assign n20003 = n19992 & ~n20002;
  assign n20004 = n19375 & n19641;
  assign n20005 = ~n19642 & ~n20004;
  assign n20006 = n9725 & n12677;
  assign n20007 = n10702 & n12674;
  assign n20008 = n9719 & n13785;
  assign n20009 = n11267 & n12671;
  assign n20010 = ~n20008 & ~n20009;
  assign n20011 = ~n20007 & n20010;
  assign n20012 = ~n20006 & n20011;
  assign n20013 = pi5  & n20012;
  assign n20014 = ~pi5  & ~n20012;
  assign n20015 = ~n20013 & ~n20014;
  assign n20016 = n20005 & ~n20015;
  assign n20017 = n9725 & n12680;
  assign n20018 = n10702 & n12677;
  assign n20019 = n9719 & n14164;
  assign n20020 = n11267 & n12674;
  assign n20021 = ~n20019 & ~n20020;
  assign n20022 = ~n20018 & n20021;
  assign n20023 = ~n20017 & n20022;
  assign n20024 = ~pi5  & ~n20023;
  assign n20025 = pi5  & n20023;
  assign n20026 = ~n20024 & ~n20025;
  assign n20027 = n19637 & ~n19639;
  assign n20028 = ~n19640 & ~n20027;
  assign n20029 = ~n20026 & n20028;
  assign n20030 = ~n20026 & ~n20028;
  assign n20031 = n20026 & n20028;
  assign n20032 = ~n20030 & ~n20031;
  assign n20033 = n9725 & n12683;
  assign n20034 = n10702 & n12680;
  assign n20035 = n9719 & n13929;
  assign n20036 = n11267 & n12677;
  assign n20037 = ~n20035 & ~n20036;
  assign n20038 = ~n20034 & n20037;
  assign n20039 = ~n20033 & n20038;
  assign n20040 = ~pi5  & ~n20039;
  assign n20041 = pi5  & n20039;
  assign n20042 = ~n20040 & ~n20041;
  assign n20043 = ~n19632 & n19635;
  assign n20044 = n19632 & ~n19635;
  assign n20045 = ~n20043 & ~n20044;
  assign n20046 = ~n20042 & ~n20045;
  assign n20047 = n9725 & n12686;
  assign n20048 = n10702 & n12683;
  assign n20049 = n9719 & n14402;
  assign n20050 = n11267 & n12680;
  assign n20051 = ~n20049 & ~n20050;
  assign n20052 = ~n20048 & n20051;
  assign n20053 = ~n20047 & n20052;
  assign n20054 = ~pi5  & ~n20053;
  assign n20055 = pi5  & n20053;
  assign n20056 = ~n20054 & ~n20055;
  assign n20057 = n19627 & n19630;
  assign n20058 = ~n19631 & ~n20057;
  assign n20059 = ~n20056 & n20058;
  assign n20060 = ~n20056 & ~n20058;
  assign n20061 = n20056 & n20058;
  assign n20062 = ~n20060 & ~n20061;
  assign n20063 = n19430 & n19625;
  assign n20064 = ~n19626 & ~n20063;
  assign n20065 = n9725 & n12689;
  assign n20066 = n10702 & n12686;
  assign n20067 = n9719 & n14552;
  assign n20068 = n11267 & n12683;
  assign n20069 = ~n20067 & ~n20068;
  assign n20070 = ~n20066 & n20069;
  assign n20071 = ~n20065 & n20070;
  assign n20072 = pi5  & n20071;
  assign n20073 = ~pi5  & ~n20071;
  assign n20074 = ~n20072 & ~n20073;
  assign n20075 = n20064 & ~n20074;
  assign n20076 = n19446 & n19623;
  assign n20077 = ~n19624 & ~n20076;
  assign n20078 = n9725 & n12692;
  assign n20079 = n10702 & n12689;
  assign n20080 = n9719 & n14382;
  assign n20081 = n11267 & n12686;
  assign n20082 = ~n20080 & ~n20081;
  assign n20083 = ~n20079 & n20082;
  assign n20084 = ~n20078 & n20083;
  assign n20085 = pi5  & n20084;
  assign n20086 = ~pi5  & ~n20084;
  assign n20087 = ~n20085 & ~n20086;
  assign n20088 = n20077 & ~n20087;
  assign n20089 = n19619 & ~n19621;
  assign n20090 = ~n19622 & ~n20089;
  assign n20091 = n9725 & n12695;
  assign n20092 = n10702 & n12692;
  assign n20093 = n9719 & n14677;
  assign n20094 = n11267 & n12689;
  assign n20095 = ~n20093 & ~n20094;
  assign n20096 = ~n20092 & n20095;
  assign n20097 = ~n20091 & n20096;
  assign n20098 = pi5  & n20097;
  assign n20099 = ~pi5  & ~n20097;
  assign n20100 = ~n20098 & ~n20099;
  assign n20101 = n20090 & ~n20100;
  assign n20102 = n9725 & n12698;
  assign n20103 = n10702 & n12695;
  assign n20104 = n9719 & n14976;
  assign n20105 = n11267 & n12692;
  assign n20106 = ~n20104 & ~n20105;
  assign n20107 = ~n20103 & n20106;
  assign n20108 = ~n20102 & n20107;
  assign n20109 = ~pi5  & ~n20108;
  assign n20110 = pi5  & n20108;
  assign n20111 = ~n20109 & ~n20110;
  assign n20112 = n19615 & ~n19617;
  assign n20113 = ~n19618 & ~n20112;
  assign n20114 = ~n20111 & n20113;
  assign n20115 = ~n20111 & ~n20113;
  assign n20116 = n20111 & n20113;
  assign n20117 = ~n20115 & ~n20116;
  assign n20118 = n9725 & n12701;
  assign n20119 = n10702 & n12698;
  assign n20120 = n9719 & n14991;
  assign n20121 = n11267 & n12695;
  assign n20122 = ~n20120 & ~n20121;
  assign n20123 = ~n20119 & n20122;
  assign n20124 = ~n20118 & n20123;
  assign n20125 = ~pi5  & ~n20124;
  assign n20126 = pi5  & n20124;
  assign n20127 = ~n20125 & ~n20126;
  assign n20128 = n19610 & n19613;
  assign n20129 = ~n19614 & ~n20128;
  assign n20130 = ~n20127 & n20129;
  assign n20131 = ~n20127 & ~n20129;
  assign n20132 = n20127 & n20129;
  assign n20133 = ~n20131 & ~n20132;
  assign n20134 = n9725 & n12704;
  assign n20135 = n10702 & n12701;
  assign n20136 = n9719 & n14655;
  assign n20137 = n11267 & n12698;
  assign n20138 = ~n20136 & ~n20137;
  assign n20139 = ~n20135 & n20138;
  assign n20140 = ~n20134 & n20139;
  assign n20141 = ~pi5  & ~n20140;
  assign n20142 = pi5  & n20140;
  assign n20143 = ~n20141 & ~n20142;
  assign n20144 = ~n19605 & n19608;
  assign n20145 = n19605 & ~n19608;
  assign n20146 = ~n20144 & ~n20145;
  assign n20147 = ~n20143 & ~n20146;
  assign n20148 = n19515 & n19603;
  assign n20149 = ~n19604 & ~n20148;
  assign n20150 = n9725 & n12707;
  assign n20151 = n10702 & n12704;
  assign n20152 = n9719 & n15024;
  assign n20153 = n11267 & n12701;
  assign n20154 = ~n20152 & ~n20153;
  assign n20155 = ~n20151 & n20154;
  assign n20156 = ~n20150 & n20155;
  assign n20157 = pi5  & n20156;
  assign n20158 = ~pi5  & ~n20156;
  assign n20159 = ~n20157 & ~n20158;
  assign n20160 = n20149 & ~n20159;
  assign n20161 = n19599 & ~n19601;
  assign n20162 = ~n19602 & ~n20161;
  assign n20163 = n9725 & n12710;
  assign n20164 = n10702 & n12707;
  assign n20165 = n9719 & n15050;
  assign n20166 = n11267 & n12704;
  assign n20167 = ~n20165 & ~n20166;
  assign n20168 = ~n20164 & n20167;
  assign n20169 = ~n20163 & n20168;
  assign n20170 = pi5  & n20169;
  assign n20171 = ~pi5  & ~n20169;
  assign n20172 = ~n20170 & ~n20171;
  assign n20173 = n20162 & ~n20172;
  assign n20174 = n19546 & n19597;
  assign n20175 = ~n19598 & ~n20174;
  assign n20176 = n9725 & n12713;
  assign n20177 = n10702 & n12710;
  assign n20178 = n9719 & n15074;
  assign n20179 = n11267 & n12707;
  assign n20180 = ~n20178 & ~n20179;
  assign n20181 = ~n20177 & n20180;
  assign n20182 = ~n20176 & n20181;
  assign n20183 = pi5  & n20182;
  assign n20184 = ~pi5  & ~n20182;
  assign n20185 = ~n20183 & ~n20184;
  assign n20186 = n20175 & ~n20185;
  assign n20187 = n9725 & n12716;
  assign n20188 = n10702 & n12713;
  assign n20189 = n9719 & n15105;
  assign n20190 = n11267 & n12710;
  assign n20191 = ~n20189 & ~n20190;
  assign n20192 = ~n20188 & n20191;
  assign n20193 = ~n20187 & n20192;
  assign n20194 = ~pi5  & ~n20193;
  assign n20195 = pi5  & n20193;
  assign n20196 = ~n20194 & ~n20195;
  assign n20197 = n19593 & ~n19595;
  assign n20198 = ~n19596 & ~n20197;
  assign n20199 = ~n20196 & n20198;
  assign n20200 = ~n20196 & ~n20198;
  assign n20201 = n20196 & n20198;
  assign n20202 = ~n20200 & ~n20201;
  assign n20203 = n9725 & n12719;
  assign n20204 = n10702 & n12716;
  assign n20205 = n9719 & n15161;
  assign n20206 = n11267 & n12713;
  assign n20207 = ~n20205 & ~n20206;
  assign n20208 = ~n20204 & n20207;
  assign n20209 = ~n20203 & n20208;
  assign n20210 = pi5  & n20209;
  assign n20211 = ~pi5  & ~n20209;
  assign n20212 = ~n20210 & ~n20211;
  assign n20213 = n19581 & n19591;
  assign n20214 = ~n19592 & ~n20213;
  assign n20215 = ~n20212 & n20214;
  assign n20216 = n9725 & n12722;
  assign n20217 = n10702 & n12719;
  assign n20218 = n9719 & n15199;
  assign n20219 = n11267 & n12716;
  assign n20220 = ~n20218 & ~n20219;
  assign n20221 = ~n20217 & n20220;
  assign n20222 = ~n20216 & n20221;
  assign n20223 = ~pi5  & ~n20222;
  assign n20224 = pi5  & n20222;
  assign n20225 = ~n20223 & ~n20224;
  assign n20226 = pi8  & ~n19569;
  assign n20227 = n19576 & ~n20226;
  assign n20228 = ~n19576 & n20226;
  assign n20229 = ~n20227 & ~n20228;
  assign n20230 = ~n20225 & n20229;
  assign n20231 = ~n20225 & ~n20229;
  assign n20232 = n20225 & n20229;
  assign n20233 = ~n20231 & ~n20232;
  assign n20234 = n9725 & n12725;
  assign n20235 = n10702 & n12722;
  assign n20236 = n9719 & n15243;
  assign n20237 = n11267 & n12719;
  assign n20238 = ~n20236 & ~n20237;
  assign n20239 = ~n20235 & n20238;
  assign n20240 = ~n20234 & n20239;
  assign n20241 = pi5  & n20240;
  assign n20242 = ~pi5  & ~n20240;
  assign n20243 = ~n20241 & ~n20242;
  assign n20244 = pi8  & n19567;
  assign n20245 = ~n19566 & n20244;
  assign n20246 = n19566 & ~n20244;
  assign n20247 = ~n20245 & ~n20246;
  assign n20248 = ~n20243 & n20247;
  assign n20249 = n9719 & ~n15312;
  assign n20250 = n11267 & n12730;
  assign n20251 = n10702 & n12732;
  assign n20252 = ~n20250 & ~n20251;
  assign n20253 = ~n20249 & n20252;
  assign n20254 = ~n9715 & n12732;
  assign n20255 = pi5  & ~n20254;
  assign n20256 = n20253 & n20255;
  assign n20257 = n9725 & n12732;
  assign n20258 = n10702 & n12730;
  assign n20259 = n9719 & ~n15356;
  assign n20260 = n11267 & n12725;
  assign n20261 = ~n20259 & ~n20260;
  assign n20262 = ~n20258 & n20261;
  assign n20263 = ~n20257 & n20262;
  assign n20264 = n20256 & n20263;
  assign n20265 = n19567 & n20264;
  assign n20266 = ~n19567 & n20264;
  assign n20267 = n19567 & ~n20264;
  assign n20268 = ~n20266 & ~n20267;
  assign n20269 = n9725 & n12730;
  assign n20270 = n10702 & n12725;
  assign n20271 = n9719 & n15267;
  assign n20272 = n11267 & n12722;
  assign n20273 = ~n20271 & ~n20272;
  assign n20274 = ~n20270 & n20273;
  assign n20275 = ~n20269 & n20274;
  assign n20276 = pi5  & n20275;
  assign n20277 = ~pi5  & ~n20275;
  assign n20278 = ~n20276 & ~n20277;
  assign n20279 = ~n20268 & ~n20278;
  assign n20280 = ~n20265 & ~n20279;
  assign n20281 = n20243 & ~n20247;
  assign n20282 = ~n20248 & ~n20281;
  assign n20283 = ~n20280 & n20282;
  assign n20284 = ~n20248 & ~n20283;
  assign n20285 = ~n20233 & ~n20284;
  assign n20286 = ~n20230 & ~n20285;
  assign n20287 = n20212 & ~n20214;
  assign n20288 = ~n20215 & ~n20287;
  assign n20289 = ~n20286 & n20288;
  assign n20290 = ~n20215 & ~n20289;
  assign n20291 = ~n20202 & ~n20290;
  assign n20292 = ~n20199 & ~n20291;
  assign n20293 = n20175 & n20185;
  assign n20294 = ~n20175 & ~n20185;
  assign n20295 = ~n20293 & ~n20294;
  assign n20296 = ~n20292 & ~n20295;
  assign n20297 = ~n20186 & ~n20296;
  assign n20298 = n20162 & n20172;
  assign n20299 = ~n20162 & ~n20172;
  assign n20300 = ~n20298 & ~n20299;
  assign n20301 = ~n20297 & ~n20300;
  assign n20302 = ~n20173 & ~n20301;
  assign n20303 = ~n20149 & n20159;
  assign n20304 = ~n20160 & ~n20303;
  assign n20305 = ~n20302 & n20304;
  assign n20306 = ~n20160 & ~n20305;
  assign n20307 = n20143 & n20146;
  assign n20308 = ~n20147 & ~n20307;
  assign n20309 = ~n20306 & n20308;
  assign n20310 = ~n20147 & ~n20309;
  assign n20311 = ~n20133 & ~n20310;
  assign n20312 = ~n20130 & ~n20311;
  assign n20313 = ~n20117 & ~n20312;
  assign n20314 = ~n20114 & ~n20313;
  assign n20315 = n20090 & n20100;
  assign n20316 = ~n20090 & ~n20100;
  assign n20317 = ~n20315 & ~n20316;
  assign n20318 = ~n20314 & ~n20317;
  assign n20319 = ~n20101 & ~n20318;
  assign n20320 = n20077 & n20087;
  assign n20321 = ~n20077 & ~n20087;
  assign n20322 = ~n20320 & ~n20321;
  assign n20323 = ~n20319 & ~n20322;
  assign n20324 = ~n20088 & ~n20323;
  assign n20325 = ~n20064 & n20074;
  assign n20326 = ~n20075 & ~n20325;
  assign n20327 = ~n20324 & n20326;
  assign n20328 = ~n20075 & ~n20327;
  assign n20329 = ~n20062 & ~n20328;
  assign n20330 = ~n20059 & ~n20329;
  assign n20331 = n20042 & n20045;
  assign n20332 = ~n20046 & ~n20331;
  assign n20333 = ~n20330 & n20332;
  assign n20334 = ~n20046 & ~n20333;
  assign n20335 = ~n20032 & ~n20334;
  assign n20336 = ~n20029 & ~n20335;
  assign n20337 = n20005 & n20015;
  assign n20338 = ~n20005 & ~n20015;
  assign n20339 = ~n20337 & ~n20338;
  assign n20340 = ~n20336 & ~n20339;
  assign n20341 = ~n20016 & ~n20340;
  assign n20342 = n19992 & n20002;
  assign n20343 = ~n19992 & ~n20002;
  assign n20344 = ~n20342 & ~n20343;
  assign n20345 = ~n20341 & ~n20344;
  assign n20346 = ~n20003 & ~n20345;
  assign n20347 = ~n19979 & n19989;
  assign n20348 = ~n19990 & ~n20347;
  assign n20349 = ~n20346 & n20348;
  assign n20350 = ~n19990 & ~n20349;
  assign n20351 = n19973 & n19976;
  assign n20352 = ~n19977 & ~n20351;
  assign n20353 = ~n20350 & n20352;
  assign n20354 = ~n19977 & ~n20353;
  assign n20355 = ~n19963 & ~n20354;
  assign n20356 = ~n19960 & ~n20355;
  assign n20357 = ~n19947 & ~n20356;
  assign n20358 = ~n19944 & ~n20357;
  assign n20359 = n19920 & n19930;
  assign n20360 = ~n19920 & ~n19930;
  assign n20361 = ~n20359 & ~n20360;
  assign n20362 = ~n20358 & ~n20361;
  assign n20363 = ~n19931 & ~n20362;
  assign n20364 = ~n19907 & n19917;
  assign n20365 = ~n19918 & ~n20364;
  assign n20366 = ~n20363 & n20365;
  assign n20367 = ~n19918 & ~n20366;
  assign n20368 = n19901 & n19904;
  assign n20369 = ~n19905 & ~n20368;
  assign n20370 = ~n20367 & n20369;
  assign n20371 = ~n19905 & ~n20370;
  assign n20372 = n19887 & n19890;
  assign n20373 = ~n19891 & ~n20372;
  assign n20374 = ~n20371 & n20373;
  assign n20375 = ~n19891 & ~n20374;
  assign n20376 = ~n19877 & ~n20375;
  assign n20377 = ~n19874 & ~n20376;
  assign n20378 = ~n19861 & ~n20377;
  assign n20379 = ~n19858 & ~n20378;
  assign n20380 = ~n19845 & ~n20379;
  assign n20381 = ~n19842 & ~n20380;
  assign n20382 = n19825 & n19828;
  assign n20383 = ~n19829 & ~n20382;
  assign n20384 = ~n20381 & n20383;
  assign n20385 = ~n19829 & ~n20384;
  assign n20386 = n19811 & n19814;
  assign n20387 = ~n19815 & ~n20386;
  assign n20388 = ~n20385 & n20387;
  assign n20389 = ~n19815 & ~n20388;
  assign n20390 = n19797 & n19800;
  assign n20391 = ~n19801 & ~n20390;
  assign n20392 = ~n20389 & n20391;
  assign n20393 = ~n19801 & ~n20392;
  assign n20394 = n19783 & n19786;
  assign n20395 = ~n19787 & ~n20394;
  assign n20396 = ~n20393 & n20395;
  assign n20397 = ~n19787 & ~n20396;
  assign n20398 = n19755 & n19764;
  assign n20399 = ~n19765 & ~n20398;
  assign n20400 = ~n20397 & n20399;
  assign n20401 = n20397 & ~n20399;
  assign n20402 = ~n20400 & ~n20401;
  assign n20403 = n20393 & ~n20395;
  assign n20404 = ~n20396 & ~n20403;
  assign n20405 = n11288 & n12606;
  assign n20406 = n11894 & n12616;
  assign n20407 = n11289 & ~n13483;
  assign n20408 = n11908 & ~n12608;
  assign n20409 = ~n20407 & ~n20408;
  assign n20410 = ~n20406 & n20409;
  assign n20411 = ~n20405 & n20410;
  assign n20412 = pi2  & n20411;
  assign n20413 = ~pi2  & ~n20411;
  assign n20414 = ~n20412 & ~n20413;
  assign n20415 = n20404 & ~n20414;
  assign n20416 = n20389 & ~n20391;
  assign n20417 = ~n20392 & ~n20416;
  assign n20418 = n11894 & n12606;
  assign n20419 = ~n12611 & n20408;
  assign n20420 = n11288 & n12614;
  assign n20421 = n11289 & n12868;
  assign n20422 = ~n20420 & ~n20421;
  assign n20423 = ~n20419 & n20422;
  assign n20424 = ~n20418 & n20423;
  assign n20425 = pi2  & n20424;
  assign n20426 = ~pi2  & ~n20424;
  assign n20427 = ~n20425 & ~n20426;
  assign n20428 = n20417 & ~n20427;
  assign n20429 = n20385 & ~n20387;
  assign n20430 = ~n20388 & ~n20429;
  assign n20431 = n11288 & n12622;
  assign n20432 = n11894 & n12614;
  assign n20433 = n11289 & ~n13310;
  assign n20434 = n11908 & n12606;
  assign n20435 = ~n20433 & ~n20434;
  assign n20436 = ~n20432 & n20435;
  assign n20437 = ~n20431 & n20436;
  assign n20438 = pi2  & n20437;
  assign n20439 = ~pi2  & ~n20437;
  assign n20440 = ~n20438 & ~n20439;
  assign n20441 = n20430 & ~n20440;
  assign n20442 = n20381 & ~n20383;
  assign n20443 = ~n20384 & ~n20442;
  assign n20444 = n11288 & n12625;
  assign n20445 = n11894 & n12622;
  assign n20446 = n11289 & n13463;
  assign n20447 = n11908 & n12614;
  assign n20448 = ~n20446 & ~n20447;
  assign n20449 = ~n20445 & n20448;
  assign n20450 = ~n20444 & n20449;
  assign n20451 = pi2  & n20450;
  assign n20452 = ~pi2  & ~n20450;
  assign n20453 = ~n20451 & ~n20452;
  assign n20454 = n20443 & ~n20453;
  assign n20455 = n19845 & n20379;
  assign n20456 = ~n20380 & ~n20455;
  assign n20457 = n11288 & n12630;
  assign n20458 = n11894 & n12625;
  assign n20459 = n11289 & n13325;
  assign n20460 = n11908 & n12622;
  assign n20461 = ~n20459 & ~n20460;
  assign n20462 = ~n20458 & n20461;
  assign n20463 = ~n20457 & n20462;
  assign n20464 = pi2  & n20463;
  assign n20465 = ~pi2  & ~n20463;
  assign n20466 = ~n20464 & ~n20465;
  assign n20467 = n20456 & ~n20466;
  assign n20468 = n19861 & n20377;
  assign n20469 = ~n20378 & ~n20468;
  assign n20470 = n11288 & n12633;
  assign n20471 = n11894 & n12630;
  assign n20472 = n11289 & ~n13227;
  assign n20473 = n11908 & n12625;
  assign n20474 = ~n20472 & ~n20473;
  assign n20475 = ~n20471 & n20474;
  assign n20476 = ~n20470 & n20475;
  assign n20477 = pi2  & n20476;
  assign n20478 = ~pi2  & ~n20476;
  assign n20479 = ~n20477 & ~n20478;
  assign n20480 = n20469 & ~n20479;
  assign n20481 = n19877 & n20375;
  assign n20482 = ~n20376 & ~n20481;
  assign n20483 = n11288 & n12636;
  assign n20484 = n11894 & n12633;
  assign n20485 = n11289 & n13292;
  assign n20486 = n11908 & n12630;
  assign n20487 = ~n20485 & ~n20486;
  assign n20488 = ~n20484 & n20487;
  assign n20489 = ~n20483 & n20488;
  assign n20490 = pi2  & n20489;
  assign n20491 = ~pi2  & ~n20489;
  assign n20492 = ~n20490 & ~n20491;
  assign n20493 = n20482 & ~n20492;
  assign n20494 = n20371 & ~n20373;
  assign n20495 = ~n20374 & ~n20494;
  assign n20496 = n11288 & n12639;
  assign n20497 = n11894 & n12636;
  assign n20498 = n11289 & n13396;
  assign n20499 = n11908 & n12633;
  assign n20500 = ~n20498 & ~n20499;
  assign n20501 = ~n20497 & n20500;
  assign n20502 = ~n20496 & n20501;
  assign n20503 = pi2  & n20502;
  assign n20504 = ~pi2  & ~n20502;
  assign n20505 = ~n20503 & ~n20504;
  assign n20506 = n20495 & ~n20505;
  assign n20507 = n20367 & ~n20369;
  assign n20508 = ~n20370 & ~n20507;
  assign n20509 = n11288 & n12644;
  assign n20510 = n11894 & n12639;
  assign n20511 = n11289 & n13210;
  assign n20512 = n11908 & n12636;
  assign n20513 = ~n20511 & ~n20512;
  assign n20514 = ~n20510 & n20513;
  assign n20515 = ~n20509 & n20514;
  assign n20516 = pi2  & n20515;
  assign n20517 = ~pi2  & ~n20515;
  assign n20518 = ~n20516 & ~n20517;
  assign n20519 = n20508 & ~n20518;
  assign n20520 = n20508 & n20518;
  assign n20521 = ~n20508 & ~n20518;
  assign n20522 = ~n20520 & ~n20521;
  assign n20523 = n20363 & ~n20365;
  assign n20524 = ~n20366 & ~n20523;
  assign n20525 = n20358 & n20361;
  assign n20526 = ~n20362 & ~n20525;
  assign n20527 = n11288 & n12653;
  assign n20528 = n11894 & n12650;
  assign n20529 = n11289 & n13042;
  assign n20530 = n11908 & n12647;
  assign n20531 = ~n20529 & ~n20530;
  assign n20532 = ~n20528 & n20531;
  assign n20533 = ~n20527 & n20532;
  assign n20534 = pi2  & n20533;
  assign n20535 = ~pi2  & ~n20533;
  assign n20536 = ~n20534 & ~n20535;
  assign n20537 = n11288 & n12656;
  assign n20538 = n11894 & n12653;
  assign n20539 = n11289 & n12991;
  assign n20540 = n11908 & n12650;
  assign n20541 = ~n20539 & ~n20540;
  assign n20542 = ~n20538 & n20541;
  assign n20543 = ~n20537 & n20542;
  assign n20544 = pi2  & n20543;
  assign n20545 = ~pi2  & ~n20543;
  assign n20546 = ~n20544 & ~n20545;
  assign n20547 = n11288 & n12659;
  assign n20548 = n11894 & n12656;
  assign n20549 = n11289 & n13059;
  assign n20550 = n11908 & n12653;
  assign n20551 = ~n20549 & ~n20550;
  assign n20552 = ~n20548 & n20551;
  assign n20553 = ~n20547 & n20552;
  assign n20554 = pi2  & n20553;
  assign n20555 = ~pi2  & ~n20553;
  assign n20556 = ~n20554 & ~n20555;
  assign n20557 = n20346 & ~n20348;
  assign n20558 = ~n20349 & ~n20557;
  assign n20559 = n20341 & n20344;
  assign n20560 = ~n20345 & ~n20559;
  assign n20561 = n20336 & n20339;
  assign n20562 = ~n20340 & ~n20561;
  assign n20563 = n11288 & n12671;
  assign n20564 = n11894 & n12668;
  assign n20565 = n11289 & n13578;
  assign n20566 = n11908 & n12665;
  assign n20567 = ~n20565 & ~n20566;
  assign n20568 = ~n20564 & n20567;
  assign n20569 = ~n20563 & n20568;
  assign n20570 = pi2  & n20569;
  assign n20571 = ~pi2  & ~n20569;
  assign n20572 = ~n20570 & ~n20571;
  assign n20573 = n11288 & n12674;
  assign n20574 = n11894 & n12671;
  assign n20575 = n11289 & n13764;
  assign n20576 = n11908 & n12668;
  assign n20577 = ~n20575 & ~n20576;
  assign n20578 = ~n20574 & n20577;
  assign n20579 = ~n20573 & n20578;
  assign n20580 = pi2  & n20579;
  assign n20581 = ~pi2  & ~n20579;
  assign n20582 = ~n20580 & ~n20581;
  assign n20583 = n11288 & n12677;
  assign n20584 = n11894 & n12674;
  assign n20585 = n11289 & n13785;
  assign n20586 = n11908 & n12671;
  assign n20587 = ~n20585 & ~n20586;
  assign n20588 = ~n20584 & n20587;
  assign n20589 = ~n20583 & n20588;
  assign n20590 = pi2  & n20589;
  assign n20591 = ~pi2  & ~n20589;
  assign n20592 = ~n20590 & ~n20591;
  assign n20593 = n20324 & ~n20326;
  assign n20594 = ~n20327 & ~n20593;
  assign n20595 = n20319 & n20322;
  assign n20596 = ~n20323 & ~n20595;
  assign n20597 = n20314 & n20317;
  assign n20598 = ~n20318 & ~n20597;
  assign n20599 = n11288 & n12689;
  assign n20600 = n11894 & n12686;
  assign n20601 = n11289 & n14552;
  assign n20602 = n11908 & n12683;
  assign n20603 = ~n20601 & ~n20602;
  assign n20604 = ~n20600 & n20603;
  assign n20605 = ~n20599 & n20604;
  assign n20606 = pi2  & n20605;
  assign n20607 = ~pi2  & ~n20605;
  assign n20608 = ~n20606 & ~n20607;
  assign n20609 = n11288 & n12692;
  assign n20610 = n11894 & n12689;
  assign n20611 = n11289 & n14382;
  assign n20612 = n11908 & n12686;
  assign n20613 = ~n20611 & ~n20612;
  assign n20614 = ~n20610 & n20613;
  assign n20615 = ~n20609 & n20614;
  assign n20616 = pi2  & n20615;
  assign n20617 = ~pi2  & ~n20615;
  assign n20618 = ~n20616 & ~n20617;
  assign n20619 = n11288 & n12695;
  assign n20620 = n11894 & n12692;
  assign n20621 = n11289 & n14677;
  assign n20622 = n11908 & n12689;
  assign n20623 = ~n20621 & ~n20622;
  assign n20624 = ~n20620 & n20623;
  assign n20625 = ~n20619 & n20624;
  assign n20626 = pi2  & n20625;
  assign n20627 = ~pi2  & ~n20625;
  assign n20628 = ~n20626 & ~n20627;
  assign n20629 = n20302 & ~n20304;
  assign n20630 = ~n20305 & ~n20629;
  assign n20631 = n20297 & n20300;
  assign n20632 = ~n20301 & ~n20631;
  assign n20633 = n20292 & n20295;
  assign n20634 = ~n20296 & ~n20633;
  assign n20635 = n11288 & n12707;
  assign n20636 = n11894 & n12704;
  assign n20637 = n11289 & n15024;
  assign n20638 = n11908 & n12701;
  assign n20639 = ~n20637 & ~n20638;
  assign n20640 = ~n20636 & n20639;
  assign n20641 = ~n20635 & n20640;
  assign n20642 = pi2  & n20641;
  assign n20643 = ~pi2  & ~n20641;
  assign n20644 = ~n20642 & ~n20643;
  assign n20645 = n11288 & n12710;
  assign n20646 = n11894 & n12707;
  assign n20647 = n11289 & n15050;
  assign n20648 = n11908 & n12704;
  assign n20649 = ~n20647 & ~n20648;
  assign n20650 = ~n20646 & n20649;
  assign n20651 = ~n20645 & n20650;
  assign n20652 = pi2  & n20651;
  assign n20653 = ~pi2  & ~n20651;
  assign n20654 = ~n20652 & ~n20653;
  assign n20655 = n11288 & n12713;
  assign n20656 = n11894 & n12710;
  assign n20657 = n11289 & n15074;
  assign n20658 = n11908 & n12707;
  assign n20659 = ~n20657 & ~n20658;
  assign n20660 = ~n20656 & n20659;
  assign n20661 = ~n20655 & n20660;
  assign n20662 = pi2  & n20661;
  assign n20663 = ~pi2  & ~n20661;
  assign n20664 = ~n20662 & ~n20663;
  assign n20665 = n20280 & ~n20282;
  assign n20666 = ~n20283 & ~n20665;
  assign n20667 = n11288 & n12719;
  assign n20668 = n11894 & n12716;
  assign n20669 = n11289 & n15161;
  assign n20670 = n11908 & n12713;
  assign n20671 = ~n20669 & ~n20670;
  assign n20672 = ~n20668 & n20671;
  assign n20673 = ~n20667 & n20672;
  assign n20674 = pi2  & n20673;
  assign n20675 = ~pi2  & ~n20673;
  assign n20676 = ~n20674 & ~n20675;
  assign n20677 = pi5  & ~n20256;
  assign n20678 = n20263 & ~n20677;
  assign n20679 = ~n20263 & n20677;
  assign n20680 = ~n20678 & ~n20679;
  assign n20681 = n11288 & n12725;
  assign n20682 = n11894 & n12722;
  assign n20683 = n11289 & n15243;
  assign n20684 = n11908 & n12719;
  assign n20685 = ~n20683 & ~n20684;
  assign n20686 = ~n20682 & n20685;
  assign n20687 = ~n20681 & n20686;
  assign n20688 = pi2  & n20687;
  assign n20689 = ~pi2  & ~n20687;
  assign n20690 = ~n20688 & ~n20689;
  assign n20691 = ~n11287 & n12732;
  assign n20692 = n11908 & n12730;
  assign n20693 = n12139 & ~n15356;
  assign n20694 = n11288 & n12732;
  assign n20695 = n11894 & n12730;
  assign n20696 = n11908 & n12725;
  assign n20697 = ~n20695 & ~n20696;
  assign n20698 = ~n20694 & n20697;
  assign n20699 = pi2  & ~n20698;
  assign n20700 = n12139 & ~n15312;
  assign n20701 = pi2  & ~n20700;
  assign n20702 = ~n20699 & n20701;
  assign n20703 = ~n20693 & n20702;
  assign n20704 = ~n20692 & n20703;
  assign n20705 = ~n20691 & n20704;
  assign n20706 = n20254 & n20705;
  assign n20707 = ~n20254 & ~n20705;
  assign n20708 = n11288 & n12730;
  assign n20709 = n11894 & n12725;
  assign n20710 = n11289 & n15267;
  assign n20711 = n11908 & n12722;
  assign n20712 = ~n20710 & ~n20711;
  assign n20713 = ~n20709 & n20712;
  assign n20714 = ~n20708 & n20713;
  assign n20715 = pi2  & ~n20714;
  assign n20716 = ~pi2  & n20714;
  assign n20717 = ~n20715 & ~n20716;
  assign n20718 = ~n20707 & n20717;
  assign n20719 = ~n20706 & ~n20718;
  assign n20720 = ~n20690 & ~n20719;
  assign n20721 = n20690 & n20719;
  assign n20722 = pi5  & n20254;
  assign n20723 = ~n20253 & n20722;
  assign n20724 = n20253 & ~n20722;
  assign n20725 = ~n20723 & ~n20724;
  assign n20726 = ~n20721 & n20725;
  assign n20727 = ~n20720 & ~n20726;
  assign n20728 = n20680 & ~n20727;
  assign n20729 = ~n20680 & n20727;
  assign n20730 = n11288 & n12722;
  assign n20731 = n11894 & n12719;
  assign n20732 = n11289 & n15199;
  assign n20733 = n11908 & n12716;
  assign n20734 = ~n20732 & ~n20733;
  assign n20735 = ~n20731 & n20734;
  assign n20736 = ~n20730 & n20735;
  assign n20737 = pi2  & ~n20736;
  assign n20738 = ~pi2  & n20736;
  assign n20739 = ~n20737 & ~n20738;
  assign n20740 = ~n20729 & n20739;
  assign n20741 = ~n20728 & ~n20740;
  assign n20742 = ~n20676 & ~n20741;
  assign n20743 = n20676 & n20741;
  assign n20744 = n20268 & n20278;
  assign n20745 = ~n20279 & ~n20744;
  assign n20746 = ~n20743 & n20745;
  assign n20747 = ~n20742 & ~n20746;
  assign n20748 = n20666 & ~n20747;
  assign n20749 = ~n20666 & n20747;
  assign n20750 = n11288 & n12716;
  assign n20751 = n11894 & n12713;
  assign n20752 = n11289 & n15105;
  assign n20753 = n11908 & n12710;
  assign n20754 = ~n20752 & ~n20753;
  assign n20755 = ~n20751 & n20754;
  assign n20756 = ~n20750 & n20755;
  assign n20757 = pi2  & ~n20756;
  assign n20758 = ~pi2  & n20756;
  assign n20759 = ~n20757 & ~n20758;
  assign n20760 = ~n20749 & n20759;
  assign n20761 = ~n20748 & ~n20760;
  assign n20762 = ~n20664 & ~n20761;
  assign n20763 = n20664 & n20761;
  assign n20764 = n20233 & n20284;
  assign n20765 = ~n20285 & ~n20764;
  assign n20766 = ~n20763 & n20765;
  assign n20767 = ~n20762 & ~n20766;
  assign n20768 = ~n20654 & ~n20767;
  assign n20769 = n20654 & n20767;
  assign n20770 = n20286 & ~n20288;
  assign n20771 = ~n20289 & ~n20770;
  assign n20772 = ~n20769 & n20771;
  assign n20773 = ~n20768 & ~n20772;
  assign n20774 = ~n20644 & ~n20773;
  assign n20775 = n20644 & n20773;
  assign n20776 = n20202 & n20290;
  assign n20777 = ~n20291 & ~n20776;
  assign n20778 = ~n20775 & n20777;
  assign n20779 = ~n20774 & ~n20778;
  assign n20780 = n20634 & ~n20779;
  assign n20781 = ~n20634 & n20779;
  assign n20782 = n11288 & n12704;
  assign n20783 = n11894 & n12701;
  assign n20784 = n11289 & n14655;
  assign n20785 = n11908 & n12698;
  assign n20786 = ~n20784 & ~n20785;
  assign n20787 = ~n20783 & n20786;
  assign n20788 = ~n20782 & n20787;
  assign n20789 = pi2  & ~n20788;
  assign n20790 = ~pi2  & n20788;
  assign n20791 = ~n20789 & ~n20790;
  assign n20792 = ~n20781 & n20791;
  assign n20793 = ~n20780 & ~n20792;
  assign n20794 = n20632 & ~n20793;
  assign n20795 = ~n20632 & n20793;
  assign n20796 = n11288 & n12701;
  assign n20797 = n11894 & n12698;
  assign n20798 = n11289 & n14991;
  assign n20799 = n11908 & n12695;
  assign n20800 = ~n20798 & ~n20799;
  assign n20801 = ~n20797 & n20800;
  assign n20802 = ~n20796 & n20801;
  assign n20803 = pi2  & ~n20802;
  assign n20804 = ~pi2  & n20802;
  assign n20805 = ~n20803 & ~n20804;
  assign n20806 = ~n20795 & n20805;
  assign n20807 = ~n20794 & ~n20806;
  assign n20808 = n20630 & ~n20807;
  assign n20809 = ~n20630 & n20807;
  assign n20810 = n11288 & n12698;
  assign n20811 = n11894 & n12695;
  assign n20812 = n11289 & n14976;
  assign n20813 = n11908 & n12692;
  assign n20814 = ~n20812 & ~n20813;
  assign n20815 = ~n20811 & n20814;
  assign n20816 = ~n20810 & n20815;
  assign n20817 = pi2  & ~n20816;
  assign n20818 = ~pi2  & n20816;
  assign n20819 = ~n20817 & ~n20818;
  assign n20820 = ~n20809 & n20819;
  assign n20821 = ~n20808 & ~n20820;
  assign n20822 = ~n20628 & ~n20821;
  assign n20823 = n20628 & n20821;
  assign n20824 = n20306 & ~n20308;
  assign n20825 = ~n20309 & ~n20824;
  assign n20826 = ~n20823 & n20825;
  assign n20827 = ~n20822 & ~n20826;
  assign n20828 = ~n20618 & ~n20827;
  assign n20829 = n20618 & n20827;
  assign n20830 = n20133 & n20310;
  assign n20831 = ~n20311 & ~n20830;
  assign n20832 = ~n20829 & n20831;
  assign n20833 = ~n20828 & ~n20832;
  assign n20834 = ~n20608 & ~n20833;
  assign n20835 = n20608 & n20833;
  assign n20836 = n20117 & n20312;
  assign n20837 = ~n20313 & ~n20836;
  assign n20838 = ~n20835 & n20837;
  assign n20839 = ~n20834 & ~n20838;
  assign n20840 = n20598 & ~n20839;
  assign n20841 = ~n20598 & n20839;
  assign n20842 = n11288 & n12686;
  assign n20843 = n11894 & n12683;
  assign n20844 = n11289 & n14402;
  assign n20845 = n11908 & n12680;
  assign n20846 = ~n20844 & ~n20845;
  assign n20847 = ~n20843 & n20846;
  assign n20848 = ~n20842 & n20847;
  assign n20849 = pi2  & ~n20848;
  assign n20850 = ~pi2  & n20848;
  assign n20851 = ~n20849 & ~n20850;
  assign n20852 = ~n20841 & n20851;
  assign n20853 = ~n20840 & ~n20852;
  assign n20854 = n20596 & ~n20853;
  assign n20855 = ~n20596 & n20853;
  assign n20856 = n11288 & n12683;
  assign n20857 = n11894 & n12680;
  assign n20858 = n11289 & n13929;
  assign n20859 = n11908 & n12677;
  assign n20860 = ~n20858 & ~n20859;
  assign n20861 = ~n20857 & n20860;
  assign n20862 = ~n20856 & n20861;
  assign n20863 = pi2  & ~n20862;
  assign n20864 = ~pi2  & n20862;
  assign n20865 = ~n20863 & ~n20864;
  assign n20866 = ~n20855 & n20865;
  assign n20867 = ~n20854 & ~n20866;
  assign n20868 = n20594 & ~n20867;
  assign n20869 = ~n20594 & n20867;
  assign n20870 = n11288 & n12680;
  assign n20871 = n11894 & n12677;
  assign n20872 = n11289 & n14164;
  assign n20873 = n11908 & n12674;
  assign n20874 = ~n20872 & ~n20873;
  assign n20875 = ~n20871 & n20874;
  assign n20876 = ~n20870 & n20875;
  assign n20877 = pi2  & ~n20876;
  assign n20878 = ~pi2  & n20876;
  assign n20879 = ~n20877 & ~n20878;
  assign n20880 = ~n20869 & n20879;
  assign n20881 = ~n20868 & ~n20880;
  assign n20882 = ~n20592 & ~n20881;
  assign n20883 = n20592 & n20881;
  assign n20884 = n20062 & n20328;
  assign n20885 = ~n20329 & ~n20884;
  assign n20886 = ~n20883 & n20885;
  assign n20887 = ~n20882 & ~n20886;
  assign n20888 = ~n20582 & ~n20887;
  assign n20889 = n20582 & n20887;
  assign n20890 = n20330 & ~n20332;
  assign n20891 = ~n20333 & ~n20890;
  assign n20892 = ~n20889 & n20891;
  assign n20893 = ~n20888 & ~n20892;
  assign n20894 = ~n20572 & ~n20893;
  assign n20895 = n20572 & n20893;
  assign n20896 = n20032 & n20334;
  assign n20897 = ~n20335 & ~n20896;
  assign n20898 = ~n20895 & n20897;
  assign n20899 = ~n20894 & ~n20898;
  assign n20900 = n20562 & ~n20899;
  assign n20901 = ~n20562 & n20899;
  assign n20902 = n11288 & n12668;
  assign n20903 = n11894 & n12665;
  assign n20904 = n11289 & n13591;
  assign n20905 = n11908 & n12662;
  assign n20906 = ~n20904 & ~n20905;
  assign n20907 = ~n20903 & n20906;
  assign n20908 = ~n20902 & n20907;
  assign n20909 = pi2  & ~n20908;
  assign n20910 = ~pi2  & n20908;
  assign n20911 = ~n20909 & ~n20910;
  assign n20912 = ~n20901 & n20911;
  assign n20913 = ~n20900 & ~n20912;
  assign n20914 = n20560 & ~n20913;
  assign n20915 = ~n20560 & n20913;
  assign n20916 = n11288 & n12665;
  assign n20917 = n11894 & n12662;
  assign n20918 = n11289 & n13165;
  assign n20919 = n11908 & n12659;
  assign n20920 = ~n20918 & ~n20919;
  assign n20921 = ~n20917 & n20920;
  assign n20922 = ~n20916 & n20921;
  assign n20923 = pi2  & ~n20922;
  assign n20924 = ~pi2  & n20922;
  assign n20925 = ~n20923 & ~n20924;
  assign n20926 = ~n20915 & n20925;
  assign n20927 = ~n20914 & ~n20926;
  assign n20928 = n20558 & ~n20927;
  assign n20929 = ~n20558 & n20927;
  assign n20930 = n11288 & n12662;
  assign n20931 = n11894 & n12659;
  assign n20932 = n11289 & n13246;
  assign n20933 = n11908 & n12656;
  assign n20934 = ~n20932 & ~n20933;
  assign n20935 = ~n20931 & n20934;
  assign n20936 = ~n20930 & n20935;
  assign n20937 = pi2  & ~n20936;
  assign n20938 = ~pi2  & n20936;
  assign n20939 = ~n20937 & ~n20938;
  assign n20940 = ~n20929 & n20939;
  assign n20941 = ~n20928 & ~n20940;
  assign n20942 = ~n20556 & ~n20941;
  assign n20943 = n20556 & n20941;
  assign n20944 = n20350 & ~n20352;
  assign n20945 = ~n20353 & ~n20944;
  assign n20946 = ~n20943 & n20945;
  assign n20947 = ~n20942 & ~n20946;
  assign n20948 = ~n20546 & ~n20947;
  assign n20949 = n20546 & n20947;
  assign n20950 = n19963 & n20354;
  assign n20951 = ~n20355 & ~n20950;
  assign n20952 = ~n20949 & n20951;
  assign n20953 = ~n20948 & ~n20952;
  assign n20954 = ~n20536 & ~n20953;
  assign n20955 = n20536 & n20953;
  assign n20956 = n19947 & n20356;
  assign n20957 = ~n20357 & ~n20956;
  assign n20958 = ~n20955 & n20957;
  assign n20959 = ~n20954 & ~n20958;
  assign n20960 = n20526 & ~n20959;
  assign n20961 = ~n20526 & n20959;
  assign n20962 = n11288 & n12650;
  assign n20963 = n11894 & n12647;
  assign n20964 = n11289 & n13275;
  assign n20965 = n11908 & n12644;
  assign n20966 = ~n20964 & ~n20965;
  assign n20967 = ~n20963 & n20966;
  assign n20968 = ~n20962 & n20967;
  assign n20969 = pi2  & ~n20968;
  assign n20970 = ~pi2  & n20968;
  assign n20971 = ~n20969 & ~n20970;
  assign n20972 = ~n20961 & n20971;
  assign n20973 = ~n20960 & ~n20972;
  assign n20974 = n20524 & ~n20973;
  assign n20975 = ~n20524 & n20973;
  assign n20976 = n11288 & n12647;
  assign n20977 = n11894 & n12644;
  assign n20978 = n11289 & ~n13193;
  assign n20979 = n11908 & n12639;
  assign n20980 = ~n20978 & ~n20979;
  assign n20981 = ~n20977 & n20980;
  assign n20982 = ~n20976 & n20981;
  assign n20983 = pi2  & ~n20982;
  assign n20984 = ~pi2  & n20982;
  assign n20985 = ~n20983 & ~n20984;
  assign n20986 = ~n20975 & n20985;
  assign n20987 = ~n20974 & ~n20986;
  assign n20988 = ~n20522 & ~n20987;
  assign n20989 = ~n20519 & ~n20988;
  assign n20990 = ~n20495 & n20505;
  assign n20991 = ~n20506 & ~n20990;
  assign n20992 = ~n20989 & n20991;
  assign n20993 = ~n20506 & ~n20992;
  assign n20994 = ~n20482 & n20492;
  assign n20995 = ~n20493 & ~n20994;
  assign n20996 = ~n20993 & n20995;
  assign n20997 = ~n20493 & ~n20996;
  assign n20998 = ~n20469 & n20479;
  assign n20999 = ~n20480 & ~n20998;
  assign n21000 = ~n20997 & n20999;
  assign n21001 = ~n20480 & ~n21000;
  assign n21002 = ~n20456 & n20466;
  assign n21003 = ~n20467 & ~n21002;
  assign n21004 = ~n21001 & n21003;
  assign n21005 = ~n20467 & ~n21004;
  assign n21006 = ~n20443 & n20453;
  assign n21007 = ~n20454 & ~n21006;
  assign n21008 = ~n21005 & n21007;
  assign n21009 = ~n20454 & ~n21008;
  assign n21010 = ~n20430 & n20440;
  assign n21011 = ~n20441 & ~n21010;
  assign n21012 = ~n21009 & n21011;
  assign n21013 = ~n20441 & ~n21012;
  assign n21014 = ~n20417 & n20427;
  assign n21015 = ~n20428 & ~n21014;
  assign n21016 = ~n21013 & n21015;
  assign n21017 = ~n20428 & ~n21016;
  assign n21018 = ~n20404 & n20414;
  assign n21019 = ~n20415 & ~n21018;
  assign n21020 = ~n21017 & n21019;
  assign n21021 = ~n20415 & ~n21020;
  assign n21022 = n20402 & ~n21021;
  assign n21023 = ~n20400 & ~n21022;
  assign n21024 = n19773 & ~n21023;
  assign n21025 = ~n19771 & ~n21024;
  assign n21026 = n19739 & ~n21025;
  assign n21027 = ~n19737 & ~n21026;
  assign n21028 = n19126 & ~n21027;
  assign n21029 = ~n19124 & ~n21028;
  assign n21030 = ~n18013 & n18547;
  assign n21031 = ~n18548 & ~n21030;
  assign n21032 = ~n21029 & n21031;
  assign n21033 = ~n18548 & ~n21032;
  assign n21034 = ~n18011 & ~n21033;
  assign n21035 = ~n18008 & ~n21034;
  assign n21036 = n17503 & ~n21035;
  assign n21037 = ~n17501 & ~n21036;
  assign n21038 = ~n16603 & n17031;
  assign n21039 = ~n17032 & ~n21038;
  assign n21040 = ~n21037 & n21039;
  assign n21041 = ~n17032 & ~n21040;
  assign n21042 = ~n16601 & ~n21041;
  assign n21043 = ~n16598 & ~n21042;
  assign n21044 = n16199 & ~n21043;
  assign n21045 = ~n16197 & ~n21044;
  assign n21046 = ~n15689 & n15841;
  assign n21047 = ~n15842 & ~n21046;
  assign n21048 = ~n21045 & n21047;
  assign n21049 = ~n15842 & ~n21048;
  assign n21050 = ~n15687 & ~n21049;
  assign n21051 = ~n15684 & ~n21050;
  assign n21052 = n15524 & ~n21051;
  assign n21053 = ~n15522 & ~n21052;
  assign n21054 = ~n14789 & n14924;
  assign n21055 = ~n14925 & ~n21054;
  assign n21056 = ~n21053 & n21055;
  assign n21057 = ~n14925 & ~n21056;
  assign n21058 = ~n14787 & ~n21057;
  assign n21059 = ~n14784 & ~n21058;
  assign n21060 = n14497 & ~n21059;
  assign n21061 = ~n14495 & ~n21060;
  assign n21062 = ~n14129 & n14258;
  assign n21063 = ~n14259 & ~n21062;
  assign n21064 = ~n21061 & n21063;
  assign n21065 = ~n14259 & ~n21064;
  assign n21066 = ~n14127 & ~n21065;
  assign n21067 = ~n14124 & ~n21066;
  assign n21068 = n14019 & ~n21067;
  assign n21069 = ~n14017 & ~n21068;
  assign n21070 = ~n13498 & n13657;
  assign n21071 = ~n13658 & ~n21070;
  assign n21072 = ~n21069 & n21071;
  assign n21073 = ~n13658 & ~n21072;
  assign n21074 = ~n13496 & ~n21073;
  assign n21075 = n13496 & n21073;
  assign n21076 = ~n21074 & ~n21075;
  assign n21077 = n9725 & n21076;
  assign n21078 = n5239 & ~n13499;
  assign n21079 = n5238 & ~n12611;
  assign n21080 = ~n71 & ~n5326;
  assign n21081 = ~n21079 & n21080;
  assign n21082 = ~n12608 & ~n21081;
  assign n21083 = ~n21078 & ~n21082;
  assign n21084 = pi23  & n21083;
  assign n21085 = ~pi23  & ~n21083;
  assign n21086 = ~n21084 & ~n21085;
  assign n21087 = ~n13458 & ~n13471;
  assign n21088 = ~n13457 & ~n21087;
  assign n21089 = ~n21086 & ~n21088;
  assign n21090 = n21086 & n21088;
  assign n21091 = ~n21089 & ~n21090;
  assign n21092 = ~n13439 & ~n13452;
  assign n21093 = n4006 & n12633;
  assign n21094 = n4133 & n12630;
  assign n21095 = n4002 & ~n13227;
  assign n21096 = n4555 & n12625;
  assign n21097 = ~n21095 & ~n21096;
  assign n21098 = ~n21094 & n21097;
  assign n21099 = ~n21093 & n21098;
  assign n21100 = pi29  & n21099;
  assign n21101 = ~pi29  & ~n21099;
  assign n21102 = ~n21100 & ~n21101;
  assign n21103 = ~n13424 & ~n13434;
  assign n21104 = n977 & n5163;
  assign n21105 = ~n548 & n21104;
  assign n21106 = n6361 & n12904;
  assign n21107 = n765 & n21106;
  assign n21108 = ~n326 & n21107;
  assign n21109 = n21105 & n21108;
  assign n21110 = n1401 & n4084;
  assign n21111 = ~n203 & n21110;
  assign n21112 = n1859 & n3045;
  assign n21113 = ~n477 & n21112;
  assign n21114 = ~n636 & n21113;
  assign n21115 = n21111 & n21114;
  assign n21116 = ~n455 & n21115;
  assign n21117 = ~n294 & n1024;
  assign n21118 = ~n385 & n21117;
  assign n21119 = n878 & n21118;
  assign n21120 = n21116 & n21119;
  assign n21121 = n1025 & n21120;
  assign n21122 = n1784 & n21121;
  assign n21123 = ~n134 & n21122;
  assign n21124 = n1181 & n4274;
  assign n21125 = ~n180 & n21124;
  assign n21126 = ~n612 & n21125;
  assign n21127 = n21123 & n21126;
  assign n21128 = n21109 & n21127;
  assign n21129 = ~n12593 & n21128;
  assign n21130 = n12593 & ~n21128;
  assign n21131 = ~n21129 & ~n21130;
  assign n21132 = n21103 & n21131;
  assign n21133 = ~n21103 & ~n21131;
  assign n21134 = ~n21132 & ~n21133;
  assign n21135 = n3641 & n12644;
  assign n21136 = n3740 & n12639;
  assign n21137 = n556 & n13210;
  assign n21138 = n3961 & n12636;
  assign n21139 = ~n21137 & ~n21138;
  assign n21140 = ~n21136 & n21139;
  assign n21141 = ~n21135 & n21140;
  assign n21142 = ~n21134 & ~n21141;
  assign n21143 = n21134 & n21141;
  assign n21144 = ~n21142 & ~n21143;
  assign n21145 = ~n21102 & n21144;
  assign n21146 = n21102 & ~n21144;
  assign n21147 = ~n21145 & ~n21146;
  assign n21148 = ~n21092 & n21147;
  assign n21149 = n21092 & ~n21147;
  assign n21150 = ~n21148 & ~n21149;
  assign n21151 = n4601 & n12622;
  assign n21152 = n4783 & n12614;
  assign n21153 = n4602 & ~n13310;
  assign n21154 = n4801 & n12606;
  assign n21155 = ~n21153 & ~n21154;
  assign n21156 = ~n21152 & n21155;
  assign n21157 = ~n21151 & n21156;
  assign n21158 = pi26  & n21157;
  assign n21159 = ~pi26  & ~n21157;
  assign n21160 = ~n21158 & ~n21159;
  assign n21161 = n21150 & ~n21160;
  assign n21162 = ~n21150 & n21160;
  assign n21163 = ~n21161 & ~n21162;
  assign n21164 = n21091 & n21163;
  assign n21165 = ~n21091 & ~n21163;
  assign n21166 = ~n21164 & ~n21165;
  assign n21167 = ~n13476 & ~n13490;
  assign n21168 = ~n13475 & ~n21167;
  assign n21169 = n21166 & ~n21168;
  assign n21170 = ~n21166 & n21168;
  assign n21171 = ~n21169 & ~n21170;
  assign n21172 = ~n13420 & n13493;
  assign n21173 = ~n21074 & ~n21172;
  assign n21174 = n21171 & ~n21173;
  assign n21175 = ~n21171 & n21173;
  assign n21176 = ~n21174 & ~n21175;
  assign n21177 = n10702 & n21176;
  assign n21178 = n21076 & n21176;
  assign n21179 = n21069 & ~n21071;
  assign n21180 = ~n21072 & ~n21179;
  assign n21181 = n21076 & n21180;
  assign n21182 = ~n14019 & n21067;
  assign n21183 = ~n21068 & ~n21182;
  assign n21184 = n21180 & n21183;
  assign n21185 = n14127 & n21065;
  assign n21186 = ~n21066 & ~n21185;
  assign n21187 = n21183 & n21186;
  assign n21188 = n21061 & ~n21063;
  assign n21189 = ~n21064 & ~n21188;
  assign n21190 = n21186 & n21189;
  assign n21191 = ~n14497 & n21059;
  assign n21192 = ~n21060 & ~n21191;
  assign n21193 = n21189 & n21192;
  assign n21194 = n14787 & n21057;
  assign n21195 = ~n21058 & ~n21194;
  assign n21196 = n21192 & n21195;
  assign n21197 = n21053 & ~n21055;
  assign n21198 = ~n21056 & ~n21197;
  assign n21199 = n21195 & n21198;
  assign n21200 = ~n15524 & n21051;
  assign n21201 = ~n21052 & ~n21200;
  assign n21202 = n21198 & n21201;
  assign n21203 = n15687 & n21049;
  assign n21204 = ~n21050 & ~n21203;
  assign n21205 = n21201 & n21204;
  assign n21206 = n21045 & ~n21047;
  assign n21207 = ~n21048 & ~n21206;
  assign n21208 = n21204 & n21207;
  assign n21209 = ~n16199 & n21043;
  assign n21210 = ~n21044 & ~n21209;
  assign n21211 = n21207 & n21210;
  assign n21212 = n16601 & n21041;
  assign n21213 = ~n21042 & ~n21212;
  assign n21214 = n21210 & n21213;
  assign n21215 = n21037 & ~n21039;
  assign n21216 = ~n21040 & ~n21215;
  assign n21217 = n21213 & n21216;
  assign n21218 = ~n17503 & n21035;
  assign n21219 = ~n21036 & ~n21218;
  assign n21220 = n21216 & n21219;
  assign n21221 = n18011 & n21033;
  assign n21222 = ~n21034 & ~n21221;
  assign n21223 = n21219 & n21222;
  assign n21224 = n21029 & ~n21031;
  assign n21225 = ~n21032 & ~n21224;
  assign n21226 = n21222 & n21225;
  assign n21227 = ~n19126 & n21027;
  assign n21228 = ~n21028 & ~n21227;
  assign n21229 = n21225 & n21228;
  assign n21230 = ~n19739 & n21025;
  assign n21231 = ~n21026 & ~n21230;
  assign n21232 = n21228 & n21231;
  assign n21233 = ~n19773 & n21023;
  assign n21234 = ~n21024 & ~n21233;
  assign n21235 = n21231 & n21234;
  assign n21236 = ~n20402 & n21021;
  assign n21237 = ~n21022 & ~n21236;
  assign n21238 = n21234 & n21237;
  assign n21239 = n21017 & ~n21019;
  assign n21240 = ~n21020 & ~n21239;
  assign n21241 = n21237 & n21240;
  assign n21242 = n21013 & ~n21015;
  assign n21243 = ~n21016 & ~n21242;
  assign n21244 = n21240 & n21243;
  assign n21245 = n21009 & ~n21011;
  assign n21246 = ~n21012 & ~n21245;
  assign n21247 = n21243 & n21246;
  assign n21248 = n21005 & ~n21007;
  assign n21249 = ~n21008 & ~n21248;
  assign n21250 = n21246 & n21249;
  assign n21251 = n21001 & ~n21003;
  assign n21252 = ~n21004 & ~n21251;
  assign n21253 = n21249 & n21252;
  assign n21254 = n20997 & ~n20999;
  assign n21255 = ~n21000 & ~n21254;
  assign n21256 = n21252 & n21255;
  assign n21257 = n20993 & ~n20995;
  assign n21258 = ~n20996 & ~n21257;
  assign n21259 = n21255 & n21258;
  assign n21260 = ~n21255 & ~n21258;
  assign n21261 = ~n21259 & ~n21260;
  assign n21262 = n20989 & ~n20991;
  assign n21263 = ~n20992 & ~n21262;
  assign n21264 = n20522 & n20987;
  assign n21265 = ~n20988 & ~n21264;
  assign n21266 = ~n21258 & ~n21265;
  assign n21267 = n21263 & ~n21266;
  assign n21268 = n21261 & n21267;
  assign n21269 = ~n21259 & ~n21268;
  assign n21270 = ~n21252 & ~n21255;
  assign n21271 = ~n21256 & ~n21270;
  assign n21272 = ~n21269 & n21271;
  assign n21273 = ~n21256 & ~n21272;
  assign n21274 = ~n21249 & ~n21252;
  assign n21275 = ~n21253 & ~n21274;
  assign n21276 = ~n21273 & n21275;
  assign n21277 = ~n21253 & ~n21276;
  assign n21278 = ~n21246 & ~n21249;
  assign n21279 = ~n21250 & ~n21278;
  assign n21280 = ~n21277 & n21279;
  assign n21281 = ~n21250 & ~n21280;
  assign n21282 = ~n21243 & ~n21246;
  assign n21283 = ~n21247 & ~n21282;
  assign n21284 = ~n21281 & n21283;
  assign n21285 = ~n21247 & ~n21284;
  assign n21286 = ~n21240 & ~n21243;
  assign n21287 = ~n21244 & ~n21286;
  assign n21288 = ~n21285 & n21287;
  assign n21289 = ~n21244 & ~n21288;
  assign n21290 = ~n21237 & ~n21240;
  assign n21291 = ~n21241 & ~n21290;
  assign n21292 = ~n21289 & n21291;
  assign n21293 = ~n21241 & ~n21292;
  assign n21294 = ~n21234 & ~n21237;
  assign n21295 = ~n21238 & ~n21294;
  assign n21296 = ~n21293 & n21295;
  assign n21297 = ~n21238 & ~n21296;
  assign n21298 = ~n21231 & ~n21234;
  assign n21299 = ~n21235 & ~n21298;
  assign n21300 = ~n21297 & n21299;
  assign n21301 = ~n21235 & ~n21300;
  assign n21302 = ~n21228 & ~n21231;
  assign n21303 = ~n21232 & ~n21302;
  assign n21304 = ~n21301 & n21303;
  assign n21305 = ~n21232 & ~n21304;
  assign n21306 = ~n21225 & ~n21228;
  assign n21307 = ~n21229 & ~n21306;
  assign n21308 = ~n21305 & n21307;
  assign n21309 = ~n21229 & ~n21308;
  assign n21310 = ~n21222 & ~n21225;
  assign n21311 = ~n21226 & ~n21310;
  assign n21312 = ~n21309 & n21311;
  assign n21313 = ~n21226 & ~n21312;
  assign n21314 = ~n21219 & ~n21222;
  assign n21315 = ~n21223 & ~n21314;
  assign n21316 = ~n21313 & n21315;
  assign n21317 = ~n21223 & ~n21316;
  assign n21318 = ~n21216 & ~n21219;
  assign n21319 = ~n21220 & ~n21318;
  assign n21320 = ~n21317 & n21319;
  assign n21321 = ~n21220 & ~n21320;
  assign n21322 = ~n21213 & ~n21216;
  assign n21323 = ~n21217 & ~n21322;
  assign n21324 = ~n21321 & n21323;
  assign n21325 = ~n21217 & ~n21324;
  assign n21326 = ~n21210 & ~n21213;
  assign n21327 = ~n21214 & ~n21326;
  assign n21328 = ~n21325 & n21327;
  assign n21329 = ~n21214 & ~n21328;
  assign n21330 = ~n21207 & ~n21210;
  assign n21331 = ~n21211 & ~n21330;
  assign n21332 = ~n21329 & n21331;
  assign n21333 = ~n21211 & ~n21332;
  assign n21334 = ~n21204 & ~n21207;
  assign n21335 = ~n21208 & ~n21334;
  assign n21336 = ~n21333 & n21335;
  assign n21337 = ~n21208 & ~n21336;
  assign n21338 = ~n21201 & ~n21204;
  assign n21339 = ~n21205 & ~n21338;
  assign n21340 = ~n21337 & n21339;
  assign n21341 = ~n21205 & ~n21340;
  assign n21342 = ~n21198 & ~n21201;
  assign n21343 = ~n21202 & ~n21342;
  assign n21344 = ~n21341 & n21343;
  assign n21345 = ~n21202 & ~n21344;
  assign n21346 = ~n21195 & ~n21198;
  assign n21347 = ~n21199 & ~n21346;
  assign n21348 = ~n21345 & n21347;
  assign n21349 = ~n21199 & ~n21348;
  assign n21350 = ~n21192 & ~n21195;
  assign n21351 = ~n21196 & ~n21350;
  assign n21352 = ~n21349 & n21351;
  assign n21353 = ~n21196 & ~n21352;
  assign n21354 = ~n21189 & ~n21192;
  assign n21355 = ~n21193 & ~n21354;
  assign n21356 = ~n21353 & n21355;
  assign n21357 = ~n21193 & ~n21356;
  assign n21358 = ~n21186 & ~n21189;
  assign n21359 = ~n21190 & ~n21358;
  assign n21360 = ~n21357 & n21359;
  assign n21361 = ~n21190 & ~n21360;
  assign n21362 = ~n21183 & ~n21186;
  assign n21363 = ~n21187 & ~n21362;
  assign n21364 = ~n21361 & n21363;
  assign n21365 = ~n21187 & ~n21364;
  assign n21366 = ~n21180 & ~n21183;
  assign n21367 = ~n21184 & ~n21366;
  assign n21368 = ~n21365 & n21367;
  assign n21369 = ~n21184 & ~n21368;
  assign n21370 = ~n21076 & ~n21180;
  assign n21371 = ~n21181 & ~n21370;
  assign n21372 = ~n21369 & n21371;
  assign n21373 = ~n21181 & ~n21372;
  assign n21374 = ~n21076 & ~n21176;
  assign n21375 = ~n21178 & ~n21374;
  assign n21376 = ~n21373 & n21375;
  assign n21377 = ~n21178 & ~n21376;
  assign n21378 = ~n21169 & ~n21174;
  assign n21379 = n4783 & n12606;
  assign n21380 = n4801 & ~n12608;
  assign n21381 = ~n12611 & n21380;
  assign n21382 = n4601 & n12614;
  assign n21383 = n4602 & n12868;
  assign n21384 = ~n21382 & ~n21383;
  assign n21385 = ~n21381 & n21384;
  assign n21386 = ~n21379 & n21385;
  assign n21387 = pi26  & n21386;
  assign n21388 = ~pi26  & ~n21386;
  assign n21389 = ~n21387 & ~n21388;
  assign n21390 = ~n21148 & n21160;
  assign n21391 = ~n21149 & ~n21390;
  assign n21392 = n21389 & n21391;
  assign n21393 = ~n21389 & ~n21391;
  assign n21394 = ~n21392 & ~n21393;
  assign n21395 = ~n21142 & ~n21145;
  assign n21396 = n5236 & n5237;
  assign n21397 = ~n12608 & ~n21396;
  assign n21398 = pi23  & ~n21397;
  assign n21399 = ~pi23  & n21397;
  assign n21400 = ~n21398 & ~n21399;
  assign n21401 = n848 & n13877;
  assign n21402 = ~n612 & n21401;
  assign n21403 = ~n362 & n15344;
  assign n21404 = ~n668 & n21403;
  assign n21405 = n21402 & n21404;
  assign n21406 = n5527 & n13087;
  assign n21407 = n1186 & n21406;
  assign n21408 = ~n334 & n21407;
  assign n21409 = n1086 & n7113;
  assign n21410 = n4353 & n21409;
  assign n21411 = n1652 & n21410;
  assign n21412 = n386 & n21411;
  assign n21413 = ~n441 & n21412;
  assign n21414 = ~n150 & n21413;
  assign n21415 = n21408 & n21414;
  assign n21416 = n21405 & n21415;
  assign n21417 = n21128 & n21416;
  assign n21418 = ~n21128 & ~n21416;
  assign n21419 = ~n21417 & ~n21418;
  assign n21420 = n21400 & n21419;
  assign n21421 = ~n21400 & ~n21419;
  assign n21422 = ~n21420 & ~n21421;
  assign n21423 = n21103 & ~n21129;
  assign n21424 = ~n21130 & ~n21423;
  assign n21425 = n21422 & n21424;
  assign n21426 = ~n21422 & ~n21424;
  assign n21427 = ~n21425 & ~n21426;
  assign n21428 = n3641 & n12639;
  assign n21429 = n3740 & n12636;
  assign n21430 = n556 & n13396;
  assign n21431 = n3961 & n12633;
  assign n21432 = ~n21430 & ~n21431;
  assign n21433 = ~n21429 & n21432;
  assign n21434 = ~n21428 & n21433;
  assign n21435 = n21427 & ~n21434;
  assign n21436 = ~n21427 & n21434;
  assign n21437 = ~n21435 & ~n21436;
  assign n21438 = n21395 & ~n21437;
  assign n21439 = ~n21395 & n21437;
  assign n21440 = ~n21438 & ~n21439;
  assign n21441 = n4006 & n12630;
  assign n21442 = n4133 & n12625;
  assign n21443 = n4002 & n13325;
  assign n21444 = n4555 & n12622;
  assign n21445 = ~n21443 & ~n21444;
  assign n21446 = ~n21442 & n21445;
  assign n21447 = ~n21441 & n21446;
  assign n21448 = pi29  & n21447;
  assign n21449 = ~pi29  & ~n21447;
  assign n21450 = ~n21448 & ~n21449;
  assign n21451 = n21440 & ~n21450;
  assign n21452 = ~n21440 & n21450;
  assign n21453 = ~n21451 & ~n21452;
  assign n21454 = ~n21394 & n21453;
  assign n21455 = n21394 & ~n21453;
  assign n21456 = ~n21454 & ~n21455;
  assign n21457 = ~n21089 & ~n21163;
  assign n21458 = ~n21090 & ~n21457;
  assign n21459 = n21456 & n21458;
  assign n21460 = ~n21456 & ~n21458;
  assign n21461 = ~n21459 & ~n21460;
  assign n21462 = ~n21378 & n21461;
  assign n21463 = n21378 & ~n21461;
  assign n21464 = ~n21462 & ~n21463;
  assign n21465 = n21176 & n21464;
  assign n21466 = ~n21176 & ~n21464;
  assign n21467 = ~n21465 & ~n21466;
  assign n21468 = n21377 & n21467;
  assign n21469 = ~n21377 & ~n21467;
  assign n21470 = ~n21468 & ~n21469;
  assign n21471 = n9719 & ~n21470;
  assign n21472 = n11267 & n21464;
  assign n21473 = ~n21471 & ~n21472;
  assign n21474 = ~n21177 & n21473;
  assign n21475 = ~n21077 & n21474;
  assign n21476 = ~pi5  & ~n21475;
  assign n21477 = pi5  & n21475;
  assign n21478 = ~n21476 & ~n21477;
  assign n21479 = n7654 & n21201;
  assign n21480 = n8091 & n21198;
  assign n21481 = n21345 & ~n21347;
  assign n21482 = ~n21348 & ~n21481;
  assign n21483 = n7648 & n21482;
  assign n21484 = n8120 & n21195;
  assign n21485 = ~n21483 & ~n21484;
  assign n21486 = ~n21480 & n21485;
  assign n21487 = ~n21479 & n21486;
  assign n21488 = ~pi11  & ~n21487;
  assign n21489 = pi11  & n21487;
  assign n21490 = ~n21488 & ~n21489;
  assign n21491 = n5435 & n21234;
  assign n21492 = n6055 & n21231;
  assign n21493 = n21301 & ~n21303;
  assign n21494 = ~n21304 & ~n21493;
  assign n21495 = n5429 & n21494;
  assign n21496 = n6071 & n21228;
  assign n21497 = ~n21495 & ~n21496;
  assign n21498 = ~n21492 & n21497;
  assign n21499 = ~n21491 & n21498;
  assign n21500 = ~pi20  & ~n21499;
  assign n21501 = pi20  & n21499;
  assign n21502 = ~n21500 & ~n21501;
  assign n21503 = n4601 & n21255;
  assign n21504 = n4783 & n21252;
  assign n21505 = n21273 & ~n21275;
  assign n21506 = ~n21276 & ~n21505;
  assign n21507 = n4602 & n21506;
  assign n21508 = n4801 & n21249;
  assign n21509 = ~n21507 & ~n21508;
  assign n21510 = ~n21504 & n21509;
  assign n21511 = ~n21503 & n21510;
  assign n21512 = ~pi26  & ~n21511;
  assign n21513 = pi26  & n21511;
  assign n21514 = ~n21512 & ~n21513;
  assign n21515 = ~n3998 & n21265;
  assign n21516 = pi29  & ~n21515;
  assign n21517 = n21263 & ~n21265;
  assign n21518 = ~n21263 & n21265;
  assign n21519 = ~n21517 & ~n21518;
  assign n21520 = n4002 & ~n21519;
  assign n21521 = n4555 & n21263;
  assign n21522 = n4133 & n21265;
  assign n21523 = ~n21521 & ~n21522;
  assign n21524 = ~n21520 & n21523;
  assign n21525 = n21516 & n21524;
  assign n21526 = pi29  & ~n21525;
  assign n21527 = n4006 & n21265;
  assign n21528 = n4133 & n21263;
  assign n21529 = n21258 & ~n21517;
  assign n21530 = ~n21258 & n21517;
  assign n21531 = ~n21529 & ~n21530;
  assign n21532 = n4002 & ~n21531;
  assign n21533 = n4555 & n21258;
  assign n21534 = ~n21532 & ~n21533;
  assign n21535 = ~n21528 & n21534;
  assign n21536 = ~n21527 & n21535;
  assign n21537 = ~n21526 & n21536;
  assign n21538 = n21526 & ~n21536;
  assign n21539 = ~n21537 & ~n21538;
  assign n21540 = ~n21514 & ~n21539;
  assign n21541 = n21514 & n21539;
  assign n21542 = ~n21540 & ~n21541;
  assign n21543 = n4601 & n21258;
  assign n21544 = n4783 & n21255;
  assign n21545 = n21269 & ~n21271;
  assign n21546 = ~n21272 & ~n21545;
  assign n21547 = n4602 & n21546;
  assign n21548 = n4801 & n21252;
  assign n21549 = ~n21547 & ~n21548;
  assign n21550 = ~n21544 & n21549;
  assign n21551 = ~n21543 & n21550;
  assign n21552 = pi26  & n21551;
  assign n21553 = ~pi26  & ~n21551;
  assign n21554 = ~n21552 & ~n21553;
  assign n21555 = pi29  & n21515;
  assign n21556 = ~n21524 & n21555;
  assign n21557 = n21524 & ~n21555;
  assign n21558 = ~n21556 & ~n21557;
  assign n21559 = ~n21554 & n21558;
  assign n21560 = ~n4598 & n21265;
  assign n21561 = pi26  & ~n21560;
  assign n21562 = n4602 & ~n21519;
  assign n21563 = n4801 & n21263;
  assign n21564 = n4783 & n21265;
  assign n21565 = ~n21563 & ~n21564;
  assign n21566 = ~n21562 & n21565;
  assign n21567 = n21561 & n21566;
  assign n21568 = n4601 & n21265;
  assign n21569 = n4783 & n21263;
  assign n21570 = n4602 & ~n21531;
  assign n21571 = n4801 & n21258;
  assign n21572 = ~n21570 & ~n21571;
  assign n21573 = ~n21569 & n21572;
  assign n21574 = ~n21568 & n21573;
  assign n21575 = n21567 & n21574;
  assign n21576 = n21515 & n21575;
  assign n21577 = ~n21515 & n21575;
  assign n21578 = n21515 & ~n21575;
  assign n21579 = ~n21577 & ~n21578;
  assign n21580 = n4601 & n21263;
  assign n21581 = n4783 & n21258;
  assign n21582 = ~n21261 & ~n21267;
  assign n21583 = ~n21268 & ~n21582;
  assign n21584 = n4602 & n21583;
  assign n21585 = n4801 & n21255;
  assign n21586 = ~n21584 & ~n21585;
  assign n21587 = ~n21581 & n21586;
  assign n21588 = ~n21580 & n21587;
  assign n21589 = pi26  & n21588;
  assign n21590 = ~pi26  & ~n21588;
  assign n21591 = ~n21589 & ~n21590;
  assign n21592 = ~n21579 & ~n21591;
  assign n21593 = ~n21576 & ~n21592;
  assign n21594 = n21554 & ~n21558;
  assign n21595 = ~n21559 & ~n21594;
  assign n21596 = ~n21593 & n21595;
  assign n21597 = ~n21559 & ~n21596;
  assign n21598 = ~n21542 & ~n21597;
  assign n21599 = n21542 & n21597;
  assign n21600 = ~n21598 & ~n21599;
  assign n21601 = n5238 & n21246;
  assign n21602 = n71 & n21243;
  assign n21603 = n21285 & ~n21287;
  assign n21604 = ~n21288 & ~n21603;
  assign n21605 = n5239 & n21604;
  assign n21606 = n5326 & n21240;
  assign n21607 = ~n21605 & ~n21606;
  assign n21608 = ~n21602 & n21607;
  assign n21609 = ~n21601 & n21608;
  assign n21610 = pi23  & n21609;
  assign n21611 = ~pi23  & ~n21609;
  assign n21612 = ~n21610 & ~n21611;
  assign n21613 = n21600 & ~n21612;
  assign n21614 = n5238 & n21249;
  assign n21615 = n71 & n21246;
  assign n21616 = n21281 & ~n21283;
  assign n21617 = ~n21284 & ~n21616;
  assign n21618 = n5239 & n21617;
  assign n21619 = n5326 & n21243;
  assign n21620 = ~n21618 & ~n21619;
  assign n21621 = ~n21615 & n21620;
  assign n21622 = ~n21614 & n21621;
  assign n21623 = ~pi23  & ~n21622;
  assign n21624 = pi23  & n21622;
  assign n21625 = ~n21623 & ~n21624;
  assign n21626 = n21593 & ~n21595;
  assign n21627 = ~n21596 & ~n21626;
  assign n21628 = ~n21625 & n21627;
  assign n21629 = ~n21625 & ~n21627;
  assign n21630 = n21625 & n21627;
  assign n21631 = ~n21629 & ~n21630;
  assign n21632 = n5238 & n21252;
  assign n21633 = n71 & n21249;
  assign n21634 = n21277 & ~n21279;
  assign n21635 = ~n21280 & ~n21634;
  assign n21636 = n5239 & n21635;
  assign n21637 = n5326 & n21246;
  assign n21638 = ~n21636 & ~n21637;
  assign n21639 = ~n21633 & n21638;
  assign n21640 = ~n21632 & n21639;
  assign n21641 = pi23  & n21640;
  assign n21642 = ~pi23  & ~n21640;
  assign n21643 = ~n21641 & ~n21642;
  assign n21644 = n21579 & n21591;
  assign n21645 = ~n21592 & ~n21644;
  assign n21646 = ~n21643 & n21645;
  assign n21647 = n5238 & n21255;
  assign n21648 = n71 & n21252;
  assign n21649 = n5239 & n21506;
  assign n21650 = n5326 & n21249;
  assign n21651 = ~n21649 & ~n21650;
  assign n21652 = ~n21648 & n21651;
  assign n21653 = ~n21647 & n21652;
  assign n21654 = ~pi23  & ~n21653;
  assign n21655 = pi23  & n21653;
  assign n21656 = ~n21654 & ~n21655;
  assign n21657 = pi26  & ~n21567;
  assign n21658 = n21574 & ~n21657;
  assign n21659 = ~n21574 & n21657;
  assign n21660 = ~n21658 & ~n21659;
  assign n21661 = ~n21656 & n21660;
  assign n21662 = ~n21656 & ~n21660;
  assign n21663 = n21656 & n21660;
  assign n21664 = ~n21662 & ~n21663;
  assign n21665 = n5238 & n21258;
  assign n21666 = n71 & n21255;
  assign n21667 = n5239 & n21546;
  assign n21668 = n5326 & n21252;
  assign n21669 = ~n21667 & ~n21668;
  assign n21670 = ~n21666 & n21669;
  assign n21671 = ~n21665 & n21670;
  assign n21672 = pi23  & n21671;
  assign n21673 = ~pi23  & ~n21671;
  assign n21674 = ~n21672 & ~n21673;
  assign n21675 = pi26  & n21560;
  assign n21676 = ~n21566 & n21675;
  assign n21677 = n21566 & ~n21675;
  assign n21678 = ~n21676 & ~n21677;
  assign n21679 = ~n21674 & n21678;
  assign n21680 = ~n70 & n21265;
  assign n21681 = pi23  & ~n21680;
  assign n21682 = n5239 & ~n21519;
  assign n21683 = n5326 & n21263;
  assign n21684 = n71 & n21265;
  assign n21685 = ~n21683 & ~n21684;
  assign n21686 = ~n21682 & n21685;
  assign n21687 = n21681 & n21686;
  assign n21688 = n5238 & n21265;
  assign n21689 = n71 & n21263;
  assign n21690 = n5239 & ~n21531;
  assign n21691 = n5326 & n21258;
  assign n21692 = ~n21690 & ~n21691;
  assign n21693 = ~n21689 & n21692;
  assign n21694 = ~n21688 & n21693;
  assign n21695 = n21687 & n21694;
  assign n21696 = n21560 & n21695;
  assign n21697 = ~n21560 & n21695;
  assign n21698 = n21560 & ~n21695;
  assign n21699 = ~n21697 & ~n21698;
  assign n21700 = n5238 & n21263;
  assign n21701 = n71 & n21258;
  assign n21702 = n5239 & n21583;
  assign n21703 = n5326 & n21255;
  assign n21704 = ~n21702 & ~n21703;
  assign n21705 = ~n21701 & n21704;
  assign n21706 = ~n21700 & n21705;
  assign n21707 = pi23  & n21706;
  assign n21708 = ~pi23  & ~n21706;
  assign n21709 = ~n21707 & ~n21708;
  assign n21710 = ~n21699 & ~n21709;
  assign n21711 = ~n21696 & ~n21710;
  assign n21712 = n21674 & ~n21678;
  assign n21713 = ~n21679 & ~n21712;
  assign n21714 = ~n21711 & n21713;
  assign n21715 = ~n21679 & ~n21714;
  assign n21716 = ~n21664 & ~n21715;
  assign n21717 = ~n21661 & ~n21716;
  assign n21718 = n21643 & ~n21645;
  assign n21719 = ~n21646 & ~n21718;
  assign n21720 = ~n21717 & n21719;
  assign n21721 = ~n21646 & ~n21720;
  assign n21722 = ~n21631 & ~n21721;
  assign n21723 = ~n21628 & ~n21722;
  assign n21724 = n21600 & n21612;
  assign n21725 = ~n21600 & ~n21612;
  assign n21726 = ~n21724 & ~n21725;
  assign n21727 = ~n21723 & ~n21726;
  assign n21728 = ~n21613 & ~n21727;
  assign n21729 = n4601 & n21252;
  assign n21730 = n4783 & n21249;
  assign n21731 = n4602 & n21635;
  assign n21732 = n4801 & n21246;
  assign n21733 = ~n21731 & ~n21732;
  assign n21734 = ~n21730 & n21733;
  assign n21735 = ~n21729 & n21734;
  assign n21736 = ~pi26  & ~n21735;
  assign n21737 = pi26  & n21735;
  assign n21738 = ~n21736 & ~n21737;
  assign n21739 = n4006 & n21263;
  assign n21740 = n4133 & n21258;
  assign n21741 = n4002 & n21583;
  assign n21742 = n4555 & n21255;
  assign n21743 = ~n21741 & ~n21742;
  assign n21744 = ~n21740 & n21743;
  assign n21745 = ~n21739 & n21744;
  assign n21746 = ~pi29  & ~n21745;
  assign n21747 = pi29  & n21745;
  assign n21748 = ~n21746 & ~n21747;
  assign n21749 = n21525 & n21536;
  assign n21750 = ~n555 & n21265;
  assign n21751 = n21749 & ~n21750;
  assign n21752 = ~n21749 & n21750;
  assign n21753 = ~n21751 & ~n21752;
  assign n21754 = ~n21748 & ~n21753;
  assign n21755 = n21748 & n21753;
  assign n21756 = ~n21754 & ~n21755;
  assign n21757 = ~n21738 & ~n21756;
  assign n21758 = n21738 & n21756;
  assign n21759 = ~n21757 & ~n21758;
  assign n21760 = ~n21514 & n21539;
  assign n21761 = ~n21598 & ~n21760;
  assign n21762 = ~n21759 & ~n21761;
  assign n21763 = n21759 & n21761;
  assign n21764 = ~n21762 & ~n21763;
  assign n21765 = n5238 & n21243;
  assign n21766 = n71 & n21240;
  assign n21767 = n21289 & ~n21291;
  assign n21768 = ~n21292 & ~n21767;
  assign n21769 = n5239 & n21768;
  assign n21770 = n5326 & n21237;
  assign n21771 = ~n21769 & ~n21770;
  assign n21772 = ~n21766 & n21771;
  assign n21773 = ~n21765 & n21772;
  assign n21774 = pi23  & n21773;
  assign n21775 = ~pi23  & ~n21773;
  assign n21776 = ~n21774 & ~n21775;
  assign n21777 = n21764 & ~n21776;
  assign n21778 = ~n21764 & n21776;
  assign n21779 = ~n21777 & ~n21778;
  assign n21780 = ~n21728 & n21779;
  assign n21781 = n21728 & ~n21779;
  assign n21782 = ~n21780 & ~n21781;
  assign n21783 = ~n21502 & ~n21782;
  assign n21784 = n21502 & n21782;
  assign n21785 = ~n21783 & ~n21784;
  assign n21786 = n5435 & n21237;
  assign n21787 = n6055 & n21234;
  assign n21788 = n21297 & ~n21299;
  assign n21789 = ~n21300 & ~n21788;
  assign n21790 = n5429 & n21789;
  assign n21791 = n6071 & n21231;
  assign n21792 = ~n21790 & ~n21791;
  assign n21793 = ~n21787 & n21792;
  assign n21794 = ~n21786 & n21793;
  assign n21795 = ~pi20  & ~n21794;
  assign n21796 = pi20  & n21794;
  assign n21797 = ~n21795 & ~n21796;
  assign n21798 = ~n21723 & n21726;
  assign n21799 = n21723 & ~n21726;
  assign n21800 = ~n21798 & ~n21799;
  assign n21801 = ~n21797 & ~n21800;
  assign n21802 = n21631 & n21721;
  assign n21803 = ~n21722 & ~n21802;
  assign n21804 = n5435 & n21240;
  assign n21805 = n6055 & n21237;
  assign n21806 = n21293 & ~n21295;
  assign n21807 = ~n21296 & ~n21806;
  assign n21808 = n5429 & n21807;
  assign n21809 = n6071 & n21234;
  assign n21810 = ~n21808 & ~n21809;
  assign n21811 = ~n21805 & n21810;
  assign n21812 = ~n21804 & n21811;
  assign n21813 = pi20  & n21812;
  assign n21814 = ~pi20  & ~n21812;
  assign n21815 = ~n21813 & ~n21814;
  assign n21816 = n21803 & ~n21815;
  assign n21817 = n21717 & ~n21719;
  assign n21818 = ~n21720 & ~n21817;
  assign n21819 = n5435 & n21243;
  assign n21820 = n6055 & n21240;
  assign n21821 = n5429 & n21768;
  assign n21822 = n6071 & n21237;
  assign n21823 = ~n21821 & ~n21822;
  assign n21824 = ~n21820 & n21823;
  assign n21825 = ~n21819 & n21824;
  assign n21826 = pi20  & n21825;
  assign n21827 = ~pi20  & ~n21825;
  assign n21828 = ~n21826 & ~n21827;
  assign n21829 = n21818 & ~n21828;
  assign n21830 = n21664 & n21715;
  assign n21831 = ~n21716 & ~n21830;
  assign n21832 = n5435 & n21246;
  assign n21833 = n6055 & n21243;
  assign n21834 = n5429 & n21604;
  assign n21835 = n6071 & n21240;
  assign n21836 = ~n21834 & ~n21835;
  assign n21837 = ~n21833 & n21836;
  assign n21838 = ~n21832 & n21837;
  assign n21839 = pi20  & n21838;
  assign n21840 = ~pi20  & ~n21838;
  assign n21841 = ~n21839 & ~n21840;
  assign n21842 = n21831 & ~n21841;
  assign n21843 = n5435 & n21249;
  assign n21844 = n6055 & n21246;
  assign n21845 = n5429 & n21617;
  assign n21846 = n6071 & n21243;
  assign n21847 = ~n21845 & ~n21846;
  assign n21848 = ~n21844 & n21847;
  assign n21849 = ~n21843 & n21848;
  assign n21850 = ~pi20  & ~n21849;
  assign n21851 = pi20  & n21849;
  assign n21852 = ~n21850 & ~n21851;
  assign n21853 = n21711 & ~n21713;
  assign n21854 = ~n21714 & ~n21853;
  assign n21855 = ~n21852 & n21854;
  assign n21856 = ~n21852 & ~n21854;
  assign n21857 = n21852 & n21854;
  assign n21858 = ~n21856 & ~n21857;
  assign n21859 = n5435 & n21252;
  assign n21860 = n6055 & n21249;
  assign n21861 = n5429 & n21635;
  assign n21862 = n6071 & n21246;
  assign n21863 = ~n21861 & ~n21862;
  assign n21864 = ~n21860 & n21863;
  assign n21865 = ~n21859 & n21864;
  assign n21866 = pi20  & n21865;
  assign n21867 = ~pi20  & ~n21865;
  assign n21868 = ~n21866 & ~n21867;
  assign n21869 = n21699 & n21709;
  assign n21870 = ~n21710 & ~n21869;
  assign n21871 = ~n21868 & n21870;
  assign n21872 = n5435 & n21255;
  assign n21873 = n6055 & n21252;
  assign n21874 = n5429 & n21506;
  assign n21875 = n6071 & n21249;
  assign n21876 = ~n21874 & ~n21875;
  assign n21877 = ~n21873 & n21876;
  assign n21878 = ~n21872 & n21877;
  assign n21879 = ~pi20  & ~n21878;
  assign n21880 = pi20  & n21878;
  assign n21881 = ~n21879 & ~n21880;
  assign n21882 = pi23  & ~n21687;
  assign n21883 = n21694 & ~n21882;
  assign n21884 = ~n21694 & n21882;
  assign n21885 = ~n21883 & ~n21884;
  assign n21886 = ~n21881 & n21885;
  assign n21887 = ~n21881 & ~n21885;
  assign n21888 = n21881 & n21885;
  assign n21889 = ~n21887 & ~n21888;
  assign n21890 = n5435 & n21258;
  assign n21891 = n6055 & n21255;
  assign n21892 = n5429 & n21546;
  assign n21893 = n6071 & n21252;
  assign n21894 = ~n21892 & ~n21893;
  assign n21895 = ~n21891 & n21894;
  assign n21896 = ~n21890 & n21895;
  assign n21897 = pi20  & n21896;
  assign n21898 = ~pi20  & ~n21896;
  assign n21899 = ~n21897 & ~n21898;
  assign n21900 = pi23  & n21680;
  assign n21901 = ~n21686 & n21900;
  assign n21902 = n21686 & ~n21900;
  assign n21903 = ~n21901 & ~n21902;
  assign n21904 = ~n21899 & n21903;
  assign n21905 = n5429 & ~n21519;
  assign n21906 = n6071 & n21263;
  assign n21907 = n6055 & n21265;
  assign n21908 = ~n21906 & ~n21907;
  assign n21909 = ~n21905 & n21908;
  assign n21910 = ~n5425 & n21265;
  assign n21911 = pi20  & ~n21910;
  assign n21912 = n21909 & n21911;
  assign n21913 = n5435 & n21265;
  assign n21914 = n6055 & n21263;
  assign n21915 = n5429 & ~n21531;
  assign n21916 = n6071 & n21258;
  assign n21917 = ~n21915 & ~n21916;
  assign n21918 = ~n21914 & n21917;
  assign n21919 = ~n21913 & n21918;
  assign n21920 = n21912 & n21919;
  assign n21921 = n21680 & n21920;
  assign n21922 = ~n21680 & n21920;
  assign n21923 = n21680 & ~n21920;
  assign n21924 = ~n21922 & ~n21923;
  assign n21925 = n5435 & n21263;
  assign n21926 = n6055 & n21258;
  assign n21927 = n5429 & n21583;
  assign n21928 = n6071 & n21255;
  assign n21929 = ~n21927 & ~n21928;
  assign n21930 = ~n21926 & n21929;
  assign n21931 = ~n21925 & n21930;
  assign n21932 = pi20  & n21931;
  assign n21933 = ~pi20  & ~n21931;
  assign n21934 = ~n21932 & ~n21933;
  assign n21935 = ~n21924 & ~n21934;
  assign n21936 = ~n21921 & ~n21935;
  assign n21937 = n21899 & ~n21903;
  assign n21938 = ~n21904 & ~n21937;
  assign n21939 = ~n21936 & n21938;
  assign n21940 = ~n21904 & ~n21939;
  assign n21941 = ~n21889 & ~n21940;
  assign n21942 = ~n21886 & ~n21941;
  assign n21943 = n21868 & ~n21870;
  assign n21944 = ~n21871 & ~n21943;
  assign n21945 = ~n21942 & n21944;
  assign n21946 = ~n21871 & ~n21945;
  assign n21947 = ~n21858 & ~n21946;
  assign n21948 = ~n21855 & ~n21947;
  assign n21949 = n21831 & n21841;
  assign n21950 = ~n21831 & ~n21841;
  assign n21951 = ~n21949 & ~n21950;
  assign n21952 = ~n21948 & ~n21951;
  assign n21953 = ~n21842 & ~n21952;
  assign n21954 = n21818 & n21828;
  assign n21955 = ~n21818 & ~n21828;
  assign n21956 = ~n21954 & ~n21955;
  assign n21957 = ~n21953 & ~n21956;
  assign n21958 = ~n21829 & ~n21957;
  assign n21959 = ~n21803 & n21815;
  assign n21960 = ~n21816 & ~n21959;
  assign n21961 = ~n21958 & n21960;
  assign n21962 = ~n21816 & ~n21961;
  assign n21963 = n21797 & n21800;
  assign n21964 = ~n21801 & ~n21963;
  assign n21965 = ~n21962 & n21964;
  assign n21966 = ~n21801 & ~n21965;
  assign n21967 = ~n21785 & ~n21966;
  assign n21968 = n21785 & n21966;
  assign n21969 = ~n21967 & ~n21968;
  assign n21970 = n6184 & n21225;
  assign n21971 = n6527 & n21222;
  assign n21972 = n21313 & ~n21315;
  assign n21973 = ~n21316 & ~n21972;
  assign n21974 = n6185 & n21973;
  assign n21975 = n6543 & n21219;
  assign n21976 = ~n21974 & ~n21975;
  assign n21977 = ~n21971 & n21976;
  assign n21978 = ~n21970 & n21977;
  assign n21979 = pi17  & n21978;
  assign n21980 = ~pi17  & ~n21978;
  assign n21981 = ~n21979 & ~n21980;
  assign n21982 = n21969 & ~n21981;
  assign n21983 = n21962 & ~n21964;
  assign n21984 = ~n21965 & ~n21983;
  assign n21985 = n6184 & n21228;
  assign n21986 = n6527 & n21225;
  assign n21987 = n21309 & ~n21311;
  assign n21988 = ~n21312 & ~n21987;
  assign n21989 = n6185 & n21988;
  assign n21990 = n6543 & n21222;
  assign n21991 = ~n21989 & ~n21990;
  assign n21992 = ~n21986 & n21991;
  assign n21993 = ~n21985 & n21992;
  assign n21994 = pi17  & n21993;
  assign n21995 = ~pi17  & ~n21993;
  assign n21996 = ~n21994 & ~n21995;
  assign n21997 = n21984 & ~n21996;
  assign n21998 = n6184 & n21231;
  assign n21999 = n6527 & n21228;
  assign n22000 = n21305 & ~n21307;
  assign n22001 = ~n21308 & ~n22000;
  assign n22002 = n6185 & n22001;
  assign n22003 = n6543 & n21225;
  assign n22004 = ~n22002 & ~n22003;
  assign n22005 = ~n21999 & n22004;
  assign n22006 = ~n21998 & n22005;
  assign n22007 = ~pi17  & ~n22006;
  assign n22008 = pi17  & n22006;
  assign n22009 = ~n22007 & ~n22008;
  assign n22010 = n21958 & ~n21960;
  assign n22011 = ~n21961 & ~n22010;
  assign n22012 = ~n22009 & n22011;
  assign n22013 = ~n22009 & ~n22011;
  assign n22014 = n22009 & n22011;
  assign n22015 = ~n22013 & ~n22014;
  assign n22016 = n6184 & n21234;
  assign n22017 = n6527 & n21231;
  assign n22018 = n6185 & n21494;
  assign n22019 = n6543 & n21228;
  assign n22020 = ~n22018 & ~n22019;
  assign n22021 = ~n22017 & n22020;
  assign n22022 = ~n22016 & n22021;
  assign n22023 = ~pi17  & ~n22022;
  assign n22024 = pi17  & n22022;
  assign n22025 = ~n22023 & ~n22024;
  assign n22026 = n21953 & n21956;
  assign n22027 = ~n21957 & ~n22026;
  assign n22028 = ~n22025 & n22027;
  assign n22029 = ~n22025 & ~n22027;
  assign n22030 = n22025 & n22027;
  assign n22031 = ~n22029 & ~n22030;
  assign n22032 = n6184 & n21237;
  assign n22033 = n6527 & n21234;
  assign n22034 = n6185 & n21789;
  assign n22035 = n6543 & n21231;
  assign n22036 = ~n22034 & ~n22035;
  assign n22037 = ~n22033 & n22036;
  assign n22038 = ~n22032 & n22037;
  assign n22039 = ~pi17  & ~n22038;
  assign n22040 = pi17  & n22038;
  assign n22041 = ~n22039 & ~n22040;
  assign n22042 = ~n21948 & n21951;
  assign n22043 = n21948 & ~n21951;
  assign n22044 = ~n22042 & ~n22043;
  assign n22045 = ~n22041 & ~n22044;
  assign n22046 = n21858 & n21946;
  assign n22047 = ~n21947 & ~n22046;
  assign n22048 = n6184 & n21240;
  assign n22049 = n6527 & n21237;
  assign n22050 = n6185 & n21807;
  assign n22051 = n6543 & n21234;
  assign n22052 = ~n22050 & ~n22051;
  assign n22053 = ~n22049 & n22052;
  assign n22054 = ~n22048 & n22053;
  assign n22055 = pi17  & n22054;
  assign n22056 = ~pi17  & ~n22054;
  assign n22057 = ~n22055 & ~n22056;
  assign n22058 = n22047 & ~n22057;
  assign n22059 = n21942 & ~n21944;
  assign n22060 = ~n21945 & ~n22059;
  assign n22061 = n6184 & n21243;
  assign n22062 = n6527 & n21240;
  assign n22063 = n6185 & n21768;
  assign n22064 = n6543 & n21237;
  assign n22065 = ~n22063 & ~n22064;
  assign n22066 = ~n22062 & n22065;
  assign n22067 = ~n22061 & n22066;
  assign n22068 = pi17  & n22067;
  assign n22069 = ~pi17  & ~n22067;
  assign n22070 = ~n22068 & ~n22069;
  assign n22071 = n22060 & ~n22070;
  assign n22072 = n21889 & n21940;
  assign n22073 = ~n21941 & ~n22072;
  assign n22074 = n6184 & n21246;
  assign n22075 = n6527 & n21243;
  assign n22076 = n6185 & n21604;
  assign n22077 = n6543 & n21240;
  assign n22078 = ~n22076 & ~n22077;
  assign n22079 = ~n22075 & n22078;
  assign n22080 = ~n22074 & n22079;
  assign n22081 = pi17  & n22080;
  assign n22082 = ~pi17  & ~n22080;
  assign n22083 = ~n22081 & ~n22082;
  assign n22084 = n22073 & ~n22083;
  assign n22085 = n6184 & n21249;
  assign n22086 = n6527 & n21246;
  assign n22087 = n6185 & n21617;
  assign n22088 = n6543 & n21243;
  assign n22089 = ~n22087 & ~n22088;
  assign n22090 = ~n22086 & n22089;
  assign n22091 = ~n22085 & n22090;
  assign n22092 = ~pi17  & ~n22091;
  assign n22093 = pi17  & n22091;
  assign n22094 = ~n22092 & ~n22093;
  assign n22095 = n21936 & ~n21938;
  assign n22096 = ~n21939 & ~n22095;
  assign n22097 = ~n22094 & n22096;
  assign n22098 = ~n22094 & ~n22096;
  assign n22099 = n22094 & n22096;
  assign n22100 = ~n22098 & ~n22099;
  assign n22101 = n6184 & n21252;
  assign n22102 = n6527 & n21249;
  assign n22103 = n6185 & n21635;
  assign n22104 = n6543 & n21246;
  assign n22105 = ~n22103 & ~n22104;
  assign n22106 = ~n22102 & n22105;
  assign n22107 = ~n22101 & n22106;
  assign n22108 = pi17  & n22107;
  assign n22109 = ~pi17  & ~n22107;
  assign n22110 = ~n22108 & ~n22109;
  assign n22111 = n21924 & n21934;
  assign n22112 = ~n21935 & ~n22111;
  assign n22113 = ~n22110 & n22112;
  assign n22114 = n6184 & n21255;
  assign n22115 = n6527 & n21252;
  assign n22116 = n6185 & n21506;
  assign n22117 = n6543 & n21249;
  assign n22118 = ~n22116 & ~n22117;
  assign n22119 = ~n22115 & n22118;
  assign n22120 = ~n22114 & n22119;
  assign n22121 = ~pi17  & ~n22120;
  assign n22122 = pi17  & n22120;
  assign n22123 = ~n22121 & ~n22122;
  assign n22124 = pi20  & ~n21912;
  assign n22125 = n21919 & ~n22124;
  assign n22126 = ~n21919 & n22124;
  assign n22127 = ~n22125 & ~n22126;
  assign n22128 = ~n22123 & n22127;
  assign n22129 = ~n22123 & ~n22127;
  assign n22130 = n22123 & n22127;
  assign n22131 = ~n22129 & ~n22130;
  assign n22132 = n6184 & n21258;
  assign n22133 = n6527 & n21255;
  assign n22134 = n6185 & n21546;
  assign n22135 = n6543 & n21252;
  assign n22136 = ~n22134 & ~n22135;
  assign n22137 = ~n22133 & n22136;
  assign n22138 = ~n22132 & n22137;
  assign n22139 = pi17  & n22138;
  assign n22140 = ~pi17  & ~n22138;
  assign n22141 = ~n22139 & ~n22140;
  assign n22142 = pi20  & n21910;
  assign n22143 = ~n21909 & n22142;
  assign n22144 = n21909 & ~n22142;
  assign n22145 = ~n22143 & ~n22144;
  assign n22146 = ~n22141 & n22145;
  assign n22147 = n6185 & ~n21519;
  assign n22148 = n6543 & n21263;
  assign n22149 = n6527 & n21265;
  assign n22150 = ~n22148 & ~n22149;
  assign n22151 = ~n22147 & n22150;
  assign n22152 = ~n6182 & n21265;
  assign n22153 = pi17  & ~n22152;
  assign n22154 = n22151 & n22153;
  assign n22155 = n6184 & n21265;
  assign n22156 = n6527 & n21263;
  assign n22157 = n6185 & ~n21531;
  assign n22158 = n6543 & n21258;
  assign n22159 = ~n22157 & ~n22158;
  assign n22160 = ~n22156 & n22159;
  assign n22161 = ~n22155 & n22160;
  assign n22162 = n22154 & n22161;
  assign n22163 = n21910 & n22162;
  assign n22164 = ~n21910 & n22162;
  assign n22165 = n21910 & ~n22162;
  assign n22166 = ~n22164 & ~n22165;
  assign n22167 = n6184 & n21263;
  assign n22168 = n6527 & n21258;
  assign n22169 = n6185 & n21583;
  assign n22170 = n6543 & n21255;
  assign n22171 = ~n22169 & ~n22170;
  assign n22172 = ~n22168 & n22171;
  assign n22173 = ~n22167 & n22172;
  assign n22174 = pi17  & n22173;
  assign n22175 = ~pi17  & ~n22173;
  assign n22176 = ~n22174 & ~n22175;
  assign n22177 = ~n22166 & ~n22176;
  assign n22178 = ~n22163 & ~n22177;
  assign n22179 = n22141 & ~n22145;
  assign n22180 = ~n22146 & ~n22179;
  assign n22181 = ~n22178 & n22180;
  assign n22182 = ~n22146 & ~n22181;
  assign n22183 = ~n22131 & ~n22182;
  assign n22184 = ~n22128 & ~n22183;
  assign n22185 = n22110 & ~n22112;
  assign n22186 = ~n22113 & ~n22185;
  assign n22187 = ~n22184 & n22186;
  assign n22188 = ~n22113 & ~n22187;
  assign n22189 = ~n22100 & ~n22188;
  assign n22190 = ~n22097 & ~n22189;
  assign n22191 = n22073 & n22083;
  assign n22192 = ~n22073 & ~n22083;
  assign n22193 = ~n22191 & ~n22192;
  assign n22194 = ~n22190 & ~n22193;
  assign n22195 = ~n22084 & ~n22194;
  assign n22196 = n22060 & n22070;
  assign n22197 = ~n22060 & ~n22070;
  assign n22198 = ~n22196 & ~n22197;
  assign n22199 = ~n22195 & ~n22198;
  assign n22200 = ~n22071 & ~n22199;
  assign n22201 = ~n22047 & n22057;
  assign n22202 = ~n22058 & ~n22201;
  assign n22203 = ~n22200 & n22202;
  assign n22204 = ~n22058 & ~n22203;
  assign n22205 = n22041 & n22044;
  assign n22206 = ~n22045 & ~n22205;
  assign n22207 = ~n22204 & n22206;
  assign n22208 = ~n22045 & ~n22207;
  assign n22209 = ~n22031 & ~n22208;
  assign n22210 = ~n22028 & ~n22209;
  assign n22211 = ~n22015 & ~n22210;
  assign n22212 = ~n22012 & ~n22211;
  assign n22213 = n21984 & n21996;
  assign n22214 = ~n21984 & ~n21996;
  assign n22215 = ~n22213 & ~n22214;
  assign n22216 = ~n22212 & ~n22215;
  assign n22217 = ~n21997 & ~n22216;
  assign n22218 = ~n21969 & n21981;
  assign n22219 = ~n21982 & ~n22218;
  assign n22220 = ~n22217 & n22219;
  assign n22221 = ~n21982 & ~n22220;
  assign n22222 = n6184 & n21222;
  assign n22223 = n6527 & n21219;
  assign n22224 = n21317 & ~n21319;
  assign n22225 = ~n21320 & ~n22224;
  assign n22226 = n6185 & n22225;
  assign n22227 = n6543 & n21216;
  assign n22228 = ~n22226 & ~n22227;
  assign n22229 = ~n22223 & n22228;
  assign n22230 = ~n22222 & n22229;
  assign n22231 = ~pi17  & ~n22230;
  assign n22232 = pi17  & n22230;
  assign n22233 = ~n22231 & ~n22232;
  assign n22234 = ~n21502 & n21782;
  assign n22235 = ~n21967 & ~n22234;
  assign n22236 = n5238 & n21240;
  assign n22237 = n71 & n21237;
  assign n22238 = n5239 & n21807;
  assign n22239 = n5326 & n21234;
  assign n22240 = ~n22238 & ~n22239;
  assign n22241 = ~n22237 & n22240;
  assign n22242 = ~n22236 & n22241;
  assign n22243 = ~pi23  & ~n22242;
  assign n22244 = pi23  & n22242;
  assign n22245 = ~n22243 & ~n22244;
  assign n22246 = ~n21738 & n21756;
  assign n22247 = ~n21762 & ~n22246;
  assign n22248 = n4601 & n21249;
  assign n22249 = n4783 & n21246;
  assign n22250 = n4602 & n21617;
  assign n22251 = n4801 & n21243;
  assign n22252 = ~n22250 & ~n22251;
  assign n22253 = ~n22249 & n22252;
  assign n22254 = ~n22248 & n22253;
  assign n22255 = pi26  & n22254;
  assign n22256 = ~pi26  & ~n22254;
  assign n22257 = ~n22255 & ~n22256;
  assign n22258 = n21749 & n21750;
  assign n22259 = ~n21754 & ~n22258;
  assign n22260 = n4006 & n21258;
  assign n22261 = n4133 & n21255;
  assign n22262 = n4002 & n21546;
  assign n22263 = n4555 & n21252;
  assign n22264 = ~n22262 & ~n22263;
  assign n22265 = ~n22261 & n22264;
  assign n22266 = ~n22260 & n22265;
  assign n22267 = ~pi29  & ~n22266;
  assign n22268 = pi29  & n22266;
  assign n22269 = ~n22267 & ~n22268;
  assign n22270 = n3443 & n4874;
  assign n22271 = n1272 & n22270;
  assign n22272 = ~n204 & n22271;
  assign n22273 = n691 & n4260;
  assign n22274 = n1132 & n22273;
  assign n22275 = ~n400 & n22274;
  assign n22276 = n22272 & n22275;
  assign n22277 = n675 & n2929;
  assign n22278 = ~n161 & n22277;
  assign n22279 = n1641 & n13555;
  assign n22280 = n327 & n22279;
  assign n22281 = ~n112 & n22280;
  assign n22282 = n22278 & n22281;
  assign n22283 = n22276 & n22282;
  assign n22284 = n1186 & n22283;
  assign n22285 = n2056 & n22284;
  assign n22286 = n954 & n22285;
  assign n22287 = ~n154 & n22286;
  assign n22288 = ~n117 & n1791;
  assign n22289 = ~n533 & n22288;
  assign n22290 = n1111 & n1394;
  assign n22291 = ~n217 & n22290;
  assign n22292 = ~n132 & n22291;
  assign n22293 = n22289 & n22292;
  assign n22294 = ~n166 & n22293;
  assign n22295 = ~n337 & n1116;
  assign n22296 = ~n260 & n22295;
  assign n22297 = n257 & n22296;
  assign n22298 = n22294 & n22297;
  assign n22299 = n1368 & n22298;
  assign n22300 = ~n384 & n22299;
  assign n22301 = n22287 & n22300;
  assign n22302 = n1895 & n2829;
  assign n22303 = n1923 & n22302;
  assign n22304 = ~n152 & n22303;
  assign n22305 = n1700 & n15213;
  assign n22306 = n15136 & n22305;
  assign n22307 = n1902 & n22306;
  assign n22308 = n4085 & n22307;
  assign n22309 = n22304 & n22308;
  assign n22310 = n22301 & n22309;
  assign n22311 = n556 & ~n21519;
  assign n22312 = n3740 & n21265;
  assign n22313 = n3961 & n21263;
  assign n22314 = ~n22312 & ~n22313;
  assign n22315 = ~n22311 & n22314;
  assign n22316 = ~n22310 & n22315;
  assign n22317 = n22310 & ~n22315;
  assign n22318 = ~n22316 & ~n22317;
  assign n22319 = ~n22269 & ~n22318;
  assign n22320 = n22269 & n22318;
  assign n22321 = ~n22319 & ~n22320;
  assign n22322 = ~n22259 & n22321;
  assign n22323 = n22259 & ~n22321;
  assign n22324 = ~n22322 & ~n22323;
  assign n22325 = n22257 & n22324;
  assign n22326 = ~n22257 & ~n22324;
  assign n22327 = ~n22325 & ~n22326;
  assign n22328 = ~n22247 & ~n22327;
  assign n22329 = n22247 & n22327;
  assign n22330 = ~n22328 & ~n22329;
  assign n22331 = ~n22245 & ~n22330;
  assign n22332 = n22245 & n22330;
  assign n22333 = ~n22331 & ~n22332;
  assign n22334 = ~n21777 & ~n21780;
  assign n22335 = n22333 & n22334;
  assign n22336 = ~n22333 & ~n22334;
  assign n22337 = ~n22335 & ~n22336;
  assign n22338 = n5435 & n21231;
  assign n22339 = n6055 & n21228;
  assign n22340 = n5429 & n22001;
  assign n22341 = n6071 & n21225;
  assign n22342 = ~n22340 & ~n22341;
  assign n22343 = ~n22339 & n22342;
  assign n22344 = ~n22338 & n22343;
  assign n22345 = pi20  & n22344;
  assign n22346 = ~pi20  & ~n22344;
  assign n22347 = ~n22345 & ~n22346;
  assign n22348 = n22337 & n22347;
  assign n22349 = ~n22337 & ~n22347;
  assign n22350 = ~n22348 & ~n22349;
  assign n22351 = ~n22235 & n22350;
  assign n22352 = n22235 & ~n22350;
  assign n22353 = ~n22351 & ~n22352;
  assign n22354 = ~n22233 & ~n22353;
  assign n22355 = n22233 & n22353;
  assign n22356 = ~n22354 & ~n22355;
  assign n22357 = ~n22221 & n22356;
  assign n22358 = n22221 & ~n22356;
  assign n22359 = ~n22357 & ~n22358;
  assign n22360 = n6835 & n21213;
  assign n22361 = n7460 & n21210;
  assign n22362 = n21329 & ~n21331;
  assign n22363 = ~n21332 & ~n22362;
  assign n22364 = n6836 & n22363;
  assign n22365 = n7487 & n21207;
  assign n22366 = ~n22364 & ~n22365;
  assign n22367 = ~n22361 & n22366;
  assign n22368 = ~n22360 & n22367;
  assign n22369 = pi14  & n22368;
  assign n22370 = ~pi14  & ~n22368;
  assign n22371 = ~n22369 & ~n22370;
  assign n22372 = n22359 & ~n22371;
  assign n22373 = n6835 & n21216;
  assign n22374 = n7460 & n21213;
  assign n22375 = n21325 & ~n21327;
  assign n22376 = ~n21328 & ~n22375;
  assign n22377 = n6836 & n22376;
  assign n22378 = n7487 & n21210;
  assign n22379 = ~n22377 & ~n22378;
  assign n22380 = ~n22374 & n22379;
  assign n22381 = ~n22373 & n22380;
  assign n22382 = ~pi14  & ~n22381;
  assign n22383 = pi14  & n22381;
  assign n22384 = ~n22382 & ~n22383;
  assign n22385 = n22217 & ~n22219;
  assign n22386 = ~n22220 & ~n22385;
  assign n22387 = ~n22384 & n22386;
  assign n22388 = ~n22384 & ~n22386;
  assign n22389 = n22384 & n22386;
  assign n22390 = ~n22388 & ~n22389;
  assign n22391 = n6835 & n21219;
  assign n22392 = n7460 & n21216;
  assign n22393 = n21321 & ~n21323;
  assign n22394 = ~n21324 & ~n22393;
  assign n22395 = n6836 & n22394;
  assign n22396 = n7487 & n21213;
  assign n22397 = ~n22395 & ~n22396;
  assign n22398 = ~n22392 & n22397;
  assign n22399 = ~n22391 & n22398;
  assign n22400 = ~pi14  & ~n22399;
  assign n22401 = pi14  & n22399;
  assign n22402 = ~n22400 & ~n22401;
  assign n22403 = n22212 & n22215;
  assign n22404 = ~n22216 & ~n22403;
  assign n22405 = ~n22402 & n22404;
  assign n22406 = ~n22402 & ~n22404;
  assign n22407 = n22402 & n22404;
  assign n22408 = ~n22406 & ~n22407;
  assign n22409 = n22015 & n22210;
  assign n22410 = ~n22211 & ~n22409;
  assign n22411 = n6835 & n21222;
  assign n22412 = n7460 & n21219;
  assign n22413 = n6836 & n22225;
  assign n22414 = n7487 & n21216;
  assign n22415 = ~n22413 & ~n22414;
  assign n22416 = ~n22412 & n22415;
  assign n22417 = ~n22411 & n22416;
  assign n22418 = pi14  & n22417;
  assign n22419 = ~pi14  & ~n22417;
  assign n22420 = ~n22418 & ~n22419;
  assign n22421 = n22410 & ~n22420;
  assign n22422 = n22031 & n22208;
  assign n22423 = ~n22209 & ~n22422;
  assign n22424 = n6835 & n21225;
  assign n22425 = n7460 & n21222;
  assign n22426 = n6836 & n21973;
  assign n22427 = n7487 & n21219;
  assign n22428 = ~n22426 & ~n22427;
  assign n22429 = ~n22425 & n22428;
  assign n22430 = ~n22424 & n22429;
  assign n22431 = pi14  & n22430;
  assign n22432 = ~pi14  & ~n22430;
  assign n22433 = ~n22431 & ~n22432;
  assign n22434 = n22423 & ~n22433;
  assign n22435 = n22204 & ~n22206;
  assign n22436 = ~n22207 & ~n22435;
  assign n22437 = n6835 & n21228;
  assign n22438 = n7460 & n21225;
  assign n22439 = n6836 & n21988;
  assign n22440 = n7487 & n21222;
  assign n22441 = ~n22439 & ~n22440;
  assign n22442 = ~n22438 & n22441;
  assign n22443 = ~n22437 & n22442;
  assign n22444 = pi14  & n22443;
  assign n22445 = ~pi14  & ~n22443;
  assign n22446 = ~n22444 & ~n22445;
  assign n22447 = n22436 & ~n22446;
  assign n22448 = n6835 & n21231;
  assign n22449 = n7460 & n21228;
  assign n22450 = n6836 & n22001;
  assign n22451 = n7487 & n21225;
  assign n22452 = ~n22450 & ~n22451;
  assign n22453 = ~n22449 & n22452;
  assign n22454 = ~n22448 & n22453;
  assign n22455 = ~pi14  & ~n22454;
  assign n22456 = pi14  & n22454;
  assign n22457 = ~n22455 & ~n22456;
  assign n22458 = n22200 & ~n22202;
  assign n22459 = ~n22203 & ~n22458;
  assign n22460 = ~n22457 & n22459;
  assign n22461 = ~n22457 & ~n22459;
  assign n22462 = n22457 & n22459;
  assign n22463 = ~n22461 & ~n22462;
  assign n22464 = n6835 & n21234;
  assign n22465 = n7460 & n21231;
  assign n22466 = n6836 & n21494;
  assign n22467 = n7487 & n21228;
  assign n22468 = ~n22466 & ~n22467;
  assign n22469 = ~n22465 & n22468;
  assign n22470 = ~n22464 & n22469;
  assign n22471 = ~pi14  & ~n22470;
  assign n22472 = pi14  & n22470;
  assign n22473 = ~n22471 & ~n22472;
  assign n22474 = n22195 & n22198;
  assign n22475 = ~n22199 & ~n22474;
  assign n22476 = ~n22473 & n22475;
  assign n22477 = ~n22473 & ~n22475;
  assign n22478 = n22473 & n22475;
  assign n22479 = ~n22477 & ~n22478;
  assign n22480 = n6835 & n21237;
  assign n22481 = n7460 & n21234;
  assign n22482 = n6836 & n21789;
  assign n22483 = n7487 & n21231;
  assign n22484 = ~n22482 & ~n22483;
  assign n22485 = ~n22481 & n22484;
  assign n22486 = ~n22480 & n22485;
  assign n22487 = ~pi14  & ~n22486;
  assign n22488 = pi14  & n22486;
  assign n22489 = ~n22487 & ~n22488;
  assign n22490 = ~n22190 & n22193;
  assign n22491 = n22190 & ~n22193;
  assign n22492 = ~n22490 & ~n22491;
  assign n22493 = ~n22489 & ~n22492;
  assign n22494 = n22100 & n22188;
  assign n22495 = ~n22189 & ~n22494;
  assign n22496 = n6835 & n21240;
  assign n22497 = n7460 & n21237;
  assign n22498 = n6836 & n21807;
  assign n22499 = n7487 & n21234;
  assign n22500 = ~n22498 & ~n22499;
  assign n22501 = ~n22497 & n22500;
  assign n22502 = ~n22496 & n22501;
  assign n22503 = pi14  & n22502;
  assign n22504 = ~pi14  & ~n22502;
  assign n22505 = ~n22503 & ~n22504;
  assign n22506 = n22495 & ~n22505;
  assign n22507 = n22184 & ~n22186;
  assign n22508 = ~n22187 & ~n22507;
  assign n22509 = n6835 & n21243;
  assign n22510 = n7460 & n21240;
  assign n22511 = n6836 & n21768;
  assign n22512 = n7487 & n21237;
  assign n22513 = ~n22511 & ~n22512;
  assign n22514 = ~n22510 & n22513;
  assign n22515 = ~n22509 & n22514;
  assign n22516 = pi14  & n22515;
  assign n22517 = ~pi14  & ~n22515;
  assign n22518 = ~n22516 & ~n22517;
  assign n22519 = n22508 & ~n22518;
  assign n22520 = n22131 & n22182;
  assign n22521 = ~n22183 & ~n22520;
  assign n22522 = n6835 & n21246;
  assign n22523 = n7460 & n21243;
  assign n22524 = n6836 & n21604;
  assign n22525 = n7487 & n21240;
  assign n22526 = ~n22524 & ~n22525;
  assign n22527 = ~n22523 & n22526;
  assign n22528 = ~n22522 & n22527;
  assign n22529 = pi14  & n22528;
  assign n22530 = ~pi14  & ~n22528;
  assign n22531 = ~n22529 & ~n22530;
  assign n22532 = n22521 & ~n22531;
  assign n22533 = n6835 & n21249;
  assign n22534 = n7460 & n21246;
  assign n22535 = n6836 & n21617;
  assign n22536 = n7487 & n21243;
  assign n22537 = ~n22535 & ~n22536;
  assign n22538 = ~n22534 & n22537;
  assign n22539 = ~n22533 & n22538;
  assign n22540 = ~pi14  & ~n22539;
  assign n22541 = pi14  & n22539;
  assign n22542 = ~n22540 & ~n22541;
  assign n22543 = n22178 & ~n22180;
  assign n22544 = ~n22181 & ~n22543;
  assign n22545 = ~n22542 & n22544;
  assign n22546 = ~n22542 & ~n22544;
  assign n22547 = n22542 & n22544;
  assign n22548 = ~n22546 & ~n22547;
  assign n22549 = n6835 & n21252;
  assign n22550 = n7460 & n21249;
  assign n22551 = n6836 & n21635;
  assign n22552 = n7487 & n21246;
  assign n22553 = ~n22551 & ~n22552;
  assign n22554 = ~n22550 & n22553;
  assign n22555 = ~n22549 & n22554;
  assign n22556 = pi14  & n22555;
  assign n22557 = ~pi14  & ~n22555;
  assign n22558 = ~n22556 & ~n22557;
  assign n22559 = n22166 & n22176;
  assign n22560 = ~n22177 & ~n22559;
  assign n22561 = ~n22558 & n22560;
  assign n22562 = n6835 & n21255;
  assign n22563 = n7460 & n21252;
  assign n22564 = n6836 & n21506;
  assign n22565 = n7487 & n21249;
  assign n22566 = ~n22564 & ~n22565;
  assign n22567 = ~n22563 & n22566;
  assign n22568 = ~n22562 & n22567;
  assign n22569 = ~pi14  & ~n22568;
  assign n22570 = pi14  & n22568;
  assign n22571 = ~n22569 & ~n22570;
  assign n22572 = pi17  & ~n22154;
  assign n22573 = n22161 & ~n22572;
  assign n22574 = ~n22161 & n22572;
  assign n22575 = ~n22573 & ~n22574;
  assign n22576 = ~n22571 & n22575;
  assign n22577 = ~n22571 & ~n22575;
  assign n22578 = n22571 & n22575;
  assign n22579 = ~n22577 & ~n22578;
  assign n22580 = n6835 & n21258;
  assign n22581 = n7460 & n21255;
  assign n22582 = n6836 & n21546;
  assign n22583 = n7487 & n21252;
  assign n22584 = ~n22582 & ~n22583;
  assign n22585 = ~n22581 & n22584;
  assign n22586 = ~n22580 & n22585;
  assign n22587 = pi14  & n22586;
  assign n22588 = ~pi14  & ~n22586;
  assign n22589 = ~n22587 & ~n22588;
  assign n22590 = pi17  & n22152;
  assign n22591 = ~n22151 & n22590;
  assign n22592 = n22151 & ~n22590;
  assign n22593 = ~n22591 & ~n22592;
  assign n22594 = ~n22589 & n22593;
  assign n22595 = n6836 & ~n21519;
  assign n22596 = n7487 & n21263;
  assign n22597 = n7460 & n21265;
  assign n22598 = ~n22596 & ~n22597;
  assign n22599 = ~n22595 & n22598;
  assign n22600 = ~n6833 & n21265;
  assign n22601 = pi14  & ~n22600;
  assign n22602 = n22599 & n22601;
  assign n22603 = n6835 & n21265;
  assign n22604 = n7460 & n21263;
  assign n22605 = n6836 & ~n21531;
  assign n22606 = n7487 & n21258;
  assign n22607 = ~n22605 & ~n22606;
  assign n22608 = ~n22604 & n22607;
  assign n22609 = ~n22603 & n22608;
  assign n22610 = n22602 & n22609;
  assign n22611 = n22152 & n22610;
  assign n22612 = ~n22152 & n22610;
  assign n22613 = n22152 & ~n22610;
  assign n22614 = ~n22612 & ~n22613;
  assign n22615 = n6835 & n21263;
  assign n22616 = n7460 & n21258;
  assign n22617 = n6836 & n21583;
  assign n22618 = n7487 & n21255;
  assign n22619 = ~n22617 & ~n22618;
  assign n22620 = ~n22616 & n22619;
  assign n22621 = ~n22615 & n22620;
  assign n22622 = pi14  & n22621;
  assign n22623 = ~pi14  & ~n22621;
  assign n22624 = ~n22622 & ~n22623;
  assign n22625 = ~n22614 & ~n22624;
  assign n22626 = ~n22611 & ~n22625;
  assign n22627 = n22589 & ~n22593;
  assign n22628 = ~n22594 & ~n22627;
  assign n22629 = ~n22626 & n22628;
  assign n22630 = ~n22594 & ~n22629;
  assign n22631 = ~n22579 & ~n22630;
  assign n22632 = ~n22576 & ~n22631;
  assign n22633 = n22558 & ~n22560;
  assign n22634 = ~n22561 & ~n22633;
  assign n22635 = ~n22632 & n22634;
  assign n22636 = ~n22561 & ~n22635;
  assign n22637 = ~n22548 & ~n22636;
  assign n22638 = ~n22545 & ~n22637;
  assign n22639 = n22521 & n22531;
  assign n22640 = ~n22521 & ~n22531;
  assign n22641 = ~n22639 & ~n22640;
  assign n22642 = ~n22638 & ~n22641;
  assign n22643 = ~n22532 & ~n22642;
  assign n22644 = n22508 & n22518;
  assign n22645 = ~n22508 & ~n22518;
  assign n22646 = ~n22644 & ~n22645;
  assign n22647 = ~n22643 & ~n22646;
  assign n22648 = ~n22519 & ~n22647;
  assign n22649 = ~n22495 & n22505;
  assign n22650 = ~n22506 & ~n22649;
  assign n22651 = ~n22648 & n22650;
  assign n22652 = ~n22506 & ~n22651;
  assign n22653 = n22489 & n22492;
  assign n22654 = ~n22493 & ~n22653;
  assign n22655 = ~n22652 & n22654;
  assign n22656 = ~n22493 & ~n22655;
  assign n22657 = ~n22479 & ~n22656;
  assign n22658 = ~n22476 & ~n22657;
  assign n22659 = ~n22463 & ~n22658;
  assign n22660 = ~n22460 & ~n22659;
  assign n22661 = n22436 & n22446;
  assign n22662 = ~n22436 & ~n22446;
  assign n22663 = ~n22661 & ~n22662;
  assign n22664 = ~n22660 & ~n22663;
  assign n22665 = ~n22447 & ~n22664;
  assign n22666 = n22423 & n22433;
  assign n22667 = ~n22423 & ~n22433;
  assign n22668 = ~n22666 & ~n22667;
  assign n22669 = ~n22665 & ~n22668;
  assign n22670 = ~n22434 & ~n22669;
  assign n22671 = ~n22410 & n22420;
  assign n22672 = ~n22421 & ~n22671;
  assign n22673 = ~n22670 & n22672;
  assign n22674 = ~n22421 & ~n22673;
  assign n22675 = ~n22408 & ~n22674;
  assign n22676 = ~n22405 & ~n22675;
  assign n22677 = ~n22390 & ~n22676;
  assign n22678 = ~n22387 & ~n22677;
  assign n22679 = n22359 & n22371;
  assign n22680 = ~n22359 & ~n22371;
  assign n22681 = ~n22679 & ~n22680;
  assign n22682 = ~n22678 & ~n22681;
  assign n22683 = ~n22372 & ~n22682;
  assign n22684 = ~n22354 & ~n22357;
  assign n22685 = n6184 & n21219;
  assign n22686 = n6527 & n21216;
  assign n22687 = n6185 & n22394;
  assign n22688 = n6543 & n21213;
  assign n22689 = ~n22687 & ~n22688;
  assign n22690 = ~n22686 & n22689;
  assign n22691 = ~n22685 & n22690;
  assign n22692 = ~pi17  & ~n22691;
  assign n22693 = pi17  & n22691;
  assign n22694 = ~n22692 & ~n22693;
  assign n22695 = n22337 & ~n22347;
  assign n22696 = ~n22235 & ~n22350;
  assign n22697 = ~n22695 & ~n22696;
  assign n22698 = n5238 & n21237;
  assign n22699 = n71 & n21234;
  assign n22700 = n5239 & n21789;
  assign n22701 = n5326 & n21231;
  assign n22702 = ~n22700 & ~n22701;
  assign n22703 = ~n22699 & n22702;
  assign n22704 = ~n22698 & n22703;
  assign n22705 = ~pi23  & ~n22704;
  assign n22706 = pi23  & n22704;
  assign n22707 = ~n22705 & ~n22706;
  assign n22708 = ~n22257 & n22324;
  assign n22709 = ~n22328 & ~n22708;
  assign n22710 = ~n22319 & ~n22322;
  assign n22711 = n4006 & n21255;
  assign n22712 = n4133 & n21252;
  assign n22713 = n4002 & n21506;
  assign n22714 = n4555 & n21249;
  assign n22715 = ~n22713 & ~n22714;
  assign n22716 = ~n22712 & n22715;
  assign n22717 = ~n22711 & n22716;
  assign n22718 = ~pi29  & ~n22717;
  assign n22719 = pi29  & n22717;
  assign n22720 = ~n22718 & ~n22719;
  assign n22721 = ~n22310 & ~n22315;
  assign n22722 = n5849 & n7148;
  assign n22723 = n1708 & n22722;
  assign n22724 = ~n166 & n22723;
  assign n22725 = ~n310 & ~n439;
  assign n22726 = ~n383 & n22725;
  assign n22727 = n759 & n22726;
  assign n22728 = n1409 & n22727;
  assign n22729 = n1934 & n22728;
  assign n22730 = ~n601 & n22729;
  assign n22731 = ~n242 & n22730;
  assign n22732 = n22724 & n22731;
  assign n22733 = n189 & n4277;
  assign n22734 = n13073 & n22733;
  assign n22735 = n15136 & n22734;
  assign n22736 = ~n413 & n22735;
  assign n22737 = n1876 & n4672;
  assign n22738 = ~n320 & n22737;
  assign n22739 = ~n132 & n22738;
  assign n22740 = n22736 & n22739;
  assign n22741 = n22732 & n22740;
  assign n22742 = n22721 & ~n22741;
  assign n22743 = ~n22721 & n22741;
  assign n22744 = ~n22742 & ~n22743;
  assign n22745 = n3641 & n21265;
  assign n22746 = n3740 & n21263;
  assign n22747 = n556 & ~n21531;
  assign n22748 = n3961 & n21258;
  assign n22749 = ~n22747 & ~n22748;
  assign n22750 = ~n22746 & n22749;
  assign n22751 = ~n22745 & n22750;
  assign n22752 = n22744 & ~n22751;
  assign n22753 = ~n22744 & n22751;
  assign n22754 = ~n22752 & ~n22753;
  assign n22755 = ~n22720 & n22754;
  assign n22756 = n22720 & ~n22754;
  assign n22757 = ~n22755 & ~n22756;
  assign n22758 = n22710 & ~n22757;
  assign n22759 = ~n22710 & n22757;
  assign n22760 = ~n22758 & ~n22759;
  assign n22761 = n4601 & n21246;
  assign n22762 = n4783 & n21243;
  assign n22763 = n4602 & n21604;
  assign n22764 = n4801 & n21240;
  assign n22765 = ~n22763 & ~n22764;
  assign n22766 = ~n22762 & n22765;
  assign n22767 = ~n22761 & n22766;
  assign n22768 = pi26  & n22767;
  assign n22769 = ~pi26  & ~n22767;
  assign n22770 = ~n22768 & ~n22769;
  assign n22771 = n22760 & n22770;
  assign n22772 = ~n22760 & ~n22770;
  assign n22773 = ~n22771 & ~n22772;
  assign n22774 = ~n22709 & ~n22773;
  assign n22775 = n22709 & n22773;
  assign n22776 = ~n22774 & ~n22775;
  assign n22777 = ~n22707 & ~n22776;
  assign n22778 = n22707 & n22776;
  assign n22779 = ~n22777 & ~n22778;
  assign n22780 = ~n22245 & n22330;
  assign n22781 = ~n22336 & ~n22780;
  assign n22782 = n22779 & n22781;
  assign n22783 = ~n22779 & ~n22781;
  assign n22784 = ~n22782 & ~n22783;
  assign n22785 = n5435 & n21228;
  assign n22786 = n6055 & n21225;
  assign n22787 = n5429 & n21988;
  assign n22788 = n6071 & n21222;
  assign n22789 = ~n22787 & ~n22788;
  assign n22790 = ~n22786 & n22789;
  assign n22791 = ~n22785 & n22790;
  assign n22792 = pi20  & n22791;
  assign n22793 = ~pi20  & ~n22791;
  assign n22794 = ~n22792 & ~n22793;
  assign n22795 = n22784 & n22794;
  assign n22796 = ~n22784 & ~n22794;
  assign n22797 = ~n22795 & ~n22796;
  assign n22798 = ~n22697 & n22797;
  assign n22799 = n22697 & ~n22797;
  assign n22800 = ~n22798 & ~n22799;
  assign n22801 = ~n22694 & ~n22800;
  assign n22802 = n22694 & n22800;
  assign n22803 = ~n22801 & ~n22802;
  assign n22804 = n22684 & ~n22803;
  assign n22805 = ~n22684 & n22803;
  assign n22806 = ~n22804 & ~n22805;
  assign n22807 = n6835 & n21210;
  assign n22808 = n7460 & n21207;
  assign n22809 = n21333 & ~n21335;
  assign n22810 = ~n21336 & ~n22809;
  assign n22811 = n6836 & n22810;
  assign n22812 = n7487 & n21204;
  assign n22813 = ~n22811 & ~n22812;
  assign n22814 = ~n22808 & n22813;
  assign n22815 = ~n22807 & n22814;
  assign n22816 = pi14  & n22815;
  assign n22817 = ~pi14  & ~n22815;
  assign n22818 = ~n22816 & ~n22817;
  assign n22819 = n22806 & n22818;
  assign n22820 = ~n22806 & ~n22818;
  assign n22821 = ~n22819 & ~n22820;
  assign n22822 = ~n22683 & ~n22821;
  assign n22823 = n22683 & n22821;
  assign n22824 = ~n22822 & ~n22823;
  assign n22825 = ~n21490 & n22824;
  assign n22826 = ~n21490 & ~n22824;
  assign n22827 = n21490 & n22824;
  assign n22828 = ~n22826 & ~n22827;
  assign n22829 = n7654 & n21204;
  assign n22830 = n8091 & n21201;
  assign n22831 = n21341 & ~n21343;
  assign n22832 = ~n21344 & ~n22831;
  assign n22833 = n7648 & n22832;
  assign n22834 = n8120 & n21198;
  assign n22835 = ~n22833 & ~n22834;
  assign n22836 = ~n22830 & n22835;
  assign n22837 = ~n22829 & n22836;
  assign n22838 = ~pi11  & ~n22837;
  assign n22839 = pi11  & n22837;
  assign n22840 = ~n22838 & ~n22839;
  assign n22841 = n22678 & n22681;
  assign n22842 = ~n22682 & ~n22841;
  assign n22843 = ~n22840 & n22842;
  assign n22844 = ~n22840 & ~n22842;
  assign n22845 = n22840 & n22842;
  assign n22846 = ~n22844 & ~n22845;
  assign n22847 = n22390 & n22676;
  assign n22848 = ~n22677 & ~n22847;
  assign n22849 = n7654 & n21207;
  assign n22850 = n8091 & n21204;
  assign n22851 = n21337 & ~n21339;
  assign n22852 = ~n21340 & ~n22851;
  assign n22853 = n7648 & n22852;
  assign n22854 = n8120 & n21201;
  assign n22855 = ~n22853 & ~n22854;
  assign n22856 = ~n22850 & n22855;
  assign n22857 = ~n22849 & n22856;
  assign n22858 = pi11  & n22857;
  assign n22859 = ~pi11  & ~n22857;
  assign n22860 = ~n22858 & ~n22859;
  assign n22861 = n22848 & ~n22860;
  assign n22862 = n22408 & n22674;
  assign n22863 = ~n22675 & ~n22862;
  assign n22864 = n7654 & n21210;
  assign n22865 = n8091 & n21207;
  assign n22866 = n7648 & n22810;
  assign n22867 = n8120 & n21204;
  assign n22868 = ~n22866 & ~n22867;
  assign n22869 = ~n22865 & n22868;
  assign n22870 = ~n22864 & n22869;
  assign n22871 = pi11  & n22870;
  assign n22872 = ~pi11  & ~n22870;
  assign n22873 = ~n22871 & ~n22872;
  assign n22874 = n22863 & ~n22873;
  assign n22875 = n7654 & n21213;
  assign n22876 = n8091 & n21210;
  assign n22877 = n7648 & n22363;
  assign n22878 = n8120 & n21207;
  assign n22879 = ~n22877 & ~n22878;
  assign n22880 = ~n22876 & n22879;
  assign n22881 = ~n22875 & n22880;
  assign n22882 = ~pi11  & ~n22881;
  assign n22883 = pi11  & n22881;
  assign n22884 = ~n22882 & ~n22883;
  assign n22885 = n22670 & ~n22672;
  assign n22886 = ~n22673 & ~n22885;
  assign n22887 = ~n22884 & n22886;
  assign n22888 = ~n22884 & ~n22886;
  assign n22889 = n22884 & n22886;
  assign n22890 = ~n22888 & ~n22889;
  assign n22891 = n7654 & n21216;
  assign n22892 = n8091 & n21213;
  assign n22893 = n7648 & n22376;
  assign n22894 = n8120 & n21210;
  assign n22895 = ~n22893 & ~n22894;
  assign n22896 = ~n22892 & n22895;
  assign n22897 = ~n22891 & n22896;
  assign n22898 = ~pi11  & ~n22897;
  assign n22899 = pi11  & n22897;
  assign n22900 = ~n22898 & ~n22899;
  assign n22901 = ~n22665 & n22668;
  assign n22902 = n22665 & ~n22668;
  assign n22903 = ~n22901 & ~n22902;
  assign n22904 = ~n22900 & ~n22903;
  assign n22905 = n7654 & n21219;
  assign n22906 = n8091 & n21216;
  assign n22907 = n7648 & n22394;
  assign n22908 = n8120 & n21213;
  assign n22909 = ~n22907 & ~n22908;
  assign n22910 = ~n22906 & n22909;
  assign n22911 = ~n22905 & n22910;
  assign n22912 = ~pi11  & ~n22911;
  assign n22913 = pi11  & n22911;
  assign n22914 = ~n22912 & ~n22913;
  assign n22915 = n22660 & n22663;
  assign n22916 = ~n22664 & ~n22915;
  assign n22917 = ~n22914 & n22916;
  assign n22918 = ~n22914 & ~n22916;
  assign n22919 = n22914 & n22916;
  assign n22920 = ~n22918 & ~n22919;
  assign n22921 = n22463 & n22658;
  assign n22922 = ~n22659 & ~n22921;
  assign n22923 = n7654 & n21222;
  assign n22924 = n8091 & n21219;
  assign n22925 = n7648 & n22225;
  assign n22926 = n8120 & n21216;
  assign n22927 = ~n22925 & ~n22926;
  assign n22928 = ~n22924 & n22927;
  assign n22929 = ~n22923 & n22928;
  assign n22930 = pi11  & n22929;
  assign n22931 = ~pi11  & ~n22929;
  assign n22932 = ~n22930 & ~n22931;
  assign n22933 = n22922 & ~n22932;
  assign n22934 = n22479 & n22656;
  assign n22935 = ~n22657 & ~n22934;
  assign n22936 = n7654 & n21225;
  assign n22937 = n8091 & n21222;
  assign n22938 = n7648 & n21973;
  assign n22939 = n8120 & n21219;
  assign n22940 = ~n22938 & ~n22939;
  assign n22941 = ~n22937 & n22940;
  assign n22942 = ~n22936 & n22941;
  assign n22943 = pi11  & n22942;
  assign n22944 = ~pi11  & ~n22942;
  assign n22945 = ~n22943 & ~n22944;
  assign n22946 = n22935 & ~n22945;
  assign n22947 = n22652 & ~n22654;
  assign n22948 = ~n22655 & ~n22947;
  assign n22949 = n7654 & n21228;
  assign n22950 = n8091 & n21225;
  assign n22951 = n7648 & n21988;
  assign n22952 = n8120 & n21222;
  assign n22953 = ~n22951 & ~n22952;
  assign n22954 = ~n22950 & n22953;
  assign n22955 = ~n22949 & n22954;
  assign n22956 = pi11  & n22955;
  assign n22957 = ~pi11  & ~n22955;
  assign n22958 = ~n22956 & ~n22957;
  assign n22959 = n22948 & ~n22958;
  assign n22960 = n7654 & n21231;
  assign n22961 = n8091 & n21228;
  assign n22962 = n7648 & n22001;
  assign n22963 = n8120 & n21225;
  assign n22964 = ~n22962 & ~n22963;
  assign n22965 = ~n22961 & n22964;
  assign n22966 = ~n22960 & n22965;
  assign n22967 = ~pi11  & ~n22966;
  assign n22968 = pi11  & n22966;
  assign n22969 = ~n22967 & ~n22968;
  assign n22970 = n22648 & ~n22650;
  assign n22971 = ~n22651 & ~n22970;
  assign n22972 = ~n22969 & n22971;
  assign n22973 = ~n22969 & ~n22971;
  assign n22974 = n22969 & n22971;
  assign n22975 = ~n22973 & ~n22974;
  assign n22976 = n7654 & n21234;
  assign n22977 = n8091 & n21231;
  assign n22978 = n7648 & n21494;
  assign n22979 = n8120 & n21228;
  assign n22980 = ~n22978 & ~n22979;
  assign n22981 = ~n22977 & n22980;
  assign n22982 = ~n22976 & n22981;
  assign n22983 = ~pi11  & ~n22982;
  assign n22984 = pi11  & n22982;
  assign n22985 = ~n22983 & ~n22984;
  assign n22986 = n22643 & n22646;
  assign n22987 = ~n22647 & ~n22986;
  assign n22988 = ~n22985 & n22987;
  assign n22989 = ~n22985 & ~n22987;
  assign n22990 = n22985 & n22987;
  assign n22991 = ~n22989 & ~n22990;
  assign n22992 = n7654 & n21237;
  assign n22993 = n8091 & n21234;
  assign n22994 = n7648 & n21789;
  assign n22995 = n8120 & n21231;
  assign n22996 = ~n22994 & ~n22995;
  assign n22997 = ~n22993 & n22996;
  assign n22998 = ~n22992 & n22997;
  assign n22999 = ~pi11  & ~n22998;
  assign n23000 = pi11  & n22998;
  assign n23001 = ~n22999 & ~n23000;
  assign n23002 = ~n22638 & n22641;
  assign n23003 = n22638 & ~n22641;
  assign n23004 = ~n23002 & ~n23003;
  assign n23005 = ~n23001 & ~n23004;
  assign n23006 = n22548 & n22636;
  assign n23007 = ~n22637 & ~n23006;
  assign n23008 = n7654 & n21240;
  assign n23009 = n8091 & n21237;
  assign n23010 = n7648 & n21807;
  assign n23011 = n8120 & n21234;
  assign n23012 = ~n23010 & ~n23011;
  assign n23013 = ~n23009 & n23012;
  assign n23014 = ~n23008 & n23013;
  assign n23015 = pi11  & n23014;
  assign n23016 = ~pi11  & ~n23014;
  assign n23017 = ~n23015 & ~n23016;
  assign n23018 = n23007 & ~n23017;
  assign n23019 = n22632 & ~n22634;
  assign n23020 = ~n22635 & ~n23019;
  assign n23021 = n7654 & n21243;
  assign n23022 = n8091 & n21240;
  assign n23023 = n7648 & n21768;
  assign n23024 = n8120 & n21237;
  assign n23025 = ~n23023 & ~n23024;
  assign n23026 = ~n23022 & n23025;
  assign n23027 = ~n23021 & n23026;
  assign n23028 = pi11  & n23027;
  assign n23029 = ~pi11  & ~n23027;
  assign n23030 = ~n23028 & ~n23029;
  assign n23031 = n23020 & ~n23030;
  assign n23032 = n22579 & n22630;
  assign n23033 = ~n22631 & ~n23032;
  assign n23034 = n7654 & n21246;
  assign n23035 = n8091 & n21243;
  assign n23036 = n7648 & n21604;
  assign n23037 = n8120 & n21240;
  assign n23038 = ~n23036 & ~n23037;
  assign n23039 = ~n23035 & n23038;
  assign n23040 = ~n23034 & n23039;
  assign n23041 = pi11  & n23040;
  assign n23042 = ~pi11  & ~n23040;
  assign n23043 = ~n23041 & ~n23042;
  assign n23044 = n23033 & ~n23043;
  assign n23045 = n7654 & n21249;
  assign n23046 = n8091 & n21246;
  assign n23047 = n7648 & n21617;
  assign n23048 = n8120 & n21243;
  assign n23049 = ~n23047 & ~n23048;
  assign n23050 = ~n23046 & n23049;
  assign n23051 = ~n23045 & n23050;
  assign n23052 = ~pi11  & ~n23051;
  assign n23053 = pi11  & n23051;
  assign n23054 = ~n23052 & ~n23053;
  assign n23055 = n22626 & ~n22628;
  assign n23056 = ~n22629 & ~n23055;
  assign n23057 = ~n23054 & n23056;
  assign n23058 = ~n23054 & ~n23056;
  assign n23059 = n23054 & n23056;
  assign n23060 = ~n23058 & ~n23059;
  assign n23061 = n7654 & n21252;
  assign n23062 = n8091 & n21249;
  assign n23063 = n7648 & n21635;
  assign n23064 = n8120 & n21246;
  assign n23065 = ~n23063 & ~n23064;
  assign n23066 = ~n23062 & n23065;
  assign n23067 = ~n23061 & n23066;
  assign n23068 = pi11  & n23067;
  assign n23069 = ~pi11  & ~n23067;
  assign n23070 = ~n23068 & ~n23069;
  assign n23071 = n22614 & n22624;
  assign n23072 = ~n22625 & ~n23071;
  assign n23073 = ~n23070 & n23072;
  assign n23074 = n7654 & n21255;
  assign n23075 = n8091 & n21252;
  assign n23076 = n7648 & n21506;
  assign n23077 = n8120 & n21249;
  assign n23078 = ~n23076 & ~n23077;
  assign n23079 = ~n23075 & n23078;
  assign n23080 = ~n23074 & n23079;
  assign n23081 = ~pi11  & ~n23080;
  assign n23082 = pi11  & n23080;
  assign n23083 = ~n23081 & ~n23082;
  assign n23084 = pi14  & ~n22602;
  assign n23085 = n22609 & ~n23084;
  assign n23086 = ~n22609 & n23084;
  assign n23087 = ~n23085 & ~n23086;
  assign n23088 = ~n23083 & n23087;
  assign n23089 = ~n23083 & ~n23087;
  assign n23090 = n23083 & n23087;
  assign n23091 = ~n23089 & ~n23090;
  assign n23092 = n7654 & n21258;
  assign n23093 = n8091 & n21255;
  assign n23094 = n7648 & n21546;
  assign n23095 = n8120 & n21252;
  assign n23096 = ~n23094 & ~n23095;
  assign n23097 = ~n23093 & n23096;
  assign n23098 = ~n23092 & n23097;
  assign n23099 = pi11  & n23098;
  assign n23100 = ~pi11  & ~n23098;
  assign n23101 = ~n23099 & ~n23100;
  assign n23102 = pi14  & n22600;
  assign n23103 = ~n22599 & n23102;
  assign n23104 = n22599 & ~n23102;
  assign n23105 = ~n23103 & ~n23104;
  assign n23106 = ~n23101 & n23105;
  assign n23107 = n7648 & ~n21519;
  assign n23108 = n8120 & n21263;
  assign n23109 = n8091 & n21265;
  assign n23110 = ~n23108 & ~n23109;
  assign n23111 = ~n23107 & n23110;
  assign n23112 = ~n7644 & n21265;
  assign n23113 = pi11  & ~n23112;
  assign n23114 = n23111 & n23113;
  assign n23115 = n7654 & n21265;
  assign n23116 = n8091 & n21263;
  assign n23117 = n7648 & ~n21531;
  assign n23118 = n8120 & n21258;
  assign n23119 = ~n23117 & ~n23118;
  assign n23120 = ~n23116 & n23119;
  assign n23121 = ~n23115 & n23120;
  assign n23122 = n23114 & n23121;
  assign n23123 = n22600 & n23122;
  assign n23124 = ~n22600 & n23122;
  assign n23125 = n22600 & ~n23122;
  assign n23126 = ~n23124 & ~n23125;
  assign n23127 = n7654 & n21263;
  assign n23128 = n8091 & n21258;
  assign n23129 = n7648 & n21583;
  assign n23130 = n8120 & n21255;
  assign n23131 = ~n23129 & ~n23130;
  assign n23132 = ~n23128 & n23131;
  assign n23133 = ~n23127 & n23132;
  assign n23134 = pi11  & n23133;
  assign n23135 = ~pi11  & ~n23133;
  assign n23136 = ~n23134 & ~n23135;
  assign n23137 = ~n23126 & ~n23136;
  assign n23138 = ~n23123 & ~n23137;
  assign n23139 = n23101 & ~n23105;
  assign n23140 = ~n23106 & ~n23139;
  assign n23141 = ~n23138 & n23140;
  assign n23142 = ~n23106 & ~n23141;
  assign n23143 = ~n23091 & ~n23142;
  assign n23144 = ~n23088 & ~n23143;
  assign n23145 = n23070 & ~n23072;
  assign n23146 = ~n23073 & ~n23145;
  assign n23147 = ~n23144 & n23146;
  assign n23148 = ~n23073 & ~n23147;
  assign n23149 = ~n23060 & ~n23148;
  assign n23150 = ~n23057 & ~n23149;
  assign n23151 = n23033 & n23043;
  assign n23152 = ~n23033 & ~n23043;
  assign n23153 = ~n23151 & ~n23152;
  assign n23154 = ~n23150 & ~n23153;
  assign n23155 = ~n23044 & ~n23154;
  assign n23156 = n23020 & n23030;
  assign n23157 = ~n23020 & ~n23030;
  assign n23158 = ~n23156 & ~n23157;
  assign n23159 = ~n23155 & ~n23158;
  assign n23160 = ~n23031 & ~n23159;
  assign n23161 = ~n23007 & n23017;
  assign n23162 = ~n23018 & ~n23161;
  assign n23163 = ~n23160 & n23162;
  assign n23164 = ~n23018 & ~n23163;
  assign n23165 = n23001 & n23004;
  assign n23166 = ~n23005 & ~n23165;
  assign n23167 = ~n23164 & n23166;
  assign n23168 = ~n23005 & ~n23167;
  assign n23169 = ~n22991 & ~n23168;
  assign n23170 = ~n22988 & ~n23169;
  assign n23171 = ~n22975 & ~n23170;
  assign n23172 = ~n22972 & ~n23171;
  assign n23173 = n22948 & n22958;
  assign n23174 = ~n22948 & ~n22958;
  assign n23175 = ~n23173 & ~n23174;
  assign n23176 = ~n23172 & ~n23175;
  assign n23177 = ~n22959 & ~n23176;
  assign n23178 = n22935 & n22945;
  assign n23179 = ~n22935 & ~n22945;
  assign n23180 = ~n23178 & ~n23179;
  assign n23181 = ~n23177 & ~n23180;
  assign n23182 = ~n22946 & ~n23181;
  assign n23183 = ~n22922 & n22932;
  assign n23184 = ~n22933 & ~n23183;
  assign n23185 = ~n23182 & n23184;
  assign n23186 = ~n22933 & ~n23185;
  assign n23187 = ~n22920 & ~n23186;
  assign n23188 = ~n22917 & ~n23187;
  assign n23189 = n22900 & n22903;
  assign n23190 = ~n22904 & ~n23189;
  assign n23191 = ~n23188 & n23190;
  assign n23192 = ~n22904 & ~n23191;
  assign n23193 = ~n22890 & ~n23192;
  assign n23194 = ~n22887 & ~n23193;
  assign n23195 = n22863 & n22873;
  assign n23196 = ~n22863 & ~n22873;
  assign n23197 = ~n23195 & ~n23196;
  assign n23198 = ~n23194 & ~n23197;
  assign n23199 = ~n22874 & ~n23198;
  assign n23200 = ~n22848 & n22860;
  assign n23201 = ~n22861 & ~n23200;
  assign n23202 = ~n23199 & n23201;
  assign n23203 = ~n22861 & ~n23202;
  assign n23204 = ~n22846 & ~n23203;
  assign n23205 = ~n22843 & ~n23204;
  assign n23206 = ~n22828 & ~n23205;
  assign n23207 = ~n22825 & ~n23206;
  assign n23208 = n7654 & n21198;
  assign n23209 = n8091 & n21195;
  assign n23210 = n21349 & ~n21351;
  assign n23211 = ~n21352 & ~n23210;
  assign n23212 = n7648 & n23211;
  assign n23213 = n8120 & n21192;
  assign n23214 = ~n23212 & ~n23213;
  assign n23215 = ~n23209 & n23214;
  assign n23216 = ~n23208 & n23215;
  assign n23217 = ~pi11  & ~n23216;
  assign n23218 = pi11  & n23216;
  assign n23219 = ~n23217 & ~n23218;
  assign n23220 = n22806 & ~n22818;
  assign n23221 = ~n22822 & ~n23220;
  assign n23222 = n6184 & n21216;
  assign n23223 = n6527 & n21213;
  assign n23224 = n6185 & n22376;
  assign n23225 = n6543 & n21210;
  assign n23226 = ~n23224 & ~n23225;
  assign n23227 = ~n23223 & n23226;
  assign n23228 = ~n23222 & n23227;
  assign n23229 = ~pi17  & ~n23228;
  assign n23230 = pi17  & n23228;
  assign n23231 = ~n23229 & ~n23230;
  assign n23232 = n22784 & ~n22794;
  assign n23233 = ~n22697 & ~n22797;
  assign n23234 = ~n23232 & ~n23233;
  assign n23235 = ~n22707 & n22776;
  assign n23236 = ~n22783 & ~n23235;
  assign n23237 = n5238 & n21234;
  assign n23238 = n71 & n21231;
  assign n23239 = n5239 & n21494;
  assign n23240 = n5326 & n21228;
  assign n23241 = ~n23239 & ~n23240;
  assign n23242 = ~n23238 & n23241;
  assign n23243 = ~n23237 & n23242;
  assign n23244 = ~pi23  & ~n23243;
  assign n23245 = pi23  & n23243;
  assign n23246 = ~n23244 & ~n23245;
  assign n23247 = n22760 & ~n22770;
  assign n23248 = ~n22774 & ~n23247;
  assign n23249 = n4006 & n21252;
  assign n23250 = n4133 & n21249;
  assign n23251 = n4002 & n21635;
  assign n23252 = n4555 & n21246;
  assign n23253 = ~n23251 & ~n23252;
  assign n23254 = ~n23250 & n23253;
  assign n23255 = ~n23249 & n23254;
  assign n23256 = ~pi29  & ~n23255;
  assign n23257 = pi29  & n23255;
  assign n23258 = ~n23256 & ~n23257;
  assign n23259 = n2444 & n4653;
  assign n23260 = ~n131 & n23259;
  assign n23261 = ~n309 & n901;
  assign n23262 = ~n593 & n23261;
  assign n23263 = n3695 & n23262;
  assign n23264 = n5704 & n23263;
  assign n23265 = n467 & n23264;
  assign n23266 = ~n442 & n23265;
  assign n23267 = n23260 & n23266;
  assign n23268 = n1805 & n5959;
  assign n23269 = n974 & n23268;
  assign n23270 = n386 & n23269;
  assign n23271 = ~n277 & n23270;
  assign n23272 = n515 & n2681;
  assign n23273 = n787 & n23272;
  assign n23274 = ~n533 & n23273;
  assign n23275 = n23271 & n23274;
  assign n23276 = n23267 & n23275;
  assign n23277 = n3641 & n21263;
  assign n23278 = n556 & n21583;
  assign n23279 = n3961 & n21255;
  assign n23280 = n3740 & n21258;
  assign n23281 = ~n23279 & ~n23280;
  assign n23282 = ~n23278 & n23281;
  assign n23283 = ~n23277 & n23282;
  assign n23284 = ~n23276 & n23283;
  assign n23285 = n23276 & ~n23283;
  assign n23286 = ~n23284 & ~n23285;
  assign n23287 = ~n22742 & n22751;
  assign n23288 = ~n22743 & ~n23287;
  assign n23289 = ~n23286 & n23288;
  assign n23290 = n23286 & ~n23288;
  assign n23291 = ~n23289 & ~n23290;
  assign n23292 = ~n23258 & ~n23291;
  assign n23293 = n23258 & n23291;
  assign n23294 = ~n23292 & ~n23293;
  assign n23295 = ~n22755 & ~n22759;
  assign n23296 = n23294 & n23295;
  assign n23297 = ~n23294 & ~n23295;
  assign n23298 = ~n23296 & ~n23297;
  assign n23299 = n4601 & n21243;
  assign n23300 = n4783 & n21240;
  assign n23301 = n4602 & n21768;
  assign n23302 = n4801 & n21237;
  assign n23303 = ~n23301 & ~n23302;
  assign n23304 = ~n23300 & n23303;
  assign n23305 = ~n23299 & n23304;
  assign n23306 = pi26  & n23305;
  assign n23307 = ~pi26  & ~n23305;
  assign n23308 = ~n23306 & ~n23307;
  assign n23309 = n23298 & n23308;
  assign n23310 = ~n23298 & ~n23308;
  assign n23311 = ~n23309 & ~n23310;
  assign n23312 = ~n23248 & n23311;
  assign n23313 = n23248 & ~n23311;
  assign n23314 = ~n23312 & ~n23313;
  assign n23315 = ~n23246 & ~n23314;
  assign n23316 = n23246 & n23314;
  assign n23317 = ~n23315 & ~n23316;
  assign n23318 = n23236 & ~n23317;
  assign n23319 = ~n23236 & n23317;
  assign n23320 = ~n23318 & ~n23319;
  assign n23321 = n5435 & n21225;
  assign n23322 = n6055 & n21222;
  assign n23323 = n5429 & n21973;
  assign n23324 = n6071 & n21219;
  assign n23325 = ~n23323 & ~n23324;
  assign n23326 = ~n23322 & n23325;
  assign n23327 = ~n23321 & n23326;
  assign n23328 = pi20  & n23327;
  assign n23329 = ~pi20  & ~n23327;
  assign n23330 = ~n23328 & ~n23329;
  assign n23331 = n23320 & n23330;
  assign n23332 = ~n23320 & ~n23330;
  assign n23333 = ~n23331 & ~n23332;
  assign n23334 = ~n23234 & ~n23333;
  assign n23335 = n23234 & n23333;
  assign n23336 = ~n23334 & ~n23335;
  assign n23337 = ~n23231 & ~n23336;
  assign n23338 = n23231 & n23336;
  assign n23339 = ~n23337 & ~n23338;
  assign n23340 = ~n22801 & ~n22805;
  assign n23341 = n23339 & n23340;
  assign n23342 = ~n23339 & ~n23340;
  assign n23343 = ~n23341 & ~n23342;
  assign n23344 = n6835 & n21207;
  assign n23345 = n7460 & n21204;
  assign n23346 = n6836 & n22852;
  assign n23347 = n7487 & n21201;
  assign n23348 = ~n23346 & ~n23347;
  assign n23349 = ~n23345 & n23348;
  assign n23350 = ~n23344 & n23349;
  assign n23351 = pi14  & n23350;
  assign n23352 = ~pi14  & ~n23350;
  assign n23353 = ~n23351 & ~n23352;
  assign n23354 = n23343 & n23353;
  assign n23355 = ~n23343 & ~n23353;
  assign n23356 = ~n23354 & ~n23355;
  assign n23357 = ~n23221 & n23356;
  assign n23358 = n23221 & ~n23356;
  assign n23359 = ~n23357 & ~n23358;
  assign n23360 = ~n23219 & ~n23359;
  assign n23361 = n23219 & n23359;
  assign n23362 = ~n23360 & ~n23361;
  assign n23363 = n23207 & ~n23362;
  assign n23364 = ~n23207 & n23362;
  assign n23365 = ~n23363 & ~n23364;
  assign n23366 = n8474 & n21189;
  assign n23367 = n9238 & n21186;
  assign n23368 = n21361 & ~n21363;
  assign n23369 = ~n21364 & ~n23368;
  assign n23370 = n8468 & n23369;
  assign n23371 = n9265 & n21183;
  assign n23372 = ~n23370 & ~n23371;
  assign n23373 = ~n23367 & n23372;
  assign n23374 = ~n23366 & n23373;
  assign n23375 = pi8  & n23374;
  assign n23376 = ~pi8  & ~n23374;
  assign n23377 = ~n23375 & ~n23376;
  assign n23378 = n23365 & ~n23377;
  assign n23379 = n22828 & n23205;
  assign n23380 = ~n23206 & ~n23379;
  assign n23381 = n8474 & n21192;
  assign n23382 = n9238 & n21189;
  assign n23383 = n21357 & ~n21359;
  assign n23384 = ~n21360 & ~n23383;
  assign n23385 = n8468 & n23384;
  assign n23386 = n9265 & n21186;
  assign n23387 = ~n23385 & ~n23386;
  assign n23388 = ~n23382 & n23387;
  assign n23389 = ~n23381 & n23388;
  assign n23390 = pi8  & n23389;
  assign n23391 = ~pi8  & ~n23389;
  assign n23392 = ~n23390 & ~n23391;
  assign n23393 = n23380 & ~n23392;
  assign n23394 = n22846 & n23203;
  assign n23395 = ~n23204 & ~n23394;
  assign n23396 = n8474 & n21195;
  assign n23397 = n9238 & n21192;
  assign n23398 = n21353 & ~n21355;
  assign n23399 = ~n21356 & ~n23398;
  assign n23400 = n8468 & n23399;
  assign n23401 = n9265 & n21189;
  assign n23402 = ~n23400 & ~n23401;
  assign n23403 = ~n23397 & n23402;
  assign n23404 = ~n23396 & n23403;
  assign n23405 = pi8  & n23404;
  assign n23406 = ~pi8  & ~n23404;
  assign n23407 = ~n23405 & ~n23406;
  assign n23408 = n23395 & ~n23407;
  assign n23409 = n8474 & n21198;
  assign n23410 = n9238 & n21195;
  assign n23411 = n8468 & n23211;
  assign n23412 = n9265 & n21192;
  assign n23413 = ~n23411 & ~n23412;
  assign n23414 = ~n23410 & n23413;
  assign n23415 = ~n23409 & n23414;
  assign n23416 = ~pi8  & ~n23415;
  assign n23417 = pi8  & n23415;
  assign n23418 = ~n23416 & ~n23417;
  assign n23419 = n23199 & ~n23201;
  assign n23420 = ~n23202 & ~n23419;
  assign n23421 = ~n23418 & n23420;
  assign n23422 = ~n23418 & ~n23420;
  assign n23423 = n23418 & n23420;
  assign n23424 = ~n23422 & ~n23423;
  assign n23425 = n8474 & n21201;
  assign n23426 = n9238 & n21198;
  assign n23427 = n8468 & n21482;
  assign n23428 = n9265 & n21195;
  assign n23429 = ~n23427 & ~n23428;
  assign n23430 = ~n23426 & n23429;
  assign n23431 = ~n23425 & n23430;
  assign n23432 = ~pi8  & ~n23431;
  assign n23433 = pi8  & n23431;
  assign n23434 = ~n23432 & ~n23433;
  assign n23435 = ~n23194 & n23197;
  assign n23436 = n23194 & ~n23197;
  assign n23437 = ~n23435 & ~n23436;
  assign n23438 = ~n23434 & ~n23437;
  assign n23439 = n22890 & n23192;
  assign n23440 = ~n23193 & ~n23439;
  assign n23441 = n8474 & n21204;
  assign n23442 = n9238 & n21201;
  assign n23443 = n8468 & n22832;
  assign n23444 = n9265 & n21198;
  assign n23445 = ~n23443 & ~n23444;
  assign n23446 = ~n23442 & n23445;
  assign n23447 = ~n23441 & n23446;
  assign n23448 = pi8  & n23447;
  assign n23449 = ~pi8  & ~n23447;
  assign n23450 = ~n23448 & ~n23449;
  assign n23451 = n23440 & ~n23450;
  assign n23452 = n23188 & ~n23190;
  assign n23453 = ~n23191 & ~n23452;
  assign n23454 = n8474 & n21207;
  assign n23455 = n9238 & n21204;
  assign n23456 = n8468 & n22852;
  assign n23457 = n9265 & n21201;
  assign n23458 = ~n23456 & ~n23457;
  assign n23459 = ~n23455 & n23458;
  assign n23460 = ~n23454 & n23459;
  assign n23461 = pi8  & n23460;
  assign n23462 = ~pi8  & ~n23460;
  assign n23463 = ~n23461 & ~n23462;
  assign n23464 = n23453 & ~n23463;
  assign n23465 = n22920 & n23186;
  assign n23466 = ~n23187 & ~n23465;
  assign n23467 = n8474 & n21210;
  assign n23468 = n9238 & n21207;
  assign n23469 = n8468 & n22810;
  assign n23470 = n9265 & n21204;
  assign n23471 = ~n23469 & ~n23470;
  assign n23472 = ~n23468 & n23471;
  assign n23473 = ~n23467 & n23472;
  assign n23474 = pi8  & n23473;
  assign n23475 = ~pi8  & ~n23473;
  assign n23476 = ~n23474 & ~n23475;
  assign n23477 = n23466 & ~n23476;
  assign n23478 = n8474 & n21213;
  assign n23479 = n9238 & n21210;
  assign n23480 = n8468 & n22363;
  assign n23481 = n9265 & n21207;
  assign n23482 = ~n23480 & ~n23481;
  assign n23483 = ~n23479 & n23482;
  assign n23484 = ~n23478 & n23483;
  assign n23485 = ~pi8  & ~n23484;
  assign n23486 = pi8  & n23484;
  assign n23487 = ~n23485 & ~n23486;
  assign n23488 = n23182 & ~n23184;
  assign n23489 = ~n23185 & ~n23488;
  assign n23490 = ~n23487 & n23489;
  assign n23491 = ~n23487 & ~n23489;
  assign n23492 = n23487 & n23489;
  assign n23493 = ~n23491 & ~n23492;
  assign n23494 = n8474 & n21216;
  assign n23495 = n9238 & n21213;
  assign n23496 = n8468 & n22376;
  assign n23497 = n9265 & n21210;
  assign n23498 = ~n23496 & ~n23497;
  assign n23499 = ~n23495 & n23498;
  assign n23500 = ~n23494 & n23499;
  assign n23501 = ~pi8  & ~n23500;
  assign n23502 = pi8  & n23500;
  assign n23503 = ~n23501 & ~n23502;
  assign n23504 = ~n23177 & n23180;
  assign n23505 = n23177 & ~n23180;
  assign n23506 = ~n23504 & ~n23505;
  assign n23507 = ~n23503 & ~n23506;
  assign n23508 = n8474 & n21219;
  assign n23509 = n9238 & n21216;
  assign n23510 = n8468 & n22394;
  assign n23511 = n9265 & n21213;
  assign n23512 = ~n23510 & ~n23511;
  assign n23513 = ~n23509 & n23512;
  assign n23514 = ~n23508 & n23513;
  assign n23515 = ~pi8  & ~n23514;
  assign n23516 = pi8  & n23514;
  assign n23517 = ~n23515 & ~n23516;
  assign n23518 = n23172 & n23175;
  assign n23519 = ~n23176 & ~n23518;
  assign n23520 = ~n23517 & n23519;
  assign n23521 = ~n23517 & ~n23519;
  assign n23522 = n23517 & n23519;
  assign n23523 = ~n23521 & ~n23522;
  assign n23524 = n22975 & n23170;
  assign n23525 = ~n23171 & ~n23524;
  assign n23526 = n8474 & n21222;
  assign n23527 = n9238 & n21219;
  assign n23528 = n8468 & n22225;
  assign n23529 = n9265 & n21216;
  assign n23530 = ~n23528 & ~n23529;
  assign n23531 = ~n23527 & n23530;
  assign n23532 = ~n23526 & n23531;
  assign n23533 = pi8  & n23532;
  assign n23534 = ~pi8  & ~n23532;
  assign n23535 = ~n23533 & ~n23534;
  assign n23536 = n23525 & ~n23535;
  assign n23537 = n22991 & n23168;
  assign n23538 = ~n23169 & ~n23537;
  assign n23539 = n8474 & n21225;
  assign n23540 = n9238 & n21222;
  assign n23541 = n8468 & n21973;
  assign n23542 = n9265 & n21219;
  assign n23543 = ~n23541 & ~n23542;
  assign n23544 = ~n23540 & n23543;
  assign n23545 = ~n23539 & n23544;
  assign n23546 = pi8  & n23545;
  assign n23547 = ~pi8  & ~n23545;
  assign n23548 = ~n23546 & ~n23547;
  assign n23549 = n23538 & ~n23548;
  assign n23550 = n23164 & ~n23166;
  assign n23551 = ~n23167 & ~n23550;
  assign n23552 = n8474 & n21228;
  assign n23553 = n9238 & n21225;
  assign n23554 = n8468 & n21988;
  assign n23555 = n9265 & n21222;
  assign n23556 = ~n23554 & ~n23555;
  assign n23557 = ~n23553 & n23556;
  assign n23558 = ~n23552 & n23557;
  assign n23559 = pi8  & n23558;
  assign n23560 = ~pi8  & ~n23558;
  assign n23561 = ~n23559 & ~n23560;
  assign n23562 = n23551 & ~n23561;
  assign n23563 = n8474 & n21231;
  assign n23564 = n9238 & n21228;
  assign n23565 = n8468 & n22001;
  assign n23566 = n9265 & n21225;
  assign n23567 = ~n23565 & ~n23566;
  assign n23568 = ~n23564 & n23567;
  assign n23569 = ~n23563 & n23568;
  assign n23570 = ~pi8  & ~n23569;
  assign n23571 = pi8  & n23569;
  assign n23572 = ~n23570 & ~n23571;
  assign n23573 = n23160 & ~n23162;
  assign n23574 = ~n23163 & ~n23573;
  assign n23575 = ~n23572 & n23574;
  assign n23576 = ~n23572 & ~n23574;
  assign n23577 = n23572 & n23574;
  assign n23578 = ~n23576 & ~n23577;
  assign n23579 = n8474 & n21234;
  assign n23580 = n9238 & n21231;
  assign n23581 = n8468 & n21494;
  assign n23582 = n9265 & n21228;
  assign n23583 = ~n23581 & ~n23582;
  assign n23584 = ~n23580 & n23583;
  assign n23585 = ~n23579 & n23584;
  assign n23586 = ~pi8  & ~n23585;
  assign n23587 = pi8  & n23585;
  assign n23588 = ~n23586 & ~n23587;
  assign n23589 = n23155 & n23158;
  assign n23590 = ~n23159 & ~n23589;
  assign n23591 = ~n23588 & n23590;
  assign n23592 = ~n23588 & ~n23590;
  assign n23593 = n23588 & n23590;
  assign n23594 = ~n23592 & ~n23593;
  assign n23595 = n8474 & n21237;
  assign n23596 = n9238 & n21234;
  assign n23597 = n8468 & n21789;
  assign n23598 = n9265 & n21231;
  assign n23599 = ~n23597 & ~n23598;
  assign n23600 = ~n23596 & n23599;
  assign n23601 = ~n23595 & n23600;
  assign n23602 = ~pi8  & ~n23601;
  assign n23603 = pi8  & n23601;
  assign n23604 = ~n23602 & ~n23603;
  assign n23605 = ~n23150 & n23153;
  assign n23606 = n23150 & ~n23153;
  assign n23607 = ~n23605 & ~n23606;
  assign n23608 = ~n23604 & ~n23607;
  assign n23609 = n23060 & n23148;
  assign n23610 = ~n23149 & ~n23609;
  assign n23611 = n8474 & n21240;
  assign n23612 = n9238 & n21237;
  assign n23613 = n8468 & n21807;
  assign n23614 = n9265 & n21234;
  assign n23615 = ~n23613 & ~n23614;
  assign n23616 = ~n23612 & n23615;
  assign n23617 = ~n23611 & n23616;
  assign n23618 = pi8  & n23617;
  assign n23619 = ~pi8  & ~n23617;
  assign n23620 = ~n23618 & ~n23619;
  assign n23621 = n23610 & ~n23620;
  assign n23622 = n23144 & ~n23146;
  assign n23623 = ~n23147 & ~n23622;
  assign n23624 = n8474 & n21243;
  assign n23625 = n9238 & n21240;
  assign n23626 = n8468 & n21768;
  assign n23627 = n9265 & n21237;
  assign n23628 = ~n23626 & ~n23627;
  assign n23629 = ~n23625 & n23628;
  assign n23630 = ~n23624 & n23629;
  assign n23631 = pi8  & n23630;
  assign n23632 = ~pi8  & ~n23630;
  assign n23633 = ~n23631 & ~n23632;
  assign n23634 = n23623 & ~n23633;
  assign n23635 = n23091 & n23142;
  assign n23636 = ~n23143 & ~n23635;
  assign n23637 = n8474 & n21246;
  assign n23638 = n9238 & n21243;
  assign n23639 = n8468 & n21604;
  assign n23640 = n9265 & n21240;
  assign n23641 = ~n23639 & ~n23640;
  assign n23642 = ~n23638 & n23641;
  assign n23643 = ~n23637 & n23642;
  assign n23644 = pi8  & n23643;
  assign n23645 = ~pi8  & ~n23643;
  assign n23646 = ~n23644 & ~n23645;
  assign n23647 = n23636 & ~n23646;
  assign n23648 = n8474 & n21249;
  assign n23649 = n9238 & n21246;
  assign n23650 = n8468 & n21617;
  assign n23651 = n9265 & n21243;
  assign n23652 = ~n23650 & ~n23651;
  assign n23653 = ~n23649 & n23652;
  assign n23654 = ~n23648 & n23653;
  assign n23655 = ~pi8  & ~n23654;
  assign n23656 = pi8  & n23654;
  assign n23657 = ~n23655 & ~n23656;
  assign n23658 = n23138 & ~n23140;
  assign n23659 = ~n23141 & ~n23658;
  assign n23660 = ~n23657 & n23659;
  assign n23661 = ~n23657 & ~n23659;
  assign n23662 = n23657 & n23659;
  assign n23663 = ~n23661 & ~n23662;
  assign n23664 = n8474 & n21252;
  assign n23665 = n9238 & n21249;
  assign n23666 = n8468 & n21635;
  assign n23667 = n9265 & n21246;
  assign n23668 = ~n23666 & ~n23667;
  assign n23669 = ~n23665 & n23668;
  assign n23670 = ~n23664 & n23669;
  assign n23671 = pi8  & n23670;
  assign n23672 = ~pi8  & ~n23670;
  assign n23673 = ~n23671 & ~n23672;
  assign n23674 = n23126 & n23136;
  assign n23675 = ~n23137 & ~n23674;
  assign n23676 = ~n23673 & n23675;
  assign n23677 = n8474 & n21255;
  assign n23678 = n9238 & n21252;
  assign n23679 = n8468 & n21506;
  assign n23680 = n9265 & n21249;
  assign n23681 = ~n23679 & ~n23680;
  assign n23682 = ~n23678 & n23681;
  assign n23683 = ~n23677 & n23682;
  assign n23684 = ~pi8  & ~n23683;
  assign n23685 = pi8  & n23683;
  assign n23686 = ~n23684 & ~n23685;
  assign n23687 = pi11  & ~n23114;
  assign n23688 = n23121 & ~n23687;
  assign n23689 = ~n23121 & n23687;
  assign n23690 = ~n23688 & ~n23689;
  assign n23691 = ~n23686 & n23690;
  assign n23692 = ~n23686 & ~n23690;
  assign n23693 = n23686 & n23690;
  assign n23694 = ~n23692 & ~n23693;
  assign n23695 = n8474 & n21258;
  assign n23696 = n9238 & n21255;
  assign n23697 = n8468 & n21546;
  assign n23698 = n9265 & n21252;
  assign n23699 = ~n23697 & ~n23698;
  assign n23700 = ~n23696 & n23699;
  assign n23701 = ~n23695 & n23700;
  assign n23702 = pi8  & n23701;
  assign n23703 = ~pi8  & ~n23701;
  assign n23704 = ~n23702 & ~n23703;
  assign n23705 = pi11  & n23112;
  assign n23706 = ~n23111 & n23705;
  assign n23707 = n23111 & ~n23705;
  assign n23708 = ~n23706 & ~n23707;
  assign n23709 = ~n23704 & n23708;
  assign n23710 = n8468 & ~n21519;
  assign n23711 = n9265 & n21263;
  assign n23712 = n9238 & n21265;
  assign n23713 = ~n23711 & ~n23712;
  assign n23714 = ~n23710 & n23713;
  assign n23715 = ~n8464 & n21265;
  assign n23716 = pi8  & ~n23715;
  assign n23717 = n23714 & n23716;
  assign n23718 = n8474 & n21265;
  assign n23719 = n9238 & n21263;
  assign n23720 = n8468 & ~n21531;
  assign n23721 = n9265 & n21258;
  assign n23722 = ~n23720 & ~n23721;
  assign n23723 = ~n23719 & n23722;
  assign n23724 = ~n23718 & n23723;
  assign n23725 = n23717 & n23724;
  assign n23726 = n23112 & n23725;
  assign n23727 = ~n23112 & n23725;
  assign n23728 = n23112 & ~n23725;
  assign n23729 = ~n23727 & ~n23728;
  assign n23730 = n8474 & n21263;
  assign n23731 = n9238 & n21258;
  assign n23732 = n8468 & n21583;
  assign n23733 = n9265 & n21255;
  assign n23734 = ~n23732 & ~n23733;
  assign n23735 = ~n23731 & n23734;
  assign n23736 = ~n23730 & n23735;
  assign n23737 = pi8  & n23736;
  assign n23738 = ~pi8  & ~n23736;
  assign n23739 = ~n23737 & ~n23738;
  assign n23740 = ~n23729 & ~n23739;
  assign n23741 = ~n23726 & ~n23740;
  assign n23742 = n23704 & ~n23708;
  assign n23743 = ~n23709 & ~n23742;
  assign n23744 = ~n23741 & n23743;
  assign n23745 = ~n23709 & ~n23744;
  assign n23746 = ~n23694 & ~n23745;
  assign n23747 = ~n23691 & ~n23746;
  assign n23748 = n23673 & ~n23675;
  assign n23749 = ~n23676 & ~n23748;
  assign n23750 = ~n23747 & n23749;
  assign n23751 = ~n23676 & ~n23750;
  assign n23752 = ~n23663 & ~n23751;
  assign n23753 = ~n23660 & ~n23752;
  assign n23754 = n23636 & n23646;
  assign n23755 = ~n23636 & ~n23646;
  assign n23756 = ~n23754 & ~n23755;
  assign n23757 = ~n23753 & ~n23756;
  assign n23758 = ~n23647 & ~n23757;
  assign n23759 = n23623 & n23633;
  assign n23760 = ~n23623 & ~n23633;
  assign n23761 = ~n23759 & ~n23760;
  assign n23762 = ~n23758 & ~n23761;
  assign n23763 = ~n23634 & ~n23762;
  assign n23764 = ~n23610 & n23620;
  assign n23765 = ~n23621 & ~n23764;
  assign n23766 = ~n23763 & n23765;
  assign n23767 = ~n23621 & ~n23766;
  assign n23768 = n23604 & n23607;
  assign n23769 = ~n23608 & ~n23768;
  assign n23770 = ~n23767 & n23769;
  assign n23771 = ~n23608 & ~n23770;
  assign n23772 = ~n23594 & ~n23771;
  assign n23773 = ~n23591 & ~n23772;
  assign n23774 = ~n23578 & ~n23773;
  assign n23775 = ~n23575 & ~n23774;
  assign n23776 = n23551 & n23561;
  assign n23777 = ~n23551 & ~n23561;
  assign n23778 = ~n23776 & ~n23777;
  assign n23779 = ~n23775 & ~n23778;
  assign n23780 = ~n23562 & ~n23779;
  assign n23781 = n23538 & n23548;
  assign n23782 = ~n23538 & ~n23548;
  assign n23783 = ~n23781 & ~n23782;
  assign n23784 = ~n23780 & ~n23783;
  assign n23785 = ~n23549 & ~n23784;
  assign n23786 = ~n23525 & n23535;
  assign n23787 = ~n23536 & ~n23786;
  assign n23788 = ~n23785 & n23787;
  assign n23789 = ~n23536 & ~n23788;
  assign n23790 = ~n23523 & ~n23789;
  assign n23791 = ~n23520 & ~n23790;
  assign n23792 = n23503 & n23506;
  assign n23793 = ~n23507 & ~n23792;
  assign n23794 = ~n23791 & n23793;
  assign n23795 = ~n23507 & ~n23794;
  assign n23796 = ~n23493 & ~n23795;
  assign n23797 = ~n23490 & ~n23796;
  assign n23798 = n23466 & n23476;
  assign n23799 = ~n23466 & ~n23476;
  assign n23800 = ~n23798 & ~n23799;
  assign n23801 = ~n23797 & ~n23800;
  assign n23802 = ~n23477 & ~n23801;
  assign n23803 = n23453 & n23463;
  assign n23804 = ~n23453 & ~n23463;
  assign n23805 = ~n23803 & ~n23804;
  assign n23806 = ~n23802 & ~n23805;
  assign n23807 = ~n23464 & ~n23806;
  assign n23808 = ~n23440 & n23450;
  assign n23809 = ~n23451 & ~n23808;
  assign n23810 = ~n23807 & n23809;
  assign n23811 = ~n23451 & ~n23810;
  assign n23812 = n23434 & n23437;
  assign n23813 = ~n23438 & ~n23812;
  assign n23814 = ~n23811 & n23813;
  assign n23815 = ~n23438 & ~n23814;
  assign n23816 = ~n23424 & ~n23815;
  assign n23817 = ~n23421 & ~n23816;
  assign n23818 = n23395 & n23407;
  assign n23819 = ~n23395 & ~n23407;
  assign n23820 = ~n23818 & ~n23819;
  assign n23821 = ~n23817 & ~n23820;
  assign n23822 = ~n23408 & ~n23821;
  assign n23823 = n23380 & n23392;
  assign n23824 = ~n23380 & ~n23392;
  assign n23825 = ~n23823 & ~n23824;
  assign n23826 = ~n23822 & ~n23825;
  assign n23827 = ~n23393 & ~n23826;
  assign n23828 = n23365 & n23377;
  assign n23829 = ~n23365 & ~n23377;
  assign n23830 = ~n23828 & ~n23829;
  assign n23831 = ~n23827 & ~n23830;
  assign n23832 = ~n23378 & ~n23831;
  assign n23833 = ~n23360 & ~n23364;
  assign n23834 = n7654 & n21195;
  assign n23835 = n8091 & n21192;
  assign n23836 = n7648 & n23399;
  assign n23837 = n8120 & n21189;
  assign n23838 = ~n23836 & ~n23837;
  assign n23839 = ~n23835 & n23838;
  assign n23840 = ~n23834 & n23839;
  assign n23841 = ~pi11  & ~n23840;
  assign n23842 = pi11  & n23840;
  assign n23843 = ~n23841 & ~n23842;
  assign n23844 = n23343 & ~n23353;
  assign n23845 = ~n23221 & ~n23356;
  assign n23846 = ~n23844 & ~n23845;
  assign n23847 = n6184 & n21213;
  assign n23848 = n6527 & n21210;
  assign n23849 = n6185 & n22363;
  assign n23850 = n6543 & n21207;
  assign n23851 = ~n23849 & ~n23850;
  assign n23852 = ~n23848 & n23851;
  assign n23853 = ~n23847 & n23852;
  assign n23854 = ~pi17  & ~n23853;
  assign n23855 = pi17  & n23853;
  assign n23856 = ~n23854 & ~n23855;
  assign n23857 = n23320 & ~n23330;
  assign n23858 = ~n23334 & ~n23857;
  assign n23859 = ~n23315 & ~n23319;
  assign n23860 = n5238 & n21231;
  assign n23861 = n71 & n21228;
  assign n23862 = n5239 & n22001;
  assign n23863 = n5326 & n21225;
  assign n23864 = ~n23862 & ~n23863;
  assign n23865 = ~n23861 & n23864;
  assign n23866 = ~n23860 & n23865;
  assign n23867 = ~pi23  & ~n23866;
  assign n23868 = pi23  & n23866;
  assign n23869 = ~n23867 & ~n23868;
  assign n23870 = n23298 & ~n23308;
  assign n23871 = ~n23248 & ~n23311;
  assign n23872 = ~n23870 & ~n23871;
  assign n23873 = n4006 & n21249;
  assign n23874 = n4133 & n21246;
  assign n23875 = n4002 & n21617;
  assign n23876 = n4555 & n21243;
  assign n23877 = ~n23875 & ~n23876;
  assign n23878 = ~n23874 & n23877;
  assign n23879 = ~n23873 & n23878;
  assign n23880 = ~pi29  & ~n23879;
  assign n23881 = pi29  & n23879;
  assign n23882 = ~n23880 & ~n23881;
  assign n23883 = ~n23276 & ~n23283;
  assign n23884 = ~n23289 & ~n23883;
  assign n23885 = n5150 & n12921;
  assign n23886 = ~n442 & n23885;
  assign n23887 = n1063 & n12902;
  assign n23888 = n1575 & n23887;
  assign n23889 = n777 & n23888;
  assign n23890 = ~n678 & n23889;
  assign n23891 = n23886 & n23890;
  assign n23892 = n6377 & n15191;
  assign n23893 = ~n154 & n23892;
  assign n23894 = n2436 & n21120;
  assign n23895 = ~n698 & n23894;
  assign n23896 = ~n536 & n23895;
  assign n23897 = n23893 & n23896;
  assign n23898 = n23891 & n23897;
  assign n23899 = n3641 & n21258;
  assign n23900 = n556 & n21546;
  assign n23901 = n3961 & n21252;
  assign n23902 = n3740 & n21255;
  assign n23903 = ~n23901 & ~n23902;
  assign n23904 = ~n23900 & n23903;
  assign n23905 = ~n23899 & n23904;
  assign n23906 = ~n23898 & n23905;
  assign n23907 = n23898 & ~n23905;
  assign n23908 = ~n23906 & ~n23907;
  assign n23909 = ~n23884 & ~n23908;
  assign n23910 = n23884 & n23908;
  assign n23911 = ~n23909 & ~n23910;
  assign n23912 = ~n23882 & ~n23911;
  assign n23913 = n23882 & n23911;
  assign n23914 = ~n23912 & ~n23913;
  assign n23915 = ~n23258 & n23291;
  assign n23916 = ~n23297 & ~n23915;
  assign n23917 = n23914 & n23916;
  assign n23918 = ~n23914 & ~n23916;
  assign n23919 = ~n23917 & ~n23918;
  assign n23920 = n4601 & n21240;
  assign n23921 = n4783 & n21237;
  assign n23922 = n4602 & n21807;
  assign n23923 = n4801 & n21234;
  assign n23924 = ~n23922 & ~n23923;
  assign n23925 = ~n23921 & n23924;
  assign n23926 = ~n23920 & n23925;
  assign n23927 = pi26  & n23926;
  assign n23928 = ~pi26  & ~n23926;
  assign n23929 = ~n23927 & ~n23928;
  assign n23930 = n23919 & n23929;
  assign n23931 = ~n23919 & ~n23929;
  assign n23932 = ~n23930 & ~n23931;
  assign n23933 = ~n23872 & n23932;
  assign n23934 = n23872 & ~n23932;
  assign n23935 = ~n23933 & ~n23934;
  assign n23936 = ~n23869 & ~n23935;
  assign n23937 = n23869 & n23935;
  assign n23938 = ~n23936 & ~n23937;
  assign n23939 = n23859 & ~n23938;
  assign n23940 = ~n23859 & n23938;
  assign n23941 = ~n23939 & ~n23940;
  assign n23942 = n5435 & n21222;
  assign n23943 = n6055 & n21219;
  assign n23944 = n5429 & n22225;
  assign n23945 = n6071 & n21216;
  assign n23946 = ~n23944 & ~n23945;
  assign n23947 = ~n23943 & n23946;
  assign n23948 = ~n23942 & n23947;
  assign n23949 = pi20  & n23948;
  assign n23950 = ~pi20  & ~n23948;
  assign n23951 = ~n23949 & ~n23950;
  assign n23952 = n23941 & n23951;
  assign n23953 = ~n23941 & ~n23951;
  assign n23954 = ~n23952 & ~n23953;
  assign n23955 = ~n23858 & ~n23954;
  assign n23956 = n23858 & n23954;
  assign n23957 = ~n23955 & ~n23956;
  assign n23958 = ~n23856 & ~n23957;
  assign n23959 = n23856 & n23957;
  assign n23960 = ~n23958 & ~n23959;
  assign n23961 = ~n23231 & n23336;
  assign n23962 = ~n23342 & ~n23961;
  assign n23963 = n23960 & n23962;
  assign n23964 = ~n23960 & ~n23962;
  assign n23965 = ~n23963 & ~n23964;
  assign n23966 = n6835 & n21204;
  assign n23967 = n7460 & n21201;
  assign n23968 = n6836 & n22832;
  assign n23969 = n7487 & n21198;
  assign n23970 = ~n23968 & ~n23969;
  assign n23971 = ~n23967 & n23970;
  assign n23972 = ~n23966 & n23971;
  assign n23973 = pi14  & n23972;
  assign n23974 = ~pi14  & ~n23972;
  assign n23975 = ~n23973 & ~n23974;
  assign n23976 = n23965 & n23975;
  assign n23977 = ~n23965 & ~n23975;
  assign n23978 = ~n23976 & ~n23977;
  assign n23979 = ~n23846 & n23978;
  assign n23980 = n23846 & ~n23978;
  assign n23981 = ~n23979 & ~n23980;
  assign n23982 = ~n23843 & ~n23981;
  assign n23983 = n23843 & n23981;
  assign n23984 = ~n23982 & ~n23983;
  assign n23985 = n23833 & ~n23984;
  assign n23986 = ~n23833 & n23984;
  assign n23987 = ~n23985 & ~n23986;
  assign n23988 = n8474 & n21186;
  assign n23989 = n9238 & n21183;
  assign n23990 = n21365 & ~n21367;
  assign n23991 = ~n21368 & ~n23990;
  assign n23992 = n8468 & n23991;
  assign n23993 = n9265 & n21180;
  assign n23994 = ~n23992 & ~n23993;
  assign n23995 = ~n23989 & n23994;
  assign n23996 = ~n23988 & n23995;
  assign n23997 = pi8  & n23996;
  assign n23998 = ~pi8  & ~n23996;
  assign n23999 = ~n23997 & ~n23998;
  assign n24000 = n23987 & n23999;
  assign n24001 = ~n23987 & ~n23999;
  assign n24002 = ~n24000 & ~n24001;
  assign n24003 = ~n23832 & ~n24002;
  assign n24004 = n23832 & n24002;
  assign n24005 = ~n24003 & ~n24004;
  assign n24006 = ~n21478 & ~n24005;
  assign n24007 = n21478 & n24005;
  assign n24008 = ~n24006 & ~n24007;
  assign n24009 = n9725 & n21180;
  assign n24010 = n10702 & n21076;
  assign n24011 = n21373 & ~n21375;
  assign n24012 = ~n21376 & ~n24011;
  assign n24013 = n9719 & n24012;
  assign n24014 = n11267 & n21176;
  assign n24015 = ~n24013 & ~n24014;
  assign n24016 = ~n24010 & n24015;
  assign n24017 = ~n24009 & n24016;
  assign n24018 = ~pi5  & ~n24017;
  assign n24019 = pi5  & n24017;
  assign n24020 = ~n24018 & ~n24019;
  assign n24021 = n23827 & n23830;
  assign n24022 = ~n23831 & ~n24021;
  assign n24023 = ~n24020 & n24022;
  assign n24024 = ~n24020 & ~n24022;
  assign n24025 = n24020 & n24022;
  assign n24026 = ~n24024 & ~n24025;
  assign n24027 = n9725 & n21183;
  assign n24028 = n10702 & n21180;
  assign n24029 = n21369 & ~n21371;
  assign n24030 = ~n21372 & ~n24029;
  assign n24031 = n9719 & n24030;
  assign n24032 = n11267 & n21076;
  assign n24033 = ~n24031 & ~n24032;
  assign n24034 = ~n24028 & n24033;
  assign n24035 = ~n24027 & n24034;
  assign n24036 = ~pi5  & ~n24035;
  assign n24037 = pi5  & n24035;
  assign n24038 = ~n24036 & ~n24037;
  assign n24039 = ~n23822 & n23825;
  assign n24040 = n23822 & ~n23825;
  assign n24041 = ~n24039 & ~n24040;
  assign n24042 = ~n24038 & ~n24041;
  assign n24043 = n9725 & n21186;
  assign n24044 = n10702 & n21183;
  assign n24045 = n9719 & n23991;
  assign n24046 = n11267 & n21180;
  assign n24047 = ~n24045 & ~n24046;
  assign n24048 = ~n24044 & n24047;
  assign n24049 = ~n24043 & n24048;
  assign n24050 = ~pi5  & ~n24049;
  assign n24051 = pi5  & n24049;
  assign n24052 = ~n24050 & ~n24051;
  assign n24053 = ~n23817 & n23820;
  assign n24054 = n23817 & ~n23820;
  assign n24055 = ~n24053 & ~n24054;
  assign n24056 = ~n24052 & ~n24055;
  assign n24057 = n23424 & n23815;
  assign n24058 = ~n23816 & ~n24057;
  assign n24059 = n9725 & n21189;
  assign n24060 = n10702 & n21186;
  assign n24061 = n9719 & n23369;
  assign n24062 = n11267 & n21183;
  assign n24063 = ~n24061 & ~n24062;
  assign n24064 = ~n24060 & n24063;
  assign n24065 = ~n24059 & n24064;
  assign n24066 = pi5  & n24065;
  assign n24067 = ~pi5  & ~n24065;
  assign n24068 = ~n24066 & ~n24067;
  assign n24069 = n24058 & ~n24068;
  assign n24070 = n23811 & ~n23813;
  assign n24071 = ~n23814 & ~n24070;
  assign n24072 = n9725 & n21192;
  assign n24073 = n10702 & n21189;
  assign n24074 = n9719 & n23384;
  assign n24075 = n11267 & n21186;
  assign n24076 = ~n24074 & ~n24075;
  assign n24077 = ~n24073 & n24076;
  assign n24078 = ~n24072 & n24077;
  assign n24079 = pi5  & n24078;
  assign n24080 = ~pi5  & ~n24078;
  assign n24081 = ~n24079 & ~n24080;
  assign n24082 = n24071 & ~n24081;
  assign n24083 = n9725 & n21195;
  assign n24084 = n10702 & n21192;
  assign n24085 = n9719 & n23399;
  assign n24086 = n11267 & n21189;
  assign n24087 = ~n24085 & ~n24086;
  assign n24088 = ~n24084 & n24087;
  assign n24089 = ~n24083 & n24088;
  assign n24090 = ~pi5  & ~n24089;
  assign n24091 = pi5  & n24089;
  assign n24092 = ~n24090 & ~n24091;
  assign n24093 = n23807 & ~n23809;
  assign n24094 = ~n23810 & ~n24093;
  assign n24095 = ~n24092 & n24094;
  assign n24096 = ~n24092 & ~n24094;
  assign n24097 = n24092 & n24094;
  assign n24098 = ~n24096 & ~n24097;
  assign n24099 = n9725 & n21198;
  assign n24100 = n10702 & n21195;
  assign n24101 = n9719 & n23211;
  assign n24102 = n11267 & n21192;
  assign n24103 = ~n24101 & ~n24102;
  assign n24104 = ~n24100 & n24103;
  assign n24105 = ~n24099 & n24104;
  assign n24106 = ~pi5  & ~n24105;
  assign n24107 = pi5  & n24105;
  assign n24108 = ~n24106 & ~n24107;
  assign n24109 = n23802 & n23805;
  assign n24110 = ~n23806 & ~n24109;
  assign n24111 = ~n24108 & n24110;
  assign n24112 = ~n24108 & ~n24110;
  assign n24113 = n24108 & n24110;
  assign n24114 = ~n24112 & ~n24113;
  assign n24115 = n9725 & n21201;
  assign n24116 = n10702 & n21198;
  assign n24117 = n9719 & n21482;
  assign n24118 = n11267 & n21195;
  assign n24119 = ~n24117 & ~n24118;
  assign n24120 = ~n24116 & n24119;
  assign n24121 = ~n24115 & n24120;
  assign n24122 = ~pi5  & ~n24121;
  assign n24123 = pi5  & n24121;
  assign n24124 = ~n24122 & ~n24123;
  assign n24125 = ~n23797 & n23800;
  assign n24126 = n23797 & ~n23800;
  assign n24127 = ~n24125 & ~n24126;
  assign n24128 = ~n24124 & ~n24127;
  assign n24129 = n23493 & n23795;
  assign n24130 = ~n23796 & ~n24129;
  assign n24131 = n9725 & n21204;
  assign n24132 = n10702 & n21201;
  assign n24133 = n9719 & n22832;
  assign n24134 = n11267 & n21198;
  assign n24135 = ~n24133 & ~n24134;
  assign n24136 = ~n24132 & n24135;
  assign n24137 = ~n24131 & n24136;
  assign n24138 = pi5  & n24137;
  assign n24139 = ~pi5  & ~n24137;
  assign n24140 = ~n24138 & ~n24139;
  assign n24141 = n24130 & ~n24140;
  assign n24142 = n23791 & ~n23793;
  assign n24143 = ~n23794 & ~n24142;
  assign n24144 = n9725 & n21207;
  assign n24145 = n10702 & n21204;
  assign n24146 = n9719 & n22852;
  assign n24147 = n11267 & n21201;
  assign n24148 = ~n24146 & ~n24147;
  assign n24149 = ~n24145 & n24148;
  assign n24150 = ~n24144 & n24149;
  assign n24151 = pi5  & n24150;
  assign n24152 = ~pi5  & ~n24150;
  assign n24153 = ~n24151 & ~n24152;
  assign n24154 = n24143 & ~n24153;
  assign n24155 = n23523 & n23789;
  assign n24156 = ~n23790 & ~n24155;
  assign n24157 = n9725 & n21210;
  assign n24158 = n10702 & n21207;
  assign n24159 = n9719 & n22810;
  assign n24160 = n11267 & n21204;
  assign n24161 = ~n24159 & ~n24160;
  assign n24162 = ~n24158 & n24161;
  assign n24163 = ~n24157 & n24162;
  assign n24164 = pi5  & n24163;
  assign n24165 = ~pi5  & ~n24163;
  assign n24166 = ~n24164 & ~n24165;
  assign n24167 = n24156 & ~n24166;
  assign n24168 = n9725 & n21213;
  assign n24169 = n10702 & n21210;
  assign n24170 = n9719 & n22363;
  assign n24171 = n11267 & n21207;
  assign n24172 = ~n24170 & ~n24171;
  assign n24173 = ~n24169 & n24172;
  assign n24174 = ~n24168 & n24173;
  assign n24175 = ~pi5  & ~n24174;
  assign n24176 = pi5  & n24174;
  assign n24177 = ~n24175 & ~n24176;
  assign n24178 = n23785 & ~n23787;
  assign n24179 = ~n23788 & ~n24178;
  assign n24180 = ~n24177 & n24179;
  assign n24181 = ~n24177 & ~n24179;
  assign n24182 = n24177 & n24179;
  assign n24183 = ~n24181 & ~n24182;
  assign n24184 = n9725 & n21216;
  assign n24185 = n10702 & n21213;
  assign n24186 = n9719 & n22376;
  assign n24187 = n11267 & n21210;
  assign n24188 = ~n24186 & ~n24187;
  assign n24189 = ~n24185 & n24188;
  assign n24190 = ~n24184 & n24189;
  assign n24191 = ~pi5  & ~n24190;
  assign n24192 = pi5  & n24190;
  assign n24193 = ~n24191 & ~n24192;
  assign n24194 = ~n23780 & n23783;
  assign n24195 = n23780 & ~n23783;
  assign n24196 = ~n24194 & ~n24195;
  assign n24197 = ~n24193 & ~n24196;
  assign n24198 = n9725 & n21219;
  assign n24199 = n10702 & n21216;
  assign n24200 = n9719 & n22394;
  assign n24201 = n11267 & n21213;
  assign n24202 = ~n24200 & ~n24201;
  assign n24203 = ~n24199 & n24202;
  assign n24204 = ~n24198 & n24203;
  assign n24205 = ~pi5  & ~n24204;
  assign n24206 = pi5  & n24204;
  assign n24207 = ~n24205 & ~n24206;
  assign n24208 = n23775 & n23778;
  assign n24209 = ~n23779 & ~n24208;
  assign n24210 = ~n24207 & n24209;
  assign n24211 = ~n24207 & ~n24209;
  assign n24212 = n24207 & n24209;
  assign n24213 = ~n24211 & ~n24212;
  assign n24214 = n23578 & n23773;
  assign n24215 = ~n23774 & ~n24214;
  assign n24216 = n9725 & n21222;
  assign n24217 = n10702 & n21219;
  assign n24218 = n9719 & n22225;
  assign n24219 = n11267 & n21216;
  assign n24220 = ~n24218 & ~n24219;
  assign n24221 = ~n24217 & n24220;
  assign n24222 = ~n24216 & n24221;
  assign n24223 = pi5  & n24222;
  assign n24224 = ~pi5  & ~n24222;
  assign n24225 = ~n24223 & ~n24224;
  assign n24226 = n24215 & ~n24225;
  assign n24227 = n23594 & n23771;
  assign n24228 = ~n23772 & ~n24227;
  assign n24229 = n9725 & n21225;
  assign n24230 = n10702 & n21222;
  assign n24231 = n9719 & n21973;
  assign n24232 = n11267 & n21219;
  assign n24233 = ~n24231 & ~n24232;
  assign n24234 = ~n24230 & n24233;
  assign n24235 = ~n24229 & n24234;
  assign n24236 = pi5  & n24235;
  assign n24237 = ~pi5  & ~n24235;
  assign n24238 = ~n24236 & ~n24237;
  assign n24239 = n24228 & ~n24238;
  assign n24240 = n23767 & ~n23769;
  assign n24241 = ~n23770 & ~n24240;
  assign n24242 = n9725 & n21228;
  assign n24243 = n10702 & n21225;
  assign n24244 = n9719 & n21988;
  assign n24245 = n11267 & n21222;
  assign n24246 = ~n24244 & ~n24245;
  assign n24247 = ~n24243 & n24246;
  assign n24248 = ~n24242 & n24247;
  assign n24249 = pi5  & n24248;
  assign n24250 = ~pi5  & ~n24248;
  assign n24251 = ~n24249 & ~n24250;
  assign n24252 = n24241 & ~n24251;
  assign n24253 = n9725 & n21231;
  assign n24254 = n10702 & n21228;
  assign n24255 = n9719 & n22001;
  assign n24256 = n11267 & n21225;
  assign n24257 = ~n24255 & ~n24256;
  assign n24258 = ~n24254 & n24257;
  assign n24259 = ~n24253 & n24258;
  assign n24260 = ~pi5  & ~n24259;
  assign n24261 = pi5  & n24259;
  assign n24262 = ~n24260 & ~n24261;
  assign n24263 = n23763 & ~n23765;
  assign n24264 = ~n23766 & ~n24263;
  assign n24265 = ~n24262 & n24264;
  assign n24266 = ~n24262 & ~n24264;
  assign n24267 = n24262 & n24264;
  assign n24268 = ~n24266 & ~n24267;
  assign n24269 = n9725 & n21234;
  assign n24270 = n10702 & n21231;
  assign n24271 = n9719 & n21494;
  assign n24272 = n11267 & n21228;
  assign n24273 = ~n24271 & ~n24272;
  assign n24274 = ~n24270 & n24273;
  assign n24275 = ~n24269 & n24274;
  assign n24276 = ~pi5  & ~n24275;
  assign n24277 = pi5  & n24275;
  assign n24278 = ~n24276 & ~n24277;
  assign n24279 = n23758 & n23761;
  assign n24280 = ~n23762 & ~n24279;
  assign n24281 = ~n24278 & n24280;
  assign n24282 = ~n24278 & ~n24280;
  assign n24283 = n24278 & n24280;
  assign n24284 = ~n24282 & ~n24283;
  assign n24285 = n9725 & n21237;
  assign n24286 = n10702 & n21234;
  assign n24287 = n9719 & n21789;
  assign n24288 = n11267 & n21231;
  assign n24289 = ~n24287 & ~n24288;
  assign n24290 = ~n24286 & n24289;
  assign n24291 = ~n24285 & n24290;
  assign n24292 = ~pi5  & ~n24291;
  assign n24293 = pi5  & n24291;
  assign n24294 = ~n24292 & ~n24293;
  assign n24295 = ~n23753 & n23756;
  assign n24296 = n23753 & ~n23756;
  assign n24297 = ~n24295 & ~n24296;
  assign n24298 = ~n24294 & ~n24297;
  assign n24299 = n23663 & n23751;
  assign n24300 = ~n23752 & ~n24299;
  assign n24301 = n9725 & n21240;
  assign n24302 = n10702 & n21237;
  assign n24303 = n9719 & n21807;
  assign n24304 = n11267 & n21234;
  assign n24305 = ~n24303 & ~n24304;
  assign n24306 = ~n24302 & n24305;
  assign n24307 = ~n24301 & n24306;
  assign n24308 = pi5  & n24307;
  assign n24309 = ~pi5  & ~n24307;
  assign n24310 = ~n24308 & ~n24309;
  assign n24311 = n24300 & ~n24310;
  assign n24312 = n23747 & ~n23749;
  assign n24313 = ~n23750 & ~n24312;
  assign n24314 = n9725 & n21243;
  assign n24315 = n10702 & n21240;
  assign n24316 = n9719 & n21768;
  assign n24317 = n11267 & n21237;
  assign n24318 = ~n24316 & ~n24317;
  assign n24319 = ~n24315 & n24318;
  assign n24320 = ~n24314 & n24319;
  assign n24321 = pi5  & n24320;
  assign n24322 = ~pi5  & ~n24320;
  assign n24323 = ~n24321 & ~n24322;
  assign n24324 = n24313 & ~n24323;
  assign n24325 = n23694 & n23745;
  assign n24326 = ~n23746 & ~n24325;
  assign n24327 = n9725 & n21246;
  assign n24328 = n10702 & n21243;
  assign n24329 = n9719 & n21604;
  assign n24330 = n11267 & n21240;
  assign n24331 = ~n24329 & ~n24330;
  assign n24332 = ~n24328 & n24331;
  assign n24333 = ~n24327 & n24332;
  assign n24334 = pi5  & n24333;
  assign n24335 = ~pi5  & ~n24333;
  assign n24336 = ~n24334 & ~n24335;
  assign n24337 = n24326 & ~n24336;
  assign n24338 = n9725 & n21249;
  assign n24339 = n10702 & n21246;
  assign n24340 = n9719 & n21617;
  assign n24341 = n11267 & n21243;
  assign n24342 = ~n24340 & ~n24341;
  assign n24343 = ~n24339 & n24342;
  assign n24344 = ~n24338 & n24343;
  assign n24345 = ~pi5  & ~n24344;
  assign n24346 = pi5  & n24344;
  assign n24347 = ~n24345 & ~n24346;
  assign n24348 = n23741 & ~n23743;
  assign n24349 = ~n23744 & ~n24348;
  assign n24350 = ~n24347 & n24349;
  assign n24351 = ~n24347 & ~n24349;
  assign n24352 = n24347 & n24349;
  assign n24353 = ~n24351 & ~n24352;
  assign n24354 = n9725 & n21252;
  assign n24355 = n10702 & n21249;
  assign n24356 = n9719 & n21635;
  assign n24357 = n11267 & n21246;
  assign n24358 = ~n24356 & ~n24357;
  assign n24359 = ~n24355 & n24358;
  assign n24360 = ~n24354 & n24359;
  assign n24361 = pi5  & n24360;
  assign n24362 = ~pi5  & ~n24360;
  assign n24363 = ~n24361 & ~n24362;
  assign n24364 = n23729 & n23739;
  assign n24365 = ~n23740 & ~n24364;
  assign n24366 = ~n24363 & n24365;
  assign n24367 = n9725 & n21255;
  assign n24368 = n10702 & n21252;
  assign n24369 = n9719 & n21506;
  assign n24370 = n11267 & n21249;
  assign n24371 = ~n24369 & ~n24370;
  assign n24372 = ~n24368 & n24371;
  assign n24373 = ~n24367 & n24372;
  assign n24374 = ~pi5  & ~n24373;
  assign n24375 = pi5  & n24373;
  assign n24376 = ~n24374 & ~n24375;
  assign n24377 = pi8  & ~n23717;
  assign n24378 = n23724 & ~n24377;
  assign n24379 = ~n23724 & n24377;
  assign n24380 = ~n24378 & ~n24379;
  assign n24381 = ~n24376 & n24380;
  assign n24382 = ~n24376 & ~n24380;
  assign n24383 = n24376 & n24380;
  assign n24384 = ~n24382 & ~n24383;
  assign n24385 = n9725 & n21258;
  assign n24386 = n10702 & n21255;
  assign n24387 = n9719 & n21546;
  assign n24388 = n11267 & n21252;
  assign n24389 = ~n24387 & ~n24388;
  assign n24390 = ~n24386 & n24389;
  assign n24391 = ~n24385 & n24390;
  assign n24392 = pi5  & n24391;
  assign n24393 = ~pi5  & ~n24391;
  assign n24394 = ~n24392 & ~n24393;
  assign n24395 = pi8  & n23715;
  assign n24396 = ~n23714 & n24395;
  assign n24397 = n23714 & ~n24395;
  assign n24398 = ~n24396 & ~n24397;
  assign n24399 = ~n24394 & n24398;
  assign n24400 = n9719 & ~n21519;
  assign n24401 = n11267 & n21263;
  assign n24402 = n10702 & n21265;
  assign n24403 = ~n24401 & ~n24402;
  assign n24404 = ~n24400 & n24403;
  assign n24405 = ~n9715 & n21265;
  assign n24406 = pi5  & ~n24405;
  assign n24407 = n24404 & n24406;
  assign n24408 = n9725 & n21265;
  assign n24409 = n10702 & n21263;
  assign n24410 = n9719 & ~n21531;
  assign n24411 = n11267 & n21258;
  assign n24412 = ~n24410 & ~n24411;
  assign n24413 = ~n24409 & n24412;
  assign n24414 = ~n24408 & n24413;
  assign n24415 = n24407 & n24414;
  assign n24416 = n23715 & n24415;
  assign n24417 = ~n23715 & n24415;
  assign n24418 = n23715 & ~n24415;
  assign n24419 = ~n24417 & ~n24418;
  assign n24420 = n9725 & n21263;
  assign n24421 = n10702 & n21258;
  assign n24422 = n9719 & n21583;
  assign n24423 = n11267 & n21255;
  assign n24424 = ~n24422 & ~n24423;
  assign n24425 = ~n24421 & n24424;
  assign n24426 = ~n24420 & n24425;
  assign n24427 = pi5  & n24426;
  assign n24428 = ~pi5  & ~n24426;
  assign n24429 = ~n24427 & ~n24428;
  assign n24430 = ~n24419 & ~n24429;
  assign n24431 = ~n24416 & ~n24430;
  assign n24432 = n24394 & ~n24398;
  assign n24433 = ~n24399 & ~n24432;
  assign n24434 = ~n24431 & n24433;
  assign n24435 = ~n24399 & ~n24434;
  assign n24436 = ~n24384 & ~n24435;
  assign n24437 = ~n24381 & ~n24436;
  assign n24438 = n24363 & ~n24365;
  assign n24439 = ~n24366 & ~n24438;
  assign n24440 = ~n24437 & n24439;
  assign n24441 = ~n24366 & ~n24440;
  assign n24442 = ~n24353 & ~n24441;
  assign n24443 = ~n24350 & ~n24442;
  assign n24444 = n24326 & n24336;
  assign n24445 = ~n24326 & ~n24336;
  assign n24446 = ~n24444 & ~n24445;
  assign n24447 = ~n24443 & ~n24446;
  assign n24448 = ~n24337 & ~n24447;
  assign n24449 = n24313 & n24323;
  assign n24450 = ~n24313 & ~n24323;
  assign n24451 = ~n24449 & ~n24450;
  assign n24452 = ~n24448 & ~n24451;
  assign n24453 = ~n24324 & ~n24452;
  assign n24454 = ~n24300 & n24310;
  assign n24455 = ~n24311 & ~n24454;
  assign n24456 = ~n24453 & n24455;
  assign n24457 = ~n24311 & ~n24456;
  assign n24458 = n24294 & n24297;
  assign n24459 = ~n24298 & ~n24458;
  assign n24460 = ~n24457 & n24459;
  assign n24461 = ~n24298 & ~n24460;
  assign n24462 = ~n24284 & ~n24461;
  assign n24463 = ~n24281 & ~n24462;
  assign n24464 = ~n24268 & ~n24463;
  assign n24465 = ~n24265 & ~n24464;
  assign n24466 = n24241 & n24251;
  assign n24467 = ~n24241 & ~n24251;
  assign n24468 = ~n24466 & ~n24467;
  assign n24469 = ~n24465 & ~n24468;
  assign n24470 = ~n24252 & ~n24469;
  assign n24471 = n24228 & n24238;
  assign n24472 = ~n24228 & ~n24238;
  assign n24473 = ~n24471 & ~n24472;
  assign n24474 = ~n24470 & ~n24473;
  assign n24475 = ~n24239 & ~n24474;
  assign n24476 = ~n24215 & n24225;
  assign n24477 = ~n24226 & ~n24476;
  assign n24478 = ~n24475 & n24477;
  assign n24479 = ~n24226 & ~n24478;
  assign n24480 = ~n24213 & ~n24479;
  assign n24481 = ~n24210 & ~n24480;
  assign n24482 = n24193 & n24196;
  assign n24483 = ~n24197 & ~n24482;
  assign n24484 = ~n24481 & n24483;
  assign n24485 = ~n24197 & ~n24484;
  assign n24486 = ~n24183 & ~n24485;
  assign n24487 = ~n24180 & ~n24486;
  assign n24488 = n24156 & n24166;
  assign n24489 = ~n24156 & ~n24166;
  assign n24490 = ~n24488 & ~n24489;
  assign n24491 = ~n24487 & ~n24490;
  assign n24492 = ~n24167 & ~n24491;
  assign n24493 = n24143 & n24153;
  assign n24494 = ~n24143 & ~n24153;
  assign n24495 = ~n24493 & ~n24494;
  assign n24496 = ~n24492 & ~n24495;
  assign n24497 = ~n24154 & ~n24496;
  assign n24498 = ~n24130 & n24140;
  assign n24499 = ~n24141 & ~n24498;
  assign n24500 = ~n24497 & n24499;
  assign n24501 = ~n24141 & ~n24500;
  assign n24502 = n24124 & n24127;
  assign n24503 = ~n24128 & ~n24502;
  assign n24504 = ~n24501 & n24503;
  assign n24505 = ~n24128 & ~n24504;
  assign n24506 = ~n24114 & ~n24505;
  assign n24507 = ~n24111 & ~n24506;
  assign n24508 = ~n24098 & ~n24507;
  assign n24509 = ~n24095 & ~n24508;
  assign n24510 = n24071 & n24081;
  assign n24511 = ~n24071 & ~n24081;
  assign n24512 = ~n24510 & ~n24511;
  assign n24513 = ~n24509 & ~n24512;
  assign n24514 = ~n24082 & ~n24513;
  assign n24515 = ~n24058 & n24068;
  assign n24516 = ~n24069 & ~n24515;
  assign n24517 = ~n24514 & n24516;
  assign n24518 = ~n24069 & ~n24517;
  assign n24519 = n24052 & n24055;
  assign n24520 = ~n24056 & ~n24519;
  assign n24521 = ~n24518 & n24520;
  assign n24522 = ~n24056 & ~n24521;
  assign n24523 = n24038 & n24041;
  assign n24524 = ~n24042 & ~n24523;
  assign n24525 = ~n24522 & n24524;
  assign n24526 = ~n24042 & ~n24525;
  assign n24527 = ~n24026 & ~n24526;
  assign n24528 = ~n24023 & ~n24527;
  assign n24529 = n24008 & n24528;
  assign n24530 = ~n24008 & ~n24528;
  assign n24531 = ~n24529 & ~n24530;
  assign n24532 = ~n21459 & ~n21462;
  assign n24533 = ~n21418 & ~n21420;
  assign n24534 = n140 & n985;
  assign n24535 = n1120 & n24534;
  assign n24536 = ~n207 & n24535;
  assign n24537 = n1110 & n2929;
  assign n24538 = ~n628 & n24537;
  assign n24539 = n24536 & n24538;
  assign n24540 = n257 & n24539;
  assign n24541 = ~n203 & n754;
  assign n24542 = ~n160 & n24541;
  assign n24543 = ~n527 & n1652;
  assign n24544 = ~n186 & n7305;
  assign n24545 = n24543 & n24544;
  assign n24546 = n765 & n24545;
  assign n24547 = n24542 & n24546;
  assign n24548 = n929 & n24547;
  assign n24549 = ~n500 & n24548;
  assign n24550 = n889 & n24549;
  assign n24551 = n24540 & n24550;
  assign n24552 = ~n24533 & n24551;
  assign n24553 = n24533 & ~n24551;
  assign n24554 = ~n24552 & ~n24553;
  assign n24555 = n3641 & n12636;
  assign n24556 = n556 & n13292;
  assign n24557 = n3961 & n12630;
  assign n24558 = n3740 & n12633;
  assign n24559 = ~n24557 & ~n24558;
  assign n24560 = ~n24556 & n24559;
  assign n24561 = ~n24555 & n24560;
  assign n24562 = n24554 & ~n24561;
  assign n24563 = ~n24554 & n24561;
  assign n24564 = ~n24562 & ~n24563;
  assign n24565 = ~n21425 & n21434;
  assign n24566 = ~n21426 & ~n24565;
  assign n24567 = n24564 & n24566;
  assign n24568 = ~n24564 & ~n24566;
  assign n24569 = ~n24567 & ~n24568;
  assign n24570 = n4006 & n12625;
  assign n24571 = n4133 & n12622;
  assign n24572 = n4002 & n13463;
  assign n24573 = n4555 & n12614;
  assign n24574 = ~n24572 & ~n24573;
  assign n24575 = ~n24571 & n24574;
  assign n24576 = ~n24570 & n24575;
  assign n24577 = pi29  & n24576;
  assign n24578 = ~pi29  & ~n24576;
  assign n24579 = ~n24577 & ~n24578;
  assign n24580 = n24569 & ~n24579;
  assign n24581 = ~n24569 & n24579;
  assign n24582 = ~n24580 & ~n24581;
  assign n24583 = ~n21439 & n21450;
  assign n24584 = ~n21438 & ~n24583;
  assign n24585 = n24582 & n24584;
  assign n24586 = ~n24582 & ~n24584;
  assign n24587 = ~n24585 & ~n24586;
  assign n24588 = n4601 & n12606;
  assign n24589 = n4783 & n12616;
  assign n24590 = n4602 & ~n13483;
  assign n24591 = ~n21380 & ~n24590;
  assign n24592 = ~n24589 & n24591;
  assign n24593 = ~n24588 & n24592;
  assign n24594 = pi26  & n24593;
  assign n24595 = ~pi26  & ~n24593;
  assign n24596 = ~n24594 & ~n24595;
  assign n24597 = n24587 & n24596;
  assign n24598 = ~n24587 & ~n24596;
  assign n24599 = ~n24597 & ~n24598;
  assign n24600 = ~n21389 & n21391;
  assign n24601 = ~n21454 & ~n24600;
  assign n24602 = ~n24599 & ~n24601;
  assign n24603 = n24599 & n24601;
  assign n24604 = ~n24602 & ~n24603;
  assign n24605 = ~n24532 & n24604;
  assign n24606 = n24532 & ~n24604;
  assign n24607 = ~n24605 & ~n24606;
  assign n24608 = n11288 & n24607;
  assign n24609 = ~n24602 & ~n24605;
  assign n24610 = ~n24552 & ~n24562;
  assign n24611 = n661 & n1880;
  assign n24612 = n167 & n24611;
  assign n24613 = ~n171 & n24612;
  assign n24614 = n748 & n1507;
  assign n24615 = ~n500 & n24614;
  assign n24616 = ~n535 & n24615;
  assign n24617 = n24613 & n24616;
  assign n24618 = n831 & n876;
  assign n24619 = ~n537 & n24618;
  assign n24620 = n140 & ~n578;
  assign n24621 = ~n414 & n24620;
  assign n24622 = n24619 & n24621;
  assign n24623 = n24617 & n24622;
  assign n24624 = ~n24551 & n24623;
  assign n24625 = n24551 & ~n24623;
  assign n24626 = ~n24624 & ~n24625;
  assign n24627 = n3641 & n12633;
  assign n24628 = n3740 & n12630;
  assign n24629 = n556 & ~n13227;
  assign n24630 = n3961 & n12625;
  assign n24631 = ~n24629 & ~n24630;
  assign n24632 = ~n24628 & n24631;
  assign n24633 = ~n24627 & n24632;
  assign n24634 = ~n24626 & n24633;
  assign n24635 = n24626 & ~n24633;
  assign n24636 = ~n24634 & ~n24635;
  assign n24637 = n24610 & ~n24636;
  assign n24638 = ~n24610 & n24636;
  assign n24639 = ~n24637 & ~n24638;
  assign n24640 = ~n24567 & ~n24580;
  assign n24641 = ~n24639 & n24640;
  assign n24642 = n24639 & ~n24640;
  assign n24643 = ~n24641 & ~n24642;
  assign n24644 = n4602 & ~n13499;
  assign n24645 = n4601 & ~n12611;
  assign n24646 = ~n4783 & ~n4801;
  assign n24647 = ~n24645 & n24646;
  assign n24648 = ~n12608 & ~n24647;
  assign n24649 = ~n24644 & ~n24648;
  assign n24650 = ~pi26  & ~n24649;
  assign n24651 = pi26  & n24649;
  assign n24652 = ~n24650 & ~n24651;
  assign n24653 = n4006 & n12622;
  assign n24654 = n4133 & n12614;
  assign n24655 = n4002 & ~n13310;
  assign n24656 = n4555 & n12606;
  assign n24657 = ~n24655 & ~n24656;
  assign n24658 = ~n24654 & n24657;
  assign n24659 = ~n24653 & n24658;
  assign n24660 = pi29  & n24659;
  assign n24661 = ~pi29  & ~n24659;
  assign n24662 = ~n24660 & ~n24661;
  assign n24663 = ~n24652 & n24662;
  assign n24664 = n24652 & ~n24662;
  assign n24665 = ~n24663 & ~n24664;
  assign n24666 = ~n24643 & n24665;
  assign n24667 = n24643 & ~n24665;
  assign n24668 = ~n24666 & ~n24667;
  assign n24669 = ~n24586 & ~n24596;
  assign n24670 = ~n24585 & ~n24669;
  assign n24671 = n24668 & ~n24670;
  assign n24672 = ~n24668 & n24670;
  assign n24673 = ~n24671 & ~n24672;
  assign n24674 = ~n24609 & n24673;
  assign n24675 = n24609 & ~n24673;
  assign n24676 = ~n24674 & ~n24675;
  assign n24677 = n11894 & n24676;
  assign n24678 = n24607 & n24676;
  assign n24679 = n21464 & n24607;
  assign n24680 = ~n21464 & ~n24607;
  assign n24681 = ~n24679 & ~n24680;
  assign n24682 = n21377 & ~n21465;
  assign n24683 = ~n21466 & ~n24682;
  assign n24684 = n24681 & n24683;
  assign n24685 = ~n24679 & ~n24684;
  assign n24686 = ~n24607 & ~n24676;
  assign n24687 = ~n24678 & ~n24686;
  assign n24688 = ~n24685 & n24687;
  assign n24689 = ~n24678 & ~n24688;
  assign n24690 = ~n24671 & ~n24674;
  assign n24691 = ~n24638 & ~n24642;
  assign n24692 = n4133 & n12606;
  assign n24693 = n4555 & ~n12608;
  assign n24694 = ~n12611 & n24693;
  assign n24695 = n4006 & n12614;
  assign n24696 = n4002 & n12868;
  assign n24697 = ~n24695 & ~n24696;
  assign n24698 = ~n24694 & n24697;
  assign n24699 = ~n24692 & n24698;
  assign n24700 = pi29  & n24699;
  assign n24701 = ~pi29  & ~n24699;
  assign n24702 = ~n24700 & ~n24701;
  assign n24703 = n4595 & n4600;
  assign n24704 = ~n12608 & ~n24703;
  assign n24705 = pi26  & ~n24704;
  assign n24706 = ~pi26  & n24704;
  assign n24707 = ~n24705 & ~n24706;
  assign n24708 = n510 & n716;
  assign n24709 = ~n666 & n24708;
  assign n24710 = n788 & n24709;
  assign n24711 = ~n414 & n24710;
  assign n24712 = n380 & n572;
  assign n24713 = n24711 & n24712;
  assign n24714 = n24551 & n24713;
  assign n24715 = ~n24551 & ~n24713;
  assign n24716 = ~n24714 & ~n24715;
  assign n24717 = n24707 & n24716;
  assign n24718 = ~n24707 & ~n24716;
  assign n24719 = ~n24717 & ~n24718;
  assign n24720 = ~n24625 & n24633;
  assign n24721 = ~n24624 & ~n24720;
  assign n24722 = n24719 & n24721;
  assign n24723 = ~n24719 & ~n24721;
  assign n24724 = ~n24722 & ~n24723;
  assign n24725 = n3641 & n12630;
  assign n24726 = n3740 & n12625;
  assign n24727 = n556 & n13325;
  assign n24728 = n3961 & n12622;
  assign n24729 = ~n24727 & ~n24728;
  assign n24730 = ~n24726 & n24729;
  assign n24731 = ~n24725 & n24730;
  assign n24732 = n24724 & ~n24731;
  assign n24733 = ~n24724 & n24731;
  assign n24734 = ~n24732 & ~n24733;
  assign n24735 = ~n24702 & n24734;
  assign n24736 = n24702 & ~n24734;
  assign n24737 = ~n24735 & ~n24736;
  assign n24738 = n24691 & ~n24737;
  assign n24739 = ~n24691 & n24737;
  assign n24740 = ~n24738 & ~n24739;
  assign n24741 = ~n24652 & ~n24662;
  assign n24742 = ~n24667 & ~n24741;
  assign n24743 = n24740 & ~n24742;
  assign n24744 = ~n24740 & n24742;
  assign n24745 = ~n24743 & ~n24744;
  assign n24746 = n24690 & ~n24745;
  assign n24747 = ~n24690 & n24745;
  assign n24748 = ~n24746 & ~n24747;
  assign n24749 = n24676 & n24748;
  assign n24750 = ~n24676 & ~n24748;
  assign n24751 = ~n24749 & ~n24750;
  assign n24752 = n24689 & n24751;
  assign n24753 = ~n24689 & ~n24751;
  assign n24754 = ~n24752 & ~n24753;
  assign n24755 = n11289 & ~n24754;
  assign n24756 = n11908 & n24748;
  assign n24757 = ~n24755 & ~n24756;
  assign n24758 = ~n24677 & n24757;
  assign n24759 = ~n24608 & n24758;
  assign n24760 = pi2  & n24759;
  assign n24761 = ~pi2  & ~n24759;
  assign n24762 = ~n24760 & ~n24761;
  assign n24763 = n24531 & ~n24762;
  assign n24764 = n24531 & n24762;
  assign n24765 = ~n24531 & ~n24762;
  assign n24766 = ~n24764 & ~n24765;
  assign n24767 = n11288 & n21464;
  assign n24768 = n11894 & n24607;
  assign n24769 = n24685 & ~n24687;
  assign n24770 = ~n24688 & ~n24769;
  assign n24771 = n11289 & n24770;
  assign n24772 = n11908 & n24676;
  assign n24773 = ~n24771 & ~n24772;
  assign n24774 = ~n24768 & n24773;
  assign n24775 = ~n24767 & n24774;
  assign n24776 = pi2  & n24775;
  assign n24777 = ~pi2  & ~n24775;
  assign n24778 = ~n24776 & ~n24777;
  assign n24779 = n11288 & n21176;
  assign n24780 = n11894 & n21464;
  assign n24781 = ~n24681 & ~n24683;
  assign n24782 = ~n24684 & ~n24781;
  assign n24783 = n11289 & n24782;
  assign n24784 = n11908 & n24607;
  assign n24785 = ~n24783 & ~n24784;
  assign n24786 = ~n24780 & n24785;
  assign n24787 = ~n24779 & n24786;
  assign n24788 = pi2  & n24787;
  assign n24789 = ~pi2  & ~n24787;
  assign n24790 = ~n24788 & ~n24789;
  assign n24791 = n11288 & n21076;
  assign n24792 = n11894 & n21176;
  assign n24793 = n11289 & ~n21470;
  assign n24794 = n11908 & n21464;
  assign n24795 = ~n24793 & ~n24794;
  assign n24796 = ~n24792 & n24795;
  assign n24797 = ~n24791 & n24796;
  assign n24798 = pi2  & n24797;
  assign n24799 = ~pi2  & ~n24797;
  assign n24800 = ~n24798 & ~n24799;
  assign n24801 = n24514 & ~n24516;
  assign n24802 = ~n24517 & ~n24801;
  assign n24803 = n24509 & n24512;
  assign n24804 = ~n24513 & ~n24803;
  assign n24805 = n11288 & n21186;
  assign n24806 = n11894 & n21183;
  assign n24807 = n11289 & n23991;
  assign n24808 = n11908 & n21180;
  assign n24809 = ~n24807 & ~n24808;
  assign n24810 = ~n24806 & n24809;
  assign n24811 = ~n24805 & n24810;
  assign n24812 = pi2  & n24811;
  assign n24813 = ~pi2  & ~n24811;
  assign n24814 = ~n24812 & ~n24813;
  assign n24815 = n11288 & n21189;
  assign n24816 = n11894 & n21186;
  assign n24817 = n11289 & n23369;
  assign n24818 = n11908 & n21183;
  assign n24819 = ~n24817 & ~n24818;
  assign n24820 = ~n24816 & n24819;
  assign n24821 = ~n24815 & n24820;
  assign n24822 = pi2  & n24821;
  assign n24823 = ~pi2  & ~n24821;
  assign n24824 = ~n24822 & ~n24823;
  assign n24825 = n11288 & n21192;
  assign n24826 = n11894 & n21189;
  assign n24827 = n11289 & n23384;
  assign n24828 = n11908 & n21186;
  assign n24829 = ~n24827 & ~n24828;
  assign n24830 = ~n24826 & n24829;
  assign n24831 = ~n24825 & n24830;
  assign n24832 = pi2  & n24831;
  assign n24833 = ~pi2  & ~n24831;
  assign n24834 = ~n24832 & ~n24833;
  assign n24835 = n24497 & ~n24499;
  assign n24836 = ~n24500 & ~n24835;
  assign n24837 = n24492 & n24495;
  assign n24838 = ~n24496 & ~n24837;
  assign n24839 = n24487 & n24490;
  assign n24840 = ~n24491 & ~n24839;
  assign n24841 = n11288 & n21204;
  assign n24842 = n11894 & n21201;
  assign n24843 = n11289 & n22832;
  assign n24844 = n11908 & n21198;
  assign n24845 = ~n24843 & ~n24844;
  assign n24846 = ~n24842 & n24845;
  assign n24847 = ~n24841 & n24846;
  assign n24848 = pi2  & n24847;
  assign n24849 = ~pi2  & ~n24847;
  assign n24850 = ~n24848 & ~n24849;
  assign n24851 = n11288 & n21207;
  assign n24852 = n11894 & n21204;
  assign n24853 = n11289 & n22852;
  assign n24854 = n11908 & n21201;
  assign n24855 = ~n24853 & ~n24854;
  assign n24856 = ~n24852 & n24855;
  assign n24857 = ~n24851 & n24856;
  assign n24858 = pi2  & n24857;
  assign n24859 = ~pi2  & ~n24857;
  assign n24860 = ~n24858 & ~n24859;
  assign n24861 = n11288 & n21210;
  assign n24862 = n11894 & n21207;
  assign n24863 = n11289 & n22810;
  assign n24864 = n11908 & n21204;
  assign n24865 = ~n24863 & ~n24864;
  assign n24866 = ~n24862 & n24865;
  assign n24867 = ~n24861 & n24866;
  assign n24868 = pi2  & n24867;
  assign n24869 = ~pi2  & ~n24867;
  assign n24870 = ~n24868 & ~n24869;
  assign n24871 = n24475 & ~n24477;
  assign n24872 = ~n24478 & ~n24871;
  assign n24873 = n24470 & n24473;
  assign n24874 = ~n24474 & ~n24873;
  assign n24875 = n24465 & n24468;
  assign n24876 = ~n24469 & ~n24875;
  assign n24877 = n11288 & n21222;
  assign n24878 = n11894 & n21219;
  assign n24879 = n11289 & n22225;
  assign n24880 = n11908 & n21216;
  assign n24881 = ~n24879 & ~n24880;
  assign n24882 = ~n24878 & n24881;
  assign n24883 = ~n24877 & n24882;
  assign n24884 = pi2  & n24883;
  assign n24885 = ~pi2  & ~n24883;
  assign n24886 = ~n24884 & ~n24885;
  assign n24887 = n11288 & n21225;
  assign n24888 = n11894 & n21222;
  assign n24889 = n11289 & n21973;
  assign n24890 = n11908 & n21219;
  assign n24891 = ~n24889 & ~n24890;
  assign n24892 = ~n24888 & n24891;
  assign n24893 = ~n24887 & n24892;
  assign n24894 = pi2  & n24893;
  assign n24895 = ~pi2  & ~n24893;
  assign n24896 = ~n24894 & ~n24895;
  assign n24897 = n11288 & n21228;
  assign n24898 = n11894 & n21225;
  assign n24899 = n11289 & n21988;
  assign n24900 = n11908 & n21222;
  assign n24901 = ~n24899 & ~n24900;
  assign n24902 = ~n24898 & n24901;
  assign n24903 = ~n24897 & n24902;
  assign n24904 = pi2  & n24903;
  assign n24905 = ~pi2  & ~n24903;
  assign n24906 = ~n24904 & ~n24905;
  assign n24907 = n24453 & ~n24455;
  assign n24908 = ~n24456 & ~n24907;
  assign n24909 = n24448 & n24451;
  assign n24910 = ~n24452 & ~n24909;
  assign n24911 = n24443 & n24446;
  assign n24912 = ~n24447 & ~n24911;
  assign n24913 = n11288 & n21240;
  assign n24914 = n11894 & n21237;
  assign n24915 = n11289 & n21807;
  assign n24916 = n11908 & n21234;
  assign n24917 = ~n24915 & ~n24916;
  assign n24918 = ~n24914 & n24917;
  assign n24919 = ~n24913 & n24918;
  assign n24920 = pi2  & n24919;
  assign n24921 = ~pi2  & ~n24919;
  assign n24922 = ~n24920 & ~n24921;
  assign n24923 = n11288 & n21243;
  assign n24924 = n11894 & n21240;
  assign n24925 = n11289 & n21768;
  assign n24926 = n11908 & n21237;
  assign n24927 = ~n24925 & ~n24926;
  assign n24928 = ~n24924 & n24927;
  assign n24929 = ~n24923 & n24928;
  assign n24930 = pi2  & n24929;
  assign n24931 = ~pi2  & ~n24929;
  assign n24932 = ~n24930 & ~n24931;
  assign n24933 = n11288 & n21246;
  assign n24934 = n11894 & n21243;
  assign n24935 = n11289 & n21604;
  assign n24936 = n11908 & n21240;
  assign n24937 = ~n24935 & ~n24936;
  assign n24938 = ~n24934 & n24937;
  assign n24939 = ~n24933 & n24938;
  assign n24940 = pi2  & n24939;
  assign n24941 = ~pi2  & ~n24939;
  assign n24942 = ~n24940 & ~n24941;
  assign n24943 = n24431 & ~n24433;
  assign n24944 = ~n24434 & ~n24943;
  assign n24945 = n11288 & n21252;
  assign n24946 = n11894 & n21249;
  assign n24947 = n11289 & n21635;
  assign n24948 = n11908 & n21246;
  assign n24949 = ~n24947 & ~n24948;
  assign n24950 = ~n24946 & n24949;
  assign n24951 = ~n24945 & n24950;
  assign n24952 = pi2  & n24951;
  assign n24953 = ~pi2  & ~n24951;
  assign n24954 = ~n24952 & ~n24953;
  assign n24955 = pi5  & ~n24407;
  assign n24956 = n24414 & ~n24955;
  assign n24957 = ~n24414 & n24955;
  assign n24958 = ~n24956 & ~n24957;
  assign n24959 = n11288 & n21258;
  assign n24960 = n11894 & n21255;
  assign n24961 = n11289 & n21546;
  assign n24962 = n11908 & n21252;
  assign n24963 = ~n24961 & ~n24962;
  assign n24964 = ~n24960 & n24963;
  assign n24965 = ~n24959 & n24964;
  assign n24966 = pi2  & n24965;
  assign n24967 = ~pi2  & ~n24965;
  assign n24968 = ~n24966 & ~n24967;
  assign n24969 = ~n11287 & n21265;
  assign n24970 = n11908 & n21263;
  assign n24971 = n12139 & ~n21531;
  assign n24972 = n11288 & n21265;
  assign n24973 = n11894 & n21263;
  assign n24974 = n11908 & n21258;
  assign n24975 = ~n24973 & ~n24974;
  assign n24976 = ~n24972 & n24975;
  assign n24977 = pi2  & ~n24976;
  assign n24978 = n12139 & ~n21519;
  assign n24979 = pi2  & ~n24978;
  assign n24980 = ~n24977 & n24979;
  assign n24981 = ~n24971 & n24980;
  assign n24982 = ~n24970 & n24981;
  assign n24983 = ~n24969 & n24982;
  assign n24984 = n24405 & n24983;
  assign n24985 = ~n24405 & ~n24983;
  assign n24986 = n11288 & n21263;
  assign n24987 = n11894 & n21258;
  assign n24988 = n11289 & n21583;
  assign n24989 = n11908 & n21255;
  assign n24990 = ~n24988 & ~n24989;
  assign n24991 = ~n24987 & n24990;
  assign n24992 = ~n24986 & n24991;
  assign n24993 = pi2  & ~n24992;
  assign n24994 = ~pi2  & n24992;
  assign n24995 = ~n24993 & ~n24994;
  assign n24996 = ~n24985 & n24995;
  assign n24997 = ~n24984 & ~n24996;
  assign n24998 = ~n24968 & ~n24997;
  assign n24999 = n24968 & n24997;
  assign n25000 = pi5  & n24405;
  assign n25001 = ~n24404 & n25000;
  assign n25002 = n24404 & ~n25000;
  assign n25003 = ~n25001 & ~n25002;
  assign n25004 = ~n24999 & n25003;
  assign n25005 = ~n24998 & ~n25004;
  assign n25006 = n24958 & ~n25005;
  assign n25007 = ~n24958 & n25005;
  assign n25008 = n11288 & n21255;
  assign n25009 = n11894 & n21252;
  assign n25010 = n11289 & n21506;
  assign n25011 = n11908 & n21249;
  assign n25012 = ~n25010 & ~n25011;
  assign n25013 = ~n25009 & n25012;
  assign n25014 = ~n25008 & n25013;
  assign n25015 = pi2  & ~n25014;
  assign n25016 = ~pi2  & n25014;
  assign n25017 = ~n25015 & ~n25016;
  assign n25018 = ~n25007 & n25017;
  assign n25019 = ~n25006 & ~n25018;
  assign n25020 = ~n24954 & ~n25019;
  assign n25021 = n24954 & n25019;
  assign n25022 = n24419 & n24429;
  assign n25023 = ~n24430 & ~n25022;
  assign n25024 = ~n25021 & n25023;
  assign n25025 = ~n25020 & ~n25024;
  assign n25026 = n24944 & ~n25025;
  assign n25027 = ~n24944 & n25025;
  assign n25028 = n11288 & n21249;
  assign n25029 = n11894 & n21246;
  assign n25030 = n11289 & n21617;
  assign n25031 = n11908 & n21243;
  assign n25032 = ~n25030 & ~n25031;
  assign n25033 = ~n25029 & n25032;
  assign n25034 = ~n25028 & n25033;
  assign n25035 = pi2  & ~n25034;
  assign n25036 = ~pi2  & n25034;
  assign n25037 = ~n25035 & ~n25036;
  assign n25038 = ~n25027 & n25037;
  assign n25039 = ~n25026 & ~n25038;
  assign n25040 = ~n24942 & ~n25039;
  assign n25041 = n24942 & n25039;
  assign n25042 = n24384 & n24435;
  assign n25043 = ~n24436 & ~n25042;
  assign n25044 = ~n25041 & n25043;
  assign n25045 = ~n25040 & ~n25044;
  assign n25046 = ~n24932 & ~n25045;
  assign n25047 = n24932 & n25045;
  assign n25048 = n24437 & ~n24439;
  assign n25049 = ~n24440 & ~n25048;
  assign n25050 = ~n25047 & n25049;
  assign n25051 = ~n25046 & ~n25050;
  assign n25052 = ~n24922 & ~n25051;
  assign n25053 = n24922 & n25051;
  assign n25054 = n24353 & n24441;
  assign n25055 = ~n24442 & ~n25054;
  assign n25056 = ~n25053 & n25055;
  assign n25057 = ~n25052 & ~n25056;
  assign n25058 = n24912 & ~n25057;
  assign n25059 = ~n24912 & n25057;
  assign n25060 = n11288 & n21237;
  assign n25061 = n11894 & n21234;
  assign n25062 = n11289 & n21789;
  assign n25063 = n11908 & n21231;
  assign n25064 = ~n25062 & ~n25063;
  assign n25065 = ~n25061 & n25064;
  assign n25066 = ~n25060 & n25065;
  assign n25067 = pi2  & ~n25066;
  assign n25068 = ~pi2  & n25066;
  assign n25069 = ~n25067 & ~n25068;
  assign n25070 = ~n25059 & n25069;
  assign n25071 = ~n25058 & ~n25070;
  assign n25072 = n24910 & ~n25071;
  assign n25073 = ~n24910 & n25071;
  assign n25074 = n11288 & n21234;
  assign n25075 = n11894 & n21231;
  assign n25076 = n11289 & n21494;
  assign n25077 = n11908 & n21228;
  assign n25078 = ~n25076 & ~n25077;
  assign n25079 = ~n25075 & n25078;
  assign n25080 = ~n25074 & n25079;
  assign n25081 = pi2  & ~n25080;
  assign n25082 = ~pi2  & n25080;
  assign n25083 = ~n25081 & ~n25082;
  assign n25084 = ~n25073 & n25083;
  assign n25085 = ~n25072 & ~n25084;
  assign n25086 = n24908 & ~n25085;
  assign n25087 = ~n24908 & n25085;
  assign n25088 = n11288 & n21231;
  assign n25089 = n11894 & n21228;
  assign n25090 = n11289 & n22001;
  assign n25091 = n11908 & n21225;
  assign n25092 = ~n25090 & ~n25091;
  assign n25093 = ~n25089 & n25092;
  assign n25094 = ~n25088 & n25093;
  assign n25095 = pi2  & ~n25094;
  assign n25096 = ~pi2  & n25094;
  assign n25097 = ~n25095 & ~n25096;
  assign n25098 = ~n25087 & n25097;
  assign n25099 = ~n25086 & ~n25098;
  assign n25100 = ~n24906 & ~n25099;
  assign n25101 = n24906 & n25099;
  assign n25102 = n24457 & ~n24459;
  assign n25103 = ~n24460 & ~n25102;
  assign n25104 = ~n25101 & n25103;
  assign n25105 = ~n25100 & ~n25104;
  assign n25106 = ~n24896 & ~n25105;
  assign n25107 = n24896 & n25105;
  assign n25108 = n24284 & n24461;
  assign n25109 = ~n24462 & ~n25108;
  assign n25110 = ~n25107 & n25109;
  assign n25111 = ~n25106 & ~n25110;
  assign n25112 = ~n24886 & ~n25111;
  assign n25113 = n24886 & n25111;
  assign n25114 = n24268 & n24463;
  assign n25115 = ~n24464 & ~n25114;
  assign n25116 = ~n25113 & n25115;
  assign n25117 = ~n25112 & ~n25116;
  assign n25118 = n24876 & ~n25117;
  assign n25119 = ~n24876 & n25117;
  assign n25120 = n11288 & n21219;
  assign n25121 = n11894 & n21216;
  assign n25122 = n11289 & n22394;
  assign n25123 = n11908 & n21213;
  assign n25124 = ~n25122 & ~n25123;
  assign n25125 = ~n25121 & n25124;
  assign n25126 = ~n25120 & n25125;
  assign n25127 = pi2  & ~n25126;
  assign n25128 = ~pi2  & n25126;
  assign n25129 = ~n25127 & ~n25128;
  assign n25130 = ~n25119 & n25129;
  assign n25131 = ~n25118 & ~n25130;
  assign n25132 = n24874 & ~n25131;
  assign n25133 = ~n24874 & n25131;
  assign n25134 = n11288 & n21216;
  assign n25135 = n11894 & n21213;
  assign n25136 = n11289 & n22376;
  assign n25137 = n11908 & n21210;
  assign n25138 = ~n25136 & ~n25137;
  assign n25139 = ~n25135 & n25138;
  assign n25140 = ~n25134 & n25139;
  assign n25141 = pi2  & ~n25140;
  assign n25142 = ~pi2  & n25140;
  assign n25143 = ~n25141 & ~n25142;
  assign n25144 = ~n25133 & n25143;
  assign n25145 = ~n25132 & ~n25144;
  assign n25146 = n24872 & ~n25145;
  assign n25147 = ~n24872 & n25145;
  assign n25148 = n11288 & n21213;
  assign n25149 = n11894 & n21210;
  assign n25150 = n11289 & n22363;
  assign n25151 = n11908 & n21207;
  assign n25152 = ~n25150 & ~n25151;
  assign n25153 = ~n25149 & n25152;
  assign n25154 = ~n25148 & n25153;
  assign n25155 = pi2  & ~n25154;
  assign n25156 = ~pi2  & n25154;
  assign n25157 = ~n25155 & ~n25156;
  assign n25158 = ~n25147 & n25157;
  assign n25159 = ~n25146 & ~n25158;
  assign n25160 = ~n24870 & ~n25159;
  assign n25161 = n24870 & n25159;
  assign n25162 = n24213 & n24479;
  assign n25163 = ~n24480 & ~n25162;
  assign n25164 = ~n25161 & n25163;
  assign n25165 = ~n25160 & ~n25164;
  assign n25166 = ~n24860 & ~n25165;
  assign n25167 = n24860 & n25165;
  assign n25168 = n24481 & ~n24483;
  assign n25169 = ~n24484 & ~n25168;
  assign n25170 = ~n25167 & n25169;
  assign n25171 = ~n25166 & ~n25170;
  assign n25172 = ~n24850 & ~n25171;
  assign n25173 = n24850 & n25171;
  assign n25174 = n24183 & n24485;
  assign n25175 = ~n24486 & ~n25174;
  assign n25176 = ~n25173 & n25175;
  assign n25177 = ~n25172 & ~n25176;
  assign n25178 = n24840 & ~n25177;
  assign n25179 = ~n24840 & n25177;
  assign n25180 = n11288 & n21201;
  assign n25181 = n11894 & n21198;
  assign n25182 = n11289 & n21482;
  assign n25183 = n11908 & n21195;
  assign n25184 = ~n25182 & ~n25183;
  assign n25185 = ~n25181 & n25184;
  assign n25186 = ~n25180 & n25185;
  assign n25187 = pi2  & ~n25186;
  assign n25188 = ~pi2  & n25186;
  assign n25189 = ~n25187 & ~n25188;
  assign n25190 = ~n25179 & n25189;
  assign n25191 = ~n25178 & ~n25190;
  assign n25192 = n24838 & ~n25191;
  assign n25193 = ~n24838 & n25191;
  assign n25194 = n11288 & n21198;
  assign n25195 = n11894 & n21195;
  assign n25196 = n11289 & n23211;
  assign n25197 = n11908 & n21192;
  assign n25198 = ~n25196 & ~n25197;
  assign n25199 = ~n25195 & n25198;
  assign n25200 = ~n25194 & n25199;
  assign n25201 = pi2  & ~n25200;
  assign n25202 = ~pi2  & n25200;
  assign n25203 = ~n25201 & ~n25202;
  assign n25204 = ~n25193 & n25203;
  assign n25205 = ~n25192 & ~n25204;
  assign n25206 = n24836 & ~n25205;
  assign n25207 = ~n24836 & n25205;
  assign n25208 = n11288 & n21195;
  assign n25209 = n11894 & n21192;
  assign n25210 = n11289 & n23399;
  assign n25211 = n11908 & n21189;
  assign n25212 = ~n25210 & ~n25211;
  assign n25213 = ~n25209 & n25212;
  assign n25214 = ~n25208 & n25213;
  assign n25215 = pi2  & ~n25214;
  assign n25216 = ~pi2  & n25214;
  assign n25217 = ~n25215 & ~n25216;
  assign n25218 = ~n25207 & n25217;
  assign n25219 = ~n25206 & ~n25218;
  assign n25220 = ~n24834 & ~n25219;
  assign n25221 = n24834 & n25219;
  assign n25222 = n24501 & ~n24503;
  assign n25223 = ~n24504 & ~n25222;
  assign n25224 = ~n25221 & n25223;
  assign n25225 = ~n25220 & ~n25224;
  assign n25226 = ~n24824 & ~n25225;
  assign n25227 = n24824 & n25225;
  assign n25228 = n24114 & n24505;
  assign n25229 = ~n24506 & ~n25228;
  assign n25230 = ~n25227 & n25229;
  assign n25231 = ~n25226 & ~n25230;
  assign n25232 = ~n24814 & ~n25231;
  assign n25233 = n24814 & n25231;
  assign n25234 = n24098 & n24507;
  assign n25235 = ~n24508 & ~n25234;
  assign n25236 = ~n25233 & n25235;
  assign n25237 = ~n25232 & ~n25236;
  assign n25238 = n24804 & ~n25237;
  assign n25239 = ~n24804 & n25237;
  assign n25240 = n11288 & n21183;
  assign n25241 = n11894 & n21180;
  assign n25242 = n11289 & n24030;
  assign n25243 = n11908 & n21076;
  assign n25244 = ~n25242 & ~n25243;
  assign n25245 = ~n25241 & n25244;
  assign n25246 = ~n25240 & n25245;
  assign n25247 = pi2  & ~n25246;
  assign n25248 = ~pi2  & n25246;
  assign n25249 = ~n25247 & ~n25248;
  assign n25250 = ~n25239 & n25249;
  assign n25251 = ~n25238 & ~n25250;
  assign n25252 = n24802 & ~n25251;
  assign n25253 = ~n24802 & n25251;
  assign n25254 = n11288 & n21180;
  assign n25255 = n11894 & n21076;
  assign n25256 = n11289 & n24012;
  assign n25257 = n11908 & n21176;
  assign n25258 = ~n25256 & ~n25257;
  assign n25259 = ~n25255 & n25258;
  assign n25260 = ~n25254 & n25259;
  assign n25261 = pi2  & ~n25260;
  assign n25262 = ~pi2  & n25260;
  assign n25263 = ~n25261 & ~n25262;
  assign n25264 = ~n25253 & n25263;
  assign n25265 = ~n25252 & ~n25264;
  assign n25266 = ~n24800 & ~n25265;
  assign n25267 = n24800 & n25265;
  assign n25268 = n24518 & ~n24520;
  assign n25269 = ~n24521 & ~n25268;
  assign n25270 = ~n25267 & n25269;
  assign n25271 = ~n25266 & ~n25270;
  assign n25272 = ~n24790 & ~n25271;
  assign n25273 = n24790 & n25271;
  assign n25274 = n24522 & ~n24524;
  assign n25275 = ~n24525 & ~n25274;
  assign n25276 = ~n25273 & n25275;
  assign n25277 = ~n25272 & ~n25276;
  assign n25278 = ~n24778 & ~n25277;
  assign n25279 = n24778 & n25277;
  assign n25280 = n24026 & n24526;
  assign n25281 = ~n24527 & ~n25280;
  assign n25282 = ~n25279 & n25281;
  assign n25283 = ~n25278 & ~n25282;
  assign n25284 = ~n24766 & ~n25283;
  assign n25285 = ~n24763 & ~n25284;
  assign n25286 = n9725 & n21176;
  assign n25287 = n10702 & n21464;
  assign n25288 = n9719 & n24782;
  assign n25289 = n11267 & n24607;
  assign n25290 = ~n25288 & ~n25289;
  assign n25291 = ~n25287 & n25290;
  assign n25292 = ~n25286 & n25291;
  assign n25293 = ~pi5  & ~n25292;
  assign n25294 = pi5  & n25292;
  assign n25295 = ~n25293 & ~n25294;
  assign n25296 = n23987 & ~n23999;
  assign n25297 = ~n24003 & ~n25296;
  assign n25298 = ~n23982 & ~n23986;
  assign n25299 = n7654 & n21192;
  assign n25300 = n8091 & n21189;
  assign n25301 = n7648 & n23384;
  assign n25302 = n8120 & n21186;
  assign n25303 = ~n25301 & ~n25302;
  assign n25304 = ~n25300 & n25303;
  assign n25305 = ~n25299 & n25304;
  assign n25306 = ~pi11  & ~n25305;
  assign n25307 = pi11  & n25305;
  assign n25308 = ~n25306 & ~n25307;
  assign n25309 = n23965 & ~n23975;
  assign n25310 = ~n23846 & ~n23978;
  assign n25311 = ~n25309 & ~n25310;
  assign n25312 = n6184 & n21210;
  assign n25313 = n6527 & n21207;
  assign n25314 = n6185 & n22810;
  assign n25315 = n6543 & n21204;
  assign n25316 = ~n25314 & ~n25315;
  assign n25317 = ~n25313 & n25316;
  assign n25318 = ~n25312 & n25317;
  assign n25319 = ~pi17  & ~n25318;
  assign n25320 = pi17  & n25318;
  assign n25321 = ~n25319 & ~n25320;
  assign n25322 = n23941 & ~n23951;
  assign n25323 = ~n23955 & ~n25322;
  assign n25324 = ~n23936 & ~n23940;
  assign n25325 = n5238 & n21228;
  assign n25326 = n71 & n21225;
  assign n25327 = n5239 & n21988;
  assign n25328 = n5326 & n21222;
  assign n25329 = ~n25327 & ~n25328;
  assign n25330 = ~n25326 & n25329;
  assign n25331 = ~n25325 & n25330;
  assign n25332 = ~pi23  & ~n25331;
  assign n25333 = pi23  & n25331;
  assign n25334 = ~n25332 & ~n25333;
  assign n25335 = n23919 & ~n23929;
  assign n25336 = ~n23872 & ~n23932;
  assign n25337 = ~n25335 & ~n25336;
  assign n25338 = n4006 & n21246;
  assign n25339 = n4133 & n21243;
  assign n25340 = n4002 & n21604;
  assign n25341 = n4555 & n21240;
  assign n25342 = ~n25340 & ~n25341;
  assign n25343 = ~n25339 & n25342;
  assign n25344 = ~n25338 & n25343;
  assign n25345 = ~pi29  & ~n25344;
  assign n25346 = pi29  & n25344;
  assign n25347 = ~n25345 & ~n25346;
  assign n25348 = ~n23898 & ~n23905;
  assign n25349 = ~n23909 & ~n25348;
  assign n25350 = n4501 & n12948;
  assign n25351 = n3693 & n13089;
  assign n25352 = n1265 & n25351;
  assign n25353 = n25350 & n25352;
  assign n25354 = ~n173 & n25353;
  assign n25355 = ~n218 & n25354;
  assign n25356 = ~n534 & n2060;
  assign n25357 = n2662 & n5109;
  assign n25358 = n1089 & n5497;
  assign n25359 = n1767 & n25358;
  assign n25360 = n25357 & n25359;
  assign n25361 = ~n289 & n25360;
  assign n25362 = n25356 & n25361;
  assign n25363 = n901 & n25362;
  assign n25364 = n25355 & n25363;
  assign n25365 = n3641 & n21255;
  assign n25366 = n556 & n21506;
  assign n25367 = n3961 & n21249;
  assign n25368 = n3740 & n21252;
  assign n25369 = ~n25367 & ~n25368;
  assign n25370 = ~n25366 & n25369;
  assign n25371 = ~n25365 & n25370;
  assign n25372 = ~n25364 & n25371;
  assign n25373 = n25364 & ~n25371;
  assign n25374 = ~n25372 & ~n25373;
  assign n25375 = ~n25349 & ~n25374;
  assign n25376 = n25349 & n25374;
  assign n25377 = ~n25375 & ~n25376;
  assign n25378 = ~n25347 & ~n25377;
  assign n25379 = n25347 & n25377;
  assign n25380 = ~n25378 & ~n25379;
  assign n25381 = ~n23882 & n23911;
  assign n25382 = ~n23918 & ~n25381;
  assign n25383 = n25380 & n25382;
  assign n25384 = ~n25380 & ~n25382;
  assign n25385 = ~n25383 & ~n25384;
  assign n25386 = n4601 & n21237;
  assign n25387 = n4783 & n21234;
  assign n25388 = n4602 & n21789;
  assign n25389 = n4801 & n21231;
  assign n25390 = ~n25388 & ~n25389;
  assign n25391 = ~n25387 & n25390;
  assign n25392 = ~n25386 & n25391;
  assign n25393 = pi26  & n25392;
  assign n25394 = ~pi26  & ~n25392;
  assign n25395 = ~n25393 & ~n25394;
  assign n25396 = n25385 & n25395;
  assign n25397 = ~n25385 & ~n25395;
  assign n25398 = ~n25396 & ~n25397;
  assign n25399 = ~n25337 & n25398;
  assign n25400 = n25337 & ~n25398;
  assign n25401 = ~n25399 & ~n25400;
  assign n25402 = ~n25334 & ~n25401;
  assign n25403 = n25334 & n25401;
  assign n25404 = ~n25402 & ~n25403;
  assign n25405 = n25324 & ~n25404;
  assign n25406 = ~n25324 & n25404;
  assign n25407 = ~n25405 & ~n25406;
  assign n25408 = n5435 & n21219;
  assign n25409 = n6055 & n21216;
  assign n25410 = n5429 & n22394;
  assign n25411 = n6071 & n21213;
  assign n25412 = ~n25410 & ~n25411;
  assign n25413 = ~n25409 & n25412;
  assign n25414 = ~n25408 & n25413;
  assign n25415 = pi20  & n25414;
  assign n25416 = ~pi20  & ~n25414;
  assign n25417 = ~n25415 & ~n25416;
  assign n25418 = n25407 & n25417;
  assign n25419 = ~n25407 & ~n25417;
  assign n25420 = ~n25418 & ~n25419;
  assign n25421 = ~n25323 & ~n25420;
  assign n25422 = n25323 & n25420;
  assign n25423 = ~n25421 & ~n25422;
  assign n25424 = ~n25321 & ~n25423;
  assign n25425 = n25321 & n25423;
  assign n25426 = ~n25424 & ~n25425;
  assign n25427 = ~n23856 & n23957;
  assign n25428 = ~n23964 & ~n25427;
  assign n25429 = n25426 & n25428;
  assign n25430 = ~n25426 & ~n25428;
  assign n25431 = ~n25429 & ~n25430;
  assign n25432 = n6835 & n21201;
  assign n25433 = n7460 & n21198;
  assign n25434 = n6836 & n21482;
  assign n25435 = n7487 & n21195;
  assign n25436 = ~n25434 & ~n25435;
  assign n25437 = ~n25433 & n25436;
  assign n25438 = ~n25432 & n25437;
  assign n25439 = pi14  & n25438;
  assign n25440 = ~pi14  & ~n25438;
  assign n25441 = ~n25439 & ~n25440;
  assign n25442 = n25431 & n25441;
  assign n25443 = ~n25431 & ~n25441;
  assign n25444 = ~n25442 & ~n25443;
  assign n25445 = ~n25311 & n25444;
  assign n25446 = n25311 & ~n25444;
  assign n25447 = ~n25445 & ~n25446;
  assign n25448 = ~n25308 & ~n25447;
  assign n25449 = n25308 & n25447;
  assign n25450 = ~n25448 & ~n25449;
  assign n25451 = n25298 & ~n25450;
  assign n25452 = ~n25298 & n25450;
  assign n25453 = ~n25451 & ~n25452;
  assign n25454 = n8474 & n21183;
  assign n25455 = n9238 & n21180;
  assign n25456 = n8468 & n24030;
  assign n25457 = n9265 & n21076;
  assign n25458 = ~n25456 & ~n25457;
  assign n25459 = ~n25455 & n25458;
  assign n25460 = ~n25454 & n25459;
  assign n25461 = pi8  & n25460;
  assign n25462 = ~pi8  & ~n25460;
  assign n25463 = ~n25461 & ~n25462;
  assign n25464 = n25453 & n25463;
  assign n25465 = ~n25453 & ~n25463;
  assign n25466 = ~n25464 & ~n25465;
  assign n25467 = ~n25297 & ~n25466;
  assign n25468 = n25297 & n25466;
  assign n25469 = ~n25467 & ~n25468;
  assign n25470 = ~n25295 & ~n25469;
  assign n25471 = n25295 & n25469;
  assign n25472 = ~n25470 & ~n25471;
  assign n25473 = ~n21478 & n24005;
  assign n25474 = ~n24530 & ~n25473;
  assign n25475 = n25472 & n25474;
  assign n25476 = ~n25472 & ~n25474;
  assign n25477 = ~n25475 & ~n25476;
  assign n25478 = n11288 & n24676;
  assign n25479 = n11894 & n24748;
  assign n25480 = ~n24743 & ~n24747;
  assign n25481 = ~n24735 & ~n24739;
  assign n25482 = ~n24715 & ~n24717;
  assign n25483 = n650 & n24709;
  assign n25484 = n524 & n25483;
  assign n25485 = ~n25482 & n25484;
  assign n25486 = n25482 & ~n25484;
  assign n25487 = ~n25485 & ~n25486;
  assign n25488 = n3641 & n12625;
  assign n25489 = n3740 & n12622;
  assign n25490 = n556 & n13463;
  assign n25491 = n3961 & n12614;
  assign n25492 = ~n25490 & ~n25491;
  assign n25493 = ~n25489 & n25492;
  assign n25494 = ~n25488 & n25493;
  assign n25495 = n25487 & ~n25494;
  assign n25496 = ~n25487 & n25494;
  assign n25497 = ~n25495 & ~n25496;
  assign n25498 = ~n24722 & n24731;
  assign n25499 = ~n24723 & ~n25498;
  assign n25500 = ~n25497 & ~n25499;
  assign n25501 = n25497 & n25499;
  assign n25502 = ~n25500 & ~n25501;
  assign n25503 = n4006 & n12606;
  assign n25504 = n4133 & ~n12608;
  assign n25505 = ~n12611 & n25504;
  assign n25506 = n4002 & ~n13483;
  assign n25507 = ~n24693 & ~n25506;
  assign n25508 = ~n25505 & n25507;
  assign n25509 = ~n25503 & n25508;
  assign n25510 = pi29  & n25509;
  assign n25511 = ~pi29  & ~n25509;
  assign n25512 = ~n25510 & ~n25511;
  assign n25513 = n25502 & ~n25512;
  assign n25514 = ~n25502 & n25512;
  assign n25515 = ~n25513 & ~n25514;
  assign n25516 = ~n25481 & n25515;
  assign n25517 = n25481 & ~n25515;
  assign n25518 = ~n25516 & ~n25517;
  assign n25519 = ~n25480 & n25518;
  assign n25520 = n25480 & ~n25518;
  assign n25521 = ~n25519 & ~n25520;
  assign n25522 = n24748 & n25521;
  assign n25523 = ~n24748 & ~n25521;
  assign n25524 = ~n25522 & ~n25523;
  assign n25525 = n24689 & ~n24749;
  assign n25526 = ~n24750 & ~n25525;
  assign n25527 = n25524 & ~n25526;
  assign n25528 = ~n25524 & n25526;
  assign n25529 = ~n25527 & ~n25528;
  assign n25530 = n11289 & ~n25529;
  assign n25531 = n11908 & n25521;
  assign n25532 = ~n25530 & ~n25531;
  assign n25533 = ~n25479 & n25532;
  assign n25534 = ~n25478 & n25533;
  assign n25535 = pi2  & n25534;
  assign n25536 = ~pi2  & ~n25534;
  assign n25537 = ~n25535 & ~n25536;
  assign n25538 = n25477 & ~n25537;
  assign n25539 = ~n25477 & n25537;
  assign n25540 = ~n25538 & ~n25539;
  assign n25541 = ~n25285 & n25540;
  assign n25542 = n25285 & ~n25540;
  assign n25543 = ~n25541 & ~n25542;
  assign n25544 = n24766 & ~n25283;
  assign n25545 = ~n24766 & n25283;
  assign n25546 = ~n25544 & ~n25545;
  assign n25547 = n25543 & ~n25546;
  assign n25548 = ~n25543 & n25546;
  assign po0  = ~n25547 & ~n25548;
  assign n25550 = ~n25538 & ~n25541;
  assign n25551 = ~n25295 & n25469;
  assign n25552 = ~n25476 & ~n25551;
  assign n25553 = n9725 & n21464;
  assign n25554 = n10702 & n24607;
  assign n25555 = n9719 & n24770;
  assign n25556 = n11267 & n24676;
  assign n25557 = ~n25555 & ~n25556;
  assign n25558 = ~n25554 & n25557;
  assign n25559 = ~n25553 & n25558;
  assign n25560 = ~pi5  & ~n25559;
  assign n25561 = pi5  & n25559;
  assign n25562 = ~n25560 & ~n25561;
  assign n25563 = n25453 & ~n25463;
  assign n25564 = ~n25467 & ~n25563;
  assign n25565 = n7654 & n21189;
  assign n25566 = n8091 & n21186;
  assign n25567 = n7648 & n23369;
  assign n25568 = n8120 & n21183;
  assign n25569 = ~n25567 & ~n25568;
  assign n25570 = ~n25566 & n25569;
  assign n25571 = ~n25565 & n25570;
  assign n25572 = ~pi11  & ~n25571;
  assign n25573 = pi11  & n25571;
  assign n25574 = ~n25572 & ~n25573;
  assign n25575 = n25431 & ~n25441;
  assign n25576 = ~n25311 & ~n25444;
  assign n25577 = ~n25575 & ~n25576;
  assign n25578 = ~n25321 & n25423;
  assign n25579 = ~n25430 & ~n25578;
  assign n25580 = n6184 & n21207;
  assign n25581 = n6527 & n21204;
  assign n25582 = n6185 & n22852;
  assign n25583 = n6543 & n21201;
  assign n25584 = ~n25582 & ~n25583;
  assign n25585 = ~n25581 & n25584;
  assign n25586 = ~n25580 & n25585;
  assign n25587 = ~pi17  & ~n25586;
  assign n25588 = pi17  & n25586;
  assign n25589 = ~n25587 & ~n25588;
  assign n25590 = n25407 & ~n25417;
  assign n25591 = ~n25421 & ~n25590;
  assign n25592 = n5238 & n21225;
  assign n25593 = n71 & n21222;
  assign n25594 = n5239 & n21973;
  assign n25595 = n5326 & n21219;
  assign n25596 = ~n25594 & ~n25595;
  assign n25597 = ~n25593 & n25596;
  assign n25598 = ~n25592 & n25597;
  assign n25599 = ~pi23  & ~n25598;
  assign n25600 = pi23  & n25598;
  assign n25601 = ~n25599 & ~n25600;
  assign n25602 = n25385 & ~n25395;
  assign n25603 = ~n25337 & ~n25398;
  assign n25604 = ~n25602 & ~n25603;
  assign n25605 = ~n25347 & n25377;
  assign n25606 = ~n25384 & ~n25605;
  assign n25607 = n4006 & n21243;
  assign n25608 = n4133 & n21240;
  assign n25609 = n4002 & n21768;
  assign n25610 = n4555 & n21237;
  assign n25611 = ~n25609 & ~n25610;
  assign n25612 = ~n25608 & n25611;
  assign n25613 = ~n25607 & n25612;
  assign n25614 = pi29  & n25613;
  assign n25615 = ~pi29  & ~n25613;
  assign n25616 = ~n25614 & ~n25615;
  assign n25617 = ~n25364 & ~n25371;
  assign n25618 = ~n25375 & ~n25617;
  assign n25619 = n3157 & n7238;
  assign n25620 = ~n401 & n25619;
  assign n25621 = n1024 & n13867;
  assign n25622 = ~n88 & n25621;
  assign n25623 = ~n349 & n25622;
  assign n25624 = n25620 & n25623;
  assign n25625 = n2427 & n7153;
  assign n25626 = n2409 & n25625;
  assign n25627 = n2340 & n25626;
  assign n25628 = ~n155 & n25627;
  assign n25629 = n1215 & n2757;
  assign n25630 = n1258 & n25629;
  assign n25631 = n148 & n25630;
  assign n25632 = n2060 & n25631;
  assign n25633 = ~n500 & n25632;
  assign n25634 = ~n259 & n25633;
  assign n25635 = n25628 & n25634;
  assign n25636 = n25624 & n25635;
  assign n25637 = n3641 & n21252;
  assign n25638 = n556 & n21635;
  assign n25639 = n3961 & n21246;
  assign n25640 = n3740 & n21249;
  assign n25641 = ~n25639 & ~n25640;
  assign n25642 = ~n25638 & n25641;
  assign n25643 = ~n25637 & n25642;
  assign n25644 = ~n25636 & n25643;
  assign n25645 = n25636 & ~n25643;
  assign n25646 = ~n25644 & ~n25645;
  assign n25647 = ~n25618 & ~n25646;
  assign n25648 = n25618 & n25646;
  assign n25649 = ~n25647 & ~n25648;
  assign n25650 = ~n25616 & n25649;
  assign n25651 = n25616 & ~n25649;
  assign n25652 = ~n25650 & ~n25651;
  assign n25653 = ~n25606 & n25652;
  assign n25654 = n25606 & ~n25652;
  assign n25655 = ~n25653 & ~n25654;
  assign n25656 = n4601 & n21234;
  assign n25657 = n4783 & n21231;
  assign n25658 = n4602 & n21494;
  assign n25659 = n4801 & n21228;
  assign n25660 = ~n25658 & ~n25659;
  assign n25661 = ~n25657 & n25660;
  assign n25662 = ~n25656 & n25661;
  assign n25663 = pi26  & n25662;
  assign n25664 = ~pi26  & ~n25662;
  assign n25665 = ~n25663 & ~n25664;
  assign n25666 = n25655 & n25665;
  assign n25667 = ~n25655 & ~n25665;
  assign n25668 = ~n25666 & ~n25667;
  assign n25669 = ~n25604 & ~n25668;
  assign n25670 = n25604 & n25668;
  assign n25671 = ~n25669 & ~n25670;
  assign n25672 = ~n25601 & ~n25671;
  assign n25673 = n25601 & n25671;
  assign n25674 = ~n25672 & ~n25673;
  assign n25675 = ~n25402 & ~n25406;
  assign n25676 = n25674 & n25675;
  assign n25677 = ~n25674 & ~n25675;
  assign n25678 = ~n25676 & ~n25677;
  assign n25679 = n5435 & n21216;
  assign n25680 = n6055 & n21213;
  assign n25681 = n5429 & n22376;
  assign n25682 = n6071 & n21210;
  assign n25683 = ~n25681 & ~n25682;
  assign n25684 = ~n25680 & n25683;
  assign n25685 = ~n25679 & n25684;
  assign n25686 = pi20  & n25685;
  assign n25687 = ~pi20  & ~n25685;
  assign n25688 = ~n25686 & ~n25687;
  assign n25689 = n25678 & n25688;
  assign n25690 = ~n25678 & ~n25688;
  assign n25691 = ~n25689 & ~n25690;
  assign n25692 = ~n25591 & n25691;
  assign n25693 = n25591 & ~n25691;
  assign n25694 = ~n25692 & ~n25693;
  assign n25695 = ~n25589 & ~n25694;
  assign n25696 = n25589 & n25694;
  assign n25697 = ~n25695 & ~n25696;
  assign n25698 = n25579 & ~n25697;
  assign n25699 = ~n25579 & n25697;
  assign n25700 = ~n25698 & ~n25699;
  assign n25701 = n6835 & n21198;
  assign n25702 = n7460 & n21195;
  assign n25703 = n6836 & n23211;
  assign n25704 = n7487 & n21192;
  assign n25705 = ~n25703 & ~n25704;
  assign n25706 = ~n25702 & n25705;
  assign n25707 = ~n25701 & n25706;
  assign n25708 = pi14  & n25707;
  assign n25709 = ~pi14  & ~n25707;
  assign n25710 = ~n25708 & ~n25709;
  assign n25711 = n25700 & n25710;
  assign n25712 = ~n25700 & ~n25710;
  assign n25713 = ~n25711 & ~n25712;
  assign n25714 = ~n25577 & ~n25713;
  assign n25715 = n25577 & n25713;
  assign n25716 = ~n25714 & ~n25715;
  assign n25717 = ~n25574 & ~n25716;
  assign n25718 = n25574 & n25716;
  assign n25719 = ~n25717 & ~n25718;
  assign n25720 = ~n25448 & ~n25452;
  assign n25721 = n25719 & n25720;
  assign n25722 = ~n25719 & ~n25720;
  assign n25723 = ~n25721 & ~n25722;
  assign n25724 = n8474 & n21180;
  assign n25725 = n9238 & n21076;
  assign n25726 = n8468 & n24012;
  assign n25727 = n9265 & n21176;
  assign n25728 = ~n25726 & ~n25727;
  assign n25729 = ~n25725 & n25728;
  assign n25730 = ~n25724 & n25729;
  assign n25731 = pi8  & n25730;
  assign n25732 = ~pi8  & ~n25730;
  assign n25733 = ~n25731 & ~n25732;
  assign n25734 = n25723 & n25733;
  assign n25735 = ~n25723 & ~n25733;
  assign n25736 = ~n25734 & ~n25735;
  assign n25737 = ~n25564 & n25736;
  assign n25738 = n25564 & ~n25736;
  assign n25739 = ~n25737 & ~n25738;
  assign n25740 = ~n25562 & ~n25739;
  assign n25741 = n25562 & n25739;
  assign n25742 = ~n25740 & ~n25741;
  assign n25743 = n25552 & ~n25742;
  assign n25744 = ~n25552 & n25742;
  assign n25745 = ~n25743 & ~n25744;
  assign n25746 = n11288 & n24748;
  assign n25747 = n11894 & n25521;
  assign n25748 = ~n25516 & ~n25519;
  assign n25749 = ~n25501 & ~n25513;
  assign n25750 = n4006 & n12616;
  assign n25751 = ~n24693 & ~n25750;
  assign n25752 = n4002 & ~n13499;
  assign n25753 = ~n25504 & ~n25752;
  assign n25754 = n25751 & n25753;
  assign n25755 = ~pi29  & ~n25754;
  assign n25756 = pi29  & n25754;
  assign n25757 = ~n25755 & ~n25756;
  assign n25758 = n3641 & n12622;
  assign n25759 = n3740 & n12614;
  assign n25760 = n556 & ~n13310;
  assign n25761 = n3961 & n12606;
  assign n25762 = ~n25760 & ~n25761;
  assign n25763 = ~n25759 & n25762;
  assign n25764 = ~n25758 & n25763;
  assign n25765 = ~n25757 & n25764;
  assign n25766 = n25757 & ~n25764;
  assign n25767 = ~n25765 & ~n25766;
  assign n25768 = n486 & n526;
  assign n25769 = n25484 & ~n25768;
  assign n25770 = ~n25484 & n25768;
  assign n25771 = ~n25769 & ~n25770;
  assign n25772 = ~n25485 & n25494;
  assign n25773 = ~n25486 & ~n25772;
  assign n25774 = n25771 & ~n25773;
  assign n25775 = ~n25771 & n25773;
  assign n25776 = ~n25774 & ~n25775;
  assign n25777 = ~n25767 & ~n25776;
  assign n25778 = n25767 & n25776;
  assign n25779 = ~n25777 & ~n25778;
  assign n25780 = ~n25749 & n25779;
  assign n25781 = n25749 & ~n25779;
  assign n25782 = ~n25780 & ~n25781;
  assign n25783 = ~n25748 & n25782;
  assign n25784 = n25748 & ~n25782;
  assign n25785 = ~n25783 & ~n25784;
  assign n25786 = ~n25521 & ~n25785;
  assign n25787 = n25521 & n25785;
  assign n25788 = ~n25786 & ~n25787;
  assign n25789 = ~n25522 & ~n25526;
  assign n25790 = ~n25523 & ~n25789;
  assign n25791 = n25788 & n25790;
  assign n25792 = ~n25788 & ~n25790;
  assign n25793 = ~n25791 & ~n25792;
  assign n25794 = n11289 & n25793;
  assign n25795 = n11908 & n25785;
  assign n25796 = ~n25794 & ~n25795;
  assign n25797 = ~n25747 & n25796;
  assign n25798 = ~n25746 & n25797;
  assign n25799 = pi2  & n25798;
  assign n25800 = ~pi2  & ~n25798;
  assign n25801 = ~n25799 & ~n25800;
  assign n25802 = n25745 & ~n25801;
  assign n25803 = ~n25745 & n25801;
  assign n25804 = ~n25802 & ~n25803;
  assign n25805 = ~n25550 & n25804;
  assign n25806 = n25550 & ~n25804;
  assign n25807 = ~n25805 & ~n25806;
  assign n25808 = n25547 & n25807;
  assign n25809 = ~n25547 & ~n25807;
  assign po1  = ~n25808 & ~n25809;
  assign n25811 = ~n25802 & ~n25805;
  assign n25812 = ~n25740 & ~n25744;
  assign n25813 = n9725 & n24607;
  assign n25814 = n10702 & n24676;
  assign n25815 = n9719 & ~n24754;
  assign n25816 = n11267 & n24748;
  assign n25817 = ~n25815 & ~n25816;
  assign n25818 = ~n25814 & n25817;
  assign n25819 = ~n25813 & n25818;
  assign n25820 = ~pi5  & ~n25819;
  assign n25821 = pi5  & n25819;
  assign n25822 = ~n25820 & ~n25821;
  assign n25823 = n25723 & ~n25733;
  assign n25824 = ~n25564 & ~n25736;
  assign n25825 = ~n25823 & ~n25824;
  assign n25826 = n7654 & n21186;
  assign n25827 = n8091 & n21183;
  assign n25828 = n7648 & n23991;
  assign n25829 = n8120 & n21180;
  assign n25830 = ~n25828 & ~n25829;
  assign n25831 = ~n25827 & n25830;
  assign n25832 = ~n25826 & n25831;
  assign n25833 = ~pi11  & ~n25832;
  assign n25834 = pi11  & n25832;
  assign n25835 = ~n25833 & ~n25834;
  assign n25836 = n25700 & ~n25710;
  assign n25837 = ~n25714 & ~n25836;
  assign n25838 = ~n25695 & ~n25699;
  assign n25839 = n6184 & n21204;
  assign n25840 = n6527 & n21201;
  assign n25841 = n6185 & n22832;
  assign n25842 = n6543 & n21198;
  assign n25843 = ~n25841 & ~n25842;
  assign n25844 = ~n25840 & n25843;
  assign n25845 = ~n25839 & n25844;
  assign n25846 = ~pi17  & ~n25845;
  assign n25847 = pi17  & n25845;
  assign n25848 = ~n25846 & ~n25847;
  assign n25849 = n25678 & ~n25688;
  assign n25850 = ~n25591 & ~n25691;
  assign n25851 = ~n25849 & ~n25850;
  assign n25852 = n5238 & n21222;
  assign n25853 = n71 & n21219;
  assign n25854 = n5239 & n22225;
  assign n25855 = n5326 & n21216;
  assign n25856 = ~n25854 & ~n25855;
  assign n25857 = ~n25853 & n25856;
  assign n25858 = ~n25852 & n25857;
  assign n25859 = ~pi23  & ~n25858;
  assign n25860 = pi23  & n25858;
  assign n25861 = ~n25859 & ~n25860;
  assign n25862 = n25655 & ~n25665;
  assign n25863 = ~n25669 & ~n25862;
  assign n25864 = ~n25650 & ~n25653;
  assign n25865 = n4006 & n21240;
  assign n25866 = n4133 & n21237;
  assign n25867 = n4002 & n21807;
  assign n25868 = n4555 & n21234;
  assign n25869 = ~n25867 & ~n25868;
  assign n25870 = ~n25866 & n25869;
  assign n25871 = ~n25865 & n25870;
  assign n25872 = pi29  & n25871;
  assign n25873 = ~pi29  & ~n25871;
  assign n25874 = ~n25872 & ~n25873;
  assign n25875 = ~n25636 & ~n25643;
  assign n25876 = ~n25647 & ~n25875;
  assign n25877 = n3122 & n4463;
  assign n25878 = n135 & n25877;
  assign n25879 = ~n204 & n25878;
  assign n25880 = n1544 & n13891;
  assign n25881 = n2400 & n25880;
  assign n25882 = n753 & n25881;
  assign n25883 = ~n297 & n25882;
  assign n25884 = ~n535 & n25883;
  assign n25885 = n25879 & n25884;
  assign n25886 = ~n385 & n25885;
  assign n25887 = n2607 & n4486;
  assign n25888 = n7287 & n13128;
  assign n25889 = n777 & n25888;
  assign n25890 = n25887 & n25889;
  assign n25891 = ~n548 & n25890;
  assign n25892 = n1186 & n25891;
  assign n25893 = n25886 & n25892;
  assign n25894 = n3641 & n21249;
  assign n25895 = n556 & n21617;
  assign n25896 = n3961 & n21243;
  assign n25897 = n3740 & n21246;
  assign n25898 = ~n25896 & ~n25897;
  assign n25899 = ~n25895 & n25898;
  assign n25900 = ~n25894 & n25899;
  assign n25901 = ~n25893 & n25900;
  assign n25902 = n25893 & ~n25900;
  assign n25903 = ~n25901 & ~n25902;
  assign n25904 = ~n25876 & ~n25903;
  assign n25905 = n25876 & n25903;
  assign n25906 = ~n25904 & ~n25905;
  assign n25907 = ~n25874 & n25906;
  assign n25908 = n25874 & ~n25906;
  assign n25909 = ~n25907 & ~n25908;
  assign n25910 = ~n25864 & n25909;
  assign n25911 = n25864 & ~n25909;
  assign n25912 = ~n25910 & ~n25911;
  assign n25913 = n4601 & n21231;
  assign n25914 = n4783 & n21228;
  assign n25915 = n4602 & n22001;
  assign n25916 = n4801 & n21225;
  assign n25917 = ~n25915 & ~n25916;
  assign n25918 = ~n25914 & n25917;
  assign n25919 = ~n25913 & n25918;
  assign n25920 = pi26  & n25919;
  assign n25921 = ~pi26  & ~n25919;
  assign n25922 = ~n25920 & ~n25921;
  assign n25923 = n25912 & n25922;
  assign n25924 = ~n25912 & ~n25922;
  assign n25925 = ~n25923 & ~n25924;
  assign n25926 = ~n25863 & ~n25925;
  assign n25927 = n25863 & n25925;
  assign n25928 = ~n25926 & ~n25927;
  assign n25929 = ~n25861 & ~n25928;
  assign n25930 = n25861 & n25928;
  assign n25931 = ~n25929 & ~n25930;
  assign n25932 = ~n25601 & n25671;
  assign n25933 = ~n25677 & ~n25932;
  assign n25934 = n25931 & n25933;
  assign n25935 = ~n25931 & ~n25933;
  assign n25936 = ~n25934 & ~n25935;
  assign n25937 = n5435 & n21213;
  assign n25938 = n6055 & n21210;
  assign n25939 = n5429 & n22363;
  assign n25940 = n6071 & n21207;
  assign n25941 = ~n25939 & ~n25940;
  assign n25942 = ~n25938 & n25941;
  assign n25943 = ~n25937 & n25942;
  assign n25944 = pi20  & n25943;
  assign n25945 = ~pi20  & ~n25943;
  assign n25946 = ~n25944 & ~n25945;
  assign n25947 = n25936 & n25946;
  assign n25948 = ~n25936 & ~n25946;
  assign n25949 = ~n25947 & ~n25948;
  assign n25950 = ~n25851 & n25949;
  assign n25951 = n25851 & ~n25949;
  assign n25952 = ~n25950 & ~n25951;
  assign n25953 = ~n25848 & ~n25952;
  assign n25954 = n25848 & n25952;
  assign n25955 = ~n25953 & ~n25954;
  assign n25956 = n25838 & ~n25955;
  assign n25957 = ~n25838 & n25955;
  assign n25958 = ~n25956 & ~n25957;
  assign n25959 = n6835 & n21195;
  assign n25960 = n7460 & n21192;
  assign n25961 = n6836 & n23399;
  assign n25962 = n7487 & n21189;
  assign n25963 = ~n25961 & ~n25962;
  assign n25964 = ~n25960 & n25963;
  assign n25965 = ~n25959 & n25964;
  assign n25966 = pi14  & n25965;
  assign n25967 = ~pi14  & ~n25965;
  assign n25968 = ~n25966 & ~n25967;
  assign n25969 = n25958 & n25968;
  assign n25970 = ~n25958 & ~n25968;
  assign n25971 = ~n25969 & ~n25970;
  assign n25972 = ~n25837 & ~n25971;
  assign n25973 = n25837 & n25971;
  assign n25974 = ~n25972 & ~n25973;
  assign n25975 = ~n25835 & ~n25974;
  assign n25976 = n25835 & n25974;
  assign n25977 = ~n25975 & ~n25976;
  assign n25978 = ~n25574 & n25716;
  assign n25979 = ~n25722 & ~n25978;
  assign n25980 = n25977 & n25979;
  assign n25981 = ~n25977 & ~n25979;
  assign n25982 = ~n25980 & ~n25981;
  assign n25983 = n8474 & n21076;
  assign n25984 = n9238 & n21176;
  assign n25985 = n8468 & ~n21470;
  assign n25986 = n9265 & n21464;
  assign n25987 = ~n25985 & ~n25986;
  assign n25988 = ~n25984 & n25987;
  assign n25989 = ~n25983 & n25988;
  assign n25990 = pi8  & n25989;
  assign n25991 = ~pi8  & ~n25989;
  assign n25992 = ~n25990 & ~n25991;
  assign n25993 = n25982 & n25992;
  assign n25994 = ~n25982 & ~n25992;
  assign n25995 = ~n25993 & ~n25994;
  assign n25996 = ~n25825 & n25995;
  assign n25997 = n25825 & ~n25995;
  assign n25998 = ~n25996 & ~n25997;
  assign n25999 = ~n25822 & ~n25998;
  assign n26000 = n25822 & n25998;
  assign n26001 = ~n25999 & ~n26000;
  assign n26002 = n25812 & ~n26001;
  assign n26003 = ~n25812 & n26001;
  assign n26004 = ~n26002 & ~n26003;
  assign n26005 = n11288 & n25521;
  assign n26006 = n11894 & n25785;
  assign n26007 = ~n25787 & ~n25791;
  assign n26008 = ~n25780 & ~n25783;
  assign n26009 = ~n25757 & ~n25764;
  assign n26010 = ~n25777 & ~n26009;
  assign n26011 = n4001 & n4005;
  assign n26012 = ~n12608 & ~n26011;
  assign n26013 = pi29  & ~n26012;
  assign n26014 = ~pi29  & n26012;
  assign n26015 = ~n26013 & ~n26014;
  assign n26016 = n12598 & n25768;
  assign n26017 = ~n12598 & ~n25768;
  assign n26018 = ~n26016 & ~n26017;
  assign n26019 = n26015 & n26018;
  assign n26020 = ~n26015 & ~n26018;
  assign n26021 = ~n26019 & ~n26020;
  assign n26022 = n3740 & n12606;
  assign n26023 = n3961 & ~n12608;
  assign n26024 = ~n12611 & n26023;
  assign n26025 = n556 & n12868;
  assign n26026 = n3641 & n12614;
  assign n26027 = ~n26025 & ~n26026;
  assign n26028 = ~n26024 & n26027;
  assign n26029 = ~n26022 & n26028;
  assign n26030 = n26021 & n26029;
  assign n26031 = ~n26021 & ~n26029;
  assign n26032 = ~n26030 & ~n26031;
  assign n26033 = ~n25770 & ~n25773;
  assign n26034 = ~n25769 & ~n26033;
  assign n26035 = ~n26032 & n26034;
  assign n26036 = n26032 & ~n26034;
  assign n26037 = ~n26035 & ~n26036;
  assign n26038 = ~n26010 & n26037;
  assign n26039 = n26010 & ~n26037;
  assign n26040 = ~n26038 & ~n26039;
  assign n26041 = ~n26008 & n26040;
  assign n26042 = n26008 & ~n26040;
  assign n26043 = ~n26041 & ~n26042;
  assign n26044 = ~n25785 & ~n26043;
  assign n26045 = n25785 & n26043;
  assign n26046 = ~n26044 & ~n26045;
  assign n26047 = ~n26007 & n26046;
  assign n26048 = n26007 & ~n26046;
  assign n26049 = ~n26047 & ~n26048;
  assign n26050 = n11289 & n26049;
  assign n26051 = n11908 & n26043;
  assign n26052 = ~n26050 & ~n26051;
  assign n26053 = ~n26006 & n26052;
  assign n26054 = ~n26005 & n26053;
  assign n26055 = pi2  & n26054;
  assign n26056 = ~pi2  & ~n26054;
  assign n26057 = ~n26055 & ~n26056;
  assign n26058 = n26004 & ~n26057;
  assign n26059 = ~n26004 & n26057;
  assign n26060 = ~n26058 & ~n26059;
  assign n26061 = ~n25811 & n26060;
  assign n26062 = n25811 & ~n26060;
  assign n26063 = ~n26061 & ~n26062;
  assign n26064 = n25808 & n26063;
  assign n26065 = ~n25808 & ~n26063;
  assign po2  = ~n26064 & ~n26065;
  assign n26067 = ~n26058 & ~n26061;
  assign n26068 = ~n25999 & ~n26003;
  assign n26069 = n9725 & n24676;
  assign n26070 = n10702 & n24748;
  assign n26071 = n9719 & ~n25529;
  assign n26072 = n11267 & n25521;
  assign n26073 = ~n26071 & ~n26072;
  assign n26074 = ~n26070 & n26073;
  assign n26075 = ~n26069 & n26074;
  assign n26076 = ~pi5  & ~n26075;
  assign n26077 = pi5  & n26075;
  assign n26078 = ~n26076 & ~n26077;
  assign n26079 = n25982 & ~n25992;
  assign n26080 = ~n25825 & ~n25995;
  assign n26081 = ~n26079 & ~n26080;
  assign n26082 = n7654 & n21183;
  assign n26083 = n8091 & n21180;
  assign n26084 = n7648 & n24030;
  assign n26085 = n8120 & n21076;
  assign n26086 = ~n26084 & ~n26085;
  assign n26087 = ~n26083 & n26086;
  assign n26088 = ~n26082 & n26087;
  assign n26089 = ~pi11  & ~n26088;
  assign n26090 = pi11  & n26088;
  assign n26091 = ~n26089 & ~n26090;
  assign n26092 = n25958 & ~n25968;
  assign n26093 = ~n25972 & ~n26092;
  assign n26094 = ~n25953 & ~n25957;
  assign n26095 = n6184 & n21201;
  assign n26096 = n6527 & n21198;
  assign n26097 = n6185 & n21482;
  assign n26098 = n6543 & n21195;
  assign n26099 = ~n26097 & ~n26098;
  assign n26100 = ~n26096 & n26099;
  assign n26101 = ~n26095 & n26100;
  assign n26102 = ~pi17  & ~n26101;
  assign n26103 = pi17  & n26101;
  assign n26104 = ~n26102 & ~n26103;
  assign n26105 = n25936 & ~n25946;
  assign n26106 = ~n25851 & ~n25949;
  assign n26107 = ~n26105 & ~n26106;
  assign n26108 = n5238 & n21219;
  assign n26109 = n71 & n21216;
  assign n26110 = n5239 & n22394;
  assign n26111 = n5326 & n21213;
  assign n26112 = ~n26110 & ~n26111;
  assign n26113 = ~n26109 & n26112;
  assign n26114 = ~n26108 & n26113;
  assign n26115 = ~pi23  & ~n26114;
  assign n26116 = pi23  & n26114;
  assign n26117 = ~n26115 & ~n26116;
  assign n26118 = n25912 & ~n25922;
  assign n26119 = ~n25926 & ~n26118;
  assign n26120 = ~n25907 & ~n25910;
  assign n26121 = n4006 & n21237;
  assign n26122 = n4133 & n21234;
  assign n26123 = n4002 & n21789;
  assign n26124 = n4555 & n21231;
  assign n26125 = ~n26123 & ~n26124;
  assign n26126 = ~n26122 & n26125;
  assign n26127 = ~n26121 & n26126;
  assign n26128 = pi29  & n26127;
  assign n26129 = ~pi29  & ~n26127;
  assign n26130 = ~n26128 & ~n26129;
  assign n26131 = ~n25893 & ~n25900;
  assign n26132 = ~n25904 & ~n26131;
  assign n26133 = n1057 & n1246;
  assign n26134 = n376 & n26133;
  assign n26135 = n3122 & n26134;
  assign n26136 = n2962 & n26135;
  assign n26137 = n896 & n26136;
  assign n26138 = n2469 & n2539;
  assign n26139 = n5506 & n26138;
  assign n26140 = n7311 & n26139;
  assign n26141 = n1482 & n26140;
  assign n26142 = ~n198 & n26141;
  assign n26143 = n26137 & n26142;
  assign n26144 = ~n545 & n26143;
  assign n26145 = n1076 & n4256;
  assign n26146 = n15007 & n26145;
  assign n26147 = n26144 & n26146;
  assign n26148 = n3641 & n21246;
  assign n26149 = n556 & n21604;
  assign n26150 = n3961 & n21240;
  assign n26151 = n3740 & n21243;
  assign n26152 = ~n26150 & ~n26151;
  assign n26153 = ~n26149 & n26152;
  assign n26154 = ~n26148 & n26153;
  assign n26155 = ~n26147 & n26154;
  assign n26156 = n26147 & ~n26154;
  assign n26157 = ~n26155 & ~n26156;
  assign n26158 = ~n26132 & ~n26157;
  assign n26159 = n26132 & n26157;
  assign n26160 = ~n26158 & ~n26159;
  assign n26161 = ~n26130 & n26160;
  assign n26162 = n26130 & ~n26160;
  assign n26163 = ~n26161 & ~n26162;
  assign n26164 = ~n26120 & n26163;
  assign n26165 = n26120 & ~n26163;
  assign n26166 = ~n26164 & ~n26165;
  assign n26167 = n4601 & n21228;
  assign n26168 = n4783 & n21225;
  assign n26169 = n4602 & n21988;
  assign n26170 = n4801 & n21222;
  assign n26171 = ~n26169 & ~n26170;
  assign n26172 = ~n26168 & n26171;
  assign n26173 = ~n26167 & n26172;
  assign n26174 = pi26  & n26173;
  assign n26175 = ~pi26  & ~n26173;
  assign n26176 = ~n26174 & ~n26175;
  assign n26177 = n26166 & n26176;
  assign n26178 = ~n26166 & ~n26176;
  assign n26179 = ~n26177 & ~n26178;
  assign n26180 = ~n26119 & ~n26179;
  assign n26181 = n26119 & n26179;
  assign n26182 = ~n26180 & ~n26181;
  assign n26183 = ~n26117 & ~n26182;
  assign n26184 = n26117 & n26182;
  assign n26185 = ~n26183 & ~n26184;
  assign n26186 = ~n25861 & n25928;
  assign n26187 = ~n25935 & ~n26186;
  assign n26188 = n26185 & n26187;
  assign n26189 = ~n26185 & ~n26187;
  assign n26190 = ~n26188 & ~n26189;
  assign n26191 = n5435 & n21210;
  assign n26192 = n6055 & n21207;
  assign n26193 = n5429 & n22810;
  assign n26194 = n6071 & n21204;
  assign n26195 = ~n26193 & ~n26194;
  assign n26196 = ~n26192 & n26195;
  assign n26197 = ~n26191 & n26196;
  assign n26198 = pi20  & n26197;
  assign n26199 = ~pi20  & ~n26197;
  assign n26200 = ~n26198 & ~n26199;
  assign n26201 = n26190 & n26200;
  assign n26202 = ~n26190 & ~n26200;
  assign n26203 = ~n26201 & ~n26202;
  assign n26204 = ~n26107 & n26203;
  assign n26205 = n26107 & ~n26203;
  assign n26206 = ~n26204 & ~n26205;
  assign n26207 = ~n26104 & ~n26206;
  assign n26208 = n26104 & n26206;
  assign n26209 = ~n26207 & ~n26208;
  assign n26210 = n26094 & ~n26209;
  assign n26211 = ~n26094 & n26209;
  assign n26212 = ~n26210 & ~n26211;
  assign n26213 = n6835 & n21192;
  assign n26214 = n7460 & n21189;
  assign n26215 = n6836 & n23384;
  assign n26216 = n7487 & n21186;
  assign n26217 = ~n26215 & ~n26216;
  assign n26218 = ~n26214 & n26217;
  assign n26219 = ~n26213 & n26218;
  assign n26220 = pi14  & n26219;
  assign n26221 = ~pi14  & ~n26219;
  assign n26222 = ~n26220 & ~n26221;
  assign n26223 = n26212 & n26222;
  assign n26224 = ~n26212 & ~n26222;
  assign n26225 = ~n26223 & ~n26224;
  assign n26226 = ~n26093 & ~n26225;
  assign n26227 = n26093 & n26225;
  assign n26228 = ~n26226 & ~n26227;
  assign n26229 = ~n26091 & ~n26228;
  assign n26230 = n26091 & n26228;
  assign n26231 = ~n26229 & ~n26230;
  assign n26232 = ~n25835 & n25974;
  assign n26233 = ~n25981 & ~n26232;
  assign n26234 = n26231 & n26233;
  assign n26235 = ~n26231 & ~n26233;
  assign n26236 = ~n26234 & ~n26235;
  assign n26237 = n8474 & n21176;
  assign n26238 = n9238 & n21464;
  assign n26239 = n8468 & n24782;
  assign n26240 = n9265 & n24607;
  assign n26241 = ~n26239 & ~n26240;
  assign n26242 = ~n26238 & n26241;
  assign n26243 = ~n26237 & n26242;
  assign n26244 = pi8  & n26243;
  assign n26245 = ~pi8  & ~n26243;
  assign n26246 = ~n26244 & ~n26245;
  assign n26247 = n26236 & n26246;
  assign n26248 = ~n26236 & ~n26246;
  assign n26249 = ~n26247 & ~n26248;
  assign n26250 = ~n26081 & n26249;
  assign n26251 = n26081 & ~n26249;
  assign n26252 = ~n26250 & ~n26251;
  assign n26253 = ~n26078 & ~n26252;
  assign n26254 = n26078 & n26252;
  assign n26255 = ~n26253 & ~n26254;
  assign n26256 = n26068 & ~n26255;
  assign n26257 = ~n26068 & n26255;
  assign n26258 = ~n26256 & ~n26257;
  assign n26259 = n11288 & n25785;
  assign n26260 = n11894 & n26043;
  assign n26261 = ~n26045 & ~n26047;
  assign n26262 = n26021 & ~n26029;
  assign n26263 = ~n26035 & ~n26262;
  assign n26264 = ~n26017 & ~n26019;
  assign n26265 = n553 & ~n26264;
  assign n26266 = ~n553 & n26264;
  assign n26267 = ~n26265 & ~n26266;
  assign n26268 = n3641 & n12606;
  assign n26269 = n3740 & ~n12608;
  assign n26270 = ~n12611 & n26269;
  assign n26271 = n556 & ~n13483;
  assign n26272 = ~n26023 & ~n26271;
  assign n26273 = ~n26270 & n26272;
  assign n26274 = ~n26268 & n26273;
  assign n26275 = n26267 & ~n26274;
  assign n26276 = ~n26267 & n26274;
  assign n26277 = ~n26275 & ~n26276;
  assign n26278 = n26263 & ~n26277;
  assign n26279 = ~n26263 & n26277;
  assign n26280 = ~n26278 & ~n26279;
  assign n26281 = ~n26038 & ~n26041;
  assign n26282 = ~n26280 & n26281;
  assign n26283 = n26280 & ~n26281;
  assign n26284 = ~n26282 & ~n26283;
  assign n26285 = n26043 & n26284;
  assign n26286 = ~n26043 & ~n26284;
  assign n26287 = ~n26285 & ~n26286;
  assign n26288 = n26261 & n26287;
  assign n26289 = ~n26261 & ~n26287;
  assign n26290 = ~n26288 & ~n26289;
  assign n26291 = n11289 & ~n26290;
  assign n26292 = n11908 & n26284;
  assign n26293 = ~n26291 & ~n26292;
  assign n26294 = ~n26260 & n26293;
  assign n26295 = ~n26259 & n26294;
  assign n26296 = pi2  & n26295;
  assign n26297 = ~pi2  & ~n26295;
  assign n26298 = ~n26296 & ~n26297;
  assign n26299 = n26258 & ~n26298;
  assign n26300 = ~n26258 & n26298;
  assign n26301 = ~n26299 & ~n26300;
  assign n26302 = ~n26067 & n26301;
  assign n26303 = n26067 & ~n26301;
  assign n26304 = ~n26302 & ~n26303;
  assign n26305 = n26064 & n26304;
  assign n26306 = ~n26064 & ~n26304;
  assign po3  = ~n26305 & ~n26306;
  assign n26308 = ~n26299 & ~n26302;
  assign n26309 = ~n26253 & ~n26257;
  assign n26310 = n9725 & n24748;
  assign n26311 = n10702 & n25521;
  assign n26312 = n9719 & n25793;
  assign n26313 = n11267 & n25785;
  assign n26314 = ~n26312 & ~n26313;
  assign n26315 = ~n26311 & n26314;
  assign n26316 = ~n26310 & n26315;
  assign n26317 = ~pi5  & ~n26316;
  assign n26318 = pi5  & n26316;
  assign n26319 = ~n26317 & ~n26318;
  assign n26320 = n26236 & ~n26246;
  assign n26321 = ~n26081 & ~n26249;
  assign n26322 = ~n26320 & ~n26321;
  assign n26323 = n7654 & n21180;
  assign n26324 = n8091 & n21076;
  assign n26325 = n7648 & n24012;
  assign n26326 = n8120 & n21176;
  assign n26327 = ~n26325 & ~n26326;
  assign n26328 = ~n26324 & n26327;
  assign n26329 = ~n26323 & n26328;
  assign n26330 = ~pi11  & ~n26329;
  assign n26331 = pi11  & n26329;
  assign n26332 = ~n26330 & ~n26331;
  assign n26333 = n26212 & ~n26222;
  assign n26334 = ~n26226 & ~n26333;
  assign n26335 = ~n26207 & ~n26211;
  assign n26336 = n6184 & n21198;
  assign n26337 = n6527 & n21195;
  assign n26338 = n6185 & n23211;
  assign n26339 = n6543 & n21192;
  assign n26340 = ~n26338 & ~n26339;
  assign n26341 = ~n26337 & n26340;
  assign n26342 = ~n26336 & n26341;
  assign n26343 = ~pi17  & ~n26342;
  assign n26344 = pi17  & n26342;
  assign n26345 = ~n26343 & ~n26344;
  assign n26346 = n26190 & ~n26200;
  assign n26347 = ~n26107 & ~n26203;
  assign n26348 = ~n26346 & ~n26347;
  assign n26349 = n5238 & n21216;
  assign n26350 = n71 & n21213;
  assign n26351 = n5239 & n22376;
  assign n26352 = n5326 & n21210;
  assign n26353 = ~n26351 & ~n26352;
  assign n26354 = ~n26350 & n26353;
  assign n26355 = ~n26349 & n26354;
  assign n26356 = ~pi23  & ~n26355;
  assign n26357 = pi23  & n26355;
  assign n26358 = ~n26356 & ~n26357;
  assign n26359 = n26166 & ~n26176;
  assign n26360 = ~n26180 & ~n26359;
  assign n26361 = ~n26161 & ~n26164;
  assign n26362 = n4006 & n21234;
  assign n26363 = n4133 & n21231;
  assign n26364 = n4002 & n21494;
  assign n26365 = n4555 & n21228;
  assign n26366 = ~n26364 & ~n26365;
  assign n26367 = ~n26363 & n26366;
  assign n26368 = ~n26362 & n26367;
  assign n26369 = pi29  & n26368;
  assign n26370 = ~pi29  & ~n26368;
  assign n26371 = ~n26369 & ~n26370;
  assign n26372 = ~n26147 & ~n26154;
  assign n26373 = ~n26158 & ~n26372;
  assign n26374 = n881 & n2153;
  assign n26375 = n2529 & n26374;
  assign n26376 = n4398 & n26375;
  assign n26377 = n1388 & n26376;
  assign n26378 = ~n297 & n26377;
  assign n26379 = ~n232 & n1024;
  assign n26380 = ~n363 & n26379;
  assign n26381 = ~n430 & n1253;
  assign n26382 = ~n533 & n26381;
  assign n26383 = n26380 & n26382;
  assign n26384 = ~n334 & n2409;
  assign n26385 = ~n610 & n26384;
  assign n26386 = ~n204 & n2842;
  assign n26387 = ~n473 & n26386;
  assign n26388 = n26385 & n26387;
  assign n26389 = n26383 & n26388;
  assign n26390 = n2837 & n26389;
  assign n26391 = n1109 & n26390;
  assign n26392 = ~n670 & n26391;
  assign n26393 = n26378 & n26392;
  assign n26394 = n184 & n5038;
  assign n26395 = n1091 & n26394;
  assign n26396 = n230 & n26395;
  assign n26397 = ~n535 & n26396;
  assign n26398 = n1925 & n2784;
  assign n26399 = ~n590 & n26398;
  assign n26400 = ~n259 & n26399;
  assign n26401 = n26397 & n26400;
  assign n26402 = n26393 & n26401;
  assign n26403 = n3641 & n21243;
  assign n26404 = n556 & n21768;
  assign n26405 = n3961 & n21237;
  assign n26406 = n3740 & n21240;
  assign n26407 = ~n26405 & ~n26406;
  assign n26408 = ~n26404 & n26407;
  assign n26409 = ~n26403 & n26408;
  assign n26410 = ~n26402 & n26409;
  assign n26411 = n26402 & ~n26409;
  assign n26412 = ~n26410 & ~n26411;
  assign n26413 = ~n26373 & ~n26412;
  assign n26414 = n26373 & n26412;
  assign n26415 = ~n26413 & ~n26414;
  assign n26416 = ~n26371 & n26415;
  assign n26417 = n26371 & ~n26415;
  assign n26418 = ~n26416 & ~n26417;
  assign n26419 = ~n26361 & n26418;
  assign n26420 = n26361 & ~n26418;
  assign n26421 = ~n26419 & ~n26420;
  assign n26422 = n4601 & n21225;
  assign n26423 = n4783 & n21222;
  assign n26424 = n4602 & n21973;
  assign n26425 = n4801 & n21219;
  assign n26426 = ~n26424 & ~n26425;
  assign n26427 = ~n26423 & n26426;
  assign n26428 = ~n26422 & n26427;
  assign n26429 = pi26  & n26428;
  assign n26430 = ~pi26  & ~n26428;
  assign n26431 = ~n26429 & ~n26430;
  assign n26432 = n26421 & n26431;
  assign n26433 = ~n26421 & ~n26431;
  assign n26434 = ~n26432 & ~n26433;
  assign n26435 = ~n26360 & ~n26434;
  assign n26436 = n26360 & n26434;
  assign n26437 = ~n26435 & ~n26436;
  assign n26438 = ~n26358 & ~n26437;
  assign n26439 = n26358 & n26437;
  assign n26440 = ~n26438 & ~n26439;
  assign n26441 = ~n26117 & n26182;
  assign n26442 = ~n26189 & ~n26441;
  assign n26443 = n26440 & n26442;
  assign n26444 = ~n26440 & ~n26442;
  assign n26445 = ~n26443 & ~n26444;
  assign n26446 = n5435 & n21207;
  assign n26447 = n6055 & n21204;
  assign n26448 = n5429 & n22852;
  assign n26449 = n6071 & n21201;
  assign n26450 = ~n26448 & ~n26449;
  assign n26451 = ~n26447 & n26450;
  assign n26452 = ~n26446 & n26451;
  assign n26453 = pi20  & n26452;
  assign n26454 = ~pi20  & ~n26452;
  assign n26455 = ~n26453 & ~n26454;
  assign n26456 = n26445 & n26455;
  assign n26457 = ~n26445 & ~n26455;
  assign n26458 = ~n26456 & ~n26457;
  assign n26459 = ~n26348 & n26458;
  assign n26460 = n26348 & ~n26458;
  assign n26461 = ~n26459 & ~n26460;
  assign n26462 = ~n26345 & ~n26461;
  assign n26463 = n26345 & n26461;
  assign n26464 = ~n26462 & ~n26463;
  assign n26465 = n26335 & ~n26464;
  assign n26466 = ~n26335 & n26464;
  assign n26467 = ~n26465 & ~n26466;
  assign n26468 = n6835 & n21189;
  assign n26469 = n7460 & n21186;
  assign n26470 = n6836 & n23369;
  assign n26471 = n7487 & n21183;
  assign n26472 = ~n26470 & ~n26471;
  assign n26473 = ~n26469 & n26472;
  assign n26474 = ~n26468 & n26473;
  assign n26475 = pi14  & n26474;
  assign n26476 = ~pi14  & ~n26474;
  assign n26477 = ~n26475 & ~n26476;
  assign n26478 = n26467 & n26477;
  assign n26479 = ~n26467 & ~n26477;
  assign n26480 = ~n26478 & ~n26479;
  assign n26481 = ~n26334 & ~n26480;
  assign n26482 = n26334 & n26480;
  assign n26483 = ~n26481 & ~n26482;
  assign n26484 = ~n26332 & ~n26483;
  assign n26485 = n26332 & n26483;
  assign n26486 = ~n26484 & ~n26485;
  assign n26487 = ~n26091 & n26228;
  assign n26488 = ~n26235 & ~n26487;
  assign n26489 = n26486 & n26488;
  assign n26490 = ~n26486 & ~n26488;
  assign n26491 = ~n26489 & ~n26490;
  assign n26492 = n8474 & n21464;
  assign n26493 = n9238 & n24607;
  assign n26494 = n8468 & n24770;
  assign n26495 = n9265 & n24676;
  assign n26496 = ~n26494 & ~n26495;
  assign n26497 = ~n26493 & n26496;
  assign n26498 = ~n26492 & n26497;
  assign n26499 = pi8  & n26498;
  assign n26500 = ~pi8  & ~n26498;
  assign n26501 = ~n26499 & ~n26500;
  assign n26502 = n26491 & n26501;
  assign n26503 = ~n26491 & ~n26501;
  assign n26504 = ~n26502 & ~n26503;
  assign n26505 = ~n26322 & n26504;
  assign n26506 = n26322 & ~n26504;
  assign n26507 = ~n26505 & ~n26506;
  assign n26508 = ~n26319 & ~n26507;
  assign n26509 = n26319 & n26507;
  assign n26510 = ~n26508 & ~n26509;
  assign n26511 = n26309 & ~n26510;
  assign n26512 = ~n26309 & n26510;
  assign n26513 = ~n26511 & ~n26512;
  assign n26514 = n11288 & n26043;
  assign n26515 = n11894 & n26284;
  assign n26516 = n3641 & n12616;
  assign n26517 = ~n26023 & ~n26516;
  assign n26518 = n556 & ~n13499;
  assign n26519 = ~n26269 & ~n26518;
  assign n26520 = n26517 & n26519;
  assign n26521 = n553 & n26520;
  assign n26522 = ~n553 & ~n26520;
  assign n26523 = ~n26521 & ~n26522;
  assign n26524 = ~n26265 & n26274;
  assign n26525 = ~n26266 & ~n26524;
  assign n26526 = n26523 & ~n26525;
  assign n26527 = ~n26523 & n26525;
  assign n26528 = ~n26526 & ~n26527;
  assign n26529 = ~n26279 & ~n26283;
  assign n26530 = ~n26528 & n26529;
  assign n26531 = n26528 & ~n26529;
  assign n26532 = ~n26530 & ~n26531;
  assign n26533 = ~n26284 & ~n26532;
  assign n26534 = n26284 & n26532;
  assign n26535 = ~n26533 & ~n26534;
  assign n26536 = n26261 & ~n26285;
  assign n26537 = ~n26286 & ~n26536;
  assign n26538 = n26535 & n26537;
  assign n26539 = ~n26535 & ~n26537;
  assign n26540 = ~n26538 & ~n26539;
  assign n26541 = n11289 & n26540;
  assign n26542 = n11908 & n26532;
  assign n26543 = ~n26541 & ~n26542;
  assign n26544 = ~n26515 & n26543;
  assign n26545 = ~n26514 & n26544;
  assign n26546 = pi2  & n26545;
  assign n26547 = ~pi2  & ~n26545;
  assign n26548 = ~n26546 & ~n26547;
  assign n26549 = n26513 & ~n26548;
  assign n26550 = ~n26513 & n26548;
  assign n26551 = ~n26549 & ~n26550;
  assign n26552 = ~n26308 & n26551;
  assign n26553 = n26308 & ~n26551;
  assign n26554 = ~n26552 & ~n26553;
  assign n26555 = n26305 & n26554;
  assign n26556 = ~n26305 & ~n26554;
  assign po4  = ~n26555 & ~n26556;
  assign n26558 = ~n26549 & ~n26552;
  assign n26559 = ~n26508 & ~n26512;
  assign n26560 = n9725 & n25521;
  assign n26561 = n10702 & n25785;
  assign n26562 = n9719 & n26049;
  assign n26563 = n11267 & n26043;
  assign n26564 = ~n26562 & ~n26563;
  assign n26565 = ~n26561 & n26564;
  assign n26566 = ~n26560 & n26565;
  assign n26567 = ~pi5  & ~n26566;
  assign n26568 = pi5  & n26566;
  assign n26569 = ~n26567 & ~n26568;
  assign n26570 = n26491 & ~n26501;
  assign n26571 = ~n26322 & ~n26504;
  assign n26572 = ~n26570 & ~n26571;
  assign n26573 = n7654 & n21076;
  assign n26574 = n8091 & n21176;
  assign n26575 = n7648 & ~n21470;
  assign n26576 = n8120 & n21464;
  assign n26577 = ~n26575 & ~n26576;
  assign n26578 = ~n26574 & n26577;
  assign n26579 = ~n26573 & n26578;
  assign n26580 = ~pi11  & ~n26579;
  assign n26581 = pi11  & n26579;
  assign n26582 = ~n26580 & ~n26581;
  assign n26583 = n26467 & ~n26477;
  assign n26584 = ~n26481 & ~n26583;
  assign n26585 = ~n26462 & ~n26466;
  assign n26586 = n6184 & n21195;
  assign n26587 = n6527 & n21192;
  assign n26588 = n6185 & n23399;
  assign n26589 = n6543 & n21189;
  assign n26590 = ~n26588 & ~n26589;
  assign n26591 = ~n26587 & n26590;
  assign n26592 = ~n26586 & n26591;
  assign n26593 = ~pi17  & ~n26592;
  assign n26594 = pi17  & n26592;
  assign n26595 = ~n26593 & ~n26594;
  assign n26596 = n26445 & ~n26455;
  assign n26597 = ~n26348 & ~n26458;
  assign n26598 = ~n26596 & ~n26597;
  assign n26599 = n5238 & n21213;
  assign n26600 = n71 & n21210;
  assign n26601 = n5239 & n22363;
  assign n26602 = n5326 & n21207;
  assign n26603 = ~n26601 & ~n26602;
  assign n26604 = ~n26600 & n26603;
  assign n26605 = ~n26599 & n26604;
  assign n26606 = ~pi23  & ~n26605;
  assign n26607 = pi23  & n26605;
  assign n26608 = ~n26606 & ~n26607;
  assign n26609 = n26421 & ~n26431;
  assign n26610 = ~n26435 & ~n26609;
  assign n26611 = ~n26416 & ~n26419;
  assign n26612 = n4006 & n21231;
  assign n26613 = n4133 & n21228;
  assign n26614 = n4002 & n22001;
  assign n26615 = n4555 & n21225;
  assign n26616 = ~n26614 & ~n26615;
  assign n26617 = ~n26613 & n26616;
  assign n26618 = ~n26612 & n26617;
  assign n26619 = pi29  & n26618;
  assign n26620 = ~pi29  & ~n26618;
  assign n26621 = ~n26619 & ~n26620;
  assign n26622 = ~n26402 & ~n26409;
  assign n26623 = ~n26413 & ~n26622;
  assign n26624 = n1058 & n4229;
  assign n26625 = n1576 & n26624;
  assign n26626 = n519 & n26625;
  assign n26627 = ~n173 & n26626;
  assign n26628 = ~n672 & n26627;
  assign n26629 = n1081 & n4200;
  assign n26630 = ~n81 & n26629;
  assign n26631 = ~n474 & n26630;
  assign n26632 = ~n414 & n26631;
  assign n26633 = n26628 & n26632;
  assign n26634 = ~n613 & n15231;
  assign n26635 = ~n238 & n26634;
  assign n26636 = ~n610 & n26635;
  assign n26637 = ~n163 & n5934;
  assign n26638 = ~n441 & n26637;
  assign n26639 = ~n638 & n26638;
  assign n26640 = n26636 & n26639;
  assign n26641 = n26633 & n26640;
  assign n26642 = n3641 & n21240;
  assign n26643 = n556 & n21807;
  assign n26644 = n3961 & n21234;
  assign n26645 = n3740 & n21237;
  assign n26646 = ~n26644 & ~n26645;
  assign n26647 = ~n26643 & n26646;
  assign n26648 = ~n26642 & n26647;
  assign n26649 = ~n26641 & n26648;
  assign n26650 = n26641 & ~n26648;
  assign n26651 = ~n26649 & ~n26650;
  assign n26652 = ~n26623 & ~n26651;
  assign n26653 = n26623 & n26651;
  assign n26654 = ~n26652 & ~n26653;
  assign n26655 = ~n26621 & n26654;
  assign n26656 = n26621 & ~n26654;
  assign n26657 = ~n26655 & ~n26656;
  assign n26658 = ~n26611 & n26657;
  assign n26659 = n26611 & ~n26657;
  assign n26660 = ~n26658 & ~n26659;
  assign n26661 = n4601 & n21222;
  assign n26662 = n4783 & n21219;
  assign n26663 = n4602 & n22225;
  assign n26664 = n4801 & n21216;
  assign n26665 = ~n26663 & ~n26664;
  assign n26666 = ~n26662 & n26665;
  assign n26667 = ~n26661 & n26666;
  assign n26668 = pi26  & n26667;
  assign n26669 = ~pi26  & ~n26667;
  assign n26670 = ~n26668 & ~n26669;
  assign n26671 = n26660 & n26670;
  assign n26672 = ~n26660 & ~n26670;
  assign n26673 = ~n26671 & ~n26672;
  assign n26674 = ~n26610 & ~n26673;
  assign n26675 = n26610 & n26673;
  assign n26676 = ~n26674 & ~n26675;
  assign n26677 = ~n26608 & ~n26676;
  assign n26678 = n26608 & n26676;
  assign n26679 = ~n26677 & ~n26678;
  assign n26680 = ~n26358 & n26437;
  assign n26681 = ~n26444 & ~n26680;
  assign n26682 = n26679 & n26681;
  assign n26683 = ~n26679 & ~n26681;
  assign n26684 = ~n26682 & ~n26683;
  assign n26685 = n5435 & n21204;
  assign n26686 = n6055 & n21201;
  assign n26687 = n5429 & n22832;
  assign n26688 = n6071 & n21198;
  assign n26689 = ~n26687 & ~n26688;
  assign n26690 = ~n26686 & n26689;
  assign n26691 = ~n26685 & n26690;
  assign n26692 = pi20  & n26691;
  assign n26693 = ~pi20  & ~n26691;
  assign n26694 = ~n26692 & ~n26693;
  assign n26695 = n26684 & n26694;
  assign n26696 = ~n26684 & ~n26694;
  assign n26697 = ~n26695 & ~n26696;
  assign n26698 = ~n26598 & n26697;
  assign n26699 = n26598 & ~n26697;
  assign n26700 = ~n26698 & ~n26699;
  assign n26701 = ~n26595 & ~n26700;
  assign n26702 = n26595 & n26700;
  assign n26703 = ~n26701 & ~n26702;
  assign n26704 = n26585 & ~n26703;
  assign n26705 = ~n26585 & n26703;
  assign n26706 = ~n26704 & ~n26705;
  assign n26707 = n6835 & n21186;
  assign n26708 = n7460 & n21183;
  assign n26709 = n6836 & n23991;
  assign n26710 = n7487 & n21180;
  assign n26711 = ~n26709 & ~n26710;
  assign n26712 = ~n26708 & n26711;
  assign n26713 = ~n26707 & n26712;
  assign n26714 = pi14  & n26713;
  assign n26715 = ~pi14  & ~n26713;
  assign n26716 = ~n26714 & ~n26715;
  assign n26717 = n26706 & n26716;
  assign n26718 = ~n26706 & ~n26716;
  assign n26719 = ~n26717 & ~n26718;
  assign n26720 = ~n26584 & ~n26719;
  assign n26721 = n26584 & n26719;
  assign n26722 = ~n26720 & ~n26721;
  assign n26723 = ~n26582 & ~n26722;
  assign n26724 = n26582 & n26722;
  assign n26725 = ~n26723 & ~n26724;
  assign n26726 = ~n26332 & n26483;
  assign n26727 = ~n26490 & ~n26726;
  assign n26728 = n26725 & n26727;
  assign n26729 = ~n26725 & ~n26727;
  assign n26730 = ~n26728 & ~n26729;
  assign n26731 = n8474 & n24607;
  assign n26732 = n9238 & n24676;
  assign n26733 = n8468 & ~n24754;
  assign n26734 = n9265 & n24748;
  assign n26735 = ~n26733 & ~n26734;
  assign n26736 = ~n26732 & n26735;
  assign n26737 = ~n26731 & n26736;
  assign n26738 = pi8  & n26737;
  assign n26739 = ~pi8  & ~n26737;
  assign n26740 = ~n26738 & ~n26739;
  assign n26741 = n26730 & n26740;
  assign n26742 = ~n26730 & ~n26740;
  assign n26743 = ~n26741 & ~n26742;
  assign n26744 = ~n26572 & n26743;
  assign n26745 = n26572 & ~n26743;
  assign n26746 = ~n26744 & ~n26745;
  assign n26747 = ~n26569 & ~n26746;
  assign n26748 = n26569 & n26746;
  assign n26749 = ~n26747 & ~n26748;
  assign n26750 = n26559 & ~n26749;
  assign n26751 = ~n26559 & n26749;
  assign n26752 = ~n26750 & ~n26751;
  assign n26753 = n11288 & n26284;
  assign n26754 = n11894 & n26532;
  assign n26755 = ~n26534 & ~n26538;
  assign n26756 = ~n26527 & ~n26531;
  assign n26757 = ~pi31  & n95;
  assign n26758 = ~n12608 & ~n26757;
  assign n26759 = n26521 & ~n26758;
  assign n26760 = ~n26521 & n26758;
  assign n26761 = ~n26759 & ~n26760;
  assign n26762 = n26756 & n26761;
  assign n26763 = ~n26756 & ~n26761;
  assign n26764 = ~n26762 & ~n26763;
  assign n26765 = n26532 & n26764;
  assign n26766 = ~n26532 & ~n26764;
  assign n26767 = ~n26765 & ~n26766;
  assign n26768 = n26755 & n26767;
  assign n26769 = ~n26755 & ~n26767;
  assign n26770 = ~n26768 & ~n26769;
  assign n26771 = n11289 & ~n26770;
  assign n26772 = n11908 & n26764;
  assign n26773 = ~n26771 & ~n26772;
  assign n26774 = ~n26754 & n26773;
  assign n26775 = ~n26753 & n26774;
  assign n26776 = pi2  & n26775;
  assign n26777 = ~pi2  & ~n26775;
  assign n26778 = ~n26776 & ~n26777;
  assign n26779 = n26752 & ~n26778;
  assign n26780 = ~n26752 & n26778;
  assign n26781 = ~n26779 & ~n26780;
  assign n26782 = ~n26558 & n26781;
  assign n26783 = n26558 & ~n26781;
  assign n26784 = ~n26782 & ~n26783;
  assign n26785 = n26555 & n26784;
  assign n26786 = ~n26555 & ~n26784;
  assign po5  = ~n26785 & ~n26786;
  assign n26788 = ~n26747 & ~n26751;
  assign n26789 = n9725 & n25785;
  assign n26790 = n10702 & n26043;
  assign n26791 = n9719 & ~n26290;
  assign n26792 = n11267 & n26284;
  assign n26793 = ~n26791 & ~n26792;
  assign n26794 = ~n26790 & n26793;
  assign n26795 = ~n26789 & n26794;
  assign n26796 = ~pi5  & ~n26795;
  assign n26797 = pi5  & n26795;
  assign n26798 = ~n26796 & ~n26797;
  assign n26799 = n26730 & ~n26740;
  assign n26800 = ~n26572 & ~n26743;
  assign n26801 = ~n26799 & ~n26800;
  assign n26802 = n7654 & n21176;
  assign n26803 = n8091 & n21464;
  assign n26804 = n7648 & n24782;
  assign n26805 = n8120 & n24607;
  assign n26806 = ~n26804 & ~n26805;
  assign n26807 = ~n26803 & n26806;
  assign n26808 = ~n26802 & n26807;
  assign n26809 = ~pi11  & ~n26808;
  assign n26810 = pi11  & n26808;
  assign n26811 = ~n26809 & ~n26810;
  assign n26812 = n26706 & ~n26716;
  assign n26813 = ~n26720 & ~n26812;
  assign n26814 = n6184 & n21192;
  assign n26815 = n6527 & n21189;
  assign n26816 = n6185 & n23384;
  assign n26817 = n6543 & n21186;
  assign n26818 = ~n26816 & ~n26817;
  assign n26819 = ~n26815 & n26818;
  assign n26820 = ~n26814 & n26819;
  assign n26821 = ~pi17  & ~n26820;
  assign n26822 = pi17  & n26820;
  assign n26823 = ~n26821 & ~n26822;
  assign n26824 = n26684 & ~n26694;
  assign n26825 = ~n26598 & ~n26697;
  assign n26826 = ~n26824 & ~n26825;
  assign n26827 = n5238 & n21210;
  assign n26828 = n71 & n21207;
  assign n26829 = n5239 & n22810;
  assign n26830 = n5326 & n21204;
  assign n26831 = ~n26829 & ~n26830;
  assign n26832 = ~n26828 & n26831;
  assign n26833 = ~n26827 & n26832;
  assign n26834 = ~pi23  & ~n26833;
  assign n26835 = pi23  & n26833;
  assign n26836 = ~n26834 & ~n26835;
  assign n26837 = n26660 & ~n26670;
  assign n26838 = ~n26674 & ~n26837;
  assign n26839 = ~n26655 & ~n26658;
  assign n26840 = n4006 & n21228;
  assign n26841 = n4133 & n21225;
  assign n26842 = n4002 & n21988;
  assign n26843 = n4555 & n21222;
  assign n26844 = ~n26842 & ~n26843;
  assign n26845 = ~n26841 & n26844;
  assign n26846 = ~n26840 & n26845;
  assign n26847 = pi29  & n26846;
  assign n26848 = ~pi29  & ~n26846;
  assign n26849 = ~n26847 & ~n26848;
  assign n26850 = ~n26641 & ~n26648;
  assign n26851 = ~n26652 & ~n26850;
  assign n26852 = n881 & n14333;
  assign n26853 = n1478 & n26852;
  assign n26854 = n1111 & n26134;
  assign n26855 = n1402 & n26854;
  assign n26856 = n3157 & n26855;
  assign n26857 = n26853 & n26856;
  assign n26858 = n1343 & n26857;
  assign n26859 = ~n298 & n26858;
  assign n26860 = ~n464 & n26859;
  assign n26861 = ~n458 & n2281;
  assign n26862 = n845 & n26861;
  assign n26863 = ~n441 & n26862;
  assign n26864 = n2502 & n3270;
  assign n26865 = n26863 & n26864;
  assign n26866 = n5712 & n13895;
  assign n26867 = n230 & n26866;
  assign n26868 = n26865 & n26867;
  assign n26869 = ~n398 & n26868;
  assign n26870 = ~n349 & n26869;
  assign n26871 = n26860 & n26870;
  assign n26872 = ~n473 & n26871;
  assign n26873 = ~n518 & n901;
  assign n26874 = ~n260 & n26873;
  assign n26875 = ~n218 & n26874;
  assign n26876 = n26872 & n26875;
  assign n26877 = n3641 & n21237;
  assign n26878 = n556 & n21789;
  assign n26879 = n3961 & n21231;
  assign n26880 = n3740 & n21234;
  assign n26881 = ~n26879 & ~n26880;
  assign n26882 = ~n26878 & n26881;
  assign n26883 = ~n26877 & n26882;
  assign n26884 = ~n26876 & n26883;
  assign n26885 = n26876 & ~n26883;
  assign n26886 = ~n26884 & ~n26885;
  assign n26887 = ~n26851 & ~n26886;
  assign n26888 = n26851 & n26886;
  assign n26889 = ~n26887 & ~n26888;
  assign n26890 = ~n26849 & n26889;
  assign n26891 = n26849 & ~n26889;
  assign n26892 = ~n26890 & ~n26891;
  assign n26893 = ~n26839 & n26892;
  assign n26894 = n26839 & ~n26892;
  assign n26895 = ~n26893 & ~n26894;
  assign n26896 = n4601 & n21219;
  assign n26897 = n4783 & n21216;
  assign n26898 = n4602 & n22394;
  assign n26899 = n4801 & n21213;
  assign n26900 = ~n26898 & ~n26899;
  assign n26901 = ~n26897 & n26900;
  assign n26902 = ~n26896 & n26901;
  assign n26903 = pi26  & n26902;
  assign n26904 = ~pi26  & ~n26902;
  assign n26905 = ~n26903 & ~n26904;
  assign n26906 = n26895 & ~n26905;
  assign n26907 = ~n26895 & n26905;
  assign n26908 = ~n26906 & ~n26907;
  assign n26909 = ~n26838 & n26908;
  assign n26910 = n26838 & ~n26908;
  assign n26911 = ~n26909 & ~n26910;
  assign n26912 = ~n26836 & ~n26911;
  assign n26913 = n26836 & n26911;
  assign n26914 = ~n26912 & ~n26913;
  assign n26915 = ~n26608 & n26676;
  assign n26916 = ~n26683 & ~n26915;
  assign n26917 = n26914 & n26916;
  assign n26918 = ~n26914 & ~n26916;
  assign n26919 = ~n26917 & ~n26918;
  assign n26920 = n5435 & n21201;
  assign n26921 = n6055 & n21198;
  assign n26922 = n5429 & n21482;
  assign n26923 = n6071 & n21195;
  assign n26924 = ~n26922 & ~n26923;
  assign n26925 = ~n26921 & n26924;
  assign n26926 = ~n26920 & n26925;
  assign n26927 = pi20  & n26926;
  assign n26928 = ~pi20  & ~n26926;
  assign n26929 = ~n26927 & ~n26928;
  assign n26930 = n26919 & ~n26929;
  assign n26931 = ~n26919 & n26929;
  assign n26932 = ~n26930 & ~n26931;
  assign n26933 = ~n26826 & n26932;
  assign n26934 = n26826 & ~n26932;
  assign n26935 = ~n26933 & ~n26934;
  assign n26936 = ~n26823 & ~n26935;
  assign n26937 = n26823 & n26935;
  assign n26938 = ~n26936 & ~n26937;
  assign n26939 = ~n26701 & ~n26705;
  assign n26940 = n26938 & n26939;
  assign n26941 = ~n26938 & ~n26939;
  assign n26942 = ~n26940 & ~n26941;
  assign n26943 = n6835 & n21183;
  assign n26944 = n7460 & n21180;
  assign n26945 = n6836 & n24030;
  assign n26946 = n7487 & n21076;
  assign n26947 = ~n26945 & ~n26946;
  assign n26948 = ~n26944 & n26947;
  assign n26949 = ~n26943 & n26948;
  assign n26950 = pi14  & n26949;
  assign n26951 = ~pi14  & ~n26949;
  assign n26952 = ~n26950 & ~n26951;
  assign n26953 = n26942 & ~n26952;
  assign n26954 = ~n26942 & n26952;
  assign n26955 = ~n26953 & ~n26954;
  assign n26956 = ~n26813 & n26955;
  assign n26957 = n26813 & ~n26955;
  assign n26958 = ~n26956 & ~n26957;
  assign n26959 = ~n26811 & ~n26958;
  assign n26960 = n26811 & n26958;
  assign n26961 = ~n26959 & ~n26960;
  assign n26962 = ~n26582 & n26722;
  assign n26963 = ~n26729 & ~n26962;
  assign n26964 = n26961 & n26963;
  assign n26965 = ~n26961 & ~n26963;
  assign n26966 = ~n26964 & ~n26965;
  assign n26967 = n8474 & n24676;
  assign n26968 = n9238 & n24748;
  assign n26969 = n8468 & ~n25529;
  assign n26970 = n9265 & n25521;
  assign n26971 = ~n26969 & ~n26970;
  assign n26972 = ~n26968 & n26971;
  assign n26973 = ~n26967 & n26972;
  assign n26974 = pi8  & n26973;
  assign n26975 = ~pi8  & ~n26973;
  assign n26976 = ~n26974 & ~n26975;
  assign n26977 = n26966 & ~n26976;
  assign n26978 = ~n26966 & n26976;
  assign n26979 = ~n26977 & ~n26978;
  assign n26980 = ~n26801 & n26979;
  assign n26981 = n26801 & ~n26979;
  assign n26982 = ~n26980 & ~n26981;
  assign n26983 = ~n26798 & ~n26982;
  assign n26984 = n26798 & n26982;
  assign n26985 = ~n26983 & ~n26984;
  assign n26986 = n26755 & ~n26765;
  assign n26987 = ~n26766 & ~n26986;
  assign n26988 = n11289 & n26987;
  assign n26989 = n11288 & n26532;
  assign n26990 = n19757 & n26764;
  assign n26991 = ~n26989 & ~n26990;
  assign n26992 = ~n26988 & n26991;
  assign n26993 = pi2  & n26992;
  assign n26994 = ~pi2  & ~n26992;
  assign n26995 = ~n26993 & ~n26994;
  assign n26996 = ~n26985 & ~n26995;
  assign n26997 = n26985 & n26995;
  assign n26998 = ~n26996 & ~n26997;
  assign n26999 = n26788 & ~n26998;
  assign n27000 = ~n26788 & n26998;
  assign n27001 = ~n26999 & ~n27000;
  assign n27002 = ~n26779 & ~n26782;
  assign n27003 = ~n27001 & n27002;
  assign n27004 = n27001 & ~n27002;
  assign n27005 = ~n27003 & ~n27004;
  assign n27006 = n26785 & n27005;
  assign n27007 = ~n26785 & ~n27005;
  assign po6  = ~n27006 & ~n27007;
  assign n27009 = ~n26798 & n26982;
  assign n27010 = ~n26996 & ~n27009;
  assign n27011 = ~n26977 & ~n26980;
  assign n27012 = ~n26811 & n26958;
  assign n27013 = ~n26965 & ~n27012;
  assign n27014 = ~n26953 & ~n26956;
  assign n27015 = ~n26823 & n26935;
  assign n27016 = ~n26941 & ~n27015;
  assign n27017 = ~n26930 & ~n26933;
  assign n27018 = ~n26836 & n26911;
  assign n27019 = ~n26918 & ~n27018;
  assign n27020 = ~n26906 & ~n26909;
  assign n27021 = ~n26890 & ~n26893;
  assign n27022 = ~n26876 & ~n26883;
  assign n27023 = ~n26887 & ~n27022;
  assign n27024 = n3117 & n12911;
  assign n27025 = n562 & n27024;
  assign n27026 = n3201 & n27025;
  assign n27027 = ~n252 & n27026;
  assign n27028 = n2653 & n12970;
  assign n27029 = n1011 & n27028;
  assign n27030 = ~n203 & n27029;
  assign n27031 = ~n325 & n27030;
  assign n27032 = n27027 & n27031;
  assign n27033 = n1169 & n7312;
  assign n27034 = n876 & n27033;
  assign n27035 = n306 & n27034;
  assign n27036 = ~n612 & n27035;
  assign n27037 = n138 & n2862;
  assign n27038 = ~n149 & n27037;
  assign n27039 = ~n414 & n27038;
  assign n27040 = n27036 & n27039;
  assign n27041 = n27032 & n27040;
  assign n27042 = pi2  & ~n26764;
  assign n27043 = n14362 & n26764;
  assign n27044 = ~n27042 & ~n27043;
  assign n27045 = ~n27041 & ~n27044;
  assign n27046 = n27041 & n27044;
  assign n27047 = ~n27045 & ~n27046;
  assign n27048 = n3641 & n21234;
  assign n27049 = n3740 & n21231;
  assign n27050 = n556 & n21494;
  assign n27051 = n3961 & n21228;
  assign n27052 = ~n27050 & ~n27051;
  assign n27053 = ~n27049 & n27052;
  assign n27054 = ~n27048 & n27053;
  assign n27055 = ~n27047 & n27054;
  assign n27056 = n27047 & ~n27054;
  assign n27057 = ~n27055 & ~n27056;
  assign n27058 = n27023 & ~n27057;
  assign n27059 = ~n27023 & n27057;
  assign n27060 = ~n27058 & ~n27059;
  assign n27061 = n4006 & n21225;
  assign n27062 = n4133 & n21222;
  assign n27063 = n4002 & n21973;
  assign n27064 = n4555 & n21219;
  assign n27065 = ~n27063 & ~n27064;
  assign n27066 = ~n27062 & n27065;
  assign n27067 = ~n27061 & n27066;
  assign n27068 = pi29  & n27067;
  assign n27069 = ~pi29  & ~n27067;
  assign n27070 = ~n27068 & ~n27069;
  assign n27071 = n27060 & ~n27070;
  assign n27072 = ~n27060 & n27070;
  assign n27073 = ~n27071 & ~n27072;
  assign n27074 = ~n27021 & n27073;
  assign n27075 = n27021 & ~n27073;
  assign n27076 = ~n27074 & ~n27075;
  assign n27077 = n4601 & n21216;
  assign n27078 = n4783 & n21213;
  assign n27079 = n4602 & n22376;
  assign n27080 = n4801 & n21210;
  assign n27081 = ~n27079 & ~n27080;
  assign n27082 = ~n27078 & n27081;
  assign n27083 = ~n27077 & n27082;
  assign n27084 = pi26  & n27083;
  assign n27085 = ~pi26  & ~n27083;
  assign n27086 = ~n27084 & ~n27085;
  assign n27087 = n27076 & ~n27086;
  assign n27088 = ~n27076 & n27086;
  assign n27089 = ~n27087 & ~n27088;
  assign n27090 = n27020 & ~n27089;
  assign n27091 = ~n27020 & n27089;
  assign n27092 = ~n27090 & ~n27091;
  assign n27093 = n5238 & n21207;
  assign n27094 = n71 & n21204;
  assign n27095 = n5239 & n22852;
  assign n27096 = n5326 & n21201;
  assign n27097 = ~n27095 & ~n27096;
  assign n27098 = ~n27094 & n27097;
  assign n27099 = ~n27093 & n27098;
  assign n27100 = pi23  & n27099;
  assign n27101 = ~pi23  & ~n27099;
  assign n27102 = ~n27100 & ~n27101;
  assign n27103 = n27092 & ~n27102;
  assign n27104 = ~n27092 & n27102;
  assign n27105 = ~n27103 & ~n27104;
  assign n27106 = n27019 & ~n27105;
  assign n27107 = ~n27019 & n27105;
  assign n27108 = ~n27106 & ~n27107;
  assign n27109 = n5435 & n21198;
  assign n27110 = n6055 & n21195;
  assign n27111 = n5429 & n23211;
  assign n27112 = n6071 & n21192;
  assign n27113 = ~n27111 & ~n27112;
  assign n27114 = ~n27110 & n27113;
  assign n27115 = ~n27109 & n27114;
  assign n27116 = pi20  & n27115;
  assign n27117 = ~pi20  & ~n27115;
  assign n27118 = ~n27116 & ~n27117;
  assign n27119 = n27108 & ~n27118;
  assign n27120 = ~n27108 & n27118;
  assign n27121 = ~n27119 & ~n27120;
  assign n27122 = n27017 & ~n27121;
  assign n27123 = ~n27017 & n27121;
  assign n27124 = ~n27122 & ~n27123;
  assign n27125 = n6184 & n21189;
  assign n27126 = n6527 & n21186;
  assign n27127 = n6185 & n23369;
  assign n27128 = n6543 & n21183;
  assign n27129 = ~n27127 & ~n27128;
  assign n27130 = ~n27126 & n27129;
  assign n27131 = ~n27125 & n27130;
  assign n27132 = pi17  & n27131;
  assign n27133 = ~pi17  & ~n27131;
  assign n27134 = ~n27132 & ~n27133;
  assign n27135 = n27124 & ~n27134;
  assign n27136 = ~n27124 & n27134;
  assign n27137 = ~n27135 & ~n27136;
  assign n27138 = n27016 & ~n27137;
  assign n27139 = ~n27016 & n27137;
  assign n27140 = ~n27138 & ~n27139;
  assign n27141 = n6835 & n21180;
  assign n27142 = n7460 & n21076;
  assign n27143 = n6836 & n24012;
  assign n27144 = n7487 & n21176;
  assign n27145 = ~n27143 & ~n27144;
  assign n27146 = ~n27142 & n27145;
  assign n27147 = ~n27141 & n27146;
  assign n27148 = pi14  & n27147;
  assign n27149 = ~pi14  & ~n27147;
  assign n27150 = ~n27148 & ~n27149;
  assign n27151 = n27140 & ~n27150;
  assign n27152 = ~n27140 & n27150;
  assign n27153 = ~n27151 & ~n27152;
  assign n27154 = n27014 & ~n27153;
  assign n27155 = ~n27014 & n27153;
  assign n27156 = ~n27154 & ~n27155;
  assign n27157 = n7654 & n21464;
  assign n27158 = n8091 & n24607;
  assign n27159 = n7648 & n24770;
  assign n27160 = n8120 & n24676;
  assign n27161 = ~n27159 & ~n27160;
  assign n27162 = ~n27158 & n27161;
  assign n27163 = ~n27157 & n27162;
  assign n27164 = pi11  & n27163;
  assign n27165 = ~pi11  & ~n27163;
  assign n27166 = ~n27164 & ~n27165;
  assign n27167 = n27156 & ~n27166;
  assign n27168 = ~n27156 & n27166;
  assign n27169 = ~n27167 & ~n27168;
  assign n27170 = n27013 & ~n27169;
  assign n27171 = ~n27013 & n27169;
  assign n27172 = ~n27170 & ~n27171;
  assign n27173 = n8474 & n24748;
  assign n27174 = n9238 & n25521;
  assign n27175 = n8468 & n25793;
  assign n27176 = n9265 & n25785;
  assign n27177 = ~n27175 & ~n27176;
  assign n27178 = ~n27174 & n27177;
  assign n27179 = ~n27173 & n27178;
  assign n27180 = pi8  & n27179;
  assign n27181 = ~pi8  & ~n27179;
  assign n27182 = ~n27180 & ~n27181;
  assign n27183 = n27172 & ~n27182;
  assign n27184 = ~n27172 & n27182;
  assign n27185 = ~n27183 & ~n27184;
  assign n27186 = n27011 & ~n27185;
  assign n27187 = ~n27011 & n27185;
  assign n27188 = ~n27186 & ~n27187;
  assign n27189 = n9725 & n26043;
  assign n27190 = n10702 & n26284;
  assign n27191 = n9719 & n26540;
  assign n27192 = n11267 & n26532;
  assign n27193 = ~n27191 & ~n27192;
  assign n27194 = ~n27190 & n27193;
  assign n27195 = ~n27189 & n27194;
  assign n27196 = pi5  & n27195;
  assign n27197 = ~pi5  & ~n27195;
  assign n27198 = ~n27196 & ~n27197;
  assign n27199 = n27188 & ~n27198;
  assign n27200 = ~n27188 & n27198;
  assign n27201 = ~n27199 & ~n27200;
  assign n27202 = n27010 & ~n27201;
  assign n27203 = ~n27010 & n27201;
  assign n27204 = ~n27202 & ~n27203;
  assign n27205 = ~n27000 & ~n27004;
  assign n27206 = ~n27204 & n27205;
  assign n27207 = n27204 & ~n27205;
  assign n27208 = ~n27206 & ~n27207;
  assign n27209 = n27006 & n27208;
  assign n27210 = ~n27006 & ~n27208;
  assign po7  = ~n27209 & ~n27210;
  assign n27212 = ~n27046 & ~n27054;
  assign n27213 = ~n27045 & ~n27212;
  assign n27214 = n364 & n22726;
  assign n27215 = n2192 & n27214;
  assign n27216 = n1435 & n27215;
  assign n27217 = n148 & n27216;
  assign n27218 = ~n324 & n27217;
  assign n27219 = n2143 & n3122;
  assign n27220 = n2566 & n27219;
  assign n27221 = n4260 & n27220;
  assign n27222 = ~n374 & n27221;
  assign n27223 = n27218 & n27222;
  assign n27224 = ~n308 & n476;
  assign n27225 = ~n632 & n15340;
  assign n27226 = ~n473 & n27225;
  assign n27227 = n27224 & n27226;
  assign n27228 = n2833 & n27227;
  assign n27229 = ~n466 & n27228;
  assign n27230 = n1775 & n15298;
  assign n27231 = n684 & n27230;
  assign n27232 = n1395 & n27231;
  assign n27233 = ~n219 & n27232;
  assign n27234 = n27229 & n27233;
  assign n27235 = n27223 & n27234;
  assign n27236 = ~n27044 & ~n27235;
  assign n27237 = n27044 & n27235;
  assign n27238 = ~n27236 & ~n27237;
  assign n27239 = n27213 & ~n27238;
  assign n27240 = ~n27213 & n27238;
  assign n27241 = ~n27239 & ~n27240;
  assign n27242 = n3641 & n21231;
  assign n27243 = n3740 & n21228;
  assign n27244 = n556 & n22001;
  assign n27245 = n3961 & n21225;
  assign n27246 = ~n27244 & ~n27245;
  assign n27247 = ~n27243 & n27246;
  assign n27248 = ~n27242 & n27247;
  assign n27249 = n27241 & n27248;
  assign n27250 = ~n27241 & ~n27248;
  assign n27251 = ~n27249 & ~n27250;
  assign n27252 = ~n27059 & ~n27071;
  assign n27253 = n27251 & n27252;
  assign n27254 = ~n27251 & ~n27252;
  assign n27255 = ~n27253 & ~n27254;
  assign n27256 = n4006 & n21222;
  assign n27257 = n4133 & n21219;
  assign n27258 = n4002 & n22225;
  assign n27259 = n4555 & n21216;
  assign n27260 = ~n27258 & ~n27259;
  assign n27261 = ~n27257 & n27260;
  assign n27262 = ~n27256 & n27261;
  assign n27263 = pi29  & n27262;
  assign n27264 = ~pi29  & ~n27262;
  assign n27265 = ~n27263 & ~n27264;
  assign n27266 = n27255 & n27265;
  assign n27267 = ~n27255 & ~n27265;
  assign n27268 = ~n27266 & ~n27267;
  assign n27269 = n4601 & n21213;
  assign n27270 = n4783 & n21210;
  assign n27271 = n4602 & n22363;
  assign n27272 = n4801 & n21207;
  assign n27273 = ~n27271 & ~n27272;
  assign n27274 = ~n27270 & n27273;
  assign n27275 = ~n27269 & n27274;
  assign n27276 = pi26  & n27275;
  assign n27277 = ~pi26  & ~n27275;
  assign n27278 = ~n27276 & ~n27277;
  assign n27279 = ~n27268 & n27278;
  assign n27280 = n27268 & ~n27278;
  assign n27281 = ~n27279 & ~n27280;
  assign n27282 = ~n27074 & n27086;
  assign n27283 = ~n27075 & ~n27282;
  assign n27284 = n27281 & ~n27283;
  assign n27285 = ~n27281 & n27283;
  assign n27286 = ~n27284 & ~n27285;
  assign n27287 = n5238 & n21204;
  assign n27288 = n71 & n21201;
  assign n27289 = n5239 & n22832;
  assign n27290 = n5326 & n21198;
  assign n27291 = ~n27289 & ~n27290;
  assign n27292 = ~n27288 & n27291;
  assign n27293 = ~n27287 & n27292;
  assign n27294 = pi23  & n27293;
  assign n27295 = ~pi23  & ~n27293;
  assign n27296 = ~n27294 & ~n27295;
  assign n27297 = n27286 & ~n27296;
  assign n27298 = ~n27286 & n27296;
  assign n27299 = ~n27297 & ~n27298;
  assign n27300 = ~n27091 & n27102;
  assign n27301 = ~n27090 & ~n27300;
  assign n27302 = ~n27299 & ~n27301;
  assign n27303 = n27299 & n27301;
  assign n27304 = ~n27302 & ~n27303;
  assign n27305 = n5435 & n21195;
  assign n27306 = n6055 & n21192;
  assign n27307 = n5429 & n23399;
  assign n27308 = n6071 & n21189;
  assign n27309 = ~n27307 & ~n27308;
  assign n27310 = ~n27306 & n27309;
  assign n27311 = ~n27305 & n27310;
  assign n27312 = pi20  & n27311;
  assign n27313 = ~pi20  & ~n27311;
  assign n27314 = ~n27312 & ~n27313;
  assign n27315 = n27304 & ~n27314;
  assign n27316 = ~n27304 & n27314;
  assign n27317 = ~n27315 & ~n27316;
  assign n27318 = ~n27107 & n27118;
  assign n27319 = ~n27106 & ~n27318;
  assign n27320 = ~n27317 & ~n27319;
  assign n27321 = n27317 & n27319;
  assign n27322 = ~n27320 & ~n27321;
  assign n27323 = n6184 & n21186;
  assign n27324 = n6527 & n21183;
  assign n27325 = n6185 & n23991;
  assign n27326 = n6543 & n21180;
  assign n27327 = ~n27325 & ~n27326;
  assign n27328 = ~n27324 & n27327;
  assign n27329 = ~n27323 & n27328;
  assign n27330 = pi17  & n27329;
  assign n27331 = ~pi17  & ~n27329;
  assign n27332 = ~n27330 & ~n27331;
  assign n27333 = n27322 & ~n27332;
  assign n27334 = ~n27322 & n27332;
  assign n27335 = ~n27333 & ~n27334;
  assign n27336 = ~n27123 & n27134;
  assign n27337 = ~n27122 & ~n27336;
  assign n27338 = ~n27335 & ~n27337;
  assign n27339 = n27335 & n27337;
  assign n27340 = ~n27338 & ~n27339;
  assign n27341 = n6835 & n21076;
  assign n27342 = n7460 & n21176;
  assign n27343 = n6836 & ~n21470;
  assign n27344 = n7487 & n21464;
  assign n27345 = ~n27343 & ~n27344;
  assign n27346 = ~n27342 & n27345;
  assign n27347 = ~n27341 & n27346;
  assign n27348 = pi14  & n27347;
  assign n27349 = ~pi14  & ~n27347;
  assign n27350 = ~n27348 & ~n27349;
  assign n27351 = n27340 & ~n27350;
  assign n27352 = ~n27340 & n27350;
  assign n27353 = ~n27351 & ~n27352;
  assign n27354 = ~n27139 & n27150;
  assign n27355 = ~n27138 & ~n27354;
  assign n27356 = ~n27353 & ~n27355;
  assign n27357 = n27353 & n27355;
  assign n27358 = ~n27356 & ~n27357;
  assign n27359 = n7654 & n24607;
  assign n27360 = n8091 & n24676;
  assign n27361 = n7648 & ~n24754;
  assign n27362 = n8120 & n24748;
  assign n27363 = ~n27361 & ~n27362;
  assign n27364 = ~n27360 & n27363;
  assign n27365 = ~n27359 & n27364;
  assign n27366 = pi11  & n27365;
  assign n27367 = ~pi11  & ~n27365;
  assign n27368 = ~n27366 & ~n27367;
  assign n27369 = n27358 & ~n27368;
  assign n27370 = ~n27358 & n27368;
  assign n27371 = ~n27369 & ~n27370;
  assign n27372 = ~n27155 & n27166;
  assign n27373 = ~n27154 & ~n27372;
  assign n27374 = ~n27371 & ~n27373;
  assign n27375 = n27371 & n27373;
  assign n27376 = ~n27374 & ~n27375;
  assign n27377 = n8474 & n25521;
  assign n27378 = n9238 & n25785;
  assign n27379 = n8468 & n26049;
  assign n27380 = n9265 & n26043;
  assign n27381 = ~n27379 & ~n27380;
  assign n27382 = ~n27378 & n27381;
  assign n27383 = ~n27377 & n27382;
  assign n27384 = pi8  & n27383;
  assign n27385 = ~pi8  & ~n27383;
  assign n27386 = ~n27384 & ~n27385;
  assign n27387 = n27376 & ~n27386;
  assign n27388 = ~n27376 & n27386;
  assign n27389 = ~n27387 & ~n27388;
  assign n27390 = ~n27171 & n27182;
  assign n27391 = ~n27170 & ~n27390;
  assign n27392 = ~n27389 & ~n27391;
  assign n27393 = n27389 & n27391;
  assign n27394 = ~n27392 & ~n27393;
  assign n27395 = n9725 & n26284;
  assign n27396 = n10702 & n26532;
  assign n27397 = n9719 & ~n26770;
  assign n27398 = n11267 & n26764;
  assign n27399 = ~n27397 & ~n27398;
  assign n27400 = ~n27396 & n27399;
  assign n27401 = ~n27395 & n27400;
  assign n27402 = pi5  & n27401;
  assign n27403 = ~pi5  & ~n27401;
  assign n27404 = ~n27402 & ~n27403;
  assign n27405 = n27394 & ~n27404;
  assign n27406 = ~n27394 & n27404;
  assign n27407 = ~n27405 & ~n27406;
  assign n27408 = ~n27187 & n27198;
  assign n27409 = ~n27186 & ~n27408;
  assign n27410 = ~n27407 & ~n27409;
  assign n27411 = n27407 & n27409;
  assign n27412 = ~n27410 & ~n27411;
  assign n27413 = ~n27203 & ~n27207;
  assign n27414 = ~n27412 & n27413;
  assign n27415 = n27412 & ~n27413;
  assign n27416 = ~n27414 & ~n27415;
  assign n27417 = n27209 & n27416;
  assign n27418 = ~n27209 & ~n27416;
  assign po8  = ~n27417 & ~n27418;
  assign n27420 = n9719 & n26987;
  assign n27421 = n9725 & n26532;
  assign n27422 = n18016 & n26764;
  assign n27423 = ~n27421 & ~n27422;
  assign n27424 = ~n27420 & n27423;
  assign n27425 = pi5  & n27424;
  assign n27426 = ~pi5  & ~n27424;
  assign n27427 = ~n27425 & ~n27426;
  assign n27428 = ~n27375 & n27386;
  assign n27429 = ~n27374 & ~n27428;
  assign n27430 = ~n27427 & n27429;
  assign n27431 = n27427 & ~n27429;
  assign n27432 = ~n27430 & ~n27431;
  assign n27433 = ~n27213 & ~n27237;
  assign n27434 = ~n27236 & ~n27433;
  assign n27435 = n1440 & n4155;
  assign n27436 = ~n391 & n27435;
  assign n27437 = n5837 & n14585;
  assign n27438 = n2915 & n27437;
  assign n27439 = ~n692 & n27438;
  assign n27440 = n27436 & n27439;
  assign n27441 = n1716 & n3460;
  assign n27442 = n797 & n27441;
  assign n27443 = ~n579 & n27442;
  assign n27444 = n1908 & n3113;
  assign n27445 = n896 & n27444;
  assign n27446 = n3159 & n27445;
  assign n27447 = ~n588 & n27446;
  assign n27448 = ~n197 & n27447;
  assign n27449 = n27443 & n27448;
  assign n27450 = n27440 & n27449;
  assign n27451 = ~n27044 & ~n27450;
  assign n27452 = n27044 & n27450;
  assign n27453 = ~n27451 & ~n27452;
  assign n27454 = n27434 & ~n27453;
  assign n27455 = ~n27434 & n27453;
  assign n27456 = ~n27454 & ~n27455;
  assign n27457 = n3641 & n21228;
  assign n27458 = n3740 & n21225;
  assign n27459 = n556 & n21988;
  assign n27460 = n3961 & n21222;
  assign n27461 = ~n27459 & ~n27460;
  assign n27462 = ~n27458 & n27461;
  assign n27463 = ~n27457 & n27462;
  assign n27464 = n27456 & n27463;
  assign n27465 = ~n27456 & ~n27463;
  assign n27466 = ~n27464 & ~n27465;
  assign n27467 = n27241 & ~n27248;
  assign n27468 = ~n27254 & ~n27467;
  assign n27469 = n27466 & n27468;
  assign n27470 = ~n27466 & ~n27468;
  assign n27471 = ~n27469 & ~n27470;
  assign n27472 = n4006 & n21219;
  assign n27473 = n4133 & n21216;
  assign n27474 = n4002 & n22394;
  assign n27475 = n4555 & n21213;
  assign n27476 = ~n27474 & ~n27475;
  assign n27477 = ~n27473 & n27476;
  assign n27478 = ~n27472 & n27477;
  assign n27479 = pi29  & n27478;
  assign n27480 = ~pi29  & ~n27478;
  assign n27481 = ~n27479 & ~n27480;
  assign n27482 = n27471 & n27481;
  assign n27483 = ~n27471 & ~n27481;
  assign n27484 = ~n27482 & ~n27483;
  assign n27485 = n4601 & n21210;
  assign n27486 = n4783 & n21207;
  assign n27487 = n4602 & n22810;
  assign n27488 = n4801 & n21204;
  assign n27489 = ~n27487 & ~n27488;
  assign n27490 = ~n27486 & n27489;
  assign n27491 = ~n27485 & n27490;
  assign n27492 = pi26  & n27491;
  assign n27493 = ~pi26  & ~n27491;
  assign n27494 = ~n27492 & ~n27493;
  assign n27495 = ~n27484 & n27494;
  assign n27496 = n27484 & ~n27494;
  assign n27497 = ~n27495 & ~n27496;
  assign n27498 = n27255 & ~n27265;
  assign n27499 = ~n27268 & ~n27278;
  assign n27500 = ~n27498 & ~n27499;
  assign n27501 = n27497 & n27500;
  assign n27502 = ~n27497 & ~n27500;
  assign n27503 = ~n27501 & ~n27502;
  assign n27504 = n5238 & n21201;
  assign n27505 = n71 & n21198;
  assign n27506 = n5239 & n21482;
  assign n27507 = n5326 & n21195;
  assign n27508 = ~n27506 & ~n27507;
  assign n27509 = ~n27505 & n27508;
  assign n27510 = ~n27504 & n27509;
  assign n27511 = pi23  & n27510;
  assign n27512 = ~pi23  & ~n27510;
  assign n27513 = ~n27511 & ~n27512;
  assign n27514 = n27503 & ~n27513;
  assign n27515 = ~n27503 & n27513;
  assign n27516 = ~n27514 & ~n27515;
  assign n27517 = ~n27285 & n27296;
  assign n27518 = ~n27284 & ~n27517;
  assign n27519 = ~n27516 & ~n27518;
  assign n27520 = n27516 & n27518;
  assign n27521 = ~n27519 & ~n27520;
  assign n27522 = n5435 & n21192;
  assign n27523 = n6055 & n21189;
  assign n27524 = n5429 & n23384;
  assign n27525 = n6071 & n21186;
  assign n27526 = ~n27524 & ~n27525;
  assign n27527 = ~n27523 & n27526;
  assign n27528 = ~n27522 & n27527;
  assign n27529 = pi20  & n27528;
  assign n27530 = ~pi20  & ~n27528;
  assign n27531 = ~n27529 & ~n27530;
  assign n27532 = n27521 & ~n27531;
  assign n27533 = ~n27521 & n27531;
  assign n27534 = ~n27532 & ~n27533;
  assign n27535 = ~n27303 & n27314;
  assign n27536 = ~n27302 & ~n27535;
  assign n27537 = ~n27534 & ~n27536;
  assign n27538 = n27534 & n27536;
  assign n27539 = ~n27537 & ~n27538;
  assign n27540 = n6184 & n21183;
  assign n27541 = n6527 & n21180;
  assign n27542 = n6185 & n24030;
  assign n27543 = n6543 & n21076;
  assign n27544 = ~n27542 & ~n27543;
  assign n27545 = ~n27541 & n27544;
  assign n27546 = ~n27540 & n27545;
  assign n27547 = pi17  & n27546;
  assign n27548 = ~pi17  & ~n27546;
  assign n27549 = ~n27547 & ~n27548;
  assign n27550 = n27539 & ~n27549;
  assign n27551 = ~n27539 & n27549;
  assign n27552 = ~n27550 & ~n27551;
  assign n27553 = ~n27321 & n27332;
  assign n27554 = ~n27320 & ~n27553;
  assign n27555 = ~n27552 & ~n27554;
  assign n27556 = n27552 & n27554;
  assign n27557 = ~n27555 & ~n27556;
  assign n27558 = n6835 & n21176;
  assign n27559 = n7460 & n21464;
  assign n27560 = n6836 & n24782;
  assign n27561 = n7487 & n24607;
  assign n27562 = ~n27560 & ~n27561;
  assign n27563 = ~n27559 & n27562;
  assign n27564 = ~n27558 & n27563;
  assign n27565 = pi14  & n27564;
  assign n27566 = ~pi14  & ~n27564;
  assign n27567 = ~n27565 & ~n27566;
  assign n27568 = n27557 & ~n27567;
  assign n27569 = ~n27557 & n27567;
  assign n27570 = ~n27568 & ~n27569;
  assign n27571 = ~n27339 & n27350;
  assign n27572 = ~n27338 & ~n27571;
  assign n27573 = ~n27570 & ~n27572;
  assign n27574 = n27570 & n27572;
  assign n27575 = ~n27573 & ~n27574;
  assign n27576 = n7654 & n24676;
  assign n27577 = n8091 & n24748;
  assign n27578 = n7648 & ~n25529;
  assign n27579 = n8120 & n25521;
  assign n27580 = ~n27578 & ~n27579;
  assign n27581 = ~n27577 & n27580;
  assign n27582 = ~n27576 & n27581;
  assign n27583 = pi11  & n27582;
  assign n27584 = ~pi11  & ~n27582;
  assign n27585 = ~n27583 & ~n27584;
  assign n27586 = n27575 & ~n27585;
  assign n27587 = ~n27575 & n27585;
  assign n27588 = ~n27586 & ~n27587;
  assign n27589 = ~n27357 & n27368;
  assign n27590 = ~n27356 & ~n27589;
  assign n27591 = ~n27588 & ~n27590;
  assign n27592 = n27588 & n27590;
  assign n27593 = ~n27591 & ~n27592;
  assign n27594 = n8474 & n25785;
  assign n27595 = n9238 & n26043;
  assign n27596 = n8468 & ~n26290;
  assign n27597 = n9265 & n26284;
  assign n27598 = ~n27596 & ~n27597;
  assign n27599 = ~n27595 & n27598;
  assign n27600 = ~n27594 & n27599;
  assign n27601 = pi8  & n27600;
  assign n27602 = ~pi8  & ~n27600;
  assign n27603 = ~n27601 & ~n27602;
  assign n27604 = n27593 & ~n27603;
  assign n27605 = ~n27593 & n27603;
  assign n27606 = ~n27604 & ~n27605;
  assign n27607 = n27432 & n27606;
  assign n27608 = ~n27432 & ~n27606;
  assign n27609 = ~n27607 & ~n27608;
  assign n27610 = ~n27393 & n27404;
  assign n27611 = ~n27392 & ~n27610;
  assign n27612 = ~n27609 & ~n27611;
  assign n27613 = n27609 & n27611;
  assign n27614 = ~n27612 & ~n27613;
  assign n27615 = ~n27411 & ~n27415;
  assign n27616 = ~n27614 & n27615;
  assign n27617 = n27614 & ~n27615;
  assign n27618 = ~n27616 & ~n27617;
  assign n27619 = n27417 & n27618;
  assign n27620 = ~n27417 & ~n27618;
  assign po9  = ~n27619 & ~n27620;
  assign n27622 = ~n27613 & ~n27617;
  assign n27623 = n27471 & ~n27481;
  assign n27624 = ~n27484 & ~n27494;
  assign n27625 = ~n27623 & ~n27624;
  assign n27626 = n4601 & n21207;
  assign n27627 = n4783 & n21204;
  assign n27628 = n4602 & n22852;
  assign n27629 = n4801 & n21201;
  assign n27630 = ~n27628 & ~n27629;
  assign n27631 = ~n27627 & n27630;
  assign n27632 = ~n27626 & n27631;
  assign n27633 = pi26  & n27632;
  assign n27634 = ~pi26  & ~n27632;
  assign n27635 = ~n27633 & ~n27634;
  assign n27636 = n27456 & ~n27463;
  assign n27637 = ~n27470 & ~n27636;
  assign n27638 = ~n27434 & ~n27452;
  assign n27639 = ~n27451 & ~n27638;
  assign n27640 = n5056 & n5087;
  assign n27641 = ~n601 & n27640;
  assign n27642 = n765 & n13119;
  assign n27643 = n437 & n27642;
  assign n27644 = ~n463 & n27643;
  assign n27645 = n27641 & n27644;
  assign n27646 = n2613 & n4368;
  assign n27647 = n3187 & n27646;
  assign n27648 = ~n578 & n27647;
  assign n27649 = n1872 & n1982;
  assign n27650 = n184 & n27649;
  assign n27651 = n22298 & n27650;
  assign n27652 = ~n468 & n27651;
  assign n27653 = n27648 & n27652;
  assign n27654 = n27645 & n27653;
  assign n27655 = n27044 & n27654;
  assign n27656 = ~n27044 & ~n27654;
  assign n27657 = ~n27655 & ~n27656;
  assign n27658 = ~n14370 & n26764;
  assign n27659 = ~pi5  & n27658;
  assign n27660 = pi5  & ~n27658;
  assign n27661 = ~n27659 & ~n27660;
  assign n27662 = ~n27657 & n27661;
  assign n27663 = n27657 & ~n27661;
  assign n27664 = ~n27662 & ~n27663;
  assign n27665 = ~n27639 & n27664;
  assign n27666 = n27639 & ~n27664;
  assign n27667 = ~n27665 & ~n27666;
  assign n27668 = n3641 & n21225;
  assign n27669 = n3740 & n21222;
  assign n27670 = n556 & n21973;
  assign n27671 = n3961 & n21219;
  assign n27672 = ~n27670 & ~n27671;
  assign n27673 = ~n27669 & n27672;
  assign n27674 = ~n27668 & n27673;
  assign n27675 = n27667 & ~n27674;
  assign n27676 = ~n27667 & n27674;
  assign n27677 = ~n27675 & ~n27676;
  assign n27678 = n27637 & ~n27677;
  assign n27679 = ~n27637 & n27677;
  assign n27680 = ~n27678 & ~n27679;
  assign n27681 = n4006 & n21216;
  assign n27682 = n4133 & n21213;
  assign n27683 = n4002 & n22376;
  assign n27684 = n4555 & n21210;
  assign n27685 = ~n27683 & ~n27684;
  assign n27686 = ~n27682 & n27685;
  assign n27687 = ~n27681 & n27686;
  assign n27688 = pi29  & n27687;
  assign n27689 = ~pi29  & ~n27687;
  assign n27690 = ~n27688 & ~n27689;
  assign n27691 = n27680 & ~n27690;
  assign n27692 = ~n27680 & n27690;
  assign n27693 = ~n27691 & ~n27692;
  assign n27694 = ~n27635 & n27693;
  assign n27695 = n27635 & ~n27693;
  assign n27696 = ~n27694 & ~n27695;
  assign n27697 = n27625 & ~n27696;
  assign n27698 = ~n27625 & n27696;
  assign n27699 = ~n27697 & ~n27698;
  assign n27700 = n5238 & n21198;
  assign n27701 = n71 & n21195;
  assign n27702 = n5239 & n23211;
  assign n27703 = n5326 & n21192;
  assign n27704 = ~n27702 & ~n27703;
  assign n27705 = ~n27701 & n27704;
  assign n27706 = ~n27700 & n27705;
  assign n27707 = pi23  & n27706;
  assign n27708 = ~pi23  & ~n27706;
  assign n27709 = ~n27707 & ~n27708;
  assign n27710 = n27699 & n27709;
  assign n27711 = ~n27699 & ~n27709;
  assign n27712 = ~n27710 & ~n27711;
  assign n27713 = ~n27502 & n27513;
  assign n27714 = ~n27501 & ~n27713;
  assign n27715 = n27712 & ~n27714;
  assign n27716 = ~n27712 & n27714;
  assign n27717 = ~n27715 & ~n27716;
  assign n27718 = n5435 & n21189;
  assign n27719 = n6055 & n21186;
  assign n27720 = n5429 & n23369;
  assign n27721 = n6071 & n21183;
  assign n27722 = ~n27720 & ~n27721;
  assign n27723 = ~n27719 & n27722;
  assign n27724 = ~n27718 & n27723;
  assign n27725 = pi20  & n27724;
  assign n27726 = ~pi20  & ~n27724;
  assign n27727 = ~n27725 & ~n27726;
  assign n27728 = n27717 & n27727;
  assign n27729 = ~n27717 & ~n27727;
  assign n27730 = ~n27728 & ~n27729;
  assign n27731 = ~n27520 & n27531;
  assign n27732 = ~n27519 & ~n27731;
  assign n27733 = n27730 & ~n27732;
  assign n27734 = ~n27730 & n27732;
  assign n27735 = ~n27733 & ~n27734;
  assign n27736 = n6184 & n21180;
  assign n27737 = n6527 & n21076;
  assign n27738 = n6185 & n24012;
  assign n27739 = n6543 & n21176;
  assign n27740 = ~n27738 & ~n27739;
  assign n27741 = ~n27737 & n27740;
  assign n27742 = ~n27736 & n27741;
  assign n27743 = pi17  & n27742;
  assign n27744 = ~pi17  & ~n27742;
  assign n27745 = ~n27743 & ~n27744;
  assign n27746 = n27735 & n27745;
  assign n27747 = ~n27735 & ~n27745;
  assign n27748 = ~n27746 & ~n27747;
  assign n27749 = ~n27538 & n27549;
  assign n27750 = ~n27537 & ~n27749;
  assign n27751 = n27748 & ~n27750;
  assign n27752 = ~n27748 & n27750;
  assign n27753 = ~n27751 & ~n27752;
  assign n27754 = n6835 & n21464;
  assign n27755 = n7460 & n24607;
  assign n27756 = n6836 & n24770;
  assign n27757 = n7487 & n24676;
  assign n27758 = ~n27756 & ~n27757;
  assign n27759 = ~n27755 & n27758;
  assign n27760 = ~n27754 & n27759;
  assign n27761 = pi14  & n27760;
  assign n27762 = ~pi14  & ~n27760;
  assign n27763 = ~n27761 & ~n27762;
  assign n27764 = ~n27556 & n27567;
  assign n27765 = ~n27555 & ~n27764;
  assign n27766 = n27763 & n27765;
  assign n27767 = ~n27763 & ~n27765;
  assign n27768 = ~n27766 & ~n27767;
  assign n27769 = ~n27753 & n27768;
  assign n27770 = n27753 & ~n27768;
  assign n27771 = ~n27769 & ~n27770;
  assign n27772 = n7654 & n24748;
  assign n27773 = n8091 & n25521;
  assign n27774 = n7648 & n25793;
  assign n27775 = n8120 & n25785;
  assign n27776 = ~n27774 & ~n27775;
  assign n27777 = ~n27773 & n27776;
  assign n27778 = ~n27772 & n27777;
  assign n27779 = pi11  & n27778;
  assign n27780 = ~pi11  & ~n27778;
  assign n27781 = ~n27779 & ~n27780;
  assign n27782 = n27771 & n27781;
  assign n27783 = ~n27771 & ~n27781;
  assign n27784 = ~n27782 & ~n27783;
  assign n27785 = ~n27574 & n27585;
  assign n27786 = ~n27573 & ~n27785;
  assign n27787 = n27784 & ~n27786;
  assign n27788 = ~n27784 & n27786;
  assign n27789 = ~n27787 & ~n27788;
  assign n27790 = n8474 & n26043;
  assign n27791 = n9238 & n26284;
  assign n27792 = n8468 & n26540;
  assign n27793 = n9265 & n26532;
  assign n27794 = ~n27792 & ~n27793;
  assign n27795 = ~n27791 & n27794;
  assign n27796 = ~n27790 & n27795;
  assign n27797 = pi8  & n27796;
  assign n27798 = ~pi8  & ~n27796;
  assign n27799 = ~n27797 & ~n27798;
  assign n27800 = ~n27592 & n27603;
  assign n27801 = ~n27591 & ~n27800;
  assign n27802 = n27799 & n27801;
  assign n27803 = ~n27799 & ~n27801;
  assign n27804 = ~n27802 & ~n27803;
  assign n27805 = ~n27789 & n27804;
  assign n27806 = n27789 & ~n27804;
  assign n27807 = ~n27805 & ~n27806;
  assign n27808 = ~n27430 & ~n27606;
  assign n27809 = ~n27431 & ~n27808;
  assign n27810 = n27807 & n27809;
  assign n27811 = ~n27807 & ~n27809;
  assign n27812 = ~n27810 & ~n27811;
  assign n27813 = ~n27622 & n27812;
  assign n27814 = n27622 & ~n27812;
  assign n27815 = ~n27813 & ~n27814;
  assign n27816 = ~n27619 & ~n27815;
  assign n27817 = n27619 & n27815;
  assign po10  = ~n27816 & ~n27817;
  assign n27819 = ~n27810 & ~n27813;
  assign n27820 = ~n27799 & n27801;
  assign n27821 = ~n27806 & ~n27820;
  assign n27822 = n27771 & ~n27781;
  assign n27823 = ~n27788 & ~n27822;
  assign n27824 = ~n27763 & n27765;
  assign n27825 = ~n27770 & ~n27824;
  assign n27826 = n27735 & ~n27745;
  assign n27827 = ~n27752 & ~n27826;
  assign n27828 = n27717 & ~n27727;
  assign n27829 = ~n27734 & ~n27828;
  assign n27830 = n27699 & ~n27709;
  assign n27831 = ~n27716 & ~n27830;
  assign n27832 = ~n27694 & ~n27698;
  assign n27833 = ~n27665 & ~n27675;
  assign n27834 = n27044 & ~n27654;
  assign n27835 = ~n27662 & ~n27834;
  assign n27836 = n2340 & n3470;
  assign n27837 = ~n372 & n27836;
  assign n27838 = n2123 & n6639;
  assign n27839 = ~n232 & n27838;
  assign n27840 = n1123 & n2105;
  assign n27841 = n1775 & n27840;
  assign n27842 = ~n374 & n27841;
  assign n27843 = n27839 & n27842;
  assign n27844 = n1565 & n2037;
  assign n27845 = ~n307 & n27844;
  assign n27846 = n857 & n7284;
  assign n27847 = ~n85 & n27846;
  assign n27848 = n27845 & n27847;
  assign n27849 = n27843 & n27848;
  assign n27850 = n1526 & n27849;
  assign n27851 = ~n430 & n27850;
  assign n27852 = ~n106 & n27851;
  assign n27853 = n27837 & n27852;
  assign n27854 = n1238 & n7251;
  assign n27855 = n2481 & n27854;
  assign n27856 = n4444 & n27855;
  assign n27857 = n1271 & n27856;
  assign n27858 = ~n206 & n27857;
  assign n27859 = ~n88 & n27858;
  assign n27860 = n1543 & n2262;
  assign n27861 = n1232 & n27860;
  assign n27862 = ~n173 & n27861;
  assign n27863 = ~n197 & n27862;
  assign n27864 = n27859 & n27863;
  assign n27865 = n27853 & n27864;
  assign n27866 = ~n27835 & n27865;
  assign n27867 = n27835 & ~n27865;
  assign n27868 = ~n27866 & ~n27867;
  assign n27869 = n3641 & n21222;
  assign n27870 = n3740 & n21219;
  assign n27871 = n556 & n22225;
  assign n27872 = n3961 & n21216;
  assign n27873 = ~n27871 & ~n27872;
  assign n27874 = ~n27870 & n27873;
  assign n27875 = ~n27869 & n27874;
  assign n27876 = n27868 & ~n27875;
  assign n27877 = ~n27868 & n27875;
  assign n27878 = ~n27876 & ~n27877;
  assign n27879 = n27833 & ~n27878;
  assign n27880 = ~n27833 & n27878;
  assign n27881 = ~n27879 & ~n27880;
  assign n27882 = n4006 & n21213;
  assign n27883 = n4133 & n21210;
  assign n27884 = n4002 & n22363;
  assign n27885 = n4555 & n21207;
  assign n27886 = ~n27884 & ~n27885;
  assign n27887 = ~n27883 & n27886;
  assign n27888 = ~n27882 & n27887;
  assign n27889 = pi29  & n27888;
  assign n27890 = ~pi29  & ~n27888;
  assign n27891 = ~n27889 & ~n27890;
  assign n27892 = n27881 & ~n27891;
  assign n27893 = ~n27881 & n27891;
  assign n27894 = ~n27892 & ~n27893;
  assign n27895 = ~n27679 & n27690;
  assign n27896 = ~n27678 & ~n27895;
  assign n27897 = n27894 & n27896;
  assign n27898 = ~n27894 & ~n27896;
  assign n27899 = ~n27897 & ~n27898;
  assign n27900 = n4601 & n21204;
  assign n27901 = n4783 & n21201;
  assign n27902 = n4602 & n22832;
  assign n27903 = n4801 & n21198;
  assign n27904 = ~n27902 & ~n27903;
  assign n27905 = ~n27901 & n27904;
  assign n27906 = ~n27900 & n27905;
  assign n27907 = pi26  & n27906;
  assign n27908 = ~pi26  & ~n27906;
  assign n27909 = ~n27907 & ~n27908;
  assign n27910 = n27899 & ~n27909;
  assign n27911 = ~n27899 & n27909;
  assign n27912 = ~n27910 & ~n27911;
  assign n27913 = n27832 & ~n27912;
  assign n27914 = ~n27832 & n27912;
  assign n27915 = ~n27913 & ~n27914;
  assign n27916 = n5238 & n21195;
  assign n27917 = n71 & n21192;
  assign n27918 = n5239 & n23399;
  assign n27919 = n5326 & n21189;
  assign n27920 = ~n27918 & ~n27919;
  assign n27921 = ~n27917 & n27920;
  assign n27922 = ~n27916 & n27921;
  assign n27923 = pi23  & n27922;
  assign n27924 = ~pi23  & ~n27922;
  assign n27925 = ~n27923 & ~n27924;
  assign n27926 = n27915 & ~n27925;
  assign n27927 = ~n27915 & n27925;
  assign n27928 = ~n27926 & ~n27927;
  assign n27929 = n27831 & ~n27928;
  assign n27930 = ~n27831 & n27928;
  assign n27931 = ~n27929 & ~n27930;
  assign n27932 = n5435 & n21186;
  assign n27933 = n6055 & n21183;
  assign n27934 = n5429 & n23991;
  assign n27935 = n6071 & n21180;
  assign n27936 = ~n27934 & ~n27935;
  assign n27937 = ~n27933 & n27936;
  assign n27938 = ~n27932 & n27937;
  assign n27939 = pi20  & n27938;
  assign n27940 = ~pi20  & ~n27938;
  assign n27941 = ~n27939 & ~n27940;
  assign n27942 = n27931 & ~n27941;
  assign n27943 = ~n27931 & n27941;
  assign n27944 = ~n27942 & ~n27943;
  assign n27945 = n27829 & ~n27944;
  assign n27946 = ~n27829 & n27944;
  assign n27947 = ~n27945 & ~n27946;
  assign n27948 = n6184 & n21076;
  assign n27949 = n6527 & n21176;
  assign n27950 = n6185 & ~n21470;
  assign n27951 = n6543 & n21464;
  assign n27952 = ~n27950 & ~n27951;
  assign n27953 = ~n27949 & n27952;
  assign n27954 = ~n27948 & n27953;
  assign n27955 = pi17  & n27954;
  assign n27956 = ~pi17  & ~n27954;
  assign n27957 = ~n27955 & ~n27956;
  assign n27958 = n27947 & ~n27957;
  assign n27959 = ~n27947 & n27957;
  assign n27960 = ~n27958 & ~n27959;
  assign n27961 = n27827 & ~n27960;
  assign n27962 = ~n27827 & n27960;
  assign n27963 = ~n27961 & ~n27962;
  assign n27964 = n6835 & n24607;
  assign n27965 = n7460 & n24676;
  assign n27966 = n6836 & ~n24754;
  assign n27967 = n7487 & n24748;
  assign n27968 = ~n27966 & ~n27967;
  assign n27969 = ~n27965 & n27968;
  assign n27970 = ~n27964 & n27969;
  assign n27971 = pi14  & n27970;
  assign n27972 = ~pi14  & ~n27970;
  assign n27973 = ~n27971 & ~n27972;
  assign n27974 = n27963 & ~n27973;
  assign n27975 = ~n27963 & n27973;
  assign n27976 = ~n27974 & ~n27975;
  assign n27977 = n27825 & n27976;
  assign n27978 = ~n27825 & ~n27976;
  assign n27979 = ~n27977 & ~n27978;
  assign n27980 = n7654 & n25521;
  assign n27981 = n8091 & n25785;
  assign n27982 = n7648 & n26049;
  assign n27983 = n8120 & n26043;
  assign n27984 = ~n27982 & ~n27983;
  assign n27985 = ~n27981 & n27984;
  assign n27986 = ~n27980 & n27985;
  assign n27987 = pi11  & n27986;
  assign n27988 = ~pi11  & ~n27986;
  assign n27989 = ~n27987 & ~n27988;
  assign n27990 = ~n27979 & ~n27989;
  assign n27991 = n27979 & n27989;
  assign n27992 = ~n27990 & ~n27991;
  assign n27993 = n27823 & ~n27992;
  assign n27994 = ~n27823 & n27992;
  assign n27995 = ~n27993 & ~n27994;
  assign n27996 = n8474 & n26284;
  assign n27997 = n9238 & n26532;
  assign n27998 = n8468 & ~n26770;
  assign n27999 = n9265 & n26764;
  assign n28000 = ~n27998 & ~n27999;
  assign n28001 = ~n27997 & n28000;
  assign n28002 = ~n27996 & n28001;
  assign n28003 = pi8  & n28002;
  assign n28004 = ~pi8  & ~n28002;
  assign n28005 = ~n28003 & ~n28004;
  assign n28006 = n27995 & ~n28005;
  assign n28007 = ~n27995 & n28005;
  assign n28008 = ~n28006 & ~n28007;
  assign n28009 = ~n27821 & n28008;
  assign n28010 = n27821 & ~n28008;
  assign n28011 = ~n28009 & ~n28010;
  assign n28012 = n27819 & ~n28011;
  assign n28013 = ~n27819 & n28011;
  assign n28014 = ~n28012 & ~n28013;
  assign n28015 = n27817 & n28014;
  assign n28016 = ~n27817 & ~n28014;
  assign po11  = ~n28015 & ~n28016;
  assign n28018 = ~n27825 & n27976;
  assign n28019 = ~n27990 & ~n28018;
  assign n28020 = n8468 & n26987;
  assign n28021 = n8474 & n26532;
  assign n28022 = n16606 & n26764;
  assign n28023 = ~n28021 & ~n28022;
  assign n28024 = ~n28020 & n28023;
  assign n28025 = pi8  & n28024;
  assign n28026 = ~pi8  & ~n28024;
  assign n28027 = ~n28025 & ~n28026;
  assign n28028 = ~n28019 & ~n28027;
  assign n28029 = n28019 & n28027;
  assign n28030 = ~n28028 & ~n28029;
  assign n28031 = ~n27880 & ~n27892;
  assign n28032 = ~n685 & n3836;
  assign n28033 = ~n361 & n28032;
  assign n28034 = ~n545 & n28033;
  assign n28035 = n1778 & n3158;
  assign n28036 = n3138 & n28035;
  assign n28037 = n5105 & n28036;
  assign n28038 = ~n475 & n28037;
  assign n28039 = n519 & n1791;
  assign n28040 = ~n535 & n28039;
  assign n28041 = n28038 & n28040;
  assign n28042 = n3125 & n28041;
  assign n28043 = n28034 & n28042;
  assign n28044 = ~n611 & n28043;
  assign n28045 = ~n458 & n28044;
  assign n28046 = ~n134 & ~n430;
  assign n28047 = ~n275 & n28046;
  assign n28048 = ~n345 & ~n668;
  assign n28049 = n28047 & n28048;
  assign n28050 = ~n692 & n28049;
  assign n28051 = ~n239 & ~n501;
  assign n28052 = ~n382 & n28051;
  assign n28053 = n28050 & n28052;
  assign n28054 = n4339 & n28053;
  assign n28055 = ~n422 & n28054;
  assign n28056 = ~n325 & n28055;
  assign n28057 = n28045 & n28056;
  assign n28058 = n12878 & n13136;
  assign n28059 = ~n427 & n28058;
  assign n28060 = ~n350 & n28059;
  assign n28061 = n4283 & n7103;
  assign n28062 = ~n383 & n28061;
  assign n28063 = ~n582 & n28062;
  assign n28064 = n28060 & n28063;
  assign n28065 = n28057 & n28064;
  assign n28066 = ~n27865 & n28065;
  assign n28067 = n27865 & ~n28065;
  assign n28068 = ~n28066 & ~n28067;
  assign n28069 = ~n27866 & n27875;
  assign n28070 = ~n27867 & ~n28069;
  assign n28071 = n28068 & ~n28070;
  assign n28072 = ~n28068 & n28070;
  assign n28073 = ~n28071 & ~n28072;
  assign n28074 = n3641 & n21219;
  assign n28075 = n3740 & n21216;
  assign n28076 = n556 & n22394;
  assign n28077 = n3961 & n21213;
  assign n28078 = ~n28076 & ~n28077;
  assign n28079 = ~n28075 & n28078;
  assign n28080 = ~n28074 & n28079;
  assign n28081 = ~n28073 & ~n28080;
  assign n28082 = n28073 & n28080;
  assign n28083 = ~n28081 & ~n28082;
  assign n28084 = n28031 & ~n28083;
  assign n28085 = ~n28031 & n28083;
  assign n28086 = ~n28084 & ~n28085;
  assign n28087 = n4006 & n21210;
  assign n28088 = n4133 & n21207;
  assign n28089 = n4002 & n22810;
  assign n28090 = n4555 & n21204;
  assign n28091 = ~n28089 & ~n28090;
  assign n28092 = ~n28088 & n28091;
  assign n28093 = ~n28087 & n28092;
  assign n28094 = pi29  & n28093;
  assign n28095 = ~pi29  & ~n28093;
  assign n28096 = ~n28094 & ~n28095;
  assign n28097 = n28086 & n28096;
  assign n28098 = ~n28086 & ~n28096;
  assign n28099 = ~n28097 & ~n28098;
  assign n28100 = n4601 & n21201;
  assign n28101 = n4783 & n21198;
  assign n28102 = n4602 & n21482;
  assign n28103 = n4801 & n21195;
  assign n28104 = ~n28102 & ~n28103;
  assign n28105 = ~n28101 & n28104;
  assign n28106 = ~n28100 & n28105;
  assign n28107 = pi26  & n28106;
  assign n28108 = ~pi26  & ~n28106;
  assign n28109 = ~n28107 & ~n28108;
  assign n28110 = ~n28099 & ~n28109;
  assign n28111 = n28099 & n28109;
  assign n28112 = ~n28110 & ~n28111;
  assign n28113 = ~n27897 & n27909;
  assign n28114 = ~n27898 & ~n28113;
  assign n28115 = ~n28112 & ~n28114;
  assign n28116 = n28112 & n28114;
  assign n28117 = ~n28115 & ~n28116;
  assign n28118 = n5238 & n21192;
  assign n28119 = n71 & n21189;
  assign n28120 = n5239 & n23384;
  assign n28121 = n5326 & n21186;
  assign n28122 = ~n28120 & ~n28121;
  assign n28123 = ~n28119 & n28122;
  assign n28124 = ~n28118 & n28123;
  assign n28125 = pi23  & n28124;
  assign n28126 = ~pi23  & ~n28124;
  assign n28127 = ~n28125 & ~n28126;
  assign n28128 = n28117 & ~n28127;
  assign n28129 = ~n28117 & n28127;
  assign n28130 = ~n28128 & ~n28129;
  assign n28131 = ~n27914 & n27925;
  assign n28132 = ~n27913 & ~n28131;
  assign n28133 = ~n28130 & ~n28132;
  assign n28134 = n28130 & n28132;
  assign n28135 = ~n28133 & ~n28134;
  assign n28136 = n5435 & n21183;
  assign n28137 = n6055 & n21180;
  assign n28138 = n5429 & n24030;
  assign n28139 = n6071 & n21076;
  assign n28140 = ~n28138 & ~n28139;
  assign n28141 = ~n28137 & n28140;
  assign n28142 = ~n28136 & n28141;
  assign n28143 = pi20  & n28142;
  assign n28144 = ~pi20  & ~n28142;
  assign n28145 = ~n28143 & ~n28144;
  assign n28146 = n28135 & ~n28145;
  assign n28147 = ~n28135 & n28145;
  assign n28148 = ~n28146 & ~n28147;
  assign n28149 = ~n27930 & n27941;
  assign n28150 = ~n27929 & ~n28149;
  assign n28151 = ~n28148 & ~n28150;
  assign n28152 = n28148 & n28150;
  assign n28153 = ~n28151 & ~n28152;
  assign n28154 = n6184 & n21176;
  assign n28155 = n6527 & n21464;
  assign n28156 = n6185 & n24782;
  assign n28157 = n6543 & n24607;
  assign n28158 = ~n28156 & ~n28157;
  assign n28159 = ~n28155 & n28158;
  assign n28160 = ~n28154 & n28159;
  assign n28161 = pi17  & n28160;
  assign n28162 = ~pi17  & ~n28160;
  assign n28163 = ~n28161 & ~n28162;
  assign n28164 = n28153 & ~n28163;
  assign n28165 = ~n28153 & n28163;
  assign n28166 = ~n28164 & ~n28165;
  assign n28167 = ~n27946 & n27957;
  assign n28168 = ~n27945 & ~n28167;
  assign n28169 = ~n28166 & ~n28168;
  assign n28170 = n28166 & n28168;
  assign n28171 = ~n28169 & ~n28170;
  assign n28172 = n6835 & n24676;
  assign n28173 = n7460 & n24748;
  assign n28174 = n6836 & ~n25529;
  assign n28175 = n7487 & n25521;
  assign n28176 = ~n28174 & ~n28175;
  assign n28177 = ~n28173 & n28176;
  assign n28178 = ~n28172 & n28177;
  assign n28179 = pi14  & n28178;
  assign n28180 = ~pi14  & ~n28178;
  assign n28181 = ~n28179 & ~n28180;
  assign n28182 = n28171 & ~n28181;
  assign n28183 = ~n28171 & n28181;
  assign n28184 = ~n28182 & ~n28183;
  assign n28185 = ~n27962 & n27973;
  assign n28186 = ~n27961 & ~n28185;
  assign n28187 = ~n28184 & ~n28186;
  assign n28188 = n28184 & n28186;
  assign n28189 = ~n28187 & ~n28188;
  assign n28190 = n7654 & n25785;
  assign n28191 = n8091 & n26043;
  assign n28192 = n7648 & ~n26290;
  assign n28193 = n8120 & n26284;
  assign n28194 = ~n28192 & ~n28193;
  assign n28195 = ~n28191 & n28194;
  assign n28196 = ~n28190 & n28195;
  assign n28197 = pi11  & n28196;
  assign n28198 = ~pi11  & ~n28196;
  assign n28199 = ~n28197 & ~n28198;
  assign n28200 = n28189 & ~n28199;
  assign n28201 = ~n28189 & n28199;
  assign n28202 = ~n28200 & ~n28201;
  assign n28203 = n28030 & n28202;
  assign n28204 = ~n28030 & ~n28202;
  assign n28205 = ~n28203 & ~n28204;
  assign n28206 = ~n27994 & n28005;
  assign n28207 = ~n27993 & ~n28206;
  assign n28208 = ~n28205 & ~n28207;
  assign n28209 = n28205 & n28207;
  assign n28210 = ~n28208 & ~n28209;
  assign n28211 = ~n28009 & ~n28013;
  assign n28212 = ~n28210 & n28211;
  assign n28213 = n28210 & ~n28211;
  assign n28214 = ~n28212 & ~n28213;
  assign n28215 = n28015 & n28214;
  assign n28216 = ~n28015 & ~n28214;
  assign po12  = ~n28215 & ~n28216;
  assign n28218 = ~n28209 & ~n28213;
  assign n28219 = ~n28081 & ~n28085;
  assign n28220 = n4006 & n21207;
  assign n28221 = n4133 & n21204;
  assign n28222 = n4002 & n22852;
  assign n28223 = n4555 & n21201;
  assign n28224 = ~n28222 & ~n28223;
  assign n28225 = ~n28221 & n28224;
  assign n28226 = ~n28220 & n28225;
  assign n28227 = pi29  & n28226;
  assign n28228 = ~pi29  & ~n28226;
  assign n28229 = ~n28227 & ~n28228;
  assign n28230 = ~n13915 & n26764;
  assign n28231 = pi8  & ~n28230;
  assign n28232 = ~pi8  & n28230;
  assign n28233 = ~n28231 & ~n28232;
  assign n28234 = n910 & n2779;
  assign n28235 = n1872 & n28234;
  assign n28236 = n167 & n28235;
  assign n28237 = n2242 & n2409;
  assign n28238 = n1316 & n28237;
  assign n28239 = ~n326 & n28238;
  assign n28240 = n28236 & n28239;
  assign n28241 = n1353 & n3495;
  assign n28242 = n1057 & n28241;
  assign n28243 = n1134 & n13081;
  assign n28244 = n3215 & n28243;
  assign n28245 = ~n700 & n28244;
  assign n28246 = n28242 & n28245;
  assign n28247 = n28240 & n28246;
  assign n28248 = n27865 & n28247;
  assign n28249 = ~n27865 & ~n28247;
  assign n28250 = ~n28248 & ~n28249;
  assign n28251 = n28233 & n28250;
  assign n28252 = ~n28233 & ~n28250;
  assign n28253 = ~n28251 & ~n28252;
  assign n28254 = ~n28067 & ~n28070;
  assign n28255 = ~n28066 & ~n28254;
  assign n28256 = n28253 & n28255;
  assign n28257 = ~n28253 & ~n28255;
  assign n28258 = ~n28256 & ~n28257;
  assign n28259 = n3641 & n21216;
  assign n28260 = n3740 & n21213;
  assign n28261 = n556 & n22376;
  assign n28262 = n3961 & n21210;
  assign n28263 = ~n28261 & ~n28262;
  assign n28264 = ~n28260 & n28263;
  assign n28265 = ~n28259 & n28264;
  assign n28266 = n28258 & ~n28265;
  assign n28267 = ~n28258 & n28265;
  assign n28268 = ~n28266 & ~n28267;
  assign n28269 = ~n28229 & n28268;
  assign n28270 = n28229 & ~n28268;
  assign n28271 = ~n28269 & ~n28270;
  assign n28272 = n28219 & ~n28271;
  assign n28273 = ~n28219 & n28271;
  assign n28274 = ~n28272 & ~n28273;
  assign n28275 = n4601 & n21198;
  assign n28276 = n4783 & n21195;
  assign n28277 = n4602 & n23211;
  assign n28278 = n4801 & n21192;
  assign n28279 = ~n28277 & ~n28278;
  assign n28280 = ~n28276 & n28279;
  assign n28281 = ~n28275 & n28280;
  assign n28282 = pi26  & n28281;
  assign n28283 = ~pi26  & ~n28281;
  assign n28284 = ~n28282 & ~n28283;
  assign n28285 = n28274 & n28284;
  assign n28286 = ~n28274 & ~n28284;
  assign n28287 = ~n28285 & ~n28286;
  assign n28288 = n28086 & ~n28096;
  assign n28289 = ~n28110 & ~n28288;
  assign n28290 = n28287 & n28289;
  assign n28291 = ~n28287 & ~n28289;
  assign n28292 = ~n28290 & ~n28291;
  assign n28293 = n5238 & n21189;
  assign n28294 = n71 & n21186;
  assign n28295 = n5239 & n23369;
  assign n28296 = n5326 & n21183;
  assign n28297 = ~n28295 & ~n28296;
  assign n28298 = ~n28294 & n28297;
  assign n28299 = ~n28293 & n28298;
  assign n28300 = pi23  & n28299;
  assign n28301 = ~pi23  & ~n28299;
  assign n28302 = ~n28300 & ~n28301;
  assign n28303 = n28292 & n28302;
  assign n28304 = ~n28292 & ~n28302;
  assign n28305 = ~n28303 & ~n28304;
  assign n28306 = ~n28116 & n28127;
  assign n28307 = ~n28115 & ~n28306;
  assign n28308 = n28305 & ~n28307;
  assign n28309 = ~n28305 & n28307;
  assign n28310 = ~n28308 & ~n28309;
  assign n28311 = n5435 & n21180;
  assign n28312 = n6055 & n21076;
  assign n28313 = n5429 & n24012;
  assign n28314 = n6071 & n21176;
  assign n28315 = ~n28313 & ~n28314;
  assign n28316 = ~n28312 & n28315;
  assign n28317 = ~n28311 & n28316;
  assign n28318 = pi20  & n28317;
  assign n28319 = ~pi20  & ~n28317;
  assign n28320 = ~n28318 & ~n28319;
  assign n28321 = n28310 & n28320;
  assign n28322 = ~n28310 & ~n28320;
  assign n28323 = ~n28321 & ~n28322;
  assign n28324 = ~n28134 & n28145;
  assign n28325 = ~n28133 & ~n28324;
  assign n28326 = n28323 & ~n28325;
  assign n28327 = ~n28323 & n28325;
  assign n28328 = ~n28326 & ~n28327;
  assign n28329 = n6184 & n21464;
  assign n28330 = n6527 & n24607;
  assign n28331 = n6185 & n24770;
  assign n28332 = n6543 & n24676;
  assign n28333 = ~n28331 & ~n28332;
  assign n28334 = ~n28330 & n28333;
  assign n28335 = ~n28329 & n28334;
  assign n28336 = pi17  & n28335;
  assign n28337 = ~pi17  & ~n28335;
  assign n28338 = ~n28336 & ~n28337;
  assign n28339 = ~n28152 & n28163;
  assign n28340 = ~n28151 & ~n28339;
  assign n28341 = n28338 & n28340;
  assign n28342 = ~n28338 & ~n28340;
  assign n28343 = ~n28341 & ~n28342;
  assign n28344 = ~n28328 & n28343;
  assign n28345 = n28328 & ~n28343;
  assign n28346 = ~n28344 & ~n28345;
  assign n28347 = n6835 & n24748;
  assign n28348 = n7460 & n25521;
  assign n28349 = n6836 & n25793;
  assign n28350 = n7487 & n25785;
  assign n28351 = ~n28349 & ~n28350;
  assign n28352 = ~n28348 & n28351;
  assign n28353 = ~n28347 & n28352;
  assign n28354 = pi14  & n28353;
  assign n28355 = ~pi14  & ~n28353;
  assign n28356 = ~n28354 & ~n28355;
  assign n28357 = n28346 & n28356;
  assign n28358 = ~n28346 & ~n28356;
  assign n28359 = ~n28357 & ~n28358;
  assign n28360 = ~n28170 & n28181;
  assign n28361 = ~n28169 & ~n28360;
  assign n28362 = n28359 & ~n28361;
  assign n28363 = ~n28359 & n28361;
  assign n28364 = ~n28362 & ~n28363;
  assign n28365 = n7654 & n26043;
  assign n28366 = n8091 & n26284;
  assign n28367 = n7648 & n26540;
  assign n28368 = n8120 & n26532;
  assign n28369 = ~n28367 & ~n28368;
  assign n28370 = ~n28366 & n28369;
  assign n28371 = ~n28365 & n28370;
  assign n28372 = pi11  & n28371;
  assign n28373 = ~pi11  & ~n28371;
  assign n28374 = ~n28372 & ~n28373;
  assign n28375 = ~n28188 & n28199;
  assign n28376 = ~n28187 & ~n28375;
  assign n28377 = n28374 & n28376;
  assign n28378 = ~n28374 & ~n28376;
  assign n28379 = ~n28377 & ~n28378;
  assign n28380 = ~n28364 & n28379;
  assign n28381 = n28364 & ~n28379;
  assign n28382 = ~n28380 & ~n28381;
  assign n28383 = ~n28028 & ~n28202;
  assign n28384 = ~n28029 & ~n28383;
  assign n28385 = n28382 & n28384;
  assign n28386 = ~n28382 & ~n28384;
  assign n28387 = ~n28385 & ~n28386;
  assign n28388 = ~n28218 & n28387;
  assign n28389 = n28218 & ~n28387;
  assign n28390 = ~n28388 & ~n28389;
  assign n28391 = ~n28215 & ~n28390;
  assign n28392 = n28215 & n28390;
  assign po13  = ~n28391 & ~n28392;
  assign n28394 = ~n28385 & ~n28388;
  assign n28395 = ~n28374 & n28376;
  assign n28396 = ~n28381 & ~n28395;
  assign n28397 = n28346 & ~n28356;
  assign n28398 = ~n28363 & ~n28397;
  assign n28399 = ~n28338 & n28340;
  assign n28400 = ~n28345 & ~n28399;
  assign n28401 = n28310 & ~n28320;
  assign n28402 = ~n28327 & ~n28401;
  assign n28403 = n28292 & ~n28302;
  assign n28404 = ~n28309 & ~n28403;
  assign n28405 = n28274 & ~n28284;
  assign n28406 = ~n28291 & ~n28405;
  assign n28407 = ~n28269 & ~n28273;
  assign n28408 = ~n28249 & ~n28251;
  assign n28409 = n3282 & n5488;
  assign n28410 = ~n166 & n28409;
  assign n28411 = n3820 & n13741;
  assign n28412 = n2533 & n28411;
  assign n28413 = ~n206 & n28412;
  assign n28414 = ~n668 & n28413;
  assign n28415 = n28410 & n28414;
  assign n28416 = n909 & n15123;
  assign n28417 = ~n548 & n28416;
  assign n28418 = ~n81 & n28417;
  assign n28419 = n1029 & n2301;
  assign n28420 = ~n588 & n28419;
  assign n28421 = ~n261 & n28420;
  assign n28422 = n28418 & n28421;
  assign n28423 = n28415 & n28422;
  assign n28424 = ~n28408 & n28423;
  assign n28425 = n28408 & ~n28423;
  assign n28426 = ~n28424 & ~n28425;
  assign n28427 = n3641 & n21213;
  assign n28428 = n3740 & n21210;
  assign n28429 = n556 & n22363;
  assign n28430 = n3961 & n21207;
  assign n28431 = ~n28429 & ~n28430;
  assign n28432 = ~n28428 & n28431;
  assign n28433 = ~n28427 & n28432;
  assign n28434 = n28426 & ~n28433;
  assign n28435 = ~n28426 & n28433;
  assign n28436 = ~n28434 & ~n28435;
  assign n28437 = ~n28256 & n28265;
  assign n28438 = ~n28257 & ~n28437;
  assign n28439 = ~n28436 & ~n28438;
  assign n28440 = n28436 & n28438;
  assign n28441 = ~n28439 & ~n28440;
  assign n28442 = n4006 & n21204;
  assign n28443 = n4133 & n21201;
  assign n28444 = n4002 & n22832;
  assign n28445 = n4555 & n21198;
  assign n28446 = ~n28444 & ~n28445;
  assign n28447 = ~n28443 & n28446;
  assign n28448 = ~n28442 & n28447;
  assign n28449 = pi29  & n28448;
  assign n28450 = ~pi29  & ~n28448;
  assign n28451 = ~n28449 & ~n28450;
  assign n28452 = n28441 & ~n28451;
  assign n28453 = ~n28441 & n28451;
  assign n28454 = ~n28452 & ~n28453;
  assign n28455 = ~n28407 & n28454;
  assign n28456 = n28407 & ~n28454;
  assign n28457 = ~n28455 & ~n28456;
  assign n28458 = n4601 & n21195;
  assign n28459 = n4783 & n21192;
  assign n28460 = n4602 & n23399;
  assign n28461 = n4801 & n21189;
  assign n28462 = ~n28460 & ~n28461;
  assign n28463 = ~n28459 & n28462;
  assign n28464 = ~n28458 & n28463;
  assign n28465 = pi26  & n28464;
  assign n28466 = ~pi26  & ~n28464;
  assign n28467 = ~n28465 & ~n28466;
  assign n28468 = n28457 & ~n28467;
  assign n28469 = ~n28457 & n28467;
  assign n28470 = ~n28468 & ~n28469;
  assign n28471 = n28406 & ~n28470;
  assign n28472 = ~n28406 & n28470;
  assign n28473 = ~n28471 & ~n28472;
  assign n28474 = n5238 & n21186;
  assign n28475 = n71 & n21183;
  assign n28476 = n5239 & n23991;
  assign n28477 = n5326 & n21180;
  assign n28478 = ~n28476 & ~n28477;
  assign n28479 = ~n28475 & n28478;
  assign n28480 = ~n28474 & n28479;
  assign n28481 = pi23  & n28480;
  assign n28482 = ~pi23  & ~n28480;
  assign n28483 = ~n28481 & ~n28482;
  assign n28484 = n28473 & ~n28483;
  assign n28485 = ~n28473 & n28483;
  assign n28486 = ~n28484 & ~n28485;
  assign n28487 = n28404 & ~n28486;
  assign n28488 = ~n28404 & n28486;
  assign n28489 = ~n28487 & ~n28488;
  assign n28490 = n5435 & n21076;
  assign n28491 = n6055 & n21176;
  assign n28492 = n5429 & ~n21470;
  assign n28493 = n6071 & n21464;
  assign n28494 = ~n28492 & ~n28493;
  assign n28495 = ~n28491 & n28494;
  assign n28496 = ~n28490 & n28495;
  assign n28497 = pi20  & n28496;
  assign n28498 = ~pi20  & ~n28496;
  assign n28499 = ~n28497 & ~n28498;
  assign n28500 = n28489 & ~n28499;
  assign n28501 = ~n28489 & n28499;
  assign n28502 = ~n28500 & ~n28501;
  assign n28503 = n28402 & ~n28502;
  assign n28504 = ~n28402 & n28502;
  assign n28505 = ~n28503 & ~n28504;
  assign n28506 = n6184 & n24607;
  assign n28507 = n6527 & n24676;
  assign n28508 = n6185 & ~n24754;
  assign n28509 = n6543 & n24748;
  assign n28510 = ~n28508 & ~n28509;
  assign n28511 = ~n28507 & n28510;
  assign n28512 = ~n28506 & n28511;
  assign n28513 = pi17  & n28512;
  assign n28514 = ~pi17  & ~n28512;
  assign n28515 = ~n28513 & ~n28514;
  assign n28516 = n28505 & ~n28515;
  assign n28517 = ~n28505 & n28515;
  assign n28518 = ~n28516 & ~n28517;
  assign n28519 = n28400 & n28518;
  assign n28520 = ~n28400 & ~n28518;
  assign n28521 = ~n28519 & ~n28520;
  assign n28522 = n6835 & n25521;
  assign n28523 = n7460 & n25785;
  assign n28524 = n6836 & n26049;
  assign n28525 = n7487 & n26043;
  assign n28526 = ~n28524 & ~n28525;
  assign n28527 = ~n28523 & n28526;
  assign n28528 = ~n28522 & n28527;
  assign n28529 = pi14  & n28528;
  assign n28530 = ~pi14  & ~n28528;
  assign n28531 = ~n28529 & ~n28530;
  assign n28532 = ~n28521 & ~n28531;
  assign n28533 = n28521 & n28531;
  assign n28534 = ~n28532 & ~n28533;
  assign n28535 = n28398 & ~n28534;
  assign n28536 = ~n28398 & n28534;
  assign n28537 = ~n28535 & ~n28536;
  assign n28538 = n7654 & n26284;
  assign n28539 = n8091 & n26532;
  assign n28540 = n7648 & ~n26770;
  assign n28541 = n8120 & n26764;
  assign n28542 = ~n28540 & ~n28541;
  assign n28543 = ~n28539 & n28542;
  assign n28544 = ~n28538 & n28543;
  assign n28545 = pi11  & n28544;
  assign n28546 = ~pi11  & ~n28544;
  assign n28547 = ~n28545 & ~n28546;
  assign n28548 = n28537 & ~n28547;
  assign n28549 = ~n28537 & n28547;
  assign n28550 = ~n28548 & ~n28549;
  assign n28551 = ~n28396 & n28550;
  assign n28552 = n28396 & ~n28550;
  assign n28553 = ~n28551 & ~n28552;
  assign n28554 = n28394 & ~n28553;
  assign n28555 = ~n28394 & n28553;
  assign n28556 = ~n28554 & ~n28555;
  assign n28557 = n28392 & n28556;
  assign n28558 = ~n28392 & ~n28556;
  assign po14  = ~n28557 & ~n28558;
  assign n28560 = ~n28400 & n28518;
  assign n28561 = ~n28532 & ~n28560;
  assign n28562 = n7648 & n26987;
  assign n28563 = n7654 & n26532;
  assign n28564 = n15692 & n26764;
  assign n28565 = ~n28563 & ~n28564;
  assign n28566 = ~n28562 & n28565;
  assign n28567 = pi11  & n28566;
  assign n28568 = ~pi11  & ~n28566;
  assign n28569 = ~n28567 & ~n28568;
  assign n28570 = ~n28561 & ~n28569;
  assign n28571 = n28561 & n28569;
  assign n28572 = ~n28570 & ~n28571;
  assign n28573 = ~n28440 & ~n28452;
  assign n28574 = n4006 & n21201;
  assign n28575 = n4133 & n21198;
  assign n28576 = n4002 & n21482;
  assign n28577 = n4555 & n21195;
  assign n28578 = ~n28576 & ~n28577;
  assign n28579 = ~n28575 & n28578;
  assign n28580 = ~n28574 & n28579;
  assign n28581 = pi29  & n28580;
  assign n28582 = ~pi29  & ~n28580;
  assign n28583 = ~n28581 & ~n28582;
  assign n28584 = n1148 & n3454;
  assign n28585 = n974 & n28584;
  assign n28586 = n1079 & n28585;
  assign n28587 = ~n252 & n28586;
  assign n28588 = n1012 & n14619;
  assign n28589 = n2064 & n28588;
  assign n28590 = ~n131 & n28589;
  assign n28591 = n28587 & n28590;
  assign n28592 = n3388 & n5934;
  assign n28593 = n1708 & n28592;
  assign n28594 = ~n598 & n28593;
  assign n28595 = n1742 & n13107;
  assign n28596 = n1830 & n28595;
  assign n28597 = n27849 & n28596;
  assign n28598 = ~n534 & n28597;
  assign n28599 = ~n323 & n28598;
  assign n28600 = n28594 & n28599;
  assign n28601 = n28591 & n28600;
  assign n28602 = ~n28423 & n28601;
  assign n28603 = n28423 & ~n28601;
  assign n28604 = ~n28602 & ~n28603;
  assign n28605 = ~n28424 & n28433;
  assign n28606 = ~n28425 & ~n28605;
  assign n28607 = n28604 & ~n28606;
  assign n28608 = ~n28604 & n28606;
  assign n28609 = ~n28607 & ~n28608;
  assign n28610 = n3641 & n21210;
  assign n28611 = n3740 & n21207;
  assign n28612 = n556 & n22810;
  assign n28613 = n3961 & n21204;
  assign n28614 = ~n28612 & ~n28613;
  assign n28615 = ~n28611 & n28614;
  assign n28616 = ~n28610 & n28615;
  assign n28617 = ~n28609 & ~n28616;
  assign n28618 = n28609 & n28616;
  assign n28619 = ~n28617 & ~n28618;
  assign n28620 = ~n28583 & n28619;
  assign n28621 = n28583 & ~n28619;
  assign n28622 = ~n28620 & ~n28621;
  assign n28623 = ~n28573 & n28622;
  assign n28624 = n28573 & ~n28622;
  assign n28625 = ~n28623 & ~n28624;
  assign n28626 = n4601 & n21192;
  assign n28627 = n4783 & n21189;
  assign n28628 = n4602 & n23384;
  assign n28629 = n4801 & n21186;
  assign n28630 = ~n28628 & ~n28629;
  assign n28631 = ~n28627 & n28630;
  assign n28632 = ~n28626 & n28631;
  assign n28633 = pi26  & n28632;
  assign n28634 = ~pi26  & ~n28632;
  assign n28635 = ~n28633 & ~n28634;
  assign n28636 = n28625 & ~n28635;
  assign n28637 = ~n28625 & n28635;
  assign n28638 = ~n28636 & ~n28637;
  assign n28639 = ~n28455 & n28467;
  assign n28640 = ~n28456 & ~n28639;
  assign n28641 = ~n28638 & ~n28640;
  assign n28642 = n28638 & n28640;
  assign n28643 = ~n28641 & ~n28642;
  assign n28644 = n5238 & n21183;
  assign n28645 = n71 & n21180;
  assign n28646 = n5239 & n24030;
  assign n28647 = n5326 & n21076;
  assign n28648 = ~n28646 & ~n28647;
  assign n28649 = ~n28645 & n28648;
  assign n28650 = ~n28644 & n28649;
  assign n28651 = pi23  & n28650;
  assign n28652 = ~pi23  & ~n28650;
  assign n28653 = ~n28651 & ~n28652;
  assign n28654 = n28643 & ~n28653;
  assign n28655 = ~n28643 & n28653;
  assign n28656 = ~n28654 & ~n28655;
  assign n28657 = ~n28472 & n28483;
  assign n28658 = ~n28471 & ~n28657;
  assign n28659 = ~n28656 & ~n28658;
  assign n28660 = n28656 & n28658;
  assign n28661 = ~n28659 & ~n28660;
  assign n28662 = n5435 & n21176;
  assign n28663 = n6055 & n21464;
  assign n28664 = n5429 & n24782;
  assign n28665 = n6071 & n24607;
  assign n28666 = ~n28664 & ~n28665;
  assign n28667 = ~n28663 & n28666;
  assign n28668 = ~n28662 & n28667;
  assign n28669 = pi20  & n28668;
  assign n28670 = ~pi20  & ~n28668;
  assign n28671 = ~n28669 & ~n28670;
  assign n28672 = n28661 & ~n28671;
  assign n28673 = ~n28661 & n28671;
  assign n28674 = ~n28672 & ~n28673;
  assign n28675 = ~n28488 & n28499;
  assign n28676 = ~n28487 & ~n28675;
  assign n28677 = ~n28674 & ~n28676;
  assign n28678 = n28674 & n28676;
  assign n28679 = ~n28677 & ~n28678;
  assign n28680 = n6184 & n24676;
  assign n28681 = n6527 & n24748;
  assign n28682 = n6185 & ~n25529;
  assign n28683 = n6543 & n25521;
  assign n28684 = ~n28682 & ~n28683;
  assign n28685 = ~n28681 & n28684;
  assign n28686 = ~n28680 & n28685;
  assign n28687 = pi17  & n28686;
  assign n28688 = ~pi17  & ~n28686;
  assign n28689 = ~n28687 & ~n28688;
  assign n28690 = n28679 & ~n28689;
  assign n28691 = ~n28679 & n28689;
  assign n28692 = ~n28690 & ~n28691;
  assign n28693 = ~n28504 & n28515;
  assign n28694 = ~n28503 & ~n28693;
  assign n28695 = ~n28692 & ~n28694;
  assign n28696 = n28692 & n28694;
  assign n28697 = ~n28695 & ~n28696;
  assign n28698 = n6835 & n25785;
  assign n28699 = n7460 & n26043;
  assign n28700 = n6836 & ~n26290;
  assign n28701 = n7487 & n26284;
  assign n28702 = ~n28700 & ~n28701;
  assign n28703 = ~n28699 & n28702;
  assign n28704 = ~n28698 & n28703;
  assign n28705 = pi14  & n28704;
  assign n28706 = ~pi14  & ~n28704;
  assign n28707 = ~n28705 & ~n28706;
  assign n28708 = n28697 & ~n28707;
  assign n28709 = ~n28697 & n28707;
  assign n28710 = ~n28708 & ~n28709;
  assign n28711 = n28572 & n28710;
  assign n28712 = ~n28572 & ~n28710;
  assign n28713 = ~n28711 & ~n28712;
  assign n28714 = ~n28536 & n28547;
  assign n28715 = ~n28535 & ~n28714;
  assign n28716 = ~n28713 & ~n28715;
  assign n28717 = n28713 & n28715;
  assign n28718 = ~n28716 & ~n28717;
  assign n28719 = ~n28551 & ~n28555;
  assign n28720 = ~n28718 & n28719;
  assign n28721 = n28718 & ~n28719;
  assign n28722 = ~n28720 & ~n28721;
  assign n28723 = n28557 & n28722;
  assign n28724 = ~n28557 & ~n28722;
  assign po15  = ~n28723 & ~n28724;
  assign n28726 = ~n28717 & ~n28721;
  assign n28727 = n4601 & n21189;
  assign n28728 = n4783 & n21186;
  assign n28729 = n4602 & n23369;
  assign n28730 = n4801 & n21183;
  assign n28731 = ~n28729 & ~n28730;
  assign n28732 = ~n28728 & n28731;
  assign n28733 = ~n28727 & n28732;
  assign n28734 = pi26  & n28733;
  assign n28735 = ~pi26  & ~n28733;
  assign n28736 = ~n28734 & ~n28735;
  assign n28737 = n4006 & n21198;
  assign n28738 = n4133 & n21195;
  assign n28739 = n4002 & n23211;
  assign n28740 = n4555 & n21192;
  assign n28741 = ~n28739 & ~n28740;
  assign n28742 = ~n28738 & n28741;
  assign n28743 = ~n28737 & n28742;
  assign n28744 = pi29  & n28743;
  assign n28745 = ~pi29  & ~n28743;
  assign n28746 = ~n28744 & ~n28745;
  assign n28747 = ~n28617 & ~n28620;
  assign n28748 = ~n13750 & n26764;
  assign n28749 = pi11  & ~n28748;
  assign n28750 = ~pi11  & n28748;
  assign n28751 = ~n28749 & ~n28750;
  assign n28752 = n2203 & n2917;
  assign n28753 = ~n254 & n28752;
  assign n28754 = n2239 & n5682;
  assign n28755 = n765 & n28754;
  assign n28756 = ~n81 & n28755;
  assign n28757 = n28753 & n28756;
  assign n28758 = n1545 & n3442;
  assign n28759 = n1211 & n28758;
  assign n28760 = n1138 & n28759;
  assign n28761 = n2066 & n28760;
  assign n28762 = ~n350 & n28761;
  assign n28763 = n1348 & n5714;
  assign n28764 = n673 & n28763;
  assign n28765 = ~n219 & n28764;
  assign n28766 = n28762 & n28765;
  assign n28767 = n28757 & n28766;
  assign n28768 = n28423 & n28767;
  assign n28769 = ~n28423 & ~n28767;
  assign n28770 = ~n28768 & ~n28769;
  assign n28771 = n28751 & n28770;
  assign n28772 = ~n28751 & ~n28770;
  assign n28773 = ~n28771 & ~n28772;
  assign n28774 = n3641 & n21207;
  assign n28775 = n3740 & n21204;
  assign n28776 = n556 & n22852;
  assign n28777 = n3961 & n21201;
  assign n28778 = ~n28776 & ~n28777;
  assign n28779 = ~n28775 & n28778;
  assign n28780 = ~n28774 & n28779;
  assign n28781 = n28773 & n28780;
  assign n28782 = ~n28773 & ~n28780;
  assign n28783 = ~n28781 & ~n28782;
  assign n28784 = ~n28603 & ~n28606;
  assign n28785 = ~n28602 & ~n28784;
  assign n28786 = ~n28783 & n28785;
  assign n28787 = n28783 & ~n28785;
  assign n28788 = ~n28786 & ~n28787;
  assign n28789 = ~n28747 & n28788;
  assign n28790 = n28747 & ~n28788;
  assign n28791 = ~n28789 & ~n28790;
  assign n28792 = n28746 & ~n28791;
  assign n28793 = ~n28746 & n28791;
  assign n28794 = ~n28792 & ~n28793;
  assign n28795 = n28736 & n28794;
  assign n28796 = ~n28736 & ~n28794;
  assign n28797 = ~n28795 & ~n28796;
  assign n28798 = ~n28623 & n28635;
  assign n28799 = ~n28624 & ~n28798;
  assign n28800 = n28797 & ~n28799;
  assign n28801 = ~n28797 & n28799;
  assign n28802 = ~n28800 & ~n28801;
  assign n28803 = n5238 & n21180;
  assign n28804 = n71 & n21076;
  assign n28805 = n5239 & n24012;
  assign n28806 = n5326 & n21176;
  assign n28807 = ~n28805 & ~n28806;
  assign n28808 = ~n28804 & n28807;
  assign n28809 = ~n28803 & n28808;
  assign n28810 = pi23  & n28809;
  assign n28811 = ~pi23  & ~n28809;
  assign n28812 = ~n28810 & ~n28811;
  assign n28813 = n28802 & n28812;
  assign n28814 = ~n28802 & ~n28812;
  assign n28815 = ~n28813 & ~n28814;
  assign n28816 = ~n28642 & n28653;
  assign n28817 = ~n28641 & ~n28816;
  assign n28818 = n28815 & ~n28817;
  assign n28819 = ~n28815 & n28817;
  assign n28820 = ~n28818 & ~n28819;
  assign n28821 = n5435 & n21464;
  assign n28822 = n6055 & n24607;
  assign n28823 = n5429 & n24770;
  assign n28824 = n6071 & n24676;
  assign n28825 = ~n28823 & ~n28824;
  assign n28826 = ~n28822 & n28825;
  assign n28827 = ~n28821 & n28826;
  assign n28828 = pi20  & n28827;
  assign n28829 = ~pi20  & ~n28827;
  assign n28830 = ~n28828 & ~n28829;
  assign n28831 = ~n28660 & n28671;
  assign n28832 = ~n28659 & ~n28831;
  assign n28833 = n28830 & n28832;
  assign n28834 = ~n28830 & ~n28832;
  assign n28835 = ~n28833 & ~n28834;
  assign n28836 = ~n28820 & n28835;
  assign n28837 = n28820 & ~n28835;
  assign n28838 = ~n28836 & ~n28837;
  assign n28839 = n6184 & n24748;
  assign n28840 = n6527 & n25521;
  assign n28841 = n6185 & n25793;
  assign n28842 = n6543 & n25785;
  assign n28843 = ~n28841 & ~n28842;
  assign n28844 = ~n28840 & n28843;
  assign n28845 = ~n28839 & n28844;
  assign n28846 = pi17  & n28845;
  assign n28847 = ~pi17  & ~n28845;
  assign n28848 = ~n28846 & ~n28847;
  assign n28849 = n28838 & n28848;
  assign n28850 = ~n28838 & ~n28848;
  assign n28851 = ~n28849 & ~n28850;
  assign n28852 = ~n28678 & n28689;
  assign n28853 = ~n28677 & ~n28852;
  assign n28854 = n28851 & ~n28853;
  assign n28855 = ~n28851 & n28853;
  assign n28856 = ~n28854 & ~n28855;
  assign n28857 = n6835 & n26043;
  assign n28858 = n7460 & n26284;
  assign n28859 = n6836 & n26540;
  assign n28860 = n7487 & n26532;
  assign n28861 = ~n28859 & ~n28860;
  assign n28862 = ~n28858 & n28861;
  assign n28863 = ~n28857 & n28862;
  assign n28864 = pi14  & n28863;
  assign n28865 = ~pi14  & ~n28863;
  assign n28866 = ~n28864 & ~n28865;
  assign n28867 = ~n28696 & n28707;
  assign n28868 = ~n28695 & ~n28867;
  assign n28869 = n28866 & n28868;
  assign n28870 = ~n28866 & ~n28868;
  assign n28871 = ~n28869 & ~n28870;
  assign n28872 = ~n28856 & n28871;
  assign n28873 = n28856 & ~n28871;
  assign n28874 = ~n28872 & ~n28873;
  assign n28875 = ~n28570 & ~n28710;
  assign n28876 = ~n28571 & ~n28875;
  assign n28877 = n28874 & n28876;
  assign n28878 = ~n28874 & ~n28876;
  assign n28879 = ~n28877 & ~n28878;
  assign n28880 = ~n28726 & n28879;
  assign n28881 = n28726 & ~n28879;
  assign n28882 = ~n28880 & ~n28881;
  assign n28883 = ~n28723 & ~n28882;
  assign n28884 = n28723 & n28882;
  assign po16  = ~n28883 & ~n28884;
  assign n28886 = ~n28877 & ~n28880;
  assign n28887 = ~n28866 & n28868;
  assign n28888 = ~n28873 & ~n28887;
  assign n28889 = n28838 & ~n28848;
  assign n28890 = ~n28855 & ~n28889;
  assign n28891 = ~n28830 & n28832;
  assign n28892 = ~n28837 & ~n28891;
  assign n28893 = n28802 & ~n28812;
  assign n28894 = ~n28819 & ~n28893;
  assign n28895 = ~n28736 & n28794;
  assign n28896 = ~n28801 & ~n28895;
  assign n28897 = n28773 & ~n28780;
  assign n28898 = ~n28786 & ~n28897;
  assign n28899 = ~n28769 & ~n28771;
  assign n28900 = n1656 & n2291;
  assign n28901 = n2814 & n28900;
  assign n28902 = n616 & n28901;
  assign n28903 = n13006 & n28902;
  assign n28904 = n2218 & n28903;
  assign n28905 = n13362 & n14621;
  assign n28906 = ~n578 & n28905;
  assign n28907 = n28904 & n28906;
  assign n28908 = n26865 & n28907;
  assign n28909 = n954 & n26389;
  assign n28910 = ~n638 & n28909;
  assign n28911 = ~n580 & n28910;
  assign n28912 = n1037 & n28911;
  assign n28913 = n28908 & n28912;
  assign n28914 = ~n28899 & n28913;
  assign n28915 = n28899 & ~n28913;
  assign n28916 = ~n28914 & ~n28915;
  assign n28917 = n3641 & n21204;
  assign n28918 = n3740 & n21201;
  assign n28919 = n556 & n22832;
  assign n28920 = n3961 & n21198;
  assign n28921 = ~n28919 & ~n28920;
  assign n28922 = ~n28918 & n28921;
  assign n28923 = ~n28917 & n28922;
  assign n28924 = n28916 & ~n28923;
  assign n28925 = ~n28916 & n28923;
  assign n28926 = ~n28924 & ~n28925;
  assign n28927 = n28898 & ~n28926;
  assign n28928 = ~n28898 & n28926;
  assign n28929 = ~n28927 & ~n28928;
  assign n28930 = n4006 & n21195;
  assign n28931 = n4133 & n21192;
  assign n28932 = n4002 & n23399;
  assign n28933 = n4555 & n21189;
  assign n28934 = ~n28932 & ~n28933;
  assign n28935 = ~n28931 & n28934;
  assign n28936 = ~n28930 & n28935;
  assign n28937 = pi29  & n28936;
  assign n28938 = ~pi29  & ~n28936;
  assign n28939 = ~n28937 & ~n28938;
  assign n28940 = n28929 & ~n28939;
  assign n28941 = ~n28929 & n28939;
  assign n28942 = ~n28940 & ~n28941;
  assign n28943 = n28746 & ~n28789;
  assign n28944 = ~n28790 & ~n28943;
  assign n28945 = n28942 & n28944;
  assign n28946 = ~n28942 & ~n28944;
  assign n28947 = ~n28945 & ~n28946;
  assign n28948 = n4601 & n21186;
  assign n28949 = n4783 & n21183;
  assign n28950 = n4602 & n23991;
  assign n28951 = n4801 & n21180;
  assign n28952 = ~n28950 & ~n28951;
  assign n28953 = ~n28949 & n28952;
  assign n28954 = ~n28948 & n28953;
  assign n28955 = pi26  & n28954;
  assign n28956 = ~pi26  & ~n28954;
  assign n28957 = ~n28955 & ~n28956;
  assign n28958 = n28947 & ~n28957;
  assign n28959 = ~n28947 & n28957;
  assign n28960 = ~n28958 & ~n28959;
  assign n28961 = n28896 & ~n28960;
  assign n28962 = ~n28896 & n28960;
  assign n28963 = ~n28961 & ~n28962;
  assign n28964 = n5238 & n21076;
  assign n28965 = n71 & n21176;
  assign n28966 = n5239 & ~n21470;
  assign n28967 = n5326 & n21464;
  assign n28968 = ~n28966 & ~n28967;
  assign n28969 = ~n28965 & n28968;
  assign n28970 = ~n28964 & n28969;
  assign n28971 = pi23  & n28970;
  assign n28972 = ~pi23  & ~n28970;
  assign n28973 = ~n28971 & ~n28972;
  assign n28974 = n28963 & ~n28973;
  assign n28975 = ~n28963 & n28973;
  assign n28976 = ~n28974 & ~n28975;
  assign n28977 = n28894 & ~n28976;
  assign n28978 = ~n28894 & n28976;
  assign n28979 = ~n28977 & ~n28978;
  assign n28980 = n5435 & n24607;
  assign n28981 = n6055 & n24676;
  assign n28982 = n5429 & ~n24754;
  assign n28983 = n6071 & n24748;
  assign n28984 = ~n28982 & ~n28983;
  assign n28985 = ~n28981 & n28984;
  assign n28986 = ~n28980 & n28985;
  assign n28987 = pi20  & n28986;
  assign n28988 = ~pi20  & ~n28986;
  assign n28989 = ~n28987 & ~n28988;
  assign n28990 = n28979 & ~n28989;
  assign n28991 = ~n28979 & n28989;
  assign n28992 = ~n28990 & ~n28991;
  assign n28993 = n28892 & n28992;
  assign n28994 = ~n28892 & ~n28992;
  assign n28995 = ~n28993 & ~n28994;
  assign n28996 = n6184 & n25521;
  assign n28997 = n6527 & n25785;
  assign n28998 = n6185 & n26049;
  assign n28999 = n6543 & n26043;
  assign n29000 = ~n28998 & ~n28999;
  assign n29001 = ~n28997 & n29000;
  assign n29002 = ~n28996 & n29001;
  assign n29003 = pi17  & n29002;
  assign n29004 = ~pi17  & ~n29002;
  assign n29005 = ~n29003 & ~n29004;
  assign n29006 = ~n28995 & ~n29005;
  assign n29007 = n28995 & n29005;
  assign n29008 = ~n29006 & ~n29007;
  assign n29009 = n28890 & ~n29008;
  assign n29010 = ~n28890 & n29008;
  assign n29011 = ~n29009 & ~n29010;
  assign n29012 = n6835 & n26284;
  assign n29013 = n7460 & n26532;
  assign n29014 = n6836 & ~n26770;
  assign n29015 = n7487 & n26764;
  assign n29016 = ~n29014 & ~n29015;
  assign n29017 = ~n29013 & n29016;
  assign n29018 = ~n29012 & n29017;
  assign n29019 = pi14  & n29018;
  assign n29020 = ~pi14  & ~n29018;
  assign n29021 = ~n29019 & ~n29020;
  assign n29022 = n29011 & ~n29021;
  assign n29023 = ~n29011 & n29021;
  assign n29024 = ~n29022 & ~n29023;
  assign n29025 = ~n28888 & n29024;
  assign n29026 = n28888 & ~n29024;
  assign n29027 = ~n29025 & ~n29026;
  assign n29028 = n28886 & ~n29027;
  assign n29029 = ~n28886 & n29027;
  assign n29030 = ~n29028 & ~n29029;
  assign n29031 = n28884 & n29030;
  assign n29032 = ~n28884 & ~n29030;
  assign po17  = ~n29031 & ~n29032;
  assign n29034 = ~n28892 & n28992;
  assign n29035 = ~n29006 & ~n29034;
  assign n29036 = n6836 & n26987;
  assign n29037 = n6835 & n26532;
  assign n29038 = ~n14792 & n26764;
  assign n29039 = ~n29037 & ~n29038;
  assign n29040 = ~n29036 & n29039;
  assign n29041 = pi14  & n29040;
  assign n29042 = ~pi14  & ~n29040;
  assign n29043 = ~n29041 & ~n29042;
  assign n29044 = ~n29035 & ~n29043;
  assign n29045 = n29035 & n29043;
  assign n29046 = ~n29044 & ~n29045;
  assign n29047 = n1605 & n2896;
  assign n29048 = n4422 & n29047;
  assign n29049 = n3919 & n29048;
  assign n29050 = ~n595 & n29049;
  assign n29051 = ~n423 & n29050;
  assign n29052 = n963 & n5849;
  assign n29053 = ~n307 & n29052;
  assign n29054 = ~n245 & n29053;
  assign n29055 = n29051 & n29054;
  assign n29056 = n3183 & n3702;
  assign n29057 = ~n206 & n29056;
  assign n29058 = ~n580 & n29057;
  assign n29059 = n300 & n3849;
  assign n29060 = ~n243 & n29059;
  assign n29061 = ~n361 & n29060;
  assign n29062 = n29058 & n29061;
  assign n29063 = n29055 & n29062;
  assign n29064 = ~n28913 & n29063;
  assign n29065 = n28913 & ~n29063;
  assign n29066 = ~n29064 & ~n29065;
  assign n29067 = n3641 & n21201;
  assign n29068 = n3740 & n21198;
  assign n29069 = n556 & n21482;
  assign n29070 = n3961 & n21195;
  assign n29071 = ~n29069 & ~n29070;
  assign n29072 = ~n29068 & n29071;
  assign n29073 = ~n29067 & n29072;
  assign n29074 = ~n29066 & n29073;
  assign n29075 = n29066 & ~n29073;
  assign n29076 = ~n29074 & ~n29075;
  assign n29077 = ~n28914 & n28923;
  assign n29078 = ~n28915 & ~n29077;
  assign n29079 = ~n29076 & ~n29078;
  assign n29080 = n29076 & n29078;
  assign n29081 = ~n29079 & ~n29080;
  assign n29082 = ~n28928 & ~n28940;
  assign n29083 = ~n29081 & n29082;
  assign n29084 = n29081 & ~n29082;
  assign n29085 = ~n29083 & ~n29084;
  assign n29086 = n4006 & n21192;
  assign n29087 = n4133 & n21189;
  assign n29088 = n4002 & n23384;
  assign n29089 = n4555 & n21186;
  assign n29090 = ~n29088 & ~n29089;
  assign n29091 = ~n29087 & n29090;
  assign n29092 = ~n29086 & n29091;
  assign n29093 = pi29  & n29092;
  assign n29094 = ~pi29  & ~n29092;
  assign n29095 = ~n29093 & ~n29094;
  assign n29096 = n29085 & n29095;
  assign n29097 = ~n29085 & ~n29095;
  assign n29098 = ~n29096 & ~n29097;
  assign n29099 = n4601 & n21183;
  assign n29100 = n4783 & n21180;
  assign n29101 = n4602 & n24030;
  assign n29102 = n4801 & n21076;
  assign n29103 = ~n29101 & ~n29102;
  assign n29104 = ~n29100 & n29103;
  assign n29105 = ~n29099 & n29104;
  assign n29106 = pi26  & n29105;
  assign n29107 = ~pi26  & ~n29105;
  assign n29108 = ~n29106 & ~n29107;
  assign n29109 = ~n29098 & ~n29108;
  assign n29110 = n29098 & n29108;
  assign n29111 = ~n29109 & ~n29110;
  assign n29112 = ~n28945 & n28957;
  assign n29113 = ~n28946 & ~n29112;
  assign n29114 = ~n29111 & ~n29113;
  assign n29115 = n29111 & n29113;
  assign n29116 = ~n29114 & ~n29115;
  assign n29117 = n5238 & n21176;
  assign n29118 = n71 & n21464;
  assign n29119 = n5239 & n24782;
  assign n29120 = n5326 & n24607;
  assign n29121 = ~n29119 & ~n29120;
  assign n29122 = ~n29118 & n29121;
  assign n29123 = ~n29117 & n29122;
  assign n29124 = pi23  & n29123;
  assign n29125 = ~pi23  & ~n29123;
  assign n29126 = ~n29124 & ~n29125;
  assign n29127 = n29116 & ~n29126;
  assign n29128 = ~n29116 & n29126;
  assign n29129 = ~n29127 & ~n29128;
  assign n29130 = ~n28962 & n28973;
  assign n29131 = ~n28961 & ~n29130;
  assign n29132 = ~n29129 & ~n29131;
  assign n29133 = n29129 & n29131;
  assign n29134 = ~n29132 & ~n29133;
  assign n29135 = n5435 & n24676;
  assign n29136 = n6055 & n24748;
  assign n29137 = n5429 & ~n25529;
  assign n29138 = n6071 & n25521;
  assign n29139 = ~n29137 & ~n29138;
  assign n29140 = ~n29136 & n29139;
  assign n29141 = ~n29135 & n29140;
  assign n29142 = pi20  & n29141;
  assign n29143 = ~pi20  & ~n29141;
  assign n29144 = ~n29142 & ~n29143;
  assign n29145 = n29134 & ~n29144;
  assign n29146 = ~n29134 & n29144;
  assign n29147 = ~n29145 & ~n29146;
  assign n29148 = ~n28978 & n28989;
  assign n29149 = ~n28977 & ~n29148;
  assign n29150 = ~n29147 & ~n29149;
  assign n29151 = n29147 & n29149;
  assign n29152 = ~n29150 & ~n29151;
  assign n29153 = n6184 & n25785;
  assign n29154 = n6527 & n26043;
  assign n29155 = n6185 & ~n26290;
  assign n29156 = n6543 & n26284;
  assign n29157 = ~n29155 & ~n29156;
  assign n29158 = ~n29154 & n29157;
  assign n29159 = ~n29153 & n29158;
  assign n29160 = pi17  & n29159;
  assign n29161 = ~pi17  & ~n29159;
  assign n29162 = ~n29160 & ~n29161;
  assign n29163 = n29152 & ~n29162;
  assign n29164 = ~n29152 & n29162;
  assign n29165 = ~n29163 & ~n29164;
  assign n29166 = n29046 & n29165;
  assign n29167 = ~n29046 & ~n29165;
  assign n29168 = ~n29166 & ~n29167;
  assign n29169 = ~n29010 & n29021;
  assign n29170 = ~n29009 & ~n29169;
  assign n29171 = ~n29168 & ~n29170;
  assign n29172 = n29168 & n29170;
  assign n29173 = ~n29171 & ~n29172;
  assign n29174 = ~n29025 & ~n29029;
  assign n29175 = ~n29173 & n29174;
  assign n29176 = n29173 & ~n29174;
  assign n29177 = ~n29175 & ~n29176;
  assign n29178 = n29031 & n29177;
  assign n29179 = ~n29031 & ~n29177;
  assign po18  = ~n29178 & ~n29179;
  assign n29181 = ~n29172 & ~n29176;
  assign n29182 = ~n29080 & ~n29084;
  assign n29183 = n4006 & n21189;
  assign n29184 = n4133 & n21186;
  assign n29185 = n4002 & n23369;
  assign n29186 = n4555 & n21183;
  assign n29187 = ~n29185 & ~n29186;
  assign n29188 = ~n29184 & n29187;
  assign n29189 = ~n29183 & n29188;
  assign n29190 = pi29  & n29189;
  assign n29191 = ~pi29  & ~n29189;
  assign n29192 = ~n29190 & ~n29191;
  assign n29193 = ~n13151 & n26764;
  assign n29194 = pi14  & ~n29193;
  assign n29195 = ~pi14  & n29193;
  assign n29196 = ~n29194 & ~n29195;
  assign n29197 = n2642 & n13809;
  assign n29198 = n1283 & n29197;
  assign n29199 = n3230 & n4350;
  assign n29200 = n2104 & n29199;
  assign n29201 = ~n527 & n29200;
  assign n29202 = n29198 & n29201;
  assign n29203 = n1888 & n7296;
  assign n29204 = ~n206 & n29203;
  assign n29205 = n1924 & n13567;
  assign n29206 = ~n229 & n29205;
  assign n29207 = n29204 & n29206;
  assign n29208 = n29202 & n29207;
  assign n29209 = n28913 & n29208;
  assign n29210 = ~n28913 & ~n29208;
  assign n29211 = ~n29209 & ~n29210;
  assign n29212 = n29196 & n29211;
  assign n29213 = ~n29196 & ~n29211;
  assign n29214 = ~n29212 & ~n29213;
  assign n29215 = ~n29065 & n29073;
  assign n29216 = ~n29064 & ~n29215;
  assign n29217 = n29214 & n29216;
  assign n29218 = ~n29214 & ~n29216;
  assign n29219 = ~n29217 & ~n29218;
  assign n29220 = n3641 & n21198;
  assign n29221 = n3740 & n21195;
  assign n29222 = n556 & n23211;
  assign n29223 = n3961 & n21192;
  assign n29224 = ~n29222 & ~n29223;
  assign n29225 = ~n29221 & n29224;
  assign n29226 = ~n29220 & n29225;
  assign n29227 = n29219 & ~n29226;
  assign n29228 = ~n29219 & n29226;
  assign n29229 = ~n29227 & ~n29228;
  assign n29230 = ~n29192 & n29229;
  assign n29231 = n29192 & ~n29229;
  assign n29232 = ~n29230 & ~n29231;
  assign n29233 = n29182 & ~n29232;
  assign n29234 = ~n29182 & n29232;
  assign n29235 = ~n29233 & ~n29234;
  assign n29236 = n4601 & n21180;
  assign n29237 = n4783 & n21076;
  assign n29238 = n4602 & n24012;
  assign n29239 = n4801 & n21176;
  assign n29240 = ~n29238 & ~n29239;
  assign n29241 = ~n29237 & n29240;
  assign n29242 = ~n29236 & n29241;
  assign n29243 = pi26  & n29242;
  assign n29244 = ~pi26  & ~n29242;
  assign n29245 = ~n29243 & ~n29244;
  assign n29246 = n29235 & n29245;
  assign n29247 = ~n29235 & ~n29245;
  assign n29248 = ~n29246 & ~n29247;
  assign n29249 = n29085 & ~n29095;
  assign n29250 = ~n29109 & ~n29249;
  assign n29251 = n29248 & n29250;
  assign n29252 = ~n29248 & ~n29250;
  assign n29253 = ~n29251 & ~n29252;
  assign n29254 = n5238 & n21464;
  assign n29255 = n71 & n24607;
  assign n29256 = n5239 & n24770;
  assign n29257 = n5326 & n24676;
  assign n29258 = ~n29256 & ~n29257;
  assign n29259 = ~n29255 & n29258;
  assign n29260 = ~n29254 & n29259;
  assign n29261 = pi23  & n29260;
  assign n29262 = ~pi23  & ~n29260;
  assign n29263 = ~n29261 & ~n29262;
  assign n29264 = ~n29115 & n29126;
  assign n29265 = ~n29114 & ~n29264;
  assign n29266 = n29263 & n29265;
  assign n29267 = ~n29263 & ~n29265;
  assign n29268 = ~n29266 & ~n29267;
  assign n29269 = ~n29253 & n29268;
  assign n29270 = n29253 & ~n29268;
  assign n29271 = ~n29269 & ~n29270;
  assign n29272 = n5435 & n24748;
  assign n29273 = n6055 & n25521;
  assign n29274 = n5429 & n25793;
  assign n29275 = n6071 & n25785;
  assign n29276 = ~n29274 & ~n29275;
  assign n29277 = ~n29273 & n29276;
  assign n29278 = ~n29272 & n29277;
  assign n29279 = pi20  & n29278;
  assign n29280 = ~pi20  & ~n29278;
  assign n29281 = ~n29279 & ~n29280;
  assign n29282 = n29271 & n29281;
  assign n29283 = ~n29271 & ~n29281;
  assign n29284 = ~n29282 & ~n29283;
  assign n29285 = ~n29133 & n29144;
  assign n29286 = ~n29132 & ~n29285;
  assign n29287 = n29284 & ~n29286;
  assign n29288 = ~n29284 & n29286;
  assign n29289 = ~n29287 & ~n29288;
  assign n29290 = n6184 & n26043;
  assign n29291 = n6527 & n26284;
  assign n29292 = n6185 & n26540;
  assign n29293 = n6543 & n26532;
  assign n29294 = ~n29292 & ~n29293;
  assign n29295 = ~n29291 & n29294;
  assign n29296 = ~n29290 & n29295;
  assign n29297 = pi17  & n29296;
  assign n29298 = ~pi17  & ~n29296;
  assign n29299 = ~n29297 & ~n29298;
  assign n29300 = ~n29151 & n29162;
  assign n29301 = ~n29150 & ~n29300;
  assign n29302 = n29299 & n29301;
  assign n29303 = ~n29299 & ~n29301;
  assign n29304 = ~n29302 & ~n29303;
  assign n29305 = ~n29289 & n29304;
  assign n29306 = n29289 & ~n29304;
  assign n29307 = ~n29305 & ~n29306;
  assign n29308 = ~n29044 & ~n29165;
  assign n29309 = ~n29045 & ~n29308;
  assign n29310 = n29307 & n29309;
  assign n29311 = ~n29307 & ~n29309;
  assign n29312 = ~n29310 & ~n29311;
  assign n29313 = ~n29181 & n29312;
  assign n29314 = n29181 & ~n29312;
  assign n29315 = ~n29313 & ~n29314;
  assign n29316 = ~n29178 & ~n29315;
  assign n29317 = n29178 & n29315;
  assign po19  = ~n29316 & ~n29317;
  assign n29319 = ~n29310 & ~n29313;
  assign n29320 = ~n29299 & n29301;
  assign n29321 = ~n29306 & ~n29320;
  assign n29322 = n29271 & ~n29281;
  assign n29323 = ~n29288 & ~n29322;
  assign n29324 = ~n29263 & n29265;
  assign n29325 = ~n29270 & ~n29324;
  assign n29326 = n29235 & ~n29245;
  assign n29327 = ~n29252 & ~n29326;
  assign n29328 = ~n29230 & ~n29234;
  assign n29329 = ~n29210 & ~n29212;
  assign n29330 = ~n468 & n2566;
  assign n29331 = n969 & n2260;
  assign n29332 = n515 & n29331;
  assign n29333 = n930 & n13851;
  assign n29334 = n997 & n29333;
  assign n29335 = n2021 & n29334;
  assign n29336 = n386 & n29335;
  assign n29337 = n29332 & n29336;
  assign n29338 = n5695 & n29337;
  assign n29339 = ~n238 & n29338;
  assign n29340 = n1813 & n6398;
  assign n29341 = n3495 & n29340;
  assign n29342 = ~n689 & n29341;
  assign n29343 = n29339 & n29342;
  assign n29344 = ~n332 & n29343;
  assign n29345 = n29330 & n29344;
  assign n29346 = ~n29329 & n29345;
  assign n29347 = n29329 & ~n29345;
  assign n29348 = ~n29346 & ~n29347;
  assign n29349 = n3641 & n21195;
  assign n29350 = n3740 & n21192;
  assign n29351 = n556 & n23399;
  assign n29352 = n3961 & n21189;
  assign n29353 = ~n29351 & ~n29352;
  assign n29354 = ~n29350 & n29353;
  assign n29355 = ~n29349 & n29354;
  assign n29356 = n29348 & ~n29355;
  assign n29357 = ~n29348 & n29355;
  assign n29358 = ~n29356 & ~n29357;
  assign n29359 = ~n29217 & n29226;
  assign n29360 = ~n29218 & ~n29359;
  assign n29361 = ~n29358 & ~n29360;
  assign n29362 = n29358 & n29360;
  assign n29363 = ~n29361 & ~n29362;
  assign n29364 = n4006 & n21186;
  assign n29365 = n4133 & n21183;
  assign n29366 = n4002 & n23991;
  assign n29367 = n4555 & n21180;
  assign n29368 = ~n29366 & ~n29367;
  assign n29369 = ~n29365 & n29368;
  assign n29370 = ~n29364 & n29369;
  assign n29371 = pi29  & n29370;
  assign n29372 = ~pi29  & ~n29370;
  assign n29373 = ~n29371 & ~n29372;
  assign n29374 = n29363 & ~n29373;
  assign n29375 = ~n29363 & n29373;
  assign n29376 = ~n29374 & ~n29375;
  assign n29377 = ~n29328 & n29376;
  assign n29378 = n29328 & ~n29376;
  assign n29379 = ~n29377 & ~n29378;
  assign n29380 = n4601 & n21076;
  assign n29381 = n4783 & n21176;
  assign n29382 = n4602 & ~n21470;
  assign n29383 = n4801 & n21464;
  assign n29384 = ~n29382 & ~n29383;
  assign n29385 = ~n29381 & n29384;
  assign n29386 = ~n29380 & n29385;
  assign n29387 = pi26  & n29386;
  assign n29388 = ~pi26  & ~n29386;
  assign n29389 = ~n29387 & ~n29388;
  assign n29390 = n29379 & ~n29389;
  assign n29391 = ~n29379 & n29389;
  assign n29392 = ~n29390 & ~n29391;
  assign n29393 = n29327 & ~n29392;
  assign n29394 = ~n29327 & n29392;
  assign n29395 = ~n29393 & ~n29394;
  assign n29396 = n5238 & n24607;
  assign n29397 = n71 & n24676;
  assign n29398 = n5239 & ~n24754;
  assign n29399 = n5326 & n24748;
  assign n29400 = ~n29398 & ~n29399;
  assign n29401 = ~n29397 & n29400;
  assign n29402 = ~n29396 & n29401;
  assign n29403 = pi23  & n29402;
  assign n29404 = ~pi23  & ~n29402;
  assign n29405 = ~n29403 & ~n29404;
  assign n29406 = n29395 & ~n29405;
  assign n29407 = ~n29395 & n29405;
  assign n29408 = ~n29406 & ~n29407;
  assign n29409 = n29325 & n29408;
  assign n29410 = ~n29325 & ~n29408;
  assign n29411 = ~n29409 & ~n29410;
  assign n29412 = n5435 & n25521;
  assign n29413 = n6055 & n25785;
  assign n29414 = n5429 & n26049;
  assign n29415 = n6071 & n26043;
  assign n29416 = ~n29414 & ~n29415;
  assign n29417 = ~n29413 & n29416;
  assign n29418 = ~n29412 & n29417;
  assign n29419 = pi20  & n29418;
  assign n29420 = ~pi20  & ~n29418;
  assign n29421 = ~n29419 & ~n29420;
  assign n29422 = ~n29411 & ~n29421;
  assign n29423 = n29411 & n29421;
  assign n29424 = ~n29422 & ~n29423;
  assign n29425 = n29323 & ~n29424;
  assign n29426 = ~n29323 & n29424;
  assign n29427 = ~n29425 & ~n29426;
  assign n29428 = n6184 & n26284;
  assign n29429 = n6527 & n26532;
  assign n29430 = n6185 & ~n26770;
  assign n29431 = n6543 & n26764;
  assign n29432 = ~n29430 & ~n29431;
  assign n29433 = ~n29429 & n29432;
  assign n29434 = ~n29428 & n29433;
  assign n29435 = pi17  & n29434;
  assign n29436 = ~pi17  & ~n29434;
  assign n29437 = ~n29435 & ~n29436;
  assign n29438 = n29427 & ~n29437;
  assign n29439 = ~n29427 & n29437;
  assign n29440 = ~n29438 & ~n29439;
  assign n29441 = ~n29321 & n29440;
  assign n29442 = n29321 & ~n29440;
  assign n29443 = ~n29441 & ~n29442;
  assign n29444 = n29319 & ~n29443;
  assign n29445 = ~n29319 & n29443;
  assign n29446 = ~n29444 & ~n29445;
  assign n29447 = n29317 & n29446;
  assign n29448 = ~n29317 & ~n29446;
  assign po20  = ~n29447 & ~n29448;
  assign n29450 = ~n29325 & n29408;
  assign n29451 = ~n29422 & ~n29450;
  assign n29452 = n6185 & n26987;
  assign n29453 = n6184 & n26532;
  assign n29454 = ~n14132 & n26764;
  assign n29455 = ~n29453 & ~n29454;
  assign n29456 = ~n29452 & n29455;
  assign n29457 = pi17  & n29456;
  assign n29458 = ~pi17  & ~n29456;
  assign n29459 = ~n29457 & ~n29458;
  assign n29460 = ~n29451 & ~n29459;
  assign n29461 = n29451 & n29459;
  assign n29462 = ~n29460 & ~n29461;
  assign n29463 = ~n29362 & ~n29374;
  assign n29464 = n4006 & n21183;
  assign n29465 = n4133 & n21180;
  assign n29466 = n4002 & n24030;
  assign n29467 = n4555 & n21076;
  assign n29468 = ~n29466 & ~n29467;
  assign n29469 = ~n29465 & n29468;
  assign n29470 = ~n29464 & n29469;
  assign n29471 = pi29  & n29470;
  assign n29472 = ~pi29  & ~n29470;
  assign n29473 = ~n29471 & ~n29472;
  assign n29474 = n841 & n5878;
  assign n29475 = ~n631 & n29474;
  assign n29476 = n1998 & n3916;
  assign n29477 = n1517 & n29476;
  assign n29478 = n29475 & n29477;
  assign n29479 = ~n81 & n2070;
  assign n29480 = ~n678 & n29479;
  assign n29481 = n3220 & n29480;
  assign n29482 = n2218 & n29481;
  assign n29483 = ~n462 & n29482;
  assign n29484 = n1389 & n2760;
  assign n29485 = n1238 & n29484;
  assign n29486 = n107 & n29485;
  assign n29487 = ~n429 & n29486;
  assign n29488 = ~n183 & n29487;
  assign n29489 = n29483 & n29488;
  assign n29490 = n29478 & n29489;
  assign n29491 = n29345 & ~n29490;
  assign n29492 = ~n29345 & n29490;
  assign n29493 = ~n29491 & ~n29492;
  assign n29494 = ~n29346 & n29355;
  assign n29495 = ~n29347 & ~n29494;
  assign n29496 = n29493 & ~n29495;
  assign n29497 = ~n29493 & n29495;
  assign n29498 = ~n29496 & ~n29497;
  assign n29499 = n3641 & n21192;
  assign n29500 = n3740 & n21189;
  assign n29501 = n556 & n23384;
  assign n29502 = n3961 & n21186;
  assign n29503 = ~n29501 & ~n29502;
  assign n29504 = ~n29500 & n29503;
  assign n29505 = ~n29499 & n29504;
  assign n29506 = ~n29498 & ~n29505;
  assign n29507 = n29498 & n29505;
  assign n29508 = ~n29506 & ~n29507;
  assign n29509 = ~n29473 & n29508;
  assign n29510 = n29473 & ~n29508;
  assign n29511 = ~n29509 & ~n29510;
  assign n29512 = ~n29463 & n29511;
  assign n29513 = n29463 & ~n29511;
  assign n29514 = ~n29512 & ~n29513;
  assign n29515 = n4601 & n21176;
  assign n29516 = n4783 & n21464;
  assign n29517 = n4602 & n24782;
  assign n29518 = n4801 & n24607;
  assign n29519 = ~n29517 & ~n29518;
  assign n29520 = ~n29516 & n29519;
  assign n29521 = ~n29515 & n29520;
  assign n29522 = pi26  & n29521;
  assign n29523 = ~pi26  & ~n29521;
  assign n29524 = ~n29522 & ~n29523;
  assign n29525 = n29514 & ~n29524;
  assign n29526 = ~n29514 & n29524;
  assign n29527 = ~n29525 & ~n29526;
  assign n29528 = ~n29377 & n29389;
  assign n29529 = ~n29378 & ~n29528;
  assign n29530 = ~n29527 & ~n29529;
  assign n29531 = n29527 & n29529;
  assign n29532 = ~n29530 & ~n29531;
  assign n29533 = n5238 & n24676;
  assign n29534 = n71 & n24748;
  assign n29535 = n5239 & ~n25529;
  assign n29536 = n5326 & n25521;
  assign n29537 = ~n29535 & ~n29536;
  assign n29538 = ~n29534 & n29537;
  assign n29539 = ~n29533 & n29538;
  assign n29540 = pi23  & n29539;
  assign n29541 = ~pi23  & ~n29539;
  assign n29542 = ~n29540 & ~n29541;
  assign n29543 = n29532 & ~n29542;
  assign n29544 = ~n29532 & n29542;
  assign n29545 = ~n29543 & ~n29544;
  assign n29546 = ~n29394 & n29405;
  assign n29547 = ~n29393 & ~n29546;
  assign n29548 = ~n29545 & ~n29547;
  assign n29549 = n29545 & n29547;
  assign n29550 = ~n29548 & ~n29549;
  assign n29551 = n5435 & n25785;
  assign n29552 = n6055 & n26043;
  assign n29553 = n5429 & ~n26290;
  assign n29554 = n6071 & n26284;
  assign n29555 = ~n29553 & ~n29554;
  assign n29556 = ~n29552 & n29555;
  assign n29557 = ~n29551 & n29556;
  assign n29558 = pi20  & n29557;
  assign n29559 = ~pi20  & ~n29557;
  assign n29560 = ~n29558 & ~n29559;
  assign n29561 = n29550 & ~n29560;
  assign n29562 = ~n29550 & n29560;
  assign n29563 = ~n29561 & ~n29562;
  assign n29564 = n29462 & n29563;
  assign n29565 = ~n29462 & ~n29563;
  assign n29566 = ~n29564 & ~n29565;
  assign n29567 = ~n29426 & n29437;
  assign n29568 = ~n29425 & ~n29567;
  assign n29569 = ~n29566 & ~n29568;
  assign n29570 = n29566 & n29568;
  assign n29571 = ~n29569 & ~n29570;
  assign n29572 = ~n29441 & ~n29445;
  assign n29573 = ~n29571 & n29572;
  assign n29574 = n29571 & ~n29572;
  assign n29575 = ~n29573 & ~n29574;
  assign n29576 = n29447 & n29575;
  assign n29577 = ~n29447 & ~n29575;
  assign po21  = ~n29576 & ~n29577;
  assign n29579 = ~n29570 & ~n29574;
  assign n29580 = n5238 & n24748;
  assign n29581 = n71 & n25521;
  assign n29582 = n5239 & n25793;
  assign n29583 = n5326 & n25785;
  assign n29584 = ~n29582 & ~n29583;
  assign n29585 = ~n29581 & n29584;
  assign n29586 = ~n29580 & n29585;
  assign n29587 = pi23  & n29586;
  assign n29588 = ~pi23  & ~n29586;
  assign n29589 = ~n29587 & ~n29588;
  assign n29590 = n4601 & n21464;
  assign n29591 = n4783 & n24607;
  assign n29592 = n4602 & n24770;
  assign n29593 = n4801 & n24676;
  assign n29594 = ~n29592 & ~n29593;
  assign n29595 = ~n29591 & n29594;
  assign n29596 = ~n29590 & n29595;
  assign n29597 = pi26  & n29596;
  assign n29598 = ~pi26  & ~n29596;
  assign n29599 = ~n29597 & ~n29598;
  assign n29600 = ~n29512 & n29524;
  assign n29601 = ~n29513 & ~n29600;
  assign n29602 = n29599 & n29601;
  assign n29603 = ~n29599 & ~n29601;
  assign n29604 = ~n29602 & ~n29603;
  assign n29605 = n4006 & n21180;
  assign n29606 = n4133 & n21076;
  assign n29607 = n4002 & n24012;
  assign n29608 = n4555 & n21176;
  assign n29609 = ~n29607 & ~n29608;
  assign n29610 = ~n29606 & n29609;
  assign n29611 = ~n29605 & n29610;
  assign n29612 = pi29  & n29611;
  assign n29613 = ~pi29  & ~n29611;
  assign n29614 = ~n29612 & ~n29613;
  assign n29615 = ~n29506 & ~n29509;
  assign n29616 = ~n12977 & n26764;
  assign n29617 = pi17  & ~n29616;
  assign n29618 = ~pi17  & n29616;
  assign n29619 = ~n29617 & ~n29618;
  assign n29620 = n1945 & n3473;
  assign n29621 = ~n275 & n29620;
  assign n29622 = n1748 & n23262;
  assign n29623 = n1395 & n29622;
  assign n29624 = ~n401 & n29623;
  assign n29625 = n29621 & n29624;
  assign n29626 = n1503 & n12889;
  assign n29627 = ~n183 & n29626;
  assign n29628 = n4698 & n5511;
  assign n29629 = ~n583 & n29628;
  assign n29630 = ~n85 & n29629;
  assign n29631 = n29627 & n29630;
  assign n29632 = n29625 & n29631;
  assign n29633 = n29490 & n29632;
  assign n29634 = ~n29490 & ~n29632;
  assign n29635 = ~n29633 & ~n29634;
  assign n29636 = n29619 & n29635;
  assign n29637 = ~n29619 & ~n29635;
  assign n29638 = ~n29636 & ~n29637;
  assign n29639 = n3641 & n21189;
  assign n29640 = n3740 & n21186;
  assign n29641 = n556 & n23369;
  assign n29642 = n3961 & n21183;
  assign n29643 = ~n29641 & ~n29642;
  assign n29644 = ~n29640 & n29643;
  assign n29645 = ~n29639 & n29644;
  assign n29646 = n29638 & n29645;
  assign n29647 = ~n29638 & ~n29645;
  assign n29648 = ~n29646 & ~n29647;
  assign n29649 = ~n29492 & ~n29495;
  assign n29650 = ~n29491 & ~n29649;
  assign n29651 = ~n29648 & n29650;
  assign n29652 = n29648 & ~n29650;
  assign n29653 = ~n29651 & ~n29652;
  assign n29654 = ~n29615 & n29653;
  assign n29655 = n29615 & ~n29653;
  assign n29656 = ~n29654 & ~n29655;
  assign n29657 = n29614 & ~n29656;
  assign n29658 = ~n29614 & n29656;
  assign n29659 = ~n29657 & ~n29658;
  assign n29660 = ~n29604 & n29659;
  assign n29661 = n29604 & ~n29659;
  assign n29662 = ~n29660 & ~n29661;
  assign n29663 = ~n29589 & n29662;
  assign n29664 = n29589 & ~n29662;
  assign n29665 = ~n29663 & ~n29664;
  assign n29666 = ~n29531 & n29542;
  assign n29667 = ~n29530 & ~n29666;
  assign n29668 = ~n29665 & ~n29667;
  assign n29669 = n29665 & n29667;
  assign n29670 = ~n29668 & ~n29669;
  assign n29671 = n5435 & n26043;
  assign n29672 = n6055 & n26284;
  assign n29673 = n5429 & n26540;
  assign n29674 = n6071 & n26532;
  assign n29675 = ~n29673 & ~n29674;
  assign n29676 = ~n29672 & n29675;
  assign n29677 = ~n29671 & n29676;
  assign n29678 = pi20  & n29677;
  assign n29679 = ~pi20  & ~n29677;
  assign n29680 = ~n29678 & ~n29679;
  assign n29681 = ~n29549 & n29560;
  assign n29682 = ~n29548 & ~n29681;
  assign n29683 = n29680 & n29682;
  assign n29684 = ~n29680 & ~n29682;
  assign n29685 = ~n29683 & ~n29684;
  assign n29686 = ~n29670 & n29685;
  assign n29687 = n29670 & ~n29685;
  assign n29688 = ~n29686 & ~n29687;
  assign n29689 = ~n29460 & ~n29563;
  assign n29690 = ~n29461 & ~n29689;
  assign n29691 = n29688 & n29690;
  assign n29692 = ~n29688 & ~n29690;
  assign n29693 = ~n29691 & ~n29692;
  assign n29694 = ~n29579 & n29693;
  assign n29695 = n29579 & ~n29693;
  assign n29696 = ~n29694 & ~n29695;
  assign n29697 = ~n29576 & ~n29696;
  assign n29698 = n29576 & n29696;
  assign po22  = ~n29697 & ~n29698;
  assign n29700 = ~n29680 & n29682;
  assign n29701 = ~n29687 & ~n29700;
  assign n29702 = ~n29663 & ~n29669;
  assign n29703 = n5238 & n25521;
  assign n29704 = n71 & n25785;
  assign n29705 = n5239 & n26049;
  assign n29706 = n5326 & n26043;
  assign n29707 = ~n29705 & ~n29706;
  assign n29708 = ~n29704 & n29707;
  assign n29709 = ~n29703 & n29708;
  assign n29710 = pi23  & n29709;
  assign n29711 = ~pi23  & ~n29709;
  assign n29712 = ~n29710 & ~n29711;
  assign n29713 = ~n29599 & n29601;
  assign n29714 = ~n29660 & ~n29713;
  assign n29715 = n29638 & ~n29645;
  assign n29716 = ~n29651 & ~n29715;
  assign n29717 = ~n29634 & ~n29636;
  assign n29718 = n1207 & n3236;
  assign n29719 = n1132 & n29718;
  assign n29720 = ~n690 & n29719;
  assign n29721 = n3341 & n7060;
  assign n29722 = n1516 & n29721;
  assign n29723 = ~n305 & n29722;
  assign n29724 = ~n193 & n29723;
  assign n29725 = n29720 & n29724;
  assign n29726 = n4888 & n12586;
  assign n29727 = ~n203 & n29726;
  assign n29728 = n1588 & n28043;
  assign n29729 = ~n601 & n29728;
  assign n29730 = ~n259 & n29729;
  assign n29731 = n29727 & n29730;
  assign n29732 = n29725 & n29731;
  assign n29733 = ~n29717 & n29732;
  assign n29734 = n29717 & ~n29732;
  assign n29735 = ~n29733 & ~n29734;
  assign n29736 = n3641 & n21186;
  assign n29737 = n3740 & n21183;
  assign n29738 = n556 & n23991;
  assign n29739 = n3961 & n21180;
  assign n29740 = ~n29738 & ~n29739;
  assign n29741 = ~n29737 & n29740;
  assign n29742 = ~n29736 & n29741;
  assign n29743 = n29735 & ~n29742;
  assign n29744 = ~n29735 & n29742;
  assign n29745 = ~n29743 & ~n29744;
  assign n29746 = n29716 & ~n29745;
  assign n29747 = ~n29716 & n29745;
  assign n29748 = ~n29746 & ~n29747;
  assign n29749 = n4006 & n21076;
  assign n29750 = n4133 & n21176;
  assign n29751 = n4002 & ~n21470;
  assign n29752 = n4555 & n21464;
  assign n29753 = ~n29751 & ~n29752;
  assign n29754 = ~n29750 & n29753;
  assign n29755 = ~n29749 & n29754;
  assign n29756 = pi29  & n29755;
  assign n29757 = ~pi29  & ~n29755;
  assign n29758 = ~n29756 & ~n29757;
  assign n29759 = n29748 & ~n29758;
  assign n29760 = ~n29748 & n29758;
  assign n29761 = ~n29759 & ~n29760;
  assign n29762 = n29614 & ~n29654;
  assign n29763 = ~n29655 & ~n29762;
  assign n29764 = n29761 & n29763;
  assign n29765 = ~n29761 & ~n29763;
  assign n29766 = ~n29764 & ~n29765;
  assign n29767 = n4601 & n24607;
  assign n29768 = n4783 & n24676;
  assign n29769 = n4602 & ~n24754;
  assign n29770 = n4801 & n24748;
  assign n29771 = ~n29769 & ~n29770;
  assign n29772 = ~n29768 & n29771;
  assign n29773 = ~n29767 & n29772;
  assign n29774 = pi26  & n29773;
  assign n29775 = ~pi26  & ~n29773;
  assign n29776 = ~n29774 & ~n29775;
  assign n29777 = n29766 & ~n29776;
  assign n29778 = ~n29766 & n29776;
  assign n29779 = ~n29777 & ~n29778;
  assign n29780 = ~n29714 & n29779;
  assign n29781 = n29714 & ~n29779;
  assign n29782 = ~n29780 & ~n29781;
  assign n29783 = n29712 & ~n29782;
  assign n29784 = ~n29712 & n29782;
  assign n29785 = ~n29783 & ~n29784;
  assign n29786 = n29702 & ~n29785;
  assign n29787 = ~n29702 & n29785;
  assign n29788 = ~n29786 & ~n29787;
  assign n29789 = n5435 & n26284;
  assign n29790 = n6055 & n26532;
  assign n29791 = n5429 & ~n26770;
  assign n29792 = n6071 & n26764;
  assign n29793 = ~n29791 & ~n29792;
  assign n29794 = ~n29790 & n29793;
  assign n29795 = ~n29789 & n29794;
  assign n29796 = pi20  & n29795;
  assign n29797 = ~pi20  & ~n29795;
  assign n29798 = ~n29796 & ~n29797;
  assign n29799 = n29788 & ~n29798;
  assign n29800 = ~n29788 & n29798;
  assign n29801 = ~n29799 & ~n29800;
  assign n29802 = n29701 & n29801;
  assign n29803 = ~n29701 & ~n29801;
  assign n29804 = ~n29802 & ~n29803;
  assign n29805 = ~n29691 & ~n29694;
  assign n29806 = n29804 & n29805;
  assign n29807 = ~n29804 & ~n29805;
  assign n29808 = ~n29806 & ~n29807;
  assign n29809 = n29698 & n29808;
  assign n29810 = ~n29698 & ~n29808;
  assign po23  = ~n29809 & ~n29810;
  assign n29812 = n5429 & n26987;
  assign n29813 = n5435 & n26532;
  assign n29814 = n13502 & n26764;
  assign n29815 = ~n29813 & ~n29814;
  assign n29816 = ~n29812 & n29815;
  assign n29817 = pi20  & n29816;
  assign n29818 = ~pi20  & ~n29816;
  assign n29819 = ~n29817 & ~n29818;
  assign n29820 = n29712 & ~n29780;
  assign n29821 = ~n29781 & ~n29820;
  assign n29822 = ~n29819 & n29821;
  assign n29823 = n29819 & ~n29821;
  assign n29824 = ~n29822 & ~n29823;
  assign n29825 = n3478 & n29480;
  assign n29826 = n1341 & n29825;
  assign n29827 = ~n455 & n29826;
  assign n29828 = n4693 & n12908;
  assign n29829 = n1526 & n29828;
  assign n29830 = ~n590 & n29829;
  assign n29831 = n29827 & n29830;
  assign n29832 = n1148 & n27227;
  assign n29833 = ~n537 & n29832;
  assign n29834 = n5061 & n7111;
  assign n29835 = ~n289 & n29834;
  assign n29836 = n29833 & n29835;
  assign n29837 = n29831 & n29836;
  assign n29838 = ~n29732 & n29837;
  assign n29839 = n29732 & ~n29837;
  assign n29840 = ~n29838 & ~n29839;
  assign n29841 = n3641 & n21183;
  assign n29842 = n3740 & n21180;
  assign n29843 = n556 & n24030;
  assign n29844 = n3961 & n21076;
  assign n29845 = ~n29843 & ~n29844;
  assign n29846 = ~n29842 & n29845;
  assign n29847 = ~n29841 & n29846;
  assign n29848 = ~n29840 & n29847;
  assign n29849 = n29840 & ~n29847;
  assign n29850 = ~n29848 & ~n29849;
  assign n29851 = ~n29733 & n29742;
  assign n29852 = ~n29734 & ~n29851;
  assign n29853 = ~n29850 & ~n29852;
  assign n29854 = n29850 & n29852;
  assign n29855 = ~n29853 & ~n29854;
  assign n29856 = ~n29747 & ~n29759;
  assign n29857 = ~n29855 & n29856;
  assign n29858 = n29855 & ~n29856;
  assign n29859 = ~n29857 & ~n29858;
  assign n29860 = n4006 & n21176;
  assign n29861 = n4133 & n21464;
  assign n29862 = n4002 & n24782;
  assign n29863 = n4555 & n24607;
  assign n29864 = ~n29862 & ~n29863;
  assign n29865 = ~n29861 & n29864;
  assign n29866 = ~n29860 & n29865;
  assign n29867 = pi29  & n29866;
  assign n29868 = ~pi29  & ~n29866;
  assign n29869 = ~n29867 & ~n29868;
  assign n29870 = n29859 & n29869;
  assign n29871 = ~n29859 & ~n29869;
  assign n29872 = ~n29870 & ~n29871;
  assign n29873 = n4601 & n24676;
  assign n29874 = n4783 & n24748;
  assign n29875 = n4602 & ~n25529;
  assign n29876 = n4801 & n25521;
  assign n29877 = ~n29875 & ~n29876;
  assign n29878 = ~n29874 & n29877;
  assign n29879 = ~n29873 & n29878;
  assign n29880 = pi26  & n29879;
  assign n29881 = ~pi26  & ~n29879;
  assign n29882 = ~n29880 & ~n29881;
  assign n29883 = ~n29872 & ~n29882;
  assign n29884 = n29872 & n29882;
  assign n29885 = ~n29883 & ~n29884;
  assign n29886 = ~n29764 & n29776;
  assign n29887 = ~n29765 & ~n29886;
  assign n29888 = ~n29885 & ~n29887;
  assign n29889 = n29885 & n29887;
  assign n29890 = ~n29888 & ~n29889;
  assign n29891 = n5238 & n25785;
  assign n29892 = n71 & n26043;
  assign n29893 = n5239 & ~n26290;
  assign n29894 = n5326 & n26284;
  assign n29895 = ~n29893 & ~n29894;
  assign n29896 = ~n29892 & n29895;
  assign n29897 = ~n29891 & n29896;
  assign n29898 = pi23  & n29897;
  assign n29899 = ~pi23  & ~n29897;
  assign n29900 = ~n29898 & ~n29899;
  assign n29901 = n29890 & ~n29900;
  assign n29902 = ~n29890 & n29900;
  assign n29903 = ~n29901 & ~n29902;
  assign n29904 = n29824 & n29903;
  assign n29905 = ~n29824 & ~n29903;
  assign n29906 = ~n29904 & ~n29905;
  assign n29907 = ~n29787 & n29798;
  assign n29908 = ~n29786 & ~n29907;
  assign n29909 = ~n29906 & ~n29908;
  assign n29910 = n29906 & n29908;
  assign n29911 = ~n29909 & ~n29910;
  assign n29912 = ~n29701 & n29801;
  assign n29913 = ~n29807 & ~n29912;
  assign n29914 = ~n29911 & n29913;
  assign n29915 = n29911 & ~n29913;
  assign n29916 = ~n29914 & ~n29915;
  assign n29917 = n29809 & n29916;
  assign n29918 = ~n29809 & ~n29916;
  assign po24  = ~n29917 & ~n29918;
  assign n29920 = ~n29910 & ~n29915;
  assign n29921 = n4601 & n24748;
  assign n29922 = n4783 & n25521;
  assign n29923 = n4602 & n25793;
  assign n29924 = n4801 & n25785;
  assign n29925 = ~n29923 & ~n29924;
  assign n29926 = ~n29922 & n29925;
  assign n29927 = ~n29921 & n29926;
  assign n29928 = pi26  & n29927;
  assign n29929 = ~pi26  & ~n29927;
  assign n29930 = ~n29928 & ~n29929;
  assign n29931 = ~n29854 & ~n29858;
  assign n29932 = ~n13335 & n26764;
  assign n29933 = pi20  & ~n29932;
  assign n29934 = ~pi20  & n29932;
  assign n29935 = ~n29933 & ~n29934;
  assign n29936 = n935 & n3422;
  assign n29937 = n1870 & n29936;
  assign n29938 = n1131 & n29937;
  assign n29939 = n1222 & n14345;
  assign n29940 = n3220 & n29939;
  assign n29941 = ~n595 & n29940;
  assign n29942 = n29938 & n29941;
  assign n29943 = n1617 & n5163;
  assign n29944 = n1011 & n29943;
  assign n29945 = ~n320 & n29944;
  assign n29946 = n491 & n15223;
  assign n29947 = ~n527 & n29946;
  assign n29948 = ~n600 & n29947;
  assign n29949 = n29945 & n29948;
  assign n29950 = n29942 & n29949;
  assign n29951 = n1955 & n29950;
  assign n29952 = n29732 & n29951;
  assign n29953 = ~n29732 & ~n29951;
  assign n29954 = ~n29952 & ~n29953;
  assign n29955 = n29935 & n29954;
  assign n29956 = ~n29935 & ~n29954;
  assign n29957 = ~n29955 & ~n29956;
  assign n29958 = ~n29839 & n29847;
  assign n29959 = ~n29838 & ~n29958;
  assign n29960 = n29957 & n29959;
  assign n29961 = ~n29957 & ~n29959;
  assign n29962 = ~n29960 & ~n29961;
  assign n29963 = n3641 & n21180;
  assign n29964 = n3740 & n21076;
  assign n29965 = n556 & n24012;
  assign n29966 = n3961 & n21176;
  assign n29967 = ~n29965 & ~n29966;
  assign n29968 = ~n29964 & n29967;
  assign n29969 = ~n29963 & n29968;
  assign n29970 = n29962 & ~n29969;
  assign n29971 = ~n29962 & n29969;
  assign n29972 = ~n29970 & ~n29971;
  assign n29973 = n29931 & ~n29972;
  assign n29974 = ~n29931 & n29972;
  assign n29975 = ~n29973 & ~n29974;
  assign n29976 = n4006 & n21464;
  assign n29977 = n4133 & n24607;
  assign n29978 = n4002 & n24770;
  assign n29979 = n4555 & n24676;
  assign n29980 = ~n29978 & ~n29979;
  assign n29981 = ~n29977 & n29980;
  assign n29982 = ~n29976 & n29981;
  assign n29983 = pi29  & n29982;
  assign n29984 = ~pi29  & ~n29982;
  assign n29985 = ~n29983 & ~n29984;
  assign n29986 = n29975 & ~n29985;
  assign n29987 = ~n29975 & n29985;
  assign n29988 = ~n29986 & ~n29987;
  assign n29989 = n29930 & n29988;
  assign n29990 = ~n29930 & ~n29988;
  assign n29991 = ~n29989 & ~n29990;
  assign n29992 = n29859 & ~n29869;
  assign n29993 = ~n29883 & ~n29992;
  assign n29994 = n29991 & n29993;
  assign n29995 = ~n29991 & ~n29993;
  assign n29996 = ~n29994 & ~n29995;
  assign n29997 = n5238 & n26043;
  assign n29998 = n71 & n26284;
  assign n29999 = n5239 & n26540;
  assign n30000 = n5326 & n26532;
  assign n30001 = ~n29999 & ~n30000;
  assign n30002 = ~n29998 & n30001;
  assign n30003 = ~n29997 & n30002;
  assign n30004 = pi23  & n30003;
  assign n30005 = ~pi23  & ~n30003;
  assign n30006 = ~n30004 & ~n30005;
  assign n30007 = ~n29889 & n29900;
  assign n30008 = ~n29888 & ~n30007;
  assign n30009 = n30006 & n30008;
  assign n30010 = ~n30006 & ~n30008;
  assign n30011 = ~n30009 & ~n30010;
  assign n30012 = ~n29996 & n30011;
  assign n30013 = n29996 & ~n30011;
  assign n30014 = ~n30012 & ~n30013;
  assign n30015 = ~n29822 & ~n29903;
  assign n30016 = ~n29823 & ~n30015;
  assign n30017 = n30014 & n30016;
  assign n30018 = ~n30014 & ~n30016;
  assign n30019 = ~n30017 & ~n30018;
  assign n30020 = ~n29920 & n30019;
  assign n30021 = n29920 & ~n30019;
  assign n30022 = ~n30020 & ~n30021;
  assign n30023 = ~n29917 & ~n30022;
  assign n30024 = n29917 & n30022;
  assign po25  = ~n30023 & ~n30024;
  assign n30026 = ~n30006 & n30008;
  assign n30027 = ~n30013 & ~n30026;
  assign n30028 = ~n29930 & n29988;
  assign n30029 = ~n29995 & ~n30028;
  assign n30030 = ~n29953 & ~n29955;
  assign n30031 = n2516 & n4362;
  assign n30032 = ~n672 & n30031;
  assign n30033 = n2375 & n2428;
  assign n30034 = n2467 & n30033;
  assign n30035 = n4698 & n30034;
  assign n30036 = n2066 & n30035;
  assign n30037 = ~n424 & n30036;
  assign n30038 = n30032 & n30037;
  assign n30039 = n5493 & n13877;
  assign n30040 = ~n590 & n30039;
  assign n30041 = n1221 & n15286;
  assign n30042 = ~n246 & n30041;
  assign n30043 = ~n88 & n30042;
  assign n30044 = n30040 & n30043;
  assign n30045 = n30038 & n30044;
  assign n30046 = ~n30030 & n30045;
  assign n30047 = n30030 & ~n30045;
  assign n30048 = ~n30046 & ~n30047;
  assign n30049 = n3641 & n21076;
  assign n30050 = n3740 & n21176;
  assign n30051 = n556 & ~n21470;
  assign n30052 = n3961 & n21464;
  assign n30053 = ~n30051 & ~n30052;
  assign n30054 = ~n30050 & n30053;
  assign n30055 = ~n30049 & n30054;
  assign n30056 = n30048 & ~n30055;
  assign n30057 = ~n30048 & n30055;
  assign n30058 = ~n30056 & ~n30057;
  assign n30059 = ~n29960 & n29969;
  assign n30060 = ~n29961 & ~n30059;
  assign n30061 = ~n30058 & ~n30060;
  assign n30062 = n30058 & n30060;
  assign n30063 = ~n30061 & ~n30062;
  assign n30064 = n4006 & n24607;
  assign n30065 = n4133 & n24676;
  assign n30066 = n4002 & ~n24754;
  assign n30067 = n4555 & n24748;
  assign n30068 = ~n30066 & ~n30067;
  assign n30069 = ~n30065 & n30068;
  assign n30070 = ~n30064 & n30069;
  assign n30071 = pi29  & n30070;
  assign n30072 = ~pi29  & ~n30070;
  assign n30073 = ~n30071 & ~n30072;
  assign n30074 = n30063 & ~n30073;
  assign n30075 = ~n30063 & n30073;
  assign n30076 = ~n30074 & ~n30075;
  assign n30077 = ~n29974 & n29985;
  assign n30078 = ~n29973 & ~n30077;
  assign n30079 = n30076 & n30078;
  assign n30080 = ~n30076 & ~n30078;
  assign n30081 = ~n30079 & ~n30080;
  assign n30082 = n4601 & n25521;
  assign n30083 = n4783 & n25785;
  assign n30084 = n4602 & n26049;
  assign n30085 = n4801 & n26043;
  assign n30086 = ~n30084 & ~n30085;
  assign n30087 = ~n30083 & n30086;
  assign n30088 = ~n30082 & n30087;
  assign n30089 = pi26  & n30088;
  assign n30090 = ~pi26  & ~n30088;
  assign n30091 = ~n30089 & ~n30090;
  assign n30092 = n30081 & ~n30091;
  assign n30093 = ~n30081 & n30091;
  assign n30094 = ~n30092 & ~n30093;
  assign n30095 = n30029 & ~n30094;
  assign n30096 = ~n30029 & n30094;
  assign n30097 = ~n30095 & ~n30096;
  assign n30098 = n5238 & n26284;
  assign n30099 = n71 & n26532;
  assign n30100 = n5239 & ~n26770;
  assign n30101 = n5326 & n26764;
  assign n30102 = ~n30100 & ~n30101;
  assign n30103 = ~n30099 & n30102;
  assign n30104 = ~n30098 & n30103;
  assign n30105 = pi23  & n30104;
  assign n30106 = ~pi23  & ~n30104;
  assign n30107 = ~n30105 & ~n30106;
  assign n30108 = n30097 & ~n30107;
  assign n30109 = ~n30097 & n30107;
  assign n30110 = ~n30108 & ~n30109;
  assign n30111 = n30027 & n30110;
  assign n30112 = ~n30027 & ~n30110;
  assign n30113 = ~n30111 & ~n30112;
  assign n30114 = ~n30017 & ~n30020;
  assign n30115 = n30113 & n30114;
  assign n30116 = ~n30113 & ~n30114;
  assign n30117 = ~n30115 & ~n30116;
  assign n30118 = n30024 & n30117;
  assign n30119 = ~n30024 & ~n30117;
  assign po26  = ~n30118 & ~n30119;
  assign n30121 = n5239 & n26987;
  assign n30122 = n5238 & n26532;
  assign n30123 = ~n21080 & n26764;
  assign n30124 = ~n30122 & ~n30123;
  assign n30125 = ~n30121 & n30124;
  assign n30126 = pi23  & n30125;
  assign n30127 = ~pi23  & ~n30125;
  assign n30128 = ~n30126 & ~n30127;
  assign n30129 = ~n30079 & n30091;
  assign n30130 = ~n30080 & ~n30129;
  assign n30131 = ~n30128 & n30130;
  assign n30132 = n30128 & ~n30130;
  assign n30133 = ~n30131 & ~n30132;
  assign n30134 = ~n30062 & ~n30074;
  assign n30135 = ~n428 & n476;
  assign n30136 = n1976 & n3806;
  assign n30137 = n1148 & n30136;
  assign n30138 = n1163 & n15153;
  assign n30139 = n1401 & n30138;
  assign n30140 = n2066 & n30139;
  assign n30141 = n30137 & n30140;
  assign n30142 = ~n299 & n30141;
  assign n30143 = n22283 & n28053;
  assign n30144 = ~n310 & n30143;
  assign n30145 = n12574 & n24547;
  assign n30146 = ~n231 & n30145;
  assign n30147 = n30144 & n30146;
  assign n30148 = n30142 & n30147;
  assign n30149 = n30135 & n30148;
  assign n30150 = n30045 & ~n30149;
  assign n30151 = ~n30045 & n30149;
  assign n30152 = ~n30150 & ~n30151;
  assign n30153 = ~n30046 & n30055;
  assign n30154 = ~n30047 & ~n30153;
  assign n30155 = n30152 & ~n30154;
  assign n30156 = ~n30152 & n30154;
  assign n30157 = ~n30155 & ~n30156;
  assign n30158 = n3641 & n21176;
  assign n30159 = n3740 & n21464;
  assign n30160 = n556 & n24782;
  assign n30161 = n3961 & n24607;
  assign n30162 = ~n30160 & ~n30161;
  assign n30163 = ~n30159 & n30162;
  assign n30164 = ~n30158 & n30163;
  assign n30165 = ~n30157 & ~n30164;
  assign n30166 = n30157 & n30164;
  assign n30167 = ~n30165 & ~n30166;
  assign n30168 = n30134 & ~n30167;
  assign n30169 = ~n30134 & n30167;
  assign n30170 = ~n30168 & ~n30169;
  assign n30171 = n4006 & n24676;
  assign n30172 = n4133 & n24748;
  assign n30173 = n4002 & ~n25529;
  assign n30174 = n4555 & n25521;
  assign n30175 = ~n30173 & ~n30174;
  assign n30176 = ~n30172 & n30175;
  assign n30177 = ~n30171 & n30176;
  assign n30178 = pi29  & n30177;
  assign n30179 = ~pi29  & ~n30177;
  assign n30180 = ~n30178 & ~n30179;
  assign n30181 = n30170 & n30180;
  assign n30182 = ~n30170 & ~n30180;
  assign n30183 = ~n30181 & ~n30182;
  assign n30184 = n4601 & n25785;
  assign n30185 = n4783 & n26043;
  assign n30186 = n4602 & ~n26290;
  assign n30187 = n4801 & n26284;
  assign n30188 = ~n30186 & ~n30187;
  assign n30189 = ~n30185 & n30188;
  assign n30190 = ~n30184 & n30189;
  assign n30191 = pi26  & n30190;
  assign n30192 = ~pi26  & ~n30190;
  assign n30193 = ~n30191 & ~n30192;
  assign n30194 = ~n30183 & ~n30193;
  assign n30195 = n30183 & n30193;
  assign n30196 = ~n30194 & ~n30195;
  assign n30197 = n30133 & n30196;
  assign n30198 = ~n30133 & ~n30196;
  assign n30199 = ~n30197 & ~n30198;
  assign n30200 = ~n30096 & n30107;
  assign n30201 = ~n30095 & ~n30200;
  assign n30202 = ~n30199 & ~n30201;
  assign n30203 = n30199 & n30201;
  assign n30204 = ~n30202 & ~n30203;
  assign n30205 = ~n30027 & n30110;
  assign n30206 = ~n30116 & ~n30205;
  assign n30207 = ~n30204 & n30206;
  assign n30208 = n30204 & ~n30206;
  assign n30209 = ~n30207 & ~n30208;
  assign n30210 = n30118 & n30209;
  assign n30211 = ~n30118 & ~n30209;
  assign po27  = ~n30210 & ~n30211;
  assign n30213 = ~n30203 & ~n30208;
  assign n30214 = n30170 & ~n30180;
  assign n30215 = ~n30194 & ~n30214;
  assign n30216 = n4601 & n26043;
  assign n30217 = n4783 & n26284;
  assign n30218 = n4602 & n26540;
  assign n30219 = n4801 & n26532;
  assign n30220 = ~n30218 & ~n30219;
  assign n30221 = ~n30217 & n30220;
  assign n30222 = ~n30216 & n30221;
  assign n30223 = pi26  & n30222;
  assign n30224 = ~pi26  & ~n30222;
  assign n30225 = ~n30223 & ~n30224;
  assign n30226 = ~n30215 & n30225;
  assign n30227 = n30215 & ~n30225;
  assign n30228 = ~n30226 & ~n30227;
  assign n30229 = ~n30165 & ~n30169;
  assign n30230 = ~n21396 & n26764;
  assign n30231 = pi23  & ~n30230;
  assign n30232 = ~pi23  & n30230;
  assign n30233 = ~n30231 & ~n30232;
  assign n30234 = ~n197 & n5475;
  assign n30235 = ~n395 & n30234;
  assign n30236 = n119 & n369;
  assign n30237 = ~n104 & n30236;
  assign n30238 = n30235 & n30237;
  assign n30239 = n263 & n710;
  assign n30240 = n546 & n30239;
  assign n30241 = ~n144 & n30240;
  assign n30242 = n1252 & n3717;
  assign n30243 = n797 & n30242;
  assign n30244 = ~n536 & n30243;
  assign n30245 = ~n132 & n30244;
  assign n30246 = n30241 & n30245;
  assign n30247 = n30238 & n30246;
  assign n30248 = n30149 & n30247;
  assign n30249 = ~n30149 & ~n30247;
  assign n30250 = ~n30248 & ~n30249;
  assign n30251 = n30233 & n30250;
  assign n30252 = ~n30233 & ~n30250;
  assign n30253 = ~n30251 & ~n30252;
  assign n30254 = ~n30151 & ~n30154;
  assign n30255 = ~n30150 & ~n30254;
  assign n30256 = n30253 & n30255;
  assign n30257 = ~n30253 & ~n30255;
  assign n30258 = ~n30256 & ~n30257;
  assign n30259 = n3641 & n21464;
  assign n30260 = n3740 & n24607;
  assign n30261 = n556 & n24770;
  assign n30262 = n3961 & n24676;
  assign n30263 = ~n30261 & ~n30262;
  assign n30264 = ~n30260 & n30263;
  assign n30265 = ~n30259 & n30264;
  assign n30266 = n30258 & ~n30265;
  assign n30267 = ~n30258 & n30265;
  assign n30268 = ~n30266 & ~n30267;
  assign n30269 = n30229 & ~n30268;
  assign n30270 = ~n30229 & n30268;
  assign n30271 = ~n30269 & ~n30270;
  assign n30272 = n4006 & n24748;
  assign n30273 = n4133 & n25521;
  assign n30274 = n4002 & n25793;
  assign n30275 = n4555 & n25785;
  assign n30276 = ~n30274 & ~n30275;
  assign n30277 = ~n30273 & n30276;
  assign n30278 = ~n30272 & n30277;
  assign n30279 = pi29  & n30278;
  assign n30280 = ~pi29  & ~n30278;
  assign n30281 = ~n30279 & ~n30280;
  assign n30282 = n30271 & ~n30281;
  assign n30283 = ~n30271 & n30281;
  assign n30284 = ~n30282 & ~n30283;
  assign n30285 = ~n30228 & n30284;
  assign n30286 = n30228 & ~n30284;
  assign n30287 = ~n30285 & ~n30286;
  assign n30288 = ~n30131 & ~n30196;
  assign n30289 = ~n30132 & ~n30288;
  assign n30290 = n30287 & n30289;
  assign n30291 = ~n30287 & ~n30289;
  assign n30292 = ~n30290 & ~n30291;
  assign n30293 = ~n30213 & n30292;
  assign n30294 = n30213 & ~n30292;
  assign n30295 = ~n30293 & ~n30294;
  assign n30296 = ~n30210 & ~n30295;
  assign n30297 = n30210 & n30295;
  assign po28  = ~n30296 & ~n30297;
  assign n30299 = ~n30290 & ~n30293;
  assign n30300 = ~n30215 & ~n30225;
  assign n30301 = ~n30285 & ~n30300;
  assign n30302 = ~n30249 & ~n30251;
  assign n30303 = n348 & n14304;
  assign n30304 = n2021 & n30303;
  assign n30305 = ~n246 & n30304;
  assign n30306 = n998 & n7134;
  assign n30307 = n2474 & n30306;
  assign n30308 = n276 & n30307;
  assign n30309 = ~n320 & n30308;
  assign n30310 = n30305 & n30309;
  assign n30311 = n467 & n730;
  assign n30312 = n2180 & n30311;
  assign n30313 = ~n427 & n30312;
  assign n30314 = n15149 & n24708;
  assign n30315 = n1340 & n30314;
  assign n30316 = ~n474 & n30315;
  assign n30317 = n30313 & n30316;
  assign n30318 = n30310 & n30317;
  assign n30319 = ~n30302 & n30318;
  assign n30320 = n30302 & ~n30318;
  assign n30321 = ~n30319 & ~n30320;
  assign n30322 = n3641 & n24607;
  assign n30323 = n3740 & n24676;
  assign n30324 = n556 & ~n24754;
  assign n30325 = n3961 & n24748;
  assign n30326 = ~n30324 & ~n30325;
  assign n30327 = ~n30323 & n30326;
  assign n30328 = ~n30322 & n30327;
  assign n30329 = n30321 & ~n30328;
  assign n30330 = ~n30321 & n30328;
  assign n30331 = ~n30329 & ~n30330;
  assign n30332 = ~n30256 & n30265;
  assign n30333 = ~n30257 & ~n30332;
  assign n30334 = ~n30331 & ~n30333;
  assign n30335 = n30331 & n30333;
  assign n30336 = ~n30334 & ~n30335;
  assign n30337 = n4006 & n25521;
  assign n30338 = n4133 & n25785;
  assign n30339 = n4002 & n26049;
  assign n30340 = n4555 & n26043;
  assign n30341 = ~n30339 & ~n30340;
  assign n30342 = ~n30338 & n30341;
  assign n30343 = ~n30337 & n30342;
  assign n30344 = pi29  & n30343;
  assign n30345 = ~pi29  & ~n30343;
  assign n30346 = ~n30344 & ~n30345;
  assign n30347 = n30336 & ~n30346;
  assign n30348 = ~n30336 & n30346;
  assign n30349 = ~n30347 & ~n30348;
  assign n30350 = ~n30270 & n30281;
  assign n30351 = ~n30269 & ~n30350;
  assign n30352 = n30349 & n30351;
  assign n30353 = ~n30349 & ~n30351;
  assign n30354 = ~n30352 & ~n30353;
  assign n30355 = n4601 & n26284;
  assign n30356 = n4783 & n26532;
  assign n30357 = n4602 & ~n26770;
  assign n30358 = n4801 & n26764;
  assign n30359 = ~n30357 & ~n30358;
  assign n30360 = ~n30356 & n30359;
  assign n30361 = ~n30355 & n30360;
  assign n30362 = pi26  & n30361;
  assign n30363 = ~pi26  & ~n30361;
  assign n30364 = ~n30362 & ~n30363;
  assign n30365 = n30354 & ~n30364;
  assign n30366 = ~n30354 & n30364;
  assign n30367 = ~n30365 & ~n30366;
  assign n30368 = ~n30301 & n30367;
  assign n30369 = n30301 & ~n30367;
  assign n30370 = ~n30368 & ~n30369;
  assign n30371 = n30299 & ~n30370;
  assign n30372 = ~n30299 & n30370;
  assign n30373 = ~n30371 & ~n30372;
  assign n30374 = n30297 & n30373;
  assign n30375 = ~n30297 & ~n30373;
  assign po29  = ~n30374 & ~n30375;
  assign n30377 = ~n30368 & ~n30372;
  assign n30378 = ~n30335 & ~n30347;
  assign n30379 = n3650 & n24708;
  assign n30380 = ~n104 & n30379;
  assign n30381 = n451 & n553;
  assign n30382 = n138 & n407;
  assign n30383 = n30381 & n30382;
  assign n30384 = n319 & n30383;
  assign n30385 = n30380 & n30384;
  assign n30386 = ~n30318 & n30385;
  assign n30387 = n30318 & ~n30385;
  assign n30388 = ~n30386 & ~n30387;
  assign n30389 = ~n30319 & n30328;
  assign n30390 = ~n30320 & ~n30389;
  assign n30391 = n30388 & ~n30390;
  assign n30392 = ~n30388 & n30390;
  assign n30393 = ~n30391 & ~n30392;
  assign n30394 = n3641 & n24676;
  assign n30395 = n3740 & n24748;
  assign n30396 = n556 & ~n25529;
  assign n30397 = n3961 & n25521;
  assign n30398 = ~n30396 & ~n30397;
  assign n30399 = ~n30395 & n30398;
  assign n30400 = ~n30394 & n30399;
  assign n30401 = ~n30393 & ~n30400;
  assign n30402 = n30393 & n30400;
  assign n30403 = ~n30401 & ~n30402;
  assign n30404 = n30378 & ~n30403;
  assign n30405 = ~n30378 & n30403;
  assign n30406 = ~n30404 & ~n30405;
  assign n30407 = n4602 & n26987;
  assign n30408 = n4601 & n26532;
  assign n30409 = ~n24646 & n26764;
  assign n30410 = ~n30408 & ~n30409;
  assign n30411 = ~n30407 & n30410;
  assign n30412 = ~pi26  & ~n30411;
  assign n30413 = pi26  & n30411;
  assign n30414 = ~n30412 & ~n30413;
  assign n30415 = n4006 & n25785;
  assign n30416 = n4133 & n26043;
  assign n30417 = n4002 & ~n26290;
  assign n30418 = n4555 & n26284;
  assign n30419 = ~n30417 & ~n30418;
  assign n30420 = ~n30416 & n30419;
  assign n30421 = ~n30415 & n30420;
  assign n30422 = pi29  & n30421;
  assign n30423 = ~pi29  & ~n30421;
  assign n30424 = ~n30422 & ~n30423;
  assign n30425 = ~n30414 & n30424;
  assign n30426 = n30414 & ~n30424;
  assign n30427 = ~n30425 & ~n30426;
  assign n30428 = ~n30406 & n30427;
  assign n30429 = n30406 & ~n30427;
  assign n30430 = ~n30428 & ~n30429;
  assign n30431 = ~n30352 & n30364;
  assign n30432 = ~n30353 & ~n30431;
  assign n30433 = n30430 & n30432;
  assign n30434 = ~n30430 & ~n30432;
  assign n30435 = ~n30433 & ~n30434;
  assign n30436 = ~n30377 & n30435;
  assign n30437 = n30377 & ~n30435;
  assign n30438 = ~n30436 & ~n30437;
  assign n30439 = ~n30374 & ~n30438;
  assign n30440 = n30374 & n30438;
  assign po30  = ~n30439 & ~n30440;
  assign n30442 = ~n24703 & n26764;
  assign n30443 = n30440 & ~n30442;
  assign n30444 = ~n30440 & n30442;
  assign n30445 = ~n30443 & ~n30444;
  assign n30446 = ~n30414 & ~n30424;
  assign n30447 = ~n30429 & ~n30446;
  assign n30448 = ~n30433 & ~n30436;
  assign n30449 = n30318 & ~n30448;
  assign n30450 = ~n30318 & n30448;
  assign n30451 = ~n30449 & ~n30450;
  assign n30452 = n30447 & n30451;
  assign n30453 = ~n30447 & ~n30451;
  assign n30454 = ~n30452 & ~n30453;
  assign n30455 = n525 & n717;
  assign n30456 = pi26  & ~n30455;
  assign n30457 = ~pi26  & n30455;
  assign n30458 = ~n30456 & ~n30457;
  assign n30459 = ~n30401 & ~n30405;
  assign n30460 = ~n30387 & ~n30390;
  assign n30461 = ~n30386 & ~n30460;
  assign n30462 = n30459 & ~n30461;
  assign n30463 = ~n30459 & n30461;
  assign n30464 = ~n30462 & ~n30463;
  assign n30465 = n4006 & n26043;
  assign n30466 = n4133 & n26284;
  assign n30467 = n4002 & n26540;
  assign n30468 = n4555 & n26532;
  assign n30469 = ~n30467 & ~n30468;
  assign n30470 = ~n30466 & n30469;
  assign n30471 = ~n30465 & n30470;
  assign n30472 = pi29  & ~n30471;
  assign n30473 = ~pi29  & n30471;
  assign n30474 = ~n30472 & ~n30473;
  assign n30475 = n3641 & n24748;
  assign n30476 = n3740 & n25521;
  assign n30477 = n556 & n25793;
  assign n30478 = n3961 & n25785;
  assign n30479 = ~n30477 & ~n30478;
  assign n30480 = ~n30476 & n30479;
  assign n30481 = ~n30475 & n30480;
  assign n30482 = n30474 & ~n30481;
  assign n30483 = ~n30474 & n30481;
  assign n30484 = ~n30482 & ~n30483;
  assign n30485 = n30464 & n30484;
  assign n30486 = ~n30464 & ~n30484;
  assign n30487 = ~n30485 & ~n30486;
  assign n30488 = n30458 & ~n30487;
  assign n30489 = ~n30458 & n30487;
  assign n30490 = ~n30488 & ~n30489;
  assign n30491 = n30454 & ~n30490;
  assign n30492 = ~n30454 & n30490;
  assign n30493 = ~n30491 & ~n30492;
  assign n30494 = n30445 & n30493;
  assign n30495 = ~n30445 & ~n30493;
  assign po31  = ~n30494 & ~n30495;
endmodule
