module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n405, n406, n407, n408, n409, n410, n412,
    n413, n414, n415, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n498,
    n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n583,
    n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n632, n633,
    n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n669,
    n670, n671, n672;
  assign n22 = ~pi3  & ~pi5 ;
  assign n23 = ~pi1  & pi9 ;
  assign n24 = ~pi0  & pi9 ;
  assign n25 = pi1  & ~n24;
  assign n26 = ~n23 & ~n25;
  assign n27 = n22 & n26;
  assign n28 = pi0  & ~pi9 ;
  assign n29 = ~pi1  & ~n28;
  assign n30 = pi1  & ~pi9 ;
  assign n31 = ~pi7  & ~n30;
  assign n32 = ~n29 & n31;
  assign n33 = ~n27 & ~n32;
  assign n34 = ~pi2  & ~n33;
  assign n35 = ~pi2  & ~pi5 ;
  assign n36 = ~pi0  & ~n35;
  assign n37 = pi1  & pi2 ;
  assign n38 = ~n36 & ~n37;
  assign n39 = ~pi9  & ~n38;
  assign n40 = ~pi2  & ~pi3 ;
  assign n41 = pi9  & ~n40;
  assign n42 = pi0  & pi3 ;
  assign n43 = ~n41 & ~n42;
  assign n44 = ~pi1  & ~n43;
  assign n45 = pi1  & ~pi3 ;
  assign n46 = ~n44 & ~n45;
  assign n47 = ~n39 & n46;
  assign n48 = ~pi7  & ~n47;
  assign n49 = ~n34 & ~n48;
  assign n50 = ~pi8  & ~n49;
  assign n51 = pi7  & pi8 ;
  assign n52 = ~pi5  & n51;
  assign n53 = ~pi7  & pi9 ;
  assign n54 = ~n52 & ~n53;
  assign n55 = pi1  & ~n54;
  assign n56 = pi1  & ~pi7 ;
  assign n57 = ~pi5  & ~pi9 ;
  assign n58 = ~n56 & n57;
  assign n59 = ~n55 & ~n58;
  assign n60 = pi0  & ~pi2 ;
  assign n61 = ~n59 & n60;
  assign n62 = pi2  & ~pi9 ;
  assign n63 = ~pi0  & ~pi1 ;
  assign n64 = n62 & n63;
  assign n65 = n52 & n64;
  assign n66 = ~n61 & ~n65;
  assign n67 = ~pi3  & ~n66;
  assign n68 = ~n50 & ~n67;
  assign n69 = ~pi6  & ~n68;
  assign n70 = ~n24 & ~n28;
  assign n71 = pi1  & n70;
  assign n72 = pi2  & n71;
  assign n73 = pi5  & n72;
  assign n74 = pi5  & pi6 ;
  assign n75 = pi6  & pi9 ;
  assign n76 = ~pi1  & ~pi2 ;
  assign n77 = ~pi0  & n76;
  assign n78 = n75 & n77;
  assign n79 = ~n74 & ~n78;
  assign n80 = ~n73 & n79;
  assign n81 = pi8  & ~n80;
  assign n82 = ~pi1  & ~n24;
  assign n83 = ~pi8  & ~n82;
  assign n84 = ~pi1  & pi2 ;
  assign n85 = n28 & n84;
  assign n86 = ~n83 & ~n85;
  assign n87 = ~pi5  & ~n86;
  assign n88 = ~n81 & ~n87;
  assign n89 = pi3  & ~n88;
  assign n90 = ~pi2  & ~n28;
  assign n91 = pi6  & ~n90;
  assign n92 = n40 & n71;
  assign n93 = ~n91 & ~n92;
  assign n94 = pi5  & ~n93;
  assign n95 = pi2  & pi9 ;
  assign n96 = ~pi2  & n30;
  assign n97 = ~n95 & ~n96;
  assign n98 = ~pi0  & ~pi3 ;
  assign n99 = ~n97 & n98;
  assign n100 = pi6  & n99;
  assign n101 = ~n94 & ~n100;
  assign n102 = pi8  & ~n101;
  assign n103 = pi2  & ~pi3 ;
  assign n104 = n23 & n103;
  assign n105 = pi1  & ~pi8 ;
  assign n106 = ~n104 & ~n105;
  assign n107 = ~pi0  & ~n106;
  assign n108 = ~pi1  & ~pi9 ;
  assign n109 = pi3  & ~pi6 ;
  assign n110 = pi2  & pi3 ;
  assign n111 = ~n109 & ~n110;
  assign n112 = n108 & n111;
  assign n113 = ~n95 & ~n112;
  assign n114 = ~pi8  & ~n113;
  assign n115 = ~n107 & ~n114;
  assign n116 = ~pi5  & ~n115;
  assign n117 = ~pi3  & ~pi8 ;
  assign n118 = pi1  & pi9 ;
  assign n119 = ~n108 & ~n118;
  assign n120 = n117 & ~n119;
  assign n121 = n77 & n120;
  assign n122 = ~n116 & ~n121;
  assign n123 = ~n102 & n122;
  assign n124 = ~n89 & n123;
  assign n125 = ~pi7  & ~n124;
  assign n126 = ~n69 & ~n125;
  assign n127 = ~pi4  & ~n126;
  assign n128 = ~pi8  & ~pi9 ;
  assign n129 = ~pi6  & n128;
  assign n130 = pi4  & pi8 ;
  assign n131 = pi6  & n130;
  assign n132 = ~n129 & ~n131;
  assign n133 = pi5  & ~n132;
  assign n134 = pi6  & ~pi9 ;
  assign n135 = pi4  & pi9 ;
  assign n136 = ~n134 & ~n135;
  assign n137 = ~n74 & ~n136;
  assign n138 = ~pi8  & n137;
  assign n139 = ~n133 & ~n138;
  assign n140 = ~pi7  & ~n139;
  assign n141 = ~pi1  & ~pi3 ;
  assign n142 = ~pi2  & n141;
  assign n143 = n140 & n142;
  assign n144 = ~pi0  & n143;
  assign po0  = n127 | n144;
  assign n146 = ~pi5  & pi8 ;
  assign n147 = ~n75 & ~n146;
  assign n148 = ~pi0  & ~n147;
  assign n149 = pi8  & n75;
  assign n150 = ~pi8  & n57;
  assign n151 = ~n149 & ~n150;
  assign n152 = ~n148 & n151;
  assign n153 = pi2  & ~n152;
  assign n154 = pi8  & pi9 ;
  assign n155 = pi0  & n154;
  assign n156 = ~n128 & ~n155;
  assign n157 = pi5  & ~n156;
  assign n158 = ~n60 & ~n62;
  assign n159 = n157 & n158;
  assign n160 = ~n153 & ~n159;
  assign n161 = ~pi4  & ~n160;
  assign n162 = ~pi0  & ~pi2 ;
  assign n163 = ~pi6  & pi9 ;
  assign n164 = pi5  & ~pi8 ;
  assign n165 = ~n130 & ~n164;
  assign n166 = ~pi6  & ~n165;
  assign n167 = ~n135 & ~n166;
  assign n168 = ~n163 & ~n167;
  assign n169 = n162 & n168;
  assign n170 = ~n161 & ~n169;
  assign n171 = ~pi1  & ~n170;
  assign n172 = pi6  & pi8 ;
  assign n173 = ~n147 & ~n172;
  assign n174 = pi0  & n173;
  assign n175 = ~pi0  & pi5 ;
  assign n176 = ~pi8  & pi9 ;
  assign n177 = n175 & n176;
  assign n178 = ~n174 & ~n177;
  assign n179 = ~pi2  & ~n178;
  assign n180 = ~pi6  & ~pi8 ;
  assign n181 = pi2  & ~pi5 ;
  assign n182 = ~pi6  & ~n181;
  assign n183 = ~n60 & n146;
  assign n184 = ~n182 & n183;
  assign n185 = ~n180 & ~n184;
  assign n186 = ~pi9  & ~n185;
  assign n187 = ~n179 & ~n186;
  assign n188 = pi1  & ~n187;
  assign n189 = ~pi6  & pi8 ;
  assign n190 = n62 & n189;
  assign n191 = ~n188 & ~n190;
  assign n192 = ~pi4  & ~n191;
  assign n193 = ~n171 & ~n192;
  assign n194 = ~pi3  & ~n193;
  assign n195 = ~pi2  & ~pi8 ;
  assign n196 = pi5  & n195;
  assign n197 = ~n117 & ~n146;
  assign n198 = pi0  & n197;
  assign n199 = ~n196 & ~n198;
  assign n200 = ~pi1  & ~n199;
  assign n201 = ~n40 & ~n195;
  assign n202 = ~pi0  & n201;
  assign n203 = ~pi2  & pi8 ;
  assign n204 = pi0  & n203;
  assign n205 = pi0  & ~pi5 ;
  assign n206 = ~n175 & ~n205;
  assign n207 = ~n204 & n206;
  assign n208 = pi1  & ~n207;
  assign n209 = ~n202 & ~n208;
  assign n210 = ~n200 & n209;
  assign n211 = ~pi6  & ~n210;
  assign n212 = ~pi1  & pi6 ;
  assign n213 = pi2  & ~n212;
  assign n214 = ~pi1  & ~pi8 ;
  assign n215 = ~n213 & ~n214;
  assign n216 = pi3  & n215;
  assign n217 = ~pi0  & pi8 ;
  assign n218 = ~pi1  & ~pi6 ;
  assign n219 = pi0  & pi1 ;
  assign n220 = ~n218 & ~n219;
  assign n221 = ~n217 & n220;
  assign n222 = ~pi2  & n221;
  assign n223 = ~n216 & ~n222;
  assign n224 = ~pi5  & ~n223;
  assign n225 = ~n211 & ~n224;
  assign n226 = ~pi9  & ~n225;
  assign n227 = pi1  & pi5 ;
  assign n228 = pi3  & ~pi8 ;
  assign n229 = n76 & n228;
  assign n230 = ~n227 & ~n229;
  assign n231 = pi0  & ~n230;
  assign n232 = pi5  & ~n40;
  assign n233 = pi3  & n37;
  assign n234 = ~n232 & ~n233;
  assign n235 = ~n231 & n234;
  assign n236 = pi6  & ~n235;
  assign n237 = n164 & n233;
  assign n238 = ~n236 & ~n237;
  assign n239 = pi9  & ~n238;
  assign n240 = ~n226 & ~n239;
  assign n241 = ~pi4  & ~n240;
  assign n242 = ~n194 & ~n241;
  assign n243 = ~pi7  & ~n242;
  assign n244 = pi2  & ~n63;
  assign n245 = n90 & ~n219;
  assign n246 = ~n244 & ~n245;
  assign n247 = ~pi8  & n246;
  assign n248 = n30 & n203;
  assign n249 = ~n247 & ~n248;
  assign n250 = pi7  & ~n249;
  assign n251 = ~n64 & ~n250;
  assign n252 = ~pi4  & ~n251;
  assign n253 = ~pi6  & n252;
  assign n254 = n22 & n253;
  assign po1  = n243 | n254;
  assign n256 = ~pi3  & pi9 ;
  assign n257 = ~n45 & ~n176;
  assign n258 = ~n256 & ~n257;
  assign n259 = ~pi6  & n258;
  assign n260 = pi3  & ~n203;
  assign n261 = pi5  & ~n260;
  assign n262 = pi3  & ~n181;
  assign n263 = pi8  & ~n262;
  assign n264 = ~n261 & ~n263;
  assign n265 = pi1  & ~n264;
  assign n266 = ~pi5  & pi6 ;
  assign n267 = ~pi8  & n266;
  assign n268 = n141 & n267;
  assign n269 = ~n265 & ~n268;
  assign n270 = ~pi9  & ~n269;
  assign n271 = ~pi1  & n201;
  assign n272 = pi2  & ~n189;
  assign n273 = ~n271 & ~n272;
  assign n274 = pi5  & ~n273;
  assign n275 = pi6  & ~pi8 ;
  assign n276 = ~n212 & ~n275;
  assign n277 = ~pi9  & n276;
  assign n278 = ~pi2  & ~n277;
  assign n279 = ~pi1  & n176;
  assign n280 = ~n278 & ~n279;
  assign n281 = pi3  & ~n280;
  assign n282 = pi6  & ~n23;
  assign n283 = pi8  & ~n30;
  assign n284 = n282 & ~n283;
  assign n285 = n256 & n284;
  assign n286 = ~n281 & ~n285;
  assign n287 = ~n274 & n286;
  assign n288 = ~n270 & n287;
  assign n289 = ~n259 & n288;
  assign n290 = ~pi4  & ~n289;
  assign n291 = ~n154 & ~n275;
  assign n292 = ~pi5  & ~n291;
  assign n293 = ~pi3  & pi4 ;
  assign n294 = ~pi1  & n293;
  assign n295 = ~n292 & n294;
  assign n296 = ~pi2  & n295;
  assign n297 = ~n290 & ~n296;
  assign n298 = ~pi0  & ~n297;
  assign n299 = ~pi5  & n95;
  assign n300 = ~n157 & ~n299;
  assign n301 = pi1  & ~n300;
  assign n302 = ~n128 & ~n154;
  assign n303 = ~n108 & ~n302;
  assign n304 = pi2  & ~n303;
  assign n305 = ~n301 & ~n304;
  assign n306 = ~pi3  & ~n305;
  assign n307 = ~pi1  & pi8 ;
  assign n308 = n41 & n307;
  assign n309 = ~n35 & ~n229;
  assign n310 = n128 & ~n309;
  assign n311 = ~n308 & ~n310;
  assign n312 = pi0  & ~n311;
  assign n313 = ~n306 & ~n312;
  assign n314 = ~pi6  & ~n313;
  assign n315 = pi2  & n118;
  assign n316 = ~n307 & ~n315;
  assign n317 = pi6  & ~n316;
  assign n318 = pi2  & n302;
  assign n319 = ~n195 & ~n318;
  assign n320 = ~n317 & ~n319;
  assign n321 = pi3  & ~n320;
  assign n322 = ~n30 & ~n282;
  assign n323 = pi8  & ~n322;
  assign n324 = ~n120 & ~n323;
  assign n325 = ~pi2  & ~n324;
  assign n326 = ~n321 & ~n325;
  assign n327 = n205 & ~n326;
  assign n328 = ~n314 & ~n327;
  assign n329 = ~pi4  & ~n328;
  assign n330 = ~n298 & ~n329;
  assign n331 = ~pi7  & ~n330;
  assign n332 = ~pi5  & ~pi6 ;
  assign n333 = n28 & n214;
  assign n334 = ~n53 & ~n176;
  assign n335 = n71 & n334;
  assign n336 = ~n333 & ~n335;
  assign n337 = ~pi4  & ~n336;
  assign n338 = n40 & n337;
  assign n339 = n332 & n338;
  assign po2  = n331 | n339;
  assign n341 = pi3  & ~n163;
  assign n342 = pi2  & pi6 ;
  assign n343 = ~n341 & ~n342;
  assign n344 = ~pi4  & ~n343;
  assign n345 = n154 & n332;
  assign n346 = ~n74 & ~n345;
  assign n347 = ~pi2  & n293;
  assign n348 = ~n346 & n347;
  assign n349 = ~n344 & ~n348;
  assign n350 = ~pi1  & ~n349;
  assign n351 = pi5  & pi8 ;
  assign n352 = n163 & n351;
  assign n353 = ~n150 & ~n352;
  assign n354 = pi2  & ~n353;
  assign n355 = ~pi6  & ~n228;
  assign n356 = pi3  & ~pi5 ;
  assign n357 = ~n355 & ~n356;
  assign n358 = pi3  & ~n357;
  assign n359 = ~n267 & ~n358;
  assign n360 = ~n354 & n359;
  assign n361 = pi1  & ~n360;
  assign n362 = pi2  & n266;
  assign n363 = ~n361 & ~n362;
  assign n364 = ~pi4  & ~n363;
  assign n365 = ~n350 & ~n364;
  assign n366 = ~pi0  & ~n365;
  assign n367 = pi2  & ~n197;
  assign n368 = ~pi2  & n351;
  assign n369 = ~n367 & ~n368;
  assign n370 = ~pi9  & ~n369;
  assign n371 = ~pi2  & pi3 ;
  assign n372 = pi9  & n196;
  assign n373 = ~n371 & ~n372;
  assign n374 = ~n357 & n373;
  assign n375 = ~n370 & n374;
  assign n376 = pi1  & ~n375;
  assign n377 = ~pi3  & n266;
  assign n378 = n196 & n218;
  assign n379 = ~n377 & ~n378;
  assign n380 = ~pi9  & ~n379;
  assign n381 = ~n376 & ~n380;
  assign n382 = pi0  & ~n381;
  assign n383 = pi2  & n109;
  assign n384 = ~n266 & ~n383;
  assign n385 = n41 & ~n384;
  assign n386 = n147 & ~n355;
  assign n387 = n346 & n386;
  assign n388 = ~n385 & ~n387;
  assign n389 = ~pi1  & ~n388;
  assign n390 = ~n57 & ~n180;
  assign n391 = ~pi2  & ~n390;
  assign n392 = pi5  & pi9 ;
  assign n393 = ~pi6  & ~n392;
  assign n394 = ~n118 & ~n351;
  assign n395 = n393 & ~n394;
  assign n396 = ~n391 & ~n395;
  assign n397 = pi3  & ~n396;
  assign n398 = n266 & n277;
  assign n399 = ~n397 & ~n398;
  assign n400 = ~n389 & n399;
  assign n401 = ~n382 & n400;
  assign n402 = ~pi4  & ~n401;
  assign n403 = ~n366 & ~n402;
  assign po3  = ~pi7  & ~n403;
  assign n405 = ~pi4  & n244;
  assign n406 = pi3  & ~pi4 ;
  assign n407 = ~n293 & ~n406;
  assign n408 = n77 & ~n407;
  assign n409 = ~n405 & ~n408;
  assign n410 = ~pi7  & ~n409;
  assign po4  = n74 & n410;
  assign n412 = ~n77 & n406;
  assign n413 = pi4  & n408;
  assign n414 = ~n412 & ~n413;
  assign n415 = ~pi7  & ~n414;
  assign po5  = n74 & n415;
  assign n417 = ~pi1  & ~pi5 ;
  assign n418 = pi2  & ~n417;
  assign n419 = ~pi9  & ~n418;
  assign n420 = ~pi6  & n419;
  assign n421 = pi5  & n118;
  assign n422 = ~n420 & ~n421;
  assign n423 = pi0  & ~n422;
  assign n424 = ~pi0  & ~n57;
  assign n425 = pi2  & n424;
  assign n426 = ~n423 & ~n425;
  assign n427 = pi8  & ~n426;
  assign n428 = ~pi8  & n108;
  assign n429 = pi2  & n24;
  assign n430 = ~n428 & ~n429;
  assign n431 = pi5  & ~n430;
  assign n432 = ~n427 & ~n431;
  assign n433 = pi6  & ~n302;
  assign n434 = ~pi2  & pi9 ;
  assign n435 = ~n62 & ~n434;
  assign n436 = n433 & n435;
  assign n437 = n432 & ~n436;
  assign n438 = ~pi7  & ~n437;
  assign n439 = ~pi9  & n51;
  assign n440 = pi8  & ~n439;
  assign n441 = n84 & ~n440;
  assign n442 = ~n96 & ~n441;
  assign n443 = ~pi0  & ~n442;
  assign n444 = ~n156 & ~n307;
  assign n445 = pi7  & n444;
  assign n446 = ~pi2  & n445;
  assign n447 = ~n443 & ~n446;
  assign n448 = n332 & ~n447;
  assign n449 = ~n438 & ~n448;
  assign n450 = ~pi3  & ~n449;
  assign n451 = ~pi0  & ~pi6 ;
  assign n452 = n119 & ~n214;
  assign n453 = n451 & n452;
  assign n454 = ~pi8  & ~n29;
  assign n455 = ~n25 & ~n454;
  assign n456 = ~n24 & ~n96;
  assign n457 = ~n455 & n456;
  assign n458 = ~n453 & ~n457;
  assign n459 = ~pi5  & ~n458;
  assign n460 = ~pi8  & n219;
  assign n461 = pi0  & n172;
  assign n462 = ~n105 & ~n461;
  assign n463 = ~pi2  & ~n462;
  assign n464 = ~n460 & ~n463;
  assign n465 = pi9  & ~n464;
  assign n466 = ~pi0  & ~pi8 ;
  assign n467 = ~n205 & ~n466;
  assign n468 = n30 & n467;
  assign n469 = ~n465 & ~n468;
  assign n470 = ~n459 & n469;
  assign n471 = pi3  & ~n470;
  assign n472 = ~pi2  & pi5 ;
  assign n473 = n70 & n472;
  assign n474 = n24 & ~n182;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~pi8  & ~n475;
  assign n477 = pi2  & ~n128;
  assign n478 = ~n155 & ~n477;
  assign n479 = pi6  & ~n478;
  assign n480 = ~n476 & ~n479;
  assign n481 = pi1  & ~n480;
  assign n482 = ~pi9  & n275;
  assign n483 = n28 & ~n390;
  assign n484 = ~n482 & ~n483;
  assign n485 = ~pi2  & ~n484;
  assign n486 = pi2  & pi8 ;
  assign n487 = n24 & n486;
  assign n488 = ~n485 & ~n487;
  assign n489 = ~pi1  & ~n488;
  assign n490 = ~n481 & ~n489;
  assign n491 = ~n471 & n490;
  assign n492 = ~pi7  & ~n491;
  assign n493 = ~n450 & ~n492;
  assign n494 = ~pi4  & ~n493;
  assign n495 = ~n74 & ~n413;
  assign n496 = ~pi7  & ~n495;
  assign po6  = ~n494 & ~n496;
  assign n498 = ~pi3  & pi8 ;
  assign n499 = ~n75 & ~n498;
  assign n500 = pi0  & ~n499;
  assign n501 = ~pi3  & n154;
  assign n502 = pi0  & pi8 ;
  assign n503 = pi3  & ~n154;
  assign n504 = ~n502 & ~n503;
  assign n505 = ~pi6  & ~n504;
  assign n506 = ~n501 & ~n505;
  assign n507 = ~pi6  & ~n154;
  assign n508 = ~n433 & ~n507;
  assign n509 = n506 & n508;
  assign n510 = ~n500 & ~n509;
  assign n511 = ~pi2  & ~n510;
  assign n512 = pi2  & ~n506;
  assign n513 = ~pi3  & n129;
  assign n514 = ~n512 & ~n513;
  assign n515 = ~n511 & n514;
  assign n516 = pi1  & ~n515;
  assign n517 = ~pi0  & n433;
  assign n518 = n90 & n507;
  assign n519 = ~n517 & ~n518;
  assign n520 = pi3  & ~n519;
  assign n521 = ~pi0  & n195;
  assign n522 = ~n461 & ~n521;
  assign n523 = ~pi9  & ~n522;
  assign n524 = ~pi6  & ~n117;
  assign n525 = n477 & ~n524;
  assign n526 = ~n523 & ~n525;
  assign n527 = ~n520 & n526;
  assign n528 = ~pi1  & ~n527;
  assign n529 = n371 & n482;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~n516 & n530;
  assign n532 = ~pi5  & ~n531;
  assign n533 = pi0  & ~n435;
  assign n534 = pi5  & ~pi9 ;
  assign n535 = ~pi0  & n534;
  assign n536 = ~n533 & ~n535;
  assign n537 = pi8  & ~n536;
  assign n538 = n95 & n164;
  assign n539 = ~n537 & ~n538;
  assign n540 = ~pi3  & ~n539;
  assign n541 = pi3  & pi5 ;
  assign n542 = ~n62 & ~n541;
  assign n543 = ~pi0  & ~n542;
  assign n544 = pi3  & n472;
  assign n545 = ~n543 & ~n544;
  assign n546 = ~pi8  & ~n545;
  assign n547 = n371 & n534;
  assign n548 = ~n546 & ~n547;
  assign n549 = ~n540 & n548;
  assign n550 = pi1  & ~n549;
  assign n551 = ~pi2  & ~n42;
  assign n552 = ~n302 & ~n551;
  assign n553 = ~n110 & ~n552;
  assign n554 = pi5  & ~n553;
  assign n555 = pi2  & n128;
  assign n556 = n42 & n555;
  assign n557 = ~n554 & ~n556;
  assign n558 = ~pi1  & ~n557;
  assign n559 = pi8  & n392;
  assign n560 = n110 & n559;
  assign n561 = ~n558 & ~n560;
  assign n562 = ~n550 & n561;
  assign n563 = ~pi6  & ~n562;
  assign n564 = ~n532 & ~n563;
  assign n565 = ~pi7  & ~n564;
  assign n566 = ~n195 & ~n486;
  assign n567 = ~pi0  & ~n566;
  assign n568 = ~n204 & ~n567;
  assign n569 = ~pi9  & ~n568;
  assign n570 = n95 & n466;
  assign n571 = ~n569 & ~n570;
  assign n572 = ~pi2  & ~n51;
  assign n573 = ~n571 & ~n572;
  assign n574 = n218 & n573;
  assign n575 = n22 & n574;
  assign n576 = ~n565 & ~n575;
  assign n577 = ~pi4  & ~n576;
  assign n578 = pi4  & ~pi7 ;
  assign n579 = n22 & n578;
  assign n580 = n162 & n218;
  assign n581 = n579 & n580;
  assign po7  = ~n577 & ~n581;
  assign n583 = ~n108 & ~n256;
  assign n584 = ~n227 & ~n356;
  assign n585 = n583 & n584;
  assign n586 = ~pi2  & n585;
  assign n587 = n119 & ~n417;
  assign n588 = n103 & ~n587;
  assign n589 = ~n586 & ~n588;
  assign n590 = n26 & n158;
  assign n591 = ~n47 & n590;
  assign n592 = n589 & ~n591;
  assign n593 = ~pi8  & ~n592;
  assign n594 = ~n98 & n584;
  assign n595 = ~pi2  & n594;
  assign n596 = n141 & n205;
  assign n597 = ~n595 & ~n596;
  assign n598 = pi8  & ~n597;
  assign n599 = pi2  & ~n205;
  assign n600 = n265 & n599;
  assign n601 = ~n598 & ~n600;
  assign n602 = ~pi9  & ~n601;
  assign n603 = ~n181 & ~n541;
  assign n604 = ~n260 & ~n603;
  assign n605 = pi1  & n604;
  assign n606 = ~pi2  & ~n175;
  assign n607 = n271 & n606;
  assign n608 = ~n605 & ~n607;
  assign n609 = pi9  & ~n608;
  assign n610 = ~n602 & ~n609;
  assign n611 = ~n593 & n610;
  assign n612 = ~pi6  & ~n611;
  assign n613 = ~pi1  & ~n128;
  assign n614 = pi2  & ~n613;
  assign n615 = ~n282 & ~n614;
  assign n616 = pi0  & ~n615;
  assign n617 = ~n218 & n272;
  assign n618 = ~n284 & ~n617;
  assign n619 = ~n616 & n618;
  assign n620 = n356 & ~n619;
  assign n621 = ~n612 & ~n620;
  assign n622 = ~pi7  & ~n621;
  assign n623 = ~pi1  & ~n571;
  assign n624 = n118 & n521;
  assign n625 = ~n623 & ~n624;
  assign n626 = n22 & ~n625;
  assign n627 = ~pi6  & n626;
  assign n628 = ~n622 & ~n627;
  assign n629 = ~pi4  & ~n628;
  assign n630 = n77 & n579;
  assign po8  = ~n629 & ~n630;
  assign n632 = pi4  & ~n142;
  assign n633 = n205 & n383;
  assign n634 = ~pi7  & ~n633;
  assign n635 = ~n613 & ~n634;
  assign n636 = ~pi7  & ~n142;
  assign n637 = pi0  & ~n636;
  assign n638 = pi7  & ~n103;
  assign n639 = ~pi3  & ~n57;
  assign n640 = n217 & ~n499;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~pi2  & ~n641;
  assign n643 = ~n154 & n383;
  assign n644 = ~pi5  & n643;
  assign n645 = ~pi6  & ~n559;
  assign n646 = ~pi3  & ~n645;
  assign n647 = ~n644 & ~n646;
  assign n648 = ~n642 & n647;
  assign n649 = pi1  & ~n648;
  assign n650 = n217 & ~n393;
  assign n651 = ~n75 & ~n650;
  assign n652 = pi3  & ~n651;
  assign n653 = pi4  & ~n332;
  assign n654 = ~pi3  & ~n653;
  assign n655 = ~n652 & ~n654;
  assign n656 = ~pi2  & ~n655;
  assign n657 = n477 & n639;
  assign n658 = ~n264 & n657;
  assign n659 = ~n656 & ~n658;
  assign n660 = ~pi1  & ~n659;
  assign n661 = ~pi5  & ~n103;
  assign n662 = pi6  & ~n661;
  assign n663 = ~n660 & ~n662;
  assign n664 = ~n649 & n663;
  assign n665 = ~n638 & n664;
  assign n666 = ~n637 & n665;
  assign n667 = ~n635 & n666;
  assign po9  = ~n632 & n667;
  assign n669 = n406 & ~n455;
  assign n670 = pi2  & n669;
  assign n671 = ~n413 & ~n670;
  assign n672 = ~pi7  & ~n671;
  assign po10  = n332 & n672;
endmodule
