module mem_ctrl ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17,
    pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26,
    pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44,
    pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53,
    pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62,
    pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80,
    pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107,
    pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116,
    pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125,
    pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134,
    pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143,
    pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152,
    pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161,
    pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170,
    pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197,
    pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215,
    pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224,
    pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233,
    pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242,
    pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251,
    pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260,
    pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287,
    pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296,
    pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305,
    pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314,
    pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323,
    pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332,
    pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341,
    pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350,
    pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377,
    pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386,
    pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395,
    pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404,
    pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413,
    pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422,
    pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431,
    pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440,
    pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467,
    pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476,
    pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485,
    pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494,
    pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503,
    pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, pi512,
    pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520, pi521,
    pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529, pi530,
    pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539,
    pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548,
    pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557,
    pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566,
    pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574, pi575,
    pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583, pi584,
    pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592, pi593,
    pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601, pi602,
    pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610, pi611,
    pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619, pi620,
    pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629,
    pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638,
    pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647,
    pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656,
    pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664, pi665,
    pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673, pi674,
    pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682, pi683,
    pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691, pi692,
    pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700, pi701,
    pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709, pi710,
    pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719,
    pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728,
    pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737,
    pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746,
    pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754, pi755,
    pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763, pi764,
    pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772, pi773,
    pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781, pi782,
    pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790, pi791,
    pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799, pi800,
    pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808, pi809,
    pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818,
    pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827,
    pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835, pi836,
    pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844, pi845,
    pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853, pi854,
    pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862, pi863,
    pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871, pi872,
    pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880, pi881,
    pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889, pi890,
    pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898, pi899,
    pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907, pi908,
    pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916, pi917,
    pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925, pi926,
    pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934, pi935,
    pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943, pi944,
    pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952, pi953,
    pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961, pi962,
    pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970, pi971,
    pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979, pi980,
    pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988, pi989,
    pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997, pi998,
    pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0, po1, po2, po3, po4, po5, po6, po7, po8,
    po9, po10, po11, po12, po13, po14, po15, po16, po17,
    po18, po19, po20, po21, po22, po23, po24, po25, po26,
    po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44,
    po45, po46, po47, po48, po49, po50, po51, po52, po53,
    po54, po55, po56, po57, po58, po59, po60, po61, po62,
    po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80,
    po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98,
    po99, po100, po101, po102, po103, po104, po105, po106, po107,
    po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125,
    po126, po127, po128, po129, po130, po131, po132, po133, po134,
    po135, po136, po137, po138, po139, po140, po141, po142, po143,
    po144, po145, po146, po147, po148, po149, po150, po151, po152,
    po153, po154, po155, po156, po157, po158, po159, po160, po161,
    po162, po163, po164, po165, po166, po167, po168, po169, po170,
    po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188,
    po189, po190, po191, po192, po193, po194, po195, po196, po197,
    po198, po199, po200, po201, po202, po203, po204, po205, po206,
    po207, po208, po209, po210, po211, po212, po213, po214, po215,
    po216, po217, po218, po219, po220, po221, po222, po223, po224,
    po225, po226, po227, po228, po229, po230, po231, po232, po233,
    po234, po235, po236, po237, po238, po239, po240, po241, po242,
    po243, po244, po245, po246, po247, po248, po249, po250, po251,
    po252, po253, po254, po255, po256, po257, po258, po259, po260,
    po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278,
    po279, po280, po281, po282, po283, po284, po285, po286, po287,
    po288, po289, po290, po291, po292, po293, po294, po295, po296,
    po297, po298, po299, po300, po301, po302, po303, po304, po305,
    po306, po307, po308, po309, po310, po311, po312, po313, po314,
    po315, po316, po317, po318, po319, po320, po321, po322, po323,
    po324, po325, po326, po327, po328, po329, po330, po331, po332,
    po333, po334, po335, po336, po337, po338, po339, po340, po341,
    po342, po343, po344, po345, po346, po347, po348, po349, po350,
    po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368,
    po369, po370, po371, po372, po373, po374, po375, po376, po377,
    po378, po379, po380, po381, po382, po383, po384, po385, po386,
    po387, po388, po389, po390, po391, po392, po393, po394, po395,
    po396, po397, po398, po399, po400, po401, po402, po403, po404,
    po405, po406, po407, po408, po409, po410, po411, po412, po413,
    po414, po415, po416, po417, po418, po419, po420, po421, po422,
    po423, po424, po425, po426, po427, po428, po429, po430, po431,
    po432, po433, po434, po435, po436, po437, po438, po439, po440,
    po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458,
    po459, po460, po461, po462, po463, po464, po465, po466, po467,
    po468, po469, po470, po471, po472, po473, po474, po475, po476,
    po477, po478, po479, po480, po481, po482, po483, po484, po485,
    po486, po487, po488, po489, po490, po491, po492, po493, po494,
    po495, po496, po497, po498, po499, po500, po501, po502, po503,
    po504, po505, po506, po507, po508, po509, po510, po511, po512,
    po513, po514, po515, po516, po517, po518, po519, po520, po521,
    po522, po523, po524, po525, po526, po527, po528, po529, po530,
    po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548,
    po549, po550, po551, po552, po553, po554, po555, po556, po557,
    po558, po559, po560, po561, po562, po563, po564, po565, po566,
    po567, po568, po569, po570, po571, po572, po573, po574, po575,
    po576, po577, po578, po579, po580, po581, po582, po583, po584,
    po585, po586, po587, po588, po589, po590, po591, po592, po593,
    po594, po595, po596, po597, po598, po599, po600, po601, po602,
    po603, po604, po605, po606, po607, po608, po609, po610, po611,
    po612, po613, po614, po615, po616, po617, po618, po619, po620,
    po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638,
    po639, po640, po641, po642, po643, po644, po645, po646, po647,
    po648, po649, po650, po651, po652, po653, po654, po655, po656,
    po657, po658, po659, po660, po661, po662, po663, po664, po665,
    po666, po667, po668, po669, po670, po671, po672, po673, po674,
    po675, po676, po677, po678, po679, po680, po681, po682, po683,
    po684, po685, po686, po687, po688, po689, po690, po691, po692,
    po693, po694, po695, po696, po697, po698, po699, po700, po701,
    po702, po703, po704, po705, po706, po707, po708, po709, po710,
    po711, po712, po713, po714, po715, po716, po717, po718, po719,
    po720, po721, po722, po723, po724, po725, po726, po727, po728,
    po729, po730, po731, po732, po733, po734, po735, po736, po737,
    po738, po739, po740, po741, po742, po743, po744, po745, po746,
    po747, po748, po749, po750, po751, po752, po753, po754, po755,
    po756, po757, po758, po759, po760, po761, po762, po763, po764,
    po765, po766, po767, po768, po769, po770, po771, po772, po773,
    po774, po775, po776, po777, po778, po779, po780, po781, po782,
    po783, po784, po785, po786, po787, po788, po789, po790, po791,
    po792, po793, po794, po795, po796, po797, po798, po799, po800,
    po801, po802, po803, po804, po805, po806, po807, po808, po809,
    po810, po811, po812, po813, po814, po815, po816, po817, po818,
    po819, po820, po821, po822, po823, po824, po825, po826, po827,
    po828, po829, po830, po831, po832, po833, po834, po835, po836,
    po837, po838, po839, po840, po841, po842, po843, po844, po845,
    po846, po847, po848, po849, po850, po851, po852, po853, po854,
    po855, po856, po857, po858, po859, po860, po861, po862, po863,
    po864, po865, po866, po867, po868, po869, po870, po871, po872,
    po873, po874, po875, po876, po877, po878, po879, po880, po881,
    po882, po883, po884, po885, po886, po887, po888, po889, po890,
    po891, po892, po893, po894, po895, po896, po897, po898, po899,
    po900, po901, po902, po903, po904, po905, po906, po907, po908,
    po909, po910, po911, po912, po913, po914, po915, po916, po917,
    po918, po919, po920, po921, po922, po923, po924, po925, po926,
    po927, po928, po929, po930, po931, po932, po933, po934, po935,
    po936, po937, po938, po939, po940, po941, po942, po943, po944,
    po945, po946, po947, po948, po949, po950, po951, po952, po953,
    po954, po955, po956, po957, po958, po959, po960, po961, po962,
    po963, po964, po965, po966, po967, po968, po969, po970, po971,
    po972, po973, po974, po975, po976, po977, po978, po979, po980,
    po981, po982, po983, po984, po985, po986, po987, po988, po989,
    po990, po991, po992, po993, po994, po995, po996, po997, po998,
    po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7,
    pi8, pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16,
    pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25,
    pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34,
    pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43,
    pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52,
    pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61,
    pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70,
    pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97,
    pi98, pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106,
    pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115,
    pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124,
    pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133,
    pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142,
    pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151,
    pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160,
    pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187,
    pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196,
    pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205,
    pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214,
    pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223,
    pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232,
    pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241,
    pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250,
    pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277,
    pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286,
    pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295,
    pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304,
    pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313,
    pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322,
    pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331,
    pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340,
    pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367,
    pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376,
    pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385,
    pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394,
    pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403,
    pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412,
    pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421,
    pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430,
    pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457,
    pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466,
    pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475,
    pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484,
    pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493,
    pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502,
    pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511,
    pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520,
    pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529,
    pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538,
    pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547,
    pi548, pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556,
    pi557, pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565,
    pi566, pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574,
    pi575, pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583,
    pi584, pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592,
    pi593, pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601,
    pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610,
    pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619,
    pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628,
    pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637,
    pi638, pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646,
    pi647, pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655,
    pi656, pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664,
    pi665, pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673,
    pi674, pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682,
    pi683, pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691,
    pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700,
    pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709,
    pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718,
    pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727,
    pi728, pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736,
    pi737, pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745,
    pi746, pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754,
    pi755, pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763,
    pi764, pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772,
    pi773, pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781,
    pi782, pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790,
    pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799,
    pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808,
    pi809, pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817,
    pi818, pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826,
    pi827, pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835,
    pi836, pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844,
    pi845, pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853,
    pi854, pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862,
    pi863, pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871,
    pi872, pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880,
    pi881, pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889,
    pi890, pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898,
    pi899, pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907,
    pi908, pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916,
    pi917, pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925,
    pi926, pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934,
    pi935, pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943,
    pi944, pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952,
    pi953, pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961,
    pi962, pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970,
    pi971, pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979,
    pi980, pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988,
    pi989, pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997,
    pi998, pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0, po1, po2, po3, po4, po5, po6, po7,
    po8, po9, po10, po11, po12, po13, po14, po15, po16,
    po17, po18, po19, po20, po21, po22, po23, po24, po25,
    po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43,
    po44, po45, po46, po47, po48, po49, po50, po51, po52,
    po53, po54, po55, po56, po57, po58, po59, po60, po61,
    po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88,
    po89, po90, po91, po92, po93, po94, po95, po96, po97,
    po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115,
    po116, po117, po118, po119, po120, po121, po122, po123, po124,
    po125, po126, po127, po128, po129, po130, po131, po132, po133,
    po134, po135, po136, po137, po138, po139, po140, po141, po142,
    po143, po144, po145, po146, po147, po148, po149, po150, po151,
    po152, po153, po154, po155, po156, po157, po158, po159, po160,
    po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178,
    po179, po180, po181, po182, po183, po184, po185, po186, po187,
    po188, po189, po190, po191, po192, po193, po194, po195, po196,
    po197, po198, po199, po200, po201, po202, po203, po204, po205,
    po206, po207, po208, po209, po210, po211, po212, po213, po214,
    po215, po216, po217, po218, po219, po220, po221, po222, po223,
    po224, po225, po226, po227, po228, po229, po230, po231, po232,
    po233, po234, po235, po236, po237, po238, po239, po240, po241,
    po242, po243, po244, po245, po246, po247, po248, po249, po250,
    po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268,
    po269, po270, po271, po272, po273, po274, po275, po276, po277,
    po278, po279, po280, po281, po282, po283, po284, po285, po286,
    po287, po288, po289, po290, po291, po292, po293, po294, po295,
    po296, po297, po298, po299, po300, po301, po302, po303, po304,
    po305, po306, po307, po308, po309, po310, po311, po312, po313,
    po314, po315, po316, po317, po318, po319, po320, po321, po322,
    po323, po324, po325, po326, po327, po328, po329, po330, po331,
    po332, po333, po334, po335, po336, po337, po338, po339, po340,
    po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358,
    po359, po360, po361, po362, po363, po364, po365, po366, po367,
    po368, po369, po370, po371, po372, po373, po374, po375, po376,
    po377, po378, po379, po380, po381, po382, po383, po384, po385,
    po386, po387, po388, po389, po390, po391, po392, po393, po394,
    po395, po396, po397, po398, po399, po400, po401, po402, po403,
    po404, po405, po406, po407, po408, po409, po410, po411, po412,
    po413, po414, po415, po416, po417, po418, po419, po420, po421,
    po422, po423, po424, po425, po426, po427, po428, po429, po430,
    po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448,
    po449, po450, po451, po452, po453, po454, po455, po456, po457,
    po458, po459, po460, po461, po462, po463, po464, po465, po466,
    po467, po468, po469, po470, po471, po472, po473, po474, po475,
    po476, po477, po478, po479, po480, po481, po482, po483, po484,
    po485, po486, po487, po488, po489, po490, po491, po492, po493,
    po494, po495, po496, po497, po498, po499, po500, po501, po502,
    po503, po504, po505, po506, po507, po508, po509, po510, po511,
    po512, po513, po514, po515, po516, po517, po518, po519, po520,
    po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538,
    po539, po540, po541, po542, po543, po544, po545, po546, po547,
    po548, po549, po550, po551, po552, po553, po554, po555, po556,
    po557, po558, po559, po560, po561, po562, po563, po564, po565,
    po566, po567, po568, po569, po570, po571, po572, po573, po574,
    po575, po576, po577, po578, po579, po580, po581, po582, po583,
    po584, po585, po586, po587, po588, po589, po590, po591, po592,
    po593, po594, po595, po596, po597, po598, po599, po600, po601,
    po602, po603, po604, po605, po606, po607, po608, po609, po610,
    po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628,
    po629, po630, po631, po632, po633, po634, po635, po636, po637,
    po638, po639, po640, po641, po642, po643, po644, po645, po646,
    po647, po648, po649, po650, po651, po652, po653, po654, po655,
    po656, po657, po658, po659, po660, po661, po662, po663, po664,
    po665, po666, po667, po668, po669, po670, po671, po672, po673,
    po674, po675, po676, po677, po678, po679, po680, po681, po682,
    po683, po684, po685, po686, po687, po688, po689, po690, po691,
    po692, po693, po694, po695, po696, po697, po698, po699, po700,
    po701, po702, po703, po704, po705, po706, po707, po708, po709,
    po710, po711, po712, po713, po714, po715, po716, po717, po718,
    po719, po720, po721, po722, po723, po724, po725, po726, po727,
    po728, po729, po730, po731, po732, po733, po734, po735, po736,
    po737, po738, po739, po740, po741, po742, po743, po744, po745,
    po746, po747, po748, po749, po750, po751, po752, po753, po754,
    po755, po756, po757, po758, po759, po760, po761, po762, po763,
    po764, po765, po766, po767, po768, po769, po770, po771, po772,
    po773, po774, po775, po776, po777, po778, po779, po780, po781,
    po782, po783, po784, po785, po786, po787, po788, po789, po790,
    po791, po792, po793, po794, po795, po796, po797, po798, po799,
    po800, po801, po802, po803, po804, po805, po806, po807, po808,
    po809, po810, po811, po812, po813, po814, po815, po816, po817,
    po818, po819, po820, po821, po822, po823, po824, po825, po826,
    po827, po828, po829, po830, po831, po832, po833, po834, po835,
    po836, po837, po838, po839, po840, po841, po842, po843, po844,
    po845, po846, po847, po848, po849, po850, po851, po852, po853,
    po854, po855, po856, po857, po858, po859, po860, po861, po862,
    po863, po864, po865, po866, po867, po868, po869, po870, po871,
    po872, po873, po874, po875, po876, po877, po878, po879, po880,
    po881, po882, po883, po884, po885, po886, po887, po888, po889,
    po890, po891, po892, po893, po894, po895, po896, po897, po898,
    po899, po900, po901, po902, po903, po904, po905, po906, po907,
    po908, po909, po910, po911, po912, po913, po914, po915, po916,
    po917, po918, po919, po920, po921, po922, po923, po924, po925,
    po926, po927, po928, po929, po930, po931, po932, po933, po934,
    po935, po936, po937, po938, po939, po940, po941, po942, po943,
    po944, po945, po946, po947, po948, po949, po950, po951, po952,
    po953, po954, po955, po956, po957, po958, po959, po960, po961,
    po962, po963, po964, po965, po966, po967, po968, po969, po970,
    po971, po972, po973, po974, po975, po976, po977, po978, po979,
    po980, po981, po982, po983, po984, po985, po986, po987, po988,
    po989, po990, po991, po992, po993, po994, po995, po996, po997,
    po998, po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2799, n2800, n2801, n2802, n2803,
    n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821,
    n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851,
    n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2880, n2881,
    n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911,
    n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953,
    n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001,
    n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061,
    n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085,
    n3086, n3087, n3088, n3089, n3090, n3091,
    n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151,
    n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175,
    n3176, n3177, n3178, n3179, n3180, n3181,
    n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211,
    n3212, n3213, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241,
    n3242, n3243, n3244, n3245, n3246, n3247,
    n3248, n3249, n3250, n3251, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271,
    n3272, n3273, n3274, n3275, n3276, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541,
    n3542, n3543, n3544, n3545, n3546, n3547,
    n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565,
    n3566, n3567, n3568, n3569, n3570, n3571,
    n3572, n3573, n3574, n3575, n3576, n3577,
    n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601,
    n3602, n3603, n3604, n3605, n3606, n3607,
    n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631,
    n3632, n3633, n3634, n3635, n3636, n3637,
    n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661,
    n3662, n3663, n3664, n3665, n3666, n3667,
    n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691,
    n3692, n3693, n3694, n3695, n3696, n3697,
    n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721,
    n3722, n3723, n3724, n3725, n3726, n3727,
    n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751,
    n3752, n3753, n3754, n3755, n3756, n3757,
    n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775,
    n3776, n3777, n3778, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787,
    n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805,
    n3806, n3807, n3808, n3809, n3810, n3811,
    n3812, n3813, n3814, n3815, n3816, n3817,
    n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835,
    n3836, n3837, n3838, n3839, n3840, n3841,
    n3842, n3843, n3844, n3845, n3846, n3847,
    n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877,
    n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901,
    n3902, n3903, n3904, n3905, n3906, n3907,
    n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931,
    n3932, n3933, n3934, n3935, n3936, n3937,
    n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961,
    n3962, n3963, n3964, n3965, n3966, n3967,
    n3968, n3969, n3970, n3971, n3972, n3973,
    n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3991,
    n3992, n3993, n3994, n3995, n3996, n3997,
    n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057,
    n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117,
    n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141,
    n4142, n4143, n4144, n4145, n4146, n4147,
    n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171,
    n4172, n4173, n4174, n4175, n4176, n4177,
    n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195,
    n4196, n4197, n4198, n4199, n4200, n4201,
    n4202, n4203, n4204, n4205, n4206, n4207,
    n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219,
    n4220, n4221, n4222, n4223, n4224, n4225,
    n4226, n4227, n4228, n4229, n4230, n4231,
    n4232, n4233, n4234, n4235, n4236, n4237,
    n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249,
    n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4259, n4260, n4261,
    n4262, n4263, n4264, n4265, n4266, n4267,
    n4268, n4269, n4270, n4271, n4272, n4273,
    n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291,
    n4292, n4293, n4294, n4295, n4296, n4297,
    n4298, n4299, n4300, n4301, n4302, n4303,
    n4304, n4305, n4306, n4307, n4308, n4309,
    n4310, n4311, n4312, n4313, n4314, n4315,
    n4316, n4317, n4318, n4319, n4320, n4321,
    n4322, n4323, n4324, n4325, n4326, n4327,
    n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339,
    n4340, n4341, n4342, n4343, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351,
    n4352, n4353, n4354, n4355, n4356, n4357,
    n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369,
    n4370, n4371, n4372, n4373, n4374, n4375,
    n4376, n4377, n4378, n4379, n4380, n4381,
    n4382, n4383, n4384, n4385, n4386, n4387,
    n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399,
    n4400, n4401, n4402, n4403, n4404, n4405,
    n4406, n4407, n4408, n4409, n4410, n4411,
    n4412, n4413, n4414, n4415, n4416, n4417,
    n4418, n4419, n4420, n4421, n4422, n4423,
    n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435,
    n4436, n4437, n4438, n4439, n4440, n4441,
    n4442, n4443, n4444, n4445, n4446, n4447,
    n4448, n4449, n4450, n4451, n4452, n4453,
    n4454, n4455, n4456, n4457, n4458, n4459,
    n4460, n4461, n4462, n4463, n4464, n4465,
    n4466, n4467, n4468, n4469, n4470, n4471,
    n4472, n4473, n4474, n4475, n4476, n4477,
    n4478, n4479, n4480, n4481, n4482, n4483,
    n4484, n4485, n4486, n4487, n4488, n4489,
    n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501,
    n4502, n4503, n4504, n4505, n4506, n4507,
    n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531,
    n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843,
    n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861,
    n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873,
    n4874, n4875, n4876, n4877, n4878, n4879,
    n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891,
    n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137,
    n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161,
    n5162, n5163, n5164, n5165, n5166, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191,
    n5192, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209,
    n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221,
    n5222, n5223, n5224, n5225, n5226, n5227,
    n5228, n5229, n5230, n5231, n5232, n5233,
    n5234, n5235, n5236, n5237, n5238, n5239,
    n5240, n5241, n5242, n5243, n5244, n5245,
    n5246, n5247, n5248, n5249, n5250, n5251,
    n5252, n5253, n5254, n5255, n5256, n5257,
    n5258, n5259, n5260, n5261, n5262, n5263,
    n5264, n5265, n5266, n5267, n5268, n5269,
    n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281,
    n5282, n5283, n5284, n5285, n5286, n5287,
    n5288, n5289, n5290, n5291, n5292, n5293,
    n5294, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5308, n5309, n5310, n5311,
    n5312, n5313, n5314, n5315, n5316, n5317,
    n5318, n5319, n5320, n5321, n5322, n5323,
    n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335,
    n5336, n5337, n5338, n5339, n5340, n5341,
    n5342, n5343, n5344, n5345, n5346, n5347,
    n5348, n5349, n5350, n5351, n5352, n5353,
    n5354, n5355, n5356, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371,
    n5372, n5373, n5374, n5375, n5376, n5377,
    n5378, n5379, n5380, n5381, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389,
    n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401,
    n5402, n5403, n5404, n5405, n5406, n5407,
    n5408, n5409, n5410, n5411, n5412, n5413,
    n5414, n5415, n5416, n5417, n5418, n5419,
    n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431,
    n5432, n5433, n5434, n5435, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443,
    n5444, n5445, n5446, n5447, n5448, n5449,
    n5450, n5451, n5452, n5453, n5454, n5455,
    n5456, n5457, n5458, n5459, n5460, n5461,
    n5462, n5463, n5464, n5465, n5466, n5467,
    n5468, n5469, n5470, n5471, n5472, n5473,
    n5474, n5475, n5476, n5477, n5478, n5479,
    n5480, n5481, n5482, n5483, n5484, n5485,
    n5486, n5487, n5488, n5489, n5490, n5491,
    n5492, n5493, n5494, n5495, n5496, n5497,
    n5498, n5499, n5500, n5501, n5502, n5503,
    n5504, n5505, n5506, n5507, n5508, n5509,
    n5510, n5511, n5512, n5513, n5514, n5515,
    n5516, n5517, n5518, n5519, n5520, n5521,
    n5522, n5523, n5524, n5525, n5526, n5527,
    n5528, n5529, n5530, n5531, n5532, n5533,
    n5534, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551,
    n5552, n5553, n5554, n5555, n5556, n5557,
    n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581,
    n5582, n5583, n5584, n5585, n5586, n5587,
    n5588, n5589, n5590, n5591, n5592, n5593,
    n5594, n5595, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611,
    n5612, n5613, n5614, n5615, n5616, n5617,
    n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5625, n5626, n5627, n5628, n5629,
    n5630, n5631, n5632, n5633, n5634, n5635,
    n5636, n5637, n5638, n5639, n5640, n5641,
    n5642, n5643, n5644, n5645, n5646, n5647,
    n5648, n5649, n5650, n5651, n5652, n5653,
    n5654, n5655, n5656, n5657, n5658, n5659,
    n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5670, n5671,
    n5672, n5673, n5674, n5675, n5676, n5677,
    n5678, n5679, n5680, n5681, n5682, n5683,
    n5684, n5685, n5686, n5687, n5688, n5689,
    n5690, n5691, n5692, n5693, n5694, n5695,
    n5696, n5697, n5698, n5699, n5700, n5701,
    n5702, n5703, n5704, n5705, n5706, n5707,
    n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5716, n5717, n5718, n5719,
    n5720, n5721, n5722, n5723, n5724, n5725,
    n5726, n5727, n5728, n5729, n5730, n5731,
    n5732, n5733, n5734, n5735, n5736, n5737,
    n5738, n5739, n5740, n5741, n5742, n5743,
    n5744, n5745, n5746, n5747, n5748, n5749,
    n5750, n5751, n5752, n5753, n5754, n5755,
    n5756, n5757, n5758, n5759, n5760, n5761,
    n5762, n5763, n5764, n5765, n5766, n5767,
    n5768, n5769, n5770, n5771, n5772, n5773,
    n5774, n5775, n5776, n5777, n5778, n5779,
    n5780, n5781, n5782, n5783, n5784, n5785,
    n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797,
    n5798, n5799, n5800, n5801, n5802, n5803,
    n5804, n5805, n5806, n5807, n5808, n5809,
    n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5817, n5818, n5819, n5820, n5821,
    n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839,
    n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857,
    n5858, n5859, n5860, n5861, n5862, n5863,
    n5864, n5865, n5866, n5867, n5868, n5869,
    n5870, n5871, n5872, n5873, n5874, n5875,
    n5876, n5877, n5878, n5879, n5880, n5881,
    n5882, n5883, n5884, n5885, n5886, n5887,
    n5888, n5889, n5890, n5891, n5892, n5893,
    n5894, n5895, n5896, n5897, n5898, n5899,
    n5900, n5901, n5902, n5903, n5904, n5905,
    n5906, n5907, n5908, n5909, n5910, n5911,
    n5912, n5913, n5914, n5915, n5916, n5917,
    n5918, n5919, n5920, n5921, n5922, n5923,
    n5924, n5925, n5926, n5927, n5928, n5929,
    n5930, n5931, n5932, n5933, n5934, n5935,
    n5936, n5937, n5938, n5939, n5940, n5941,
    n5942, n5943, n5944, n5945, n5946, n5947,
    n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5958, n5959,
    n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977,
    n5978, n5979, n5980, n5981, n5982, n5983,
    n5984, n5985, n5986, n5987, n5988, n5989,
    n5990, n5991, n5992, n5993, n5994, n5995,
    n5996, n5997, n5998, n5999, n6000, n6001,
    n6002, n6003, n6004, n6005, n6006, n6007,
    n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019,
    n6020, n6021, n6022, n6023, n6024, n6025,
    n6026, n6027, n6028, n6029, n6030, n6031,
    n6032, n6033, n6034, n6035, n6036, n6037,
    n6038, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049,
    n6050, n6051, n6052, n6053, n6054, n6055,
    n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067,
    n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079,
    n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097,
    n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151,
    n6152, n6153, n6154, n6155, n6156, n6157,
    n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175,
    n6176, n6177, n6178, n6179, n6180, n6181,
    n6182, n6183, n6184, n6185, n6186, n6187,
    n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6203, n6204, n6205,
    n6206, n6207, n6208, n6209, n6210, n6211,
    n6212, n6213, n6214, n6215, n6216, n6217,
    n6218, n6219, n6220, n6221, n6222, n6223,
    n6224, n6225, n6226, n6227, n6228, n6229,
    n6230, n6231, n6232, n6233, n6234, n6235,
    n6236, n6237, n6238, n6239, n6240, n6241,
    n6242, n6243, n6244, n6245, n6246, n6247,
    n6248, n6249, n6250, n6251, n6252, n6253,
    n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271,
    n6272, n6273, n6274, n6275, n6276, n6277,
    n6278, n6279, n6280, n6281, n6282, n6283,
    n6284, n6285, n6286, n6287, n6288, n6289,
    n6290, n6291, n6292, n6293, n6294, n6295,
    n6296, n6297, n6298, n6299, n6300, n6301,
    n6302, n6303, n6304, n6305, n6306, n6307,
    n6308, n6309, n6310, n6311, n6312, n6313,
    n6314, n6315, n6316, n6317, n6318, n6319,
    n6320, n6321, n6322, n6323, n6324, n6325,
    n6326, n6327, n6328, n6329, n6330, n6331,
    n6332, n6333, n6334, n6335, n6336, n6337,
    n6338, n6339, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349,
    n6350, n6351, n6352, n6353, n6354, n6355,
    n6356, n6357, n6358, n6359, n6360, n6361,
    n6362, n6363, n6364, n6365, n6366, n6367,
    n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379,
    n6380, n6381, n6382, n6383, n6384, n6385,
    n6386, n6387, n6388, n6389, n6390, n6391,
    n6392, n6393, n6394, n6395, n6396, n6397,
    n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409,
    n6410, n6411, n6412, n6413, n6414, n6415,
    n6416, n6417, n6418, n6419, n6420, n6421,
    n6422, n6423, n6424, n6425, n6426, n6427,
    n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6437, n6438, n6439,
    n6440, n6441, n6442, n6443, n6444, n6445,
    n6446, n6447, n6448, n6449, n6450, n6451,
    n6452, n6453, n6454, n6455, n6456, n6457,
    n6458, n6459, n6460, n6461, n6462, n6463,
    n6464, n6465, n6466, n6467, n6468, n6469,
    n6470, n6471, n6472, n6473, n6474, n6475,
    n6476, n6477, n6478, n6479, n6480, n6481,
    n6482, n6483, n6484, n6485, n6486, n6487,
    n6488, n6489, n6490, n6491, n6492, n6493,
    n6494, n6495, n6496, n6497, n6498, n6499,
    n6500, n6501, n6502, n6503, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511,
    n6512, n6513, n6514, n6515, n6516, n6517,
    n6518, n6519, n6520, n6521, n6522, n6523,
    n6524, n6525, n6526, n6527, n6528, n6529,
    n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541,
    n6542, n6543, n6544, n6545, n6546, n6547,
    n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571,
    n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601,
    n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649,
    n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661,
    n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691,
    n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721,
    n6722, n6723, n6724, n6725, n6726, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751,
    n6752, n6753, n6754, n6755, n6756, n6757,
    n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781,
    n6782, n6783, n6784, n6785, n6786, n6787,
    n6788, n6789, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6899, n6900, n6901, n6902, n6903,
    n6904, n6905, n6906, n6907, n6908, n6909,
    n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921,
    n6922, n6923, n6924, n6925, n6926, n6927,
    n6928, n6929, n6930, n6931, n6932, n6933,
    n6934, n6935, n6936, n6937, n6938, n6939,
    n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951,
    n6952, n6953, n6954, n6955, n6956, n6957,
    n6958, n6959, n6960, n6961, n6962, n6963,
    n6964, n6965, n6966, n6967, n6968, n6969,
    n6970, n6971, n6972, n6973, n6974, n6975,
    n6976, n6977, n6978, n6979, n6980, n6981,
    n6982, n6983, n6984, n6985, n6986, n6987,
    n6988, n6989, n6990, n6991, n6992, n6993,
    n6994, n6995, n6996, n6997, n6998, n6999,
    n7000, n7001, n7002, n7003, n7004, n7005,
    n7006, n7007, n7008, n7009, n7010, n7011,
    n7012, n7013, n7014, n7015, n7016, n7017,
    n7018, n7019, n7020, n7021, n7022, n7023,
    n7024, n7025, n7026, n7027, n7028, n7029,
    n7030, n7031, n7032, n7033, n7034, n7035,
    n7036, n7037, n7038, n7039, n7040, n7041,
    n7042, n7043, n7044, n7045, n7046, n7047,
    n7048, n7049, n7050, n7051, n7052, n7053,
    n7054, n7055, n7056, n7057, n7058, n7059,
    n7060, n7061, n7062, n7063, n7064, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071,
    n7072, n7073, n7074, n7075, n7076, n7077,
    n7078, n7079, n7080, n7081, n7082, n7083,
    n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101,
    n7102, n7103, n7104, n7105, n7106, n7107,
    n7108, n7109, n7110, n7111, n7112, n7113,
    n7114, n7115, n7116, n7117, n7118, n7119,
    n7120, n7121, n7122, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131,
    n7132, n7133, n7134, n7135, n7136, n7137,
    n7138, n7139, n7140, n7141, n7142, n7143,
    n7144, n7145, n7146, n7147, n7148, n7149,
    n7150, n7151, n7152, n7153, n7154, n7155,
    n7156, n7157, n7158, n7159, n7160, n7161,
    n7162, n7163, n7164, n7165, n7166, n7167,
    n7168, n7169, n7170, n7171, n7172, n7173,
    n7174, n7175, n7176, n7177, n7178, n7179,
    n7180, n7181, n7182, n7183, n7184, n7185,
    n7186, n7187, n7188, n7189, n7190, n7191,
    n7192, n7193, n7194, n7195, n7196, n7197,
    n7198, n7199, n7200, n7201, n7202, n7203,
    n7204, n7205, n7206, n7207, n7208, n7209,
    n7210, n7211, n7212, n7213, n7214, n7215,
    n7216, n7217, n7218, n7219, n7220, n7221,
    n7222, n7223, n7224, n7225, n7226, n7227,
    n7228, n7229, n7230, n7231, n7232, n7233,
    n7234, n7235, n7236, n7237, n7238, n7239,
    n7240, n7241, n7242, n7243, n7244, n7245,
    n7246, n7247, n7248, n7249, n7250, n7251,
    n7252, n7253, n7254, n7255, n7256, n7257,
    n7258, n7259, n7260, n7261, n7262, n7263,
    n7264, n7265, n7266, n7267, n7268, n7269,
    n7270, n7271, n7272, n7273, n7274, n7275,
    n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287,
    n7288, n7289, n7290, n7291, n7292, n7293,
    n7294, n7295, n7296, n7297, n7298, n7299,
    n7300, n7301, n7302, n7303, n7304, n7305,
    n7306, n7307, n7308, n7309, n7310, n7311,
    n7312, n7313, n7314, n7315, n7316, n7317,
    n7318, n7319, n7320, n7321, n7322, n7323,
    n7324, n7325, n7326, n7327, n7328, n7329,
    n7330, n7331, n7332, n7333, n7334, n7335,
    n7336, n7337, n7338, n7339, n7340, n7341,
    n7342, n7343, n7344, n7345, n7346, n7347,
    n7348, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359,
    n7360, n7361, n7362, n7363, n7364, n7365,
    n7366, n7367, n7368, n7369, n7370, n7371,
    n7372, n7373, n7374, n7375, n7376, n7377,
    n7378, n7379, n7380, n7381, n7382, n7383,
    n7384, n7385, n7386, n7387, n7388, n7389,
    n7390, n7391, n7392, n7393, n7394, n7395,
    n7396, n7397, n7398, n7399, n7400, n7401,
    n7402, n7403, n7404, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431,
    n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443,
    n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461,
    n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479,
    n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491,
    n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503,
    n7504, n7505, n7506, n7507, n7508, n7509,
    n7510, n7511, n7512, n7513, n7514, n7515,
    n7516, n7517, n7518, n7519, n7520, n7521,
    n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551,
    n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581,
    n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725,
    n7726, n7727, n7728, n7729, n7730, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737,
    n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7746, n7747, n7748, n7749,
    n7750, n7751, n7752, n7753, n7754, n7755,
    n7756, n7757, n7758, n7759, n7760, n7761,
    n7762, n7763, n7764, n7765, n7766, n7767,
    n7768, n7769, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785,
    n7786, n7787, n7788, n7789, n7790, n7791,
    n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821,
    n7822, n7823, n7824, n7825, n7826, n7827,
    n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851,
    n7852, n7853, n7854, n7855, n7856, n7857,
    n7858, n7859, n7860, n7861, n7862, n7863,
    n7864, n7865, n7866, n7867, n7868, n7869,
    n7870, n7871, n7872, n7873, n7874, n7875,
    n7876, n7877, n7878, n7879, n7880, n7881,
    n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893,
    n7894, n7895, n7896, n7897, n7898, n7899,
    n7900, n7901, n7902, n7903, n7904, n7905,
    n7906, n7907, n7908, n7909, n7910, n7911,
    n7912, n7913, n7914, n7915, n7916, n7917,
    n7918, n7919, n7920, n7921, n7922, n7923,
    n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935,
    n7936, n7937, n7938, n7939, n7940, n7941,
    n7942, n7943, n7944, n7945, n7946, n7947,
    n7948, n7949, n7950, n7951, n7952, n7953,
    n7954, n7955, n7956, n7957, n7958, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965,
    n7966, n7967, n7968, n7969, n7970, n7971,
    n7972, n7973, n7974, n7975, n7976, n7977,
    n7978, n7979, n7980, n7981, n7982, n7983,
    n7984, n7985, n7986, n7987, n7988, n7989,
    n7990, n7991, n7992, n7993, n7994, n7995,
    n7996, n7997, n7998, n7999, n8000, n8001,
    n8002, n8003, n8004, n8005, n8006, n8007,
    n8008, n8009, n8010, n8011, n8012, n8013,
    n8014, n8015, n8016, n8017, n8018, n8019,
    n8020, n8021, n8022, n8023, n8024, n8025,
    n8026, n8027, n8028, n8029, n8030, n8031,
    n8032, n8033, n8034, n8035, n8036, n8037,
    n8038, n8039, n8040, n8041, n8042, n8043,
    n8044, n8045, n8046, n8047, n8048, n8049,
    n8050, n8051, n8052, n8053, n8054, n8055,
    n8056, n8057, n8058, n8059, n8060, n8061,
    n8062, n8063, n8064, n8065, n8066, n8067,
    n8068, n8069, n8070, n8071, n8072, n8073,
    n8074, n8075, n8076, n8077, n8078, n8079,
    n8080, n8081, n8082, n8083, n8084, n8085,
    n8086, n8087, n8088, n8089, n8090, n8091,
    n8092, n8093, n8094, n8095, n8096, n8097,
    n8098, n8099, n8100, n8101, n8102, n8103,
    n8104, n8105, n8106, n8107, n8108, n8109,
    n8110, n8111, n8112, n8113, n8114, n8115,
    n8116, n8117, n8118, n8119, n8120, n8121,
    n8122, n8123, n8124, n8125, n8126, n8127,
    n8128, n8129, n8130, n8131, n8132, n8133,
    n8134, n8135, n8136, n8137, n8138, n8139,
    n8140, n8141, n8142, n8143, n8144, n8145,
    n8146, n8147, n8148, n8149, n8150, n8151,
    n8152, n8153, n8154, n8155, n8156, n8157,
    n8158, n8159, n8160, n8161, n8162, n8163,
    n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175,
    n8176, n8177, n8178, n8179, n8180, n8181,
    n8182, n8183, n8184, n8185, n8186, n8187,
    n8188, n8189, n8190, n8191, n8192, n8193,
    n8194, n8195, n8196, n8197, n8198, n8199,
    n8200, n8201, n8202, n8203, n8204, n8205,
    n8206, n8207, n8208, n8209, n8210, n8211,
    n8212, n8213, n8214, n8215, n8216, n8217,
    n8218, n8219, n8220, n8221, n8222, n8223,
    n8224, n8225, n8226, n8227, n8228, n8229,
    n8230, n8231, n8232, n8233, n8234, n8235,
    n8236, n8237, n8238, n8239, n8240, n8241,
    n8242, n8243, n8244, n8245, n8246, n8247,
    n8248, n8249, n8250, n8251, n8252, n8253,
    n8254, n8255, n8256, n8257, n8258, n8259,
    n8260, n8261, n8262, n8263, n8264, n8265,
    n8266, n8267, n8268, n8269, n8270, n8271,
    n8272, n8273, n8274, n8275, n8276, n8277,
    n8278, n8279, n8280, n8281, n8282, n8283,
    n8284, n8285, n8286, n8287, n8288, n8289,
    n8290, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301,
    n8302, n8303, n8304, n8305, n8306, n8307,
    n8308, n8309, n8310, n8311, n8312, n8313,
    n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325,
    n8326, n8327, n8328, n8329, n8330, n8331,
    n8332, n8333, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8342, n8343,
    n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8354, n8355,
    n8356, n8357, n8358, n8359, n8360, n8361,
    n8362, n8363, n8364, n8365, n8366, n8367,
    n8368, n8369, n8370, n8371, n8372, n8373,
    n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385,
    n8386, n8387, n8388, n8389, n8390, n8391,
    n8392, n8393, n8394, n8395, n8396, n8397,
    n8398, n8399, n8400, n8401, n8402, n8403,
    n8404, n8405, n8406, n8407, n8408, n8409,
    n8410, n8411, n8412, n8413, n8414, n8415,
    n8416, n8417, n8418, n8419, n8420, n8421,
    n8422, n8423, n8424, n8425, n8426, n8427,
    n8428, n8429, n8430, n8431, n8432, n8433,
    n8434, n8435, n8436, n8437, n8438, n8439,
    n8440, n8441, n8442, n8443, n8444, n8445,
    n8446, n8447, n8448, n8449, n8450, n8451,
    n8452, n8453, n8454, n8455, n8456, n8457,
    n8458, n8459, n8460, n8461, n8462, n8463,
    n8464, n8465, n8466, n8467, n8468, n8469,
    n8470, n8471, n8472, n8473, n8474, n8475,
    n8476, n8477, n8478, n8479, n8480, n8481,
    n8482, n8483, n8484, n8485, n8486, n8487,
    n8488, n8489, n8490, n8491, n8492, n8493,
    n8494, n8495, n8496, n8497, n8498, n8499,
    n8500, n8501, n8502, n8503, n8504, n8505,
    n8506, n8507, n8508, n8509, n8510, n8511,
    n8512, n8513, n8514, n8515, n8516, n8517,
    n8518, n8519, n8520, n8521, n8522, n8523,
    n8524, n8525, n8526, n8527, n8528, n8529,
    n8530, n8531, n8532, n8533, n8534, n8535,
    n8536, n8537, n8538, n8539, n8540, n8541,
    n8542, n8543, n8544, n8545, n8546, n8547,
    n8548, n8549, n8550, n8551, n8552, n8553,
    n8554, n8555, n8556, n8557, n8558, n8559,
    n8560, n8561, n8562, n8563, n8564, n8565,
    n8566, n8567, n8568, n8569, n8570, n8571,
    n8572, n8573, n8574, n8575, n8576, n8577,
    n8578, n8579, n8580, n8581, n8582, n8583,
    n8584, n8585, n8586, n8587, n8588, n8589,
    n8590, n8591, n8592, n8593, n8594, n8595,
    n8596, n8597, n8598, n8599, n8600, n8601,
    n8602, n8603, n8604, n8605, n8606, n8607,
    n8608, n8609, n8610, n8611, n8612, n8613,
    n8614, n8615, n8616, n8617, n8618, n8619,
    n8620, n8621, n8622, n8623, n8624, n8625,
    n8626, n8627, n8628, n8629, n8630, n8631,
    n8632, n8633, n8634, n8635, n8636, n8637,
    n8638, n8639, n8640, n8641, n8642, n8643,
    n8644, n8645, n8646, n8647, n8648, n8649,
    n8650, n8651, n8652, n8653, n8654, n8655,
    n8656, n8657, n8658, n8659, n8660, n8661,
    n8662, n8663, n8664, n8665, n8666, n8667,
    n8668, n8669, n8670, n8671, n8672, n8673,
    n8674, n8675, n8676, n8677, n8678, n8679,
    n8680, n8681, n8682, n8683, n8684, n8685,
    n8686, n8687, n8688, n8689, n8690, n8691,
    n8692, n8693, n8694, n8695, n8696, n8697,
    n8698, n8699, n8700, n8701, n8702, n8703,
    n8704, n8705, n8706, n8707, n8708, n8709,
    n8710, n8711, n8712, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722,
    n8723, n8724, n8725, n8726, n8727, n8728,
    n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746,
    n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758,
    n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776,
    n8777, n8778, n8779, n8780, n8781, n8782,
    n8783, n8784, n8785, n8786, n8787, n8788,
    n8789, n8790, n8791, n8792, n8793, n8794,
    n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806,
    n8807, n8808, n8809, n8810, n8811, n8812,
    n8813, n8814, n8815, n8816, n8817, n8818,
    n8819, n8820, n8821, n8822, n8823, n8824,
    n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836,
    n8837, n8838, n8839, n8840, n8841, n8842,
    n8843, n8844, n8845, n8846, n8847, n8848,
    n8849, n8850, n8851, n8852, n8853, n8854,
    n8855, n8856, n8857, n8858, n8859, n8860,
    n8861, n8862, n8863, n8864, n8865, n8866,
    n8867, n8868, n8869, n8870, n8871, n8872,
    n8873, n8874, n8875, n8876, n8877, n8878,
    n8879, n8880, n8881, n8882, n8883, n8884,
    n8885, n8886, n8887, n8888, n8889, n8890,
    n8891, n8892, n8893, n8894, n8895, n8896,
    n8897, n8898, n8899, n8900, n8901, n8902,
    n8903, n8904, n8905, n8906, n8907, n8908,
    n8909, n8910, n8911, n8912, n8913, n8914,
    n8915, n8916, n8917, n8918, n8919, n8920,
    n8921, n8922, n8923, n8924, n8925, n8926,
    n8927, n8928, n8929, n8930, n8931, n8932,
    n8933, n8934, n8935, n8936, n8937, n8938,
    n8939, n8940, n8941, n8942, n8943, n8944,
    n8945, n8946, n8947, n8948, n8949, n8950,
    n8951, n8952, n8953, n8954, n8955, n8956,
    n8957, n8958, n8959, n8960, n8961, n8962,
    n8963, n8964, n8965, n8966, n8967, n8968,
    n8969, n8970, n8971, n8972, n8973, n8974,
    n8975, n8976, n8977, n8978, n8979, n8980,
    n8981, n8982, n8983, n8984, n8985, n8986,
    n8987, n8988, n8989, n8990, n8991, n8992,
    n8993, n8994, n8995, n8996, n8997, n8998,
    n8999, n9000, n9001, n9002, n9003, n9004,
    n9005, n9006, n9007, n9008, n9009, n9010,
    n9011, n9012, n9013, n9014, n9015, n9016,
    n9017, n9018, n9019, n9020, n9021, n9022,
    n9023, n9024, n9025, n9026, n9027, n9028,
    n9029, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040,
    n9041, n9042, n9043, n9044, n9045, n9046,
    n9047, n9048, n9049, n9050, n9051, n9052,
    n9053, n9054, n9055, n9056, n9057, n9058,
    n9059, n9060, n9061, n9062, n9063, n9064,
    n9065, n9066, n9067, n9068, n9069, n9070,
    n9071, n9072, n9073, n9074, n9075, n9076,
    n9077, n9078, n9079, n9080, n9081, n9082,
    n9083, n9084, n9085, n9086, n9087, n9088,
    n9089, n9090, n9091, n9092, n9093, n9094,
    n9095, n9096, n9097, n9098, n9099, n9100,
    n9101, n9102, n9103, n9104, n9105, n9106,
    n9107, n9108, n9109, n9110, n9111, n9112,
    n9113, n9114, n9115, n9116, n9117, n9118,
    n9119, n9120, n9121, n9122, n9123, n9124,
    n9125, n9126, n9127, n9128, n9129, n9130,
    n9131, n9132, n9133, n9134, n9135, n9136,
    n9137, n9138, n9139, n9140, n9141, n9142,
    n9143, n9144, n9145, n9146, n9147, n9148,
    n9149, n9150, n9151, n9152, n9153, n9154,
    n9155, n9156, n9157, n9158, n9159, n9160,
    n9161, n9162, n9163, n9164, n9165, n9166,
    n9167, n9168, n9169, n9170, n9171, n9172,
    n9173, n9174, n9175, n9176, n9177, n9178,
    n9179, n9180, n9181, n9182, n9183, n9184,
    n9185, n9186, n9187, n9188, n9189, n9190,
    n9191, n9192, n9193, n9194, n9195, n9196,
    n9197, n9198, n9199, n9200, n9201, n9202,
    n9203, n9204, n9205, n9206, n9207, n9208,
    n9209, n9210, n9211, n9212, n9213, n9214,
    n9215, n9216, n9217, n9218, n9219, n9220,
    n9221, n9222, n9223, n9224, n9225, n9226,
    n9227, n9228, n9229, n9230, n9231, n9232,
    n9233, n9234, n9235, n9236, n9237, n9238,
    n9239, n9240, n9241, n9242, n9243, n9244,
    n9245, n9246, n9247, n9248, n9249, n9250,
    n9251, n9252, n9253, n9254, n9255, n9256,
    n9257, n9258, n9259, n9260, n9261, n9262,
    n9263, n9264, n9265, n9266, n9267, n9268,
    n9269, n9270, n9271, n9272, n9273, n9274,
    n9275, n9276, n9277, n9278, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9286,
    n9287, n9288, n9289, n9290, n9291, n9292,
    n9293, n9294, n9295, n9296, n9297, n9298,
    n9299, n9300, n9301, n9302, n9303, n9304,
    n9305, n9306, n9307, n9308, n9309, n9310,
    n9311, n9312, n9313, n9314, n9315, n9316,
    n9317, n9318, n9319, n9320, n9321, n9322,
    n9323, n9324, n9325, n9326, n9327, n9328,
    n9329, n9330, n9331, n9332, n9333, n9334,
    n9335, n9337, n9338, n9339, n9340, n9341,
    n9342, n9343, n9344, n9345, n9346, n9347,
    n9348, n9349, n9350, n9351, n9352, n9353,
    n9354, n9355, n9356, n9357, n9358, n9359,
    n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371,
    n9372, n9373, n9374, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9382, n9383,
    n9384, n9385, n9386, n9387, n9388, n9389,
    n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401,
    n9402, n9403, n9404, n9405, n9406, n9407,
    n9408, n9409, n9410, n9411, n9412, n9413,
    n9414, n9415, n9416, n9417, n9418, n9419,
    n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431,
    n9432, n9433, n9434, n9435, n9436, n9437,
    n9438, n9439, n9440, n9441, n9442, n9443,
    n9444, n9445, n9446, n9447, n9448, n9449,
    n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461,
    n9462, n9463, n9464, n9465, n9466, n9467,
    n9468, n9469, n9470, n9471, n9472, n9473,
    n9474, n9475, n9476, n9477, n9478, n9479,
    n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491,
    n9492, n9493, n9494, n9495, n9496, n9497,
    n9498, n9499, n9500, n9501, n9502, n9503,
    n9504, n9505, n9506, n9507, n9508, n9509,
    n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521,
    n9522, n9523, n9524, n9525, n9526, n9527,
    n9528, n9529, n9530, n9531, n9532, n9533,
    n9534, n9535, n9536, n9537, n9538, n9539,
    n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551,
    n9552, n9553, n9554, n9555, n9556, n9557,
    n9558, n9559, n9560, n9561, n9562, n9563,
    n9564, n9565, n9566, n9567, n9568, n9569,
    n9570, n9571, n9572, n9573, n9574, n9575,
    n9576, n9577, n9578, n9579, n9580, n9581,
    n9582, n9583, n9584, n9585, n9586, n9587,
    n9588, n9589, n9590, n9591, n9592, n9593,
    n9594, n9595, n9596, n9597, n9598, n9599,
    n9600, n9601, n9602, n9603, n9604, n9605,
    n9606, n9607, n9608, n9609, n9610, n9611,
    n9612, n9613, n9614, n9615, n9616, n9617,
    n9618, n9619, n9620, n9621, n9622, n9623,
    n9624, n9625, n9626, n9627, n9628, n9629,
    n9630, n9631, n9632, n9633, n9634, n9635,
    n9636, n9637, n9638, n9639, n9640, n9641,
    n9642, n9643, n9644, n9645, n9646, n9647,
    n9648, n9649, n9650, n9651, n9652, n9653,
    n9654, n9655, n9656, n9657, n9658, n9659,
    n9660, n9661, n9662, n9663, n9664, n9665,
    n9666, n9667, n9668, n9669, n9670, n9671,
    n9672, n9673, n9674, n9675, n9676, n9677,
    n9678, n9679, n9680, n9681, n9682, n9683,
    n9684, n9685, n9686, n9687, n9688, n9689,
    n9690, n9691, n9692, n9693, n9694, n9695,
    n9696, n9697, n9698, n9699, n9700, n9701,
    n9702, n9703, n9704, n9705, n9706, n9707,
    n9708, n9709, n9710, n9711, n9712, n9713,
    n9714, n9715, n9716, n9717, n9718, n9719,
    n9720, n9721, n9722, n9723, n9724, n9725,
    n9726, n9727, n9728, n9729, n9730, n9731,
    n9732, n9733, n9734, n9735, n9736, n9737,
    n9738, n9739, n9740, n9741, n9742, n9743,
    n9744, n9745, n9746, n9747, n9748, n9749,
    n9750, n9751, n9752, n9753, n9754, n9755,
    n9756, n9757, n9758, n9759, n9760, n9761,
    n9762, n9763, n9764, n9765, n9766, n9767,
    n9768, n9769, n9770, n9771, n9772, n9773,
    n9774, n9775, n9776, n9777, n9778, n9779,
    n9780, n9781, n9782, n9783, n9784, n9785,
    n9786, n9787, n9788, n9789, n9790, n9791,
    n9792, n9793, n9794, n9795, n9796, n9797,
    n9798, n9799, n9800, n9801, n9802, n9803,
    n9804, n9805, n9806, n9807, n9808, n9809,
    n9810, n9811, n9812, n9813, n9814, n9815,
    n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9824, n9825, n9826, n9827,
    n9828, n9829, n9830, n9831, n9832, n9833,
    n9834, n9835, n9836, n9837, n9838, n9839,
    n9840, n9841, n9842, n9843, n9844, n9845,
    n9846, n9847, n9848, n9849, n9850, n9851,
    n9852, n9853, n9854, n9855, n9856, n9857,
    n9858, n9859, n9860, n9861, n9862, n9863,
    n9864, n9865, n9866, n9867, n9868, n9869,
    n9870, n9871, n9872, n9873, n9874, n9875,
    n9876, n9877, n9878, n9879, n9880, n9881,
    n9882, n9883, n9884, n9885, n9886, n9887,
    n9888, n9889, n9890, n9891, n9892, n9893,
    n9894, n9895, n9896, n9897, n9898, n9899,
    n9900, n9901, n9902, n9903, n9904, n9905,
    n9906, n9907, n9908, n9909, n9910, n9911,
    n9912, n9913, n9914, n9915, n9916, n9917,
    n9918, n9919, n9920, n9921, n9922, n9923,
    n9924, n9925, n9926, n9927, n9928, n9929,
    n9930, n9931, n9932, n9933, n9934, n9935,
    n9936, n9937, n9938, n9939, n9940, n9941,
    n9942, n9943, n9944, n9945, n9946, n9947,
    n9948, n9949, n9950, n9951, n9952, n9953,
    n9954, n9955, n9956, n9957, n9958, n9959,
    n9960, n9961, n9962, n9963, n9964, n9965,
    n9966, n9967, n9968, n9969, n9970, n9971,
    n9972, n9973, n9974, n9975, n9976, n9977,
    n9978, n9979, n9980, n9981, n9982, n9983,
    n9984, n9985, n9986, n9987, n9988, n9989,
    n9990, n9991, n9992, n9993, n9994, n9995,
    n9996, n9997, n9998, n9999, n10000, n10001,
    n10002, n10003, n10004, n10005, n10006, n10007,
    n10008, n10009, n10010, n10011, n10012, n10013,
    n10014, n10015, n10016, n10017, n10018, n10019,
    n10020, n10021, n10022, n10023, n10024, n10025,
    n10026, n10027, n10028, n10029, n10030, n10031,
    n10032, n10033, n10034, n10035, n10036, n10037,
    n10038, n10039, n10040, n10041, n10042, n10043,
    n10044, n10045, n10046, n10047, n10048, n10049,
    n10050, n10051, n10052, n10053, n10054, n10055,
    n10056, n10057, n10058, n10059, n10060, n10061,
    n10062, n10063, n10064, n10065, n10066, n10067,
    n10068, n10069, n10070, n10071, n10072, n10073,
    n10074, n10075, n10076, n10077, n10078, n10079,
    n10080, n10081, n10082, n10083, n10084, n10085,
    n10086, n10087, n10088, n10089, n10090, n10091,
    n10092, n10093, n10094, n10095, n10096, n10097,
    n10098, n10099, n10100, n10101, n10102, n10103,
    n10104, n10105, n10106, n10107, n10108, n10109,
    n10110, n10111, n10112, n10113, n10114, n10115,
    n10116, n10117, n10118, n10119, n10120, n10121,
    n10122, n10123, n10124, n10125, n10126, n10127,
    n10128, n10129, n10130, n10131, n10132, n10133,
    n10134, n10135, n10136, n10137, n10138, n10139,
    n10140, n10141, n10142, n10143, n10144, n10145,
    n10146, n10147, n10148, n10149, n10150, n10151,
    n10152, n10153, n10154, n10155, n10156, n10157,
    n10158, n10159, n10160, n10161, n10162, n10163,
    n10164, n10165, n10166, n10167, n10168, n10169,
    n10170, n10171, n10172, n10173, n10174, n10175,
    n10176, n10177, n10178, n10179, n10180, n10181,
    n10182, n10183, n10184, n10185, n10186, n10187,
    n10188, n10189, n10190, n10191, n10192, n10193,
    n10194, n10195, n10196, n10197, n10198, n10199,
    n10200, n10201, n10202, n10203, n10204, n10205,
    n10206, n10207, n10208, n10209, n10210, n10211,
    n10212, n10213, n10214, n10215, n10216, n10217,
    n10218, n10219, n10220, n10221, n10222, n10223,
    n10224, n10225, n10226, n10227, n10228, n10229,
    n10230, n10231, n10232, n10233, n10234, n10235,
    n10236, n10237, n10238, n10239, n10240, n10241,
    n10242, n10243, n10244, n10245, n10246, n10247,
    n10248, n10249, n10250, n10251, n10252, n10253,
    n10254, n10255, n10256, n10257, n10258, n10259,
    n10260, n10261, n10262, n10263, n10264, n10265,
    n10266, n10267, n10268, n10269, n10270, n10271,
    n10272, n10273, n10274, n10275, n10276, n10277,
    n10278, n10279, n10280, n10281, n10282, n10283,
    n10284, n10285, n10286, n10287, n10288, n10289,
    n10290, n10291, n10292, n10293, n10294, n10295,
    n10296, n10297, n10298, n10299, n10300, n10301,
    n10302, n10303, n10304, n10305, n10306, n10307,
    n10308, n10309, n10310, n10311, n10312, n10313,
    n10314, n10315, n10316, n10317, n10318, n10319,
    n10320, n10321, n10322, n10323, n10324, n10325,
    n10326, n10327, n10328, n10329, n10330, n10332,
    n10333, n10334, n10335, n10336, n10337, n10338,
    n10339, n10340, n10341, n10342, n10343, n10344,
    n10345, n10346, n10347, n10348, n10349, n10350,
    n10351, n10352, n10353, n10354, n10355, n10356,
    n10357, n10358, n10359, n10360, n10361, n10362,
    n10363, n10364, n10365, n10366, n10367, n10368,
    n10369, n10370, n10371, n10372, n10373, n10374,
    n10375, n10376, n10377, n10378, n10379, n10380,
    n10381, n10382, n10383, n10384, n10385, n10386,
    n10387, n10388, n10389, n10390, n10391, n10392,
    n10393, n10394, n10395, n10396, n10397, n10398,
    n10399, n10400, n10401, n10402, n10403, n10404,
    n10405, n10406, n10407, n10408, n10409, n10410,
    n10411, n10412, n10413, n10414, n10415, n10416,
    n10417, n10418, n10419, n10420, n10421, n10422,
    n10423, n10424, n10425, n10426, n10427, n10428,
    n10429, n10430, n10431, n10432, n10433, n10434,
    n10435, n10436, n10437, n10438, n10439, n10440,
    n10441, n10442, n10443, n10444, n10445, n10446,
    n10447, n10448, n10449, n10450, n10451, n10452,
    n10453, n10454, n10455, n10456, n10457, n10458,
    n10459, n10460, n10461, n10462, n10463, n10464,
    n10465, n10466, n10467, n10468, n10469, n10470,
    n10471, n10472, n10473, n10474, n10475, n10476,
    n10477, n10478, n10479, n10480, n10481, n10482,
    n10483, n10484, n10485, n10486, n10487, n10488,
    n10489, n10490, n10491, n10492, n10493, n10494,
    n10495, n10496, n10497, n10498, n10499, n10500,
    n10501, n10502, n10503, n10504, n10505, n10506,
    n10507, n10508, n10509, n10510, n10511, n10512,
    n10513, n10514, n10515, n10516, n10517, n10518,
    n10519, n10520, n10521, n10522, n10523, n10524,
    n10525, n10526, n10527, n10528, n10529, n10530,
    n10531, n10532, n10533, n10534, n10535, n10536,
    n10537, n10538, n10539, n10540, n10541, n10542,
    n10543, n10544, n10545, n10546, n10547, n10548,
    n10549, n10550, n10551, n10552, n10553, n10554,
    n10555, n10556, n10557, n10558, n10559, n10560,
    n10561, n10562, n10563, n10564, n10565, n10566,
    n10567, n10568, n10569, n10570, n10571, n10572,
    n10573, n10574, n10575, n10576, n10577, n10578,
    n10579, n10580, n10581, n10582, n10583, n10584,
    n10585, n10586, n10587, n10588, n10589, n10590,
    n10591, n10592, n10593, n10594, n10595, n10596,
    n10597, n10598, n10599, n10600, n10601, n10602,
    n10603, n10604, n10605, n10606, n10607, n10608,
    n10609, n10610, n10611, n10612, n10613, n10614,
    n10615, n10616, n10617, n10618, n10619, n10620,
    n10621, n10622, n10623, n10624, n10625, n10626,
    n10627, n10628, n10629, n10630, n10631, n10632,
    n10633, n10634, n10635, n10636, n10637, n10638,
    n10639, n10640, n10641, n10642, n10643, n10644,
    n10645, n10646, n10647, n10648, n10649, n10650,
    n10651, n10652, n10653, n10654, n10655, n10656,
    n10657, n10658, n10659, n10660, n10661, n10662,
    n10663, n10664, n10665, n10666, n10667, n10668,
    n10669, n10670, n10671, n10672, n10673, n10674,
    n10675, n10676, n10677, n10678, n10679, n10680,
    n10681, n10682, n10683, n10684, n10685, n10686,
    n10687, n10688, n10689, n10690, n10691, n10692,
    n10693, n10694, n10695, n10696, n10697, n10698,
    n10699, n10700, n10701, n10702, n10703, n10704,
    n10705, n10706, n10707, n10708, n10709, n10710,
    n10711, n10712, n10713, n10714, n10715, n10716,
    n10717, n10718, n10719, n10720, n10721, n10722,
    n10723, n10724, n10725, n10726, n10727, n10728,
    n10729, n10730, n10731, n10732, n10733, n10734,
    n10735, n10736, n10737, n10738, n10739, n10740,
    n10741, n10742, n10743, n10744, n10745, n10746,
    n10747, n10748, n10749, n10750, n10751, n10752,
    n10753, n10754, n10755, n10756, n10757, n10758,
    n10759, n10760, n10761, n10762, n10763, n10764,
    n10765, n10766, n10767, n10768, n10769, n10770,
    n10771, n10772, n10773, n10774, n10775, n10776,
    n10777, n10778, n10779, n10780, n10781, n10782,
    n10783, n10784, n10785, n10786, n10787, n10788,
    n10789, n10790, n10791, n10792, n10793, n10794,
    n10795, n10796, n10797, n10798, n10799, n10800,
    n10801, n10802, n10803, n10804, n10805, n10806,
    n10807, n10808, n10809, n10810, n10811, n10812,
    n10813, n10814, n10815, n10816, n10817, n10818,
    n10819, n10820, n10821, n10822, n10823, n10824,
    n10825, n10826, n10827, n10828, n10829, n10830,
    n10831, n10832, n10833, n10834, n10835, n10836,
    n10837, n10838, n10839, n10840, n10841, n10842,
    n10843, n10844, n10845, n10846, n10847, n10848,
    n10849, n10850, n10851, n10852, n10853, n10854,
    n10855, n10856, n10857, n10858, n10859, n10860,
    n10861, n10862, n10863, n10864, n10865, n10866,
    n10867, n10868, n10869, n10870, n10871, n10872,
    n10873, n10874, n10875, n10876, n10877, n10878,
    n10879, n10880, n10881, n10882, n10883, n10884,
    n10885, n10886, n10887, n10888, n10889, n10890,
    n10891, n10892, n10893, n10894, n10895, n10896,
    n10897, n10898, n10899, n10900, n10901, n10902,
    n10903, n10904, n10905, n10906, n10907, n10908,
    n10909, n10910, n10911, n10912, n10913, n10914,
    n10915, n10916, n10917, n10918, n10919, n10920,
    n10921, n10922, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10945,
    n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963,
    n10964, n10965, n10966, n10967, n10968, n10969,
    n10970, n10971, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10981,
    n10982, n10983, n10984, n10985, n10986, n10987,
    n10988, n10989, n10990, n10991, n10992, n10993,
    n10994, n10995, n10996, n10997, n10998, n10999,
    n11000, n11001, n11002, n11003, n11004, n11005,
    n11006, n11007, n11008, n11009, n11010, n11011,
    n11012, n11013, n11014, n11015, n11016, n11017,
    n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11025, n11026, n11027, n11028, n11029,
    n11030, n11031, n11032, n11033, n11034, n11035,
    n11036, n11037, n11038, n11039, n11040, n11041,
    n11042, n11043, n11044, n11045, n11046, n11047,
    n11048, n11049, n11050, n11051, n11052, n11053,
    n11054, n11055, n11056, n11057, n11058, n11059,
    n11060, n11061, n11062, n11063, n11064, n11065,
    n11066, n11067, n11068, n11069, n11070, n11071,
    n11072, n11073, n11074, n11075, n11076, n11077,
    n11078, n11079, n11080, n11081, n11082, n11083,
    n11084, n11085, n11086, n11087, n11088, n11089,
    n11090, n11091, n11092, n11093, n11094, n11095,
    n11096, n11097, n11098, n11099, n11100, n11101,
    n11102, n11103, n11104, n11105, n11106, n11107,
    n11108, n11109, n11110, n11111, n11112, n11113,
    n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125,
    n11126, n11127, n11128, n11129, n11130, n11131,
    n11132, n11133, n11134, n11135, n11136, n11137,
    n11138, n11139, n11140, n11141, n11142, n11143,
    n11144, n11145, n11146, n11147, n11148, n11149,
    n11150, n11151, n11152, n11153, n11154, n11155,
    n11156, n11157, n11158, n11159, n11160, n11161,
    n11162, n11163, n11164, n11165, n11166, n11167,
    n11168, n11169, n11170, n11171, n11172, n11173,
    n11174, n11175, n11176, n11177, n11178, n11179,
    n11180, n11181, n11182, n11183, n11184, n11185,
    n11186, n11187, n11188, n11189, n11190, n11191,
    n11192, n11193, n11194, n11195, n11196, n11197,
    n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209,
    n11210, n11211, n11212, n11213, n11214, n11215,
    n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227,
    n11228, n11229, n11230, n11231, n11232, n11233,
    n11234, n11235, n11236, n11237, n11238, n11239,
    n11240, n11241, n11242, n11243, n11244, n11245,
    n11246, n11247, n11248, n11249, n11250, n11251,
    n11252, n11253, n11254, n11255, n11256, n11257,
    n11258, n11259, n11260, n11261, n11262, n11263,
    n11264, n11265, n11266, n11267, n11268, n11269,
    n11270, n11271, n11272, n11273, n11274, n11275,
    n11276, n11277, n11278, n11279, n11280, n11281,
    n11282, n11283, n11284, n11285, n11286, n11287,
    n11288, n11289, n11290, n11291, n11292, n11293,
    n11294, n11295, n11296, n11297, n11298, n11299,
    n11300, n11301, n11302, n11303, n11304, n11305,
    n11306, n11307, n11308, n11309, n11310, n11311,
    n11312, n11313, n11314, n11315, n11316, n11317,
    n11318, n11319, n11320, n11321, n11322, n11323,
    n11324, n11325, n11326, n11327, n11328, n11329,
    n11330, n11331, n11332, n11333, n11334, n11335,
    n11336, n11337, n11338, n11339, n11340, n11341,
    n11342, n11343, n11344, n11345, n11346, n11347,
    n11348, n11349, n11350, n11351, n11352, n11353,
    n11354, n11355, n11356, n11357, n11358, n11359,
    n11360, n11361, n11362, n11363, n11364, n11365,
    n11366, n11367, n11368, n11369, n11370, n11371,
    n11372, n11373, n11374, n11375, n11376, n11377,
    n11378, n11379, n11380, n11381, n11382, n11383,
    n11384, n11385, n11386, n11387, n11388, n11389,
    n11390, n11391, n11392, n11393, n11394, n11395,
    n11396, n11397, n11398, n11399, n11400, n11401,
    n11402, n11403, n11404, n11405, n11406, n11407,
    n11408, n11409, n11410, n11411, n11412, n11413,
    n11414, n11415, n11416, n11417, n11418, n11419,
    n11420, n11421, n11422, n11423, n11424, n11425,
    n11426, n11427, n11428, n11429, n11430, n11431,
    n11432, n11433, n11434, n11435, n11436, n11437,
    n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449,
    n11450, n11451, n11452, n11453, n11454, n11455,
    n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473,
    n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497,
    n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515,
    n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527,
    n11528, n11529, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545,
    n11546, n11547, n11548, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575,
    n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11590, n11591, n11592, n11593,
    n11594, n11595, n11596, n11597, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618,
    n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630,
    n11631, n11632, n11633, n11634, n11635, n11636,
    n11637, n11638, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11648,
    n11649, n11650, n11651, n11652, n11653, n11654,
    n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666,
    n11667, n11668, n11669, n11670, n11671, n11672,
    n11673, n11674, n11675, n11676, n11677, n11678,
    n11679, n11680, n11681, n11682, n11683, n11684,
    n11685, n11686, n11687, n11688, n11689, n11690,
    n11691, n11692, n11693, n11694, n11695, n11696,
    n11697, n11698, n11699, n11700, n11701, n11702,
    n11703, n11704, n11705, n11706, n11707, n11708,
    n11709, n11710, n11711, n11712, n11713, n11714,
    n11715, n11716, n11717, n11718, n11719, n11720,
    n11721, n11722, n11723, n11724, n11725, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756,
    n11757, n11758, n11759, n11760, n11761, n11762,
    n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774,
    n11775, n11776, n11777, n11778, n11779, n11780,
    n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792,
    n11793, n11794, n11795, n11796, n11797, n11798,
    n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810,
    n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12217, n12218, n12219,
    n12220, n12221, n12222, n12223, n12224, n12225,
    n12226, n12227, n12228, n12229, n12230, n12231,
    n12232, n12233, n12234, n12235, n12236, n12237,
    n12238, n12239, n12240, n12241, n12242, n12243,
    n12244, n12245, n12246, n12247, n12248, n12249,
    n12250, n12251, n12252, n12253, n12254, n12255,
    n12256, n12257, n12258, n12259, n12260, n12261,
    n12262, n12263, n12264, n12265, n12266, n12267,
    n12268, n12269, n12270, n12271, n12272, n12273,
    n12274, n12275, n12276, n12277, n12278, n12279,
    n12280, n12281, n12282, n12283, n12284, n12285,
    n12286, n12287, n12288, n12289, n12290, n12291,
    n12292, n12293, n12294, n12295, n12296, n12297,
    n12298, n12299, n12300, n12301, n12302, n12303,
    n12304, n12305, n12306, n12307, n12308, n12309,
    n12310, n12311, n12312, n12313, n12314, n12315,
    n12316, n12317, n12318, n12319, n12320, n12321,
    n12322, n12323, n12324, n12325, n12326, n12327,
    n12328, n12329, n12330, n12331, n12332, n12333,
    n12334, n12335, n12336, n12337, n12338, n12339,
    n12340, n12341, n12342, n12343, n12344, n12345,
    n12346, n12347, n12348, n12349, n12350, n12351,
    n12352, n12353, n12354, n12355, n12356, n12357,
    n12358, n12359, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369,
    n12370, n12371, n12372, n12373, n12374, n12375,
    n12376, n12377, n12378, n12379, n12380, n12381,
    n12382, n12383, n12384, n12385, n12386, n12387,
    n12388, n12389, n12390, n12391, n12392, n12393,
    n12394, n12395, n12396, n12397, n12398, n12399,
    n12400, n12401, n12402, n12403, n12404, n12405,
    n12406, n12407, n12408, n12409, n12410, n12411,
    n12412, n12413, n12414, n12415, n12416, n12417,
    n12418, n12419, n12420, n12421, n12422, n12423,
    n12424, n12425, n12426, n12427, n12428, n12429,
    n12430, n12431, n12432, n12433, n12434, n12435,
    n12436, n12437, n12438, n12439, n12440, n12441,
    n12442, n12443, n12444, n12445, n12446, n12447,
    n12448, n12449, n12450, n12451, n12452, n12453,
    n12454, n12455, n12456, n12457, n12458, n12459,
    n12460, n12461, n12462, n12463, n12464, n12465,
    n12466, n12467, n12468, n12469, n12470, n12471,
    n12472, n12473, n12474, n12475, n12476, n12477,
    n12478, n12479, n12480, n12481, n12482, n12483,
    n12484, n12485, n12486, n12487, n12488, n12489,
    n12490, n12491, n12492, n12493, n12494, n12495,
    n12496, n12497, n12498, n12499, n12500, n12501,
    n12502, n12503, n12504, n12505, n12506, n12507,
    n12508, n12509, n12510, n12511, n12512, n12513,
    n12514, n12515, n12516, n12517, n12518, n12519,
    n12520, n12521, n12522, n12523, n12524, n12525,
    n12526, n12527, n12528, n12529, n12530, n12531,
    n12532, n12533, n12534, n12535, n12536, n12537,
    n12538, n12539, n12540, n12541, n12542, n12543,
    n12544, n12545, n12546, n12547, n12548, n12549,
    n12550, n12551, n12552, n12553, n12554, n12555,
    n12556, n12557, n12558, n12559, n12560, n12561,
    n12562, n12563, n12564, n12565, n12566, n12567,
    n12568, n12569, n12570, n12571, n12572, n12573,
    n12574, n12575, n12576, n12577, n12578, n12579,
    n12580, n12581, n12582, n12583, n12584, n12585,
    n12586, n12587, n12588, n12589, n12590, n12591,
    n12592, n12593, n12594, n12595, n12596, n12597,
    n12598, n12599, n12600, n12601, n12602, n12603,
    n12604, n12605, n12606, n12607, n12608, n12609,
    n12610, n12611, n12612, n12613, n12614, n12615,
    n12616, n12617, n12618, n12619, n12620, n12621,
    n12622, n12623, n12624, n12625, n12626, n12627,
    n12628, n12629, n12630, n12631, n12632, n12633,
    n12634, n12635, n12636, n12637, n12638, n12639,
    n12640, n12641, n12642, n12643, n12644, n12645,
    n12646, n12647, n12648, n12649, n12650, n12651,
    n12652, n12653, n12654, n12655, n12656, n12657,
    n12658, n12659, n12660, n12661, n12662, n12663,
    n12664, n12665, n12666, n12667, n12668, n12669,
    n12670, n12671, n12672, n12673, n12674, n12675,
    n12676, n12677, n12678, n12679, n12680, n12681,
    n12682, n12683, n12684, n12685, n12686, n12687,
    n12688, n12689, n12690, n12691, n12692, n12693,
    n12694, n12695, n12696, n12697, n12698, n12699,
    n12700, n12701, n12702, n12703, n12704, n12705,
    n12706, n12707, n12708, n12709, n12710, n12711,
    n12712, n12713, n12714, n12715, n12716, n12717,
    n12718, n12719, n12720, n12721, n12722, n12723,
    n12724, n12725, n12726, n12727, n12728, n12729,
    n12730, n12731, n12732, n12733, n12734, n12735,
    n12736, n12737, n12738, n12739, n12740, n12741,
    n12742, n12743, n12744, n12745, n12746, n12747,
    n12748, n12749, n12750, n12751, n12752, n12753,
    n12754, n12755, n12756, n12757, n12758, n12759,
    n12760, n12761, n12762, n12763, n12764, n12765,
    n12766, n12767, n12768, n12769, n12770, n12771,
    n12772, n12773, n12774, n12775, n12776, n12777,
    n12778, n12779, n12780, n12781, n12782, n12783,
    n12784, n12785, n12786, n12787, n12788, n12789,
    n12790, n12791, n12792, n12793, n12794, n12795,
    n12796, n12797, n12798, n12799, n12800, n12802,
    n12803, n12804, n12805, n12806, n12807, n12808,
    n12809, n12810, n12811, n12812, n12813, n12814,
    n12815, n12816, n12817, n12818, n12819, n12820,
    n12821, n12822, n12823, n12824, n12825, n12826,
    n12827, n12828, n12829, n12830, n12831, n12832,
    n12833, n12834, n12835, n12836, n12837, n12838,
    n12839, n12840, n12841, n12842, n12843, n12844,
    n12845, n12846, n12847, n12848, n12849, n12850,
    n12851, n12852, n12853, n12854, n12855, n12856,
    n12857, n12858, n12859, n12860, n12861, n12862,
    n12863, n12864, n12865, n12866, n12867, n12868,
    n12869, n12870, n12871, n12872, n12873, n12874,
    n12875, n12876, n12877, n12878, n12879, n12880,
    n12881, n12882, n12883, n12884, n12885, n12886,
    n12887, n12888, n12889, n12890, n12891, n12892,
    n12893, n12894, n12895, n12896, n12897, n12898,
    n12899, n12900, n12901, n12902, n12903, n12904,
    n12905, n12906, n12907, n12908, n12909, n12910,
    n12911, n12912, n12913, n12914, n12915, n12916,
    n12917, n12918, n12919, n12920, n12921, n12922,
    n12923, n12924, n12925, n12926, n12927, n12928,
    n12929, n12930, n12931, n12932, n12933, n12934,
    n12935, n12936, n12937, n12938, n12939, n12940,
    n12941, n12942, n12943, n12944, n12945, n12946,
    n12947, n12948, n12949, n12950, n12951, n12952,
    n12953, n12954, n12955, n12956, n12957, n12958,
    n12959, n12960, n12961, n12962, n12963, n12964,
    n12965, n12966, n12967, n12968, n12969, n12970,
    n12971, n12972, n12973, n12974, n12975, n12976,
    n12977, n12978, n12979, n12980, n12981, n12982,
    n12983, n12984, n12985, n12986, n12987, n12988,
    n12989, n12990, n12991, n12992, n12993, n12994,
    n12995, n12996, n12997, n12998, n12999, n13000,
    n13001, n13002, n13003, n13004, n13005, n13006,
    n13007, n13008, n13009, n13010, n13011, n13012,
    n13013, n13014, n13015, n13016, n13017, n13018,
    n13019, n13020, n13021, n13022, n13023, n13024,
    n13025, n13026, n13027, n13028, n13029, n13030,
    n13031, n13032, n13033, n13034, n13035, n13036,
    n13037, n13038, n13039, n13040, n13041, n13042,
    n13043, n13044, n13045, n13046, n13047, n13048,
    n13049, n13050, n13051, n13052, n13053, n13054,
    n13055, n13056, n13057, n13058, n13059, n13060,
    n13061, n13062, n13063, n13064, n13065, n13066,
    n13067, n13068, n13069, n13070, n13071, n13072,
    n13073, n13074, n13075, n13076, n13077, n13078,
    n13079, n13080, n13081, n13082, n13083, n13084,
    n13085, n13086, n13087, n13088, n13089, n13090,
    n13091, n13092, n13093, n13094, n13095, n13096,
    n13097, n13098, n13099, n13100, n13101, n13102,
    n13103, n13104, n13105, n13106, n13107, n13108,
    n13109, n13110, n13111, n13112, n13113, n13114,
    n13115, n13116, n13117, n13118, n13119, n13120,
    n13121, n13122, n13123, n13124, n13125, n13126,
    n13127, n13128, n13129, n13130, n13131, n13132,
    n13133, n13134, n13135, n13136, n13137, n13138,
    n13139, n13140, n13141, n13142, n13143, n13144,
    n13145, n13146, n13147, n13148, n13149, n13150,
    n13151, n13152, n13153, n13154, n13155, n13156,
    n13157, n13158, n13159, n13160, n13161, n13162,
    n13163, n13164, n13165, n13166, n13167, n13168,
    n13169, n13170, n13171, n13172, n13173, n13174,
    n13175, n13176, n13177, n13178, n13179, n13180,
    n13181, n13182, n13183, n13184, n13185, n13186,
    n13187, n13188, n13189, n13190, n13191, n13192,
    n13193, n13194, n13195, n13196, n13197, n13198,
    n13199, n13200, n13201, n13202, n13203, n13204,
    n13205, n13206, n13207, n13208, n13209, n13210,
    n13211, n13212, n13213, n13214, n13215, n13216,
    n13217, n13218, n13219, n13220, n13221, n13222,
    n13223, n13224, n13225, n13226, n13227, n13228,
    n13229, n13230, n13231, n13232, n13233, n13234,
    n13235, n13236, n13237, n13238, n13239, n13240,
    n13241, n13242, n13243, n13244, n13245, n13246,
    n13247, n13248, n13249, n13250, n13251, n13252,
    n13253, n13254, n13255, n13256, n13257, n13258,
    n13259, n13260, n13261, n13262, n13263, n13264,
    n13265, n13266, n13267, n13268, n13269, n13270,
    n13271, n13272, n13273, n13274, n13275, n13276,
    n13277, n13278, n13279, n13280, n13281, n13282,
    n13283, n13284, n13285, n13286, n13287, n13288,
    n13289, n13290, n13291, n13292, n13293, n13294,
    n13295, n13296, n13297, n13298, n13299, n13300,
    n13301, n13302, n13303, n13304, n13305, n13306,
    n13307, n13308, n13309, n13310, n13311, n13312,
    n13313, n13314, n13315, n13316, n13317, n13318,
    n13319, n13320, n13321, n13322, n13323, n13324,
    n13325, n13326, n13327, n13328, n13329, n13330,
    n13331, n13332, n13333, n13334, n13335, n13336,
    n13337, n13338, n13339, n13340, n13341, n13342,
    n13343, n13344, n13345, n13346, n13347, n13348,
    n13349, n13350, n13351, n13352, n13353, n13354,
    n13355, n13356, n13357, n13358, n13359, n13360,
    n13361, n13362, n13363, n13364, n13365, n13366,
    n13367, n13368, n13369, n13370, n13371, n13372,
    n13373, n13374, n13375, n13376, n13377, n13378,
    n13379, n13380, n13381, n13382, n13383, n13384,
    n13385, n13386, n13387, n13388, n13389, n13390,
    n13391, n13392, n13393, n13394, n13395, n13396,
    n13397, n13398, n13399, n13400, n13401, n13402,
    n13403, n13404, n13405, n13406, n13407, n13408,
    n13409, n13410, n13411, n13412, n13413, n13414,
    n13415, n13416, n13417, n13418, n13419, n13420,
    n13421, n13422, n13423, n13424, n13425, n13426,
    n13427, n13428, n13429, n13430, n13431, n13432,
    n13433, n13434, n13435, n13436, n13438, n13439,
    n13440, n13441, n13442, n13443, n13444, n13445,
    n13446, n13447, n13448, n13449, n13450, n13451,
    n13452, n13453, n13454, n13455, n13456, n13457,
    n13458, n13459, n13460, n13461, n13462, n13463,
    n13464, n13465, n13466, n13467, n13468, n13469,
    n13470, n13471, n13472, n13473, n13474, n13475,
    n13476, n13477, n13478, n13479, n13480, n13481,
    n13482, n13483, n13484, n13485, n13486, n13487,
    n13488, n13489, n13490, n13491, n13492, n13493,
    n13494, n13495, n13496, n13497, n13498, n13499,
    n13500, n13501, n13502, n13503, n13504, n13505,
    n13506, n13507, n13508, n13509, n13510, n13511,
    n13512, n13513, n13514, n13515, n13516, n13517,
    n13518, n13519, n13520, n13521, n13522, n13523,
    n13524, n13525, n13526, n13527, n13528, n13529,
    n13530, n13531, n13532, n13533, n13534, n13535,
    n13536, n13537, n13538, n13539, n13540, n13541,
    n13542, n13543, n13544, n13545, n13546, n13547,
    n13548, n13549, n13550, n13551, n13552, n13553,
    n13554, n13555, n13556, n13557, n13558, n13559,
    n13560, n13561, n13562, n13563, n13564, n13565,
    n13566, n13567, n13568, n13569, n13570, n13571,
    n13572, n13573, n13574, n13575, n13576, n13577,
    n13578, n13579, n13580, n13581, n13582, n13583,
    n13584, n13585, n13586, n13587, n13588, n13589,
    n13590, n13591, n13592, n13593, n13594, n13595,
    n13596, n13597, n13598, n13599, n13600, n13601,
    n13602, n13603, n13604, n13605, n13606, n13607,
    n13608, n13609, n13610, n13611, n13612, n13613,
    n13614, n13615, n13616, n13617, n13618, n13619,
    n13620, n13621, n13622, n13623, n13624, n13625,
    n13626, n13627, n13628, n13629, n13630, n13631,
    n13632, n13633, n13634, n13635, n13636, n13637,
    n13638, n13639, n13640, n13641, n13642, n13643,
    n13644, n13645, n13646, n13647, n13648, n13649,
    n13650, n13651, n13652, n13653, n13654, n13655,
    n13656, n13657, n13658, n13659, n13660, n13661,
    n13662, n13663, n13664, n13665, n13666, n13667,
    n13668, n13669, n13670, n13671, n13672, n13673,
    n13674, n13675, n13676, n13677, n13678, n13679,
    n13680, n13681, n13682, n13683, n13684, n13685,
    n13686, n13687, n13688, n13689, n13690, n13691,
    n13692, n13693, n13694, n13695, n13696, n13697,
    n13698, n13699, n13700, n13701, n13702, n13703,
    n13704, n13705, n13706, n13707, n13708, n13709,
    n13710, n13711, n13712, n13713, n13714, n13715,
    n13716, n13717, n13718, n13719, n13720, n13721,
    n13722, n13723, n13724, n13725, n13726, n13727,
    n13728, n13729, n13730, n13731, n13732, n13733,
    n13734, n13735, n13736, n13737, n13738, n13739,
    n13740, n13741, n13742, n13743, n13744, n13745,
    n13746, n13747, n13748, n13749, n13750, n13751,
    n13752, n13753, n13754, n13755, n13756, n13757,
    n13758, n13759, n13760, n13761, n13762, n13763,
    n13764, n13765, n13766, n13767, n13768, n13769,
    n13770, n13771, n13772, n13773, n13774, n13775,
    n13776, n13777, n13778, n13779, n13780, n13781,
    n13782, n13783, n13784, n13785, n13786, n13787,
    n13788, n13789, n13790, n13791, n13792, n13793,
    n13794, n13795, n13796, n13797, n13798, n13799,
    n13800, n13801, n13802, n13803, n13804, n13805,
    n13806, n13807, n13808, n13809, n13810, n13811,
    n13812, n13813, n13814, n13815, n13816, n13817,
    n13818, n13819, n13820, n13821, n13822, n13823,
    n13824, n13825, n13826, n13827, n13828, n13829,
    n13830, n13831, n13832, n13833, n13834, n13835,
    n13836, n13837, n13838, n13839, n13840, n13841,
    n13842, n13843, n13844, n13845, n13846, n13847,
    n13848, n13849, n13850, n13851, n13852, n13853,
    n13854, n13855, n13856, n13857, n13858, n13859,
    n13860, n13861, n13862, n13863, n13864, n13865,
    n13866, n13867, n13868, n13869, n13870, n13871,
    n13872, n13873, n13874, n13875, n13876, n13877,
    n13878, n13879, n13880, n13881, n13882, n13883,
    n13884, n13885, n13886, n13887, n13888, n13889,
    n13890, n13891, n13892, n13893, n13894, n13895,
    n13896, n13897, n13898, n13899, n13900, n13901,
    n13902, n13903, n13904, n13905, n13906, n13907,
    n13908, n13909, n13910, n13911, n13912, n13913,
    n13914, n13915, n13916, n13917, n13918, n13919,
    n13920, n13921, n13922, n13923, n13924, n13925,
    n13926, n13927, n13928, n13929, n13930, n13931,
    n13932, n13933, n13934, n13935, n13936, n13937,
    n13938, n13939, n13940, n13941, n13942, n13943,
    n13944, n13945, n13946, n13947, n13948, n13949,
    n13950, n13951, n13952, n13953, n13954, n13955,
    n13956, n13957, n13958, n13959, n13960, n13961,
    n13962, n13963, n13964, n13965, n13966, n13967,
    n13968, n13969, n13970, n13971, n13972, n13973,
    n13974, n13975, n13976, n13977, n13978, n13979,
    n13980, n13981, n13982, n13983, n13984, n13985,
    n13986, n13987, n13988, n13989, n13990, n13991,
    n13992, n13993, n13994, n13995, n13996, n13997,
    n13998, n13999, n14000, n14001, n14002, n14003,
    n14004, n14005, n14006, n14007, n14008, n14009,
    n14010, n14011, n14012, n14013, n14014, n14015,
    n14016, n14017, n14018, n14019, n14020, n14021,
    n14022, n14023, n14024, n14025, n14026, n14027,
    n14028, n14029, n14030, n14031, n14032, n14033,
    n14034, n14035, n14036, n14037, n14038, n14039,
    n14040, n14041, n14042, n14043, n14044, n14046,
    n14047, n14048, n14049, n14050, n14051, n14052,
    n14053, n14054, n14055, n14056, n14057, n14058,
    n14059, n14060, n14061, n14062, n14063, n14064,
    n14065, n14066, n14067, n14068, n14069, n14070,
    n14071, n14072, n14073, n14074, n14075, n14076,
    n14077, n14078, n14079, n14080, n14081, n14082,
    n14083, n14084, n14085, n14086, n14087, n14088,
    n14089, n14090, n14091, n14092, n14093, n14094,
    n14095, n14096, n14097, n14098, n14099, n14100,
    n14101, n14102, n14103, n14104, n14105, n14106,
    n14107, n14108, n14109, n14110, n14111, n14112,
    n14113, n14114, n14115, n14116, n14117, n14118,
    n14119, n14120, n14121, n14122, n14123, n14124,
    n14125, n14126, n14127, n14128, n14129, n14130,
    n14131, n14132, n14133, n14134, n14135, n14136,
    n14137, n14138, n14139, n14140, n14141, n14142,
    n14143, n14144, n14145, n14146, n14147, n14148,
    n14149, n14150, n14151, n14152, n14153, n14154,
    n14155, n14156, n14157, n14158, n14159, n14160,
    n14161, n14162, n14163, n14164, n14165, n14166,
    n14167, n14168, n14169, n14170, n14171, n14172,
    n14173, n14174, n14175, n14176, n14177, n14178,
    n14179, n14180, n14181, n14182, n14183, n14184,
    n14185, n14186, n14187, n14188, n14189, n14190,
    n14191, n14192, n14193, n14194, n14195, n14196,
    n14197, n14198, n14199, n14200, n14201, n14202,
    n14203, n14204, n14205, n14206, n14207, n14208,
    n14209, n14210, n14211, n14212, n14213, n14214,
    n14215, n14216, n14217, n14218, n14219, n14220,
    n14221, n14222, n14223, n14224, n14225, n14226,
    n14227, n14228, n14229, n14230, n14231, n14232,
    n14233, n14234, n14235, n14236, n14237, n14238,
    n14239, n14240, n14241, n14242, n14243, n14244,
    n14245, n14246, n14247, n14248, n14249, n14250,
    n14251, n14252, n14253, n14254, n14255, n14256,
    n14257, n14258, n14259, n14260, n14261, n14262,
    n14263, n14264, n14265, n14266, n14267, n14268,
    n14269, n14270, n14271, n14272, n14273, n14274,
    n14275, n14276, n14277, n14278, n14279, n14280,
    n14281, n14282, n14283, n14284, n14285, n14286,
    n14287, n14288, n14289, n14290, n14291, n14292,
    n14293, n14294, n14295, n14296, n14297, n14298,
    n14299, n14300, n14301, n14302, n14303, n14304,
    n14305, n14306, n14307, n14308, n14309, n14310,
    n14311, n14312, n14313, n14314, n14315, n14316,
    n14317, n14318, n14319, n14320, n14321, n14322,
    n14323, n14324, n14325, n14326, n14327, n14328,
    n14329, n14330, n14331, n14332, n14333, n14334,
    n14335, n14336, n14337, n14338, n14339, n14340,
    n14341, n14342, n14343, n14344, n14345, n14346,
    n14347, n14348, n14349, n14350, n14351, n14352,
    n14353, n14354, n14355, n14356, n14357, n14358,
    n14359, n14360, n14361, n14362, n14363, n14364,
    n14365, n14366, n14367, n14368, n14369, n14370,
    n14371, n14372, n14373, n14374, n14375, n14376,
    n14377, n14378, n14379, n14380, n14381, n14382,
    n14383, n14384, n14385, n14386, n14387, n14388,
    n14389, n14390, n14391, n14392, n14393, n14394,
    n14395, n14396, n14397, n14398, n14399, n14400,
    n14401, n14402, n14403, n14404, n14405, n14406,
    n14407, n14408, n14409, n14410, n14411, n14412,
    n14413, n14414, n14415, n14416, n14417, n14418,
    n14419, n14420, n14421, n14422, n14423, n14424,
    n14425, n14426, n14427, n14428, n14429, n14430,
    n14431, n14432, n14433, n14434, n14435, n14436,
    n14437, n14438, n14439, n14440, n14441, n14442,
    n14443, n14444, n14445, n14446, n14447, n14448,
    n14449, n14450, n14451, n14452, n14453, n14454,
    n14455, n14456, n14457, n14458, n14459, n14460,
    n14461, n14462, n14463, n14464, n14465, n14466,
    n14467, n14468, n14469, n14470, n14471, n14472,
    n14473, n14474, n14475, n14476, n14477, n14478,
    n14479, n14480, n14481, n14482, n14483, n14484,
    n14485, n14486, n14487, n14488, n14489, n14490,
    n14491, n14492, n14493, n14494, n14495, n14496,
    n14497, n14498, n14499, n14500, n14501, n14502,
    n14503, n14504, n14505, n14506, n14507, n14508,
    n14509, n14510, n14511, n14512, n14513, n14514,
    n14515, n14516, n14517, n14518, n14519, n14520,
    n14521, n14522, n14523, n14524, n14525, n14526,
    n14527, n14528, n14529, n14530, n14531, n14532,
    n14533, n14534, n14535, n14536, n14537, n14538,
    n14539, n14540, n14541, n14542, n14543, n14544,
    n14545, n14546, n14547, n14548, n14549, n14550,
    n14551, n14552, n14553, n14554, n14555, n14556,
    n14557, n14558, n14559, n14560, n14561, n14562,
    n14563, n14564, n14565, n14566, n14567, n14568,
    n14569, n14570, n14571, n14572, n14573, n14574,
    n14575, n14576, n14577, n14578, n14579, n14580,
    n14581, n14582, n14583, n14584, n14585, n14586,
    n14587, n14588, n14589, n14590, n14591, n14592,
    n14593, n14594, n14595, n14596, n14597, n14598,
    n14599, n14600, n14601, n14602, n14603, n14604,
    n14605, n14606, n14607, n14608, n14609, n14610,
    n14611, n14612, n14613, n14614, n14615, n14616,
    n14617, n14618, n14619, n14620, n14621, n14622,
    n14623, n14624, n14625, n14626, n14627, n14628,
    n14630, n14631, n14632, n14633, n14634, n14635,
    n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647,
    n14648, n14649, n14650, n14651, n14652, n14653,
    n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665,
    n14666, n14667, n14668, n14669, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683,
    n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701,
    n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719,
    n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731,
    n14732, n14733, n14734, n14735, n14736, n14737,
    n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749,
    n14750, n14751, n14752, n14753, n14754, n14755,
    n14756, n14757, n14758, n14759, n14760, n14761,
    n14762, n14763, n14764, n14765, n14766, n14767,
    n14768, n14769, n14770, n14771, n14772, n14773,
    n14774, n14775, n14776, n14777, n14778, n14779,
    n14780, n14781, n14782, n14783, n14784, n14785,
    n14786, n14787, n14788, n14789, n14790, n14791,
    n14792, n14793, n14794, n14795, n14796, n14797,
    n14798, n14799, n14800, n14801, n14802, n14803,
    n14804, n14805, n14806, n14807, n14808, n14809,
    n14810, n14811, n14812, n14813, n14814, n14815,
    n14816, n14817, n14818, n14819, n14820, n14821,
    n14822, n14823, n14824, n14825, n14826, n14827,
    n14828, n14829, n14830, n14831, n14832, n14833,
    n14834, n14835, n14836, n14837, n14838, n14839,
    n14840, n14841, n14842, n14843, n14844, n14845,
    n14846, n14847, n14848, n14849, n14850, n14851,
    n14852, n14853, n14854, n14855, n14856, n14857,
    n14858, n14859, n14860, n14861, n14862, n14863,
    n14864, n14865, n14866, n14867, n14868, n14869,
    n14870, n14871, n14872, n14873, n14874, n14875,
    n14876, n14877, n14878, n14879, n14880, n14881,
    n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14890, n14891, n14892, n14893,
    n14894, n14895, n14896, n14897, n14898, n14899,
    n14900, n14901, n14902, n14903, n14904, n14905,
    n14906, n14907, n14908, n14909, n14910, n14911,
    n14912, n14913, n14914, n14915, n14916, n14917,
    n14918, n14919, n14920, n14921, n14922, n14923,
    n14924, n14925, n14926, n14927, n14928, n14929,
    n14930, n14931, n14932, n14933, n14934, n14935,
    n14936, n14937, n14938, n14939, n14940, n14941,
    n14942, n14943, n14944, n14945, n14946, n14947,
    n14948, n14949, n14950, n14951, n14952, n14953,
    n14954, n14955, n14956, n14957, n14958, n14959,
    n14960, n14961, n14962, n14963, n14964, n14965,
    n14966, n14967, n14968, n14969, n14970, n14971,
    n14972, n14973, n14974, n14975, n14976, n14977,
    n14978, n14979, n14980, n14981, n14982, n14983,
    n14984, n14985, n14986, n14987, n14988, n14989,
    n14990, n14991, n14992, n14993, n14994, n14995,
    n14996, n14997, n14998, n14999, n15000, n15001,
    n15002, n15003, n15004, n15005, n15006, n15007,
    n15008, n15009, n15010, n15011, n15012, n15013,
    n15014, n15015, n15016, n15017, n15018, n15019,
    n15020, n15021, n15022, n15023, n15024, n15025,
    n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037,
    n15038, n15039, n15040, n15041, n15042, n15043,
    n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055,
    n15056, n15057, n15058, n15059, n15060, n15061,
    n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073,
    n15074, n15075, n15076, n15077, n15078, n15079,
    n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091,
    n15092, n15093, n15094, n15095, n15096, n15097,
    n15098, n15099, n15100, n15101, n15102, n15103,
    n15104, n15105, n15106, n15107, n15108, n15109,
    n15110, n15111, n15112, n15113, n15114, n15115,
    n15116, n15117, n15118, n15119, n15120, n15121,
    n15122, n15123, n15124, n15125, n15126, n15127,
    n15128, n15129, n15130, n15131, n15132, n15133,
    n15134, n15135, n15136, n15137, n15138, n15139,
    n15140, n15141, n15142, n15143, n15144, n15145,
    n15146, n15147, n15148, n15149, n15150, n15151,
    n15152, n15153, n15154, n15155, n15156, n15157,
    n15158, n15159, n15160, n15161, n15162, n15163,
    n15164, n15165, n15166, n15167, n15168, n15169,
    n15170, n15171, n15172, n15173, n15174, n15175,
    n15176, n15177, n15178, n15179, n15180, n15181,
    n15182, n15183, n15184, n15185, n15186, n15187,
    n15188, n15189, n15190, n15191, n15192, n15193,
    n15194, n15195, n15196, n15197, n15198, n15199,
    n15200, n15201, n15202, n15203, n15204, n15205,
    n15206, n15207, n15208, n15209, n15210, n15211,
    n15212, n15213, n15214, n15215, n15216, n15217,
    n15218, n15219, n15220, n15221, n15222, n15223,
    n15224, n15225, n15226, n15227, n15228, n15229,
    n15230, n15231, n15232, n15233, n15234, n15235,
    n15236, n15237, n15238, n15239, n15240, n15241,
    n15242, n15243, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253,
    n15254, n15255, n15256, n15257, n15258, n15259,
    n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271,
    n15272, n15273, n15274, n15276, n15277, n15278,
    n15279, n15280, n15281, n15282, n15283, n15284,
    n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302,
    n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314,
    n15315, n15316, n15317, n15318, n15319, n15320,
    n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338,
    n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15355, n15356,
    n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368,
    n15369, n15370, n15371, n15372, n15373, n15374,
    n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392,
    n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404,
    n15405, n15406, n15407, n15408, n15409, n15410,
    n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422,
    n15423, n15424, n15425, n15426, n15427, n15428,
    n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440,
    n15441, n15442, n15443, n15444, n15445, n15446,
    n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458,
    n15459, n15460, n15461, n15462, n15463, n15464,
    n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476,
    n15477, n15478, n15479, n15480, n15481, n15482,
    n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494,
    n15495, n15496, n15497, n15498, n15499, n15500,
    n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512,
    n15513, n15514, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530,
    n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15768, n15769, n15770,
    n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782,
    n15783, n15784, n15785, n15786, n15787, n15788,
    n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800,
    n15801, n15802, n15803, n15804, n15805, n15806,
    n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824,
    n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854,
    n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15871, n15872, n15873,
    n15874, n15875, n15876, n15877, n15878, n15879,
    n15880, n15881, n15882, n15883, n15884, n15885,
    n15886, n15887, n15888, n15889, n15890, n15891,
    n15892, n15893, n15894, n15895, n15896, n15897,
    n15898, n15899, n15900, n15901, n15902, n15903,
    n15904, n15905, n15906, n15907, n15908, n15909,
    n15910, n15911, n15912, n15913, n15914, n15915,
    n15916, n15917, n15918, n15919, n15920, n15921,
    n15922, n15923, n15924, n15925, n15926, n15927,
    n15928, n15929, n15930, n15931, n15932, n15933,
    n15934, n15935, n15936, n15937, n15938, n15939,
    n15940, n15941, n15942, n15943, n15944, n15945,
    n15946, n15947, n15948, n15949, n15950, n15951,
    n15952, n15953, n15954, n15955, n15956, n15957,
    n15958, n15959, n15960, n15961, n15962, n15963,
    n15964, n15965, n15966, n15967, n15968, n15969,
    n15970, n15971, n15972, n15973, n15974, n15975,
    n15976, n15977, n15978, n15979, n15980, n15981,
    n15982, n15983, n15984, n15985, n15986, n15987,
    n15988, n15989, n15990, n15991, n15992, n15993,
    n15994, n15995, n15996, n15997, n15998, n15999,
    n16000, n16001, n16002, n16003, n16004, n16005,
    n16006, n16007, n16008, n16009, n16010, n16011,
    n16012, n16013, n16014, n16015, n16016, n16017,
    n16018, n16019, n16020, n16021, n16022, n16023,
    n16024, n16025, n16026, n16027, n16028, n16029,
    n16030, n16031, n16032, n16033, n16034, n16035,
    n16036, n16037, n16038, n16039, n16040, n16041,
    n16042, n16043, n16044, n16045, n16046, n16047,
    n16048, n16049, n16050, n16051, n16052, n16053,
    n16054, n16055, n16056, n16057, n16058, n16059,
    n16060, n16061, n16062, n16063, n16064, n16065,
    n16066, n16067, n16068, n16069, n16070, n16071,
    n16072, n16073, n16074, n16075, n16076, n16077,
    n16078, n16079, n16080, n16081, n16082, n16083,
    n16084, n16085, n16086, n16087, n16088, n16089,
    n16090, n16091, n16092, n16093, n16094, n16095,
    n16096, n16097, n16098, n16099, n16100, n16101,
    n16102, n16103, n16104, n16105, n16106, n16107,
    n16108, n16109, n16110, n16111, n16112, n16113,
    n16114, n16115, n16116, n16117, n16118, n16119,
    n16120, n16121, n16122, n16123, n16124, n16125,
    n16126, n16127, n16128, n16129, n16130, n16131,
    n16132, n16133, n16134, n16135, n16136, n16137,
    n16138, n16139, n16140, n16141, n16142, n16143,
    n16144, n16145, n16146, n16147, n16148, n16149,
    n16150, n16151, n16152, n16153, n16154, n16155,
    n16156, n16157, n16158, n16159, n16160, n16161,
    n16162, n16163, n16164, n16165, n16166, n16167,
    n16168, n16169, n16170, n16171, n16172, n16173,
    n16174, n16175, n16176, n16177, n16178, n16179,
    n16180, n16181, n16182, n16183, n16184, n16185,
    n16186, n16187, n16188, n16189, n16190, n16191,
    n16192, n16193, n16194, n16195, n16196, n16197,
    n16198, n16199, n16200, n16201, n16202, n16203,
    n16204, n16205, n16206, n16207, n16208, n16209,
    n16210, n16211, n16212, n16213, n16214, n16215,
    n16216, n16217, n16218, n16219, n16220, n16221,
    n16222, n16223, n16224, n16225, n16226, n16227,
    n16228, n16229, n16230, n16231, n16232, n16233,
    n16234, n16235, n16236, n16237, n16238, n16239,
    n16240, n16241, n16242, n16243, n16244, n16245,
    n16246, n16247, n16248, n16249, n16250, n16251,
    n16252, n16253, n16254, n16255, n16256, n16257,
    n16258, n16259, n16260, n16261, n16262, n16263,
    n16264, n16265, n16266, n16267, n16268, n16269,
    n16270, n16271, n16272, n16273, n16274, n16275,
    n16276, n16277, n16278, n16279, n16280, n16281,
    n16282, n16283, n16284, n16285, n16286, n16287,
    n16288, n16289, n16290, n16291, n16292, n16293,
    n16294, n16295, n16296, n16297, n16298, n16299,
    n16300, n16301, n16302, n16303, n16304, n16305,
    n16306, n16307, n16308, n16309, n16310, n16311,
    n16312, n16313, n16314, n16315, n16316, n16317,
    n16318, n16319, n16320, n16321, n16322, n16323,
    n16324, n16325, n16326, n16327, n16328, n16329,
    n16330, n16331, n16332, n16333, n16334, n16335,
    n16336, n16337, n16338, n16339, n16340, n16341,
    n16342, n16343, n16344, n16345, n16346, n16347,
    n16348, n16349, n16350, n16351, n16352, n16353,
    n16354, n16355, n16356, n16357, n16358, n16359,
    n16360, n16361, n16362, n16363, n16364, n16365,
    n16366, n16367, n16368, n16369, n16370, n16371,
    n16372, n16373, n16374, n16375, n16376, n16377,
    n16378, n16379, n16380, n16381, n16382, n16383,
    n16384, n16385, n16386, n16387, n16388, n16389,
    n16390, n16391, n16392, n16393, n16394, n16395,
    n16396, n16397, n16398, n16399, n16400, n16401,
    n16402, n16403, n16404, n16405, n16406, n16407,
    n16408, n16409, n16410, n16411, n16412, n16413,
    n16414, n16415, n16416, n16417, n16418, n16419,
    n16420, n16421, n16422, n16423, n16424, n16425,
    n16426, n16427, n16428, n16429, n16430, n16431,
    n16432, n16433, n16434, n16435, n16436, n16437,
    n16438, n16439, n16440, n16441, n16442, n16443,
    n16444, n16445, n16446, n16447, n16448, n16449,
    n16450, n16451, n16452, n16453, n16454, n16455,
    n16456, n16457, n16458, n16459, n16460, n16461,
    n16462, n16463, n16464, n16465, n16466, n16467,
    n16468, n16469, n16470, n16471, n16472, n16473,
    n16474, n16475, n16476, n16477, n16478, n16479,
    n16480, n16481, n16482, n16483, n16484, n16485,
    n16486, n16487, n16488, n16489, n16490, n16491,
    n16492, n16493, n16494, n16495, n16496, n16497,
    n16498, n16499, n16500, n16501, n16502, n16503,
    n16504, n16505, n16506, n16507, n16508, n16509,
    n16510, n16511, n16512, n16513, n16514, n16515,
    n16516, n16517, n16518, n16519, n16520, n16521,
    n16522, n16523, n16524, n16525, n16526, n16527,
    n16528, n16529, n16530, n16531, n16532, n16533,
    n16534, n16535, n16536, n16537, n16538, n16539,
    n16540, n16542, n16543, n16544, n16545, n16546,
    n16547, n16548, n16549, n16550, n16551, n16552,
    n16553, n16554, n16555, n16556, n16557, n16558,
    n16559, n16560, n16561, n16562, n16563, n16564,
    n16565, n16566, n16567, n16568, n16569, n16570,
    n16571, n16572, n16573, n16574, n16575, n16576,
    n16577, n16578, n16579, n16580, n16581, n16582,
    n16583, n16584, n16585, n16586, n16587, n16588,
    n16589, n16590, n16591, n16592, n16593, n16594,
    n16595, n16596, n16597, n16598, n16599, n16600,
    n16601, n16602, n16603, n16604, n16605, n16606,
    n16607, n16608, n16609, n16610, n16611, n16612,
    n16613, n16614, n16615, n16616, n16617, n16618,
    n16619, n16620, n16621, n16622, n16623, n16624,
    n16625, n16626, n16627, n16628, n16629, n16630,
    n16631, n16632, n16633, n16634, n16635, n16636,
    n16637, n16638, n16639, n16640, n16641, n16642,
    n16643, n16644, n16645, n16646, n16647, n16648,
    n16649, n16650, n16651, n16652, n16653, n16654,
    n16655, n16656, n16657, n16658, n16659, n16660,
    n16661, n16662, n16663, n16664, n16665, n16666,
    n16667, n16668, n16669, n16670, n16671, n16672,
    n16673, n16674, n16675, n16676, n16677, n16678,
    n16679, n16680, n16681, n16682, n16683, n16684,
    n16685, n16686, n16687, n16688, n16689, n16690,
    n16691, n16692, n16693, n16694, n16695, n16696,
    n16697, n16698, n16699, n16700, n16701, n16702,
    n16703, n16704, n16705, n16706, n16707, n16708,
    n16709, n16710, n16711, n16712, n16713, n16714,
    n16715, n16716, n16717, n16718, n16719, n16720,
    n16721, n16722, n16723, n16724, n16725, n16726,
    n16727, n16728, n16729, n16730, n16731, n16732,
    n16733, n16734, n16735, n16736, n16737, n16738,
    n16739, n16740, n16741, n16742, n16743, n16744,
    n16745, n16746, n16747, n16748, n16749, n16750,
    n16751, n16752, n16753, n16754, n16755, n16756,
    n16757, n16758, n16759, n16760, n16761, n16762,
    n16763, n16764, n16765, n16766, n16767, n16768,
    n16769, n16770, n16771, n16772, n16773, n16774,
    n16775, n16776, n16777, n16778, n16779, n16780,
    n16781, n16782, n16783, n16784, n16785, n16786,
    n16787, n16788, n16789, n16790, n16791, n16792,
    n16793, n16794, n16795, n16796, n16797, n16798,
    n16799, n16800, n16801, n16802, n16803, n16804,
    n16805, n16806, n16807, n16808, n16809, n16810,
    n16811, n16812, n16813, n16814, n16815, n16816,
    n16817, n16818, n16819, n16820, n16821, n16822,
    n16823, n16824, n16825, n16826, n16827, n16828,
    n16829, n16830, n16831, n16832, n16833, n16834,
    n16835, n16836, n16837, n16838, n16839, n16840,
    n16841, n16842, n16843, n16844, n16845, n16846,
    n16847, n16848, n16849, n16850, n16851, n16852,
    n16853, n16854, n16855, n16856, n16857, n16858,
    n16859, n16860, n16861, n16862, n16863, n16864,
    n16865, n16866, n16867, n16868, n16869, n16870,
    n16871, n16872, n16873, n16874, n16875, n16876,
    n16877, n16878, n16879, n16880, n16881, n16882,
    n16883, n16884, n16885, n16886, n16887, n16888,
    n16889, n16890, n16891, n16892, n16893, n16894,
    n16895, n16896, n16897, n16898, n16899, n16900,
    n16901, n16902, n16903, n16904, n16905, n16906,
    n16907, n16908, n16909, n16910, n16911, n16912,
    n16913, n16914, n16915, n16916, n16917, n16918,
    n16919, n16920, n16921, n16922, n16923, n16924,
    n16925, n16926, n16927, n16928, n16929, n16930,
    n16931, n16932, n16933, n16934, n16935, n16936,
    n16937, n16938, n16939, n16940, n16941, n16942,
    n16943, n16944, n16945, n16946, n16947, n16948,
    n16949, n16950, n16951, n16952, n16953, n16954,
    n16955, n16956, n16957, n16958, n16959, n16960,
    n16961, n16962, n16963, n16964, n16965, n16966,
    n16967, n16968, n16969, n16970, n16971, n16972,
    n16973, n16974, n16975, n16976, n16977, n16978,
    n16979, n16980, n16981, n16982, n16983, n16984,
    n16985, n16986, n16987, n16988, n16989, n16990,
    n16991, n16992, n16993, n16994, n16995, n16996,
    n16997, n16998, n16999, n17000, n17001, n17002,
    n17003, n17004, n17005, n17006, n17007, n17008,
    n17009, n17010, n17011, n17012, n17013, n17014,
    n17015, n17016, n17017, n17018, n17019, n17020,
    n17021, n17022, n17023, n17024, n17025, n17026,
    n17027, n17028, n17029, n17030, n17031, n17032,
    n17033, n17034, n17035, n17036, n17037, n17038,
    n17039, n17040, n17041, n17042, n17043, n17044,
    n17045, n17046, n17047, n17048, n17049, n17050,
    n17051, n17052, n17053, n17054, n17055, n17056,
    n17057, n17058, n17059, n17060, n17061, n17062,
    n17063, n17064, n17065, n17066, n17067, n17068,
    n17069, n17070, n17071, n17072, n17073, n17074,
    n17075, n17076, n17077, n17078, n17079, n17080,
    n17081, n17082, n17083, n17084, n17085, n17086,
    n17087, n17088, n17089, n17090, n17091, n17092,
    n17093, n17094, n17095, n17096, n17097, n17098,
    n17099, n17100, n17101, n17102, n17103, n17104,
    n17105, n17106, n17107, n17108, n17109, n17110,
    n17111, n17112, n17113, n17114, n17115, n17116,
    n17117, n17118, n17119, n17120, n17121, n17122,
    n17123, n17124, n17125, n17126, n17127, n17128,
    n17129, n17130, n17131, n17132, n17133, n17134,
    n17135, n17137, n17138, n17139, n17140, n17141,
    n17142, n17143, n17144, n17145, n17146, n17147,
    n17148, n17149, n17150, n17151, n17152, n17153,
    n17154, n17155, n17156, n17157, n17158, n17159,
    n17160, n17161, n17162, n17163, n17164, n17165,
    n17166, n17167, n17168, n17169, n17170, n17171,
    n17172, n17173, n17174, n17175, n17176, n17177,
    n17178, n17179, n17180, n17181, n17182, n17183,
    n17184, n17185, n17186, n17187, n17188, n17189,
    n17190, n17191, n17192, n17193, n17194, n17195,
    n17196, n17197, n17198, n17199, n17200, n17201,
    n17202, n17203, n17204, n17205, n17206, n17207,
    n17208, n17209, n17210, n17211, n17212, n17213,
    n17214, n17215, n17216, n17217, n17218, n17219,
    n17220, n17221, n17222, n17223, n17224, n17225,
    n17226, n17227, n17228, n17229, n17230, n17231,
    n17232, n17233, n17234, n17235, n17236, n17237,
    n17238, n17239, n17240, n17241, n17242, n17243,
    n17244, n17245, n17246, n17247, n17248, n17249,
    n17250, n17251, n17252, n17253, n17254, n17255,
    n17256, n17257, n17258, n17259, n17260, n17261,
    n17262, n17263, n17264, n17265, n17266, n17267,
    n17268, n17269, n17270, n17271, n17272, n17273,
    n17274, n17275, n17276, n17277, n17278, n17279,
    n17280, n17281, n17282, n17283, n17284, n17285,
    n17286, n17287, n17288, n17289, n17290, n17291,
    n17292, n17293, n17294, n17295, n17296, n17297,
    n17298, n17299, n17300, n17301, n17302, n17303,
    n17304, n17305, n17306, n17307, n17308, n17309,
    n17310, n17311, n17312, n17313, n17314, n17315,
    n17316, n17317, n17318, n17319, n17320, n17321,
    n17322, n17323, n17324, n17325, n17326, n17327,
    n17328, n17329, n17330, n17331, n17332, n17333,
    n17334, n17335, n17336, n17337, n17338, n17339,
    n17340, n17341, n17342, n17343, n17344, n17345,
    n17346, n17347, n17348, n17349, n17350, n17351,
    n17352, n17353, n17354, n17355, n17356, n17357,
    n17358, n17359, n17360, n17361, n17362, n17363,
    n17364, n17365, n17366, n17367, n17368, n17369,
    n17370, n17371, n17372, n17373, n17374, n17375,
    n17376, n17377, n17378, n17379, n17380, n17381,
    n17382, n17383, n17384, n17385, n17386, n17387,
    n17388, n17389, n17390, n17391, n17392, n17393,
    n17394, n17395, n17396, n17397, n17398, n17399,
    n17400, n17401, n17402, n17403, n17404, n17405,
    n17406, n17407, n17408, n17409, n17410, n17411,
    n17412, n17413, n17414, n17415, n17416, n17417,
    n17418, n17419, n17420, n17421, n17422, n17423,
    n17424, n17425, n17426, n17427, n17428, n17429,
    n17430, n17431, n17432, n17433, n17434, n17435,
    n17436, n17437, n17438, n17439, n17440, n17441,
    n17442, n17443, n17444, n17445, n17446, n17447,
    n17448, n17449, n17450, n17451, n17452, n17453,
    n17454, n17455, n17456, n17457, n17458, n17459,
    n17460, n17461, n17462, n17463, n17464, n17465,
    n17466, n17467, n17468, n17469, n17470, n17471,
    n17472, n17473, n17474, n17475, n17476, n17477,
    n17478, n17479, n17480, n17481, n17482, n17483,
    n17484, n17485, n17486, n17487, n17488, n17489,
    n17490, n17491, n17492, n17493, n17494, n17495,
    n17496, n17497, n17498, n17499, n17500, n17501,
    n17502, n17503, n17504, n17505, n17506, n17507,
    n17508, n17509, n17510, n17511, n17512, n17513,
    n17514, n17515, n17516, n17517, n17518, n17519,
    n17520, n17521, n17522, n17523, n17524, n17525,
    n17526, n17527, n17528, n17529, n17530, n17531,
    n17532, n17533, n17534, n17535, n17536, n17537,
    n17538, n17539, n17540, n17541, n17542, n17543,
    n17544, n17545, n17546, n17547, n17548, n17549,
    n17550, n17551, n17552, n17553, n17554, n17555,
    n17556, n17557, n17558, n17559, n17560, n17561,
    n17562, n17563, n17564, n17565, n17566, n17567,
    n17568, n17569, n17570, n17571, n17572, n17573,
    n17574, n17575, n17576, n17577, n17578, n17579,
    n17580, n17581, n17582, n17583, n17584, n17585,
    n17586, n17587, n17588, n17589, n17590, n17591,
    n17592, n17593, n17594, n17595, n17596, n17597,
    n17598, n17599, n17600, n17601, n17602, n17603,
    n17604, n17605, n17606, n17607, n17608, n17609,
    n17610, n17611, n17612, n17613, n17614, n17615,
    n17616, n17617, n17618, n17619, n17620, n17621,
    n17622, n17623, n17624, n17625, n17626, n17627,
    n17628, n17629, n17630, n17631, n17632, n17633,
    n17634, n17635, n17636, n17637, n17638, n17639,
    n17640, n17641, n17642, n17643, n17644, n17645,
    n17646, n17647, n17648, n17649, n17650, n17651,
    n17652, n17653, n17654, n17655, n17656, n17657,
    n17658, n17659, n17660, n17661, n17662, n17663,
    n17664, n17665, n17666, n17667, n17668, n17669,
    n17670, n17671, n17672, n17673, n17674, n17675,
    n17676, n17677, n17678, n17679, n17680, n17681,
    n17682, n17683, n17684, n17685, n17686, n17687,
    n17688, n17689, n17690, n17691, n17692, n17693,
    n17694, n17695, n17696, n17697, n17698, n17699,
    n17700, n17701, n17702, n17703, n17704, n17705,
    n17706, n17707, n17708, n17709, n17710, n17711,
    n17712, n17713, n17714, n17715, n17716, n17717,
    n17718, n17719, n17720, n17721, n17722, n17723,
    n17724, n17725, n17726, n17727, n17728, n17729,
    n17730, n17732, n17733, n17734, n17735, n17736,
    n17737, n17738, n17739, n17740, n17741, n17742,
    n17743, n17744, n17745, n17746, n17747, n17748,
    n17749, n17750, n17751, n17752, n17753, n17754,
    n17755, n17756, n17757, n17758, n17759, n17760,
    n17761, n17762, n17763, n17764, n17765, n17766,
    n17767, n17768, n17769, n17770, n17771, n17772,
    n17773, n17774, n17775, n17776, n17777, n17778,
    n17779, n17780, n17781, n17782, n17783, n17784,
    n17785, n17786, n17787, n17788, n17789, n17790,
    n17791, n17792, n17793, n17794, n17795, n17796,
    n17797, n17798, n17799, n17800, n17801, n17802,
    n17803, n17804, n17805, n17806, n17807, n17808,
    n17809, n17810, n17811, n17812, n17813, n17814,
    n17815, n17816, n17817, n17818, n17819, n17820,
    n17821, n17822, n17823, n17824, n17825, n17826,
    n17827, n17828, n17829, n17830, n17831, n17832,
    n17833, n17834, n17835, n17836, n17837, n17838,
    n17839, n17840, n17841, n17842, n17843, n17844,
    n17845, n17846, n17847, n17848, n17849, n17850,
    n17851, n17852, n17853, n17854, n17855, n17856,
    n17857, n17858, n17859, n17860, n17861, n17862,
    n17863, n17864, n17865, n17866, n17867, n17868,
    n17869, n17870, n17871, n17872, n17873, n17874,
    n17875, n17876, n17877, n17878, n17879, n17880,
    n17881, n17882, n17883, n17884, n17885, n17886,
    n17887, n17888, n17889, n17890, n17891, n17892,
    n17893, n17894, n17895, n17896, n17897, n17898,
    n17899, n17900, n17901, n17902, n17903, n17904,
    n17905, n17906, n17907, n17908, n17909, n17910,
    n17911, n17912, n17913, n17914, n17915, n17916,
    n17917, n17918, n17919, n17920, n17921, n17922,
    n17923, n17924, n17925, n17926, n17927, n17928,
    n17929, n17930, n17931, n17932, n17933, n17934,
    n17935, n17936, n17937, n17938, n17939, n17940,
    n17941, n17942, n17943, n17944, n17945, n17946,
    n17947, n17948, n17949, n17950, n17951, n17952,
    n17953, n17954, n17955, n17956, n17957, n17958,
    n17959, n17960, n17961, n17962, n17963, n17964,
    n17965, n17966, n17967, n17968, n17969, n17970,
    n17971, n17972, n17973, n17974, n17975, n17976,
    n17977, n17978, n17979, n17980, n17981, n17982,
    n17983, n17984, n17985, n17986, n17987, n17988,
    n17989, n17990, n17991, n17992, n17993, n17994,
    n17995, n17996, n17997, n17998, n17999, n18000,
    n18001, n18002, n18003, n18004, n18005, n18006,
    n18007, n18008, n18009, n18010, n18011, n18012,
    n18013, n18014, n18015, n18016, n18017, n18018,
    n18019, n18020, n18021, n18022, n18023, n18024,
    n18025, n18026, n18027, n18028, n18029, n18030,
    n18031, n18032, n18033, n18034, n18035, n18036,
    n18037, n18038, n18039, n18040, n18041, n18042,
    n18043, n18044, n18045, n18046, n18047, n18048,
    n18049, n18050, n18051, n18052, n18053, n18054,
    n18055, n18056, n18057, n18058, n18059, n18060,
    n18061, n18062, n18063, n18064, n18065, n18066,
    n18067, n18068, n18069, n18070, n18071, n18072,
    n18073, n18074, n18075, n18076, n18077, n18078,
    n18079, n18080, n18081, n18082, n18083, n18084,
    n18085, n18086, n18087, n18088, n18089, n18090,
    n18091, n18092, n18093, n18094, n18095, n18096,
    n18097, n18098, n18099, n18100, n18101, n18102,
    n18103, n18104, n18105, n18106, n18107, n18108,
    n18109, n18110, n18111, n18112, n18113, n18114,
    n18115, n18116, n18117, n18118, n18119, n18120,
    n18121, n18122, n18123, n18124, n18125, n18126,
    n18127, n18128, n18129, n18130, n18131, n18132,
    n18133, n18134, n18135, n18136, n18137, n18138,
    n18139, n18140, n18141, n18142, n18143, n18144,
    n18145, n18146, n18147, n18148, n18149, n18150,
    n18151, n18152, n18153, n18154, n18155, n18156,
    n18157, n18158, n18159, n18160, n18161, n18162,
    n18163, n18164, n18165, n18166, n18167, n18168,
    n18169, n18170, n18171, n18172, n18173, n18174,
    n18175, n18176, n18177, n18178, n18179, n18180,
    n18181, n18182, n18183, n18184, n18185, n18186,
    n18187, n18188, n18189, n18190, n18191, n18192,
    n18193, n18194, n18195, n18196, n18197, n18198,
    n18199, n18200, n18201, n18202, n18203, n18204,
    n18205, n18206, n18207, n18208, n18209, n18210,
    n18211, n18212, n18213, n18214, n18215, n18216,
    n18217, n18218, n18219, n18220, n18221, n18222,
    n18223, n18224, n18225, n18226, n18227, n18228,
    n18229, n18230, n18231, n18232, n18233, n18234,
    n18235, n18236, n18237, n18238, n18239, n18240,
    n18241, n18242, n18243, n18244, n18245, n18246,
    n18247, n18248, n18249, n18250, n18251, n18252,
    n18253, n18254, n18255, n18256, n18257, n18258,
    n18259, n18260, n18261, n18262, n18263, n18264,
    n18265, n18266, n18267, n18268, n18269, n18270,
    n18271, n18272, n18273, n18274, n18275, n18276,
    n18277, n18278, n18279, n18280, n18281, n18282,
    n18283, n18284, n18285, n18286, n18287, n18288,
    n18289, n18290, n18291, n18292, n18293, n18294,
    n18295, n18296, n18297, n18298, n18299, n18300,
    n18301, n18302, n18303, n18304, n18305, n18306,
    n18307, n18308, n18309, n18310, n18311, n18312,
    n18313, n18314, n18315, n18316, n18317, n18318,
    n18319, n18320, n18321, n18322, n18323, n18325,
    n18326, n18327, n18328, n18329, n18330, n18331,
    n18332, n18333, n18334, n18335, n18336, n18337,
    n18338, n18339, n18340, n18341, n18342, n18343,
    n18344, n18345, n18346, n18347, n18348, n18349,
    n18350, n18351, n18352, n18353, n18354, n18355,
    n18356, n18357, n18358, n18359, n18360, n18361,
    n18362, n18363, n18364, n18365, n18366, n18367,
    n18368, n18369, n18370, n18371, n18372, n18373,
    n18374, n18375, n18376, n18377, n18378, n18379,
    n18380, n18381, n18382, n18383, n18384, n18385,
    n18386, n18387, n18388, n18389, n18390, n18391,
    n18392, n18393, n18394, n18395, n18396, n18397,
    n18398, n18399, n18400, n18401, n18402, n18403,
    n18404, n18405, n18406, n18407, n18408, n18409,
    n18410, n18411, n18412, n18413, n18414, n18415,
    n18416, n18417, n18418, n18419, n18420, n18421,
    n18422, n18423, n18424, n18425, n18426, n18427,
    n18428, n18429, n18430, n18431, n18432, n18433,
    n18434, n18435, n18436, n18437, n18438, n18439,
    n18440, n18441, n18442, n18443, n18444, n18445,
    n18446, n18447, n18448, n18449, n18450, n18451,
    n18452, n18453, n18454, n18455, n18456, n18457,
    n18458, n18459, n18460, n18461, n18462, n18463,
    n18464, n18465, n18466, n18467, n18468, n18469,
    n18470, n18471, n18472, n18473, n18474, n18475,
    n18476, n18477, n18478, n18479, n18480, n18481,
    n18482, n18483, n18484, n18485, n18486, n18487,
    n18488, n18489, n18490, n18491, n18492, n18493,
    n18494, n18495, n18496, n18497, n18498, n18499,
    n18500, n18501, n18502, n18503, n18504, n18505,
    n18506, n18507, n18508, n18509, n18510, n18511,
    n18512, n18513, n18514, n18515, n18516, n18517,
    n18518, n18519, n18520, n18521, n18522, n18523,
    n18524, n18525, n18526, n18527, n18528, n18529,
    n18530, n18531, n18532, n18533, n18534, n18535,
    n18536, n18537, n18538, n18539, n18540, n18541,
    n18542, n18543, n18544, n18545, n18546, n18547,
    n18548, n18549, n18550, n18551, n18552, n18553,
    n18554, n18555, n18556, n18557, n18558, n18559,
    n18560, n18561, n18562, n18563, n18564, n18565,
    n18566, n18567, n18568, n18569, n18570, n18571,
    n18572, n18573, n18574, n18575, n18576, n18577,
    n18578, n18579, n18580, n18581, n18582, n18583,
    n18584, n18585, n18586, n18587, n18588, n18589,
    n18590, n18591, n18592, n18593, n18594, n18595,
    n18596, n18597, n18598, n18599, n18600, n18601,
    n18602, n18603, n18604, n18605, n18606, n18607,
    n18608, n18609, n18610, n18611, n18612, n18613,
    n18614, n18615, n18616, n18617, n18618, n18619,
    n18620, n18621, n18622, n18623, n18624, n18625,
    n18626, n18627, n18628, n18629, n18630, n18631,
    n18632, n18633, n18634, n18635, n18636, n18637,
    n18638, n18639, n18640, n18641, n18642, n18643,
    n18644, n18645, n18646, n18647, n18648, n18649,
    n18650, n18651, n18652, n18653, n18654, n18655,
    n18656, n18657, n18658, n18659, n18660, n18661,
    n18662, n18663, n18664, n18665, n18666, n18667,
    n18668, n18669, n18670, n18671, n18672, n18673,
    n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685,
    n18686, n18687, n18688, n18689, n18690, n18691,
    n18692, n18693, n18694, n18695, n18696, n18697,
    n18698, n18699, n18700, n18701, n18702, n18703,
    n18704, n18705, n18706, n18707, n18708, n18709,
    n18710, n18711, n18712, n18713, n18714, n18715,
    n18716, n18717, n18718, n18719, n18720, n18721,
    n18722, n18723, n18724, n18725, n18726, n18727,
    n18728, n18729, n18730, n18731, n18732, n18733,
    n18734, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18742, n18743, n18744, n18745,
    n18746, n18747, n18748, n18749, n18750, n18751,
    n18752, n18753, n18754, n18755, n18756, n18757,
    n18758, n18759, n18760, n18761, n18762, n18763,
    n18764, n18765, n18766, n18767, n18768, n18769,
    n18770, n18771, n18772, n18773, n18774, n18775,
    n18776, n18777, n18778, n18779, n18780, n18781,
    n18782, n18783, n18784, n18785, n18786, n18787,
    n18788, n18789, n18790, n18791, n18792, n18793,
    n18794, n18795, n18796, n18797, n18798, n18799,
    n18800, n18801, n18802, n18803, n18804, n18805,
    n18806, n18807, n18808, n18809, n18810, n18811,
    n18812, n18813, n18814, n18815, n18816, n18817,
    n18818, n18819, n18820, n18821, n18822, n18823,
    n18824, n18825, n18826, n18827, n18828, n18829,
    n18830, n18831, n18832, n18833, n18834, n18835,
    n18836, n18837, n18838, n18839, n18840, n18841,
    n18842, n18843, n18844, n18845, n18846, n18847,
    n18848, n18849, n18850, n18851, n18852, n18853,
    n18854, n18855, n18856, n18857, n18858, n18859,
    n18860, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18871,
    n18872, n18873, n18874, n18875, n18876, n18877,
    n18878, n18879, n18880, n18881, n18882, n18883,
    n18884, n18885, n18886, n18887, n18888, n18889,
    n18890, n18891, n18892, n18893, n18894, n18895,
    n18896, n18897, n18898, n18899, n18900, n18901,
    n18902, n18903, n18904, n18905, n18906, n18907,
    n18908, n18909, n18910, n18911, n18912, n18913,
    n18914, n18915, n18916, n18918, n18919, n18920,
    n18921, n18922, n18923, n18924, n18925, n18926,
    n18927, n18928, n18929, n18930, n18931, n18932,
    n18933, n18934, n18935, n18936, n18937, n18938,
    n18939, n18940, n18941, n18942, n18943, n18944,
    n18945, n18946, n18947, n18948, n18949, n18950,
    n18951, n18952, n18953, n18954, n18955, n18956,
    n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968,
    n18969, n18970, n18971, n18972, n18973, n18974,
    n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986,
    n18987, n18988, n18989, n18990, n18991, n18992,
    n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004,
    n19005, n19006, n19007, n19008, n19009, n19010,
    n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022,
    n19023, n19024, n19025, n19026, n19027, n19028,
    n19029, n19030, n19031, n19032, n19033, n19034,
    n19035, n19036, n19037, n19038, n19039, n19040,
    n19041, n19042, n19043, n19044, n19045, n19046,
    n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058,
    n19059, n19060, n19061, n19062, n19063, n19064,
    n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076,
    n19077, n19078, n19079, n19080, n19081, n19082,
    n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094,
    n19095, n19096, n19097, n19098, n19099, n19100,
    n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112,
    n19113, n19114, n19115, n19116, n19117, n19118,
    n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130,
    n19131, n19132, n19133, n19134, n19135, n19136,
    n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148,
    n19149, n19150, n19151, n19152, n19153, n19154,
    n19155, n19156, n19157, n19158, n19159, n19160,
    n19161, n19162, n19163, n19164, n19165, n19166,
    n19167, n19168, n19169, n19170, n19171, n19172,
    n19173, n19174, n19175, n19176, n19177, n19178,
    n19179, n19180, n19181, n19182, n19183, n19184,
    n19185, n19186, n19187, n19188, n19189, n19190,
    n19191, n19192, n19193, n19194, n19195, n19196,
    n19197, n19198, n19199, n19200, n19201, n19202,
    n19203, n19204, n19205, n19206, n19207, n19208,
    n19209, n19210, n19211, n19212, n19213, n19214,
    n19215, n19216, n19217, n19218, n19219, n19220,
    n19221, n19222, n19223, n19224, n19225, n19226,
    n19227, n19228, n19229, n19230, n19231, n19232,
    n19233, n19234, n19235, n19236, n19237, n19238,
    n19239, n19240, n19241, n19242, n19243, n19244,
    n19245, n19246, n19247, n19248, n19249, n19250,
    n19251, n19252, n19253, n19254, n19255, n19256,
    n19257, n19258, n19259, n19260, n19261, n19262,
    n19263, n19264, n19265, n19266, n19267, n19268,
    n19269, n19270, n19271, n19272, n19273, n19274,
    n19275, n19276, n19277, n19278, n19279, n19280,
    n19281, n19282, n19283, n19284, n19285, n19286,
    n19287, n19288, n19289, n19290, n19291, n19292,
    n19293, n19294, n19295, n19296, n19297, n19298,
    n19299, n19300, n19301, n19302, n19303, n19304,
    n19305, n19306, n19307, n19308, n19309, n19310,
    n19311, n19312, n19313, n19314, n19315, n19316,
    n19317, n19318, n19319, n19320, n19321, n19322,
    n19323, n19324, n19325, n19326, n19327, n19328,
    n19329, n19330, n19331, n19332, n19333, n19334,
    n19335, n19336, n19337, n19338, n19339, n19340,
    n19341, n19342, n19343, n19344, n19345, n19346,
    n19347, n19348, n19349, n19350, n19351, n19352,
    n19353, n19354, n19355, n19356, n19357, n19358,
    n19359, n19360, n19361, n19362, n19363, n19364,
    n19365, n19366, n19367, n19368, n19369, n19370,
    n19371, n19372, n19373, n19374, n19375, n19376,
    n19377, n19378, n19379, n19380, n19381, n19382,
    n19383, n19384, n19385, n19386, n19387, n19388,
    n19389, n19390, n19391, n19392, n19393, n19394,
    n19395, n19396, n19397, n19398, n19399, n19400,
    n19401, n19402, n19403, n19404, n19405, n19406,
    n19407, n19408, n19409, n19410, n19411, n19412,
    n19413, n19414, n19415, n19416, n19417, n19418,
    n19419, n19420, n19421, n19422, n19423, n19424,
    n19425, n19426, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19435, n19436,
    n19437, n19438, n19439, n19440, n19441, n19442,
    n19443, n19444, n19445, n19446, n19447, n19448,
    n19449, n19450, n19451, n19452, n19453, n19454,
    n19455, n19456, n19457, n19458, n19459, n19460,
    n19461, n19462, n19463, n19464, n19465, n19466,
    n19467, n19468, n19469, n19470, n19471, n19472,
    n19473, n19474, n19475, n19476, n19477, n19478,
    n19479, n19480, n19481, n19482, n19483, n19484,
    n19485, n19486, n19487, n19488, n19489, n19490,
    n19491, n19492, n19493, n19494, n19495, n19496,
    n19497, n19498, n19499, n19500, n19501, n19502,
    n19503, n19504, n19505, n19506, n19507, n19508,
    n19509, n19511, n19512, n19513, n19514, n19515,
    n19516, n19517, n19518, n19519, n19520, n19521,
    n19522, n19523, n19524, n19525, n19526, n19527,
    n19528, n19529, n19530, n19531, n19532, n19533,
    n19534, n19535, n19536, n19537, n19538, n19539,
    n19540, n19541, n19542, n19543, n19544, n19545,
    n19546, n19547, n19548, n19549, n19550, n19551,
    n19552, n19553, n19554, n19555, n19556, n19557,
    n19558, n19559, n19560, n19561, n19562, n19563,
    n19564, n19565, n19566, n19567, n19568, n19569,
    n19570, n19571, n19572, n19573, n19574, n19575,
    n19576, n19577, n19578, n19579, n19580, n19581,
    n19582, n19583, n19584, n19585, n19586, n19587,
    n19588, n19589, n19590, n19591, n19592, n19593,
    n19594, n19595, n19596, n19597, n19598, n19599,
    n19600, n19601, n19602, n19603, n19604, n19605,
    n19606, n19607, n19608, n19609, n19610, n19611,
    n19612, n19613, n19614, n19615, n19616, n19617,
    n19618, n19619, n19620, n19621, n19622, n19623,
    n19624, n19625, n19626, n19627, n19628, n19629,
    n19630, n19631, n19632, n19633, n19634, n19635,
    n19636, n19637, n19638, n19639, n19640, n19641,
    n19642, n19643, n19644, n19645, n19646, n19647,
    n19648, n19649, n19650, n19651, n19652, n19653,
    n19654, n19655, n19656, n19657, n19658, n19659,
    n19660, n19661, n19662, n19663, n19664, n19665,
    n19666, n19667, n19668, n19669, n19670, n19671,
    n19672, n19673, n19674, n19675, n19676, n19677,
    n19678, n19679, n19680, n19681, n19682, n19683,
    n19684, n19685, n19686, n19687, n19688, n19689,
    n19690, n19691, n19692, n19693, n19694, n19695,
    n19696, n19697, n19698, n19699, n19700, n19701,
    n19702, n19703, n19704, n19705, n19706, n19707,
    n19708, n19709, n19710, n19711, n19712, n19713,
    n19714, n19715, n19716, n19717, n19718, n19719,
    n19720, n19721, n19722, n19723, n19724, n19725,
    n19726, n19727, n19728, n19729, n19730, n19731,
    n19732, n19733, n19734, n19735, n19736, n19737,
    n19738, n19739, n19740, n19741, n19742, n19743,
    n19744, n19745, n19746, n19747, n19748, n19749,
    n19750, n19751, n19752, n19753, n19754, n19755,
    n19756, n19757, n19758, n19759, n19760, n19761,
    n19762, n19763, n19764, n19765, n19766, n19767,
    n19768, n19769, n19770, n19771, n19772, n19773,
    n19774, n19775, n19776, n19777, n19778, n19779,
    n19780, n19781, n19782, n19783, n19784, n19785,
    n19786, n19787, n19788, n19789, n19790, n19791,
    n19792, n19793, n19794, n19795, n19796, n19797,
    n19798, n19799, n19800, n19801, n19802, n19803,
    n19804, n19805, n19806, n19807, n19808, n19809,
    n19810, n19811, n19812, n19813, n19814, n19815,
    n19816, n19817, n19818, n19819, n19820, n19821,
    n19822, n19823, n19824, n19825, n19826, n19827,
    n19828, n19829, n19830, n19831, n19832, n19833,
    n19834, n19835, n19836, n19837, n19838, n19839,
    n19840, n19841, n19842, n19843, n19844, n19845,
    n19846, n19847, n19848, n19849, n19850, n19851,
    n19852, n19853, n19854, n19855, n19856, n19857,
    n19858, n19859, n19860, n19861, n19862, n19863,
    n19864, n19865, n19866, n19867, n19868, n19869,
    n19870, n19871, n19872, n19873, n19874, n19875,
    n19876, n19877, n19878, n19879, n19880, n19881,
    n19882, n19883, n19884, n19885, n19886, n19887,
    n19888, n19889, n19890, n19891, n19892, n19893,
    n19894, n19895, n19896, n19897, n19898, n19899,
    n19900, n19901, n19902, n19903, n19904, n19905,
    n19906, n19907, n19908, n19909, n19910, n19911,
    n19912, n19913, n19914, n19915, n19916, n19917,
    n19918, n19919, n19920, n19921, n19922, n19923,
    n19924, n19925, n19926, n19927, n19928, n19929,
    n19930, n19931, n19932, n19933, n19934, n19935,
    n19936, n19937, n19938, n19939, n19940, n19941,
    n19942, n19943, n19944, n19945, n19946, n19947,
    n19948, n19949, n19950, n19951, n19952, n19953,
    n19954, n19955, n19956, n19957, n19958, n19959,
    n19960, n19961, n19962, n19963, n19964, n19965,
    n19966, n19967, n19968, n19969, n19970, n19971,
    n19972, n19973, n19974, n19975, n19976, n19977,
    n19978, n19979, n19980, n19981, n19982, n19983,
    n19984, n19985, n19986, n19987, n19988, n19989,
    n19990, n19991, n19992, n19993, n19994, n19995,
    n19996, n19997, n19998, n19999, n20000, n20001,
    n20002, n20003, n20004, n20005, n20006, n20007,
    n20008, n20009, n20010, n20011, n20012, n20013,
    n20014, n20015, n20016, n20017, n20018, n20019,
    n20020, n20021, n20022, n20023, n20024, n20025,
    n20026, n20027, n20028, n20029, n20030, n20031,
    n20032, n20033, n20034, n20035, n20036, n20037,
    n20038, n20039, n20040, n20041, n20042, n20043,
    n20044, n20045, n20046, n20047, n20048, n20049,
    n20050, n20051, n20052, n20053, n20054, n20055,
    n20056, n20057, n20058, n20059, n20060, n20061,
    n20062, n20063, n20064, n20065, n20066, n20067,
    n20068, n20069, n20070, n20071, n20072, n20073,
    n20074, n20075, n20076, n20077, n20078, n20079,
    n20080, n20081, n20082, n20083, n20084, n20085,
    n20086, n20087, n20088, n20089, n20090, n20091,
    n20092, n20093, n20094, n20095, n20096, n20097,
    n20098, n20099, n20100, n20101, n20102, n20103,
    n20104, n20106, n20107, n20108, n20109, n20110,
    n20111, n20112, n20113, n20114, n20115, n20116,
    n20117, n20118, n20119, n20120, n20121, n20122,
    n20123, n20124, n20125, n20126, n20127, n20128,
    n20129, n20130, n20131, n20132, n20133, n20134,
    n20135, n20136, n20137, n20138, n20139, n20140,
    n20141, n20142, n20143, n20144, n20145, n20146,
    n20147, n20148, n20149, n20150, n20151, n20152,
    n20153, n20154, n20155, n20156, n20157, n20158,
    n20159, n20160, n20161, n20162, n20163, n20164,
    n20165, n20166, n20167, n20168, n20169, n20170,
    n20171, n20172, n20173, n20174, n20175, n20176,
    n20177, n20178, n20179, n20180, n20181, n20182,
    n20183, n20184, n20185, n20186, n20187, n20188,
    n20189, n20190, n20191, n20192, n20193, n20194,
    n20195, n20196, n20197, n20198, n20199, n20200,
    n20201, n20202, n20203, n20204, n20205, n20206,
    n20207, n20208, n20209, n20210, n20211, n20212,
    n20213, n20214, n20215, n20216, n20217, n20218,
    n20219, n20220, n20221, n20222, n20223, n20224,
    n20225, n20226, n20227, n20228, n20229, n20230,
    n20231, n20232, n20233, n20234, n20235, n20236,
    n20237, n20238, n20239, n20240, n20241, n20242,
    n20243, n20244, n20245, n20246, n20247, n20248,
    n20249, n20250, n20251, n20252, n20253, n20254,
    n20255, n20256, n20257, n20258, n20259, n20260,
    n20261, n20262, n20263, n20264, n20265, n20266,
    n20267, n20268, n20269, n20270, n20271, n20272,
    n20273, n20274, n20275, n20276, n20277, n20278,
    n20279, n20280, n20281, n20282, n20283, n20284,
    n20285, n20286, n20287, n20288, n20289, n20290,
    n20291, n20292, n20293, n20294, n20295, n20296,
    n20297, n20298, n20299, n20300, n20301, n20302,
    n20303, n20304, n20305, n20306, n20307, n20308,
    n20309, n20310, n20311, n20312, n20313, n20314,
    n20315, n20316, n20317, n20318, n20319, n20320,
    n20321, n20322, n20323, n20324, n20325, n20326,
    n20327, n20328, n20329, n20330, n20331, n20332,
    n20333, n20334, n20335, n20336, n20337, n20338,
    n20339, n20340, n20341, n20342, n20343, n20344,
    n20345, n20346, n20347, n20348, n20349, n20350,
    n20351, n20352, n20353, n20354, n20355, n20356,
    n20357, n20358, n20359, n20360, n20361, n20362,
    n20363, n20364, n20365, n20366, n20367, n20368,
    n20369, n20370, n20371, n20372, n20373, n20374,
    n20375, n20376, n20377, n20378, n20379, n20380,
    n20381, n20382, n20383, n20384, n20385, n20386,
    n20387, n20388, n20389, n20390, n20391, n20392,
    n20393, n20394, n20395, n20396, n20397, n20398,
    n20399, n20400, n20401, n20402, n20403, n20404,
    n20405, n20406, n20407, n20408, n20409, n20410,
    n20411, n20412, n20413, n20414, n20415, n20416,
    n20417, n20418, n20419, n20420, n20421, n20422,
    n20423, n20424, n20425, n20426, n20427, n20428,
    n20429, n20430, n20431, n20432, n20433, n20434,
    n20435, n20436, n20437, n20438, n20439, n20440,
    n20441, n20442, n20443, n20444, n20445, n20446,
    n20447, n20448, n20449, n20450, n20451, n20452,
    n20453, n20454, n20455, n20456, n20457, n20458,
    n20459, n20460, n20461, n20462, n20463, n20464,
    n20465, n20466, n20467, n20468, n20469, n20470,
    n20471, n20472, n20473, n20474, n20475, n20476,
    n20477, n20478, n20479, n20480, n20481, n20482,
    n20483, n20484, n20485, n20486, n20487, n20488,
    n20489, n20490, n20491, n20492, n20493, n20494,
    n20495, n20496, n20497, n20498, n20499, n20500,
    n20501, n20502, n20503, n20504, n20505, n20506,
    n20507, n20508, n20509, n20510, n20511, n20512,
    n20513, n20514, n20515, n20516, n20517, n20518,
    n20519, n20520, n20521, n20522, n20523, n20524,
    n20525, n20526, n20527, n20528, n20529, n20530,
    n20531, n20532, n20533, n20534, n20535, n20536,
    n20537, n20538, n20539, n20540, n20541, n20542,
    n20543, n20544, n20545, n20546, n20547, n20548,
    n20549, n20550, n20551, n20552, n20553, n20554,
    n20555, n20556, n20557, n20558, n20559, n20560,
    n20561, n20562, n20563, n20564, n20565, n20566,
    n20567, n20568, n20569, n20570, n20571, n20572,
    n20573, n20574, n20575, n20576, n20577, n20578,
    n20579, n20580, n20581, n20582, n20583, n20584,
    n20585, n20586, n20587, n20588, n20589, n20590,
    n20591, n20592, n20593, n20594, n20595, n20596,
    n20597, n20598, n20599, n20600, n20601, n20602,
    n20603, n20604, n20605, n20606, n20607, n20608,
    n20609, n20610, n20611, n20612, n20613, n20614,
    n20615, n20616, n20617, n20618, n20619, n20620,
    n20621, n20622, n20623, n20624, n20625, n20626,
    n20627, n20628, n20629, n20630, n20631, n20632,
    n20633, n20634, n20635, n20636, n20637, n20638,
    n20639, n20640, n20641, n20642, n20643, n20644,
    n20645, n20646, n20647, n20648, n20649, n20650,
    n20651, n20652, n20653, n20654, n20655, n20656,
    n20657, n20658, n20659, n20660, n20661, n20662,
    n20663, n20664, n20665, n20666, n20667, n20668,
    n20669, n20670, n20671, n20672, n20673, n20674,
    n20675, n20676, n20677, n20678, n20679, n20680,
    n20681, n20682, n20683, n20684, n20685, n20686,
    n20687, n20688, n20689, n20690, n20691, n20692,
    n20693, n20694, n20695, n20696, n20697, n20698,
    n20699, n20700, n20701, n20702, n20703, n20704,
    n20705, n20706, n20707, n20708, n20709, n20710,
    n20711, n20712, n20713, n20714, n20715, n20716,
    n20717, n20718, n20719, n20720, n20721, n20722,
    n20723, n20724, n20725, n20726, n20727, n20728,
    n20729, n20730, n20731, n20732, n20733, n20734,
    n20735, n20736, n20737, n20738, n20739, n20740,
    n20741, n20742, n20743, n20744, n20745, n20746,
    n20747, n20748, n20749, n20750, n20751, n20752,
    n20754, n20755, n20756, n20757, n20758, n20759,
    n20760, n20761, n20762, n20763, n20764, n20765,
    n20766, n20767, n20768, n20769, n20770, n20771,
    n20772, n20773, n20774, n20775, n20776, n20777,
    n20778, n20779, n20780, n20781, n20782, n20783,
    n20784, n20785, n20786, n20787, n20788, n20789,
    n20790, n20791, n20792, n20793, n20794, n20795,
    n20796, n20797, n20798, n20799, n20800, n20801,
    n20802, n20803, n20804, n20805, n20806, n20807,
    n20808, n20809, n20810, n20811, n20812, n20813,
    n20814, n20815, n20816, n20817, n20818, n20819,
    n20820, n20821, n20822, n20823, n20824, n20825,
    n20826, n20827, n20828, n20829, n20830, n20831,
    n20832, n20833, n20834, n20835, n20836, n20837,
    n20838, n20839, n20840, n20841, n20842, n20843,
    n20844, n20845, n20846, n20847, n20848, n20849,
    n20850, n20851, n20852, n20853, n20854, n20855,
    n20856, n20857, n20858, n20859, n20860, n20861,
    n20862, n20863, n20864, n20865, n20866, n20867,
    n20868, n20869, n20870, n20871, n20872, n20873,
    n20874, n20875, n20876, n20877, n20878, n20879,
    n20880, n20881, n20882, n20883, n20884, n20885,
    n20886, n20887, n20888, n20889, n20890, n20891,
    n20892, n20893, n20894, n20895, n20896, n20897,
    n20898, n20899, n20900, n20901, n20902, n20903,
    n20904, n20905, n20906, n20907, n20908, n20909,
    n20910, n20911, n20912, n20913, n20914, n20915,
    n20916, n20917, n20918, n20919, n20920, n20921,
    n20922, n20923, n20924, n20925, n20926, n20927,
    n20928, n20929, n20930, n20931, n20932, n20933,
    n20934, n20935, n20936, n20937, n20938, n20939,
    n20940, n20941, n20942, n20943, n20944, n20945,
    n20946, n20947, n20948, n20949, n20950, n20951,
    n20952, n20953, n20954, n20955, n20956, n20957,
    n20958, n20959, n20960, n20961, n20962, n20963,
    n20964, n20965, n20966, n20967, n20968, n20969,
    n20970, n20971, n20972, n20973, n20974, n20975,
    n20976, n20977, n20978, n20979, n20980, n20981,
    n20982, n20983, n20984, n20985, n20986, n20987,
    n20988, n20989, n20990, n20991, n20992, n20993,
    n20994, n20995, n20996, n20997, n20998, n20999,
    n21000, n21001, n21002, n21003, n21004, n21005,
    n21006, n21007, n21008, n21009, n21010, n21011,
    n21012, n21013, n21014, n21015, n21016, n21017,
    n21018, n21019, n21020, n21021, n21022, n21023,
    n21024, n21025, n21026, n21027, n21028, n21029,
    n21030, n21031, n21032, n21033, n21034, n21035,
    n21036, n21037, n21038, n21039, n21040, n21041,
    n21042, n21043, n21044, n21045, n21046, n21047,
    n21048, n21049, n21050, n21051, n21052, n21053,
    n21054, n21055, n21056, n21057, n21058, n21059,
    n21060, n21061, n21062, n21063, n21064, n21065,
    n21066, n21067, n21068, n21069, n21070, n21071,
    n21072, n21073, n21074, n21075, n21076, n21077,
    n21078, n21079, n21080, n21081, n21082, n21083,
    n21084, n21085, n21086, n21087, n21088, n21089,
    n21090, n21091, n21092, n21093, n21094, n21095,
    n21096, n21097, n21098, n21099, n21100, n21101,
    n21102, n21103, n21104, n21105, n21106, n21107,
    n21108, n21109, n21110, n21111, n21112, n21113,
    n21114, n21115, n21116, n21117, n21118, n21119,
    n21120, n21121, n21122, n21123, n21124, n21125,
    n21126, n21127, n21128, n21129, n21130, n21131,
    n21132, n21133, n21134, n21135, n21136, n21137,
    n21138, n21139, n21140, n21141, n21142, n21143,
    n21144, n21145, n21146, n21147, n21148, n21149,
    n21150, n21151, n21152, n21153, n21154, n21155,
    n21156, n21157, n21158, n21159, n21160, n21161,
    n21162, n21163, n21164, n21165, n21166, n21167,
    n21168, n21169, n21170, n21171, n21172, n21173,
    n21174, n21175, n21176, n21177, n21178, n21179,
    n21180, n21181, n21182, n21183, n21184, n21185,
    n21186, n21187, n21188, n21189, n21190, n21191,
    n21192, n21193, n21194, n21195, n21196, n21197,
    n21198, n21199, n21200, n21201, n21202, n21203,
    n21204, n21205, n21206, n21207, n21208, n21209,
    n21210, n21211, n21212, n21213, n21214, n21215,
    n21216, n21217, n21218, n21219, n21220, n21221,
    n21222, n21223, n21224, n21225, n21226, n21227,
    n21228, n21229, n21230, n21231, n21232, n21233,
    n21234, n21235, n21236, n21237, n21238, n21239,
    n21240, n21241, n21242, n21243, n21244, n21245,
    n21246, n21247, n21248, n21249, n21250, n21251,
    n21252, n21253, n21254, n21255, n21256, n21257,
    n21258, n21259, n21260, n21261, n21262, n21263,
    n21264, n21265, n21266, n21267, n21268, n21269,
    n21270, n21271, n21272, n21273, n21274, n21275,
    n21276, n21277, n21278, n21279, n21280, n21281,
    n21282, n21283, n21284, n21285, n21286, n21287,
    n21288, n21289, n21290, n21291, n21292, n21293,
    n21294, n21295, n21296, n21297, n21298, n21299,
    n21300, n21301, n21302, n21303, n21304, n21305,
    n21306, n21307, n21308, n21309, n21310, n21311,
    n21312, n21313, n21314, n21315, n21316, n21317,
    n21318, n21319, n21320, n21321, n21322, n21323,
    n21324, n21325, n21326, n21327, n21328, n21329,
    n21330, n21331, n21332, n21333, n21334, n21335,
    n21336, n21337, n21338, n21339, n21340, n21341,
    n21342, n21343, n21344, n21345, n21346, n21347,
    n21348, n21349, n21350, n21351, n21352, n21353,
    n21354, n21355, n21356, n21357, n21358, n21359,
    n21360, n21361, n21362, n21363, n21364, n21365,
    n21366, n21367, n21368, n21369, n21370, n21371,
    n21372, n21373, n21374, n21375, n21376, n21377,
    n21378, n21379, n21380, n21381, n21382, n21383,
    n21384, n21385, n21386, n21387, n21388, n21389,
    n21390, n21391, n21392, n21393, n21394, n21395,
    n21396, n21397, n21398, n21399, n21401, n21402,
    n21403, n21404, n21405, n21406, n21407, n21408,
    n21409, n21410, n21411, n21412, n21413, n21414,
    n21415, n21416, n21417, n21418, n21419, n21420,
    n21421, n21422, n21423, n21424, n21425, n21426,
    n21427, n21428, n21429, n21430, n21431, n21432,
    n21433, n21434, n21435, n21436, n21437, n21438,
    n21439, n21440, n21441, n21442, n21443, n21444,
    n21445, n21446, n21447, n21448, n21449, n21450,
    n21451, n21452, n21453, n21454, n21455, n21456,
    n21457, n21458, n21459, n21460, n21461, n21462,
    n21463, n21464, n21465, n21466, n21467, n21468,
    n21469, n21470, n21471, n21472, n21473, n21474,
    n21475, n21476, n21477, n21478, n21479, n21480,
    n21481, n21482, n21483, n21484, n21485, n21486,
    n21487, n21488, n21489, n21490, n21491, n21492,
    n21493, n21494, n21495, n21496, n21497, n21498,
    n21499, n21500, n21501, n21502, n21503, n21504,
    n21505, n21506, n21507, n21508, n21509, n21510,
    n21511, n21512, n21513, n21514, n21515, n21516,
    n21517, n21518, n21519, n21520, n21521, n21522,
    n21523, n21524, n21525, n21526, n21527, n21528,
    n21529, n21530, n21531, n21532, n21533, n21534,
    n21535, n21536, n21537, n21538, n21539, n21540,
    n21541, n21542, n21543, n21544, n21545, n21546,
    n21547, n21548, n21549, n21550, n21551, n21552,
    n21553, n21554, n21555, n21556, n21557, n21558,
    n21559, n21560, n21561, n21562, n21563, n21564,
    n21565, n21566, n21567, n21568, n21569, n21570,
    n21571, n21572, n21573, n21574, n21575, n21576,
    n21577, n21578, n21579, n21580, n21581, n21582,
    n21583, n21584, n21585, n21586, n21587, n21588,
    n21589, n21590, n21591, n21592, n21593, n21594,
    n21595, n21596, n21597, n21598, n21599, n21600,
    n21601, n21602, n21603, n21604, n21605, n21606,
    n21607, n21608, n21609, n21610, n21611, n21612,
    n21613, n21614, n21615, n21616, n21617, n21618,
    n21619, n21620, n21621, n21622, n21623, n21624,
    n21625, n21626, n21627, n21628, n21629, n21630,
    n21631, n21632, n21633, n21634, n21635, n21636,
    n21637, n21638, n21639, n21640, n21641, n21642,
    n21643, n21644, n21645, n21646, n21647, n21648,
    n21649, n21650, n21651, n21652, n21653, n21654,
    n21655, n21656, n21657, n21658, n21659, n21660,
    n21661, n21662, n21663, n21664, n21665, n21666,
    n21667, n21668, n21669, n21670, n21671, n21672,
    n21673, n21674, n21675, n21676, n21677, n21678,
    n21679, n21680, n21681, n21682, n21683, n21684,
    n21685, n21686, n21687, n21688, n21689, n21690,
    n21691, n21692, n21693, n21694, n21695, n21696,
    n21697, n21698, n21699, n21700, n21701, n21702,
    n21703, n21704, n21705, n21706, n21707, n21708,
    n21709, n21710, n21711, n21712, n21713, n21714,
    n21715, n21716, n21717, n21718, n21719, n21720,
    n21721, n21722, n21723, n21724, n21725, n21726,
    n21727, n21728, n21729, n21730, n21731, n21732,
    n21733, n21734, n21735, n21736, n21737, n21738,
    n21739, n21740, n21741, n21742, n21743, n21744,
    n21745, n21746, n21747, n21748, n21749, n21750,
    n21751, n21752, n21753, n21754, n21755, n21756,
    n21757, n21758, n21759, n21760, n21761, n21762,
    n21763, n21764, n21765, n21766, n21767, n21768,
    n21769, n21770, n21771, n21772, n21773, n21774,
    n21775, n21776, n21777, n21778, n21779, n21780,
    n21781, n21782, n21783, n21784, n21785, n21786,
    n21787, n21788, n21789, n21790, n21791, n21792,
    n21793, n21794, n21795, n21796, n21797, n21798,
    n21799, n21800, n21801, n21802, n21803, n21804,
    n21805, n21806, n21807, n21808, n21809, n21810,
    n21811, n21812, n21813, n21814, n21815, n21816,
    n21817, n21818, n21819, n21820, n21821, n21822,
    n21823, n21824, n21825, n21826, n21827, n21828,
    n21829, n21830, n21831, n21832, n21833, n21834,
    n21835, n21836, n21837, n21838, n21839, n21840,
    n21841, n21842, n21843, n21844, n21845, n21846,
    n21847, n21848, n21849, n21850, n21851, n21852,
    n21853, n21854, n21855, n21856, n21857, n21858,
    n21859, n21860, n21861, n21862, n21863, n21864,
    n21865, n21866, n21867, n21868, n21869, n21870,
    n21871, n21872, n21873, n21874, n21875, n21876,
    n21877, n21878, n21879, n21880, n21881, n21882,
    n21883, n21884, n21885, n21886, n21887, n21888,
    n21889, n21890, n21891, n21892, n21893, n21894,
    n21895, n21896, n21897, n21898, n21899, n21900,
    n21901, n21902, n21903, n21904, n21905, n21906,
    n21907, n21908, n21909, n21910, n21911, n21912,
    n21913, n21914, n21915, n21916, n21917, n21918,
    n21919, n21920, n21921, n21922, n21923, n21924,
    n21925, n21926, n21927, n21928, n21929, n21930,
    n21931, n21932, n21933, n21934, n21935, n21936,
    n21937, n21938, n21939, n21940, n21941, n21942,
    n21943, n21944, n21945, n21946, n21947, n21948,
    n21949, n21950, n21951, n21952, n21953, n21954,
    n21955, n21956, n21957, n21958, n21959, n21960,
    n21961, n21962, n21963, n21964, n21965, n21966,
    n21967, n21968, n21969, n21970, n21971, n21972,
    n21973, n21974, n21975, n21976, n21977, n21978,
    n21979, n21980, n21981, n21982, n21983, n21984,
    n21985, n21986, n21987, n21988, n21989, n21990,
    n21991, n21992, n21993, n21994, n21995, n21996,
    n21997, n21998, n21999, n22000, n22001, n22002,
    n22003, n22004, n22005, n22006, n22007, n22008,
    n22009, n22010, n22011, n22012, n22013, n22014,
    n22015, n22016, n22017, n22018, n22019, n22020,
    n22021, n22022, n22023, n22024, n22025, n22026,
    n22027, n22028, n22029, n22030, n22031, n22032,
    n22033, n22034, n22035, n22036, n22037, n22038,
    n22039, n22040, n22041, n22042, n22043, n22044,
    n22045, n22046, n22048, n22049, n22050, n22051,
    n22052, n22053, n22054, n22055, n22056, n22057,
    n22058, n22059, n22060, n22061, n22062, n22063,
    n22064, n22065, n22066, n22067, n22068, n22069,
    n22070, n22071, n22072, n22073, n22074, n22075,
    n22076, n22077, n22078, n22079, n22080, n22081,
    n22082, n22083, n22084, n22085, n22086, n22087,
    n22088, n22089, n22090, n22091, n22092, n22093,
    n22094, n22095, n22096, n22097, n22098, n22099,
    n22100, n22101, n22102, n22103, n22104, n22105,
    n22106, n22107, n22108, n22109, n22110, n22111,
    n22112, n22113, n22114, n22115, n22116, n22117,
    n22118, n22119, n22120, n22121, n22122, n22123,
    n22124, n22125, n22126, n22127, n22128, n22129,
    n22130, n22131, n22132, n22133, n22134, n22135,
    n22136, n22137, n22138, n22139, n22140, n22141,
    n22142, n22143, n22144, n22145, n22146, n22147,
    n22148, n22149, n22150, n22151, n22152, n22153,
    n22154, n22155, n22156, n22157, n22158, n22159,
    n22160, n22161, n22162, n22163, n22164, n22165,
    n22166, n22167, n22168, n22169, n22170, n22171,
    n22172, n22173, n22174, n22175, n22176, n22177,
    n22178, n22179, n22180, n22181, n22182, n22183,
    n22184, n22185, n22186, n22187, n22188, n22189,
    n22190, n22191, n22192, n22193, n22194, n22195,
    n22196, n22197, n22198, n22199, n22200, n22201,
    n22202, n22203, n22204, n22205, n22206, n22207,
    n22208, n22209, n22210, n22211, n22212, n22213,
    n22214, n22215, n22216, n22217, n22218, n22219,
    n22220, n22221, n22222, n22223, n22224, n22225,
    n22226, n22227, n22228, n22229, n22230, n22231,
    n22232, n22233, n22234, n22235, n22236, n22237,
    n22238, n22239, n22240, n22241, n22242, n22243,
    n22244, n22245, n22246, n22247, n22248, n22249,
    n22250, n22251, n22252, n22253, n22254, n22255,
    n22256, n22257, n22258, n22259, n22260, n22261,
    n22262, n22263, n22264, n22265, n22266, n22267,
    n22268, n22269, n22270, n22271, n22272, n22273,
    n22274, n22275, n22276, n22277, n22278, n22279,
    n22280, n22281, n22282, n22283, n22284, n22285,
    n22286, n22287, n22288, n22289, n22290, n22291,
    n22292, n22293, n22294, n22295, n22296, n22297,
    n22298, n22299, n22300, n22301, n22302, n22303,
    n22304, n22305, n22306, n22307, n22308, n22309,
    n22310, n22311, n22312, n22313, n22314, n22315,
    n22316, n22317, n22318, n22319, n22320, n22321,
    n22322, n22323, n22324, n22325, n22326, n22327,
    n22328, n22329, n22330, n22331, n22332, n22333,
    n22334, n22335, n22336, n22337, n22338, n22339,
    n22340, n22341, n22342, n22343, n22344, n22345,
    n22346, n22347, n22348, n22349, n22350, n22351,
    n22352, n22353, n22354, n22355, n22356, n22357,
    n22358, n22359, n22360, n22361, n22362, n22363,
    n22364, n22365, n22366, n22367, n22368, n22369,
    n22370, n22371, n22372, n22373, n22374, n22375,
    n22376, n22377, n22378, n22379, n22380, n22381,
    n22382, n22383, n22384, n22385, n22386, n22387,
    n22388, n22389, n22390, n22391, n22392, n22393,
    n22394, n22395, n22396, n22397, n22398, n22399,
    n22400, n22401, n22402, n22403, n22404, n22405,
    n22406, n22407, n22408, n22409, n22410, n22411,
    n22412, n22413, n22414, n22415, n22416, n22417,
    n22418, n22419, n22420, n22421, n22422, n22423,
    n22424, n22425, n22426, n22427, n22428, n22429,
    n22430, n22431, n22432, n22433, n22434, n22435,
    n22436, n22437, n22438, n22439, n22440, n22441,
    n22442, n22443, n22444, n22445, n22446, n22447,
    n22448, n22449, n22450, n22451, n22452, n22453,
    n22454, n22455, n22456, n22457, n22458, n22459,
    n22460, n22461, n22462, n22463, n22464, n22465,
    n22466, n22467, n22468, n22469, n22470, n22471,
    n22472, n22473, n22474, n22475, n22476, n22477,
    n22478, n22479, n22480, n22481, n22482, n22483,
    n22484, n22485, n22486, n22487, n22488, n22489,
    n22490, n22491, n22492, n22493, n22494, n22495,
    n22496, n22497, n22498, n22499, n22500, n22501,
    n22502, n22503, n22504, n22505, n22506, n22507,
    n22508, n22509, n22510, n22511, n22512, n22513,
    n22514, n22515, n22516, n22517, n22518, n22519,
    n22520, n22521, n22522, n22523, n22524, n22525,
    n22526, n22527, n22528, n22529, n22530, n22531,
    n22532, n22533, n22534, n22535, n22536, n22537,
    n22538, n22539, n22540, n22541, n22542, n22543,
    n22544, n22545, n22546, n22547, n22548, n22549,
    n22550, n22551, n22552, n22553, n22554, n22555,
    n22556, n22557, n22558, n22559, n22560, n22561,
    n22562, n22563, n22564, n22565, n22566, n22567,
    n22568, n22569, n22570, n22571, n22572, n22573,
    n22574, n22575, n22576, n22577, n22578, n22579,
    n22580, n22581, n22582, n22583, n22584, n22585,
    n22586, n22587, n22588, n22589, n22590, n22591,
    n22592, n22593, n22594, n22595, n22596, n22597,
    n22598, n22599, n22600, n22601, n22602, n22603,
    n22604, n22605, n22606, n22607, n22608, n22609,
    n22610, n22611, n22612, n22613, n22614, n22615,
    n22616, n22617, n22618, n22619, n22620, n22621,
    n22622, n22623, n22624, n22625, n22626, n22627,
    n22628, n22629, n22630, n22631, n22632, n22633,
    n22634, n22635, n22636, n22637, n22638, n22639,
    n22640, n22641, n22642, n22643, n22644, n22645,
    n22646, n22647, n22648, n22649, n22650, n22651,
    n22652, n22653, n22654, n22655, n22656, n22657,
    n22658, n22659, n22660, n22661, n22662, n22663,
    n22664, n22665, n22666, n22667, n22668, n22669,
    n22670, n22671, n22672, n22673, n22674, n22675,
    n22676, n22677, n22678, n22679, n22680, n22681,
    n22682, n22683, n22684, n22685, n22686, n22687,
    n22688, n22689, n22690, n22691, n22692, n22693,
    n22694, n22695, n22697, n22698, n22699, n22700,
    n22701, n22702, n22703, n22704, n22705, n22706,
    n22707, n22708, n22709, n22710, n22711, n22712,
    n22713, n22714, n22715, n22716, n22717, n22718,
    n22719, n22720, n22721, n22722, n22723, n22724,
    n22725, n22726, n22727, n22728, n22729, n22730,
    n22731, n22732, n22733, n22734, n22735, n22736,
    n22737, n22738, n22739, n22740, n22741, n22742,
    n22743, n22744, n22745, n22746, n22747, n22748,
    n22749, n22750, n22751, n22752, n22753, n22754,
    n22755, n22756, n22757, n22758, n22759, n22760,
    n22761, n22762, n22763, n22764, n22765, n22766,
    n22767, n22768, n22769, n22770, n22771, n22772,
    n22773, n22774, n22775, n22776, n22777, n22778,
    n22779, n22780, n22781, n22782, n22783, n22784,
    n22785, n22786, n22787, n22788, n22789, n22790,
    n22791, n22792, n22793, n22794, n22795, n22796,
    n22797, n22798, n22799, n22800, n22801, n22802,
    n22803, n22804, n22805, n22806, n22807, n22808,
    n22809, n22810, n22811, n22812, n22813, n22814,
    n22815, n22816, n22817, n22818, n22819, n22820,
    n22821, n22822, n22823, n22824, n22825, n22826,
    n22827, n22828, n22829, n22830, n22831, n22832,
    n22833, n22834, n22835, n22836, n22837, n22838,
    n22839, n22840, n22841, n22842, n22843, n22844,
    n22845, n22846, n22847, n22848, n22849, n22850,
    n22851, n22852, n22853, n22854, n22855, n22856,
    n22857, n22858, n22859, n22860, n22861, n22862,
    n22863, n22864, n22865, n22866, n22867, n22868,
    n22869, n22870, n22871, n22872, n22873, n22874,
    n22875, n22876, n22877, n22878, n22879, n22880,
    n22881, n22882, n22883, n22884, n22885, n22886,
    n22887, n22888, n22889, n22890, n22891, n22892,
    n22893, n22894, n22895, n22896, n22897, n22898,
    n22899, n22900, n22901, n22902, n22903, n22904,
    n22905, n22906, n22907, n22908, n22909, n22910,
    n22911, n22912, n22913, n22914, n22915, n22916,
    n22917, n22918, n22919, n22920, n22921, n22922,
    n22923, n22924, n22925, n22926, n22927, n22928,
    n22929, n22930, n22931, n22932, n22933, n22934,
    n22935, n22936, n22937, n22938, n22939, n22940,
    n22941, n22942, n22943, n22944, n22945, n22946,
    n22947, n22948, n22949, n22950, n22951, n22952,
    n22953, n22954, n22955, n22956, n22957, n22958,
    n22959, n22960, n22961, n22962, n22963, n22964,
    n22965, n22966, n22967, n22968, n22969, n22970,
    n22971, n22972, n22973, n22974, n22975, n22976,
    n22977, n22978, n22979, n22980, n22981, n22982,
    n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994,
    n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012,
    n23013, n23014, n23015, n23016, n23017, n23018,
    n23019, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n23028, n23029, n23030,
    n23031, n23032, n23033, n23034, n23035, n23036,
    n23037, n23038, n23039, n23040, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048,
    n23049, n23050, n23051, n23052, n23053, n23054,
    n23055, n23056, n23057, n23058, n23059, n23060,
    n23061, n23062, n23063, n23064, n23065, n23066,
    n23067, n23068, n23069, n23070, n23071, n23072,
    n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084,
    n23085, n23086, n23087, n23088, n23089, n23090,
    n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102,
    n23103, n23104, n23105, n23106, n23107, n23108,
    n23109, n23110, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120,
    n23121, n23122, n23123, n23124, n23125, n23126,
    n23127, n23128, n23129, n23130, n23131, n23132,
    n23133, n23134, n23135, n23136, n23137, n23138,
    n23139, n23140, n23141, n23142, n23143, n23144,
    n23145, n23146, n23147, n23148, n23149, n23150,
    n23151, n23152, n23153, n23154, n23155, n23156,
    n23157, n23158, n23159, n23160, n23161, n23162,
    n23163, n23164, n23165, n23166, n23167, n23168,
    n23169, n23170, n23171, n23172, n23173, n23174,
    n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186,
    n23187, n23188, n23189, n23190, n23191, n23192,
    n23193, n23194, n23195, n23196, n23197, n23198,
    n23199, n23200, n23201, n23202, n23203, n23204,
    n23205, n23206, n23207, n23208, n23209, n23210,
    n23211, n23212, n23213, n23214, n23215, n23216,
    n23217, n23218, n23219, n23220, n23221, n23222,
    n23223, n23224, n23225, n23226, n23227, n23228,
    n23229, n23230, n23231, n23232, n23233, n23234,
    n23235, n23236, n23237, n23238, n23239, n23240,
    n23241, n23242, n23243, n23244, n23245, n23246,
    n23247, n23248, n23249, n23250, n23251, n23252,
    n23253, n23254, n23255, n23256, n23257, n23258,
    n23259, n23260, n23261, n23262, n23263, n23264,
    n23265, n23266, n23267, n23268, n23269, n23270,
    n23271, n23272, n23273, n23274, n23275, n23276,
    n23277, n23278, n23279, n23280, n23281, n23282,
    n23283, n23284, n23285, n23286, n23287, n23288,
    n23289, n23290, n23291, n23292, n23293, n23294,
    n23295, n23296, n23297, n23298, n23300, n23301,
    n23302, n23303, n23304, n23305, n23306, n23307,
    n23308, n23309, n23310, n23311, n23312, n23313,
    n23314, n23315, n23316, n23317, n23318, n23319,
    n23320, n23321, n23322, n23323, n23324, n23325,
    n23326, n23327, n23328, n23329, n23330, n23331,
    n23332, n23333, n23334, n23335, n23336, n23337,
    n23338, n23339, n23340, n23341, n23342, n23343,
    n23344, n23345, n23346, n23347, n23348, n23349,
    n23350, n23351, n23352, n23353, n23354, n23355,
    n23356, n23357, n23358, n23359, n23360, n23361,
    n23362, n23363, n23364, n23365, n23366, n23367,
    n23368, n23369, n23370, n23371, n23372, n23373,
    n23374, n23375, n23376, n23377, n23378, n23379,
    n23380, n23381, n23382, n23383, n23384, n23385,
    n23386, n23387, n23388, n23389, n23390, n23391,
    n23392, n23393, n23394, n23395, n23396, n23397,
    n23398, n23399, n23400, n23401, n23402, n23403,
    n23404, n23405, n23406, n23407, n23408, n23409,
    n23410, n23411, n23412, n23413, n23414, n23415,
    n23416, n23417, n23418, n23419, n23420, n23421,
    n23422, n23423, n23424, n23425, n23426, n23427,
    n23428, n23429, n23430, n23431, n23432, n23433,
    n23434, n23435, n23436, n23437, n23438, n23439,
    n23440, n23441, n23442, n23443, n23444, n23445,
    n23446, n23447, n23448, n23449, n23450, n23451,
    n23452, n23453, n23454, n23455, n23456, n23457,
    n23458, n23459, n23460, n23461, n23462, n23463,
    n23464, n23465, n23466, n23467, n23468, n23469,
    n23470, n23471, n23472, n23473, n23474, n23475,
    n23476, n23477, n23478, n23479, n23480, n23481,
    n23482, n23483, n23484, n23485, n23486, n23487,
    n23488, n23489, n23490, n23491, n23492, n23493,
    n23494, n23495, n23496, n23497, n23498, n23499,
    n23500, n23501, n23502, n23503, n23504, n23505,
    n23506, n23507, n23508, n23509, n23510, n23511,
    n23512, n23513, n23514, n23515, n23516, n23517,
    n23518, n23519, n23520, n23521, n23522, n23523,
    n23524, n23525, n23526, n23527, n23528, n23529,
    n23530, n23531, n23532, n23533, n23534, n23535,
    n23536, n23537, n23538, n23539, n23540, n23541,
    n23542, n23543, n23544, n23545, n23546, n23547,
    n23548, n23549, n23550, n23551, n23552, n23553,
    n23554, n23555, n23556, n23557, n23558, n23559,
    n23560, n23561, n23562, n23563, n23564, n23565,
    n23566, n23567, n23568, n23569, n23570, n23571,
    n23572, n23573, n23574, n23575, n23576, n23577,
    n23578, n23579, n23580, n23581, n23582, n23583,
    n23584, n23585, n23586, n23587, n23588, n23589,
    n23590, n23591, n23592, n23593, n23594, n23595,
    n23596, n23597, n23598, n23599, n23600, n23601,
    n23602, n23603, n23604, n23605, n23606, n23607,
    n23608, n23609, n23610, n23611, n23612, n23613,
    n23614, n23615, n23616, n23617, n23618, n23619,
    n23620, n23621, n23622, n23623, n23624, n23625,
    n23626, n23627, n23628, n23629, n23630, n23631,
    n23632, n23633, n23634, n23635, n23636, n23637,
    n23638, n23639, n23640, n23641, n23642, n23643,
    n23644, n23645, n23646, n23647, n23648, n23649,
    n23650, n23651, n23652, n23653, n23654, n23655,
    n23656, n23657, n23658, n23659, n23660, n23661,
    n23662, n23663, n23664, n23665, n23666, n23667,
    n23668, n23669, n23670, n23671, n23672, n23673,
    n23674, n23675, n23676, n23677, n23678, n23679,
    n23680, n23681, n23682, n23683, n23684, n23685,
    n23686, n23687, n23688, n23689, n23690, n23691,
    n23692, n23693, n23694, n23695, n23696, n23697,
    n23698, n23699, n23700, n23701, n23702, n23703,
    n23704, n23705, n23706, n23707, n23708, n23709,
    n23710, n23711, n23712, n23713, n23714, n23715,
    n23716, n23717, n23718, n23719, n23720, n23721,
    n23722, n23723, n23724, n23725, n23726, n23727,
    n23728, n23729, n23730, n23731, n23732, n23733,
    n23734, n23735, n23736, n23737, n23738, n23739,
    n23740, n23741, n23742, n23743, n23744, n23745,
    n23746, n23747, n23748, n23749, n23750, n23751,
    n23752, n23753, n23754, n23755, n23756, n23757,
    n23758, n23759, n23760, n23761, n23762, n23763,
    n23764, n23765, n23766, n23767, n23768, n23769,
    n23770, n23771, n23772, n23773, n23774, n23775,
    n23776, n23777, n23778, n23779, n23780, n23781,
    n23782, n23783, n23784, n23785, n23786, n23787,
    n23788, n23789, n23790, n23791, n23792, n23793,
    n23794, n23795, n23796, n23797, n23798, n23799,
    n23800, n23801, n23802, n23803, n23804, n23805,
    n23806, n23807, n23808, n23809, n23810, n23811,
    n23812, n23813, n23814, n23815, n23816, n23817,
    n23818, n23819, n23820, n23821, n23822, n23823,
    n23824, n23825, n23826, n23827, n23828, n23829,
    n23830, n23831, n23832, n23833, n23834, n23835,
    n23836, n23837, n23838, n23839, n23840, n23841,
    n23842, n23843, n23844, n23845, n23846, n23847,
    n23848, n23849, n23850, n23851, n23852, n23853,
    n23854, n23855, n23856, n23857, n23858, n23859,
    n23860, n23861, n23862, n23863, n23864, n23865,
    n23866, n23867, n23868, n23869, n23870, n23871,
    n23872, n23873, n23874, n23875, n23876, n23877,
    n23878, n23879, n23880, n23881, n23882, n23883,
    n23884, n23885, n23886, n23887, n23888, n23889,
    n23890, n23891, n23892, n23893, n23894, n23895,
    n23896, n23897, n23898, n23899, n23900, n23901,
    n23903, n23904, n23905, n23906, n23907, n23908,
    n23909, n23910, n23911, n23912, n23913, n23914,
    n23915, n23916, n23917, n23918, n23919, n23920,
    n23921, n23922, n23923, n23924, n23925, n23926,
    n23927, n23928, n23929, n23930, n23931, n23932,
    n23933, n23934, n23935, n23936, n23937, n23938,
    n23939, n23940, n23941, n23942, n23943, n23944,
    n23945, n23946, n23947, n23948, n23949, n23950,
    n23951, n23952, n23953, n23954, n23955, n23956,
    n23957, n23958, n23959, n23960, n23961, n23962,
    n23963, n23964, n23965, n23966, n23967, n23968,
    n23969, n23970, n23971, n23972, n23973, n23974,
    n23975, n23976, n23977, n23978, n23979, n23980,
    n23981, n23982, n23983, n23984, n23985, n23986,
    n23987, n23988, n23989, n23990, n23991, n23992,
    n23993, n23994, n23995, n23996, n23997, n23998,
    n23999, n24000, n24001, n24002, n24003, n24004,
    n24005, n24006, n24007, n24008, n24009, n24010,
    n24011, n24012, n24013, n24014, n24015, n24016,
    n24017, n24018, n24019, n24020, n24021, n24022,
    n24023, n24024, n24025, n24026, n24027, n24028,
    n24029, n24030, n24031, n24032, n24033, n24034,
    n24035, n24036, n24037, n24038, n24039, n24040,
    n24041, n24042, n24043, n24044, n24045, n24046,
    n24047, n24048, n24049, n24050, n24051, n24052,
    n24053, n24054, n24055, n24056, n24057, n24058,
    n24059, n24060, n24061, n24062, n24063, n24064,
    n24065, n24066, n24067, n24068, n24069, n24070,
    n24071, n24072, n24073, n24074, n24075, n24076,
    n24077, n24078, n24079, n24080, n24081, n24082,
    n24083, n24084, n24085, n24086, n24087, n24088,
    n24089, n24090, n24091, n24092, n24093, n24094,
    n24095, n24096, n24097, n24098, n24099, n24100,
    n24101, n24102, n24103, n24104, n24105, n24106,
    n24107, n24108, n24109, n24110, n24111, n24112,
    n24113, n24114, n24115, n24116, n24117, n24118,
    n24119, n24120, n24121, n24122, n24123, n24124,
    n24125, n24126, n24127, n24128, n24129, n24130,
    n24131, n24132, n24133, n24134, n24135, n24136,
    n24137, n24138, n24139, n24140, n24141, n24142,
    n24143, n24144, n24145, n24146, n24147, n24148,
    n24149, n24150, n24151, n24152, n24153, n24154,
    n24155, n24156, n24157, n24158, n24159, n24160,
    n24161, n24162, n24163, n24164, n24165, n24166,
    n24167, n24168, n24169, n24170, n24171, n24172,
    n24173, n24174, n24175, n24176, n24177, n24178,
    n24179, n24180, n24181, n24182, n24183, n24184,
    n24185, n24186, n24187, n24188, n24189, n24190,
    n24191, n24192, n24193, n24194, n24195, n24196,
    n24197, n24198, n24199, n24200, n24201, n24202,
    n24203, n24204, n24205, n24206, n24207, n24208,
    n24209, n24210, n24211, n24212, n24213, n24214,
    n24215, n24216, n24217, n24218, n24219, n24220,
    n24221, n24222, n24223, n24224, n24225, n24226,
    n24227, n24228, n24229, n24230, n24231, n24232,
    n24233, n24234, n24235, n24236, n24237, n24238,
    n24239, n24240, n24241, n24242, n24243, n24244,
    n24245, n24246, n24247, n24248, n24249, n24250,
    n24251, n24252, n24253, n24254, n24255, n24256,
    n24257, n24258, n24259, n24260, n24261, n24262,
    n24263, n24264, n24265, n24266, n24267, n24268,
    n24269, n24270, n24271, n24272, n24273, n24274,
    n24275, n24276, n24277, n24278, n24279, n24280,
    n24281, n24282, n24283, n24284, n24285, n24286,
    n24287, n24288, n24289, n24290, n24291, n24292,
    n24293, n24294, n24295, n24296, n24297, n24298,
    n24299, n24300, n24301, n24302, n24303, n24304,
    n24305, n24306, n24307, n24308, n24309, n24310,
    n24311, n24312, n24313, n24314, n24315, n24316,
    n24317, n24318, n24319, n24320, n24321, n24322,
    n24323, n24324, n24325, n24326, n24327, n24328,
    n24329, n24330, n24331, n24332, n24333, n24334,
    n24335, n24336, n24337, n24338, n24339, n24340,
    n24341, n24342, n24343, n24344, n24345, n24346,
    n24347, n24348, n24349, n24350, n24351, n24352,
    n24353, n24354, n24355, n24356, n24357, n24358,
    n24359, n24360, n24361, n24362, n24363, n24364,
    n24365, n24366, n24367, n24368, n24369, n24370,
    n24371, n24372, n24373, n24374, n24375, n24376,
    n24377, n24378, n24379, n24380, n24381, n24382,
    n24383, n24384, n24385, n24386, n24387, n24388,
    n24389, n24390, n24391, n24392, n24393, n24394,
    n24395, n24396, n24397, n24398, n24399, n24400,
    n24401, n24402, n24403, n24404, n24405, n24406,
    n24407, n24408, n24409, n24410, n24411, n24412,
    n24413, n24414, n24415, n24416, n24417, n24418,
    n24419, n24420, n24421, n24422, n24423, n24424,
    n24425, n24426, n24427, n24428, n24429, n24430,
    n24431, n24432, n24433, n24434, n24435, n24436,
    n24437, n24438, n24439, n24440, n24441, n24442,
    n24443, n24444, n24445, n24446, n24447, n24448,
    n24449, n24450, n24451, n24452, n24453, n24454,
    n24455, n24456, n24457, n24458, n24459, n24460,
    n24461, n24462, n24463, n24464, n24465, n24466,
    n24467, n24468, n24469, n24470, n24471, n24472,
    n24473, n24474, n24475, n24476, n24477, n24478,
    n24479, n24480, n24481, n24482, n24483, n24484,
    n24485, n24486, n24487, n24488, n24489, n24490,
    n24491, n24492, n24493, n24494, n24495, n24496,
    n24497, n24498, n24499, n24500, n24501, n24502,
    n24503, n24504, n24506, n24507, n24508, n24509,
    n24510, n24511, n24512, n24513, n24514, n24515,
    n24516, n24517, n24518, n24519, n24520, n24521,
    n24522, n24523, n24524, n24525, n24526, n24527,
    n24528, n24529, n24530, n24531, n24532, n24533,
    n24534, n24535, n24536, n24537, n24538, n24539,
    n24540, n24541, n24542, n24543, n24544, n24545,
    n24546, n24547, n24548, n24549, n24550, n24551,
    n24552, n24553, n24554, n24555, n24556, n24557,
    n24558, n24559, n24560, n24561, n24562, n24563,
    n24564, n24565, n24566, n24567, n24568, n24569,
    n24570, n24571, n24572, n24573, n24574, n24575,
    n24576, n24577, n24578, n24579, n24580, n24581,
    n24582, n24583, n24584, n24585, n24586, n24587,
    n24588, n24589, n24590, n24591, n24592, n24593,
    n24594, n24595, n24596, n24597, n24598, n24599,
    n24600, n24601, n24602, n24603, n24604, n24605,
    n24606, n24607, n24608, n24609, n24610, n24611,
    n24612, n24613, n24614, n24615, n24616, n24617,
    n24618, n24619, n24620, n24621, n24622, n24623,
    n24624, n24625, n24626, n24627, n24628, n24629,
    n24630, n24631, n24632, n24633, n24634, n24635,
    n24636, n24637, n24638, n24639, n24640, n24641,
    n24642, n24643, n24644, n24645, n24646, n24647,
    n24648, n24649, n24650, n24651, n24652, n24653,
    n24654, n24655, n24656, n24657, n24658, n24659,
    n24660, n24661, n24662, n24663, n24664, n24665,
    n24666, n24667, n24668, n24669, n24670, n24671,
    n24672, n24673, n24674, n24675, n24676, n24677,
    n24678, n24679, n24680, n24681, n24682, n24683,
    n24684, n24685, n24686, n24687, n24688, n24689,
    n24690, n24691, n24692, n24693, n24694, n24695,
    n24696, n24697, n24698, n24699, n24700, n24701,
    n24702, n24703, n24704, n24705, n24706, n24707,
    n24708, n24709, n24710, n24711, n24712, n24713,
    n24714, n24715, n24716, n24717, n24718, n24719,
    n24720, n24721, n24722, n24723, n24724, n24725,
    n24726, n24727, n24728, n24729, n24730, n24731,
    n24732, n24733, n24734, n24735, n24736, n24737,
    n24738, n24739, n24740, n24741, n24742, n24743,
    n24744, n24745, n24746, n24747, n24748, n24749,
    n24750, n24751, n24752, n24753, n24754, n24755,
    n24756, n24757, n24758, n24759, n24760, n24761,
    n24762, n24763, n24764, n24765, n24766, n24767,
    n24768, n24769, n24770, n24771, n24772, n24773,
    n24774, n24775, n24776, n24777, n24778, n24779,
    n24780, n24781, n24782, n24783, n24784, n24785,
    n24786, n24787, n24788, n24789, n24790, n24791,
    n24792, n24793, n24794, n24795, n24796, n24797,
    n24798, n24799, n24800, n24801, n24802, n24803,
    n24804, n24805, n24806, n24807, n24808, n24809,
    n24810, n24811, n24812, n24813, n24814, n24815,
    n24816, n24817, n24818, n24819, n24820, n24821,
    n24822, n24823, n24824, n24825, n24826, n24827,
    n24828, n24829, n24830, n24831, n24832, n24833,
    n24834, n24835, n24836, n24837, n24838, n24839,
    n24840, n24841, n24842, n24843, n24844, n24845,
    n24846, n24847, n24848, n24849, n24850, n24851,
    n24852, n24853, n24854, n24855, n24856, n24857,
    n24858, n24859, n24860, n24861, n24862, n24863,
    n24864, n24865, n24866, n24867, n24868, n24869,
    n24870, n24871, n24872, n24873, n24874, n24875,
    n24876, n24877, n24878, n24879, n24880, n24881,
    n24882, n24883, n24884, n24885, n24886, n24887,
    n24888, n24889, n24890, n24891, n24892, n24893,
    n24894, n24895, n24896, n24897, n24898, n24899,
    n24900, n24901, n24902, n24903, n24904, n24905,
    n24906, n24907, n24908, n24909, n24910, n24911,
    n24912, n24913, n24914, n24915, n24916, n24917,
    n24918, n24919, n24920, n24921, n24922, n24923,
    n24924, n24925, n24926, n24927, n24928, n24929,
    n24930, n24931, n24932, n24933, n24934, n24935,
    n24936, n24937, n24938, n24939, n24940, n24941,
    n24942, n24943, n24944, n24945, n24946, n24947,
    n24948, n24949, n24950, n24951, n24952, n24953,
    n24954, n24955, n24956, n24957, n24958, n24959,
    n24960, n24961, n24962, n24963, n24964, n24965,
    n24966, n24967, n24968, n24969, n24970, n24971,
    n24972, n24973, n24974, n24975, n24976, n24977,
    n24978, n24979, n24980, n24981, n24982, n24983,
    n24984, n24985, n24986, n24987, n24988, n24989,
    n24990, n24991, n24992, n24993, n24994, n24995,
    n24996, n24997, n24998, n24999, n25000, n25001,
    n25002, n25003, n25004, n25005, n25006, n25007,
    n25008, n25009, n25010, n25011, n25012, n25013,
    n25014, n25015, n25016, n25017, n25018, n25019,
    n25020, n25021, n25022, n25023, n25024, n25025,
    n25026, n25027, n25028, n25029, n25030, n25031,
    n25032, n25033, n25034, n25035, n25036, n25037,
    n25038, n25039, n25040, n25041, n25042, n25043,
    n25044, n25045, n25046, n25047, n25048, n25049,
    n25050, n25051, n25052, n25053, n25054, n25055,
    n25056, n25057, n25058, n25059, n25060, n25061,
    n25062, n25063, n25064, n25065, n25066, n25067,
    n25068, n25069, n25070, n25071, n25072, n25073,
    n25074, n25075, n25076, n25077, n25078, n25079,
    n25080, n25081, n25082, n25083, n25084, n25085,
    n25086, n25087, n25088, n25089, n25090, n25091,
    n25092, n25094, n25095, n25096, n25097, n25098,
    n25099, n25100, n25101, n25102, n25103, n25104,
    n25105, n25106, n25107, n25108, n25109, n25110,
    n25111, n25112, n25113, n25114, n25115, n25116,
    n25117, n25118, n25119, n25120, n25121, n25122,
    n25123, n25124, n25125, n25126, n25127, n25128,
    n25129, n25130, n25131, n25132, n25133, n25134,
    n25135, n25136, n25137, n25138, n25139, n25140,
    n25141, n25142, n25143, n25144, n25145, n25146,
    n25147, n25148, n25149, n25150, n25151, n25152,
    n25153, n25154, n25155, n25156, n25157, n25158,
    n25159, n25160, n25161, n25162, n25163, n25164,
    n25165, n25166, n25167, n25168, n25169, n25170,
    n25171, n25172, n25173, n25174, n25175, n25176,
    n25177, n25178, n25179, n25180, n25181, n25182,
    n25183, n25184, n25185, n25186, n25187, n25188,
    n25189, n25190, n25191, n25192, n25193, n25194,
    n25195, n25196, n25197, n25198, n25199, n25200,
    n25201, n25202, n25203, n25204, n25205, n25206,
    n25207, n25208, n25209, n25210, n25211, n25212,
    n25213, n25214, n25215, n25216, n25217, n25218,
    n25219, n25220, n25221, n25222, n25223, n25224,
    n25225, n25226, n25227, n25228, n25229, n25230,
    n25231, n25232, n25233, n25234, n25235, n25236,
    n25237, n25238, n25239, n25240, n25241, n25242,
    n25243, n25244, n25245, n25246, n25247, n25248,
    n25249, n25250, n25251, n25252, n25253, n25254,
    n25255, n25256, n25257, n25258, n25259, n25260,
    n25261, n25262, n25263, n25264, n25265, n25266,
    n25267, n25268, n25269, n25270, n25271, n25272,
    n25273, n25274, n25275, n25276, n25277, n25278,
    n25279, n25280, n25281, n25282, n25283, n25284,
    n25285, n25286, n25287, n25288, n25289, n25290,
    n25291, n25292, n25293, n25294, n25295, n25296,
    n25297, n25298, n25299, n25300, n25301, n25302,
    n25303, n25304, n25305, n25306, n25307, n25308,
    n25309, n25310, n25311, n25312, n25313, n25314,
    n25315, n25316, n25317, n25318, n25319, n25320,
    n25321, n25322, n25323, n25324, n25325, n25326,
    n25327, n25328, n25329, n25330, n25331, n25332,
    n25333, n25334, n25335, n25336, n25337, n25338,
    n25339, n25340, n25341, n25342, n25343, n25344,
    n25345, n25346, n25347, n25348, n25349, n25350,
    n25351, n25352, n25353, n25354, n25355, n25356,
    n25357, n25358, n25359, n25360, n25361, n25362,
    n25363, n25364, n25365, n25366, n25367, n25368,
    n25369, n25370, n25371, n25372, n25373, n25374,
    n25375, n25376, n25377, n25378, n25379, n25380,
    n25381, n25382, n25383, n25384, n25385, n25386,
    n25387, n25388, n25389, n25390, n25391, n25392,
    n25393, n25394, n25395, n25396, n25397, n25398,
    n25399, n25400, n25401, n25402, n25403, n25404,
    n25405, n25406, n25407, n25408, n25409, n25410,
    n25411, n25412, n25413, n25414, n25415, n25416,
    n25417, n25418, n25419, n25420, n25421, n25422,
    n25423, n25424, n25425, n25426, n25427, n25428,
    n25429, n25430, n25431, n25432, n25433, n25434,
    n25435, n25436, n25437, n25438, n25439, n25440,
    n25441, n25442, n25443, n25444, n25445, n25446,
    n25447, n25448, n25449, n25450, n25451, n25452,
    n25453, n25454, n25455, n25456, n25457, n25458,
    n25459, n25460, n25461, n25462, n25463, n25464,
    n25465, n25466, n25467, n25468, n25469, n25470,
    n25471, n25472, n25473, n25474, n25475, n25476,
    n25477, n25478, n25479, n25480, n25481, n25482,
    n25483, n25484, n25485, n25486, n25487, n25488,
    n25489, n25490, n25491, n25492, n25493, n25494,
    n25495, n25496, n25497, n25498, n25499, n25500,
    n25501, n25502, n25503, n25504, n25505, n25506,
    n25507, n25508, n25509, n25510, n25511, n25512,
    n25513, n25514, n25515, n25516, n25517, n25518,
    n25519, n25520, n25521, n25522, n25523, n25524,
    n25525, n25526, n25527, n25528, n25529, n25530,
    n25531, n25532, n25533, n25534, n25535, n25536,
    n25537, n25538, n25539, n25540, n25541, n25542,
    n25543, n25544, n25545, n25546, n25547, n25548,
    n25549, n25550, n25551, n25552, n25553, n25554,
    n25555, n25556, n25557, n25558, n25559, n25560,
    n25561, n25562, n25563, n25564, n25565, n25566,
    n25567, n25568, n25569, n25570, n25571, n25572,
    n25573, n25574, n25575, n25576, n25577, n25578,
    n25579, n25580, n25581, n25582, n25583, n25584,
    n25585, n25586, n25587, n25588, n25589, n25590,
    n25591, n25592, n25593, n25594, n25595, n25596,
    n25597, n25598, n25599, n25600, n25601, n25602,
    n25603, n25604, n25605, n25606, n25607, n25608,
    n25609, n25610, n25611, n25612, n25613, n25614,
    n25615, n25616, n25617, n25618, n25619, n25620,
    n25621, n25622, n25623, n25624, n25625, n25626,
    n25627, n25628, n25629, n25630, n25631, n25632,
    n25633, n25634, n25635, n25636, n25637, n25638,
    n25639, n25640, n25641, n25642, n25643, n25644,
    n25645, n25646, n25647, n25648, n25649, n25650,
    n25651, n25652, n25653, n25654, n25655, n25656,
    n25657, n25658, n25659, n25660, n25661, n25662,
    n25663, n25664, n25665, n25666, n25667, n25668,
    n25669, n25670, n25671, n25672, n25673, n25674,
    n25675, n25676, n25677, n25678, n25679, n25680,
    n25681, n25682, n25683, n25684, n25685, n25686,
    n25687, n25688, n25689, n25690, n25691, n25692,
    n25693, n25694, n25695, n25696, n25697, n25698,
    n25699, n25700, n25701, n25702, n25703, n25704,
    n25705, n25706, n25707, n25708, n25709, n25710,
    n25711, n25712, n25713, n25714, n25715, n25716,
    n25717, n25718, n25719, n25720, n25721, n25722,
    n25723, n25724, n25725, n25726, n25727, n25728,
    n25729, n25730, n25731, n25732, n25733, n25734,
    n25735, n25736, n25737, n25738, n25739, n25740,
    n25741, n25742, n25743, n25744, n25745, n25746,
    n25747, n25748, n25749, n25750, n25751, n25752,
    n25753, n25754, n25755, n25757, n25758, n25759,
    n25760, n25761, n25762, n25763, n25764, n25765,
    n25766, n25767, n25768, n25769, n25770, n25771,
    n25772, n25773, n25774, n25775, n25776, n25777,
    n25778, n25779, n25780, n25781, n25782, n25783,
    n25784, n25785, n25786, n25787, n25788, n25789,
    n25790, n25791, n25792, n25793, n25794, n25795,
    n25796, n25797, n25798, n25799, n25800, n25801,
    n25802, n25803, n25804, n25805, n25806, n25807,
    n25808, n25809, n25810, n25811, n25812, n25813,
    n25814, n25815, n25816, n25817, n25818, n25819,
    n25820, n25821, n25822, n25823, n25824, n25825,
    n25826, n25827, n25828, n25829, n25830, n25831,
    n25832, n25833, n25834, n25835, n25836, n25837,
    n25838, n25839, n25840, n25841, n25842, n25843,
    n25844, n25845, n25846, n25847, n25848, n25849,
    n25850, n25851, n25852, n25853, n25854, n25855,
    n25856, n25857, n25858, n25859, n25860, n25861,
    n25862, n25863, n25864, n25865, n25866, n25867,
    n25868, n25869, n25870, n25871, n25872, n25873,
    n25874, n25875, n25876, n25877, n25878, n25879,
    n25880, n25881, n25882, n25883, n25884, n25885,
    n25886, n25887, n25888, n25889, n25890, n25891,
    n25892, n25893, n25894, n25895, n25896, n25897,
    n25898, n25899, n25900, n25901, n25902, n25903,
    n25904, n25905, n25906, n25907, n25908, n25909,
    n25910, n25911, n25912, n25913, n25914, n25915,
    n25916, n25917, n25918, n25919, n25920, n25921,
    n25922, n25923, n25924, n25925, n25926, n25927,
    n25928, n25929, n25930, n25931, n25932, n25933,
    n25934, n25935, n25936, n25937, n25938, n25939,
    n25940, n25941, n25942, n25943, n25944, n25945,
    n25946, n25947, n25948, n25949, n25950, n25951,
    n25952, n25953, n25954, n25955, n25956, n25957,
    n25958, n25959, n25960, n25961, n25962, n25963,
    n25964, n25965, n25966, n25967, n25968, n25969,
    n25970, n25971, n25972, n25973, n25974, n25975,
    n25976, n25977, n25978, n25979, n25980, n25981,
    n25982, n25983, n25984, n25985, n25986, n25987,
    n25988, n25989, n25990, n25991, n25992, n25993,
    n25994, n25995, n25996, n25997, n25998, n25999,
    n26000, n26001, n26002, n26003, n26004, n26005,
    n26006, n26007, n26008, n26009, n26010, n26011,
    n26012, n26013, n26014, n26015, n26016, n26017,
    n26018, n26019, n26020, n26021, n26022, n26023,
    n26024, n26025, n26026, n26027, n26028, n26029,
    n26030, n26031, n26032, n26033, n26034, n26035,
    n26036, n26037, n26038, n26039, n26040, n26041,
    n26042, n26043, n26044, n26045, n26046, n26047,
    n26048, n26049, n26050, n26051, n26052, n26053,
    n26054, n26055, n26056, n26057, n26058, n26059,
    n26060, n26061, n26062, n26063, n26064, n26065,
    n26066, n26067, n26068, n26069, n26070, n26071,
    n26072, n26073, n26074, n26075, n26076, n26077,
    n26078, n26079, n26080, n26081, n26082, n26083,
    n26084, n26085, n26086, n26087, n26088, n26089,
    n26090, n26091, n26092, n26093, n26094, n26095,
    n26096, n26097, n26098, n26099, n26100, n26101,
    n26102, n26103, n26104, n26105, n26106, n26107,
    n26108, n26109, n26110, n26111, n26112, n26113,
    n26114, n26115, n26116, n26117, n26118, n26119,
    n26120, n26121, n26122, n26123, n26124, n26125,
    n26126, n26127, n26128, n26129, n26130, n26131,
    n26132, n26133, n26134, n26135, n26136, n26137,
    n26138, n26139, n26140, n26141, n26142, n26143,
    n26144, n26145, n26146, n26147, n26148, n26149,
    n26150, n26151, n26152, n26153, n26154, n26155,
    n26156, n26157, n26158, n26159, n26160, n26161,
    n26162, n26163, n26164, n26165, n26166, n26167,
    n26168, n26169, n26170, n26171, n26172, n26173,
    n26174, n26175, n26176, n26177, n26178, n26179,
    n26180, n26181, n26182, n26183, n26184, n26185,
    n26186, n26187, n26188, n26189, n26190, n26191,
    n26192, n26193, n26194, n26195, n26196, n26197,
    n26198, n26199, n26200, n26201, n26202, n26203,
    n26204, n26205, n26206, n26207, n26208, n26209,
    n26210, n26211, n26212, n26213, n26214, n26215,
    n26216, n26217, n26218, n26219, n26220, n26221,
    n26222, n26223, n26224, n26225, n26226, n26227,
    n26228, n26229, n26230, n26231, n26232, n26233,
    n26234, n26235, n26236, n26237, n26238, n26239,
    n26240, n26241, n26242, n26243, n26244, n26245,
    n26246, n26247, n26248, n26249, n26250, n26251,
    n26252, n26253, n26254, n26255, n26256, n26257,
    n26258, n26259, n26260, n26261, n26262, n26263,
    n26264, n26265, n26266, n26267, n26268, n26269,
    n26270, n26271, n26272, n26273, n26274, n26275,
    n26276, n26277, n26278, n26279, n26280, n26281,
    n26282, n26283, n26284, n26285, n26286, n26287,
    n26288, n26289, n26290, n26291, n26292, n26293,
    n26294, n26295, n26296, n26297, n26298, n26299,
    n26300, n26301, n26302, n26303, n26304, n26305,
    n26306, n26307, n26308, n26309, n26310, n26311,
    n26312, n26313, n26314, n26315, n26316, n26317,
    n26318, n26319, n26320, n26321, n26322, n26323,
    n26324, n26325, n26326, n26327, n26328, n26329,
    n26330, n26331, n26332, n26333, n26334, n26335,
    n26336, n26337, n26338, n26339, n26340, n26341,
    n26342, n26343, n26344, n26345, n26346, n26347,
    n26348, n26349, n26350, n26351, n26352, n26353,
    n26354, n26355, n26356, n26357, n26358, n26359,
    n26360, n26361, n26362, n26363, n26364, n26365,
    n26366, n26367, n26368, n26369, n26370, n26371,
    n26372, n26373, n26374, n26375, n26376, n26377,
    n26378, n26379, n26380, n26381, n26382, n26383,
    n26384, n26385, n26386, n26387, n26388, n26389,
    n26390, n26391, n26392, n26393, n26394, n26395,
    n26396, n26397, n26398, n26399, n26400, n26401,
    n26402, n26403, n26404, n26405, n26406, n26407,
    n26408, n26409, n26410, n26411, n26412, n26413,
    n26414, n26415, n26416, n26417, n26418, n26419,
    n26420, n26421, n26422, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26431,
    n26432, n26433, n26434, n26435, n26436, n26437,
    n26438, n26439, n26440, n26441, n26442, n26443,
    n26444, n26445, n26446, n26447, n26448, n26449,
    n26450, n26451, n26452, n26453, n26454, n26455,
    n26456, n26457, n26458, n26459, n26460, n26461,
    n26462, n26463, n26464, n26465, n26466, n26467,
    n26468, n26469, n26470, n26471, n26472, n26473,
    n26474, n26475, n26476, n26477, n26478, n26479,
    n26480, n26481, n26482, n26483, n26484, n26485,
    n26486, n26487, n26488, n26489, n26490, n26491,
    n26492, n26493, n26494, n26495, n26496, n26497,
    n26498, n26499, n26500, n26501, n26502, n26503,
    n26504, n26505, n26506, n26507, n26508, n26509,
    n26510, n26511, n26512, n26513, n26514, n26515,
    n26516, n26517, n26518, n26519, n26520, n26521,
    n26522, n26523, n26524, n26525, n26526, n26527,
    n26528, n26529, n26530, n26531, n26532, n26533,
    n26534, n26535, n26536, n26537, n26538, n26539,
    n26540, n26541, n26542, n26543, n26544, n26545,
    n26546, n26547, n26548, n26549, n26550, n26551,
    n26552, n26553, n26554, n26555, n26556, n26557,
    n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26571, n26572, n26573, n26574, n26575,
    n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587,
    n26588, n26589, n26590, n26591, n26592, n26593,
    n26594, n26595, n26596, n26597, n26598, n26599,
    n26600, n26601, n26602, n26603, n26604, n26605,
    n26606, n26607, n26608, n26609, n26610, n26611,
    n26612, n26613, n26614, n26615, n26616, n26617,
    n26618, n26619, n26620, n26621, n26622, n26623,
    n26624, n26625, n26626, n26627, n26628, n26629,
    n26630, n26631, n26632, n26633, n26634, n26635,
    n26636, n26637, n26638, n26639, n26640, n26641,
    n26642, n26643, n26644, n26645, n26646, n26647,
    n26648, n26649, n26650, n26651, n26652, n26653,
    n26654, n26655, n26656, n26657, n26658, n26659,
    n26660, n26661, n26662, n26663, n26664, n26665,
    n26666, n26667, n26668, n26669, n26670, n26671,
    n26672, n26673, n26674, n26675, n26676, n26677,
    n26678, n26679, n26680, n26681, n26682, n26683,
    n26684, n26685, n26686, n26687, n26688, n26689,
    n26690, n26691, n26692, n26693, n26694, n26695,
    n26696, n26697, n26698, n26699, n26700, n26701,
    n26702, n26703, n26704, n26705, n26706, n26707,
    n26708, n26709, n26710, n26711, n26712, n26713,
    n26714, n26715, n26716, n26717, n26718, n26719,
    n26720, n26721, n26722, n26723, n26724, n26725,
    n26726, n26727, n26728, n26729, n26730, n26731,
    n26732, n26733, n26734, n26735, n26736, n26737,
    n26738, n26739, n26740, n26741, n26742, n26743,
    n26744, n26745, n26746, n26747, n26748, n26749,
    n26750, n26751, n26752, n26753, n26754, n26755,
    n26756, n26757, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767,
    n26768, n26769, n26770, n26771, n26772, n26773,
    n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785,
    n26786, n26787, n26788, n26789, n26790, n26791,
    n26792, n26793, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26802, n26803,
    n26804, n26805, n26806, n26807, n26808, n26809,
    n26810, n26811, n26812, n26813, n26814, n26815,
    n26816, n26817, n26818, n26819, n26820, n26821,
    n26822, n26823, n26824, n26825, n26826, n26827,
    n26828, n26829, n26830, n26831, n26832, n26833,
    n26834, n26835, n26836, n26837, n26838, n26839,
    n26840, n26841, n26842, n26843, n26844, n26845,
    n26846, n26847, n26848, n26849, n26850, n26851,
    n26852, n26853, n26854, n26855, n26856, n26857,
    n26858, n26859, n26860, n26861, n26862, n26863,
    n26864, n26865, n26866, n26867, n26868, n26869,
    n26870, n26871, n26872, n26873, n26874, n26875,
    n26876, n26877, n26878, n26879, n26880, n26881,
    n26882, n26883, n26884, n26885, n26886, n26887,
    n26888, n26889, n26890, n26891, n26892, n26893,
    n26894, n26895, n26896, n26897, n26898, n26899,
    n26900, n26901, n26902, n26903, n26904, n26905,
    n26906, n26907, n26908, n26909, n26910, n26911,
    n26912, n26913, n26914, n26915, n26916, n26917,
    n26918, n26919, n26920, n26921, n26922, n26923,
    n26924, n26925, n26926, n26927, n26928, n26929,
    n26930, n26931, n26932, n26933, n26934, n26935,
    n26936, n26937, n26938, n26939, n26940, n26941,
    n26942, n26943, n26944, n26945, n26946, n26947,
    n26948, n26949, n26950, n26951, n26952, n26953,
    n26954, n26955, n26956, n26957, n26958, n26959,
    n26960, n26961, n26962, n26963, n26964, n26965,
    n26966, n26967, n26968, n26969, n26970, n26971,
    n26972, n26973, n26974, n26975, n26976, n26977,
    n26978, n26979, n26980, n26981, n26982, n26983,
    n26984, n26985, n26986, n26987, n26988, n26989,
    n26990, n26991, n26992, n26993, n26994, n26995,
    n26996, n26997, n26998, n26999, n27000, n27001,
    n27002, n27003, n27004, n27005, n27006, n27007,
    n27008, n27009, n27010, n27011, n27012, n27013,
    n27014, n27015, n27016, n27017, n27018, n27019,
    n27020, n27021, n27022, n27023, n27024, n27025,
    n27026, n27027, n27028, n27029, n27030, n27031,
    n27032, n27033, n27034, n27035, n27036, n27037,
    n27038, n27039, n27040, n27041, n27042, n27043,
    n27044, n27045, n27046, n27047, n27048, n27049,
    n27050, n27051, n27052, n27053, n27054, n27055,
    n27056, n27057, n27058, n27059, n27060, n27061,
    n27062, n27063, n27064, n27065, n27066, n27067,
    n27068, n27069, n27070, n27071, n27072, n27073,
    n27074, n27075, n27076, n27077, n27078, n27079,
    n27080, n27081, n27082, n27083, n27084, n27085,
    n27086, n27087, n27088, n27089, n27090, n27091,
    n27092, n27093, n27094, n27095, n27096, n27097,
    n27098, n27099, n27100, n27101, n27102, n27103,
    n27104, n27105, n27106, n27107, n27108, n27109,
    n27110, n27111, n27112, n27113, n27114, n27115,
    n27116, n27117, n27118, n27119, n27120, n27121,
    n27122, n27123, n27124, n27125, n27126, n27127,
    n27128, n27129, n27130, n27131, n27132, n27133,
    n27134, n27135, n27136, n27137, n27138, n27139,
    n27140, n27141, n27142, n27143, n27144, n27145,
    n27146, n27147, n27148, n27149, n27150, n27151,
    n27152, n27153, n27154, n27155, n27156, n27157,
    n27158, n27159, n27160, n27161, n27162, n27163,
    n27164, n27165, n27166, n27167, n27168, n27169,
    n27170, n27171, n27172, n27173, n27174, n27175,
    n27176, n27177, n27178, n27179, n27180, n27181,
    n27182, n27183, n27184, n27185, n27186, n27187,
    n27188, n27189, n27190, n27191, n27192, n27193,
    n27194, n27195, n27196, n27197, n27198, n27199,
    n27200, n27201, n27202, n27203, n27204, n27205,
    n27206, n27207, n27208, n27209, n27210, n27211,
    n27212, n27213, n27214, n27215, n27216, n27217,
    n27218, n27219, n27220, n27221, n27222, n27223,
    n27224, n27225, n27226, n27227, n27228, n27229,
    n27230, n27231, n27232, n27233, n27234, n27235,
    n27236, n27237, n27238, n27239, n27240, n27241,
    n27242, n27243, n27244, n27245, n27246, n27247,
    n27248, n27249, n27250, n27251, n27252, n27253,
    n27254, n27255, n27256, n27257, n27258, n27259,
    n27260, n27261, n27262, n27263, n27264, n27265,
    n27266, n27267, n27268, n27269, n27270, n27271,
    n27272, n27273, n27274, n27275, n27276, n27277,
    n27278, n27279, n27280, n27281, n27282, n27283,
    n27284, n27285, n27286, n27287, n27288, n27289,
    n27290, n27291, n27292, n27293, n27294, n27295,
    n27296, n27297, n27298, n27299, n27300, n27301,
    n27302, n27303, n27304, n27305, n27306, n27307,
    n27308, n27309, n27310, n27311, n27312, n27313,
    n27314, n27315, n27316, n27317, n27318, n27319,
    n27320, n27321, n27322, n27323, n27324, n27325,
    n27326, n27327, n27328, n27329, n27330, n27331,
    n27332, n27333, n27334, n27335, n27336, n27337,
    n27338, n27339, n27340, n27341, n27342, n27343,
    n27344, n27345, n27346, n27347, n27348, n27349,
    n27350, n27351, n27352, n27353, n27354, n27355,
    n27356, n27357, n27358, n27359, n27360, n27361,
    n27362, n27363, n27364, n27365, n27366, n27367,
    n27368, n27369, n27370, n27371, n27372, n27373,
    n27374, n27375, n27376, n27377, n27378, n27379,
    n27380, n27381, n27382, n27383, n27384, n27385,
    n27386, n27387, n27388, n27389, n27390, n27391,
    n27392, n27393, n27394, n27395, n27396, n27397,
    n27398, n27399, n27400, n27401, n27402, n27403,
    n27404, n27405, n27406, n27407, n27408, n27409,
    n27410, n27411, n27412, n27413, n27414, n27415,
    n27416, n27417, n27418, n27419, n27420, n27421,
    n27422, n27423, n27424, n27425, n27426, n27427,
    n27428, n27429, n27430, n27431, n27432, n27433,
    n27434, n27435, n27436, n27437, n27438, n27439,
    n27440, n27441, n27442, n27443, n27444, n27445,
    n27446, n27447, n27448, n27449, n27450, n27451,
    n27452, n27453, n27454, n27455, n27456, n27457,
    n27458, n27459, n27460, n27461, n27462, n27463,
    n27464, n27465, n27466, n27467, n27468, n27469,
    n27470, n27471, n27472, n27473, n27474, n27475,
    n27476, n27477, n27478, n27479, n27480, n27481,
    n27482, n27483, n27484, n27485, n27486, n27487,
    n27488, n27489, n27490, n27491, n27492, n27493,
    n27494, n27495, n27496, n27497, n27498, n27499,
    n27500, n27501, n27502, n27503, n27504, n27505,
    n27506, n27507, n27508, n27509, n27510, n27511,
    n27512, n27513, n27514, n27515, n27516, n27517,
    n27518, n27519, n27520, n27521, n27522, n27523,
    n27524, n27525, n27526, n27527, n27528, n27529,
    n27530, n27531, n27532, n27533, n27534, n27535,
    n27536, n27537, n27538, n27539, n27540, n27541,
    n27542, n27543, n27544, n27545, n27546, n27547,
    n27548, n27549, n27550, n27551, n27552, n27553,
    n27554, n27555, n27556, n27557, n27558, n27559,
    n27560, n27561, n27562, n27563, n27564, n27565,
    n27566, n27567, n27568, n27569, n27570, n27571,
    n27572, n27573, n27574, n27575, n27576, n27577,
    n27578, n27579, n27580, n27581, n27582, n27583,
    n27584, n27585, n27586, n27587, n27588, n27589,
    n27590, n27591, n27592, n27593, n27594, n27595,
    n27596, n27597, n27598, n27599, n27600, n27601,
    n27602, n27603, n27604, n27605, n27606, n27607,
    n27608, n27609, n27610, n27611, n27612, n27613,
    n27614, n27615, n27616, n27617, n27618, n27619,
    n27620, n27621, n27622, n27623, n27624, n27625,
    n27626, n27627, n27628, n27629, n27630, n27631,
    n27632, n27633, n27634, n27635, n27636, n27637,
    n27638, n27639, n27640, n27641, n27642, n27643,
    n27644, n27645, n27646, n27647, n27648, n27649,
    n27650, n27651, n27652, n27653, n27654, n27655,
    n27656, n27657, n27658, n27659, n27660, n27661,
    n27662, n27663, n27664, n27665, n27666, n27667,
    n27668, n27669, n27670, n27671, n27672, n27673,
    n27674, n27675, n27676, n27677, n27678, n27679,
    n27680, n27681, n27682, n27683, n27684, n27685,
    n27686, n27687, n27688, n27689, n27690, n27691,
    n27692, n27693, n27694, n27695, n27696, n27697,
    n27698, n27699, n27700, n27701, n27702, n27703,
    n27704, n27705, n27706, n27707, n27708, n27709,
    n27710, n27711, n27712, n27713, n27714, n27715,
    n27716, n27717, n27718, n27719, n27720, n27721,
    n27722, n27723, n27724, n27725, n27726, n27727,
    n27728, n27729, n27730, n27731, n27732, n27733,
    n27734, n27735, n27736, n27737, n27738, n27739,
    n27740, n27741, n27742, n27743, n27744, n27745,
    n27746, n27747, n27748, n27749, n27750, n27751,
    n27752, n27753, n27754, n27755, n27756, n27757,
    n27758, n27759, n27760, n27761, n27762, n27763,
    n27764, n27765, n27766, n27767, n27768, n27769,
    n27770, n27771, n27772, n27773, n27774, n27775,
    n27776, n27777, n27778, n27779, n27780, n27781,
    n27782, n27783, n27784, n27785, n27786, n27787,
    n27788, n27789, n27790, n27791, n27792, n27793,
    n27794, n27795, n27796, n27797, n27798, n27799,
    n27800, n27801, n27802, n27803, n27804, n27805,
    n27806, n27807, n27808, n27809, n27810, n27811,
    n27812, n27813, n27814, n27815, n27816, n27817,
    n27818, n27819, n27820, n27821, n27822, n27823,
    n27824, n27825, n27826, n27827, n27828, n27829,
    n27830, n27831, n27832, n27833, n27834, n27835,
    n27836, n27837, n27838, n27839, n27840, n27841,
    n27842, n27843, n27844, n27845, n27846, n27847,
    n27848, n27849, n27850, n27851, n27852, n27853,
    n27854, n27855, n27856, n27857, n27858, n27859,
    n27860, n27861, n27862, n27863, n27864, n27865,
    n27866, n27867, n27868, n27869, n27870, n27871,
    n27872, n27873, n27874, n27875, n27876, n27877,
    n27878, n27879, n27880, n27881, n27882, n27883,
    n27884, n27885, n27886, n27887, n27888, n27889,
    n27890, n27891, n27892, n27893, n27894, n27895,
    n27896, n27897, n27898, n27899, n27900, n27901,
    n27902, n27903, n27904, n27905, n27906, n27907,
    n27908, n27909, n27910, n27911, n27912, n27913,
    n27914, n27915, n27916, n27917, n27918, n27919,
    n27920, n27921, n27922, n27923, n27924, n27925,
    n27926, n27927, n27928, n27929, n27930, n27931,
    n27932, n27933, n27934, n27935, n27936, n27937,
    n27938, n27939, n27940, n27941, n27942, n27943,
    n27944, n27945, n27946, n27947, n27948, n27949,
    n27950, n27951, n27952, n27953, n27954, n27955,
    n27956, n27957, n27958, n27959, n27960, n27961,
    n27962, n27963, n27964, n27965, n27966, n27967,
    n27968, n27969, n27970, n27971, n27972, n27973,
    n27974, n27975, n27976, n27977, n27978, n27979,
    n27980, n27981, n27982, n27983, n27984, n27985,
    n27986, n27987, n27988, n27989, n27990, n27991,
    n27992, n27993, n27994, n27995, n27996, n27997,
    n27998, n27999, n28000, n28001, n28002, n28003,
    n28004, n28005, n28006, n28007, n28008, n28009,
    n28010, n28011, n28012, n28013, n28014, n28015,
    n28016, n28017, n28018, n28019, n28020, n28021,
    n28022, n28023, n28024, n28025, n28026, n28027,
    n28028, n28029, n28030, n28031, n28032, n28033,
    n28034, n28035, n28036, n28037, n28038, n28039,
    n28040, n28041, n28042, n28043, n28044, n28045,
    n28046, n28047, n28048, n28049, n28050, n28051,
    n28052, n28053, n28054, n28055, n28056, n28057,
    n28058, n28059, n28060, n28061, n28062, n28063,
    n28064, n28065, n28066, n28067, n28068, n28069,
    n28070, n28071, n28072, n28073, n28074, n28075,
    n28076, n28077, n28078, n28079, n28080, n28081,
    n28082, n28083, n28084, n28085, n28086, n28087,
    n28088, n28089, n28090, n28091, n28092, n28093,
    n28094, n28095, n28096, n28097, n28098, n28099,
    n28100, n28101, n28102, n28103, n28104, n28105,
    n28106, n28107, n28108, n28109, n28110, n28111,
    n28112, n28113, n28114, n28115, n28116, n28117,
    n28118, n28119, n28120, n28121, n28122, n28123,
    n28124, n28125, n28126, n28127, n28128, n28129,
    n28130, n28131, n28132, n28133, n28134, n28135,
    n28136, n28137, n28138, n28139, n28140, n28141,
    n28142, n28143, n28144, n28145, n28146, n28147,
    n28148, n28149, n28150, n28151, n28152, n28153,
    n28154, n28155, n28156, n28157, n28158, n28159,
    n28160, n28161, n28162, n28163, n28164, n28165,
    n28166, n28167, n28168, n28169, n28170, n28171,
    n28172, n28173, n28174, n28175, n28176, n28177,
    n28178, n28179, n28180, n28181, n28182, n28183,
    n28184, n28185, n28186, n28187, n28188, n28189,
    n28190, n28191, n28192, n28193, n28194, n28195,
    n28196, n28197, n28198, n28199, n28200, n28201,
    n28202, n28203, n28204, n28205, n28206, n28207,
    n28208, n28209, n28210, n28211, n28212, n28213,
    n28214, n28215, n28216, n28217, n28218, n28219,
    n28220, n28221, n28222, n28223, n28224, n28225,
    n28226, n28227, n28228, n28229, n28230, n28231,
    n28232, n28233, n28234, n28235, n28236, n28237,
    n28238, n28239, n28240, n28241, n28242, n28243,
    n28244, n28245, n28246, n28247, n28248, n28249,
    n28250, n28251, n28252, n28253, n28254, n28255,
    n28256, n28257, n28258, n28259, n28260, n28261,
    n28262, n28263, n28264, n28265, n28266, n28267,
    n28268, n28269, n28270, n28271, n28272, n28273,
    n28274, n28275, n28276, n28277, n28278, n28279,
    n28280, n28281, n28282, n28283, n28284, n28285,
    n28286, n28287, n28288, n28289, n28290, n28291,
    n28292, n28293, n28294, n28295, n28296, n28297,
    n28298, n28299, n28300, n28301, n28302, n28303,
    n28304, n28305, n28306, n28307, n28308, n28309,
    n28310, n28311, n28312, n28313, n28314, n28315,
    n28316, n28317, n28318, n28319, n28320, n28321,
    n28322, n28323, n28324, n28325, n28326, n28327,
    n28328, n28329, n28330, n28331, n28332, n28333,
    n28334, n28335, n28336, n28337, n28338, n28339,
    n28340, n28341, n28342, n28343, n28344, n28345,
    n28346, n28347, n28348, n28349, n28350, n28351,
    n28352, n28353, n28354, n28355, n28356, n28357,
    n28358, n28359, n28360, n28361, n28362, n28363,
    n28364, n28365, n28366, n28367, n28368, n28369,
    n28370, n28371, n28372, n28373, n28374, n28375,
    n28376, n28377, n28378, n28379, n28380, n28381,
    n28382, n28383, n28384, n28385, n28386, n28387,
    n28388, n28389, n28390, n28391, n28392, n28393,
    n28394, n28395, n28396, n28397, n28398, n28399,
    n28400, n28401, n28402, n28403, n28404, n28405,
    n28406, n28407, n28408, n28409, n28410, n28411,
    n28412, n28413, n28414, n28415, n28416, n28417,
    n28418, n28419, n28420, n28421, n28422, n28423,
    n28424, n28425, n28426, n28427, n28428, n28429,
    n28430, n28431, n28432, n28433, n28434, n28435,
    n28436, n28437, n28438, n28439, n28440, n28441,
    n28442, n28443, n28444, n28445, n28446, n28447,
    n28448, n28449, n28450, n28451, n28452, n28453,
    n28454, n28455, n28456, n28457, n28458, n28459,
    n28460, n28461, n28462, n28463, n28464, n28465,
    n28466, n28467, n28468, n28469, n28470, n28471,
    n28472, n28473, n28474, n28475, n28476, n28477,
    n28478, n28479, n28480, n28481, n28482, n28483,
    n28484, n28485, n28486, n28487, n28488, n28489,
    n28490, n28491, n28492, n28493, n28494, n28495,
    n28496, n28497, n28498, n28499, n28500, n28501,
    n28502, n28503, n28504, n28505, n28506, n28507,
    n28508, n28509, n28510, n28511, n28512, n28513,
    n28514, n28515, n28516, n28517, n28518, n28519,
    n28520, n28521, n28522, n28523, n28524, n28525,
    n28526, n28527, n28528, n28529, n28530, n28531,
    n28532, n28533, n28534, n28535, n28536, n28537,
    n28538, n28539, n28540, n28541, n28542, n28543,
    n28544, n28545, n28546, n28547, n28548, n28549,
    n28550, n28551, n28552, n28553, n28554, n28555,
    n28556, n28557, n28558, n28559, n28560, n28561,
    n28562, n28563, n28564, n28565, n28566, n28567,
    n28568, n28569, n28570, n28571, n28572, n28573,
    n28574, n28575, n28576, n28577, n28578, n28579,
    n28580, n28581, n28582, n28583, n28584, n28585,
    n28586, n28587, n28588, n28589, n28590, n28591,
    n28592, n28593, n28594, n28595, n28596, n28597,
    n28598, n28599, n28600, n28601, n28602, n28603,
    n28604, n28605, n28606, n28607, n28608, n28609,
    n28610, n28611, n28612, n28613, n28614, n28615,
    n28616, n28617, n28618, n28619, n28620, n28621,
    n28622, n28623, n28624, n28625, n28626, n28627,
    n28628, n28629, n28630, n28631, n28632, n28633,
    n28634, n28635, n28636, n28637, n28638, n28639,
    n28640, n28641, n28642, n28643, n28644, n28645,
    n28646, n28647, n28648, n28649, n28650, n28651,
    n28652, n28653, n28654, n28655, n28656, n28657,
    n28658, n28659, n28660, n28661, n28662, n28663,
    n28664, n28665, n28666, n28667, n28668, n28669,
    n28670, n28671, n28672, n28673, n28674, n28675,
    n28676, n28677, n28678, n28679, n28680, n28681,
    n28682, n28683, n28684, n28685, n28686, n28687,
    n28688, n28689, n28690, n28691, n28692, n28693,
    n28694, n28695, n28696, n28697, n28698, n28699,
    n28700, n28701, n28702, n28703, n28704, n28705,
    n28706, n28707, n28708, n28709, n28710, n28711,
    n28712, n28713, n28714, n28715, n28716, n28717,
    n28718, n28719, n28720, n28721, n28722, n28723,
    n28724, n28725, n28726, n28727, n28728, n28729,
    n28730, n28731, n28732, n28733, n28734, n28735,
    n28736, n28737, n28738, n28739, n28740, n28741,
    n28742, n28743, n28744, n28745, n28746, n28747,
    n28748, n28749, n28750, n28751, n28752, n28753,
    n28754, n28755, n28756, n28757, n28758, n28759,
    n28760, n28761, n28762, n28763, n28764, n28765,
    n28766, n28767, n28768, n28769, n28770, n28771,
    n28772, n28773, n28774, n28775, n28776, n28777,
    n28778, n28779, n28780, n28781, n28782, n28783,
    n28784, n28785, n28786, n28787, n28788, n28789,
    n28790, n28791, n28792, n28793, n28794, n28795,
    n28796, n28797, n28798, n28799, n28800, n28801,
    n28802, n28803, n28804, n28805, n28806, n28807,
    n28808, n28809, n28810, n28811, n28812, n28813,
    n28814, n28815, n28816, n28817, n28818, n28819,
    n28820, n28821, n28822, n28823, n28824, n28825,
    n28826, n28827, n28828, n28829, n28830, n28831,
    n28832, n28833, n28834, n28835, n28836, n28837,
    n28838, n28839, n28840, n28841, n28842, n28843,
    n28844, n28845, n28846, n28847, n28848, n28849,
    n28850, n28851, n28852, n28853, n28854, n28855,
    n28856, n28857, n28858, n28859, n28860, n28861,
    n28862, n28863, n28864, n28865, n28866, n28867,
    n28868, n28869, n28870, n28871, n28872, n28873,
    n28874, n28875, n28876, n28877, n28878, n28879,
    n28880, n28881, n28882, n28883, n28884, n28885,
    n28886, n28887, n28888, n28889, n28890, n28891,
    n28892, n28893, n28894, n28895, n28896, n28897,
    n28898, n28899, n28900, n28901, n28902, n28903,
    n28904, n28905, n28906, n28907, n28908, n28909,
    n28910, n28911, n28912, n28913, n28914, n28915,
    n28916, n28917, n28918, n28919, n28920, n28921,
    n28922, n28923, n28924, n28925, n28926, n28927,
    n28928, n28929, n28930, n28931, n28932, n28933,
    n28934, n28935, n28936, n28937, n28938, n28939,
    n28940, n28941, n28942, n28943, n28944, n28945,
    n28946, n28947, n28948, n28949, n28950, n28951,
    n28952, n28953, n28954, n28955, n28956, n28957,
    n28958, n28959, n28960, n28961, n28962, n28963,
    n28964, n28965, n28966, n28967, n28968, n28969,
    n28970, n28971, n28972, n28973, n28974, n28975,
    n28976, n28977, n28978, n28979, n28980, n28981,
    n28982, n28983, n28984, n28985, n28986, n28987,
    n28988, n28989, n28990, n28991, n28992, n28993,
    n28994, n28995, n28996, n28997, n28998, n28999,
    n29000, n29001, n29002, n29003, n29004, n29005,
    n29006, n29007, n29008, n29009, n29010, n29011,
    n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023,
    n29024, n29025, n29026, n29027, n29028, n29029,
    n29030, n29031, n29032, n29033, n29034, n29035,
    n29036, n29037, n29038, n29039, n29040, n29041,
    n29042, n29043, n29044, n29045, n29046, n29047,
    n29048, n29049, n29050, n29051, n29052, n29053,
    n29054, n29055, n29056, n29057, n29058, n29059,
    n29060, n29061, n29062, n29063, n29064, n29065,
    n29066, n29067, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077,
    n29078, n29079, n29080, n29081, n29082, n29083,
    n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095,
    n29096, n29097, n29098, n29099, n29100, n29101,
    n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113,
    n29114, n29115, n29116, n29117, n29118, n29119,
    n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131,
    n29132, n29133, n29134, n29135, n29136, n29137,
    n29138, n29139, n29140, n29141, n29142, n29143,
    n29144, n29145, n29146, n29147, n29148, n29149,
    n29150, n29151, n29152, n29153, n29154, n29155,
    n29156, n29157, n29158, n29159, n29160, n29161,
    n29162, n29163, n29164, n29165, n29166, n29167,
    n29168, n29169, n29170, n29171, n29172, n29173,
    n29174, n29175, n29176, n29177, n29178, n29179,
    n29180, n29181, n29182, n29183, n29184, n29185,
    n29186, n29187, n29188, n29189, n29190, n29191,
    n29192, n29193, n29194, n29195, n29196, n29197,
    n29198, n29199, n29200, n29201, n29202, n29203,
    n29204, n29205, n29206, n29207, n29208, n29209,
    n29210, n29211, n29212, n29213, n29214, n29215,
    n29216, n29217, n29218, n29219, n29220, n29221,
    n29222, n29223, n29224, n29225, n29226, n29227,
    n29228, n29229, n29230, n29231, n29232, n29233,
    n29234, n29235, n29236, n29237, n29238, n29239,
    n29240, n29241, n29242, n29243, n29244, n29245,
    n29246, n29247, n29248, n29249, n29250, n29251,
    n29252, n29253, n29254, n29255, n29256, n29257,
    n29258, n29259, n29260, n29261, n29262, n29263,
    n29264, n29265, n29266, n29267, n29268, n29269,
    n29270, n29271, n29272, n29273, n29274, n29275,
    n29276, n29277, n29278, n29279, n29280, n29281,
    n29282, n29283, n29284, n29285, n29286, n29287,
    n29288, n29289, n29290, n29291, n29292, n29293,
    n29294, n29295, n29296, n29297, n29298, n29299,
    n29300, n29301, n29302, n29303, n29304, n29305,
    n29306, n29307, n29308, n29309, n29310, n29311,
    n29312, n29313, n29314, n29315, n29316, n29317,
    n29318, n29319, n29320, n29321, n29322, n29323,
    n29324, n29325, n29326, n29327, n29328, n29329,
    n29330, n29331, n29332, n29333, n29334, n29335,
    n29336, n29337, n29338, n29339, n29340, n29341,
    n29342, n29343, n29344, n29345, n29346, n29347,
    n29348, n29349, n29350, n29351, n29352, n29353,
    n29354, n29355, n29356, n29357, n29358, n29359,
    n29360, n29361, n29362, n29363, n29364, n29365,
    n29366, n29367, n29368, n29369, n29370, n29371,
    n29372, n29373, n29374, n29375, n29376, n29377,
    n29378, n29379, n29380, n29381, n29382, n29383,
    n29384, n29385, n29386, n29387, n29388, n29389,
    n29390, n29391, n29392, n29393, n29394, n29395,
    n29396, n29397, n29398, n29399, n29400, n29401,
    n29402, n29403, n29404, n29405, n29406, n29407,
    n29408, n29409, n29410, n29411, n29412, n29413,
    n29414, n29415, n29416, n29417, n29418, n29419,
    n29420, n29421, n29422, n29423, n29424, n29425,
    n29426, n29427, n29428, n29429, n29430, n29431,
    n29432, n29433, n29434, n29435, n29436, n29437,
    n29438, n29439, n29440, n29441, n29442, n29443,
    n29444, n29445, n29446, n29447, n29448, n29449,
    n29450, n29451, n29452, n29453, n29454, n29455,
    n29456, n29457, n29458, n29459, n29460, n29461,
    n29462, n29463, n29464, n29465, n29466, n29467,
    n29468, n29469, n29470, n29471, n29472, n29473,
    n29474, n29475, n29476, n29477, n29478, n29479,
    n29480, n29481, n29482, n29483, n29484, n29485,
    n29486, n29487, n29488, n29489, n29490, n29491,
    n29492, n29493, n29494, n29495, n29496, n29497,
    n29498, n29499, n29500, n29501, n29502, n29503,
    n29504, n29505, n29506, n29507, n29508, n29509,
    n29510, n29511, n29512, n29513, n29514, n29515,
    n29516, n29517, n29518, n29519, n29520, n29521,
    n29522, n29523, n29524, n29525, n29526, n29527,
    n29528, n29529, n29530, n29531, n29532, n29533,
    n29534, n29535, n29536, n29537, n29538, n29539,
    n29540, n29541, n29542, n29543, n29544, n29545,
    n29546, n29547, n29548, n29549, n29550, n29551,
    n29552, n29553, n29554, n29555, n29556, n29557,
    n29558, n29559, n29560, n29561, n29562, n29563,
    n29564, n29565, n29566, n29567, n29568, n29569,
    n29570, n29571, n29572, n29573, n29574, n29575,
    n29576, n29577, n29578, n29579, n29580, n29581,
    n29582, n29583, n29584, n29585, n29586, n29587,
    n29588, n29589, n29590, n29591, n29592, n29593,
    n29594, n29595, n29596, n29597, n29598, n29599,
    n29600, n29601, n29602, n29603, n29604, n29605,
    n29606, n29607, n29608, n29609, n29610, n29611,
    n29612, n29613, n29614, n29615, n29616, n29617,
    n29618, n29619, n29620, n29621, n29622, n29623,
    n29624, n29625, n29626, n29627, n29628, n29629,
    n29630, n29631, n29632, n29633, n29634, n29635,
    n29636, n29637, n29638, n29639, n29640, n29641,
    n29642, n29643, n29644, n29645, n29646, n29647,
    n29648, n29649, n29650, n29651, n29652, n29653,
    n29654, n29655, n29656, n29657, n29658, n29659,
    n29660, n29661, n29662, n29663, n29664, n29665,
    n29666, n29667, n29668, n29669, n29670, n29671,
    n29672, n29673, n29674, n29675, n29676, n29677,
    n29678, n29679, n29680, n29681, n29682, n29683,
    n29684, n29685, n29686, n29687, n29688, n29689,
    n29690, n29691, n29692, n29693, n29694, n29695,
    n29696, n29697, n29698, n29699, n29700, n29701,
    n29702, n29703, n29704, n29705, n29706, n29707,
    n29708, n29709, n29710, n29711, n29712, n29713,
    n29714, n29715, n29716, n29717, n29718, n29719,
    n29720, n29721, n29722, n29723, n29724, n29725,
    n29726, n29727, n29728, n29729, n29730, n29731,
    n29732, n29733, n29734, n29735, n29736, n29737,
    n29738, n29739, n29740, n29741, n29742, n29743,
    n29744, n29745, n29746, n29747, n29748, n29749,
    n29750, n29751, n29752, n29753, n29754, n29755,
    n29756, n29757, n29758, n29759, n29760, n29761,
    n29762, n29763, n29764, n29765, n29766, n29767,
    n29768, n29769, n29770, n29771, n29772, n29773,
    n29774, n29775, n29776, n29777, n29778, n29779,
    n29780, n29781, n29782, n29783, n29784, n29785,
    n29786, n29787, n29788, n29789, n29790, n29791,
    n29792, n29793, n29794, n29795, n29796, n29797,
    n29798, n29799, n29800, n29801, n29802, n29803,
    n29804, n29805, n29806, n29807, n29808, n29809,
    n29810, n29811, n29812, n29813, n29814, n29815,
    n29816, n29817, n29818, n29819, n29820, n29821,
    n29822, n29823, n29824, n29825, n29826, n29827,
    n29828, n29829, n29830, n29831, n29832, n29833,
    n29834, n29835, n29836, n29837, n29838, n29839,
    n29840, n29841, n29842, n29843, n29844, n29845,
    n29846, n29847, n29848, n29849, n29850, n29851,
    n29852, n29853, n29854, n29855, n29856, n29857,
    n29858, n29859, n29860, n29861, n29862, n29863,
    n29864, n29865, n29866, n29867, n29868, n29869,
    n29870, n29871, n29872, n29873, n29874, n29875,
    n29876, n29877, n29878, n29879, n29880, n29881,
    n29882, n29883, n29884, n29885, n29886, n29887,
    n29888, n29889, n29890, n29891, n29892, n29893,
    n29894, n29895, n29896, n29897, n29898, n29899,
    n29900, n29901, n29902, n29903, n29904, n29905,
    n29906, n29907, n29908, n29909, n29910, n29911,
    n29912, n29913, n29914, n29915, n29916, n29917,
    n29918, n29919, n29920, n29921, n29922, n29923,
    n29924, n29925, n29926, n29927, n29928, n29929,
    n29930, n29931, n29932, n29933, n29934, n29935,
    n29936, n29937, n29938, n29939, n29940, n29941,
    n29942, n29943, n29944, n29945, n29946, n29947,
    n29948, n29949, n29950, n29951, n29952, n29953,
    n29954, n29955, n29956, n29957, n29958, n29959,
    n29960, n29961, n29962, n29963, n29964, n29965,
    n29966, n29967, n29968, n29969, n29970, n29971,
    n29972, n29973, n29974, n29975, n29976, n29977,
    n29978, n29979, n29980, n29981, n29982, n29983,
    n29984, n29985, n29986, n29987, n29988, n29989,
    n29990, n29991, n29992, n29993, n29994, n29995,
    n29996, n29997, n29998, n29999, n30000, n30001,
    n30002, n30003, n30004, n30005, n30006, n30007,
    n30008, n30009, n30010, n30011, n30012, n30013,
    n30014, n30015, n30016, n30017, n30018, n30019,
    n30020, n30021, n30022, n30023, n30024, n30025,
    n30026, n30027, n30028, n30029, n30030, n30031,
    n30032, n30033, n30034, n30035, n30036, n30037,
    n30038, n30039, n30040, n30041, n30042, n30043,
    n30044, n30045, n30046, n30047, n30048, n30049,
    n30050, n30051, n30052, n30053, n30054, n30055,
    n30056, n30057, n30058, n30059, n30060, n30061,
    n30062, n30063, n30064, n30065, n30066, n30067,
    n30068, n30069, n30070, n30071, n30072, n30073,
    n30074, n30075, n30076, n30077, n30078, n30079,
    n30080, n30081, n30082, n30083, n30084, n30085,
    n30086, n30087, n30088, n30089, n30090, n30091,
    n30092, n30093, n30094, n30095, n30096, n30097,
    n30098, n30099, n30100, n30101, n30102, n30103,
    n30104, n30105, n30106, n30107, n30108, n30109,
    n30110, n30111, n30112, n30113, n30114, n30115,
    n30116, n30117, n30118, n30119, n30120, n30121,
    n30122, n30123, n30124, n30125, n30126, n30127,
    n30128, n30129, n30130, n30131, n30132, n30133,
    n30134, n30135, n30136, n30137, n30138, n30139,
    n30140, n30141, n30142, n30143, n30144, n30145,
    n30146, n30147, n30148, n30149, n30150, n30151,
    n30152, n30153, n30154, n30155, n30156, n30157,
    n30158, n30159, n30160, n30161, n30162, n30163,
    n30164, n30165, n30166, n30167, n30168, n30169,
    n30170, n30171, n30172, n30173, n30174, n30175,
    n30176, n30177, n30178, n30179, n30180, n30181,
    n30182, n30183, n30184, n30185, n30186, n30187,
    n30188, n30189, n30190, n30191, n30192, n30193,
    n30194, n30195, n30196, n30197, n30198, n30199,
    n30200, n30201, n30202, n30203, n30204, n30205,
    n30206, n30207, n30208, n30209, n30210, n30211,
    n30212, n30213, n30214, n30215, n30216, n30217,
    n30218, n30219, n30220, n30221, n30222, n30223,
    n30224, n30225, n30226, n30227, n30228, n30229,
    n30230, n30231, n30232, n30233, n30234, n30235,
    n30236, n30237, n30238, n30239, n30240, n30241,
    n30242, n30243, n30244, n30245, n30246, n30247,
    n30248, n30249, n30250, n30251, n30252, n30253,
    n30254, n30255, n30256, n30257, n30258, n30259,
    n30260, n30261, n30262, n30263, n30264, n30265,
    n30266, n30267, n30268, n30269, n30270, n30271,
    n30272, n30273, n30274, n30275, n30276, n30277,
    n30278, n30279, n30280, n30281, n30282, n30283,
    n30284, n30285, n30286, n30287, n30288, n30289,
    n30290, n30291, n30292, n30293, n30294, n30295,
    n30296, n30297, n30298, n30299, n30300, n30301,
    n30302, n30303, n30304, n30305, n30306, n30307,
    n30308, n30309, n30310, n30311, n30312, n30313,
    n30314, n30315, n30316, n30317, n30318, n30319,
    n30320, n30321, n30322, n30323, n30324, n30325,
    n30326, n30327, n30328, n30329, n30330, n30331,
    n30332, n30333, n30334, n30335, n30336, n30337,
    n30338, n30339, n30340, n30341, n30342, n30343,
    n30344, n30345, n30346, n30347, n30348, n30349,
    n30350, n30351, n30352, n30353, n30354, n30355,
    n30356, n30357, n30358, n30359, n30360, n30361,
    n30362, n30363, n30364, n30365, n30366, n30367,
    n30368, n30369, n30370, n30371, n30372, n30373,
    n30374, n30375, n30376, n30377, n30378, n30379,
    n30380, n30381, n30382, n30383, n30384, n30385,
    n30386, n30387, n30388, n30389, n30390, n30391,
    n30392, n30393, n30394, n30395, n30396, n30397,
    n30398, n30399, n30400, n30401, n30402, n30403,
    n30404, n30405, n30406, n30407, n30408, n30409,
    n30410, n30411, n30412, n30413, n30414, n30415,
    n30416, n30417, n30418, n30419, n30420, n30421,
    n30422, n30423, n30424, n30425, n30426, n30427,
    n30428, n30429, n30430, n30431, n30432, n30433,
    n30434, n30435, n30436, n30437, n30438, n30439,
    n30440, n30441, n30442, n30443, n30444, n30445,
    n30446, n30447, n30448, n30449, n30450, n30451,
    n30452, n30453, n30454, n30455, n30456, n30457,
    n30458, n30459, n30460, n30461, n30462, n30463,
    n30464, n30465, n30466, n30467, n30468, n30469,
    n30470, n30471, n30472, n30473, n30474, n30475,
    n30476, n30477, n30478, n30479, n30480, n30481,
    n30482, n30483, n30484, n30485, n30486, n30487,
    n30488, n30489, n30490, n30491, n30492, n30493,
    n30494, n30495, n30496, n30497, n30498, n30499,
    n30500, n30501, n30502, n30503, n30504, n30505,
    n30506, n30507, n30508, n30509, n30510, n30511,
    n30512, n30513, n30514, n30515, n30516, n30517,
    n30518, n30519, n30520, n30521, n30522, n30523,
    n30524, n30525, n30526, n30527, n30528, n30529,
    n30530, n30531, n30532, n30533, n30534, n30535,
    n30536, n30537, n30538, n30539, n30540, n30541,
    n30542, n30543, n30544, n30545, n30546, n30547,
    n30548, n30549, n30550, n30551, n30552, n30553,
    n30554, n30555, n30556, n30557, n30558, n30559,
    n30560, n30561, n30562, n30563, n30564, n30565,
    n30566, n30567, n30568, n30570, n30571, n30572,
    n30573, n30574, n30575, n30576, n30577, n30578,
    n30579, n30580, n30581, n30582, n30583, n30584,
    n30585, n30586, n30587, n30588, n30589, n30590,
    n30591, n30592, n30593, n30594, n30595, n30596,
    n30597, n30598, n30599, n30600, n30601, n30602,
    n30603, n30604, n30605, n30606, n30607, n30608,
    n30609, n30610, n30611, n30612, n30613, n30614,
    n30615, n30616, n30617, n30618, n30619, n30620,
    n30621, n30622, n30623, n30624, n30625, n30626,
    n30627, n30628, n30629, n30630, n30631, n30632,
    n30633, n30634, n30635, n30636, n30637, n30638,
    n30639, n30640, n30641, n30642, n30643, n30644,
    n30645, n30646, n30647, n30648, n30649, n30650,
    n30651, n30652, n30653, n30654, n30655, n30656,
    n30657, n30658, n30659, n30660, n30661, n30662,
    n30663, n30664, n30665, n30666, n30667, n30668,
    n30669, n30670, n30671, n30672, n30673, n30674,
    n30675, n30676, n30677, n30678, n30679, n30680,
    n30681, n30682, n30683, n30684, n30685, n30686,
    n30687, n30688, n30689, n30690, n30691, n30692,
    n30693, n30694, n30695, n30696, n30697, n30698,
    n30699, n30700, n30701, n30702, n30703, n30704,
    n30705, n30706, n30707, n30708, n30709, n30710,
    n30711, n30712, n30713, n30714, n30715, n30716,
    n30717, n30718, n30719, n30720, n30721, n30722,
    n30723, n30724, n30725, n30726, n30727, n30728,
    n30729, n30730, n30731, n30732, n30733, n30734,
    n30735, n30736, n30737, n30738, n30739, n30740,
    n30741, n30742, n30743, n30744, n30745, n30746,
    n30747, n30748, n30749, n30750, n30751, n30752,
    n30753, n30754, n30755, n30756, n30757, n30758,
    n30759, n30760, n30761, n30762, n30763, n30764,
    n30765, n30766, n30767, n30768, n30769, n30770,
    n30771, n30772, n30773, n30774, n30775, n30776,
    n30777, n30778, n30779, n30780, n30781, n30782,
    n30783, n30784, n30785, n30786, n30787, n30788,
    n30789, n30790, n30791, n30792, n30793, n30794,
    n30795, n30796, n30797, n30798, n30799, n30800,
    n30801, n30802, n30803, n30804, n30805, n30806,
    n30807, n30808, n30809, n30810, n30811, n30812,
    n30813, n30814, n30815, n30816, n30817, n30818,
    n30819, n30820, n30821, n30822, n30823, n30824,
    n30825, n30826, n30827, n30828, n30829, n30830,
    n30831, n30832, n30833, n30834, n30835, n30836,
    n30837, n30838, n30839, n30840, n30841, n30842,
    n30843, n30844, n30845, n30846, n30847, n30848,
    n30849, n30850, n30851, n30852, n30853, n30854,
    n30855, n30856, n30857, n30858, n30859, n30860,
    n30861, n30862, n30863, n30864, n30865, n30866,
    n30867, n30868, n30869, n30870, n30871, n30872,
    n30873, n30874, n30875, n30876, n30877, n30878,
    n30879, n30880, n30881, n30882, n30883, n30884,
    n30885, n30886, n30887, n30888, n30889, n30890,
    n30891, n30892, n30893, n30894, n30895, n30896,
    n30897, n30898, n30899, n30900, n30901, n30902,
    n30903, n30904, n30905, n30906, n30907, n30909,
    n30910, n30912, n30913, n30914, n30915, n30916,
    n30917, n30918, n30919, n30920, n30921, n30922,
    n30923, n30924, n30925, n30926, n30927, n30928,
    n30929, n30930, n30931, n30932, n30933, n30934,
    n30935, n30936, n30937, n30938, n30939, n30940,
    n30941, n30942, n30943, n30944, n30945, n30946,
    n30947, n30948, n30949, n30950, n30951, n30952,
    n30953, n30954, n30955, n30956, n30957, n30958,
    n30959, n30960, n30961, n30962, n30963, n30964,
    n30965, n30966, n30967, n30968, n30969, n30970,
    n30971, n30972, n30973, n30974, n30975, n30976,
    n30977, n30978, n30979, n30980, n30981, n30982,
    n30983, n30984, n30985, n30986, n30987, n30988,
    n30989, n30990, n30991, n30992, n30993, n30994,
    n30995, n30996, n30997, n30998, n30999, n31000,
    n31001, n31002, n31003, n31004, n31005, n31006,
    n31007, n31008, n31009, n31010, n31011, n31012,
    n31013, n31014, n31015, n31016, n31017, n31018,
    n31019, n31020, n31021, n31022, n31023, n31024,
    n31025, n31026, n31027, n31028, n31029, n31030,
    n31031, n31032, n31033, n31034, n31035, n31036,
    n31037, n31038, n31039, n31040, n31041, n31042,
    n31043, n31044, n31045, n31046, n31047, n31048,
    n31049, n31050, n31051, n31052, n31053, n31054,
    n31055, n31056, n31057, n31058, n31059, n31060,
    n31061, n31062, n31063, n31064, n31065, n31066,
    n31067, n31068, n31069, n31070, n31071, n31072,
    n31073, n31074, n31075, n31076, n31077, n31078,
    n31079, n31080, n31081, n31082, n31083, n31084,
    n31085, n31086, n31087, n31088, n31089, n31090,
    n31091, n31092, n31093, n31094, n31095, n31096,
    n31097, n31098, n31099, n31100, n31101, n31102,
    n31103, n31104, n31105, n31106, n31107, n31108,
    n31109, n31110, n31111, n31112, n31113, n31114,
    n31115, n31116, n31117, n31118, n31119, n31120,
    n31121, n31122, n31123, n31124, n31125, n31126,
    n31127, n31128, n31129, n31130, n31131, n31132,
    n31133, n31134, n31135, n31136, n31137, n31138,
    n31139, n31140, n31141, n31142, n31143, n31144,
    n31145, n31146, n31147, n31148, n31149, n31150,
    n31151, n31152, n31153, n31154, n31155, n31156,
    n31157, n31158, n31159, n31160, n31161, n31162,
    n31163, n31164, n31165, n31166, n31167, n31168,
    n31169, n31170, n31171, n31172, n31173, n31174,
    n31175, n31176, n31177, n31178, n31179, n31180,
    n31181, n31182, n31183, n31184, n31185, n31186,
    n31187, n31188, n31189, n31190, n31191, n31192,
    n31193, n31194, n31195, n31196, n31197, n31198,
    n31199, n31200, n31201, n31202, n31203, n31204,
    n31205, n31206, n31207, n31208, n31209, n31210,
    n31211, n31212, n31213, n31214, n31215, n31216,
    n31217, n31218, n31219, n31220, n31221, n31222,
    n31223, n31224, n31225, n31226, n31227, n31228,
    n31229, n31230, n31231, n31232, n31233, n31234,
    n31235, n31236, n31237, n31238, n31239, n31240,
    n31241, n31242, n31243, n31244, n31245, n31246,
    n31247, n31248, n31249, n31250, n31251, n31252,
    n31253, n31254, n31255, n31256, n31257, n31258,
    n31259, n31260, n31261, n31262, n31263, n31264,
    n31265, n31266, n31267, n31268, n31269, n31270,
    n31271, n31272, n31273, n31274, n31275, n31276,
    n31277, n31278, n31279, n31280, n31281, n31282,
    n31283, n31284, n31285, n31286, n31287, n31288,
    n31289, n31290, n31291, n31292, n31293, n31294,
    n31295, n31296, n31297, n31298, n31299, n31300,
    n31301, n31302, n31303, n31304, n31305, n31306,
    n31307, n31308, n31309, n31310, n31311, n31312,
    n31313, n31314, n31315, n31316, n31317, n31318,
    n31319, n31320, n31321, n31322, n31323, n31324,
    n31325, n31326, n31327, n31328, n31329, n31330,
    n31331, n31332, n31333, n31334, n31335, n31336,
    n31337, n31338, n31339, n31340, n31341, n31342,
    n31343, n31344, n31345, n31346, n31347, n31348,
    n31349, n31350, n31351, n31352, n31353, n31354,
    n31355, n31356, n31357, n31358, n31359, n31360,
    n31361, n31362, n31363, n31364, n31365, n31366,
    n31367, n31368, n31369, n31370, n31371, n31372,
    n31373, n31374, n31375, n31376, n31377, n31378,
    n31379, n31380, n31381, n31382, n31383, n31384,
    n31385, n31386, n31387, n31388, n31389, n31390,
    n31391, n31392, n31393, n31394, n31395, n31396,
    n31397, n31398, n31399, n31400, n31401, n31402,
    n31403, n31404, n31405, n31406, n31407, n31408,
    n31409, n31410, n31411, n31412, n31413, n31414,
    n31415, n31416, n31417, n31418, n31419, n31420,
    n31421, n31422, n31423, n31424, n31425, n31426,
    n31427, n31428, n31429, n31430, n31431, n31432,
    n31433, n31434, n31435, n31436, n31437, n31438,
    n31439, n31440, n31441, n31442, n31443, n31444,
    n31445, n31446, n31447, n31448, n31449, n31450,
    n31451, n31452, n31453, n31454, n31455, n31456,
    n31457, n31458, n31459, n31460, n31461, n31462,
    n31463, n31464, n31465, n31466, n31467, n31468,
    n31469, n31470, n31471, n31472, n31473, n31474,
    n31475, n31476, n31477, n31478, n31479, n31480,
    n31481, n31482, n31483, n31484, n31485, n31486,
    n31487, n31488, n31489, n31490, n31491, n31492,
    n31493, n31494, n31495, n31496, n31497, n31498,
    n31499, n31500, n31501, n31502, n31503, n31504,
    n31505, n31506, n31507, n31508, n31509, n31510,
    n31511, n31512, n31513, n31514, n31515, n31516,
    n31517, n31518, n31519, n31520, n31521, n31522,
    n31523, n31524, n31525, n31526, n31527, n31528,
    n31529, n31530, n31531, n31532, n31533, n31534,
    n31535, n31536, n31537, n31538, n31539, n31540,
    n31541, n31542, n31543, n31544, n31545, n31546,
    n31547, n31548, n31549, n31550, n31551, n31552,
    n31553, n31554, n31555, n31556, n31557, n31558,
    n31559, n31560, n31561, n31562, n31563, n31564,
    n31565, n31566, n31567, n31568, n31569, n31570,
    n31571, n31572, n31573, n31574, n31575, n31576,
    n31577, n31578, n31579, n31580, n31581, n31582,
    n31583, n31584, n31585, n31586, n31587, n31588,
    n31589, n31590, n31591, n31592, n31593, n31594,
    n31595, n31596, n31597, n31598, n31599, n31600,
    n31601, n31602, n31603, n31604, n31605, n31606,
    n31607, n31608, n31609, n31610, n31611, n31612,
    n31613, n31614, n31615, n31616, n31617, n31618,
    n31619, n31620, n31621, n31622, n31623, n31624,
    n31625, n31626, n31627, n31628, n31629, n31630,
    n31631, n31632, n31633, n31634, n31635, n31636,
    n31637, n31638, n31639, n31640, n31641, n31642,
    n31643, n31644, n31645, n31646, n31647, n31648,
    n31649, n31650, n31651, n31652, n31653, n31654,
    n31655, n31656, n31657, n31658, n31659, n31660,
    n31661, n31662, n31663, n31664, n31665, n31666,
    n31667, n31668, n31669, n31670, n31671, n31672,
    n31673, n31674, n31675, n31676, n31677, n31678,
    n31679, n31680, n31681, n31682, n31683, n31684,
    n31685, n31686, n31687, n31688, n31689, n31690,
    n31691, n31692, n31693, n31694, n31695, n31696,
    n31697, n31698, n31699, n31700, n31701, n31702,
    n31703, n31704, n31705, n31706, n31707, n31708,
    n31709, n31710, n31711, n31712, n31713, n31714,
    n31715, n31716, n31717, n31718, n31719, n31720,
    n31721, n31722, n31723, n31724, n31725, n31726,
    n31727, n31728, n31729, n31730, n31731, n31732,
    n31733, n31734, n31735, n31736, n31737, n31738,
    n31739, n31740, n31741, n31742, n31743, n31744,
    n31745, n31746, n31747, n31748, n31749, n31750,
    n31751, n31752, n31753, n31754, n31755, n31756,
    n31757, n31758, n31759, n31760, n31761, n31762,
    n31763, n31764, n31765, n31766, n31767, n31768,
    n31769, n31770, n31771, n31772, n31773, n31774,
    n31775, n31776, n31777, n31778, n31779, n31780,
    n31781, n31782, n31783, n31784, n31785, n31786,
    n31787, n31788, n31789, n31790, n31791, n31792,
    n31793, n31794, n31795, n31796, n31797, n31798,
    n31799, n31800, n31801, n31802, n31803, n31804,
    n31805, n31806, n31807, n31808, n31809, n31810,
    n31811, n31812, n31813, n31814, n31815, n31816,
    n31817, n31818, n31819, n31820, n31821, n31822,
    n31823, n31824, n31825, n31826, n31827, n31828,
    n31829, n31830, n31831, n31832, n31833, n31834,
    n31835, n31836, n31837, n31838, n31839, n31840,
    n31841, n31842, n31843, n31844, n31845, n31846,
    n31847, n31848, n31849, n31850, n31851, n31852,
    n31853, n31854, n31855, n31856, n31857, n31858,
    n31859, n31860, n31861, n31862, n31863, n31864,
    n31865, n31866, n31867, n31868, n31869, n31870,
    n31871, n31872, n31873, n31874, n31875, n31876,
    n31877, n31878, n31879, n31880, n31881, n31882,
    n31883, n31884, n31885, n31886, n31887, n31888,
    n31889, n31890, n31891, n31892, n31893, n31894,
    n31895, n31896, n31897, n31898, n31899, n31900,
    n31901, n31902, n31903, n31904, n31905, n31906,
    n31907, n31908, n31909, n31910, n31911, n31912,
    n31913, n31914, n31915, n31916, n31917, n31918,
    n31919, n31920, n31921, n31922, n31923, n31924,
    n31925, n31926, n31927, n31928, n31929, n31930,
    n31931, n31932, n31933, n31934, n31935, n31936,
    n31937, n31938, n31939, n31940, n31941, n31942,
    n31943, n31944, n31945, n31946, n31947, n31948,
    n31949, n31950, n31951, n31952, n31953, n31954,
    n31955, n31956, n31957, n31958, n31959, n31960,
    n31961, n31962, n31963, n31964, n31965, n31966,
    n31967, n31968, n31969, n31970, n31971, n31972,
    n31973, n31974, n31975, n31976, n31977, n31978,
    n31979, n31980, n31981, n31982, n31983, n31984,
    n31985, n31986, n31987, n31988, n31989, n31990,
    n31991, n31992, n31993, n31994, n31995, n31996,
    n31997, n31998, n31999, n32000, n32001, n32002,
    n32003, n32004, n32005, n32006, n32007, n32008,
    n32009, n32010, n32011, n32012, n32013, n32014,
    n32015, n32016, n32017, n32018, n32019, n32020,
    n32021, n32022, n32023, n32024, n32025, n32026,
    n32027, n32028, n32029, n32030, n32031, n32032,
    n32033, n32034, n32035, n32036, n32037, n32038,
    n32039, n32040, n32041, n32042, n32043, n32044,
    n32045, n32046, n32047, n32048, n32049, n32050,
    n32051, n32052, n32053, n32054, n32055, n32056,
    n32057, n32058, n32059, n32060, n32061, n32062,
    n32063, n32064, n32065, n32066, n32067, n32068,
    n32069, n32070, n32071, n32072, n32073, n32074,
    n32075, n32076, n32077, n32078, n32079, n32080,
    n32081, n32082, n32083, n32084, n32085, n32086,
    n32087, n32088, n32089, n32090, n32091, n32092,
    n32093, n32094, n32095, n32096, n32097, n32098,
    n32099, n32100, n32101, n32102, n32103, n32104,
    n32105, n32106, n32107, n32108, n32109, n32110,
    n32111, n32112, n32113, n32114, n32115, n32116,
    n32117, n32118, n32119, n32120, n32121, n32122,
    n32123, n32124, n32125, n32126, n32127, n32128,
    n32129, n32130, n32131, n32132, n32133, n32134,
    n32135, n32136, n32137, n32138, n32139, n32140,
    n32141, n32142, n32143, n32144, n32145, n32146,
    n32147, n32148, n32149, n32150, n32151, n32152,
    n32153, n32154, n32155, n32156, n32157, n32158,
    n32159, n32160, n32161, n32162, n32163, n32164,
    n32165, n32166, n32167, n32168, n32169, n32170,
    n32171, n32172, n32173, n32174, n32175, n32176,
    n32177, n32178, n32179, n32180, n32181, n32182,
    n32183, n32184, n32185, n32186, n32187, n32188,
    n32189, n32190, n32191, n32192, n32193, n32194,
    n32195, n32196, n32197, n32198, n32199, n32200,
    n32201, n32202, n32203, n32204, n32205, n32206,
    n32207, n32208, n32209, n32210, n32211, n32212,
    n32213, n32214, n32215, n32216, n32217, n32218,
    n32219, n32220, n32221, n32222, n32223, n32224,
    n32225, n32226, n32227, n32228, n32229, n32230,
    n32231, n32232, n32233, n32234, n32235, n32236,
    n32237, n32238, n32239, n32240, n32241, n32242,
    n32243, n32244, n32245, n32246, n32247, n32248,
    n32249, n32250, n32251, n32252, n32253, n32254,
    n32255, n32256, n32257, n32258, n32259, n32260,
    n32261, n32262, n32263, n32264, n32265, n32266,
    n32267, n32268, n32269, n32270, n32271, n32272,
    n32273, n32274, n32275, n32276, n32277, n32278,
    n32279, n32280, n32281, n32282, n32283, n32284,
    n32285, n32286, n32287, n32288, n32289, n32290,
    n32291, n32292, n32293, n32294, n32295, n32296,
    n32297, n32298, n32299, n32300, n32301, n32303,
    n32304, n32305, n32306, n32307, n32308, n32309,
    n32310, n32311, n32312, n32313, n32314, n32315,
    n32316, n32317, n32318, n32319, n32320, n32321,
    n32322, n32323, n32324, n32325, n32326, n32327,
    n32328, n32329, n32330, n32331, n32332, n32333,
    n32334, n32335, n32336, n32337, n32338, n32339,
    n32340, n32341, n32342, n32343, n32344, n32345,
    n32346, n32347, n32348, n32349, n32350, n32351,
    n32352, n32353, n32354, n32355, n32356, n32357,
    n32358, n32359, n32360, n32361, n32362, n32363,
    n32364, n32365, n32366, n32367, n32368, n32369,
    n32370, n32371, n32372, n32373, n32374, n32375,
    n32376, n32377, n32378, n32379, n32380, n32381,
    n32382, n32383, n32384, n32385, n32386, n32387,
    n32388, n32389, n32390, n32391, n32392, n32393,
    n32394, n32395, n32396, n32397, n32398, n32399,
    n32400, n32401, n32402, n32403, n32404, n32405,
    n32406, n32407, n32408, n32409, n32410, n32411,
    n32412, n32413, n32414, n32415, n32416, n32417,
    n32418, n32419, n32420, n32421, n32422, n32423,
    n32424, n32425, n32426, n32427, n32428, n32429,
    n32430, n32431, n32432, n32433, n32434, n32435,
    n32436, n32437, n32438, n32439, n32440, n32441,
    n32442, n32443, n32444, n32445, n32446, n32447,
    n32448, n32449, n32450, n32451, n32452, n32453,
    n32454, n32455, n32456, n32457, n32458, n32459,
    n32460, n32461, n32462, n32463, n32464, n32465,
    n32466, n32467, n32468, n32469, n32470, n32471,
    n32472, n32473, n32474, n32475, n32476, n32477,
    n32478, n32479, n32480, n32481, n32482, n32483,
    n32484, n32485, n32486, n32487, n32488, n32489,
    n32490, n32491, n32492, n32493, n32494, n32495,
    n32496, n32497, n32498, n32499, n32500, n32501,
    n32502, n32503, n32504, n32505, n32506, n32507,
    n32508, n32509, n32510, n32511, n32512, n32513,
    n32514, n32515, n32516, n32517, n32518, n32519,
    n32520, n32521, n32522, n32523, n32524, n32525,
    n32526, n32527, n32528, n32529, n32530, n32531,
    n32532, n32533, n32534, n32535, n32536, n32537,
    n32538, n32539, n32540, n32541, n32542, n32543,
    n32544, n32545, n32546, n32547, n32548, n32549,
    n32550, n32551, n32552, n32553, n32554, n32555,
    n32556, n32557, n32558, n32559, n32560, n32561,
    n32562, n32563, n32564, n32565, n32566, n32567,
    n32568, n32569, n32570, n32571, n32572, n32573,
    n32574, n32575, n32576, n32577, n32578, n32579,
    n32580, n32581, n32582, n32583, n32584, n32585,
    n32586, n32587, n32588, n32589, n32590, n32591,
    n32592, n32593, n32594, n32595, n32596, n32597,
    n32598, n32599, n32600, n32601, n32602, n32603,
    n32604, n32605, n32606, n32607, n32608, n32609,
    n32610, n32611, n32612, n32613, n32614, n32615,
    n32616, n32617, n32618, n32619, n32620, n32621,
    n32622, n32623, n32624, n32625, n32626, n32627,
    n32628, n32629, n32630, n32631, n32632, n32633,
    n32634, n32635, n32636, n32637, n32638, n32639,
    n32640, n32641, n32642, n32643, n32644, n32645,
    n32646, n32647, n32648, n32649, n32650, n32651,
    n32652, n32653, n32654, n32655, n32656, n32657,
    n32658, n32659, n32660, n32661, n32662, n32663,
    n32664, n32665, n32666, n32667, n32668, n32669,
    n32670, n32671, n32672, n32673, n32674, n32675,
    n32676, n32677, n32678, n32679, n32680, n32681,
    n32682, n32683, n32684, n32685, n32686, n32687,
    n32688, n32689, n32690, n32691, n32692, n32693,
    n32694, n32695, n32696, n32697, n32698, n32699,
    n32700, n32701, n32702, n32703, n32704, n32705,
    n32706, n32707, n32708, n32709, n32710, n32711,
    n32712, n32713, n32714, n32715, n32716, n32717,
    n32718, n32719, n32720, n32721, n32722, n32723,
    n32724, n32725, n32726, n32727, n32728, n32729,
    n32730, n32731, n32732, n32733, n32734, n32735,
    n32736, n32737, n32738, n32739, n32740, n32741,
    n32742, n32743, n32744, n32745, n32746, n32747,
    n32748, n32749, n32750, n32751, n32752, n32753,
    n32754, n32755, n32756, n32757, n32758, n32759,
    n32760, n32761, n32762, n32763, n32764, n32765,
    n32766, n32767, n32768, n32769, n32770, n32771,
    n32772, n32773, n32774, n32775, n32776, n32777,
    n32778, n32779, n32780, n32781, n32782, n32783,
    n32784, n32785, n32786, n32787, n32788, n32789,
    n32790, n32791, n32792, n32793, n32794, n32795,
    n32796, n32797, n32798, n32799, n32800, n32801,
    n32802, n32803, n32804, n32805, n32806, n32807,
    n32808, n32809, n32810, n32811, n32812, n32813,
    n32814, n32815, n32816, n32817, n32818, n32819,
    n32820, n32821, n32822, n32823, n32824, n32825,
    n32826, n32827, n32828, n32829, n32830, n32831,
    n32832, n32833, n32834, n32835, n32836, n32837,
    n32838, n32839, n32840, n32841, n32842, n32843,
    n32844, n32845, n32846, n32847, n32848, n32849,
    n32850, n32851, n32852, n32853, n32854, n32855,
    n32856, n32857, n32858, n32859, n32860, n32861,
    n32862, n32863, n32864, n32865, n32866, n32867,
    n32868, n32869, n32870, n32871, n32872, n32873,
    n32874, n32875, n32876, n32877, n32878, n32879,
    n32880, n32881, n32882, n32883, n32884, n32885,
    n32886, n32887, n32888, n32889, n32890, n32891,
    n32892, n32893, n32894, n32895, n32896, n32897,
    n32898, n32899, n32900, n32901, n32902, n32903,
    n32904, n32905, n32906, n32907, n32908, n32909,
    n32910, n32911, n32912, n32913, n32914, n32915,
    n32916, n32917, n32918, n32919, n32920, n32921,
    n32922, n32923, n32924, n32925, n32926, n32927,
    n32928, n32929, n32930, n32931, n32932, n32933,
    n32934, n32935, n32936, n32937, n32938, n32939,
    n32940, n32941, n32942, n32943, n32944, n32945,
    n32946, n32947, n32948, n32949, n32950, n32951,
    n32952, n32953, n32954, n32955, n32956, n32957,
    n32958, n32959, n32960, n32961, n32962, n32963,
    n32964, n32965, n32966, n32967, n32968, n32969,
    n32970, n32971, n32972, n32973, n32974, n32975,
    n32976, n32977, n32978, n32979, n32980, n32981,
    n32982, n32983, n32984, n32985, n32986, n32987,
    n32988, n32989, n32990, n32991, n32992, n32993,
    n32994, n32995, n32996, n32997, n32998, n32999,
    n33000, n33001, n33002, n33003, n33004, n33005,
    n33006, n33007, n33008, n33009, n33010, n33011,
    n33012, n33013, n33014, n33015, n33016, n33017,
    n33018, n33019, n33020, n33021, n33022, n33023,
    n33024, n33025, n33026, n33027, n33028, n33029,
    n33030, n33031, n33032, n33033, n33034, n33035,
    n33036, n33037, n33038, n33039, n33040, n33041,
    n33042, n33043, n33044, n33045, n33046, n33047,
    n33048, n33049, n33050, n33051, n33052, n33053,
    n33054, n33055, n33056, n33057, n33058, n33059,
    n33060, n33061, n33062, n33063, n33064, n33065,
    n33066, n33067, n33068, n33069, n33070, n33071,
    n33072, n33073, n33074, n33075, n33076, n33077,
    n33078, n33079, n33080, n33081, n33082, n33083,
    n33084, n33085, n33086, n33087, n33088, n33089,
    n33090, n33091, n33092, n33093, n33094, n33095,
    n33096, n33097, n33098, n33099, n33100, n33101,
    n33102, n33103, n33104, n33105, n33106, n33107,
    n33108, n33109, n33110, n33111, n33112, n33113,
    n33114, n33115, n33116, n33117, n33118, n33119,
    n33120, n33121, n33122, n33123, n33124, n33125,
    n33126, n33127, n33128, n33129, n33130, n33131,
    n33132, n33133, n33134, n33135, n33136, n33137,
    n33138, n33139, n33140, n33141, n33142, n33143,
    n33144, n33145, n33146, n33147, n33148, n33149,
    n33150, n33151, n33152, n33153, n33154, n33155,
    n33156, n33157, n33158, n33159, n33160, n33161,
    n33162, n33163, n33164, n33165, n33166, n33167,
    n33168, n33169, n33170, n33171, n33172, n33173,
    n33174, n33175, n33176, n33177, n33178, n33179,
    n33180, n33181, n33182, n33183, n33184, n33185,
    n33186, n33187, n33188, n33189, n33190, n33191,
    n33192, n33193, n33194, n33195, n33196, n33197,
    n33198, n33199, n33200, n33201, n33202, n33203,
    n33204, n33205, n33206, n33207, n33208, n33209,
    n33210, n33211, n33212, n33213, n33214, n33215,
    n33216, n33217, n33218, n33219, n33220, n33221,
    n33222, n33223, n33224, n33225, n33226, n33227,
    n33228, n33229, n33230, n33231, n33232, n33233,
    n33234, n33235, n33236, n33237, n33238, n33239,
    n33240, n33241, n33242, n33243, n33244, n33245,
    n33246, n33247, n33248, n33249, n33250, n33251,
    n33252, n33253, n33254, n33255, n33256, n33257,
    n33258, n33259, n33260, n33261, n33262, n33263,
    n33264, n33265, n33266, n33267, n33268, n33269,
    n33270, n33271, n33272, n33273, n33274, n33275,
    n33276, n33277, n33278, n33279, n33280, n33281,
    n33282, n33283, n33284, n33285, n33286, n33287,
    n33288, n33289, n33290, n33291, n33292, n33293,
    n33294, n33295, n33296, n33297, n33298, n33299,
    n33300, n33301, n33302, n33303, n33304, n33305,
    n33306, n33307, n33308, n33309, n33310, n33311,
    n33312, n33313, n33314, n33315, n33316, n33317,
    n33318, n33319, n33320, n33321, n33322, n33323,
    n33324, n33325, n33326, n33327, n33328, n33329,
    n33330, n33331, n33332, n33333, n33334, n33335,
    n33336, n33337, n33338, n33339, n33340, n33341,
    n33342, n33343, n33344, n33345, n33346, n33347,
    n33348, n33349, n33350, n33351, n33352, n33353,
    n33354, n33355, n33356, n33357, n33358, n33359,
    n33360, n33361, n33362, n33363, n33364, n33365,
    n33366, n33367, n33368, n33369, n33370, n33371,
    n33372, n33373, n33374, n33375, n33376, n33377,
    n33378, n33379, n33380, n33381, n33382, n33383,
    n33384, n33385, n33386, n33387, n33388, n33389,
    n33390, n33391, n33392, n33393, n33394, n33395,
    n33396, n33397, n33398, n33399, n33400, n33401,
    n33402, n33403, n33404, n33405, n33406, n33407,
    n33408, n33409, n33410, n33411, n33412, n33413,
    n33414, n33415, n33416, n33417, n33418, n33419,
    n33420, n33421, n33422, n33423, n33424, n33425,
    n33426, n33427, n33428, n33429, n33430, n33431,
    n33432, n33433, n33434, n33435, n33436, n33437,
    n33438, n33439, n33440, n33441, n33442, n33443,
    n33444, n33445, n33446, n33447, n33448, n33449,
    n33450, n33451, n33452, n33453, n33454, n33455,
    n33456, n33457, n33458, n33459, n33460, n33461,
    n33462, n33463, n33464, n33465, n33466, n33467,
    n33468, n33469, n33470, n33471, n33472, n33473,
    n33474, n33475, n33476, n33477, n33478, n33479,
    n33480, n33481, n33482, n33483, n33484, n33485,
    n33486, n33487, n33488, n33489, n33490, n33491,
    n33492, n33493, n33494, n33495, n33496, n33497,
    n33498, n33499, n33500, n33501, n33502, n33503,
    n33504, n33505, n33506, n33507, n33508, n33509,
    n33510, n33511, n33512, n33513, n33514, n33515,
    n33516, n33517, n33518, n33519, n33520, n33521,
    n33522, n33523, n33524, n33525, n33526, n33527,
    n33528, n33529, n33530, n33531, n33532, n33533,
    n33534, n33535, n33536, n33537, n33538, n33539,
    n33540, n33541, n33542, n33543, n33544, n33545,
    n33546, n33547, n33548, n33549, n33550, n33551,
    n33552, n33553, n33554, n33555, n33556, n33557,
    n33558, n33559, n33560, n33561, n33562, n33563,
    n33564, n33565, n33566, n33567, n33568, n33569,
    n33570, n33571, n33572, n33573, n33574, n33575,
    n33576, n33577, n33578, n33579, n33580, n33581,
    n33582, n33583, n33584, n33585, n33586, n33587,
    n33588, n33589, n33590, n33591, n33592, n33593,
    n33594, n33595, n33596, n33597, n33598, n33599,
    n33600, n33601, n33602, n33603, n33604, n33605,
    n33606, n33607, n33608, n33609, n33610, n33611,
    n33612, n33613, n33614, n33615, n33616, n33617,
    n33618, n33619, n33620, n33621, n33622, n33623,
    n33624, n33625, n33626, n33627, n33628, n33629,
    n33630, n33631, n33632, n33633, n33634, n33635,
    n33636, n33637, n33638, n33639, n33640, n33641,
    n33642, n33643, n33644, n33645, n33646, n33647,
    n33648, n33649, n33650, n33651, n33652, n33653,
    n33654, n33655, n33656, n33657, n33658, n33659,
    n33660, n33661, n33662, n33663, n33664, n33665,
    n33666, n33667, n33668, n33669, n33670, n33671,
    n33672, n33673, n33674, n33675, n33676, n33677,
    n33678, n33679, n33680, n33681, n33682, n33683,
    n33684, n33685, n33686, n33687, n33688, n33689,
    n33690, n33691, n33692, n33693, n33694, n33695,
    n33696, n33697, n33698, n33699, n33700, n33701,
    n33702, n33703, n33704, n33705, n33706, n33707,
    n33708, n33709, n33710, n33711, n33712, n33713,
    n33714, n33715, n33716, n33717, n33718, n33719,
    n33720, n33721, n33722, n33723, n33724, n33725,
    n33726, n33727, n33728, n33729, n33730, n33731,
    n33732, n33733, n33734, n33735, n33736, n33737,
    n33738, n33739, n33740, n33741, n33742, n33743,
    n33744, n33745, n33746, n33747, n33748, n33749,
    n33750, n33751, n33752, n33753, n33754, n33755,
    n33756, n33757, n33758, n33759, n33760, n33761,
    n33762, n33763, n33764, n33765, n33766, n33767,
    n33768, n33769, n33770, n33771, n33772, n33773,
    n33774, n33775, n33776, n33777, n33778, n33779,
    n33780, n33781, n33782, n33783, n33784, n33785,
    n33786, n33787, n33788, n33789, n33790, n33791,
    n33792, n33793, n33794, n33795, n33796, n33797,
    n33798, n33799, n33800, n33801, n33802, n33803,
    n33804, n33805, n33806, n33807, n33808, n33809,
    n33810, n33811, n33812, n33813, n33814, n33815,
    n33816, n33817, n33818, n33819, n33820, n33821,
    n33822, n33823, n33824, n33825, n33826, n33827,
    n33828, n33829, n33830, n33831, n33832, n33833,
    n33834, n33835, n33836, n33837, n33838, n33839,
    n33840, n33841, n33842, n33843, n33844, n33846,
    n33847, n33848, n33849, n33850, n33851, n33852,
    n33853, n33854, n33855, n33856, n33857, n33858,
    n33859, n33860, n33861, n33862, n33863, n33864,
    n33865, n33866, n33867, n33868, n33869, n33870,
    n33871, n33872, n33873, n33874, n33875, n33876,
    n33877, n33878, n33879, n33880, n33881, n33882,
    n33883, n33884, n33885, n33886, n33887, n33888,
    n33889, n33890, n33891, n33892, n33893, n33894,
    n33895, n33896, n33897, n33898, n33899, n33900,
    n33901, n33902, n33903, n33904, n33905, n33906,
    n33907, n33908, n33909, n33910, n33911, n33912,
    n33913, n33914, n33915, n33916, n33917, n33918,
    n33919, n33920, n33921, n33922, n33923, n33924,
    n33925, n33926, n33927, n33928, n33929, n33930,
    n33931, n33932, n33933, n33934, n33935, n33936,
    n33937, n33938, n33939, n33940, n33941, n33942,
    n33943, n33944, n33945, n33946, n33947, n33948,
    n33949, n33950, n33951, n33952, n33953, n33954,
    n33955, n33956, n33957, n33958, n33959, n33960,
    n33961, n33962, n33963, n33964, n33965, n33966,
    n33967, n33968, n33969, n33970, n33971, n33972,
    n33973, n33974, n33975, n33976, n33977, n33978,
    n33979, n33980, n33981, n33982, n33983, n33984,
    n33985, n33986, n33987, n33988, n33989, n33990,
    n33991, n33992, n33993, n33994, n33995, n33996,
    n33997, n33998, n33999, n34000, n34001, n34002,
    n34003, n34004, n34005, n34006, n34007, n34008,
    n34009, n34010, n34011, n34012, n34013, n34014,
    n34015, n34016, n34017, n34018, n34019, n34020,
    n34021, n34022, n34023, n34024, n34025, n34026,
    n34027, n34028, n34029, n34030, n34031, n34032,
    n34033, n34034, n34035, n34036, n34037, n34038,
    n34039, n34040, n34041, n34042, n34043, n34044,
    n34045, n34046, n34047, n34048, n34049, n34050,
    n34051, n34053, n34054, n34055, n34056, n34057,
    n34058, n34059, n34060, n34061, n34062, n34063,
    n34064, n34065, n34066, n34067, n34068, n34069,
    n34070, n34071, n34072, n34073, n34074, n34075,
    n34076, n34077, n34078, n34079, n34080, n34081,
    n34082, n34083, n34084, n34085, n34086, n34087,
    n34088, n34089, n34090, n34091, n34092, n34093,
    n34094, n34095, n34096, n34097, n34098, n34099,
    n34100, n34101, n34102, n34103, n34104, n34105,
    n34106, n34107, n34108, n34109, n34110, n34111,
    n34112, n34113, n34114, n34115, n34116, n34117,
    n34118, n34119, n34120, n34121, n34122, n34123,
    n34124, n34125, n34126, n34127, n34128, n34129,
    n34130, n34131, n34132, n34133, n34134, n34135,
    n34136, n34137, n34138, n34139, n34140, n34141,
    n34142, n34143, n34144, n34145, n34146, n34147,
    n34148, n34149, n34150, n34151, n34152, n34153,
    n34154, n34155, n34156, n34157, n34158, n34159,
    n34160, n34161, n34162, n34163, n34164, n34165,
    n34166, n34167, n34168, n34169, n34170, n34171,
    n34172, n34173, n34174, n34175, n34176, n34177,
    n34178, n34179, n34180, n34181, n34182, n34183,
    n34184, n34185, n34186, n34187, n34188, n34189,
    n34190, n34191, n34192, n34193, n34194, n34195,
    n34196, n34197, n34198, n34199, n34200, n34201,
    n34202, n34203, n34204, n34205, n34206, n34208,
    n34209, n34210, n34211, n34212, n34213, n34214,
    n34215, n34216, n34217, n34218, n34219, n34220,
    n34221, n34222, n34223, n34224, n34225, n34226,
    n34227, n34228, n34229, n34230, n34231, n34232,
    n34233, n34234, n34235, n34236, n34237, n34238,
    n34239, n34240, n34241, n34242, n34243, n34244,
    n34245, n34246, n34247, n34248, n34249, n34250,
    n34251, n34252, n34253, n34254, n34255, n34256,
    n34257, n34258, n34259, n34260, n34261, n34262,
    n34263, n34264, n34265, n34266, n34267, n34268,
    n34269, n34270, n34271, n34272, n34273, n34274,
    n34275, n34276, n34277, n34278, n34279, n34280,
    n34281, n34282, n34283, n34284, n34285, n34286,
    n34287, n34288, n34289, n34290, n34291, n34292,
    n34293, n34294, n34295, n34296, n34297, n34298,
    n34299, n34300, n34301, n34302, n34303, n34304,
    n34305, n34306, n34307, n34308, n34309, n34310,
    n34311, n34312, n34313, n34314, n34315, n34316,
    n34317, n34318, n34319, n34320, n34321, n34322,
    n34323, n34324, n34325, n34326, n34327, n34328,
    n34329, n34330, n34331, n34332, n34333, n34334,
    n34335, n34337, n34338, n34339, n34340, n34341,
    n34342, n34343, n34344, n34345, n34346, n34347,
    n34348, n34349, n34350, n34351, n34352, n34353,
    n34354, n34355, n34356, n34357, n34358, n34359,
    n34360, n34361, n34362, n34363, n34364, n34365,
    n34366, n34367, n34368, n34369, n34370, n34371,
    n34372, n34373, n34374, n34375, n34376, n34377,
    n34378, n34379, n34380, n34381, n34382, n34383,
    n34384, n34385, n34386, n34387, n34388, n34389,
    n34390, n34391, n34392, n34393, n34394, n34395,
    n34396, n34397, n34398, n34399, n34400, n34401,
    n34402, n34403, n34404, n34405, n34406, n34407,
    n34408, n34409, n34410, n34411, n34412, n34413,
    n34414, n34415, n34416, n34417, n34418, n34419,
    n34420, n34421, n34422, n34423, n34424, n34425,
    n34426, n34427, n34428, n34429, n34430, n34431,
    n34432, n34433, n34434, n34435, n34436, n34437,
    n34438, n34439, n34440, n34441, n34442, n34443,
    n34444, n34445, n34446, n34447, n34448, n34449,
    n34450, n34451, n34452, n34453, n34454, n34455,
    n34456, n34457, n34458, n34459, n34460, n34461,
    n34462, n34463, n34465, n34466, n34467, n34468,
    n34469, n34470, n34471, n34472, n34473, n34474,
    n34475, n34476, n34477, n34478, n34479, n34480,
    n34481, n34482, n34483, n34484, n34485, n34486,
    n34487, n34488, n34489, n34490, n34491, n34492,
    n34493, n34494, n34495, n34496, n34497, n34498,
    n34499, n34500, n34501, n34502, n34503, n34504,
    n34505, n34506, n34507, n34508, n34509, n34510,
    n34511, n34512, n34513, n34514, n34515, n34516,
    n34517, n34518, n34519, n34520, n34521, n34522,
    n34523, n34524, n34525, n34526, n34527, n34528,
    n34529, n34530, n34531, n34532, n34533, n34534,
    n34535, n34536, n34537, n34538, n34539, n34540,
    n34541, n34542, n34543, n34544, n34545, n34546,
    n34547, n34548, n34549, n34550, n34551, n34552,
    n34553, n34554, n34555, n34556, n34557, n34558,
    n34559, n34561, n34562, n34563, n34564, n34565,
    n34566, n34567, n34568, n34569, n34570, n34571,
    n34572, n34573, n34574, n34575, n34576, n34577,
    n34578, n34579, n34580, n34581, n34582, n34583,
    n34584, n34585, n34586, n34587, n34588, n34589,
    n34590, n34591, n34592, n34593, n34594, n34595,
    n34596, n34597, n34598, n34599, n34600, n34601,
    n34602, n34603, n34604, n34605, n34606, n34607,
    n34608, n34609, n34610, n34611, n34612, n34613,
    n34614, n34615, n34616, n34617, n34618, n34619,
    n34620, n34621, n34622, n34623, n34624, n34625,
    n34626, n34627, n34628, n34629, n34630, n34631,
    n34632, n34633, n34634, n34635, n34636, n34637,
    n34638, n34639, n34640, n34641, n34642, n34643,
    n34644, n34645, n34646, n34647, n34648, n34649,
    n34650, n34651, n34652, n34653, n34654, n34655,
    n34657, n34658, n34659, n34660, n34661, n34662,
    n34663, n34664, n34665, n34666, n34667, n34668,
    n34669, n34670, n34671, n34672, n34673, n34674,
    n34675, n34676, n34677, n34678, n34679, n34680,
    n34681, n34682, n34683, n34684, n34685, n34686,
    n34687, n34688, n34689, n34690, n34691, n34692,
    n34693, n34694, n34695, n34696, n34697, n34698,
    n34699, n34700, n34701, n34702, n34703, n34704,
    n34705, n34706, n34707, n34708, n34709, n34710,
    n34711, n34712, n34713, n34714, n34715, n34716,
    n34717, n34718, n34719, n34720, n34721, n34722,
    n34723, n34724, n34725, n34726, n34727, n34728,
    n34729, n34730, n34731, n34732, n34733, n34734,
    n34735, n34736, n34737, n34738, n34739, n34740,
    n34741, n34742, n34743, n34744, n34745, n34746,
    n34747, n34748, n34749, n34750, n34751, n34753,
    n34754, n34755, n34756, n34757, n34758, n34759,
    n34760, n34761, n34762, n34763, n34764, n34765,
    n34766, n34767, n34768, n34769, n34770, n34771,
    n34772, n34773, n34774, n34775, n34776, n34777,
    n34778, n34779, n34780, n34781, n34782, n34783,
    n34784, n34785, n34786, n34787, n34788, n34789,
    n34790, n34791, n34792, n34793, n34794, n34795,
    n34796, n34797, n34798, n34799, n34800, n34801,
    n34802, n34803, n34804, n34805, n34806, n34807,
    n34808, n34809, n34810, n34811, n34812, n34813,
    n34814, n34815, n34816, n34817, n34818, n34819,
    n34820, n34821, n34822, n34823, n34824, n34825,
    n34826, n34827, n34828, n34829, n34830, n34831,
    n34832, n34833, n34834, n34835, n34836, n34837,
    n34838, n34839, n34840, n34841, n34842, n34843,
    n34844, n34845, n34846, n34847, n34849, n34850,
    n34851, n34852, n34853, n34854, n34855, n34856,
    n34857, n34858, n34859, n34860, n34861, n34862,
    n34863, n34864, n34865, n34866, n34867, n34868,
    n34869, n34870, n34871, n34872, n34873, n34874,
    n34875, n34876, n34877, n34878, n34879, n34880,
    n34881, n34882, n34883, n34884, n34885, n34886,
    n34887, n34888, n34889, n34890, n34891, n34892,
    n34893, n34894, n34895, n34896, n34897, n34898,
    n34899, n34900, n34901, n34902, n34903, n34904,
    n34905, n34906, n34907, n34908, n34909, n34910,
    n34911, n34912, n34913, n34914, n34915, n34916,
    n34917, n34918, n34919, n34920, n34921, n34922,
    n34923, n34924, n34925, n34926, n34927, n34928,
    n34929, n34930, n34931, n34932, n34933, n34934,
    n34935, n34936, n34937, n34938, n34939, n34941,
    n34942, n34943, n34944, n34945, n34946, n34947,
    n34948, n34949, n34950, n34951, n34952, n34953,
    n34954, n34955, n34956, n34957, n34958, n34959,
    n34960, n34961, n34962, n34963, n34964, n34965,
    n34966, n34967, n34968, n34969, n34970, n34971,
    n34972, n34973, n34974, n34975, n34976, n34977,
    n34978, n34979, n34980, n34981, n34982, n34983,
    n34984, n34985, n34986, n34987, n34988, n34989,
    n34990, n34991, n34992, n34993, n34994, n34995,
    n34996, n34997, n34998, n34999, n35000, n35001,
    n35002, n35003, n35004, n35005, n35006, n35007,
    n35008, n35009, n35010, n35011, n35012, n35013,
    n35014, n35015, n35016, n35017, n35018, n35019,
    n35020, n35021, n35022, n35023, n35024, n35025,
    n35026, n35027, n35028, n35029, n35030, n35031,
    n35032, n35033, n35034, n35035, n35036, n35037,
    n35038, n35039, n35040, n35041, n35042, n35043,
    n35044, n35045, n35046, n35047, n35048, n35049,
    n35050, n35051, n35052, n35053, n35054, n35055,
    n35056, n35057, n35058, n35059, n35060, n35061,
    n35062, n35063, n35064, n35065, n35066, n35067,
    n35068, n35069, n35070, n35071, n35072, n35073,
    n35074, n35075, n35076, n35077, n35078, n35079,
    n35080, n35081, n35082, n35083, n35084, n35085,
    n35086, n35087, n35088, n35089, n35090, n35091,
    n35092, n35093, n35094, n35095, n35096, n35097,
    n35098, n35099, n35100, n35101, n35102, n35103,
    n35104, n35105, n35106, n35107, n35108, n35109,
    n35110, n35111, n35112, n35113, n35114, n35115,
    n35116, n35117, n35118, n35119, n35120, n35121,
    n35122, n35123, n35124, n35125, n35126, n35127,
    n35128, n35129, n35131, n35132, n35133, n35134,
    n35135, n35136, n35137, n35138, n35139, n35140,
    n35141, n35142, n35143, n35144, n35145, n35146,
    n35147, n35148, n35149, n35150, n35151, n35152,
    n35153, n35154, n35155, n35156, n35157, n35158,
    n35159, n35160, n35161, n35162, n35163, n35164,
    n35165, n35166, n35167, n35168, n35169, n35170,
    n35171, n35172, n35173, n35174, n35175, n35176,
    n35177, n35178, n35179, n35180, n35181, n35182,
    n35183, n35184, n35185, n35186, n35187, n35188,
    n35189, n35190, n35191, n35192, n35193, n35194,
    n35195, n35197, n35198, n35199, n35200, n35201,
    n35202, n35203, n35204, n35205, n35206, n35207,
    n35208, n35209, n35210, n35211, n35212, n35213,
    n35214, n35215, n35216, n35217, n35218, n35219,
    n35220, n35221, n35222, n35223, n35224, n35225,
    n35226, n35227, n35228, n35229, n35230, n35231,
    n35232, n35233, n35234, n35235, n35236, n35237,
    n35238, n35239, n35240, n35241, n35242, n35243,
    n35244, n35245, n35246, n35247, n35248, n35249,
    n35250, n35251, n35252, n35253, n35254, n35255,
    n35256, n35257, n35258, n35259, n35260, n35261,
    n35262, n35263, n35264, n35265, n35266, n35267,
    n35268, n35269, n35270, n35271, n35272, n35273,
    n35274, n35275, n35276, n35277, n35278, n35279,
    n35280, n35281, n35282, n35283, n35284, n35285,
    n35286, n35287, n35288, n35289, n35290, n35291,
    n35292, n35293, n35294, n35295, n35296, n35297,
    n35298, n35299, n35300, n35301, n35302, n35303,
    n35304, n35305, n35306, n35307, n35308, n35309,
    n35310, n35311, n35312, n35313, n35314, n35315,
    n35316, n35317, n35318, n35319, n35320, n35321,
    n35322, n35323, n35324, n35325, n35326, n35327,
    n35328, n35329, n35330, n35331, n35332, n35333,
    n35334, n35335, n35336, n35337, n35338, n35339,
    n35340, n35341, n35342, n35343, n35344, n35345,
    n35346, n35347, n35348, n35349, n35350, n35351,
    n35352, n35353, n35354, n35355, n35356, n35357,
    n35358, n35359, n35360, n35361, n35362, n35363,
    n35364, n35365, n35366, n35367, n35368, n35369,
    n35370, n35371, n35372, n35373, n35374, n35375,
    n35376, n35377, n35378, n35379, n35380, n35381,
    n35382, n35383, n35384, n35385, n35386, n35387,
    n35388, n35389, n35390, n35391, n35392, n35393,
    n35394, n35395, n35396, n35397, n35398, n35399,
    n35400, n35401, n35402, n35403, n35404, n35405,
    n35406, n35407, n35408, n35409, n35410, n35411,
    n35412, n35413, n35414, n35415, n35416, n35417,
    n35418, n35419, n35420, n35421, n35422, n35423,
    n35424, n35425, n35426, n35427, n35428, n35429,
    n35430, n35431, n35432, n35433, n35434, n35435,
    n35436, n35437, n35438, n35439, n35440, n35441,
    n35442, n35443, n35444, n35445, n35446, n35447,
    n35448, n35449, n35450, n35451, n35452, n35453,
    n35454, n35455, n35456, n35457, n35458, n35459,
    n35460, n35461, n35462, n35463, n35464, n35465,
    n35466, n35467, n35468, n35469, n35470, n35471,
    n35472, n35473, n35474, n35475, n35476, n35477,
    n35478, n35479, n35480, n35481, n35482, n35483,
    n35484, n35485, n35486, n35487, n35488, n35489,
    n35490, n35491, n35492, n35493, n35494, n35495,
    n35496, n35497, n35498, n35499, n35500, n35501,
    n35502, n35503, n35504, n35505, n35506, n35507,
    n35508, n35509, n35510, n35511, n35512, n35513,
    n35514, n35515, n35516, n35517, n35518, n35519,
    n35520, n35521, n35522, n35523, n35524, n35525,
    n35526, n35527, n35528, n35529, n35530, n35531,
    n35532, n35533, n35534, n35535, n35536, n35537,
    n35538, n35539, n35540, n35541, n35542, n35543,
    n35544, n35545, n35546, n35547, n35548, n35549,
    n35550, n35551, n35552, n35553, n35554, n35555,
    n35556, n35557, n35558, n35559, n35560, n35561,
    n35562, n35563, n35564, n35565, n35566, n35567,
    n35568, n35569, n35570, n35571, n35572, n35573,
    n35574, n35575, n35576, n35577, n35578, n35579,
    n35580, n35581, n35582, n35583, n35584, n35585,
    n35586, n35587, n35588, n35589, n35590, n35591,
    n35592, n35593, n35594, n35595, n35596, n35597,
    n35598, n35599, n35600, n35601, n35602, n35603,
    n35604, n35605, n35606, n35607, n35608, n35609,
    n35610, n35611, n35612, n35613, n35614, n35615,
    n35616, n35617, n35618, n35619, n35620, n35621,
    n35622, n35623, n35624, n35625, n35626, n35627,
    n35628, n35629, n35630, n35631, n35632, n35633,
    n35634, n35635, n35636, n35637, n35638, n35639,
    n35640, n35641, n35642, n35643, n35644, n35645,
    n35646, n35647, n35648, n35649, n35650, n35651,
    n35652, n35653, n35654, n35655, n35656, n35657,
    n35658, n35659, n35660, n35661, n35662, n35663,
    n35664, n35665, n35666, n35667, n35668, n35669,
    n35670, n35671, n35672, n35673, n35674, n35675,
    n35676, n35677, n35678, n35679, n35680, n35681,
    n35682, n35683, n35684, n35685, n35686, n35687,
    n35688, n35689, n35690, n35691, n35692, n35693,
    n35694, n35695, n35696, n35697, n35698, n35699,
    n35700, n35701, n35702, n35703, n35704, n35705,
    n35706, n35707, n35708, n35709, n35710, n35711,
    n35712, n35713, n35714, n35715, n35716, n35717,
    n35718, n35719, n35720, n35721, n35722, n35723,
    n35724, n35725, n35726, n35727, n35728, n35729,
    n35730, n35731, n35732, n35733, n35734, n35735,
    n35736, n35737, n35738, n35739, n35741, n35742,
    n35743, n35744, n35745, n35746, n35747, n35748,
    n35749, n35750, n35751, n35752, n35753, n35754,
    n35755, n35756, n35757, n35758, n35759, n35760,
    n35761, n35762, n35763, n35764, n35765, n35766,
    n35767, n35768, n35769, n35770, n35771, n35772,
    n35773, n35774, n35775, n35776, n35777, n35778,
    n35779, n35780, n35781, n35782, n35783, n35784,
    n35785, n35786, n35787, n35788, n35789, n35790,
    n35791, n35792, n35793, n35794, n35795, n35796,
    n35797, n35798, n35799, n35800, n35801, n35802,
    n35803, n35804, n35805, n35806, n35807, n35808,
    n35809, n35810, n35811, n35812, n35813, n35814,
    n35815, n35816, n35817, n35818, n35819, n35820,
    n35821, n35822, n35823, n35824, n35825, n35826,
    n35827, n35828, n35829, n35830, n35831, n35832,
    n35833, n35834, n35835, n35836, n35837, n35838,
    n35839, n35840, n35841, n35842, n35843, n35844,
    n35845, n35846, n35847, n35848, n35849, n35850,
    n35851, n35852, n35853, n35854, n35855, n35856,
    n35857, n35858, n35859, n35860, n35861, n35862,
    n35863, n35864, n35865, n35866, n35867, n35868,
    n35869, n35870, n35871, n35872, n35873, n35874,
    n35875, n35876, n35877, n35878, n35879, n35880,
    n35881, n35882, n35883, n35884, n35885, n35886,
    n35887, n35888, n35889, n35890, n35891, n35892,
    n35893, n35894, n35895, n35896, n35897, n35898,
    n35899, n35901, n35902, n35903, n35904, n35905,
    n35906, n35907, n35908, n35909, n35910, n35911,
    n35912, n35913, n35914, n35915, n35916, n35917,
    n35918, n35919, n35920, n35921, n35922, n35923,
    n35924, n35925, n35926, n35927, n35928, n35929,
    n35930, n35931, n35932, n35933, n35934, n35935,
    n35936, n35937, n35938, n35939, n35940, n35941,
    n35942, n35943, n35944, n35945, n35946, n35947,
    n35948, n35949, n35950, n35951, n35952, n35953,
    n35954, n35955, n35956, n35957, n35958, n35959,
    n35960, n35961, n35962, n35963, n35964, n35965,
    n35966, n35967, n35968, n35969, n35970, n35971,
    n35972, n35973, n35974, n35975, n35977, n35978,
    n35979, n35980, n35981, n35982, n35983, n35984,
    n35985, n35986, n35987, n35988, n35989, n35990,
    n35991, n35992, n35993, n35994, n35995, n35996,
    n35997, n35998, n35999, n36000, n36001, n36002,
    n36003, n36004, n36005, n36006, n36007, n36008,
    n36009, n36010, n36011, n36012, n36013, n36014,
    n36015, n36016, n36017, n36018, n36019, n36020,
    n36021, n36022, n36023, n36024, n36025, n36026,
    n36027, n36028, n36029, n36030, n36031, n36032,
    n36033, n36034, n36035, n36036, n36037, n36038,
    n36039, n36040, n36041, n36042, n36043, n36044,
    n36045, n36046, n36047, n36048, n36049, n36050,
    n36051, n36052, n36053, n36054, n36055, n36056,
    n36057, n36058, n36059, n36060, n36061, n36062,
    n36063, n36064, n36065, n36066, n36067, n36068,
    n36070, n36071, n36072, n36073, n36074, n36075,
    n36076, n36077, n36078, n36079, n36080, n36081,
    n36082, n36083, n36084, n36085, n36086, n36087,
    n36088, n36089, n36090, n36091, n36092, n36093,
    n36094, n36095, n36096, n36097, n36098, n36099,
    n36100, n36101, n36102, n36103, n36104, n36105,
    n36106, n36107, n36108, n36109, n36110, n36111,
    n36112, n36113, n36114, n36115, n36116, n36117,
    n36118, n36119, n36120, n36121, n36122, n36123,
    n36124, n36125, n36126, n36127, n36128, n36129,
    n36130, n36131, n36132, n36133, n36134, n36135,
    n36136, n36137, n36138, n36139, n36140, n36141,
    n36142, n36143, n36144, n36145, n36146, n36147,
    n36148, n36149, n36150, n36151, n36152, n36153,
    n36154, n36155, n36156, n36157, n36158, n36159,
    n36160, n36161, n36162, n36163, n36164, n36165,
    n36166, n36167, n36168, n36169, n36170, n36171,
    n36172, n36173, n36174, n36175, n36176, n36177,
    n36178, n36179, n36180, n36181, n36182, n36183,
    n36184, n36185, n36186, n36187, n36188, n36189,
    n36190, n36191, n36192, n36193, n36194, n36195,
    n36196, n36197, n36198, n36199, n36200, n36201,
    n36202, n36203, n36204, n36205, n36206, n36207,
    n36208, n36209, n36210, n36211, n36212, n36213,
    n36214, n36215, n36216, n36217, n36218, n36219,
    n36220, n36221, n36222, n36223, n36224, n36225,
    n36226, n36227, n36228, n36229, n36230, n36231,
    n36232, n36233, n36234, n36235, n36236, n36237,
    n36238, n36239, n36240, n36241, n36242, n36243,
    n36244, n36245, n36246, n36247, n36248, n36249,
    n36250, n36251, n36252, n36253, n36254, n36255,
    n36256, n36257, n36258, n36259, n36260, n36261,
    n36262, n36263, n36264, n36265, n36266, n36267,
    n36268, n36269, n36270, n36271, n36272, n36273,
    n36274, n36275, n36276, n36277, n36278, n36279,
    n36280, n36281, n36282, n36283, n36284, n36285,
    n36286, n36287, n36288, n36289, n36290, n36291,
    n36292, n36293, n36294, n36295, n36296, n36297,
    n36298, n36299, n36300, n36301, n36302, n36303,
    n36304, n36305, n36306, n36307, n36308, n36309,
    n36310, n36311, n36312, n36313, n36314, n36315,
    n36316, n36317, n36318, n36319, n36320, n36321,
    n36322, n36323, n36324, n36325, n36326, n36327,
    n36328, n36329, n36330, n36331, n36332, n36333,
    n36334, n36335, n36336, n36337, n36338, n36339,
    n36340, n36342, n36343, n36344, n36345, n36346,
    n36347, n36348, n36349, n36350, n36351, n36352,
    n36353, n36354, n36355, n36356, n36357, n36358,
    n36359, n36360, n36361, n36362, n36363, n36364,
    n36365, n36366, n36367, n36368, n36369, n36370,
    n36371, n36372, n36373, n36374, n36375, n36376,
    n36377, n36378, n36379, n36380, n36381, n36382,
    n36383, n36384, n36385, n36386, n36387, n36388,
    n36389, n36390, n36391, n36393, n36394, n36395,
    n36396, n36397, n36398, n36399, n36400, n36401,
    n36402, n36403, n36404, n36405, n36406, n36407,
    n36408, n36409, n36410, n36411, n36412, n36413,
    n36414, n36415, n36416, n36417, n36418, n36419,
    n36420, n36421, n36422, n36423, n36424, n36426,
    n36427, n36428, n36429, n36430, n36431, n36432,
    n36433, n36434, n36435, n36436, n36437, n36438,
    n36439, n36440, n36441, n36442, n36443, n36444,
    n36445, n36446, n36447, n36448, n36449, n36450,
    n36451, n36452, n36453, n36454, n36455, n36456,
    n36457, n36458, n36459, n36460, n36461, n36462,
    n36463, n36464, n36465, n36466, n36467, n36468,
    n36469, n36470, n36471, n36472, n36473, n36474,
    n36475, n36476, n36477, n36478, n36479, n36480,
    n36481, n36482, n36483, n36484, n36485, n36486,
    n36487, n36488, n36489, n36490, n36491, n36492,
    n36493, n36494, n36495, n36496, n36497, n36498,
    n36499, n36500, n36501, n36502, n36503, n36504,
    n36505, n36506, n36507, n36508, n36509, n36510,
    n36511, n36512, n36514, n36515, n36516, n36517,
    n36518, n36519, n36520, n36521, n36522, n36523,
    n36524, n36525, n36526, n36527, n36528, n36529,
    n36530, n36531, n36532, n36533, n36534, n36535,
    n36536, n36537, n36538, n36539, n36540, n36541,
    n36542, n36543, n36544, n36545, n36546, n36547,
    n36548, n36549, n36550, n36551, n36552, n36553,
    n36554, n36555, n36556, n36557, n36558, n36559,
    n36560, n36561, n36562, n36563, n36564, n36565,
    n36566, n36567, n36568, n36569, n36570, n36571,
    n36572, n36573, n36574, n36575, n36576, n36577,
    n36578, n36579, n36580, n36581, n36582, n36583,
    n36584, n36585, n36586, n36587, n36588, n36590,
    n36591, n36592, n36593, n36594, n36595, n36596,
    n36597, n36598, n36599, n36600, n36601, n36602,
    n36603, n36604, n36605, n36606, n36607, n36608,
    n36609, n36610, n36611, n36612, n36613, n36614,
    n36615, n36616, n36617, n36618, n36619, n36620,
    n36621, n36622, n36623, n36624, n36625, n36626,
    n36627, n36628, n36629, n36630, n36631, n36632,
    n36633, n36634, n36635, n36636, n36637, n36638,
    n36639, n36640, n36641, n36642, n36643, n36644,
    n36645, n36646, n36647, n36648, n36649, n36650,
    n36651, n36652, n36653, n36654, n36655, n36656,
    n36657, n36658, n36659, n36660, n36661, n36662,
    n36663, n36664, n36666, n36667, n36668, n36669,
    n36670, n36671, n36672, n36673, n36674, n36675,
    n36676, n36677, n36678, n36679, n36680, n36681,
    n36682, n36683, n36684, n36685, n36686, n36687,
    n36688, n36689, n36690, n36691, n36692, n36693,
    n36694, n36695, n36696, n36697, n36698, n36699,
    n36700, n36701, n36702, n36703, n36704, n36705,
    n36706, n36707, n36708, n36709, n36710, n36711,
    n36712, n36713, n36714, n36715, n36716, n36717,
    n36718, n36719, n36720, n36721, n36722, n36723,
    n36724, n36725, n36726, n36727, n36728, n36729,
    n36730, n36731, n36732, n36733, n36734, n36735,
    n36736, n36737, n36738, n36739, n36740, n36741,
    n36742, n36743, n36744, n36745, n36746, n36747,
    n36748, n36749, n36751, n36752, n36753, n36754,
    n36755, n36756, n36757, n36758, n36759, n36760,
    n36761, n36762, n36763, n36764, n36765, n36766,
    n36767, n36768, n36769, n36770, n36771, n36772,
    n36773, n36774, n36775, n36776, n36777, n36778,
    n36779, n36780, n36781, n36782, n36783, n36784,
    n36785, n36786, n36787, n36788, n36789, n36790,
    n36791, n36792, n36793, n36794, n36795, n36796,
    n36797, n36798, n36799, n36800, n36801, n36802,
    n36803, n36804, n36805, n36806, n36807, n36808,
    n36809, n36810, n36811, n36812, n36813, n36814,
    n36815, n36816, n36817, n36818, n36819, n36820,
    n36821, n36822, n36823, n36824, n36825, n36826,
    n36827, n36828, n36829, n36830, n36831, n36832,
    n36833, n36834, n36835, n36836, n36837, n36838,
    n36839, n36840, n36841, n36842, n36843, n36844,
    n36845, n36846, n36847, n36848, n36849, n36850,
    n36851, n36852, n36853, n36854, n36855, n36856,
    n36857, n36858, n36859, n36860, n36861, n36862,
    n36863, n36864, n36865, n36866, n36867, n36868,
    n36869, n36870, n36871, n36872, n36873, n36874,
    n36875, n36876, n36877, n36878, n36879, n36880,
    n36881, n36882, n36883, n36884, n36885, n36886,
    n36887, n36888, n36889, n36890, n36891, n36892,
    n36893, n36894, n36895, n36896, n36897, n36898,
    n36899, n36900, n36901, n36902, n36903, n36904,
    n36905, n36906, n36907, n36908, n36909, n36910,
    n36911, n36912, n36913, n36914, n36915, n36916,
    n36917, n36918, n36919, n36920, n36921, n36922,
    n36923, n36924, n36925, n36926, n36927, n36928,
    n36929, n36930, n36931, n36932, n36933, n36934,
    n36935, n36936, n36937, n36938, n36939, n36940,
    n36941, n36942, n36943, n36944, n36946, n36947,
    n36948, n36949, n36950, n36951, n36952, n36953,
    n36954, n36955, n36956, n36957, n36958, n36959,
    n36960, n36961, n36962, n36963, n36964, n36965,
    n36966, n36967, n36968, n36969, n36970, n36971,
    n36972, n36973, n36974, n36975, n36976, n36977,
    n36978, n36979, n36980, n36981, n36982, n36983,
    n36984, n36985, n36986, n36987, n36988, n36989,
    n36990, n36991, n36992, n36993, n36994, n36995,
    n36996, n36997, n36998, n36999, n37000, n37001,
    n37002, n37003, n37004, n37005, n37006, n37007,
    n37008, n37009, n37010, n37011, n37012, n37013,
    n37014, n37015, n37016, n37017, n37018, n37019,
    n37020, n37021, n37022, n37023, n37024, n37025,
    n37026, n37027, n37028, n37029, n37031, n37032,
    n37033, n37034, n37035, n37036, n37037, n37038,
    n37039, n37040, n37041, n37042, n37043, n37044,
    n37045, n37046, n37047, n37048, n37049, n37050,
    n37051, n37052, n37053, n37054, n37055, n37056,
    n37057, n37058, n37059, n37060, n37061, n37062,
    n37063, n37064, n37065, n37066, n37067, n37068,
    n37069, n37070, n37071, n37072, n37073, n37074,
    n37076, n37077, n37078, n37079, n37080, n37081,
    n37082, n37083, n37084, n37085, n37086, n37087,
    n37088, n37089, n37090, n37091, n37092, n37093,
    n37094, n37095, n37096, n37097, n37098, n37099,
    n37100, n37101, n37102, n37103, n37104, n37105,
    n37106, n37107, n37108, n37109, n37110, n37111,
    n37112, n37113, n37114, n37115, n37116, n37117,
    n37118, n37119, n37121, n37122, n37123, n37124,
    n37125, n37126, n37127, n37128, n37129, n37130,
    n37131, n37132, n37133, n37134, n37135, n37136,
    n37137, n37138, n37139, n37140, n37141, n37142,
    n37143, n37144, n37145, n37146, n37147, n37148,
    n37149, n37150, n37151, n37152, n37153, n37154,
    n37155, n37156, n37157, n37158, n37159, n37160,
    n37161, n37162, n37163, n37164, n37165, n37166,
    n37167, n37168, n37169, n37170, n37171, n37172,
    n37173, n37174, n37175, n37176, n37177, n37178,
    n37179, n37180, n37181, n37182, n37183, n37184,
    n37185, n37186, n37187, n37188, n37189, n37190,
    n37191, n37192, n37193, n37194, n37195, n37196,
    n37197, n37198, n37199, n37200, n37201, n37202,
    n37203, n37204, n37205, n37206, n37207, n37208,
    n37209, n37210, n37211, n37212, n37213, n37214,
    n37215, n37216, n37217, n37218, n37219, n37220,
    n37221, n37222, n37223, n37224, n37225, n37226,
    n37227, n37228, n37229, n37230, n37231, n37232,
    n37233, n37234, n37235, n37236, n37237, n37238,
    n37239, n37240, n37241, n37242, n37243, n37244,
    n37245, n37246, n37247, n37248, n37249, n37250,
    n37251, n37252, n37253, n37254, n37255, n37256,
    n37257, n37258, n37259, n37260, n37261, n37262,
    n37263, n37264, n37265, n37266, n37267, n37268,
    n37269, n37270, n37271, n37272, n37273, n37274,
    n37275, n37276, n37277, n37278, n37279, n37280,
    n37281, n37282, n37283, n37284, n37286, n37287,
    n37288, n37289, n37290, n37291, n37292, n37293,
    n37294, n37295, n37296, n37297, n37298, n37299,
    n37300, n37301, n37302, n37303, n37304, n37305,
    n37306, n37307, n37308, n37309, n37310, n37311,
    n37312, n37313, n37314, n37315, n37316, n37317,
    n37318, n37319, n37320, n37321, n37322, n37323,
    n37324, n37325, n37326, n37327, n37328, n37329,
    n37330, n37331, n37332, n37333, n37334, n37335,
    n37336, n37337, n37338, n37339, n37340, n37341,
    n37342, n37343, n37344, n37345, n37346, n37347,
    n37348, n37349, n37350, n37351, n37352, n37353,
    n37354, n37355, n37356, n37357, n37358, n37359,
    n37360, n37361, n37362, n37363, n37364, n37365,
    n37366, n37367, n37368, n37369, n37370, n37371,
    n37372, n37373, n37374, n37375, n37376, n37377,
    n37378, n37379, n37380, n37381, n37382, n37383,
    n37384, n37385, n37386, n37387, n37388, n37389,
    n37390, n37391, n37392, n37393, n37394, n37395,
    n37396, n37397, n37398, n37399, n37400, n37401,
    n37402, n37403, n37404, n37405, n37406, n37407,
    n37408, n37409, n37410, n37411, n37412, n37413,
    n37414, n37415, n37416, n37417, n37418, n37419,
    n37420, n37421, n37422, n37423, n37424, n37425,
    n37426, n37427, n37428, n37429, n37430, n37431,
    n37432, n37433, n37434, n37435, n37436, n37437,
    n37438, n37439, n37440, n37441, n37442, n37443,
    n37444, n37445, n37446, n37447, n37448, n37449,
    n37450, n37451, n37452, n37453, n37454, n37455,
    n37456, n37457, n37458, n37459, n37460, n37461,
    n37462, n37463, n37464, n37465, n37466, n37467,
    n37468, n37469, n37470, n37471, n37472, n37473,
    n37474, n37475, n37476, n37477, n37478, n37479,
    n37480, n37481, n37482, n37483, n37484, n37485,
    n37486, n37487, n37488, n37489, n37490, n37491,
    n37492, n37493, n37494, n37495, n37496, n37497,
    n37498, n37499, n37500, n37501, n37502, n37503,
    n37504, n37505, n37506, n37507, n37508, n37509,
    n37510, n37511, n37512, n37513, n37514, n37515,
    n37516, n37517, n37518, n37519, n37520, n37521,
    n37522, n37523, n37524, n37525, n37526, n37527,
    n37528, n37529, n37530, n37531, n37532, n37533,
    n37534, n37535, n37536, n37537, n37538, n37539,
    n37540, n37541, n37542, n37543, n37544, n37545,
    n37546, n37547, n37548, n37549, n37550, n37551,
    n37552, n37553, n37554, n37555, n37556, n37557,
    n37558, n37559, n37560, n37561, n37562, n37563,
    n37564, n37565, n37566, n37567, n37568, n37569,
    n37570, n37571, n37572, n37573, n37574, n37575,
    n37576, n37577, n37578, n37579, n37580, n37581,
    n37582, n37583, n37584, n37585, n37586, n37587,
    n37588, n37589, n37590, n37591, n37592, n37593,
    n37594, n37595, n37596, n37597, n37598, n37599,
    n37600, n37601, n37602, n37603, n37604, n37605,
    n37606, n37607, n37608, n37609, n37610, n37611,
    n37612, n37613, n37614, n37615, n37616, n37617,
    n37618, n37619, n37620, n37621, n37622, n37623,
    n37624, n37625, n37626, n37627, n37628, n37629,
    n37630, n37631, n37632, n37633, n37634, n37635,
    n37636, n37637, n37638, n37639, n37640, n37641,
    n37642, n37643, n37644, n37645, n37646, n37647,
    n37648, n37649, n37650, n37651, n37652, n37653,
    n37654, n37655, n37656, n37657, n37658, n37659,
    n37660, n37661, n37662, n37663, n37664, n37665,
    n37666, n37667, n37668, n37669, n37670, n37671,
    n37672, n37673, n37674, n37675, n37676, n37677,
    n37678, n37679, n37680, n37681, n37682, n37683,
    n37684, n37685, n37686, n37687, n37688, n37689,
    n37690, n37691, n37692, n37693, n37694, n37695,
    n37696, n37697, n37698, n37699, n37700, n37701,
    n37702, n37703, n37704, n37705, n37706, n37707,
    n37708, n37709, n37710, n37711, n37712, n37713,
    n37714, n37715, n37716, n37717, n37718, n37719,
    n37720, n37721, n37722, n37723, n37724, n37725,
    n37726, n37727, n37728, n37729, n37730, n37731,
    n37732, n37733, n37734, n37735, n37736, n37737,
    n37738, n37739, n37740, n37741, n37742, n37743,
    n37744, n37745, n37746, n37747, n37748, n37749,
    n37750, n37751, n37752, n37753, n37754, n37755,
    n37756, n37757, n37758, n37759, n37760, n37761,
    n37762, n37763, n37764, n37765, n37766, n37767,
    n37768, n37769, n37770, n37771, n37772, n37773,
    n37774, n37775, n37776, n37777, n37778, n37779,
    n37780, n37781, n37782, n37783, n37784, n37785,
    n37786, n37787, n37788, n37789, n37790, n37791,
    n37792, n37793, n37794, n37795, n37796, n37797,
    n37798, n37799, n37800, n37801, n37802, n37803,
    n37804, n37805, n37806, n37807, n37808, n37809,
    n37810, n37811, n37812, n37813, n37814, n37815,
    n37816, n37817, n37818, n37819, n37820, n37821,
    n37822, n37823, n37824, n37825, n37826, n37827,
    n37828, n37829, n37830, n37831, n37832, n37833,
    n37834, n37835, n37836, n37837, n37838, n37839,
    n37840, n37841, n37842, n37843, n37844, n37845,
    n37846, n37847, n37848, n37849, n37850, n37851,
    n37852, n37853, n37854, n37855, n37856, n37857,
    n37858, n37859, n37860, n37861, n37862, n37863,
    n37864, n37865, n37866, n37867, n37868, n37869,
    n37870, n37871, n37872, n37873, n37874, n37875,
    n37877, n37878, n37879, n37880, n37881, n37882,
    n37883, n37884, n37885, n37886, n37887, n37888,
    n37889, n37891, n37892, n37893, n37894, n37895,
    n37896, n37897, n37898, n37899, n37900, n37901,
    n37902, n37903, n37904, n37905, n37906, n37907,
    n37908, n37909, n37910, n37911, n37912, n37913,
    n37914, n37915, n37916, n37917, n37918, n37919,
    n37920, n37921, n37922, n37923, n37924, n37925,
    n37926, n37927, n37928, n37929, n37930, n37931,
    n37932, n37933, n37934, n37935, n37936, n37937,
    n37938, n37939, n37940, n37941, n37942, n37943,
    n37944, n37945, n37946, n37947, n37948, n37949,
    n37950, n37951, n37952, n37953, n37954, n37955,
    n37956, n37957, n37958, n37959, n37960, n37961,
    n37962, n37963, n37964, n37965, n37966, n37967,
    n37968, n37969, n37970, n37971, n37972, n37973,
    n37974, n37975, n37976, n37977, n37978, n37979,
    n37980, n37981, n37982, n37983, n37984, n37985,
    n37986, n37987, n37988, n37989, n37990, n37991,
    n37992, n37993, n37994, n37995, n37996, n37997,
    n37998, n37999, n38000, n38001, n38002, n38003,
    n38004, n38005, n38006, n38007, n38008, n38009,
    n38010, n38011, n38012, n38013, n38014, n38015,
    n38016, n38017, n38018, n38019, n38020, n38021,
    n38022, n38023, n38024, n38025, n38026, n38027,
    n38028, n38029, n38030, n38031, n38032, n38033,
    n38034, n38035, n38036, n38037, n38038, n38039,
    n38040, n38041, n38042, n38043, n38044, n38045,
    n38046, n38047, n38048, n38049, n38050, n38051,
    n38052, n38053, n38054, n38055, n38056, n38057,
    n38058, n38059, n38060, n38061, n38062, n38063,
    n38064, n38065, n38066, n38067, n38068, n38069,
    n38070, n38071, n38072, n38073, n38074, n38075,
    n38076, n38077, n38078, n38079, n38080, n38081,
    n38082, n38083, n38084, n38085, n38086, n38087,
    n38088, n38089, n38090, n38091, n38092, n38093,
    n38094, n38095, n38096, n38097, n38098, n38099,
    n38100, n38101, n38102, n38103, n38104, n38105,
    n38106, n38107, n38108, n38109, n38110, n38111,
    n38112, n38113, n38114, n38115, n38116, n38117,
    n38118, n38119, n38120, n38121, n38122, n38123,
    n38124, n38125, n38126, n38127, n38128, n38129,
    n38130, n38131, n38132, n38133, n38134, n38135,
    n38136, n38137, n38138, n38139, n38140, n38141,
    n38142, n38143, n38144, n38145, n38146, n38147,
    n38148, n38149, n38150, n38151, n38152, n38153,
    n38154, n38155, n38156, n38157, n38158, n38159,
    n38160, n38161, n38162, n38163, n38164, n38165,
    n38166, n38167, n38168, n38169, n38170, n38171,
    n38172, n38173, n38174, n38175, n38176, n38178,
    n38179, n38180, n38181, n38182, n38183, n38184,
    n38185, n38186, n38187, n38188, n38189, n38190,
    n38191, n38192, n38193, n38194, n38195, n38196,
    n38197, n38198, n38199, n38200, n38201, n38202,
    n38203, n38204, n38205, n38206, n38207, n38208,
    n38209, n38210, n38212, n38213, n38214, n38215,
    n38216, n38217, n38218, n38219, n38220, n38221,
    n38222, n38223, n38224, n38225, n38226, n38227,
    n38228, n38229, n38230, n38231, n38232, n38233,
    n38234, n38235, n38236, n38237, n38238, n38239,
    n38240, n38241, n38242, n38243, n38244, n38245,
    n38246, n38247, n38248, n38249, n38250, n38251,
    n38252, n38254, n38255, n38256, n38257, n38258,
    n38259, n38260, n38261, n38262, n38263, n38264,
    n38265, n38266, n38267, n38269, n38270, n38271,
    n38272, n38273, n38274, n38275, n38276, n38277,
    n38278, n38279, n38280, n38281, n38282, n38283,
    n38284, n38285, n38286, n38287, n38288, n38289,
    n38290, n38291, n38292, n38293, n38294, n38295,
    n38296, n38297, n38298, n38299, n38300, n38301,
    n38302, n38303, n38304, n38305, n38306, n38307,
    n38308, n38309, n38310, n38311, n38312, n38313,
    n38314, n38315, n38316, n38317, n38318, n38319,
    n38320, n38321, n38322, n38323, n38324, n38325,
    n38326, n38327, n38328, n38329, n38330, n38331,
    n38332, n38333, n38334, n38335, n38336, n38337,
    n38338, n38339, n38340, n38341, n38342, n38343,
    n38344, n38345, n38346, n38347, n38348, n38349,
    n38350, n38351, n38352, n38353, n38354, n38355,
    n38356, n38357, n38358, n38359, n38360, n38361,
    n38362, n38363, n38364, n38365, n38366, n38367,
    n38368, n38369, n38370, n38371, n38372, n38373,
    n38374, n38375, n38376, n38377, n38378, n38379,
    n38380, n38381, n38382, n38383, n38384, n38385,
    n38386, n38387, n38388, n38389, n38390, n38391,
    n38392, n38393, n38394, n38395, n38396, n38397,
    n38398, n38399, n38400, n38401, n38402, n38403,
    n38404, n38405, n38406, n38407, n38408, n38409,
    n38410, n38411, n38412, n38413, n38414, n38415,
    n38416, n38417, n38418, n38419, n38420, n38421,
    n38422, n38423, n38424, n38425, n38426, n38427,
    n38428, n38429, n38430, n38431, n38432, n38433,
    n38434, n38435, n38436, n38437, n38438, n38439,
    n38440, n38441, n38442, n38443, n38444, n38445,
    n38446, n38447, n38448, n38449, n38450, n38451,
    n38452, n38453, n38454, n38455, n38456, n38457,
    n38458, n38459, n38460, n38461, n38462, n38463,
    n38464, n38465, n38466, n38467, n38468, n38469,
    n38470, n38471, n38472, n38473, n38474, n38475,
    n38476, n38477, n38478, n38479, n38480, n38481,
    n38482, n38483, n38484, n38485, n38486, n38487,
    n38488, n38489, n38490, n38491, n38492, n38493,
    n38494, n38495, n38496, n38497, n38498, n38499,
    n38500, n38501, n38502, n38503, n38504, n38505,
    n38506, n38507, n38508, n38509, n38510, n38511,
    n38512, n38513, n38514, n38515, n38516, n38517,
    n38518, n38519, n38520, n38521, n38522, n38523,
    n38524, n38525, n38526, n38527, n38528, n38529,
    n38530, n38531, n38532, n38533, n38534, n38535,
    n38536, n38537, n38538, n38539, n38540, n38541,
    n38542, n38543, n38544, n38545, n38546, n38547,
    n38548, n38549, n38550, n38551, n38552, n38553,
    n38554, n38555, n38556, n38557, n38558, n38559,
    n38560, n38561, n38562, n38563, n38564, n38565,
    n38566, n38567, n38568, n38569, n38570, n38571,
    n38572, n38573, n38574, n38575, n38576, n38577,
    n38578, n38580, n38581, n38582, n38583, n38584,
    n38585, n38586, n38587, n38588, n38589, n38590,
    n38591, n38592, n38593, n38594, n38595, n38596,
    n38597, n38598, n38599, n38600, n38601, n38602,
    n38603, n38604, n38605, n38606, n38607, n38608,
    n38609, n38610, n38611, n38612, n38613, n38614,
    n38615, n38616, n38617, n38618, n38619, n38620,
    n38621, n38622, n38623, n38624, n38625, n38626,
    n38627, n38628, n38629, n38630, n38631, n38632,
    n38633, n38634, n38635, n38636, n38637, n38638,
    n38639, n38640, n38641, n38642, n38643, n38644,
    n38645, n38646, n38647, n38648, n38649, n38650,
    n38651, n38652, n38653, n38654, n38655, n38656,
    n38657, n38658, n38659, n38660, n38661, n38662,
    n38663, n38664, n38665, n38666, n38667, n38668,
    n38669, n38670, n38671, n38672, n38673, n38674,
    n38675, n38676, n38677, n38678, n38679, n38680,
    n38681, n38682, n38683, n38684, n38685, n38686,
    n38687, n38688, n38689, n38690, n38691, n38692,
    n38693, n38694, n38695, n38696, n38697, n38698,
    n38699, n38700, n38701, n38702, n38703, n38704,
    n38705, n38706, n38707, n38708, n38709, n38710,
    n38711, n38712, n38713, n38714, n38715, n38716,
    n38717, n38718, n38719, n38720, n38721, n38722,
    n38723, n38724, n38725, n38727, n38728, n38729,
    n38730, n38731, n38732, n38733, n38734, n38735,
    n38736, n38737, n38738, n38739, n38740, n38741,
    n38742, n38743, n38744, n38745, n38746, n38747,
    n38748, n38749, n38750, n38751, n38752, n38753,
    n38754, n38755, n38756, n38757, n38758, n38759,
    n38760, n38761, n38762, n38763, n38764, n38765,
    n38766, n38767, n38768, n38769, n38770, n38771,
    n38772, n38773, n38774, n38775, n38776, n38777,
    n38778, n38779, n38780, n38781, n38782, n38783,
    n38784, n38785, n38786, n38787, n38788, n38789,
    n38790, n38791, n38792, n38793, n38794, n38795,
    n38796, n38797, n38798, n38799, n38800, n38801,
    n38802, n38803, n38804, n38805, n38806, n38807,
    n38808, n38809, n38810, n38811, n38812, n38813,
    n38814, n38815, n38816, n38817, n38818, n38819,
    n38820, n38821, n38822, n38823, n38824, n38825,
    n38826, n38827, n38828, n38829, n38830, n38831,
    n38832, n38833, n38834, n38835, n38836, n38837,
    n38838, n38839, n38840, n38841, n38842, n38843,
    n38844, n38845, n38846, n38848, n38849, n38850,
    n38851, n38852, n38853, n38854, n38855, n38856,
    n38857, n38858, n38859, n38860, n38861, n38862,
    n38863, n38864, n38865, n38866, n38867, n38868,
    n38869, n38870, n38871, n38872, n38873, n38874,
    n38875, n38876, n38877, n38878, n38879, n38880,
    n38881, n38882, n38883, n38884, n38885, n38886,
    n38887, n38888, n38889, n38890, n38891, n38892,
    n38893, n38894, n38895, n38896, n38897, n38898,
    n38899, n38900, n38901, n38902, n38903, n38904,
    n38905, n38906, n38907, n38908, n38909, n38910,
    n38911, n38912, n38913, n38914, n38915, n38916,
    n38917, n38918, n38919, n38920, n38921, n38922,
    n38923, n38924, n38925, n38926, n38928, n38929,
    n38930, n38931, n38932, n38933, n38934, n38935,
    n38936, n38937, n38938, n38939, n38940, n38941,
    n38942, n38943, n38944, n38945, n38946, n38947,
    n38948, n38949, n38950, n38951, n38952, n38953,
    n38954, n38955, n38956, n38958, n38959, n38960,
    n38961, n38962, n38963, n38964, n38965, n38966,
    n38967, n38968, n38969, n38971, n38972, n38973,
    n38974, n38975, n38976, n38977, n38978, n38979,
    n38980, n38981, n38982, n38983, n38984, n38985,
    n38986, n38987, n38988, n38989, n38990, n38991,
    n38992, n38993, n38994, n38995, n38996, n38997,
    n38998, n38999, n39000, n39001, n39002, n39003,
    n39004, n39005, n39006, n39007, n39008, n39009,
    n39010, n39011, n39012, n39013, n39014, n39015,
    n39016, n39017, n39018, n39019, n39020, n39021,
    n39022, n39023, n39024, n39025, n39026, n39027,
    n39028, n39029, n39030, n39031, n39032, n39033,
    n39034, n39035, n39036, n39037, n39038, n39039,
    n39040, n39041, n39042, n39043, n39044, n39045,
    n39046, n39047, n39048, n39049, n39050, n39051,
    n39052, n39053, n39054, n39055, n39056, n39057,
    n39058, n39059, n39060, n39061, n39062, n39063,
    n39064, n39065, n39066, n39067, n39068, n39069,
    n39070, n39071, n39072, n39073, n39074, n39075,
    n39076, n39077, n39078, n39079, n39080, n39081,
    n39082, n39083, n39084, n39085, n39086, n39087,
    n39088, n39089, n39090, n39091, n39092, n39093,
    n39094, n39095, n39096, n39097, n39098, n39099,
    n39100, n39101, n39102, n39103, n39104, n39105,
    n39106, n39107, n39108, n39109, n39110, n39111,
    n39112, n39113, n39114, n39115, n39116, n39117,
    n39118, n39119, n39120, n39121, n39122, n39123,
    n39124, n39125, n39126, n39127, n39128, n39129,
    n39130, n39131, n39132, n39133, n39134, n39135,
    n39136, n39137, n39138, n39139, n39140, n39141,
    n39142, n39143, n39144, n39145, n39146, n39147,
    n39148, n39149, n39150, n39151, n39152, n39153,
    n39154, n39155, n39156, n39157, n39158, n39159,
    n39160, n39161, n39162, n39163, n39164, n39165,
    n39166, n39167, n39168, n39169, n39170, n39171,
    n39172, n39173, n39174, n39175, n39176, n39177,
    n39178, n39179, n39180, n39181, n39182, n39183,
    n39184, n39185, n39186, n39187, n39188, n39189,
    n39190, n39191, n39192, n39193, n39194, n39195,
    n39196, n39197, n39198, n39199, n39200, n39201,
    n39202, n39203, n39204, n39205, n39206, n39207,
    n39208, n39209, n39210, n39211, n39212, n39213,
    n39214, n39215, n39216, n39217, n39218, n39219,
    n39220, n39221, n39222, n39223, n39224, n39225,
    n39226, n39227, n39228, n39229, n39230, n39231,
    n39232, n39233, n39234, n39235, n39236, n39237,
    n39238, n39239, n39240, n39241, n39242, n39243,
    n39244, n39245, n39246, n39247, n39248, n39249,
    n39250, n39251, n39252, n39253, n39254, n39255,
    n39256, n39257, n39258, n39259, n39260, n39261,
    n39262, n39263, n39264, n39265, n39266, n39267,
    n39268, n39269, n39270, n39271, n39272, n39273,
    n39274, n39275, n39276, n39277, n39278, n39279,
    n39280, n39281, n39282, n39283, n39284, n39285,
    n39286, n39287, n39288, n39289, n39290, n39291,
    n39292, n39293, n39294, n39295, n39296, n39297,
    n39298, n39299, n39300, n39301, n39302, n39303,
    n39304, n39305, n39306, n39307, n39308, n39309,
    n39310, n39311, n39312, n39313, n39314, n39315,
    n39316, n39317, n39318, n39319, n39320, n39321,
    n39322, n39323, n39324, n39325, n39326, n39327,
    n39328, n39329, n39330, n39331, n39332, n39333,
    n39334, n39335, n39336, n39337, n39338, n39339,
    n39340, n39341, n39342, n39343, n39344, n39345,
    n39346, n39347, n39348, n39349, n39350, n39351,
    n39352, n39353, n39354, n39355, n39356, n39357,
    n39358, n39359, n39360, n39361, n39362, n39363,
    n39364, n39365, n39366, n39367, n39368, n39369,
    n39370, n39371, n39372, n39373, n39374, n39375,
    n39376, n39377, n39378, n39379, n39380, n39381,
    n39382, n39383, n39384, n39385, n39386, n39387,
    n39388, n39389, n39390, n39391, n39392, n39393,
    n39394, n39395, n39396, n39397, n39398, n39399,
    n39400, n39401, n39402, n39403, n39404, n39405,
    n39406, n39407, n39408, n39409, n39410, n39411,
    n39412, n39413, n39414, n39415, n39416, n39417,
    n39418, n39419, n39420, n39421, n39422, n39423,
    n39424, n39425, n39426, n39427, n39428, n39429,
    n39430, n39431, n39432, n39433, n39434, n39435,
    n39436, n39437, n39438, n39439, n39440, n39441,
    n39442, n39443, n39444, n39445, n39446, n39447,
    n39448, n39449, n39450, n39451, n39452, n39453,
    n39454, n39455, n39456, n39457, n39458, n39459,
    n39460, n39461, n39462, n39463, n39464, n39465,
    n39466, n39467, n39468, n39469, n39470, n39471,
    n39472, n39473, n39474, n39475, n39476, n39477,
    n39478, n39479, n39480, n39481, n39482, n39483,
    n39484, n39485, n39486, n39487, n39488, n39489,
    n39490, n39491, n39492, n39493, n39494, n39495,
    n39496, n39497, n39498, n39499, n39500, n39501,
    n39502, n39503, n39504, n39505, n39506, n39507,
    n39508, n39509, n39510, n39511, n39512, n39513,
    n39514, n39515, n39516, n39517, n39518, n39519,
    n39520, n39521, n39522, n39523, n39524, n39525,
    n39526, n39527, n39528, n39529, n39530, n39531,
    n39532, n39533, n39534, n39535, n39536, n39537,
    n39538, n39539, n39540, n39541, n39542, n39543,
    n39544, n39545, n39546, n39547, n39548, n39549,
    n39550, n39551, n39552, n39553, n39554, n39555,
    n39556, n39557, n39558, n39559, n39560, n39561,
    n39562, n39563, n39564, n39565, n39566, n39567,
    n39568, n39569, n39570, n39571, n39572, n39573,
    n39574, n39575, n39576, n39577, n39578, n39579,
    n39580, n39581, n39582, n39583, n39584, n39585,
    n39586, n39587, n39588, n39589, n39590, n39591,
    n39592, n39593, n39594, n39595, n39596, n39597,
    n39598, n39599, n39600, n39601, n39602, n39603,
    n39604, n39605, n39606, n39607, n39608, n39609,
    n39610, n39611, n39612, n39613, n39614, n39615,
    n39616, n39617, n39618, n39619, n39620, n39621,
    n39622, n39623, n39624, n39625, n39626, n39627,
    n39628, n39629, n39630, n39631, n39632, n39633,
    n39634, n39635, n39636, n39637, n39638, n39639,
    n39640, n39641, n39642, n39643, n39644, n39645,
    n39646, n39647, n39648, n39649, n39650, n39651,
    n39652, n39653, n39654, n39655, n39656, n39657,
    n39658, n39659, n39660, n39661, n39662, n39663,
    n39664, n39665, n39666, n39667, n39668, n39669,
    n39670, n39671, n39672, n39673, n39674, n39675,
    n39676, n39677, n39678, n39679, n39680, n39681,
    n39682, n39683, n39684, n39685, n39686, n39687,
    n39688, n39689, n39690, n39691, n39692, n39693,
    n39694, n39695, n39696, n39697, n39698, n39699,
    n39700, n39701, n39702, n39703, n39704, n39705,
    n39706, n39707, n39708, n39709, n39710, n39711,
    n39712, n39713, n39714, n39715, n39716, n39717,
    n39718, n39719, n39720, n39721, n39722, n39723,
    n39724, n39725, n39726, n39727, n39728, n39729,
    n39730, n39731, n39732, n39733, n39734, n39735,
    n39736, n39737, n39738, n39739, n39740, n39741,
    n39742, n39743, n39744, n39745, n39746, n39747,
    n39748, n39749, n39750, n39751, n39752, n39753,
    n39754, n39755, n39756, n39757, n39758, n39759,
    n39760, n39761, n39762, n39763, n39764, n39765,
    n39766, n39767, n39768, n39769, n39770, n39771,
    n39772, n39773, n39774, n39775, n39776, n39777,
    n39778, n39779, n39780, n39781, n39782, n39783,
    n39784, n39785, n39786, n39787, n39788, n39789,
    n39790, n39791, n39792, n39793, n39794, n39795,
    n39796, n39797, n39798, n39799, n39800, n39801,
    n39802, n39803, n39804, n39805, n39806, n39807,
    n39808, n39809, n39810, n39811, n39812, n39813,
    n39814, n39815, n39816, n39817, n39818, n39819,
    n39820, n39821, n39822, n39823, n39824, n39825,
    n39826, n39827, n39828, n39829, n39830, n39831,
    n39832, n39833, n39834, n39835, n39836, n39838,
    n39839, n39840, n39841, n39842, n39843, n39844,
    n39846, n39847, n39848, n39849, n39850, n39851,
    n39852, n39853, n39854, n39855, n39856, n39857,
    n39858, n39859, n39860, n39861, n39862, n39864,
    n39865, n39866, n39867, n39868, n39869, n39870,
    n39871, n39872, n39873, n39874, n39875, n39876,
    n39877, n39878, n39879, n39880, n39881, n39882,
    n39883, n39884, n39885, n39886, n39887, n39888,
    n39889, n39890, n39891, n39892, n39893, n39894,
    n39895, n39896, n39897, n39898, n39899, n39900,
    n39901, n39902, n39903, n39904, n39905, n39906,
    n39907, n39908, n39909, n39910, n39911, n39912,
    n39913, n39914, n39915, n39916, n39917, n39918,
    n39919, n39920, n39921, n39922, n39923, n39924,
    n39925, n39926, n39927, n39928, n39929, n39930,
    n39931, n39932, n39933, n39934, n39935, n39936,
    n39937, n39938, n39939, n39940, n39941, n39942,
    n39943, n39944, n39945, n39946, n39947, n39948,
    n39949, n39950, n39951, n39952, n39953, n39954,
    n39955, n39956, n39957, n39958, n39959, n39960,
    n39961, n39962, n39963, n39964, n39965, n39966,
    n39967, n39968, n39969, n39970, n39971, n39972,
    n39973, n39974, n39975, n39976, n39977, n39978,
    n39979, n39980, n39981, n39982, n39983, n39984,
    n39985, n39986, n39987, n39988, n39989, n39990,
    n39991, n39992, n39993, n39994, n39995, n39996,
    n39997, n39998, n39999, n40000, n40001, n40002,
    n40003, n40004, n40005, n40006, n40007, n40008,
    n40009, n40010, n40011, n40012, n40013, n40014,
    n40015, n40016, n40017, n40018, n40019, n40020,
    n40021, n40022, n40023, n40024, n40025, n40026,
    n40027, n40028, n40029, n40030, n40031, n40032,
    n40033, n40034, n40035, n40036, n40037, n40038,
    n40039, n40040, n40041, n40042, n40043, n40044,
    n40045, n40046, n40047, n40048, n40050, n40051,
    n40052, n40054, n40055, n40056, n40057, n40058,
    n40059, n40060, n40061, n40062, n40063, n40064,
    n40065, n40066, n40067, n40068, n40069, n40070,
    n40071, n40072, n40073, n40074, n40075, n40076,
    n40077, n40078, n40079, n40080, n40081, n40082,
    n40083, n40084, n40085, n40086, n40087, n40088,
    n40089, n40090, n40091, n40092, n40093, n40094,
    n40095, n40096, n40097, n40098, n40099, n40100,
    n40101, n40103, n40104, n40105, n40106, n40107,
    n40108, n40109, n40110, n40111, n40112, n40113,
    n40114, n40115, n40116, n40117, n40118, n40119,
    n40120, n40121, n40122, n40123, n40124, n40125,
    n40126, n40127, n40128, n40129, n40130, n40131,
    n40132, n40133, n40134, n40135, n40136, n40137,
    n40138, n40139, n40140, n40141, n40142, n40143,
    n40144, n40145, n40146, n40147, n40148, n40149,
    n40150, n40151, n40152, n40153, n40154, n40155,
    n40156, n40157, n40158, n40159, n40160, n40161,
    n40162, n40163, n40164, n40165, n40166, n40168,
    n40169, n40170, n40171, n40172, n40173, n40174,
    n40175, n40176, n40177, n40178, n40179, n40180,
    n40181, n40182, n40183, n40184, n40185, n40186,
    n40187, n40188, n40189, n40190, n40191, n40192,
    n40193, n40194, n40195, n40196, n40197, n40198,
    n40199, n40200, n40201, n40202, n40203, n40204,
    n40205, n40206, n40207, n40208, n40209, n40210,
    n40211, n40212, n40213, n40214, n40215, n40216,
    n40217, n40218, n40219, n40220, n40221, n40222,
    n40223, n40224, n40225, n40226, n40227, n40228,
    n40229, n40230, n40231, n40232, n40233, n40234,
    n40235, n40236, n40237, n40238, n40239, n40240,
    n40241, n40242, n40244, n40245, n40246, n40247,
    n40248, n40249, n40250, n40251, n40252, n40253,
    n40254, n40255, n40256, n40257, n40258, n40259,
    n40260, n40261, n40262, n40263, n40264, n40265,
    n40266, n40267, n40268, n40269, n40270, n40271,
    n40272, n40273, n40274, n40275, n40276, n40277,
    n40278, n40279, n40280, n40281, n40282, n40283,
    n40284, n40285, n40286, n40287, n40288, n40289,
    n40290, n40291, n40292, n40293, n40294, n40295,
    n40296, n40297, n40298, n40299, n40300, n40301,
    n40302, n40303, n40304, n40305, n40306, n40307,
    n40308, n40309, n40310, n40311, n40312, n40313,
    n40314, n40315, n40316, n40317, n40318, n40319,
    n40320, n40321, n40322, n40323, n40324, n40325,
    n40326, n40327, n40328, n40329, n40330, n40331,
    n40332, n40333, n40334, n40335, n40336, n40337,
    n40338, n40339, n40341, n40342, n40343, n40344,
    n40345, n40346, n40347, n40348, n40349, n40350,
    n40351, n40352, n40353, n40354, n40355, n40356,
    n40357, n40358, n40359, n40360, n40361, n40362,
    n40363, n40364, n40365, n40366, n40367, n40368,
    n40369, n40370, n40371, n40372, n40373, n40374,
    n40375, n40376, n40377, n40378, n40379, n40380,
    n40381, n40382, n40383, n40384, n40385, n40386,
    n40387, n40388, n40389, n40390, n40391, n40392,
    n40393, n40394, n40395, n40396, n40397, n40398,
    n40399, n40400, n40401, n40402, n40403, n40404,
    n40405, n40406, n40407, n40408, n40409, n40410,
    n40411, n40412, n40413, n40414, n40415, n40416,
    n40417, n40418, n40419, n40420, n40421, n40422,
    n40423, n40424, n40425, n40426, n40427, n40428,
    n40429, n40430, n40431, n40432, n40433, n40434,
    n40435, n40436, n40437, n40438, n40439, n40440,
    n40441, n40442, n40443, n40444, n40445, n40446,
    n40447, n40448, n40449, n40450, n40451, n40452,
    n40453, n40454, n40455, n40456, n40457, n40458,
    n40459, n40460, n40461, n40462, n40463, n40464,
    n40465, n40466, n40467, n40468, n40469, n40470,
    n40471, n40472, n40473, n40474, n40475, n40476,
    n40477, n40478, n40479, n40480, n40481, n40482,
    n40483, n40484, n40485, n40486, n40487, n40488,
    n40489, n40490, n40491, n40492, n40493, n40494,
    n40495, n40496, n40497, n40498, n40499, n40500,
    n40501, n40502, n40503, n40504, n40505, n40506,
    n40507, n40508, n40509, n40510, n40511, n40512,
    n40513, n40514, n40515, n40516, n40517, n40518,
    n40519, n40520, n40521, n40522, n40523, n40524,
    n40525, n40526, n40527, n40528, n40529, n40530,
    n40531, n40532, n40533, n40534, n40535, n40536,
    n40537, n40538, n40539, n40540, n40541, n40542,
    n40543, n40544, n40545, n40546, n40547, n40548,
    n40549, n40550, n40551, n40552, n40553, n40554,
    n40555, n40556, n40557, n40558, n40559, n40560,
    n40561, n40562, n40563, n40564, n40565, n40566,
    n40567, n40568, n40569, n40570, n40571, n40572,
    n40573, n40574, n40575, n40576, n40577, n40578,
    n40579, n40580, n40581, n40582, n40583, n40584,
    n40585, n40586, n40587, n40588, n40589, n40590,
    n40591, n40592, n40593, n40594, n40595, n40596,
    n40597, n40598, n40599, n40600, n40601, n40602,
    n40603, n40604, n40605, n40606, n40607, n40608,
    n40609, n40610, n40611, n40612, n40613, n40614,
    n40615, n40616, n40617, n40618, n40619, n40620,
    n40621, n40622, n40623, n40624, n40625, n40626,
    n40627, n40628, n40629, n40630, n40631, n40632,
    n40633, n40634, n40635, n40636, n40637, n40638,
    n40639, n40640, n40641, n40642, n40643, n40644,
    n40645, n40646, n40647, n40648, n40649, n40650,
    n40651, n40652, n40653, n40654, n40655, n40656,
    n40657, n40658, n40659, n40660, n40661, n40662,
    n40663, n40664, n40665, n40666, n40667, n40668,
    n40669, n40670, n40671, n40672, n40673, n40674,
    n40675, n40676, n40677, n40678, n40679, n40680,
    n40681, n40682, n40683, n40684, n40685, n40686,
    n40687, n40688, n40689, n40690, n40691, n40692,
    n40693, n40694, n40695, n40696, n40697, n40698,
    n40699, n40700, n40701, n40702, n40703, n40704,
    n40705, n40706, n40707, n40708, n40709, n40710,
    n40711, n40712, n40713, n40714, n40715, n40716,
    n40717, n40718, n40719, n40720, n40721, n40722,
    n40723, n40724, n40725, n40726, n40727, n40728,
    n40729, n40730, n40731, n40732, n40733, n40734,
    n40735, n40736, n40737, n40738, n40739, n40740,
    n40741, n40742, n40743, n40744, n40745, n40746,
    n40747, n40748, n40749, n40750, n40751, n40752,
    n40753, n40754, n40755, n40756, n40757, n40758,
    n40759, n40760, n40761, n40762, n40763, n40764,
    n40765, n40766, n40767, n40768, n40769, n40770,
    n40771, n40772, n40773, n40774, n40775, n40776,
    n40777, n40778, n40779, n40780, n40781, n40782,
    n40783, n40784, n40785, n40786, n40787, n40788,
    n40789, n40790, n40791, n40792, n40793, n40794,
    n40795, n40796, n40797, n40798, n40799, n40800,
    n40801, n40802, n40803, n40804, n40805, n40806,
    n40807, n40808, n40809, n40810, n40811, n40812,
    n40813, n40814, n40815, n40816, n40817, n40818,
    n40819, n40820, n40821, n40822, n40823, n40824,
    n40825, n40826, n40827, n40828, n40829, n40830,
    n40831, n40832, n40833, n40834, n40835, n40836,
    n40838, n40839, n40840, n40841, n40842, n40843,
    n40844, n40845, n40846, n40847, n40848, n40849,
    n40850, n40851, n40852, n40853, n40854, n40855,
    n40856, n40857, n40858, n40859, n40860, n40861,
    n40862, n40863, n40864, n40865, n40866, n40867,
    n40868, n40869, n40870, n40871, n40872, n40873,
    n40874, n40875, n40876, n40877, n40878, n40879,
    n40880, n40881, n40882, n40883, n40884, n40885,
    n40886, n40887, n40888, n40889, n40890, n40891,
    n40892, n40893, n40894, n40895, n40897, n40898,
    n40899, n40900, n40901, n40902, n40903, n40904,
    n40905, n40906, n40907, n40908, n40909, n40910,
    n40911, n40912, n40913, n40914, n40915, n40916,
    n40917, n40918, n40919, n40920, n40921, n40922,
    n40923, n40924, n40925, n40926, n40927, n40928,
    n40929, n40930, n40931, n40932, n40933, n40934,
    n40935, n40936, n40937, n40938, n40939, n40940,
    n40941, n40942, n40943, n40944, n40945, n40947,
    n40948, n40949, n40950, n40951, n40952, n40953,
    n40954, n40955, n40956, n40957, n40958, n40959,
    n40960, n40961, n40962, n40963, n40964, n40965,
    n40966, n40967, n40968, n40969, n40970, n40971,
    n40972, n40973, n40974, n40975, n40976, n40977,
    n40978, n40979, n40980, n40981, n40982, n40983,
    n40984, n40985, n40986, n40987, n40988, n40989,
    n40990, n40991, n40992, n40993, n40994, n40995,
    n40996, n40997, n40998, n40999, n41000, n41001,
    n41002, n41003, n41004, n41006, n41007, n41008,
    n41009, n41010, n41011, n41012, n41013, n41014,
    n41015, n41016, n41017, n41018, n41019, n41020,
    n41021, n41022, n41023, n41024, n41025, n41026,
    n41027, n41028, n41029, n41030, n41031, n41032,
    n41033, n41034, n41035, n41036, n41037, n41038,
    n41039, n41040, n41041, n41042, n41043, n41044,
    n41045, n41046, n41047, n41048, n41049, n41050,
    n41051, n41052, n41053, n41054, n41055, n41056,
    n41057, n41058, n41059, n41060, n41061, n41062,
    n41063, n41064, n41065, n41066, n41067, n41068,
    n41069, n41070, n41071, n41072, n41073, n41074,
    n41075, n41076, n41077, n41078, n41079, n41080,
    n41081, n41082, n41083, n41084, n41085, n41086,
    n41087, n41088, n41089, n41090, n41091, n41092,
    n41093, n41094, n41095, n41096, n41097, n41098,
    n41099, n41100, n41101, n41102, n41103, n41104,
    n41105, n41106, n41107, n41108, n41109, n41110,
    n41111, n41112, n41113, n41114, n41115, n41116,
    n41117, n41118, n41119, n41120, n41121, n41122,
    n41123, n41124, n41125, n41126, n41127, n41128,
    n41129, n41130, n41131, n41132, n41133, n41134,
    n41135, n41136, n41137, n41138, n41139, n41140,
    n41141, n41142, n41143, n41144, n41145, n41146,
    n41147, n41148, n41149, n41150, n41151, n41152,
    n41153, n41154, n41155, n41156, n41157, n41158,
    n41159, n41160, n41161, n41162, n41163, n41164,
    n41165, n41166, n41167, n41168, n41169, n41170,
    n41171, n41172, n41173, n41174, n41175, n41176,
    n41177, n41178, n41179, n41180, n41181, n41182,
    n41183, n41184, n41185, n41186, n41187, n41188,
    n41189, n41190, n41191, n41192, n41193, n41194,
    n41195, n41196, n41197, n41198, n41199, n41200,
    n41201, n41202, n41203, n41204, n41205, n41206,
    n41207, n41208, n41209, n41210, n41211, n41212,
    n41213, n41214, n41215, n41216, n41217, n41218,
    n41219, n41220, n41221, n41222, n41223, n41224,
    n41225, n41226, n41227, n41228, n41229, n41230,
    n41231, n41232, n41233, n41234, n41235, n41236,
    n41237, n41238, n41239, n41240, n41241, n41242,
    n41243, n41244, n41245, n41246, n41247, n41248,
    n41249, n41250, n41251, n41252, n41253, n41254,
    n41255, n41256, n41257, n41258, n41259, n41260,
    n41261, n41262, n41263, n41264, n41265, n41266,
    n41267, n41268, n41269, n41270, n41271, n41272,
    n41273, n41274, n41275, n41276, n41277, n41278,
    n41279, n41280, n41281, n41282, n41283, n41284,
    n41285, n41286, n41287, n41288, n41289, n41290,
    n41291, n41292, n41293, n41294, n41295, n41296,
    n41297, n41298, n41299, n41300, n41301, n41302,
    n41303, n41304, n41305, n41306, n41307, n41308,
    n41309, n41310, n41311, n41312, n41313, n41314,
    n41315, n41316, n41317, n41318, n41319, n41320,
    n41321, n41322, n41323, n41324, n41325, n41326,
    n41327, n41328, n41329, n41330, n41331, n41332,
    n41333, n41334, n41335, n41336, n41337, n41338,
    n41339, n41340, n41341, n41342, n41343, n41344,
    n41345, n41346, n41347, n41348, n41349, n41350,
    n41351, n41352, n41353, n41354, n41355, n41356,
    n41357, n41358, n41359, n41360, n41361, n41362,
    n41363, n41364, n41365, n41366, n41367, n41368,
    n41369, n41370, n41371, n41372, n41373, n41374,
    n41375, n41376, n41377, n41378, n41379, n41380,
    n41381, n41382, n41383, n41384, n41385, n41386,
    n41387, n41388, n41389, n41390, n41391, n41392,
    n41393, n41394, n41395, n41396, n41397, n41398,
    n41399, n41400, n41401, n41402, n41403, n41404,
    n41405, n41406, n41407, n41408, n41409, n41410,
    n41411, n41412, n41413, n41414, n41415, n41416,
    n41417, n41418, n41419, n41420, n41421, n41422,
    n41423, n41424, n41425, n41426, n41427, n41428,
    n41429, n41430, n41431, n41432, n41433, n41434,
    n41435, n41436, n41437, n41438, n41439, n41440,
    n41441, n41442, n41443, n41444, n41445, n41446,
    n41447, n41448, n41449, n41450, n41451, n41452,
    n41453, n41454, n41455, n41456, n41457, n41458,
    n41459, n41460, n41461, n41462, n41463, n41464,
    n41465, n41466, n41467, n41468, n41469, n41470,
    n41471, n41472, n41473, n41474, n41475, n41476,
    n41477, n41478, n41479, n41480, n41481, n41482,
    n41483, n41484, n41485, n41486, n41487, n41488,
    n41489, n41490, n41491, n41492, n41493, n41494,
    n41495, n41496, n41497, n41498, n41499, n41500,
    n41501, n41502, n41503, n41504, n41505, n41506,
    n41507, n41508, n41509, n41510, n41511, n41512,
    n41513, n41514, n41515, n41516, n41517, n41518,
    n41519, n41520, n41521, n41522, n41523, n41524,
    n41525, n41526, n41527, n41528, n41529, n41530,
    n41531, n41532, n41533, n41534, n41535, n41536,
    n41537, n41538, n41539, n41540, n41541, n41542,
    n41543, n41544, n41545, n41546, n41547, n41548,
    n41549, n41550, n41551, n41552, n41553, n41554,
    n41555, n41556, n41557, n41558, n41559, n41560,
    n41561, n41562, n41563, n41564, n41565, n41566,
    n41567, n41568, n41569, n41570, n41571, n41572,
    n41573, n41574, n41575, n41576, n41577, n41578,
    n41579, n41580, n41581, n41582, n41583, n41584,
    n41585, n41586, n41587, n41588, n41589, n41590,
    n41591, n41592, n41593, n41594, n41595, n41596,
    n41597, n41598, n41599, n41600, n41601, n41602,
    n41603, n41604, n41605, n41606, n41607, n41608,
    n41609, n41610, n41611, n41612, n41613, n41614,
    n41615, n41616, n41617, n41618, n41619, n41620,
    n41621, n41622, n41623, n41624, n41625, n41626,
    n41627, n41628, n41629, n41630, n41631, n41632,
    n41633, n41634, n41635, n41636, n41637, n41638,
    n41639, n41640, n41641, n41642, n41643, n41644,
    n41645, n41646, n41647, n41648, n41649, n41650,
    n41651, n41652, n41653, n41654, n41655, n41656,
    n41657, n41658, n41659, n41660, n41661, n41662,
    n41663, n41664, n41665, n41666, n41667, n41668,
    n41669, n41670, n41671, n41672, n41673, n41674,
    n41675, n41676, n41677, n41678, n41679, n41680,
    n41681, n41682, n41683, n41684, n41685, n41686,
    n41687, n41688, n41689, n41690, n41691, n41692,
    n41693, n41694, n41695, n41696, n41697, n41698,
    n41699, n41700, n41701, n41702, n41703, n41704,
    n41705, n41706, n41707, n41708, n41709, n41710,
    n41711, n41712, n41713, n41714, n41715, n41716,
    n41717, n41718, n41719, n41720, n41721, n41722,
    n41723, n41724, n41725, n41726, n41727, n41728,
    n41729, n41730, n41731, n41732, n41733, n41734,
    n41735, n41736, n41737, n41738, n41739, n41740,
    n41742, n41743, n41744, n41745, n41746, n41747,
    n41748, n41749, n41750, n41751, n41752, n41753,
    n41754, n41755, n41756, n41757, n41758, n41759,
    n41760, n41762, n41763, n41764, n41765, n41766,
    n41767, n41768, n41769, n41770, n41771, n41772,
    n41773, n41774, n41775, n41776, n41777, n41778,
    n41779, n41780, n41781, n41782, n41783, n41784,
    n41785, n41786, n41787, n41788, n41789, n41790,
    n41791, n41792, n41793, n41794, n41795, n41796,
    n41797, n41798, n41799, n41800, n41801, n41802,
    n41803, n41804, n41805, n41806, n41807, n41808,
    n41809, n41810, n41811, n41812, n41813, n41814,
    n41815, n41816, n41817, n41818, n41819, n41820,
    n41821, n41822, n41823, n41824, n41825, n41826,
    n41827, n41828, n41829, n41830, n41831, n41832,
    n41833, n41834, n41835, n41836, n41837, n41838,
    n41839, n41840, n41841, n41842, n41843, n41844,
    n41845, n41846, n41847, n41848, n41849, n41850,
    n41851, n41852, n41853, n41854, n41855, n41856,
    n41857, n41858, n41859, n41860, n41861, n41862,
    n41863, n41864, n41865, n41866, n41867, n41868,
    n41869, n41870, n41871, n41872, n41873, n41874,
    n41875, n41876, n41877, n41878, n41879, n41880,
    n41881, n41882, n41883, n41884, n41885, n41886,
    n41887, n41888, n41889, n41890, n41891, n41892,
    n41893, n41894, n41895, n41896, n41897, n41898,
    n41899, n41900, n41901, n41902, n41903, n41904,
    n41905, n41906, n41907, n41908, n41909, n41910,
    n41911, n41912, n41913, n41914, n41915, n41916,
    n41917, n41918, n41919, n41920, n41921, n41922,
    n41923, n41924, n41925, n41926, n41927, n41928,
    n41929, n41930, n41931, n41932, n41933, n41934,
    n41935, n41936, n41937, n41938, n41939, n41940,
    n41941, n41942, n41943, n41944, n41945, n41946,
    n41947, n41948, n41949, n41950, n41951, n41952,
    n41953, n41954, n41955, n41956, n41957, n41958,
    n41959, n41960, n41961, n41962, n41963, n41964,
    n41965, n41966, n41967, n41968, n41969, n41970,
    n41971, n41972, n41973, n41974, n41975, n41976,
    n41977, n41978, n41979, n41980, n41981, n41982,
    n41983, n41984, n41985, n41986, n41987, n41988,
    n41989, n41990, n41991, n41992, n41993, n41994,
    n41995, n41996, n41997, n41998, n41999, n42000,
    n42001, n42002, n42003, n42004, n42005, n42006,
    n42007, n42008, n42009, n42010, n42011, n42012,
    n42013, n42014, n42015, n42016, n42017, n42018,
    n42019, n42020, n42021, n42022, n42023, n42024,
    n42025, n42026, n42027, n42028, n42029, n42030,
    n42031, n42032, n42033, n42034, n42035, n42036,
    n42037, n42038, n42039, n42040, n42041, n42042,
    n42043, n42044, n42045, n42046, n42047, n42048,
    n42049, n42050, n42051, n42052, n42053, n42054,
    n42055, n42056, n42057, n42058, n42059, n42060,
    n42061, n42062, n42063, n42064, n42065, n42066,
    n42067, n42068, n42069, n42070, n42071, n42072,
    n42073, n42074, n42075, n42076, n42077, n42078,
    n42079, n42080, n42081, n42082, n42083, n42084,
    n42085, n42086, n42087, n42088, n42089, n42090,
    n42091, n42092, n42093, n42094, n42095, n42096,
    n42097, n42098, n42099, n42100, n42101, n42102,
    n42103, n42104, n42105, n42106, n42107, n42108,
    n42109, n42110, n42111, n42112, n42113, n42114,
    n42115, n42116, n42117, n42118, n42119, n42120,
    n42121, n42122, n42123, n42124, n42125, n42126,
    n42127, n42128, n42129, n42130, n42131, n42132,
    n42133, n42134, n42135, n42136, n42137, n42138,
    n42139, n42140, n42141, n42142, n42143, n42144,
    n42145, n42146, n42147, n42148, n42149, n42150,
    n42151, n42152, n42153, n42154, n42155, n42156,
    n42157, n42158, n42159, n42160, n42161, n42162,
    n42163, n42164, n42165, n42166, n42167, n42168,
    n42169, n42170, n42171, n42172, n42173, n42174,
    n42175, n42176, n42177, n42178, n42179, n42180,
    n42181, n42182, n42183, n42184, n42185, n42186,
    n42187, n42188, n42189, n42190, n42191, n42192,
    n42193, n42194, n42195, n42196, n42197, n42198,
    n42199, n42200, n42201, n42202, n42203, n42204,
    n42205, n42206, n42207, n42208, n42209, n42210,
    n42211, n42212, n42213, n42214, n42215, n42216,
    n42217, n42218, n42219, n42220, n42221, n42222,
    n42223, n42224, n42225, n42226, n42227, n42228,
    n42229, n42230, n42231, n42232, n42233, n42234,
    n42235, n42236, n42237, n42238, n42239, n42240,
    n42241, n42242, n42243, n42244, n42245, n42246,
    n42247, n42248, n42249, n42250, n42251, n42252,
    n42253, n42254, n42255, n42256, n42257, n42258,
    n42259, n42260, n42261, n42262, n42263, n42264,
    n42265, n42266, n42267, n42268, n42269, n42270,
    n42271, n42272, n42273, n42274, n42275, n42276,
    n42277, n42278, n42279, n42280, n42281, n42282,
    n42283, n42284, n42285, n42286, n42287, n42288,
    n42289, n42290, n42291, n42292, n42293, n42294,
    n42295, n42296, n42297, n42298, n42299, n42300,
    n42301, n42302, n42303, n42304, n42305, n42306,
    n42307, n42308, n42309, n42310, n42311, n42312,
    n42313, n42314, n42315, n42316, n42317, n42318,
    n42319, n42320, n42321, n42322, n42323, n42324,
    n42325, n42326, n42327, n42328, n42329, n42330,
    n42331, n42332, n42333, n42334, n42335, n42336,
    n42337, n42338, n42339, n42340, n42341, n42342,
    n42343, n42344, n42345, n42346, n42347, n42348,
    n42349, n42350, n42351, n42352, n42353, n42354,
    n42355, n42356, n42357, n42358, n42359, n42360,
    n42361, n42362, n42363, n42364, n42365, n42366,
    n42367, n42368, n42369, n42370, n42371, n42372,
    n42373, n42374, n42375, n42376, n42377, n42378,
    n42379, n42380, n42381, n42382, n42383, n42384,
    n42385, n42386, n42387, n42388, n42389, n42390,
    n42391, n42392, n42393, n42394, n42395, n42396,
    n42397, n42398, n42399, n42400, n42401, n42402,
    n42403, n42404, n42405, n42406, n42407, n42408,
    n42409, n42410, n42411, n42412, n42413, n42414,
    n42415, n42416, n42417, n42418, n42419, n42420,
    n42421, n42422, n42423, n42424, n42425, n42426,
    n42427, n42428, n42429, n42430, n42431, n42432,
    n42433, n42434, n42435, n42436, n42437, n42438,
    n42439, n42440, n42441, n42442, n42443, n42444,
    n42445, n42446, n42447, n42448, n42449, n42450,
    n42451, n42452, n42453, n42454, n42455, n42456,
    n42457, n42458, n42459, n42460, n42461, n42462,
    n42463, n42464, n42465, n42466, n42467, n42468,
    n42469, n42470, n42471, n42472, n42473, n42474,
    n42475, n42476, n42477, n42478, n42479, n42480,
    n42481, n42482, n42483, n42484, n42485, n42486,
    n42487, n42488, n42489, n42490, n42491, n42492,
    n42493, n42494, n42495, n42496, n42497, n42498,
    n42499, n42500, n42501, n42502, n42503, n42504,
    n42505, n42506, n42507, n42508, n42509, n42510,
    n42511, n42512, n42513, n42514, n42515, n42516,
    n42517, n42518, n42519, n42520, n42521, n42522,
    n42523, n42524, n42525, n42526, n42527, n42528,
    n42529, n42530, n42531, n42532, n42533, n42534,
    n42535, n42536, n42537, n42538, n42539, n42540,
    n42541, n42542, n42543, n42544, n42545, n42546,
    n42547, n42548, n42549, n42550, n42551, n42552,
    n42553, n42554, n42555, n42556, n42557, n42558,
    n42559, n42560, n42561, n42562, n42563, n42564,
    n42565, n42566, n42567, n42568, n42569, n42570,
    n42571, n42572, n42573, n42574, n42575, n42576,
    n42577, n42578, n42579, n42580, n42581, n42582,
    n42583, n42584, n42585, n42586, n42587, n42588,
    n42589, n42590, n42591, n42592, n42593, n42594,
    n42595, n42596, n42597, n42598, n42599, n42600,
    n42601, n42602, n42603, n42604, n42605, n42606,
    n42607, n42608, n42609, n42610, n42611, n42612,
    n42613, n42614, n42615, n42616, n42617, n42618,
    n42619, n42620, n42621, n42622, n42623, n42624,
    n42625, n42626, n42627, n42628, n42629, n42630,
    n42631, n42632, n42633, n42634, n42635, n42636,
    n42637, n42638, n42639, n42640, n42641, n42642,
    n42643, n42644, n42645, n42646, n42647, n42648,
    n42649, n42650, n42651, n42652, n42653, n42654,
    n42655, n42656, n42657, n42658, n42659, n42660,
    n42661, n42662, n42663, n42664, n42665, n42666,
    n42667, n42668, n42669, n42670, n42671, n42672,
    n42673, n42674, n42675, n42676, n42677, n42678,
    n42679, n42680, n42681, n42682, n42683, n42684,
    n42685, n42686, n42687, n42688, n42689, n42690,
    n42691, n42692, n42693, n42694, n42695, n42696,
    n42697, n42698, n42699, n42700, n42701, n42702,
    n42703, n42704, n42705, n42706, n42707, n42708,
    n42709, n42710, n42711, n42712, n42713, n42714,
    n42715, n42716, n42717, n42718, n42719, n42720,
    n42721, n42722, n42723, n42724, n42725, n42726,
    n42727, n42728, n42729, n42730, n42731, n42732,
    n42733, n42734, n42735, n42736, n42737, n42738,
    n42739, n42740, n42741, n42742, n42743, n42744,
    n42745, n42746, n42747, n42748, n42749, n42750,
    n42751, n42752, n42753, n42754, n42755, n42756,
    n42757, n42758, n42759, n42760, n42761, n42762,
    n42763, n42764, n42765, n42766, n42767, n42768,
    n42769, n42770, n42771, n42772, n42773, n42774,
    n42775, n42776, n42777, n42778, n42779, n42780,
    n42781, n42782, n42783, n42784, n42785, n42786,
    n42787, n42788, n42789, n42790, n42791, n42792,
    n42793, n42794, n42795, n42796, n42797, n42798,
    n42799, n42800, n42801, n42802, n42803, n42804,
    n42805, n42806, n42807, n42808, n42809, n42810,
    n42811, n42812, n42813, n42814, n42815, n42816,
    n42817, n42818, n42819, n42820, n42821, n42822,
    n42823, n42824, n42825, n42826, n42827, n42828,
    n42829, n42830, n42831, n42832, n42833, n42834,
    n42835, n42836, n42837, n42838, n42839, n42840,
    n42841, n42842, n42843, n42844, n42845, n42846,
    n42847, n42848, n42849, n42850, n42851, n42852,
    n42853, n42854, n42855, n42856, n42857, n42858,
    n42859, n42860, n42861, n42862, n42863, n42864,
    n42865, n42866, n42867, n42868, n42869, n42870,
    n42871, n42872, n42873, n42874, n42875, n42876,
    n42877, n42878, n42879, n42880, n42881, n42882,
    n42883, n42884, n42885, n42886, n42887, n42888,
    n42889, n42890, n42891, n42892, n42893, n42894,
    n42895, n42896, n42897, n42898, n42899, n42900,
    n42901, n42902, n42903, n42904, n42905, n42906,
    n42907, n42908, n42909, n42910, n42911, n42912,
    n42913, n42914, n42915, n42916, n42917, n42918,
    n42919, n42920, n42921, n42922, n42923, n42924,
    n42925, n42926, n42927, n42928, n42929, n42930,
    n42931, n42932, n42933, n42934, n42935, n42936,
    n42937, n42938, n42939, n42940, n42941, n42942,
    n42943, n42944, n42945, n42946, n42947, n42948,
    n42949, n42950, n42951, n42952, n42953, n42954,
    n42955, n42956, n42957, n42958, n42959, n42960,
    n42961, n42962, n42963, n42964, n42965, n42966,
    n42967, n42968, n42969, n42970, n42971, n42972,
    n42973, n42974, n42975, n42976, n42977, n42978,
    n42979, n42980, n42981, n42982, n42983, n42984,
    n42985, n42986, n42987, n42988, n42989, n42990,
    n42991, n42992, n42993, n42994, n42995, n42996,
    n42997, n42998, n42999, n43000, n43001, n43002,
    n43003, n43004, n43005, n43006, n43007, n43008,
    n43009, n43010, n43011, n43012, n43013, n43014,
    n43015, n43016, n43017, n43018, n43019, n43020,
    n43021, n43022, n43023, n43024, n43025, n43026,
    n43027, n43028, n43029, n43030, n43031, n43032,
    n43033, n43034, n43035, n43036, n43037, n43038,
    n43039, n43040, n43041, n43042, n43043, n43044,
    n43045, n43046, n43047, n43048, n43049, n43050,
    n43051, n43052, n43053, n43054, n43055, n43056,
    n43057, n43058, n43059, n43060, n43061, n43062,
    n43063, n43064, n43065, n43066, n43067, n43068,
    n43069, n43070, n43071, n43072, n43073, n43074,
    n43075, n43076, n43077, n43078, n43079, n43080,
    n43081, n43082, n43083, n43084, n43085, n43086,
    n43087, n43088, n43089, n43090, n43091, n43092,
    n43093, n43094, n43095, n43096, n43097, n43098,
    n43099, n43100, n43101, n43102, n43103, n43104,
    n43105, n43106, n43107, n43108, n43109, n43110,
    n43111, n43112, n43113, n43114, n43115, n43116,
    n43117, n43118, n43119, n43120, n43121, n43122,
    n43123, n43124, n43125, n43126, n43127, n43128,
    n43129, n43130, n43131, n43132, n43133, n43134,
    n43135, n43136, n43137, n43138, n43139, n43140,
    n43141, n43142, n43143, n43144, n43145, n43146,
    n43147, n43148, n43149, n43150, n43151, n43152,
    n43153, n43154, n43155, n43156, n43157, n43158,
    n43159, n43160, n43161, n43162, n43163, n43164,
    n43165, n43166, n43167, n43168, n43169, n43170,
    n43171, n43172, n43173, n43174, n43175, n43176,
    n43177, n43178, n43179, n43180, n43181, n43182,
    n43183, n43184, n43185, n43186, n43187, n43188,
    n43189, n43190, n43191, n43192, n43193, n43194,
    n43195, n43196, n43197, n43198, n43199, n43200,
    n43201, n43202, n43203, n43204, n43205, n43206,
    n43207, n43208, n43209, n43210, n43211, n43212,
    n43213, n43214, n43215, n43216, n43217, n43218,
    n43219, n43220, n43221, n43222, n43223, n43224,
    n43225, n43226, n43227, n43228, n43229, n43230,
    n43231, n43233, n43234, n43235, n43236, n43237,
    n43238, n43239, n43240, n43241, n43242, n43243,
    n43244, n43245, n43246, n43247, n43248, n43249,
    n43250, n43251, n43252, n43253, n43254, n43255,
    n43256, n43257, n43258, n43259, n43260, n43261,
    n43262, n43263, n43264, n43265, n43266, n43267,
    n43268, n43269, n43270, n43271, n43272, n43273,
    n43274, n43275, n43276, n43277, n43278, n43279,
    n43280, n43281, n43282, n43283, n43284, n43285,
    n43286, n43287, n43288, n43289, n43290, n43291,
    n43292, n43293, n43294, n43295, n43296, n43297,
    n43298, n43299, n43300, n43301, n43302, n43303,
    n43304, n43305, n43306, n43307, n43308, n43309,
    n43310, n43311, n43312, n43313, n43314, n43315,
    n43316, n43317, n43318, n43319, n43320, n43321,
    n43322, n43323, n43324, n43325, n43326, n43327,
    n43328, n43329, n43330, n43331, n43332, n43333,
    n43334, n43335, n43336, n43337, n43338, n43339,
    n43340, n43341, n43342, n43343, n43344, n43345,
    n43346, n43347, n43348, n43349, n43350, n43351,
    n43352, n43353, n43354, n43355, n43356, n43357,
    n43358, n43359, n43360, n43361, n43362, n43363,
    n43364, n43365, n43366, n43367, n43368, n43369,
    n43370, n43371, n43372, n43373, n43374, n43375,
    n43376, n43377, n43378, n43379, n43380, n43381,
    n43382, n43383, n43384, n43385, n43386, n43387,
    n43388, n43389, n43390, n43391, n43392, n43393,
    n43394, n43395, n43396, n43397, n43398, n43399,
    n43400, n43401, n43402, n43403, n43404, n43405,
    n43406, n43407, n43408, n43409, n43410, n43411,
    n43412, n43413, n43414, n43415, n43416, n43417,
    n43418, n43419, n43420, n43421, n43422, n43423,
    n43424, n43425, n43426, n43427, n43428, n43429,
    n43430, n43431, n43432, n43433, n43434, n43435,
    n43436, n43437, n43438, n43439, n43440, n43441,
    n43442, n43443, n43444, n43445, n43446, n43447,
    n43448, n43449, n43450, n43451, n43452, n43453,
    n43454, n43455, n43456, n43457, n43458, n43459,
    n43460, n43461, n43462, n43463, n43464, n43465,
    n43466, n43467, n43468, n43469, n43470, n43471,
    n43472, n43473, n43474, n43475, n43476, n43477,
    n43478, n43479, n43480, n43481, n43482, n43483,
    n43484, n43485, n43486, n43487, n43488, n43489,
    n43490, n43491, n43492, n43493, n43494, n43495,
    n43496, n43497, n43498, n43499, n43500, n43501,
    n43502, n43503, n43504, n43505, n43506, n43507,
    n43508, n43509, n43510, n43511, n43512, n43513,
    n43514, n43515, n43516, n43517, n43518, n43519,
    n43520, n43521, n43522, n43523, n43524, n43525,
    n43526, n43527, n43528, n43529, n43530, n43531,
    n43532, n43533, n43534, n43535, n43536, n43537,
    n43538, n43539, n43540, n43541, n43542, n43543,
    n43544, n43545, n43546, n43547, n43548, n43549,
    n43550, n43551, n43552, n43553, n43554, n43555,
    n43556, n43557, n43558, n43559, n43560, n43561,
    n43562, n43563, n43564, n43565, n43566, n43567,
    n43568, n43569, n43570, n43571, n43572, n43573,
    n43574, n43575, n43576, n43577, n43578, n43579,
    n43580, n43581, n43582, n43583, n43584, n43585,
    n43586, n43587, n43588, n43589, n43590, n43591,
    n43592, n43593, n43594, n43595, n43596, n43597,
    n43598, n43599, n43600, n43601, n43602, n43603,
    n43604, n43605, n43606, n43607, n43608, n43609,
    n43610, n43611, n43612, n43613, n43614, n43615,
    n43616, n43617, n43618, n43619, n43620, n43621,
    n43622, n43623, n43624, n43625, n43626, n43627,
    n43628, n43629, n43630, n43631, n43632, n43633,
    n43634, n43635, n43636, n43637, n43638, n43639,
    n43640, n43641, n43642, n43643, n43644, n43645,
    n43646, n43647, n43648, n43649, n43650, n43651,
    n43652, n43653, n43654, n43655, n43656, n43657,
    n43658, n43659, n43660, n43661, n43662, n43663,
    n43664, n43665, n43666, n43667, n43668, n43669,
    n43670, n43671, n43672, n43673, n43674, n43675,
    n43676, n43677, n43679, n43680, n43681, n43682,
    n43683, n43684, n43685, n43686, n43687, n43688,
    n43689, n43690, n43691, n43692, n43693, n43694,
    n43696, n43697, n43698, n43699, n43700, n43701,
    n43702, n43703, n43704, n43705, n43706, n43707,
    n43708, n43709, n43710, n43711, n43712, n43713,
    n43714, n43715, n43716, n43717, n43718, n43719,
    n43720, n43721, n43722, n43723, n43724, n43725,
    n43726, n43727, n43728, n43729, n43730, n43731,
    n43732, n43733, n43734, n43735, n43737, n43738,
    n43739, n43740, n43741, n43742, n43743, n43744,
    n43745, n43746, n43747, n43748, n43749, n43750,
    n43751, n43752, n43753, n43754, n43755, n43756,
    n43757, n43758, n43759, n43760, n43761, n43762,
    n43763, n43764, n43765, n43766, n43767, n43768,
    n43769, n43770, n43771, n43772, n43773, n43774,
    n43775, n43776, n43777, n43778, n43779, n43780,
    n43781, n43782, n43783, n43784, n43785, n43786,
    n43787, n43788, n43789, n43790, n43791, n43792,
    n43793, n43794, n43795, n43796, n43797, n43798,
    n43799, n43800, n43801, n43802, n43803, n43804,
    n43805, n43806, n43807, n43808, n43809, n43810,
    n43811, n43812, n43813, n43814, n43815, n43816,
    n43817, n43818, n43819, n43820, n43821, n43822,
    n43823, n43824, n43825, n43826, n43827, n43828,
    n43829, n43830, n43831, n43832, n43833, n43834,
    n43835, n43836, n43837, n43838, n43839, n43840,
    n43841, n43842, n43843, n43844, n43845, n43846,
    n43847, n43848, n43849, n43850, n43851, n43852,
    n43853, n43854, n43855, n43856, n43857, n43858,
    n43859, n43860, n43861, n43862, n43863, n43864,
    n43865, n43866, n43867, n43868, n43869, n43870,
    n43871, n43872, n43873, n43874, n43875, n43876,
    n43877, n43878, n43880, n43881, n43882, n43883,
    n43884, n43885, n43886, n43887, n43888, n43889,
    n43890, n43891, n43892, n43893, n43894, n43895,
    n43896, n43897, n43898, n43899, n43900, n43901,
    n43902, n43903, n43904, n43905, n43906, n43907,
    n43908, n43909, n43910, n43911, n43912, n43913,
    n43914, n43915, n43916, n43917, n43918, n43919,
    n43920, n43921, n43922, n43923, n43924, n43925,
    n43926, n43927, n43928, n43929, n43930, n43931,
    n43932, n43933, n43934, n43935, n43936, n43937,
    n43938, n43939, n43940, n43941, n43942, n43943,
    n43944, n43945, n43946, n43947, n43948, n43949,
    n43950, n43951, n43952, n43953, n43954, n43955,
    n43956, n43957, n43958, n43959, n43960, n43961,
    n43962, n43963, n43964, n43965, n43966, n43967,
    n43968, n43969, n43970, n43971, n43972, n43973,
    n43974, n43975, n43976, n43977, n43978, n43979,
    n43980, n43981, n43982, n43983, n43984, n43985,
    n43986, n43987, n43988, n43989, n43990, n43991,
    n43992, n43993, n43994, n43995, n43996, n43997,
    n43998, n43999, n44000, n44001, n44002, n44003,
    n44004, n44005, n44006, n44007, n44008, n44009,
    n44010, n44011, n44012, n44013, n44014, n44015,
    n44016, n44017, n44018, n44019, n44020, n44021,
    n44022, n44023, n44024, n44025, n44026, n44027,
    n44028, n44029, n44030, n44031, n44032, n44033,
    n44034, n44035, n44036, n44037, n44038, n44039,
    n44040, n44041, n44042, n44043, n44044, n44045,
    n44046, n44047, n44048, n44049, n44050, n44051,
    n44052, n44053, n44054, n44055, n44056, n44057,
    n44058, n44059, n44060, n44061, n44062, n44063,
    n44064, n44065, n44066, n44067, n44068, n44069,
    n44070, n44071, n44072, n44073, n44074, n44075,
    n44076, n44077, n44078, n44079, n44080, n44081,
    n44082, n44083, n44084, n44085, n44086, n44087,
    n44088, n44089, n44090, n44091, n44092, n44093,
    n44094, n44095, n44096, n44097, n44098, n44099,
    n44100, n44101, n44102, n44103, n44104, n44105,
    n44106, n44107, n44108, n44109, n44110, n44111,
    n44112, n44113, n44114, n44115, n44116, n44117,
    n44118, n44119, n44120, n44121, n44122, n44123,
    n44124, n44125, n44126, n44127, n44128, n44129,
    n44130, n44131, n44132, n44133, n44134, n44135,
    n44136, n44137, n44138, n44139, n44140, n44141,
    n44142, n44143, n44144, n44145, n44146, n44147,
    n44148, n44149, n44150, n44151, n44152, n44153,
    n44154, n44155, n44156, n44157, n44158, n44159,
    n44160, n44161, n44162, n44163, n44164, n44165,
    n44166, n44167, n44168, n44169, n44170, n44171,
    n44172, n44173, n44174, n44175, n44176, n44177,
    n44178, n44179, n44180, n44181, n44182, n44183,
    n44184, n44185, n44186, n44187, n44188, n44189,
    n44190, n44191, n44192, n44193, n44194, n44195,
    n44196, n44197, n44198, n44199, n44200, n44201,
    n44202, n44203, n44204, n44205, n44206, n44207,
    n44208, n44209, n44210, n44211, n44212, n44213,
    n44214, n44215, n44216, n44217, n44218, n44219,
    n44220, n44221, n44222, n44223, n44224, n44225,
    n44226, n44227, n44228, n44229, n44230, n44231,
    n44232, n44233, n44234, n44235, n44236, n44237,
    n44238, n44239, n44240, n44241, n44242, n44243,
    n44244, n44245, n44246, n44247, n44248, n44249,
    n44250, n44251, n44252, n44253, n44254, n44255,
    n44256, n44257, n44258, n44259, n44260, n44261,
    n44262, n44263, n44264, n44265, n44266, n44267,
    n44268, n44269, n44270, n44271, n44272, n44273,
    n44274, n44275, n44276, n44277, n44278, n44279,
    n44280, n44281, n44282, n44283, n44284, n44285,
    n44286, n44287, n44288, n44289, n44290, n44291,
    n44292, n44293, n44294, n44295, n44296, n44297,
    n44298, n44299, n44300, n44301, n44302, n44303,
    n44304, n44305, n44306, n44307, n44308, n44309,
    n44310, n44311, n44312, n44313, n44314, n44315,
    n44316, n44317, n44318, n44319, n44320, n44321,
    n44322, n44323, n44324, n44325, n44326, n44327,
    n44328, n44329, n44330, n44331, n44332, n44333,
    n44334, n44335, n44336, n44337, n44338, n44339,
    n44340, n44341, n44342, n44343, n44344, n44345,
    n44346, n44347, n44348, n44349, n44350, n44351,
    n44352, n44353, n44354, n44355, n44356, n44357,
    n44358, n44359, n44360, n44361, n44362, n44363,
    n44364, n44365, n44366, n44367, n44368, n44369,
    n44370, n44371, n44372, n44373, n44374, n44375,
    n44376, n44377, n44378, n44379, n44380, n44381,
    n44382, n44383, n44384, n44385, n44386, n44387,
    n44388, n44389, n44390, n44391, n44392, n44393,
    n44394, n44395, n44396, n44397, n44398, n44399,
    n44400, n44401, n44402, n44403, n44404, n44405,
    n44406, n44407, n44408, n44409, n44410, n44411,
    n44412, n44413, n44414, n44415, n44416, n44417,
    n44418, n44419, n44420, n44421, n44422, n44423,
    n44424, n44425, n44426, n44427, n44428, n44429,
    n44430, n44431, n44432, n44433, n44434, n44435,
    n44436, n44437, n44438, n44439, n44440, n44441,
    n44442, n44443, n44444, n44445, n44446, n44447,
    n44448, n44449, n44450, n44451, n44452, n44453,
    n44454, n44455, n44456, n44457, n44458, n44459,
    n44460, n44461, n44462, n44463, n44464, n44465,
    n44466, n44467, n44468, n44469, n44470, n44471,
    n44472, n44473, n44474, n44475, n44476, n44477,
    n44478, n44479, n44480, n44481, n44482, n44483,
    n44484, n44485, n44486, n44487, n44488, n44489,
    n44490, n44491, n44492, n44493, n44494, n44495,
    n44496, n44497, n44498, n44499, n44500, n44501,
    n44502, n44503, n44504, n44505, n44506, n44507,
    n44508, n44509, n44510, n44511, n44512, n44513,
    n44514, n44515, n44516, n44517, n44518, n44519,
    n44520, n44521, n44522, n44523, n44524, n44525,
    n44526, n44527, n44528, n44529, n44530, n44531,
    n44532, n44533, n44534, n44535, n44536, n44537,
    n44538, n44539, n44540, n44541, n44542, n44543,
    n44544, n44545, n44546, n44547, n44548, n44549,
    n44550, n44551, n44552, n44553, n44554, n44555,
    n44556, n44557, n44558, n44559, n44560, n44561,
    n44562, n44563, n44564, n44565, n44566, n44567,
    n44568, n44569, n44570, n44571, n44572, n44573,
    n44574, n44575, n44576, n44577, n44578, n44579,
    n44580, n44581, n44582, n44583, n44584, n44585,
    n44586, n44587, n44588, n44589, n44590, n44591,
    n44592, n44593, n44594, n44595, n44596, n44597,
    n44598, n44599, n44600, n44601, n44602, n44603,
    n44604, n44605, n44606, n44607, n44608, n44609,
    n44610, n44611, n44612, n44613, n44614, n44615,
    n44616, n44617, n44618, n44619, n44620, n44621,
    n44622, n44623, n44624, n44625, n44626, n44627,
    n44628, n44629, n44630, n44631, n44632, n44633,
    n44634, n44635, n44636, n44637, n44638, n44639,
    n44640, n44641, n44642, n44643, n44644, n44645,
    n44646, n44647, n44648, n44649, n44650, n44651,
    n44652, n44653, n44654, n44655, n44656, n44657,
    n44658, n44659, n44660, n44661, n44662, n44663,
    n44664, n44665, n44666, n44667, n44668, n44669,
    n44670, n44671, n44672, n44673, n44674, n44675,
    n44676, n44677, n44678, n44679, n44680, n44681,
    n44682, n44683, n44684, n44685, n44686, n44687,
    n44688, n44689, n44690, n44691, n44692, n44693,
    n44694, n44695, n44696, n44697, n44698, n44699,
    n44700, n44701, n44702, n44703, n44704, n44705,
    n44706, n44707, n44708, n44709, n44710, n44711,
    n44712, n44713, n44714, n44715, n44716, n44717,
    n44718, n44719, n44720, n44721, n44722, n44723,
    n44724, n44725, n44726, n44727, n44728, n44729,
    n44730, n44731, n44732, n44733, n44734, n44735,
    n44736, n44737, n44738, n44739, n44740, n44741,
    n44742, n44743, n44744, n44745, n44746, n44747,
    n44748, n44749, n44750, n44751, n44752, n44753,
    n44754, n44755, n44756, n44757, n44758, n44759,
    n44760, n44761, n44762, n44763, n44764, n44765,
    n44766, n44767, n44768, n44769, n44770, n44771,
    n44772, n44773, n44774, n44775, n44776, n44777,
    n44778, n44779, n44780, n44781, n44782, n44783,
    n44784, n44785, n44786, n44787, n44788, n44789,
    n44790, n44791, n44792, n44793, n44794, n44795,
    n44796, n44797, n44798, n44799, n44800, n44801,
    n44802, n44803, n44804, n44805, n44806, n44807,
    n44808, n44809, n44810, n44811, n44812, n44813,
    n44814, n44815, n44816, n44817, n44818, n44819,
    n44820, n44821, n44822, n44823, n44824, n44825,
    n44826, n44827, n44828, n44829, n44830, n44831,
    n44832, n44833, n44834, n44835, n44836, n44837,
    n44838, n44839, n44840, n44841, n44842, n44843,
    n44844, n44845, n44846, n44847, n44848, n44849,
    n44850, n44851, n44852, n44853, n44854, n44855,
    n44856, n44857, n44858, n44859, n44860, n44861,
    n44862, n44863, n44864, n44865, n44866, n44867,
    n44868, n44869, n44870, n44871, n44872, n44873,
    n44874, n44875, n44876, n44877, n44878, n44879,
    n44880, n44881, n44882, n44883, n44884, n44885,
    n44886, n44887, n44888, n44889, n44890, n44891,
    n44892, n44893, n44894, n44895, n44896, n44897,
    n44898, n44899, n44900, n44901, n44902, n44903,
    n44904, n44905, n44906, n44907, n44908, n44909,
    n44910, n44911, n44912, n44913, n44914, n44915,
    n44916, n44917, n44918, n44919, n44920, n44921,
    n44922, n44923, n44924, n44925, n44926, n44927,
    n44928, n44929, n44930, n44931, n44932, n44933,
    n44934, n44935, n44936, n44937, n44938, n44939,
    n44940, n44941, n44942, n44943, n44944, n44945,
    n44946, n44947, n44948, n44949, n44950, n44951,
    n44952, n44953, n44954, n44955, n44956, n44957,
    n44958, n44959, n44960, n44961, n44962, n44963,
    n44964, n44965, n44966, n44967, n44968, n44969,
    n44970, n44971, n44972, n44973, n44974, n44975,
    n44976, n44977, n44978, n44979, n44980, n44981,
    n44982, n44983, n44984, n44985, n44986, n44987,
    n44988, n44989, n44990, n44991, n44992, n44993,
    n44994, n44995, n44996, n44997, n44998, n44999,
    n45000, n45001, n45002, n45003, n45004, n45005,
    n45006, n45007, n45008, n45009, n45010, n45011,
    n45012, n45013, n45014, n45015, n45016, n45017,
    n45018, n45019, n45020, n45021, n45022, n45023,
    n45024, n45025, n45026, n45027, n45028, n45029,
    n45030, n45031, n45032, n45033, n45034, n45035,
    n45036, n45037, n45038, n45039, n45040, n45041,
    n45042, n45043, n45044, n45045, n45046, n45047,
    n45048, n45049, n45050, n45051, n45052, n45053,
    n45054, n45055, n45056, n45057, n45058, n45059,
    n45060, n45061, n45062, n45063, n45064, n45065,
    n45066, n45067, n45068, n45069, n45070, n45071,
    n45072, n45073, n45074, n45075, n45076, n45077,
    n45078, n45079, n45080, n45081, n45082, n45083,
    n45084, n45085, n45086, n45087, n45088, n45089,
    n45090, n45091, n45092, n45093, n45094, n45095,
    n45096, n45097, n45098, n45099, n45100, n45101,
    n45102, n45103, n45104, n45105, n45106, n45107,
    n45108, n45109, n45110, n45111, n45112, n45113,
    n45114, n45115, n45116, n45117, n45118, n45119,
    n45120, n45121, n45122, n45123, n45124, n45125,
    n45126, n45127, n45128, n45129, n45130, n45131,
    n45132, n45133, n45134, n45135, n45136, n45137,
    n45138, n45139, n45140, n45141, n45142, n45143,
    n45144, n45145, n45146, n45147, n45148, n45149,
    n45150, n45151, n45152, n45153, n45154, n45155,
    n45156, n45157, n45158, n45159, n45160, n45161,
    n45162, n45163, n45164, n45165, n45166, n45167,
    n45168, n45169, n45170, n45171, n45172, n45173,
    n45174, n45175, n45176, n45177, n45178, n45179,
    n45180, n45181, n45182, n45183, n45184, n45185,
    n45186, n45187, n45188, n45189, n45190, n45191,
    n45192, n45193, n45194, n45195, n45196, n45197,
    n45198, n45199, n45200, n45201, n45202, n45203,
    n45204, n45205, n45206, n45207, n45208, n45209,
    n45210, n45211, n45212, n45213, n45214, n45215,
    n45216, n45217, n45218, n45219, n45220, n45221,
    n45222, n45223, n45224, n45225, n45226, n45227,
    n45228, n45229, n45230, n45231, n45232, n45233,
    n45234, n45235, n45236, n45237, n45238, n45239,
    n45240, n45241, n45242, n45243, n45244, n45245,
    n45246, n45247, n45248, n45249, n45250, n45251,
    n45252, n45253, n45254, n45255, n45256, n45257,
    n45258, n45259, n45260, n45261, n45262, n45263,
    n45264, n45265, n45266, n45267, n45268, n45269,
    n45270, n45271, n45272, n45273, n45274, n45275,
    n45276, n45277, n45278, n45279, n45280, n45281,
    n45282, n45283, n45284, n45285, n45286, n45287,
    n45288, n45289, n45290, n45291, n45292, n45293,
    n45294, n45295, n45296, n45297, n45298, n45299,
    n45300, n45301, n45302, n45303, n45304, n45305,
    n45306, n45307, n45308, n45309, n45310, n45311,
    n45312, n45313, n45314, n45315, n45316, n45317,
    n45318, n45319, n45320, n45321, n45322, n45323,
    n45324, n45325, n45326, n45327, n45328, n45329,
    n45330, n45331, n45332, n45333, n45334, n45335,
    n45336, n45337, n45338, n45339, n45340, n45341,
    n45342, n45343, n45344, n45345, n45346, n45347,
    n45348, n45349, n45350, n45351, n45352, n45353,
    n45354, n45355, n45356, n45357, n45358, n45359,
    n45360, n45361, n45362, n45363, n45364, n45365,
    n45366, n45367, n45368, n45369, n45370, n45371,
    n45372, n45373, n45374, n45375, n45376, n45377,
    n45378, n45379, n45380, n45381, n45382, n45383,
    n45384, n45385, n45386, n45387, n45388, n45389,
    n45390, n45391, n45392, n45393, n45394, n45395,
    n45396, n45397, n45398, n45399, n45400, n45401,
    n45402, n45403, n45404, n45405, n45406, n45407,
    n45408, n45409, n45410, n45411, n45412, n45413,
    n45414, n45415, n45416, n45417, n45418, n45419,
    n45420, n45421, n45422, n45423, n45424, n45425,
    n45426, n45427, n45428, n45429, n45430, n45431,
    n45432, n45433, n45434, n45435, n45436, n45437,
    n45438, n45439, n45440, n45441, n45442, n45443,
    n45444, n45445, n45446, n45447, n45448, n45449,
    n45450, n45451, n45452, n45453, n45454, n45455,
    n45456, n45457, n45458, n45459, n45460, n45461,
    n45462, n45463, n45464, n45465, n45466, n45467,
    n45468, n45469, n45470, n45471, n45472, n45473,
    n45474, n45475, n45476, n45477, n45478, n45479,
    n45480, n45481, n45482, n45483, n45484, n45485,
    n45486, n45487, n45488, n45489, n45490, n45491,
    n45492, n45493, n45494, n45495, n45496, n45497,
    n45498, n45499, n45500, n45501, n45502, n45503,
    n45504, n45505, n45506, n45507, n45508, n45509,
    n45510, n45511, n45512, n45513, n45514, n45515,
    n45516, n45517, n45518, n45519, n45520, n45521,
    n45522, n45523, n45524, n45525, n45526, n45527,
    n45528, n45529, n45530, n45531, n45532, n45533,
    n45534, n45535, n45536, n45537, n45538, n45539,
    n45540, n45541, n45542, n45543, n45544, n45545,
    n45546, n45547, n45548, n45549, n45550, n45551,
    n45552, n45553, n45554, n45555, n45556, n45557,
    n45558, n45559, n45560, n45561, n45562, n45563,
    n45564, n45565, n45566, n45567, n45568, n45569,
    n45570, n45571, n45572, n45573, n45574, n45575,
    n45576, n45577, n45578, n45579, n45580, n45581,
    n45582, n45583, n45584, n45585, n45586, n45587,
    n45588, n45589, n45590, n45591, n45592, n45593,
    n45594, n45595, n45596, n45597, n45598, n45599,
    n45600, n45601, n45602, n45603, n45604, n45605,
    n45606, n45607, n45608, n45609, n45610, n45611,
    n45612, n45613, n45614, n45615, n45616, n45617,
    n45618, n45619, n45620, n45621, n45622, n45623,
    n45624, n45625, n45626, n45627, n45628, n45629,
    n45630, n45631, n45632, n45633, n45634, n45635,
    n45636, n45637, n45638, n45639, n45640, n45641,
    n45642, n45643, n45644, n45645, n45646, n45647,
    n45648, n45649, n45650, n45651, n45652, n45653,
    n45654, n45655, n45656, n45657, n45658, n45659,
    n45660, n45661, n45662, n45663, n45664, n45665,
    n45666, n45667, n45668, n45669, n45670, n45671,
    n45672, n45673, n45674, n45675, n45676, n45677,
    n45678, n45679, n45680, n45681, n45682, n45683,
    n45684, n45685, n45686, n45687, n45688, n45689,
    n45690, n45691, n45692, n45693, n45694, n45695,
    n45696, n45697, n45698, n45699, n45700, n45701,
    n45702, n45703, n45704, n45705, n45706, n45707,
    n45708, n45709, n45710, n45711, n45712, n45713,
    n45714, n45715, n45716, n45717, n45718, n45719,
    n45720, n45721, n45722, n45723, n45724, n45725,
    n45726, n45727, n45728, n45729, n45730, n45731,
    n45732, n45733, n45734, n45735, n45736, n45737,
    n45738, n45739, n45740, n45741, n45742, n45743,
    n45744, n45745, n45746, n45747, n45748, n45749,
    n45750, n45751, n45752, n45753, n45754, n45755,
    n45756, n45757, n45758, n45759, n45760, n45761,
    n45762, n45763, n45764, n45765, n45766, n45767,
    n45768, n45769, n45770, n45771, n45772, n45773,
    n45774, n45775, n45776, n45777, n45778, n45779,
    n45780, n45781, n45782, n45783, n45784, n45785,
    n45786, n45787, n45788, n45789, n45790, n45791,
    n45792, n45793, n45794, n45795, n45796, n45797,
    n45798, n45799, n45800, n45801, n45802, n45803,
    n45804, n45805, n45806, n45807, n45808, n45809,
    n45810, n45811, n45812, n45813, n45814, n45815,
    n45816, n45817, n45818, n45819, n45820, n45821,
    n45822, n45823, n45824, n45825, n45826, n45827,
    n45828, n45829, n45830, n45831, n45832, n45833,
    n45834, n45835, n45836, n45837, n45838, n45839,
    n45840, n45841, n45842, n45843, n45844, n45845,
    n45846, n45847, n45848, n45849, n45850, n45851,
    n45852, n45853, n45854, n45855, n45856, n45857,
    n45858, n45859, n45860, n45861, n45862, n45863,
    n45864, n45865, n45866, n45867, n45868, n45869,
    n45870, n45871, n45872, n45873, n45874, n45875,
    n45876, n45877, n45878, n45879, n45880, n45881,
    n45882, n45883, n45884, n45885, n45886, n45887,
    n45888, n45889, n45890, n45891, n45892, n45893,
    n45894, n45895, n45896, n45897, n45898, n45899,
    n45900, n45901, n45902, n45903, n45904, n45905,
    n45906, n45907, n45908, n45909, n45910, n45911,
    n45912, n45913, n45914, n45915, n45916, n45917,
    n45918, n45919, n45920, n45921, n45922, n45923,
    n45924, n45925, n45926, n45927, n45928, n45929,
    n45930, n45931, n45932, n45933, n45934, n45935,
    n45936, n45937, n45938, n45939, n45940, n45941,
    n45942, n45943, n45944, n45945, n45946, n45947,
    n45948, n45949, n45950, n45951, n45952, n45953,
    n45954, n45955, n45956, n45957, n45958, n45960,
    n45961, n45962, n45963, n45964, n45965, n45966,
    n45967, n45968, n45969, n45970, n45971, n45972,
    n45973, n45974, n45975, n45976, n45977, n45978,
    n45979, n45980, n45981, n45982, n45983, n45984,
    n45985, n45986, n45987, n45988, n45989, n45990,
    n45991, n45992, n45993, n45994, n45995, n45996,
    n45997, n45998, n45999, n46000, n46001, n46002,
    n46003, n46004, n46005, n46006, n46007, n46008,
    n46009, n46010, n46011, n46012, n46013, n46014,
    n46015, n46016, n46017, n46018, n46019, n46020,
    n46021, n46022, n46023, n46024, n46025, n46026,
    n46027, n46028, n46029, n46030, n46031, n46032,
    n46033, n46034, n46035, n46036, n46037, n46038,
    n46039, n46040, n46041, n46042, n46043, n46044,
    n46045, n46046, n46047, n46048, n46049, n46050,
    n46051, n46052, n46053, n46054, n46055, n46056,
    n46057, n46058, n46059, n46060, n46061, n46062,
    n46063, n46064, n46065, n46066, n46067, n46068,
    n46069, n46070, n46071, n46072, n46073, n46074,
    n46075, n46076, n46077, n46078, n46079, n46080,
    n46081, n46082, n46083, n46084, n46085, n46086,
    n46087, n46088, n46089, n46090, n46091, n46092,
    n46093, n46094, n46095, n46096, n46097, n46098,
    n46099, n46100, n46101, n46102, n46103, n46104,
    n46105, n46106, n46107, n46108, n46109, n46110,
    n46111, n46112, n46113, n46114, n46115, n46116,
    n46117, n46118, n46119, n46120, n46121, n46122,
    n46123, n46124, n46125, n46126, n46127, n46128,
    n46129, n46130, n46131, n46132, n46133, n46134,
    n46135, n46136, n46137, n46138, n46139, n46140,
    n46141, n46142, n46143, n46144, n46145, n46146,
    n46147, n46148, n46149, n46150, n46151, n46152,
    n46153, n46154, n46155, n46156, n46157, n46158,
    n46159, n46160, n46161, n46162, n46163, n46164,
    n46165, n46166, n46167, n46168, n46169, n46170,
    n46171, n46172, n46173, n46174, n46175, n46176,
    n46177, n46178, n46179, n46180, n46181, n46182,
    n46183, n46184, n46185, n46186, n46187, n46188,
    n46189, n46190, n46191, n46192, n46193, n46194,
    n46195, n46196, n46197, n46198, n46199, n46200,
    n46201, n46202, n46203, n46204, n46205, n46206,
    n46207, n46208, n46209, n46210, n46211, n46212,
    n46213, n46214, n46215, n46216, n46217, n46218,
    n46219, n46220, n46221, n46222, n46223, n46224,
    n46225, n46226, n46227, n46228, n46229, n46230,
    n46231, n46232, n46233, n46234, n46235, n46236,
    n46237, n46238, n46239, n46240, n46241, n46242,
    n46243, n46244, n46245, n46246, n46247, n46248,
    n46249, n46250, n46251, n46252, n46253, n46254,
    n46255, n46256, n46257, n46258, n46259, n46260,
    n46261, n46262, n46263, n46264, n46265, n46266,
    n46267, n46268, n46269, n46270, n46271, n46272,
    n46273, n46274, n46275, n46276, n46277, n46278,
    n46279, n46280, n46281, n46282, n46283, n46284,
    n46285, n46286, n46287, n46288, n46289, n46290,
    n46291, n46292, n46293, n46294, n46295, n46296,
    n46297, n46298, n46299, n46300, n46301, n46302,
    n46303, n46304, n46305, n46306, n46307, n46308,
    n46309, n46310, n46311, n46312, n46313, n46314,
    n46315, n46316, n46317, n46318, n46319, n46320,
    n46321, n46322, n46323, n46324, n46325, n46326,
    n46327, n46328, n46329, n46330, n46331, n46332,
    n46333, n46334, n46335, n46336, n46337, n46338,
    n46339, n46340, n46341, n46342, n46343, n46344,
    n46345, n46346, n46348, n46349, n46350, n46351,
    n46352, n46353, n46354, n46355, n46356, n46357,
    n46358, n46359, n46360, n46361, n46362, n46363,
    n46364, n46365, n46366, n46367, n46368, n46369,
    n46370, n46371, n46372, n46373, n46374, n46375,
    n46376, n46377, n46378, n46379, n46380, n46381,
    n46382, n46383, n46384, n46385, n46386, n46387,
    n46388, n46389, n46390, n46391, n46392, n46393,
    n46394, n46395, n46396, n46397, n46398, n46399,
    n46400, n46401, n46402, n46403, n46404, n46405,
    n46406, n46407, n46408, n46409, n46410, n46411,
    n46412, n46413, n46414, n46415, n46416, n46417,
    n46418, n46419, n46420, n46421, n46422, n46423,
    n46424, n46425, n46426, n46427, n46428, n46429,
    n46430, n46431, n46432, n46433, n46434, n46435,
    n46436, n46437, n46438, n46439, n46440, n46441,
    n46442, n46443, n46444, n46445, n46446, n46447,
    n46448, n46449, n46450, n46451, n46452, n46453,
    n46454, n46455, n46456, n46457, n46458, n46459,
    n46460, n46461, n46462, n46463, n46464, n46465,
    n46466, n46467, n46468, n46469, n46470, n46471,
    n46472, n46473, n46474, n46475, n46476, n46477,
    n46478, n46479, n46480, n46481, n46482, n46483,
    n46484, n46485, n46486, n46487, n46488, n46489,
    n46490, n46491, n46492, n46493, n46494, n46495,
    n46496, n46497, n46498, n46499, n46500, n46501,
    n46502, n46503, n46504, n46505, n46506, n46507,
    n46508, n46509, n46510, n46511, n46512, n46513,
    n46514, n46515, n46516, n46517, n46518, n46519,
    n46520, n46521, n46522, n46523, n46524, n46525,
    n46526, n46527, n46528, n46529, n46530, n46531,
    n46532, n46533, n46534, n46535, n46536, n46537,
    n46538, n46539, n46540, n46541, n46542, n46543,
    n46544, n46545, n46546, n46547, n46548, n46549,
    n46550, n46551, n46552, n46553, n46554, n46555,
    n46556, n46557, n46558, n46559, n46560, n46561,
    n46562, n46563, n46564, n46565, n46566, n46567,
    n46568, n46569, n46570, n46571, n46572, n46573,
    n46574, n46575, n46576, n46577, n46578, n46579,
    n46580, n46581, n46582, n46583, n46584, n46585,
    n46586, n46587, n46588, n46589, n46590, n46591,
    n46592, n46593, n46594, n46595, n46596, n46597,
    n46598, n46599, n46600, n46601, n46602, n46603,
    n46604, n46605, n46606, n46607, n46608, n46609,
    n46610, n46611, n46612, n46613, n46614, n46615,
    n46616, n46617, n46618, n46619, n46620, n46621,
    n46622, n46623, n46624, n46625, n46626, n46627,
    n46628, n46629, n46630, n46631, n46632, n46633,
    n46634, n46635, n46636, n46637, n46638, n46639,
    n46640, n46641, n46642, n46643, n46644, n46645,
    n46646, n46647, n46648, n46649, n46650, n46651,
    n46652, n46653, n46654, n46655, n46656, n46657,
    n46658, n46659, n46660, n46661, n46662, n46663,
    n46664, n46665, n46666, n46667, n46668, n46669,
    n46670, n46671, n46672, n46673, n46674, n46675,
    n46676, n46677, n46678, n46679, n46680, n46681,
    n46682, n46683, n46684, n46685, n46686, n46687,
    n46688, n46689, n46690, n46691, n46692, n46693,
    n46694, n46695, n46696, n46697, n46698, n46699,
    n46700, n46701, n46702, n46703, n46704, n46705,
    n46706, n46707, n46708, n46709, n46710, n46711,
    n46712, n46713, n46714, n46715, n46716, n46717,
    n46718, n46719, n46720, n46721, n46722, n46723,
    n46724, n46725, n46726, n46727, n46728, n46729,
    n46730, n46731, n46732, n46733, n46734, n46735,
    n46736, n46737, n46738, n46739, n46740, n46741,
    n46742, n46743, n46744, n46745, n46746, n46747,
    n46748, n46749, n46750, n46751, n46752, n46753,
    n46754, n46755, n46756, n46757, n46758, n46759,
    n46760, n46761, n46762, n46763, n46764, n46765,
    n46766, n46767, n46768, n46769, n46770, n46771,
    n46772, n46773, n46774, n46775, n46776, n46777,
    n46778, n46779, n46780, n46781, n46782, n46783,
    n46784, n46785, n46786, n46787, n46788, n46789,
    n46790, n46791, n46792, n46793, n46794, n46795,
    n46796, n46797, n46798, n46799, n46800, n46801,
    n46802, n46803, n46804, n46805, n46806, n46807,
    n46808, n46809, n46810, n46811, n46812, n46813,
    n46814, n46815, n46816, n46817, n46818, n46819,
    n46820, n46821, n46822, n46823, n46824, n46825,
    n46826, n46827, n46828, n46829, n46830, n46831,
    n46832, n46833, n46834, n46835, n46836, n46837,
    n46838, n46839, n46840, n46841, n46842, n46843,
    n46844, n46845, n46846, n46847, n46848, n46849,
    n46850, n46851, n46852, n46853, n46854, n46855,
    n46856, n46857, n46858, n46859, n46860, n46861,
    n46862, n46863, n46864, n46865, n46866, n46867,
    n46868, n46869, n46870, n46871, n46872, n46873,
    n46874, n46875, n46876, n46877, n46878, n46879,
    n46880, n46881, n46882, n46883, n46884, n46885,
    n46886, n46887, n46888, n46889, n46890, n46891,
    n46892, n46893, n46894, n46895, n46896, n46897,
    n46898, n46899, n46900, n46901, n46902, n46903,
    n46904, n46905, n46906, n46907, n46908, n46909,
    n46910, n46911, n46912, n46913, n46914, n46915,
    n46916, n46917, n46918, n46919, n46920, n46921,
    n46922, n46923, n46924, n46925, n46926, n46927,
    n46928, n46929, n46930, n46931, n46932, n46933,
    n46934, n46935, n46936, n46937, n46938, n46939,
    n46940, n46941, n46942, n46943, n46944, n46945,
    n46946, n46947, n46948, n46949, n46950, n46951,
    n46952, n46953, n46954, n46955, n46956, n46957,
    n46958, n46959, n46960, n46961, n46962, n46963,
    n46964, n46965, n46966, n46967, n46968, n46969,
    n46970, n46971, n46972, n46973, n46974, n46975,
    n46976, n46977, n46978, n46979, n46980, n46981,
    n46982, n46983, n46984, n46985, n46986, n46987,
    n46988, n46989, n46990, n46991, n46992, n46993,
    n46994, n46995, n46996, n46997, n46998, n46999,
    n47000, n47001, n47002, n47003, n47004, n47005,
    n47006, n47007, n47008, n47009, n47010, n47011,
    n47012, n47013, n47014, n47015, n47016, n47017,
    n47018, n47019, n47020, n47021, n47022, n47023,
    n47024, n47025, n47026, n47027, n47028, n47029,
    n47030, n47031, n47032, n47033, n47034, n47035,
    n47036, n47037, n47038, n47039, n47040, n47041,
    n47042, n47043, n47044, n47045, n47046, n47047,
    n47048, n47049, n47050, n47051, n47052, n47053,
    n47054, n47055, n47056, n47057, n47058, n47059,
    n47060, n47061, n47062, n47063, n47064, n47065,
    n47066, n47067, n47068, n47069, n47070, n47071,
    n47072, n47073, n47074, n47075, n47076, n47077,
    n47078, n47079, n47080, n47081, n47082, n47083,
    n47084, n47085, n47086, n47087, n47088, n47089,
    n47090, n47091, n47092, n47093, n47094, n47095,
    n47096, n47097, n47098, n47099, n47100, n47101,
    n47102, n47103, n47104, n47105, n47106, n47107,
    n47108, n47109, n47110, n47111, n47112, n47113,
    n47114, n47115, n47116, n47117, n47118, n47119,
    n47120, n47121, n47122, n47123, n47124, n47125,
    n47126, n47127, n47128, n47129, n47130, n47131,
    n47132, n47133, n47134, n47135, n47136, n47137,
    n47138, n47139, n47140, n47141, n47142, n47143,
    n47144, n47145, n47146, n47147, n47148, n47149,
    n47150, n47151, n47152, n47153, n47154, n47155,
    n47156, n47157, n47158, n47159, n47160, n47161,
    n47162, n47163, n47164, n47165, n47166, n47167,
    n47168, n47169, n47170, n47171, n47172, n47173,
    n47174, n47175, n47176, n47177, n47178, n47179,
    n47180, n47181, n47182, n47183, n47184, n47185,
    n47186, n47187, n47188, n47189, n47190, n47191,
    n47192, n47193, n47194, n47195, n47196, n47197,
    n47198, n47199, n47200, n47201, n47202, n47203,
    n47204, n47205, n47206, n47207, n47208, n47209,
    n47210, n47211, n47212, n47213, n47214, n47215,
    n47216, n47217, n47218, n47219, n47220, n47221,
    n47222, n47223, n47224, n47225, n47226, n47227,
    n47228, n47229, n47230, n47231, n47232, n47233,
    n47234, n47235, n47236, n47237, n47238, n47239,
    n47240, n47241, n47242, n47243, n47244, n47245,
    n47246, n47247, n47248, n47249, n47250, n47251,
    n47252, n47253, n47254, n47255, n47256, n47257,
    n47258, n47259, n47260, n47261, n47262, n47263,
    n47264, n47265, n47266, n47267, n47268, n47269,
    n47270, n47271, n47272, n47273, n47274, n47275,
    n47276, n47277, n47278, n47279, n47280, n47281,
    n47282, n47283, n47284, n47285, n47286, n47287,
    n47288, n47289, n47290, n47291, n47292, n47293,
    n47294, n47295, n47296, n47297, n47298, n47299,
    n47300, n47301, n47302, n47303, n47304, n47305,
    n47306, n47307, n47308, n47309, n47310, n47311,
    n47312, n47313, n47314, n47315, n47316, n47317,
    n47318, n47319, n47320, n47321, n47322, n47323,
    n47324, n47325, n47326, n47327, n47328, n47329,
    n47330, n47331, n47332, n47333, n47334, n47335,
    n47336, n47337, n47338, n47339, n47340, n47341,
    n47342, n47343, n47344, n47345, n47346, n47347,
    n47348, n47349, n47350, n47351, n47352, n47353,
    n47354, n47355, n47356, n47357, n47358, n47359,
    n47360, n47361, n47362, n47363, n47364, n47365,
    n47366, n47367, n47368, n47369, n47370, n47371,
    n47372, n47373, n47374, n47375, n47376, n47377,
    n47378, n47379, n47380, n47381, n47382, n47383,
    n47384, n47385, n47386, n47387, n47388, n47389,
    n47390, n47391, n47392, n47393, n47394, n47395,
    n47396, n47397, n47398, n47399, n47400, n47401,
    n47402, n47403, n47404, n47405, n47406, n47407,
    n47408, n47409, n47410, n47411, n47412, n47413,
    n47414, n47415, n47416, n47417, n47418, n47419,
    n47420, n47421, n47422, n47423, n47424, n47425,
    n47426, n47427, n47428, n47429, n47430, n47431,
    n47432, n47433, n47434, n47435, n47436, n47437,
    n47438, n47439, n47440, n47441, n47442, n47443,
    n47444, n47445, n47446, n47447, n47448, n47449,
    n47450, n47451, n47452, n47453, n47454, n47455,
    n47456, n47457, n47458, n47459, n47460, n47461,
    n47462, n47463, n47464, n47465, n47466, n47467,
    n47468, n47469, n47470, n47471, n47472, n47473,
    n47474, n47475, n47476, n47477, n47478, n47479,
    n47480, n47481, n47482, n47483, n47484, n47486,
    n47487, n47488, n47489, n47490, n47491, n47492,
    n47493, n47494, n47495, n47496, n47497, n47498,
    n47499, n47500, n47501, n47502, n47503, n47504,
    n47505, n47506, n47507, n47508, n47509, n47510,
    n47511, n47512, n47513, n47514, n47515, n47516,
    n47517, n47518, n47519, n47520, n47521, n47522,
    n47523, n47524, n47526, n47527, n47528, n47529,
    n47530, n47531, n47532, n47533, n47534, n47535,
    n47536, n47537, n47538, n47539, n47540, n47541,
    n47542, n47543, n47544, n47545, n47546, n47548,
    n47549, n47550, n47551, n47552, n47553, n47554,
    n47555, n47556, n47557, n47558, n47559, n47560,
    n47561, n47562, n47563, n47564, n47565, n47566,
    n47567, n47568, n47569, n47570, n47571, n47572,
    n47573, n47574, n47575, n47576, n47577, n47579,
    n47580, n47581, n47582, n47583, n47584, n47585,
    n47586, n47587, n47588, n47589, n47590, n47591,
    n47592, n47593, n47594, n47595, n47596, n47597,
    n47598, n47599, n47600, n47601, n47602, n47603,
    n47604, n47605, n47606, n47607, n47608, n47609,
    n47610, n47611, n47612, n47613, n47614, n47615,
    n47616, n47617, n47618, n47619, n47620, n47621,
    n47622, n47623, n47624, n47625, n47626, n47627,
    n47628, n47629, n47630, n47631, n47632, n47633,
    n47634, n47635, n47636, n47637, n47638, n47639,
    n47640, n47641, n47642, n47643, n47644, n47645,
    n47646, n47647, n47648, n47649, n47650, n47651,
    n47652, n47653, n47654, n47655, n47656, n47657,
    n47658, n47659, n47660, n47661, n47662, n47663,
    n47664, n47665, n47666, n47667, n47668, n47669,
    n47670, n47671, n47672, n47673, n47674, n47675,
    n47676, n47677, n47678, n47679, n47680, n47681,
    n47682, n47683, n47684, n47685, n47686, n47687,
    n47688, n47689, n47690, n47691, n47692, n47693,
    n47694, n47695, n47696, n47697, n47698, n47699,
    n47700, n47701, n47702, n47703, n47704, n47705,
    n47706, n47707, n47708, n47709, n47710, n47711,
    n47712, n47713, n47714, n47715, n47716, n47717,
    n47718, n47719, n47720, n47721, n47722, n47723,
    n47724, n47725, n47726, n47727, n47728, n47729,
    n47730, n47731, n47732, n47733, n47734, n47735,
    n47736, n47737, n47738, n47739, n47740, n47741,
    n47742, n47743, n47744, n47745, n47746, n47747,
    n47748, n47749, n47750, n47751, n47752, n47753,
    n47754, n47755, n47756, n47757, n47758, n47759,
    n47760, n47761, n47762, n47763, n47764, n47765,
    n47766, n47767, n47768, n47769, n47770, n47771,
    n47772, n47773, n47774, n47775, n47776, n47777,
    n47778, n47779, n47780, n47781, n47782, n47783,
    n47784, n47785, n47786, n47787, n47788, n47789,
    n47790, n47791, n47792, n47793, n47794, n47795,
    n47796, n47797, n47798, n47799, n47800, n47801,
    n47802, n47803, n47804, n47805, n47806, n47807,
    n47808, n47809, n47810, n47811, n47812, n47813,
    n47814, n47815, n47816, n47817, n47819, n47820,
    n47821, n47822, n47823, n47824, n47825, n47827,
    n47828, n47829, n47830, n47831, n47832, n47833,
    n47835, n47836, n47837, n47838, n47839, n47840,
    n47841, n47842, n47843, n47844, n47845, n47846,
    n47847, n47848, n47849, n47850, n47851, n47852,
    n47853, n47854, n47855, n47856, n47857, n47858,
    n47859, n47860, n47861, n47862, n47863, n47864,
    n47865, n47866, n47867, n47868, n47869, n47870,
    n47871, n47872, n47873, n47874, n47875, n47876,
    n47877, n47878, n47879, n47880, n47881, n47882,
    n47883, n47884, n47885, n47886, n47887, n47888,
    n47889, n47890, n47891, n47892, n47893, n47894,
    n47895, n47896, n47897, n47898, n47899, n47900,
    n47901, n47902, n47903, n47904, n47905, n47906,
    n47907, n47908, n47909, n47910, n47911, n47912,
    n47913, n47914, n47915, n47916, n47917, n47918,
    n47919, n47920, n47921, n47922, n47923, n47924,
    n47925, n47926, n47927, n47928, n47929, n47930,
    n47931, n47932, n47933, n47934, n47935, n47936,
    n47937, n47938, n47939, n47940, n47941, n47942,
    n47943, n47944, n47945, n47946, n47947, n47948,
    n47949, n47950, n47951, n47952, n47953, n47954,
    n47956, n47957, n47958, n47959, n47960, n47961,
    n47963, n47964, n47965, n47966, n47967, n47968,
    n47969, n47971, n47972, n47973, n47974, n47975,
    n47976, n47978, n47979, n47980, n47981, n47982,
    n47983, n47985, n47986, n47987, n47988, n47989,
    n47990, n47991, n47992, n47993, n47994, n47995,
    n47996, n47997, n47998, n47999, n48000, n48001,
    n48002, n48003, n48004, n48005, n48006, n48008,
    n48009, n48010, n48011, n48012, n48013, n48014,
    n48015, n48016, n48017, n48018, n48019, n48020,
    n48021, n48022, n48023, n48024, n48025, n48026,
    n48027, n48028, n48029, n48030, n48031, n48032,
    n48033, n48034, n48035, n48036, n48037, n48038,
    n48039, n48040, n48041, n48042, n48043, n48044,
    n48045, n48046, n48047, n48048, n48049, n48050,
    n48051, n48052, n48053, n48054, n48055, n48056,
    n48057, n48058, n48059, n48060, n48061, n48062,
    n48063, n48064, n48065, n48066, n48067, n48068,
    n48069, n48070, n48071, n48072, n48073, n48074,
    n48075, n48076, n48077, n48078, n48079, n48080,
    n48081, n48082, n48083, n48084, n48085, n48086,
    n48087, n48088, n48089, n48090, n48091, n48092,
    n48093, n48094, n48095, n48096, n48097, n48098,
    n48099, n48100, n48101, n48102, n48103, n48104,
    n48105, n48106, n48107, n48108, n48109, n48110,
    n48111, n48112, n48113, n48114, n48115, n48116,
    n48117, n48119, n48120, n48121, n48122, n48123,
    n48124, n48125, n48126, n48127, n48128, n48129,
    n48130, n48131, n48132, n48133, n48134, n48135,
    n48136, n48137, n48138, n48140, n48141, n48142,
    n48143, n48144, n48145, n48146, n48147, n48148,
    n48149, n48150, n48151, n48152, n48153, n48154,
    n48155, n48156, n48157, n48158, n48159, n48160,
    n48161, n48162, n48163, n48164, n48165, n48166,
    n48167, n48168, n48169, n48171, n48172, n48173,
    n48175, n48176, n48177, n48178, n48179, n48180,
    n48181, n48182, n48183, n48184, n48185, n48187,
    n48188, n48189, n48190, n48191, n48192, n48193,
    n48194, n48195, n48196, n48197, n48198, n48199,
    n48200, n48202, n48203, n48204, n48205, n48206,
    n48207, n48208, n48209, n48210, n48211, n48212,
    n48213, n48214, n48215, n48216, n48217, n48218,
    n48219, n48220, n48221, n48222, n48223, n48224,
    n48226, n48227, n48228, n48229, n48230, n48231,
    n48232, n48233, n48234, n48235, n48236, n48237,
    n48239, n48240, n48241, n48242, n48243, n48244,
    n48245, n48246, n48247, n48248, n48249, n48250,
    n48251, n48252, n48253, n48254, n48255, n48256,
    n48257, n48258, n48259, n48260, n48261, n48262,
    n48263, n48264, n48265, n48266, n48267, n48268,
    n48269, n48270, n48271, n48272, n48273, n48274,
    n48275, n48276, n48277, n48278, n48279, n48280,
    n48281, n48282, n48283, n48284, n48285, n48286,
    n48287, n48288, n48289, n48290, n48291, n48292,
    n48293, n48294, n48295, n48296, n48297, n48298,
    n48299, n48300, n48301, n48302, n48303, n48304,
    n48305, n48306, n48307, n48308, n48309, n48310,
    n48311, n48312, n48313, n48314, n48315, n48316,
    n48317, n48318, n48319, n48320, n48321, n48322,
    n48323, n48324, n48325, n48326, n48327, n48328,
    n48329, n48330, n48331, n48332, n48333, n48334,
    n48335, n48336, n48337, n48338, n48339, n48340,
    n48341, n48342, n48343, n48344, n48345, n48346,
    n48347, n48348, n48349, n48350, n48351, n48352,
    n48353, n48354, n48355, n48356, n48357, n48358,
    n48359, n48360, n48361, n48362, n48363, n48364,
    n48365, n48366, n48367, n48368, n48369, n48370,
    n48371, n48372, n48373, n48374, n48375, n48376,
    n48377, n48378, n48379, n48380, n48381, n48382,
    n48383, n48384, n48385, n48386, n48387, n48388,
    n48389, n48390, n48391, n48392, n48393, n48394,
    n48395, n48396, n48397, n48398, n48399, n48400,
    n48401, n48402, n48403, n48404, n48405, n48406,
    n48407, n48408, n48409, n48410, n48411, n48412,
    n48413, n48414, n48415, n48416, n48417, n48418,
    n48419, n48420, n48421, n48422, n48423, n48424,
    n48425, n48426, n48427, n48428, n48429, n48430,
    n48431, n48432, n48433, n48434, n48435, n48436,
    n48437, n48438, n48439, n48440, n48441, n48442,
    n48443, n48444, n48445, n48446, n48447, n48449,
    n48450, n48451, n48452, n48453, n48454, n48455,
    n48456, n48457, n48458, n48459, n48460, n48461,
    n48462, n48463, n48464, n48465, n48467, n48469,
    n48470, n48471, n48472, n48473, n48474, n48475,
    n48476, n48477, n48478, n48479, n48480, n48481,
    n48482, n48483, n48484, n48485, n48486, n48487,
    n48488, n48490, n48491, n48492, n48493, n48494,
    n48495, n48496, n48497, n48498, n48499, n48500,
    n48501, n48502, n48504, n48505, n48506, n48507,
    n48508, n48509, n48510, n48511, n48512, n48513,
    n48514, n48515, n48516, n48517, n48518, n48519,
    n48520, n48521, n48522, n48523, n48524, n48525,
    n48526, n48527, n48528, n48529, n48530, n48531,
    n48532, n48533, n48534, n48535, n48536, n48537,
    n48538, n48539, n48540, n48541, n48542, n48543,
    n48544, n48545, n48546, n48548, n48549, n48550,
    n48551, n48552, n48553, n48554, n48555, n48556,
    n48557, n48558, n48559, n48560, n48561, n48562,
    n48563, n48564, n48565, n48566, n48567, n48568,
    n48569, n48570, n48571, n48572, n48573, n48574,
    n48575, n48577, n48578, n48579, n48580, n48581,
    n48582, n48583, n48584, n48585, n48586, n48587,
    n48588, n48589, n48590, n48591, n48592, n48593,
    n48594, n48595, n48597, n48598, n48599, n48600,
    n48601, n48602, n48603, n48604, n48605, n48606,
    n48607, n48608, n48609, n48610, n48611, n48612,
    n48613, n48614, n48615, n48616, n48617, n48618,
    n48619, n48621, n48623, n48624, n48625, n48626,
    n48627, n48628, n48629, n48630, n48631, n48632,
    n48633, n48634, n48635, n48636, n48637, n48638,
    n48639, n48641, n48642, n48643, n48644, n48645,
    n48646, n48647, n48648, n48649, n48650, n48651,
    n48652, n48653, n48654, n48655, n48656, n48658,
    n48659, n48660, n48661, n48662, n48663, n48664,
    n48665, n48666, n48667, n48668, n48669, n48670,
    n48671, n48672, n48673, n48674, n48675, n48676,
    n48677, n48678, n48680, n48681, n48682, n48683,
    n48684, n48686, n48687, n48688, n48689, n48690,
    n48691, n48692, n48693, n48694, n48695, n48696,
    n48697, n48698, n48699, n48700, n48701, n48702,
    n48703, n48704, n48705, n48706, n48707, n48708,
    n48709, n48710, n48711, n48712, n48713, n48714,
    n48715, n48716, n48718, n48719, n48720, n48721,
    n48722, n48723, n48724, n48725, n48726, n48727,
    n48728, n48729, n48730, n48732, n48733, n48734,
    n48735, n48736, n48737, n48739, n48740, n48741,
    n48743, n48744, n48745, n48746, n48747, n48748,
    n48749, n48750, n48751, n48752, n48753, n48755,
    n48756, n48757, n48758, n48759, n48760, n48761,
    n48762, n48763, n48764, n48765, n48766, n48767,
    n48768, n48769, n48770, n48772, n48773, n48774,
    n48775, n48776, n48777, n48778, n48779, n48780,
    n48781, n48782, n48783, n48784, n48785, n48786,
    n48787, n48788, n48789, n48790, n48793, n48794,
    n48795, n48796, n48797, n48798, n48799, n48800,
    n48801, n48802, n48803, n48804, n48805, n48806,
    n48807, n48808, n48809, n48810, n48811, n48812,
    n48813, n48814, n48815, n48816, n48817, n48818,
    n48819, n48820, n48821, n48822, n48823, n48824,
    n48825, n48826, n48827, n48828, n48829, n48830,
    n48831, n48832, n48833, n48834, n48836, n48837,
    n48838, n48840, n48841, n48842, n48843, n48844,
    n48845, n48846, n48847, n48848, n48849, n48851,
    n48852, n48853, n48854, n48855, n48856, n48857,
    n48858, n48859, n48861, n48862, n48863, n48864,
    n48865, n48866, n48867, n48868, n48869, n48871,
    n48872, n48873, n48874, n48876, n48877, n48878,
    n48880, n48881, n48882, n48883, n48884, n48885,
    n48886, n48889, n48890, n48891, n48892, n48893,
    n48894, n48895, n48897, n48898, n48899, n48900,
    n48902, n48903, n48904, n48905, n48906, n48907,
    n48908, n48909, n48910, n48911, n48912, n48913,
    n48914, n48915, n48916, n48917, n48918, n48919,
    n48920, n48921, n48922, n48923, n48924, n48925,
    n48926, n48927, n48928, n48929, n48930, n48931,
    n48932, n48933, n48935, n48936, n48937, n48938,
    n48940, n48941, n48942, n48943, n48944, n48945,
    n48946, n48947, n48948, n48949, n48951, n48952,
    n48953, n48954, n48955, n48958, n48959, n48961,
    n48962, n48964, n48966, n48967, n48969, n48970,
    n48971, n48972, n48973, n48974, n48975, n48976,
    n48977, n48978, n48979, n48980, n48981, n48982,
    n48983, n48984, n48985, n48986, n48987, n48988,
    n48989, n48990, n48991, n48993, n48994, n48995,
    n48996, n48997, n48998, n48999, n49000, n49001,
    n49002, n49003, n49004, n49005, n49006, n49007,
    n49008, n49009, n49010, n49011, n49012, n49013,
    n49014, n49015, n49016, n49017, n49018, n49019,
    n49020, n49021, n49022, n49023, n49024, n49025,
    n49026, n49027, n49028, n49029, n49030, n49031,
    n49032, n49033, n49035, n49036, n49037, n49038,
    n49039, n49040, n49041, n49042, n49043, n49044,
    n49045, n49046, n49047, n49048, n49049, n49050,
    n49051, n49052, n49053, n49054, n49055, n49056,
    n49057, n49058, n49059, n49060, n49061, n49062,
    n49063, n49064, n49065, n49066, n49067, n49068,
    n49069, n49070, n49071, n49072, n49073, n49074,
    n49075, n49076, n49077, n49078, n49079, n49080,
    n49081, n49082, n49083, n49084, n49085, n49086,
    n49087, n49088, n49089, n49090, n49091, n49092,
    n49093, n49094, n49095, n49096, n49097, n49098,
    n49099, n49100, n49101, n49102, n49103, n49104,
    n49105, n49106, n49107, n49108, n49109, n49110,
    n49111, n49112, n49113, n49114, n49115, n49116,
    n49117, n49118, n49119, n49120, n49121, n49122,
    n49123, n49124, n49125, n49126, n49127, n49128,
    n49129, n49130, n49131, n49132, n49133, n49134,
    n49135, n49136, n49137, n49138, n49139, n49140,
    n49141, n49142, n49143, n49144, n49145, n49146,
    n49147, n49148, n49149, n49150, n49151, n49152,
    n49153, n49154, n49155, n49156, n49157, n49158,
    n49159, n49160, n49161, n49162, n49163, n49164,
    n49165, n49166, n49167, n49168, n49169, n49170,
    n49171, n49172, n49173, n49174, n49175, n49176,
    n49177, n49178, n49179, n49180, n49181, n49182,
    n49183, n49184, n49185, n49186, n49187, n49188,
    n49189, n49190, n49191, n49192, n49193, n49194,
    n49195, n49196, n49197, n49198, n49199, n49200,
    n49201, n49202, n49203, n49204, n49205, n49206,
    n49207, n49208, n49209, n49210, n49211, n49212,
    n49213, n49214, n49215, n49216, n49217, n49218,
    n49219, n49220, n49221, n49222, n49223, n49224,
    n49225, n49226, n49227, n49228, n49229, n49230,
    n49231, n49232, n49233, n49234, n49235, n49236,
    n49237, n49238, n49239, n49240, n49241, n49242,
    n49243, n49244, n49245, n49246, n49247, n49248,
    n49249, n49250, n49251, n49252, n49253, n49254,
    n49255, n49256, n49257, n49258, n49259, n49260,
    n49261, n49262, n49263, n49264, n49265, n49266,
    n49267, n49268, n49269, n49270, n49271, n49272,
    n49273, n49274, n49275, n49276, n49277, n49278,
    n49279, n49280, n49281, n49282, n49283, n49284,
    n49285, n49286, n49287, n49288, n49289, n49290,
    n49291, n49292, n49293, n49294, n49295, n49296,
    n49297, n49298, n49299, n49300, n49301, n49302,
    n49303, n49304, n49305, n49306, n49307, n49308,
    n49309, n49310, n49311, n49312, n49313, n49314,
    n49315, n49316, n49317, n49318, n49319, n49320,
    n49321, n49322, n49323, n49324, n49325, n49326,
    n49327, n49328, n49329, n49330, n49331, n49332,
    n49333, n49334, n49335, n49336, n49337, n49338,
    n49339, n49340, n49341, n49342, n49343, n49344,
    n49345, n49346, n49347, n49348, n49349, n49350,
    n49351, n49352, n49353, n49354, n49355, n49356,
    n49357, n49358, n49359, n49360, n49361, n49362,
    n49363, n49364, n49365, n49366, n49367, n49368,
    n49369, n49370, n49371, n49372, n49373, n49374,
    n49375, n49376, n49377, n49378, n49379, n49380,
    n49381, n49382, n49383, n49384, n49385, n49386,
    n49387, n49388, n49389, n49390, n49391, n49392,
    n49393, n49394, n49395, n49396, n49397, n49398,
    n49399, n49400, n49401, n49402, n49403, n49404,
    n49405, n49406, n49407, n49408, n49409, n49410,
    n49411, n49412, n49413, n49414, n49415, n49416,
    n49417, n49418, n49419, n49420, n49421, n49422,
    n49423, n49424, n49425, n49426, n49427, n49428,
    n49429, n49430, n49431, n49432, n49433, n49434,
    n49435, n49436, n49437, n49438, n49439, n49440,
    n49441, n49442, n49443, n49444, n49445, n49446,
    n49447, n49448, n49449, n49450, n49451, n49452,
    n49453, n49454, n49455, n49456, n49457, n49458,
    n49459, n49460, n49461, n49462, n49463, n49464,
    n49465, n49466, n49467, n49468, n49469, n49470,
    n49471, n49472, n49473, n49474, n49475, n49476,
    n49477, n49478, n49479, n49480, n49481, n49482,
    n49483, n49484, n49485, n49486, n49487, n49488,
    n49489, n49490, n49491, n49492, n49493, n49494,
    n49495, n49496, n49497, n49498, n49499, n49500,
    n49501, n49502, n49503, n49504, n49505, n49506,
    n49507, n49508, n49509, n49510, n49511, n49512,
    n49513, n49514, n49515, n49516, n49517, n49518,
    n49519, n49520, n49521, n49522, n49523, n49524,
    n49525, n49526, n49527, n49528, n49529, n49530,
    n49531, n49532, n49533, n49534, n49535, n49536,
    n49537, n49538, n49539, n49540, n49541, n49542,
    n49543, n49544, n49545, n49546, n49547, n49548,
    n49549, n49550, n49551, n49552, n49553, n49554,
    n49555, n49556, n49557, n49558, n49559, n49560,
    n49561, n49562, n49563, n49564, n49565, n49566,
    n49567, n49568, n49569, n49570, n49571, n49572,
    n49573, n49574, n49575, n49576, n49577, n49578,
    n49579, n49580, n49581, n49582, n49583, n49584,
    n49585, n49586, n49587, n49588, n49589, n49590,
    n49591, n49593, n49594, n49595, n49596, n49597,
    n49598, n49599, n49600, n49601, n49602, n49603,
    n49604, n49605, n49606, n49607, n49608, n49609,
    n49610, n49611, n49612, n49613, n49614, n49615,
    n49616, n49617, n49618, n49619, n49620, n49621,
    n49622, n49623, n49624, n49625, n49626, n49627,
    n49628, n49629, n49630, n49631, n49632, n49633,
    n49634, n49635, n49636, n49637, n49638, n49639,
    n49640, n49641, n49642, n49643, n49644, n49645,
    n49646, n49647, n49648, n49649, n49650, n49651,
    n49652, n49653, n49654, n49655, n49656, n49657,
    n49658, n49659, n49660, n49661, n49662, n49663,
    n49664, n49665, n49666, n49667, n49668, n49669,
    n49670, n49671, n49672, n49673, n49674, n49675,
    n49676, n49677, n49678, n49679, n49680, n49681,
    n49682, n49683, n49684, n49685, n49686, n49687,
    n49688, n49689, n49690, n49691, n49692, n49693,
    n49694, n49695, n49696, n49697, n49698, n49699,
    n49700, n49701, n49702, n49703, n49704, n49705,
    n49706, n49707, n49708, n49709, n49710, n49711,
    n49712, n49713, n49714, n49715, n49716, n49717,
    n49718, n49719, n49720, n49721, n49722, n49723,
    n49724, n49725, n49726, n49727, n49728, n49729,
    n49730, n49731, n49732, n49733, n49734, n49735,
    n49736, n49737, n49738, n49739, n49740, n49741,
    n49742, n49743, n49744, n49745, n49746, n49747,
    n49748, n49749, n49750, n49751, n49752, n49753,
    n49754, n49755, n49756, n49757, n49758, n49759,
    n49760, n49761, n49762, n49763, n49764, n49765,
    n49766, n49767, n49768, n49769, n49770, n49771,
    n49772, n49773, n49774, n49775, n49776, n49777,
    n49778, n49779, n49780, n49781, n49782, n49783,
    n49784, n49785, n49786, n49787, n49788, n49789,
    n49790, n49791, n49792, n49793, n49794, n49795,
    n49796, n49797, n49798, n49799, n49800, n49801,
    n49802, n49803, n49804, n49805, n49806, n49807,
    n49808, n49809, n49810, n49811, n49812, n49813,
    n49814, n49815, n49816, n49817, n49818, n49819,
    n49820, n49821, n49822, n49823, n49824, n49825,
    n49826, n49827, n49828, n49829, n49830, n49831,
    n49832, n49833, n49834, n49835, n49836, n49837,
    n49838, n49839, n49840, n49841, n49842, n49843,
    n49844, n49845, n49846, n49847, n49848, n49849,
    n49850, n49851, n49852, n49853, n49854, n49855,
    n49856, n49857, n49858, n49859, n49860, n49861,
    n49862, n49863, n49864, n49865, n49866, n49867,
    n49868, n49869, n49870, n49871, n49872, n49873,
    n49874, n49875, n49876, n49877, n49878, n49879,
    n49880, n49881, n49882, n49883, n49884, n49885,
    n49886, n49887, n49888, n49889, n49890, n49891,
    n49892, n49893, n49894, n49895, n49896, n49897,
    n49898, n49899, n49900, n49901, n49902, n49903,
    n49904, n49905, n49906, n49908, n49909, n49910,
    n49911, n49912, n49913, n49914, n49915, n49916,
    n49917, n49918, n49919, n49920, n49921, n49922,
    n49923, n49924, n49925, n49926, n49927, n49928,
    n49929, n49930, n49931, n49932, n49933, n49934,
    n49935, n49936, n49937, n49938, n49939, n49940,
    n49941, n49942, n49943, n49944, n49945, n49946,
    n49947, n49948, n49949, n49950, n49951, n49952,
    n49953, n49954, n49955, n49956, n49957, n49958,
    n49959, n49960, n49961, n49962, n49963, n49964,
    n49965, n49966, n49967, n49968, n49969, n49970,
    n49971, n49972, n49973, n49974, n49975, n49976,
    n49977, n49978, n49979, n49980, n49981, n49982,
    n49983, n49984, n49985, n49986, n49987, n49988,
    n49989, n49990, n49991, n49992, n49993, n49994,
    n49995, n49996, n49997, n49998, n49999, n50000,
    n50001, n50002, n50003, n50004, n50005, n50006,
    n50007, n50008, n50009, n50010, n50011, n50012,
    n50013, n50014, n50015, n50016, n50017, n50018,
    n50019, n50020, n50021, n50022, n50023, n50024,
    n50025, n50026, n50027, n50028, n50029, n50030,
    n50031, n50032, n50033, n50034, n50035, n50036,
    n50037, n50038, n50039, n50040, n50041, n50042,
    n50043, n50044, n50045, n50046, n50047, n50048,
    n50049, n50050, n50051, n50052, n50053, n50054,
    n50055, n50056, n50057, n50058, n50059, n50060,
    n50061, n50062, n50063, n50064, n50065, n50066,
    n50067, n50068, n50069, n50070, n50071, n50072,
    n50073, n50074, n50075, n50076, n50077, n50078,
    n50079, n50080, n50081, n50082, n50083, n50084,
    n50085, n50086, n50087, n50088, n50089, n50090,
    n50091, n50092, n50093, n50094, n50095, n50096,
    n50097, n50098, n50099, n50100, n50101, n50102,
    n50103, n50104, n50105, n50106, n50107, n50108,
    n50109, n50110, n50111, n50112, n50113, n50114,
    n50115, n50116, n50117, n50118, n50119, n50120,
    n50121, n50122, n50123, n50124, n50125, n50126,
    n50127, n50128, n50129, n50130, n50131, n50132,
    n50133, n50134, n50135, n50136, n50137, n50138,
    n50139, n50140, n50141, n50142, n50143, n50144,
    n50145, n50146, n50147, n50148, n50149, n50150,
    n50151, n50152, n50153, n50154, n50155, n50156,
    n50157, n50158, n50159, n50160, n50161, n50162,
    n50163, n50164, n50165, n50166, n50167, n50168,
    n50169, n50170, n50171, n50172, n50173, n50174,
    n50175, n50176, n50177, n50178, n50179, n50180,
    n50181, n50182, n50183, n50184, n50185, n50186,
    n50187, n50188, n50189, n50190, n50191, n50192,
    n50193, n50194, n50195, n50196, n50197, n50198,
    n50199, n50200, n50201, n50202, n50203, n50204,
    n50205, n50206, n50207, n50208, n50209, n50210,
    n50211, n50212, n50213, n50214, n50215, n50216,
    n50217, n50218, n50219, n50220, n50221, n50222,
    n50223, n50224, n50225, n50226, n50227, n50228,
    n50229, n50231, n50232, n50233, n50234, n50235,
    n50236, n50237, n50238, n50239, n50240, n50241,
    n50242, n50243, n50244, n50245, n50246, n50247,
    n50248, n50249, n50250, n50251, n50252, n50253,
    n50254, n50255, n50256, n50257, n50258, n50259,
    n50260, n50261, n50262, n50263, n50264, n50265,
    n50266, n50267, n50268, n50269, n50270, n50271,
    n50272, n50273, n50274, n50275, n50276, n50277,
    n50278, n50279, n50280, n50281, n50282, n50283,
    n50284, n50285, n50286, n50287, n50288, n50289,
    n50290, n50291, n50292, n50293, n50294, n50295,
    n50296, n50297, n50298, n50299, n50300, n50301,
    n50302, n50303, n50304, n50305, n50306, n50307,
    n50308, n50309, n50310, n50311, n50312, n50313,
    n50314, n50315, n50316, n50317, n50318, n50319,
    n50320, n50321, n50322, n50323, n50324, n50325,
    n50326, n50327, n50328, n50329, n50330, n50331,
    n50332, n50333, n50334, n50335, n50336, n50337,
    n50338, n50339, n50340, n50341, n50342, n50343,
    n50344, n50345, n50346, n50347, n50348, n50349,
    n50350, n50351, n50352, n50353, n50354, n50355,
    n50356, n50357, n50358, n50359, n50360, n50361,
    n50362, n50363, n50364, n50365, n50366, n50367,
    n50368, n50369, n50370, n50371, n50372, n50373,
    n50374, n50375, n50376, n50377, n50378, n50379,
    n50380, n50381, n50382, n50383, n50384, n50385,
    n50386, n50387, n50388, n50389, n50390, n50391,
    n50392, n50393, n50394, n50395, n50396, n50397,
    n50398, n50399, n50400, n50401, n50402, n50403,
    n50404, n50405, n50406, n50407, n50408, n50409,
    n50410, n50411, n50412, n50413, n50414, n50415,
    n50416, n50417, n50418, n50419, n50420, n50421,
    n50422, n50423, n50424, n50425, n50426, n50427,
    n50428, n50429, n50430, n50431, n50432, n50433,
    n50434, n50435, n50436, n50437, n50438, n50439,
    n50440, n50441, n50442, n50443, n50444, n50445,
    n50446, n50447, n50448, n50449, n50450, n50451,
    n50452, n50453, n50454, n50455, n50456, n50457,
    n50458, n50459, n50460, n50461, n50462, n50463,
    n50464, n50465, n50466, n50467, n50468, n50469,
    n50470, n50471, n50472, n50473, n50474, n50475,
    n50476, n50477, n50478, n50479, n50480, n50481,
    n50482, n50483, n50484, n50485, n50486, n50487,
    n50488, n50489, n50490, n50491, n50492, n50493,
    n50494, n50495, n50496, n50498, n50499, n50500,
    n50501, n50502, n50503, n50504, n50505, n50506,
    n50507, n50508, n50509, n50510, n50511, n50512,
    n50513, n50514, n50515, n50516, n50517, n50518,
    n50519, n50520, n50521, n50522, n50523, n50524,
    n50525, n50526, n50527, n50528, n50529, n50530,
    n50531, n50532, n50533, n50534, n50535, n50536,
    n50537, n50538, n50539, n50540, n50541, n50542,
    n50543, n50544, n50545, n50546, n50547, n50548,
    n50549, n50550, n50551, n50552, n50553, n50554,
    n50555, n50556, n50557, n50558, n50559, n50560,
    n50561, n50562, n50563, n50564, n50565, n50566,
    n50567, n50568, n50569, n50570, n50571, n50572,
    n50573, n50574, n50575, n50576, n50577, n50578,
    n50579, n50580, n50581, n50582, n50583, n50584,
    n50585, n50586, n50587, n50588, n50589, n50590,
    n50591, n50592, n50593, n50594, n50595, n50596,
    n50597, n50598, n50599, n50600, n50601, n50602,
    n50603, n50604, n50605, n50606, n50607, n50608,
    n50609, n50610, n50611, n50612, n50613, n50614,
    n50615, n50616, n50617, n50618, n50619, n50620,
    n50621, n50622, n50623, n50624, n50625, n50626,
    n50627, n50628, n50629, n50630, n50631, n50632,
    n50633, n50634, n50635, n50636, n50637, n50638,
    n50639, n50640, n50641, n50642, n50643, n50644,
    n50645, n50646, n50647, n50648, n50649, n50650,
    n50651, n50652, n50653, n50654, n50655, n50656,
    n50657, n50658, n50659, n50660, n50661, n50662,
    n50663, n50664, n50665, n50666, n50667, n50668,
    n50669, n50670, n50671, n50672, n50673, n50674,
    n50675, n50676, n50677, n50678, n50679, n50680,
    n50681, n50682, n50683, n50684, n50685, n50686,
    n50687, n50688, n50689, n50690, n50691, n50692,
    n50693, n50694, n50695, n50696, n50697, n50698,
    n50699, n50700, n50701, n50702, n50703, n50704,
    n50705, n50706, n50707, n50708, n50709, n50710,
    n50711, n50712, n50713, n50714, n50715, n50716,
    n50717, n50718, n50719, n50720, n50721, n50722,
    n50723, n50724, n50725, n50726, n50727, n50728,
    n50729, n50730, n50731, n50732, n50733, n50734,
    n50735, n50736, n50737, n50738, n50739, n50740,
    n50741, n50742, n50743, n50744, n50745, n50746,
    n50747, n50748, n50749, n50750, n50751, n50752,
    n50753, n50754, n50755, n50756, n50757, n50758,
    n50759, n50760, n50761, n50763, n50764, n50765,
    n50766, n50767, n50768, n50769, n50770, n50771,
    n50772, n50773, n50774, n50775, n50776, n50777,
    n50778, n50779, n50780, n50781, n50782, n50783,
    n50784, n50785, n50786, n50787, n50788, n50789,
    n50790, n50791, n50792, n50793, n50794, n50795,
    n50796, n50797, n50798, n50799, n50800, n50801,
    n50802, n50803, n50804, n50805, n50806, n50807,
    n50808, n50809, n50810, n50811, n50812, n50813,
    n50814, n50815, n50816, n50817, n50818, n50819,
    n50820, n50821, n50822, n50823, n50824, n50825,
    n50826, n50827, n50828, n50829, n50830, n50831,
    n50832, n50833, n50834, n50835, n50836, n50837,
    n50838, n50839, n50840, n50841, n50842, n50843,
    n50844, n50845, n50846, n50847, n50848, n50849,
    n50850, n50851, n50852, n50853, n50854, n50855,
    n50856, n50857, n50858, n50859, n50860, n50861,
    n50862, n50863, n50864, n50865, n50866, n50867,
    n50868, n50869, n50870, n50871, n50872, n50873,
    n50874, n50875, n50876, n50877, n50878, n50879,
    n50880, n50881, n50882, n50883, n50884, n50885,
    n50886, n50887, n50888, n50889, n50890, n50891,
    n50892, n50893, n50894, n50895, n50896, n50897,
    n50898, n50899, n50900, n50901, n50902, n50903,
    n50904, n50905, n50906, n50907, n50908, n50909,
    n50910, n50911, n50912, n50913, n50914, n50915,
    n50916, n50917, n50918, n50919, n50920, n50921,
    n50922, n50923, n50924, n50925, n50926, n50927,
    n50928, n50929, n50930, n50931, n50932, n50933,
    n50934, n50935, n50936, n50937, n50938, n50939,
    n50940, n50941, n50942, n50943, n50944, n50945,
    n50946, n50947, n50948, n50949, n50950, n50951,
    n50952, n50953, n50954, n50955, n50956, n50957,
    n50958, n50959, n50960, n50961, n50962, n50963,
    n50964, n50965, n50966, n50967, n50968, n50969,
    n50970, n50971, n50972, n50973, n50974, n50975,
    n50976, n50977, n50978, n50979, n50980, n50981,
    n50982, n50983, n50984, n50985, n50986, n50987,
    n50988, n50989, n50990, n50991, n50992, n50993,
    n50994, n50995, n50996, n50997, n50998, n50999,
    n51000, n51001, n51002, n51003, n51004, n51005,
    n51006, n51007, n51008, n51009, n51010, n51011,
    n51012, n51013, n51014, n51015, n51016, n51017,
    n51018, n51019, n51020, n51021, n51022, n51023,
    n51024, n51025, n51026, n51027, n51028, n51029,
    n51030, n51031, n51032, n51033, n51034, n51035,
    n51036, n51037, n51038, n51039, n51040, n51041,
    n51042, n51043, n51044, n51045, n51046, n51047,
    n51048, n51049, n51050, n51051, n51052, n51053,
    n51054, n51055, n51056, n51057, n51058, n51059,
    n51060, n51061, n51062, n51063, n51064, n51065,
    n51066, n51067, n51068, n51069, n51070, n51071,
    n51072, n51073, n51074, n51075, n51076, n51077,
    n51078, n51079, n51080, n51081, n51082, n51083,
    n51084, n51085, n51086, n51087, n51088, n51089,
    n51090, n51091, n51092, n51093, n51094, n51095,
    n51096, n51097, n51098, n51099, n51100, n51101,
    n51102, n51103, n51104, n51105, n51106, n51107,
    n51108, n51109, n51110, n51111, n51112, n51113,
    n51114, n51115, n51116, n51117, n51118, n51119,
    n51120, n51121, n51122, n51123, n51124, n51125,
    n51126, n51127, n51128, n51129, n51130, n51131,
    n51132, n51133, n51134, n51135, n51136, n51137,
    n51138, n51139, n51140, n51141, n51142, n51143,
    n51144, n51145, n51146, n51147, n51148, n51149,
    n51150, n51151, n51152, n51153, n51154, n51155,
    n51156, n51157, n51158, n51159, n51160, n51161,
    n51162, n51163, n51164, n51165, n51166, n51167,
    n51168, n51169, n51170, n51171, n51172, n51173,
    n51174, n51175, n51176, n51177, n51178, n51179,
    n51180, n51181, n51182, n51183, n51184, n51185,
    n51186, n51187, n51188, n51189, n51190, n51191,
    n51192, n51193, n51194, n51195, n51196, n51197,
    n51198, n51199, n51200, n51201, n51202, n51203,
    n51204, n51205, n51206, n51207, n51208, n51209,
    n51210, n51211, n51212, n51213, n51214, n51215,
    n51216, n51217, n51218, n51219, n51220, n51221,
    n51222, n51223, n51224, n51225, n51226, n51227,
    n51228, n51229, n51230, n51231, n51232, n51233,
    n51234, n51235, n51236, n51237, n51238, n51239,
    n51240, n51241, n51242, n51243, n51244, n51245,
    n51246, n51247, n51248, n51249, n51250, n51251,
    n51252, n51253, n51254, n51255, n51256, n51257,
    n51258, n51259, n51260, n51261, n51262, n51263,
    n51264, n51265, n51266, n51267, n51268, n51269,
    n51270, n51271, n51272, n51273, n51274, n51275,
    n51276, n51277, n51278, n51279, n51280, n51281,
    n51282, n51283, n51284, n51285, n51286, n51287,
    n51288, n51289, n51290, n51291, n51292, n51293,
    n51294, n51295, n51296, n51297, n51298, n51299,
    n51300, n51301, n51302, n51303, n51304, n51305,
    n51306, n51307, n51308, n51309, n51310, n51311,
    n51312, n51313, n51314, n51315, n51316, n51317,
    n51318, n51319, n51320, n51321, n51322, n51323,
    n51324, n51325, n51326, n51327, n51328, n51329,
    n51331, n51332, n51333, n51334, n51335, n51336,
    n51337, n51338, n51339, n51340, n51341, n51342,
    n51343, n51344, n51345, n51346, n51347, n51348,
    n51349, n51350, n51351, n51352, n51353, n51354,
    n51355, n51356, n51357, n51358, n51359, n51360,
    n51361, n51362, n51363, n51364, n51365, n51366,
    n51367, n51368, n51369, n51370, n51371, n51372,
    n51373, n51374, n51375, n51376, n51377, n51378,
    n51379, n51380, n51381, n51382, n51383, n51384,
    n51385, n51386, n51387, n51388, n51389, n51390,
    n51391, n51392, n51393, n51394, n51395, n51396,
    n51397, n51398, n51399, n51400, n51401, n51402,
    n51403, n51404, n51405, n51406, n51407, n51408,
    n51409, n51410, n51411, n51412, n51413, n51414,
    n51415, n51416, n51417, n51418, n51419, n51420,
    n51421, n51422, n51423, n51424, n51425, n51426,
    n51427, n51428, n51429, n51430, n51431, n51432,
    n51433, n51434, n51435, n51436, n51437, n51438,
    n51439, n51440, n51441, n51442, n51443, n51444,
    n51445, n51446, n51447, n51448, n51449, n51450,
    n51451, n51452, n51453, n51454, n51455, n51456,
    n51457, n51458, n51459, n51460, n51461, n51462,
    n51463, n51464, n51465, n51466, n51467, n51468,
    n51469, n51470, n51471, n51472, n51473, n51474,
    n51475, n51476, n51477, n51478, n51479, n51480,
    n51481, n51482, n51483, n51484, n51485, n51486,
    n51487, n51488, n51489, n51490, n51491, n51492,
    n51493, n51494, n51495, n51496, n51497, n51498,
    n51499, n51500, n51501, n51502, n51503, n51504,
    n51505, n51506, n51507, n51508, n51509, n51510,
    n51511, n51512, n51513, n51514, n51515, n51516,
    n51517, n51518, n51519, n51520, n51521, n51522,
    n51523, n51524, n51525, n51526, n51527, n51528,
    n51529, n51530, n51531, n51532, n51533, n51534,
    n51535, n51536, n51537, n51538, n51539, n51540,
    n51541, n51542, n51543, n51544, n51545, n51546,
    n51547, n51548, n51549, n51550, n51551, n51552,
    n51553, n51554, n51555, n51556, n51557, n51558,
    n51559, n51560, n51561, n51562, n51563, n51565,
    n51566, n51567, n51568, n51569, n51570, n51571,
    n51572, n51573, n51574, n51575, n51576, n51577,
    n51578, n51579, n51580, n51581, n51582, n51583,
    n51584, n51585, n51586, n51587, n51588, n51589,
    n51590, n51591, n51592, n51593, n51594, n51595,
    n51596, n51597, n51598, n51599, n51600, n51601,
    n51602, n51603, n51604, n51605, n51606, n51607,
    n51608, n51609, n51610, n51611, n51612, n51613,
    n51614, n51615, n51616, n51617, n51618, n51619,
    n51620, n51621, n51622, n51623, n51624, n51625,
    n51626, n51627, n51628, n51629, n51630, n51631,
    n51632, n51633, n51634, n51635, n51636, n51637,
    n51638, n51639, n51640, n51641, n51642, n51643,
    n51644, n51645, n51646, n51647, n51648, n51649,
    n51650, n51651, n51652, n51653, n51654, n51655,
    n51656, n51658, n51659, n51660, n51661, n51662,
    n51663, n51664, n51665, n51666, n51667, n51668,
    n51669, n51670, n51671, n51672, n51673, n51674,
    n51675, n51676, n51677, n51678, n51679, n51680,
    n51681, n51682, n51683, n51684, n51685, n51686,
    n51687, n51688, n51689, n51690, n51691, n51692,
    n51693, n51694, n51695, n51696, n51697, n51698,
    n51699, n51700, n51701, n51702, n51703, n51704,
    n51705, n51706, n51707, n51708, n51709, n51710,
    n51711, n51712, n51713, n51714, n51715, n51716,
    n51717, n51718, n51719, n51720, n51721, n51722,
    n51723, n51724, n51725, n51726, n51727, n51728,
    n51729, n51730, n51731, n51732, n51733, n51734,
    n51735, n51736, n51737, n51738, n51739, n51740,
    n51741, n51742, n51743, n51744, n51745, n51746,
    n51747, n51748, n51749, n51750, n51751, n51752,
    n51753, n51754, n51755, n51756, n51757, n51758,
    n51759, n51760, n51761, n51762, n51763, n51764,
    n51765, n51766, n51767, n51768, n51769, n51770,
    n51771, n51772, n51773, n51774, n51775, n51776,
    n51777, n51778, n51779, n51780, n51781, n51782,
    n51783, n51784, n51785, n51786, n51787, n51788,
    n51789, n51790, n51791, n51792, n51793, n51794,
    n51795, n51796, n51797, n51798, n51799, n51800,
    n51801, n51802, n51803, n51804, n51805, n51806,
    n51807, n51808, n51809, n51810, n51811, n51812,
    n51813, n51814, n51815, n51816, n51817, n51818,
    n51819, n51820, n51821, n51822, n51823, n51824,
    n51825, n51826, n51827, n51828, n51829, n51830,
    n51831, n51832, n51833, n51834, n51835, n51836,
    n51837, n51838, n51839, n51840, n51841, n51842,
    n51843, n51844, n51845, n51846, n51847, n51848,
    n51849, n51850, n51851, n51852, n51853, n51854,
    n51855, n51856, n51857, n51858, n51859, n51860,
    n51861, n51862, n51863, n51864, n51865, n51866,
    n51867, n51868, n51869, n51870, n51871, n51872,
    n51873, n51874, n51875, n51876, n51877, n51878,
    n51879, n51880, n51881, n51882, n51883, n51884,
    n51885, n51886, n51887, n51888, n51889, n51890,
    n51891, n51892, n51893, n51894, n51895, n51896,
    n51897, n51898, n51899, n51900, n51901, n51902,
    n51903, n51904, n51905, n51906, n51907, n51908,
    n51909, n51910, n51911, n51912, n51913, n51914,
    n51915, n51916, n51917, n51918, n51919, n51920,
    n51921, n51922, n51923, n51924, n51925, n51926,
    n51927, n51928, n51929, n51930, n51931, n51932,
    n51933, n51934, n51935, n51936, n51937, n51938,
    n51939, n51940, n51941, n51942, n51943, n51944,
    n51945, n51946, n51947, n51948, n51949, n51950,
    n51951, n51952, n51953, n51954, n51955, n51956,
    n51957, n51958, n51959, n51960, n51961, n51962,
    n51963, n51964, n51965, n51966, n51967, n51968,
    n51969, n51970, n51971, n51972, n51973, n51974,
    n51975, n51976, n51977, n51978, n51979, n51980,
    n51981, n51982, n51983, n51984, n51985, n51986,
    n51987, n51988, n51989, n51990, n51991, n51992,
    n51993, n51994, n51995, n51996, n51997, n51998,
    n51999, n52000, n52001, n52002, n52003, n52004,
    n52005, n52006, n52007, n52008, n52009, n52010,
    n52011, n52012, n52013, n52014, n52015, n52016,
    n52017, n52018, n52019, n52020, n52021, n52022,
    n52023, n52024, n52025, n52026, n52027, n52028,
    n52029, n52030, n52031, n52032, n52033, n52034,
    n52035, n52036, n52037, n52038, n52039, n52040,
    n52041, n52042, n52043, n52044, n52045, n52046,
    n52047, n52048, n52049, n52050, n52051, n52052,
    n52053, n52054, n52055, n52056, n52057, n52058,
    n52059, n52060, n52061, n52062, n52063, n52064,
    n52065, n52066, n52067, n52068, n52069, n52070,
    n52071, n52072, n52073, n52074, n52075, n52076,
    n52077, n52078, n52079, n52080, n52081, n52082,
    n52083, n52084, n52085, n52086, n52087, n52088,
    n52089, n52090, n52091, n52092, n52093, n52094,
    n52095, n52096, n52097, n52098, n52099, n52100,
    n52101, n52102, n52103, n52104, n52105, n52106,
    n52107, n52108, n52109, n52110, n52111, n52112,
    n52113, n52114, n52115, n52116, n52117, n52118,
    n52119, n52120, n52121, n52122, n52123, n52124,
    n52125, n52126, n52127, n52128, n52129, n52130,
    n52131, n52132, n52133, n52134, n52135, n52136,
    n52137, n52138, n52139, n52140, n52141, n52142,
    n52143, n52144, n52145, n52146, n52147, n52148,
    n52149, n52150, n52151, n52152, n52153, n52154,
    n52155, n52156, n52157, n52158, n52159, n52160,
    n52161, n52162, n52163, n52164, n52165, n52166,
    n52167, n52168, n52169, n52170, n52171, n52172,
    n52173, n52174, n52175, n52176, n52177, n52178,
    n52179, n52180, n52181, n52182, n52183, n52184,
    n52185, n52186, n52187, n52188, n52189, n52190,
    n52191, n52192, n52193, n52194, n52195, n52196,
    n52197, n52198, n52199, n52200, n52201, n52202,
    n52203, n52204, n52205, n52206, n52207, n52208,
    n52209, n52210, n52211, n52212, n52213, n52214,
    n52215, n52216, n52217, n52218, n52219, n52220,
    n52221, n52222, n52223, n52224, n52225, n52226,
    n52227, n52228, n52229, n52230, n52231, n52232,
    n52233, n52234, n52235, n52236, n52237, n52238,
    n52239, n52240, n52241, n52242, n52243, n52244,
    n52245, n52246, n52247, n52248, n52249, n52250,
    n52251, n52252, n52253, n52254, n52255, n52256,
    n52257, n52258, n52259, n52260, n52261, n52262,
    n52263, n52264, n52265, n52266, n52267, n52268,
    n52269, n52270, n52271, n52272, n52273, n52274,
    n52275, n52276, n52277, n52278, n52279, n52280,
    n52281, n52282, n52283, n52284, n52285, n52286,
    n52287, n52289, n52290, n52291, n52292, n52293,
    n52294, n52295, n52296, n52297, n52298, n52299,
    n52300, n52301, n52302, n52303, n52304, n52305,
    n52306, n52307, n52308, n52309, n52310, n52311,
    n52312, n52313, n52314, n52315, n52316, n52317,
    n52318, n52319, n52320, n52321, n52322, n52323,
    n52324, n52325, n52326, n52327, n52328, n52329,
    n52330, n52331, n52332, n52333, n52334, n52335,
    n52336, n52337, n52338, n52339, n52340, n52341,
    n52342, n52343, n52344, n52345, n52346, n52347,
    n52348, n52349, n52350, n52351, n52352, n52353,
    n52354, n52355, n52356, n52357, n52358, n52359,
    n52360, n52361, n52362, n52363, n52364, n52365,
    n52366, n52367, n52368, n52369, n52370, n52371,
    n52372, n52373, n52374, n52375, n52376, n52377,
    n52378, n52379, n52380, n52381, n52382, n52383,
    n52384, n52385, n52386, n52387, n52388, n52389,
    n52390, n52391, n52392, n52393, n52394, n52395,
    n52396, n52397, n52398, n52399, n52400, n52401,
    n52402, n52403, n52404, n52405, n52406, n52407,
    n52408, n52409, n52410, n52411, n52412, n52413,
    n52414, n52415, n52416, n52417, n52418, n52419,
    n52420, n52421, n52422, n52423, n52424, n52425,
    n52426, n52427, n52428, n52429, n52430, n52431,
    n52432, n52433, n52434, n52435, n52436, n52437,
    n52438, n52439, n52440, n52441, n52442, n52443,
    n52444, n52445, n52446, n52447, n52448, n52449,
    n52450, n52451, n52452, n52453, n52454, n52455,
    n52456, n52457, n52458, n52459, n52460, n52461,
    n52462, n52463, n52464, n52465, n52466, n52467,
    n52468, n52469, n52470, n52471, n52472, n52473,
    n52474, n52475, n52476, n52477, n52478, n52479,
    n52480, n52481, n52482, n52483, n52484, n52485,
    n52486, n52487, n52488, n52489, n52490, n52491,
    n52492, n52493, n52494, n52495, n52496, n52497,
    n52498, n52499, n52500, n52501, n52502, n52503,
    n52504, n52505, n52506, n52507, n52508, n52509,
    n52510, n52511, n52512, n52513, n52514, n52515,
    n52517, n52518, n52519, n52520, n52521, n52522,
    n52523, n52524, n52525, n52526, n52527, n52528,
    n52529, n52530, n52531, n52532, n52533, n52534,
    n52535, n52536, n52537, n52538, n52539, n52540,
    n52541, n52542, n52543, n52544, n52545, n52546,
    n52547, n52548, n52549, n52550, n52551, n52552,
    n52553, n52554, n52555, n52556, n52557, n52558,
    n52559, n52560, n52561, n52562, n52563, n52564,
    n52565, n52566, n52567, n52568, n52569, n52570,
    n52571, n52572, n52573, n52574, n52575, n52576,
    n52577, n52578, n52579, n52580, n52581, n52582,
    n52583, n52584, n52585, n52586, n52587, n52588,
    n52589, n52590, n52591, n52592, n52593, n52594,
    n52595, n52596, n52597, n52598, n52599, n52600,
    n52601, n52602, n52603, n52604, n52605, n52606,
    n52607, n52608, n52609, n52610, n52611, n52612,
    n52613, n52614, n52615, n52616, n52617, n52618,
    n52619, n52620, n52621, n52622, n52623, n52624,
    n52625, n52626, n52627, n52628, n52629, n52630,
    n52631, n52632, n52633, n52634, n52635, n52636,
    n52637, n52638, n52639, n52640, n52641, n52642,
    n52643, n52644, n52645, n52646, n52647, n52648,
    n52649, n52650, n52651, n52652, n52653, n52654,
    n52655, n52656, n52657, n52658, n52659, n52660,
    n52661, n52662, n52663, n52664, n52665, n52666,
    n52667, n52668, n52669, n52670, n52671, n52672,
    n52673, n52674, n52675, n52676, n52677, n52678,
    n52679, n52680, n52681, n52682, n52683, n52684,
    n52685, n52686, n52687, n52688, n52689, n52690,
    n52691, n52692, n52693, n52694, n52695, n52696,
    n52697, n52698, n52699, n52700, n52701, n52702,
    n52703, n52704, n52705, n52706, n52707, n52708,
    n52709, n52710, n52711, n52712, n52713, n52714,
    n52715, n52716, n52717, n52718, n52719, n52720,
    n52721, n52722, n52723, n52724, n52725, n52726,
    n52727, n52728, n52729, n52730, n52731, n52732,
    n52733, n52734, n52735, n52736, n52737, n52738,
    n52739, n52740, n52741, n52742, n52743, n52744,
    n52745, n52746, n52747, n52748, n52749, n52750,
    n52751, n52752, n52753, n52754, n52755, n52756,
    n52757, n52758, n52759, n52760, n52761, n52762,
    n52763, n52764, n52765, n52766, n52767, n52768,
    n52769, n52770, n52771, n52772, n52773, n52774,
    n52775, n52776, n52777, n52778, n52779, n52780,
    n52781, n52782, n52783, n52784, n52785, n52786,
    n52787, n52788, n52789, n52790, n52791, n52792,
    n52793, n52794, n52795, n52796, n52797, n52798,
    n52799, n52800, n52801, n52802, n52803, n52804,
    n52805, n52806, n52807, n52808, n52809, n52810,
    n52811, n52812, n52813, n52814, n52815, n52816,
    n52817, n52818, n52819, n52820, n52821, n52822,
    n52823, n52824, n52825, n52826, n52827, n52828,
    n52829, n52830, n52831, n52832, n52833, n52834,
    n52835, n52836, n52837, n52838, n52839, n52840,
    n52841, n52842, n52843, n52844, n52845, n52846,
    n52847, n52848, n52849, n52850, n52851, n52852,
    n52853, n52854, n52855, n52856, n52857, n52858,
    n52859, n52860, n52861, n52862, n52863, n52864,
    n52865, n52866, n52867, n52868, n52869, n52870,
    n52871, n52872, n52873, n52874, n52875, n52876,
    n52877, n52878, n52879, n52880, n52881, n52882,
    n52883, n52884, n52885, n52886, n52887, n52888,
    n52889, n52890, n52891, n52892, n52893, n52894,
    n52895, n52896, n52897, n52898, n52899, n52900,
    n52901, n52902, n52903, n52904, n52905, n52906,
    n52907, n52908, n52909, n52910, n52911, n52912,
    n52913, n52914, n52915, n52916, n52917, n52918,
    n52919, n52920, n52921, n52922, n52923, n52924,
    n52925, n52926, n52927, n52928, n52929, n52930,
    n52931, n52932, n52933, n52934, n52935, n52936,
    n52937, n52938, n52939, n52940, n52941, n52942,
    n52943, n52944, n52945, n52946, n52947, n52948,
    n52949, n52950, n52951, n52952, n52953, n52954,
    n52955, n52956, n52957, n52958, n52959, n52960,
    n52961, n52962, n52963, n52964, n52965, n52966,
    n52967, n52968, n52969, n52970, n52971, n52972,
    n52973, n52974, n52975, n52976, n52977, n52978,
    n52979, n52980, n52981, n52982, n52983, n52984,
    n52985, n52986, n52987, n52988, n52989, n52990,
    n52991, n52992, n52993, n52994, n52995, n52996,
    n52997, n52998, n52999, n53000, n53001, n53002,
    n53003, n53004, n53005, n53006, n53007, n53008,
    n53009, n53010, n53011, n53012, n53013, n53014,
    n53015, n53016, n53017, n53018, n53019, n53020,
    n53021, n53022, n53023, n53024, n53025, n53026,
    n53027, n53028, n53029, n53030, n53031, n53032,
    n53033, n53034, n53035, n53036, n53037, n53038,
    n53039, n53040, n53041, n53042, n53043, n53044,
    n53045, n53046, n53047, n53048, n53049, n53050,
    n53051, n53052, n53053, n53054, n53055, n53056,
    n53057, n53058, n53059, n53060, n53061, n53062,
    n53063, n53064, n53065, n53066, n53067, n53068,
    n53069, n53070, n53071, n53072, n53073, n53074,
    n53075, n53076, n53077, n53078, n53079, n53080,
    n53081, n53082, n53083, n53084, n53085, n53086,
    n53087, n53088, n53089, n53090, n53091, n53092,
    n53093, n53094, n53095, n53096, n53097, n53098,
    n53099, n53100, n53101, n53102, n53103, n53104,
    n53105, n53106, n53107, n53108, n53109, n53110,
    n53111, n53112, n53113, n53114, n53115, n53116,
    n53117, n53118, n53119, n53120, n53121, n53122,
    n53123, n53124, n53125, n53126, n53127, n53128,
    n53129, n53130, n53131, n53132, n53133, n53134,
    n53135, n53136, n53137, n53138, n53139, n53140,
    n53141, n53142, n53143, n53144, n53145, n53146,
    n53147, n53148, n53149, n53150, n53151, n53152,
    n53153, n53154, n53155, n53156, n53157, n53158,
    n53159, n53160, n53161, n53162, n53163, n53164,
    n53165, n53166, n53167, n53168, n53169, n53170,
    n53171, n53172, n53173, n53174, n53175, n53176,
    n53177, n53178, n53179, n53180, n53181, n53182,
    n53183, n53184, n53185, n53186, n53187, n53188,
    n53189, n53190, n53191, n53192, n53193, n53194,
    n53195, n53196, n53197, n53198, n53199, n53200,
    n53201, n53202, n53203, n53204, n53205, n53206,
    n53207, n53208, n53209, n53210, n53211, n53212,
    n53213, n53214, n53215, n53216, n53217, n53218,
    n53219, n53220, n53221, n53222, n53223, n53224,
    n53225, n53226, n53227, n53228, n53229, n53230,
    n53231, n53232, n53233, n53234, n53235, n53236,
    n53237, n53238, n53239, n53240, n53241, n53242,
    n53243, n53244, n53245, n53246, n53247, n53248,
    n53249, n53250, n53251, n53252, n53253, n53254,
    n53255, n53256, n53257, n53258, n53259, n53260,
    n53261, n53262, n53263, n53264, n53265, n53266,
    n53267, n53268, n53269, n53270, n53271, n53272,
    n53273, n53274, n53275, n53276, n53277, n53278,
    n53279, n53280, n53281, n53282, n53283, n53284,
    n53285, n53286, n53287, n53288, n53289, n53290,
    n53291, n53292, n53293, n53294, n53295, n53296,
    n53297, n53298, n53299, n53300, n53301, n53302,
    n53303, n53304, n53305, n53306, n53307, n53308,
    n53309, n53310, n53311, n53312, n53313, n53314,
    n53315, n53316, n53317, n53318, n53319, n53320,
    n53321, n53322, n53323, n53324, n53325, n53326,
    n53327, n53328, n53329, n53330, n53331, n53332,
    n53333, n53334, n53335, n53336, n53337, n53338,
    n53339, n53340, n53341, n53342, n53343, n53344,
    n53345, n53346, n53347, n53348, n53349, n53350,
    n53351, n53352, n53353, n53354, n53355, n53356,
    n53357, n53358, n53359, n53360, n53361, n53362,
    n53363, n53364, n53365, n53366, n53367, n53368,
    n53369, n53370, n53371, n53372, n53373, n53374,
    n53375, n53376, n53377, n53378, n53379, n53380,
    n53381, n53382, n53383, n53384, n53385, n53386,
    n53387, n53388, n53389, n53390, n53391, n53392,
    n53393, n53394, n53395, n53396, n53397, n53398,
    n53399, n53400, n53401, n53402, n53403, n53404,
    n53405, n53406, n53407, n53408, n53409, n53410,
    n53411, n53412, n53413, n53414, n53415, n53416,
    n53417, n53418, n53419, n53420, n53421, n53422,
    n53423, n53424, n53425, n53426, n53427, n53428,
    n53429, n53430, n53431, n53432, n53433, n53434,
    n53435, n53436, n53437, n53438, n53439, n53440,
    n53441, n53442, n53443, n53444, n53445, n53446,
    n53447, n53448, n53449, n53450, n53451, n53452,
    n53453, n53454, n53455, n53456, n53457, n53458,
    n53459, n53460, n53461, n53462, n53463, n53464,
    n53465, n53466, n53467, n53468, n53469, n53470,
    n53471, n53472, n53473, n53474, n53475, n53476,
    n53477, n53478, n53479, n53480, n53481, n53482,
    n53483, n53484, n53485, n53486, n53487, n53488,
    n53489, n53490, n53491, n53492, n53493, n53494,
    n53495, n53496, n53497, n53498, n53499, n53500,
    n53501, n53502, n53503, n53504, n53505, n53506,
    n53507, n53508, n53509, n53510, n53511, n53512,
    n53513, n53514, n53515, n53516, n53517, n53518,
    n53519, n53520, n53521, n53522, n53523, n53524,
    n53525, n53526, n53527, n53528, n53529, n53530,
    n53531, n53532, n53533, n53534, n53535, n53536,
    n53537, n53538, n53539, n53540, n53541, n53542,
    n53543, n53544, n53545, n53546, n53547, n53548,
    n53549, n53550, n53551, n53552, n53553, n53554,
    n53555, n53556, n53557, n53558, n53559, n53560,
    n53561, n53562, n53563, n53564, n53565, n53566,
    n53567, n53568, n53569, n53570, n53571, n53572,
    n53573, n53574, n53575, n53576, n53577, n53578,
    n53579, n53580, n53581, n53582, n53583, n53584,
    n53585, n53586, n53587, n53588, n53589, n53590,
    n53591, n53592, n53593, n53594, n53595, n53596,
    n53597, n53598, n53599, n53600, n53601, n53602,
    n53603, n53604, n53605, n53606, n53607, n53608,
    n53609, n53610, n53611, n53612, n53613, n53614,
    n53615, n53616, n53617, n53618, n53619, n53620,
    n53622, n53623, n53624, n53625, n53626, n53627,
    n53628, n53629, n53630, n53631, n53632, n53633,
    n53634, n53635, n53636, n53637, n53638, n53639,
    n53640, n53641, n53642, n53643, n53644, n53645,
    n53646, n53647, n53648, n53649, n53650, n53651,
    n53652, n53653, n53654, n53655, n53656, n53657,
    n53658, n53659, n53660, n53661, n53662, n53663,
    n53664, n53665, n53666, n53667, n53668, n53669,
    n53670, n53671, n53672, n53673, n53674, n53675,
    n53676, n53677, n53678, n53679, n53680, n53681,
    n53682, n53683, n53684, n53685, n53686, n53687,
    n53688, n53689, n53690, n53691, n53692, n53693,
    n53694, n53695, n53696, n53697, n53698, n53699,
    n53700, n53701, n53702, n53703, n53704, n53705,
    n53706, n53707, n53708, n53709, n53710, n53711,
    n53712, n53713, n53714, n53715, n53716, n53717,
    n53718, n53719, n53720, n53721, n53722, n53723,
    n53724, n53725, n53726, n53727, n53728, n53729,
    n53730, n53731, n53732, n53733, n53734, n53735,
    n53736, n53738, n53739, n53740, n53741, n53742,
    n53743, n53744, n53745, n53746, n53747, n53748,
    n53749, n53750, n53751, n53752, n53753, n53754,
    n53755, n53756, n53757, n53758, n53759, n53760,
    n53761, n53762, n53763, n53764, n53765, n53766,
    n53767, n53768, n53769, n53770, n53771, n53772,
    n53773, n53774, n53775, n53776, n53777, n53778,
    n53779, n53780, n53781, n53782, n53783, n53784,
    n53785, n53786, n53787, n53788, n53789, n53790,
    n53791, n53792, n53793, n53794, n53795, n53796,
    n53797, n53798, n53799, n53800, n53801, n53802,
    n53803, n53804, n53805, n53806, n53807, n53808,
    n53809, n53810, n53811, n53812, n53813, n53814,
    n53815, n53816, n53817, n53818, n53819, n53820,
    n53821, n53822, n53823, n53824, n53825, n53826,
    n53827, n53828, n53829, n53830, n53831, n53832,
    n53833, n53834, n53835, n53836, n53837, n53838,
    n53839, n53840, n53841, n53842, n53843, n53844,
    n53845, n53846, n53847, n53848, n53849, n53850,
    n53851, n53852, n53853, n53854, n53855, n53856,
    n53857, n53858, n53859, n53860, n53861, n53862,
    n53863, n53864, n53865, n53866, n53867, n53868,
    n53869, n53870, n53871, n53872, n53873, n53874,
    n53875, n53876, n53877, n53878, n53879, n53880,
    n53881, n53882, n53883, n53884, n53885, n53886,
    n53887, n53888, n53889, n53890, n53891, n53892,
    n53893, n53894, n53895, n53896, n53897, n53898,
    n53899, n53900, n53901, n53902, n53903, n53904,
    n53905, n53906, n53907, n53908, n53909, n53910,
    n53911, n53912, n53913, n53914, n53915, n53916,
    n53917, n53918, n53919, n53920, n53921, n53922,
    n53923, n53924, n53925, n53926, n53927, n53928,
    n53929, n53930, n53931, n53932, n53933, n53934,
    n53935, n53936, n53937, n53938, n53939, n53940,
    n53941, n53942, n53943, n53944, n53945, n53946,
    n53947, n53948, n53949, n53950, n53951, n53952,
    n53953, n53954, n53955, n53956, n53957, n53958,
    n53959, n53960, n53961, n53962, n53963, n53964,
    n53965, n53966, n53967, n53968, n53969, n53970,
    n53971, n53972, n53973, n53974, n53975, n53976,
    n53977, n53978, n53979, n53980, n53981, n53982,
    n53983, n53984, n53985, n53986, n53987, n53988,
    n53989, n53990, n53991, n53992, n53993, n53994,
    n53995, n53996, n53997, n53998, n53999, n54000,
    n54001, n54002, n54003, n54004, n54005, n54006,
    n54007, n54008, n54009, n54010, n54011, n54012,
    n54013, n54014, n54015, n54016, n54017, n54018,
    n54019, n54020, n54021, n54022, n54023, n54024,
    n54025, n54026, n54027, n54028, n54029, n54030,
    n54031, n54032, n54033, n54034, n54035, n54036,
    n54037, n54038, n54039, n54040, n54041, n54042,
    n54043, n54044, n54045, n54046, n54047, n54048,
    n54049, n54050, n54051, n54052, n54053, n54054,
    n54055, n54056, n54057, n54058, n54059, n54060,
    n54061, n54062, n54063, n54064, n54065, n54066,
    n54067, n54068, n54069, n54070, n54071, n54072,
    n54073, n54074, n54075, n54076, n54077, n54078,
    n54079, n54080, n54081, n54082, n54083, n54084,
    n54085, n54086, n54087, n54088, n54089, n54090,
    n54091, n54092, n54093, n54094, n54095, n54096,
    n54097, n54098, n54099, n54100, n54101, n54102,
    n54103, n54104, n54105, n54106, n54107, n54108,
    n54109, n54110, n54111, n54112, n54113, n54114,
    n54115, n54116, n54117, n54118, n54119, n54120,
    n54121, n54122, n54123, n54124, n54125, n54126,
    n54127, n54128, n54129, n54130, n54131, n54132,
    n54133, n54134, n54135, n54136, n54137, n54138,
    n54139, n54140, n54141, n54142, n54143, n54144,
    n54145, n54146, n54147, n54148, n54149, n54150,
    n54151, n54152, n54153, n54154, n54155, n54156,
    n54157, n54158, n54159, n54160, n54161, n54162,
    n54163, n54164, n54165, n54166, n54167, n54168,
    n54169, n54170, n54171, n54172, n54173, n54174,
    n54175, n54176, n54177, n54178, n54179, n54180,
    n54181, n54182, n54183, n54184, n54185, n54186,
    n54187, n54188, n54189, n54190, n54191, n54192,
    n54193, n54194, n54195, n54196, n54197, n54198,
    n54199, n54200, n54201, n54202, n54203, n54204,
    n54205, n54206, n54207, n54208, n54209, n54210,
    n54211, n54212, n54213, n54214, n54215, n54216,
    n54217, n54218, n54219, n54220, n54221, n54222,
    n54223, n54224, n54225, n54226, n54227, n54228,
    n54229, n54230, n54231, n54232, n54233, n54234,
    n54235, n54236, n54237, n54238, n54239, n54240,
    n54241, n54242, n54243, n54244, n54245, n54246,
    n54247, n54248, n54249, n54250, n54251, n54252,
    n54253, n54254, n54255, n54256, n54257, n54258,
    n54259, n54260, n54261, n54262, n54263, n54264,
    n54265, n54266, n54267, n54268, n54269, n54270,
    n54271, n54272, n54273, n54274, n54275, n54276,
    n54277, n54279, n54280, n54281, n54282, n54283,
    n54284, n54285, n54286, n54287, n54288, n54289,
    n54290, n54291, n54292, n54293, n54294, n54295,
    n54296, n54297, n54298, n54299, n54300, n54301,
    n54302, n54303, n54304, n54305, n54306, n54307,
    n54308, n54309, n54310, n54311, n54312, n54313,
    n54314, n54315, n54316, n54317, n54318, n54319,
    n54320, n54321, n54322, n54323, n54324, n54325,
    n54326, n54327, n54328, n54329, n54330, n54331,
    n54332, n54333, n54334, n54335, n54336, n54337,
    n54338, n54339, n54340, n54341, n54342, n54343,
    n54344, n54345, n54346, n54347, n54348, n54349,
    n54350, n54351, n54352, n54353, n54354, n54355,
    n54356, n54357, n54358, n54359, n54360, n54361,
    n54362, n54363, n54364, n54365, n54366, n54367,
    n54368, n54369, n54370, n54371, n54372, n54373,
    n54374, n54375, n54376, n54377, n54378, n54379,
    n54380, n54381, n54382, n54383, n54384, n54385,
    n54386, n54387, n54388, n54389, n54390, n54391,
    n54392, n54393, n54394, n54395, n54396, n54397,
    n54398, n54399, n54400, n54401, n54402, n54403,
    n54404, n54405, n54406, n54407, n54408, n54409,
    n54410, n54411, n54412, n54413, n54414, n54415,
    n54416, n54417, n54418, n54419, n54420, n54421,
    n54422, n54423, n54424, n54425, n54426, n54427,
    n54428, n54429, n54430, n54431, n54432, n54433,
    n54434, n54435, n54436, n54437, n54438, n54439,
    n54440, n54441, n54442, n54443, n54444, n54445,
    n54446, n54447, n54448, n54449, n54450, n54451,
    n54452, n54453, n54454, n54455, n54456, n54457,
    n54458, n54459, n54460, n54461, n54462, n54463,
    n54464, n54465, n54466, n54467, n54468, n54469,
    n54470, n54471, n54472, n54473, n54474, n54475,
    n54476, n54477, n54478, n54479, n54480, n54481,
    n54482, n54483, n54484, n54485, n54486, n54487,
    n54488, n54489, n54490, n54491, n54492, n54493,
    n54494, n54495, n54496, n54497, n54498, n54499,
    n54500, n54501, n54502, n54503, n54504, n54505,
    n54506, n54507, n54508, n54509, n54510, n54511,
    n54512, n54513, n54514, n54515, n54516, n54517,
    n54518, n54519, n54520, n54521, n54522, n54523,
    n54524, n54525, n54526, n54527, n54528, n54529,
    n54530, n54531, n54532, n54533, n54534, n54535,
    n54536, n54537, n54538, n54539, n54540, n54541,
    n54542, n54543, n54544, n54545, n54546, n54547,
    n54548, n54549, n54550, n54551, n54552, n54553,
    n54554, n54555, n54556, n54557, n54558, n54559,
    n54560, n54561, n54562, n54563, n54564, n54565,
    n54566, n54567, n54568, n54569, n54570, n54571,
    n54572, n54573, n54574, n54575, n54576, n54577,
    n54578, n54579, n54580, n54581, n54582, n54583,
    n54584, n54585, n54586, n54587, n54588, n54589,
    n54590, n54591, n54592, n54593, n54594, n54595,
    n54596, n54597, n54598, n54599, n54600, n54601,
    n54602, n54603, n54604, n54605, n54606, n54607,
    n54608, n54609, n54610, n54611, n54612, n54613,
    n54614, n54615, n54616, n54617, n54618, n54619,
    n54620, n54621, n54622, n54623, n54624, n54625,
    n54626, n54627, n54628, n54629, n54630, n54631,
    n54632, n54633, n54634, n54635, n54636, n54637,
    n54638, n54639, n54640, n54641, n54642, n54643,
    n54644, n54645, n54646, n54647, n54648, n54649,
    n54650, n54651, n54652, n54653, n54654, n54655,
    n54656, n54657, n54658, n54659, n54660, n54661,
    n54662, n54663, n54664, n54665, n54666, n54667,
    n54668, n54669, n54670, n54671, n54672, n54673,
    n54674, n54675, n54676, n54677, n54678, n54679,
    n54680, n54681, n54682, n54683, n54684, n54685,
    n54686, n54687, n54688, n54689, n54690, n54691,
    n54692, n54693, n54694, n54695, n54696, n54697,
    n54698, n54699, n54700, n54701, n54702, n54703,
    n54704, n54705, n54706, n54707, n54708, n54709,
    n54710, n54711, n54712, n54713, n54714, n54715,
    n54716, n54717, n54718, n54719, n54720, n54721,
    n54722, n54723, n54724, n54725, n54726, n54727,
    n54728, n54729, n54730, n54731, n54732, n54733,
    n54734, n54735, n54736, n54737, n54738, n54739,
    n54740, n54741, n54742, n54743, n54744, n54745,
    n54746, n54747, n54748, n54749, n54750, n54751,
    n54752, n54753, n54754, n54755, n54756, n54757,
    n54758, n54759, n54761, n54762, n54763, n54764,
    n54765, n54766, n54767, n54768, n54769, n54770,
    n54771, n54772, n54773, n54774, n54775, n54776,
    n54777, n54778, n54779, n54780, n54781, n54782,
    n54783, n54784, n54785, n54786, n54787, n54788,
    n54789, n54790, n54791, n54792, n54793, n54794,
    n54795, n54796, n54797, n54798, n54799, n54800,
    n54801, n54802, n54803, n54804, n54805, n54806,
    n54807, n54808, n54809, n54810, n54811, n54812,
    n54813, n54814, n54815, n54816, n54817, n54818,
    n54819, n54820, n54821, n54822, n54823, n54824,
    n54825, n54826, n54827, n54828, n54829, n54830,
    n54831, n54832, n54833, n54834, n54835, n54836,
    n54837, n54838, n54839, n54840, n54841, n54842,
    n54843, n54844, n54845, n54846, n54847, n54848,
    n54849, n54850, n54851, n54852, n54853, n54854,
    n54855, n54856, n54857, n54858, n54859, n54860,
    n54861, n54862, n54863, n54864, n54865, n54866,
    n54867, n54868, n54869, n54870, n54871, n54872,
    n54873, n54874, n54875, n54876, n54877, n54878,
    n54879, n54880, n54881, n54882, n54883, n54884,
    n54885, n54886, n54887, n54888, n54889, n54890,
    n54891, n54892, n54893, n54894, n54895, n54896,
    n54897, n54898, n54899, n54900, n54901, n54902,
    n54903, n54904, n54905, n54906, n54907, n54908,
    n54909, n54910, n54911, n54912, n54913, n54914,
    n54915, n54916, n54917, n54918, n54919, n54920,
    n54921, n54922, n54923, n54924, n54925, n54926,
    n54927, n54928, n54929, n54930, n54931, n54932,
    n54933, n54934, n54935, n54936, n54937, n54938,
    n54939, n54940, n54941, n54942, n54943, n54944,
    n54945, n54946, n54947, n54948, n54949, n54950,
    n54951, n54952, n54953, n54954, n54955, n54956,
    n54957, n54958, n54959, n54960, n54961, n54962,
    n54963, n54964, n54965, n54966, n54967, n54968,
    n54969, n54970, n54971, n54972, n54973, n54974,
    n54975, n54976, n54977, n54978, n54979, n54980,
    n54981, n54982, n54983, n54984, n54985, n54986,
    n54987, n54988, n54989, n54990, n54991, n54992,
    n54993, n54994, n54995, n54996, n54997, n54998,
    n54999, n55000, n55001, n55002, n55003, n55004,
    n55005, n55006, n55007, n55008, n55009, n55010,
    n55011, n55012, n55013, n55014, n55015, n55016,
    n55017, n55018, n55019, n55020, n55021, n55022,
    n55023, n55024, n55025, n55026, n55027, n55028,
    n55029, n55030, n55031, n55032, n55033, n55034,
    n55035, n55036, n55037, n55038, n55039, n55040,
    n55041, n55042, n55043, n55044, n55045, n55046,
    n55047, n55048, n55049, n55050, n55051, n55052,
    n55053, n55054, n55055, n55056, n55057, n55058,
    n55059, n55060, n55061, n55062, n55063, n55064,
    n55065, n55066, n55067, n55068, n55069, n55070,
    n55071, n55072, n55073, n55074, n55075, n55076,
    n55077, n55078, n55079, n55080, n55081, n55082,
    n55083, n55084, n55085, n55086, n55087, n55088,
    n55089, n55090, n55091, n55092, n55093, n55094,
    n55095, n55096, n55097, n55098, n55099, n55100,
    n55101, n55102, n55103, n55104, n55105, n55106,
    n55107, n55108, n55109, n55110, n55111, n55112,
    n55113, n55114, n55115, n55116, n55117, n55118,
    n55119, n55120, n55121, n55122, n55123, n55124,
    n55125, n55126, n55127, n55128, n55129, n55130,
    n55131, n55132, n55133, n55134, n55135, n55136,
    n55137, n55138, n55139, n55140, n55141, n55142,
    n55143, n55144, n55145, n55146, n55147, n55148,
    n55149, n55150, n55151, n55152, n55153, n55154,
    n55155, n55156, n55157, n55158, n55159, n55160,
    n55161, n55162, n55163, n55164, n55165, n55166,
    n55167, n55168, n55169, n55170, n55171, n55172,
    n55173, n55174, n55175, n55176, n55177, n55178,
    n55179, n55180, n55181, n55182, n55183, n55184,
    n55185, n55186, n55187, n55188, n55189, n55190,
    n55191, n55192, n55193, n55194, n55195, n55196,
    n55197, n55198, n55199, n55200, n55201, n55202,
    n55203, n55204, n55205, n55206, n55207, n55208,
    n55209, n55210, n55211, n55212, n55213, n55214,
    n55215, n55216, n55217, n55218, n55219, n55220,
    n55221, n55222, n55223, n55224, n55225, n55226,
    n55227, n55228, n55229, n55230, n55231, n55232,
    n55233, n55234, n55235, n55236, n55237, n55238,
    n55239, n55240, n55241, n55242, n55243, n55244,
    n55245, n55246, n55247, n55248, n55249, n55250,
    n55251, n55252, n55253, n55254, n55255, n55256,
    n55257, n55258, n55259, n55260, n55261, n55262,
    n55263, n55264, n55265, n55266, n55267, n55268,
    n55269, n55270, n55271, n55272, n55273, n55274,
    n55275, n55276, n55277, n55278, n55279, n55280,
    n55281, n55282, n55283, n55284, n55285, n55286,
    n55287, n55288, n55289, n55290, n55291, n55292,
    n55293, n55294, n55295, n55296, n55297, n55298,
    n55299, n55300, n55301, n55302, n55303, n55304,
    n55305, n55306, n55307, n55308, n55309, n55310,
    n55311, n55312, n55313, n55314, n55315, n55316,
    n55317, n55318, n55319, n55320, n55321, n55322,
    n55323, n55324, n55325, n55326, n55327, n55328,
    n55329, n55330, n55331, n55332, n55333, n55334,
    n55335, n55336, n55337, n55338, n55339, n55340,
    n55341, n55342, n55343, n55344, n55345, n55346,
    n55347, n55348, n55349, n55350, n55351, n55352,
    n55353, n55354, n55355, n55356, n55357, n55358,
    n55359, n55360, n55361, n55362, n55363, n55364,
    n55365, n55366, n55367, n55368, n55369, n55370,
    n55371, n55372, n55373, n55374, n55375, n55376,
    n55377, n55378, n55379, n55380, n55381, n55382,
    n55383, n55384, n55385, n55386, n55387, n55388,
    n55389, n55390, n55391, n55392, n55393, n55394,
    n55395, n55396, n55397, n55398, n55399, n55400,
    n55401, n55402, n55403, n55404, n55405, n55406,
    n55407, n55408, n55409, n55410, n55411, n55412,
    n55413, n55414, n55415, n55416, n55417, n55418,
    n55419, n55420, n55421, n55422, n55423, n55424,
    n55425, n55426, n55427, n55428, n55429, n55430,
    n55431, n55432, n55433, n55434, n55435, n55436,
    n55437, n55438, n55439, n55440, n55441, n55442,
    n55443, n55444, n55445, n55446, n55447, n55448,
    n55449, n55450, n55451, n55452, n55453, n55454,
    n55455, n55456, n55457, n55458, n55459, n55460,
    n55461, n55462, n55463, n55464, n55465, n55466,
    n55467, n55468, n55469, n55470, n55471, n55472,
    n55473, n55474, n55475, n55476, n55477, n55478,
    n55479, n55480, n55481, n55482, n55483, n55484,
    n55485, n55486, n55487, n55488, n55489, n55490,
    n55491, n55492, n55493, n55494, n55495, n55496,
    n55497, n55498, n55499, n55500, n55501, n55502,
    n55503, n55504, n55505, n55506, n55507, n55508,
    n55509, n55510, n55511, n55512, n55513, n55514,
    n55515, n55516, n55517, n55518, n55519, n55520,
    n55521, n55522, n55523, n55524, n55525, n55526,
    n55527, n55528, n55529, n55530, n55531, n55532,
    n55533, n55534, n55535, n55536, n55537, n55538,
    n55539, n55540, n55541, n55542, n55543, n55544,
    n55545, n55546, n55547, n55548, n55549, n55550,
    n55551, n55552, n55553, n55554, n55555, n55556,
    n55557, n55558, n55559, n55560, n55561, n55562,
    n55563, n55564, n55565, n55566, n55567, n55568,
    n55569, n55570, n55571, n55572, n55573, n55574,
    n55575, n55576, n55577, n55578, n55579, n55580,
    n55581, n55582, n55583, n55584, n55585, n55586,
    n55587, n55588, n55589, n55590, n55591, n55592,
    n55593, n55594, n55595, n55596, n55597, n55598,
    n55599, n55600, n55601, n55602, n55603, n55604,
    n55605, n55606, n55607, n55608, n55609, n55610,
    n55611, n55612, n55613, n55614, n55615, n55616,
    n55617, n55618, n55619, n55620, n55621, n55622,
    n55623, n55624, n55625, n55626, n55627, n55628,
    n55629, n55630, n55631, n55632, n55633, n55634,
    n55635, n55636, n55637, n55638, n55639, n55640,
    n55641, n55642, n55643, n55644, n55645, n55646,
    n55647, n55648, n55649, n55650, n55651, n55652,
    n55653, n55654, n55655, n55656, n55657, n55658,
    n55659, n55660, n55661, n55662, n55663, n55664,
    n55665, n55666, n55667, n55668, n55669, n55670,
    n55671, n55672, n55673, n55674, n55675, n55676,
    n55677, n55678, n55679, n55680, n55681, n55682,
    n55683, n55684, n55685, n55686, n55687, n55688,
    n55689, n55690, n55691, n55692, n55693, n55694,
    n55695, n55696, n55697, n55698, n55699, n55700,
    n55701, n55702, n55703, n55704, n55705, n55706,
    n55707, n55708, n55709, n55710, n55711, n55712,
    n55713, n55714, n55715, n55716, n55717, n55718,
    n55719, n55720, n55721, n55722, n55723, n55724,
    n55725, n55726, n55727, n55728, n55729, n55730,
    n55731, n55732, n55733, n55734, n55735, n55736,
    n55737, n55738, n55739, n55740, n55741, n55742,
    n55743, n55744, n55745, n55746, n55747, n55748,
    n55749, n55750, n55751, n55752, n55753, n55754,
    n55755, n55756, n55757, n55758, n55759, n55760,
    n55761, n55762, n55763, n55764, n55765, n55766,
    n55767, n55768, n55769, n55770, n55771, n55772,
    n55773, n55774, n55775, n55776, n55777, n55778,
    n55779, n55780, n55781, n55782, n55783, n55784,
    n55785, n55786, n55787, n55788, n55789, n55791,
    n55792, n55793, n55794, n55795, n55796, n55797,
    n55798, n55799, n55800, n55801, n55802, n55803,
    n55804, n55805, n55806, n55807, n55808, n55809,
    n55810, n55811, n55812, n55813, n55814, n55815,
    n55816, n55817, n55818, n55819, n55820, n55821,
    n55822, n55823, n55824, n55825, n55826, n55827,
    n55828, n55829, n55830, n55831, n55832, n55833,
    n55834, n55835, n55836, n55837, n55838, n55839,
    n55840, n55841, n55842, n55843, n55844, n55845,
    n55846, n55847, n55848, n55849, n55850, n55851,
    n55853, n55854, n55855, n55856, n55857, n55858,
    n55859, n55860, n55861, n55862, n55863, n55864,
    n55865, n55866, n55867, n55868, n55869, n55870,
    n55871, n55872, n55873, n55874, n55875, n55876,
    n55877, n55878, n55879, n55880, n55881, n55882,
    n55883, n55884, n55885, n55886, n55887, n55888,
    n55889, n55890, n55891, n55892, n55893, n55894,
    n55895, n55896, n55897, n55898, n55899, n55900,
    n55901, n55902, n55903, n55904, n55905, n55906,
    n55907, n55908, n55909, n55910, n55911, n55912,
    n55913, n55914, n55915, n55916, n55917, n55918,
    n55919, n55920, n55921, n55922, n55923, n55924,
    n55925, n55926, n55927, n55928, n55929, n55930,
    n55931, n55932, n55933, n55934, n55935, n55936,
    n55937, n55938, n55939, n55940, n55941, n55942,
    n55943, n55944, n55945, n55946, n55947, n55948,
    n55949, n55950, n55951, n55952, n55953, n55954,
    n55955, n55956, n55957, n55958, n55959, n55960,
    n55961, n55962, n55963, n55964, n55965, n55966,
    n55967, n55968, n55969, n55970, n55971, n55972,
    n55973, n55974, n55975, n55976, n55977, n55978,
    n55979, n55980, n55981, n55982, n55983, n55984,
    n55985, n55986, n55987, n55988, n55989, n55990,
    n55991, n55992, n55993, n55994, n55995, n55996,
    n55997, n55998, n55999, n56000, n56001, n56002,
    n56003, n56004, n56005, n56006, n56007, n56008,
    n56009, n56010, n56011, n56012, n56013, n56014,
    n56015, n56016, n56017, n56018, n56019, n56020,
    n56021, n56022, n56023, n56024, n56025, n56026,
    n56027, n56028, n56029, n56030, n56031, n56032,
    n56033, n56034, n56035, n56036, n56037, n56038,
    n56039, n56040, n56041, n56042, n56043, n56044,
    n56045, n56046, n56047, n56048, n56049, n56050,
    n56051, n56052, n56053, n56054, n56055, n56056,
    n56057, n56058, n56059, n56060, n56061, n56062,
    n56063, n56064, n56065, n56066, n56067, n56068,
    n56069, n56070, n56071, n56072, n56073, n56074,
    n56075, n56076, n56077, n56078, n56079, n56080,
    n56081, n56082, n56083, n56084, n56085, n56086,
    n56087, n56088, n56089, n56090, n56091, n56092,
    n56093, n56094, n56095, n56096, n56097, n56098,
    n56099, n56100, n56101, n56102, n56103, n56104,
    n56105, n56106, n56107, n56108, n56109, n56110,
    n56111, n56112, n56113, n56114, n56115, n56116,
    n56117, n56118, n56119, n56120, n56121, n56122,
    n56123, n56124, n56125, n56126, n56127, n56128,
    n56129, n56130, n56131, n56132, n56133, n56134,
    n56135, n56136, n56137, n56138, n56139, n56140,
    n56141, n56142, n56143, n56144, n56145, n56146,
    n56147, n56148, n56149, n56150, n56151, n56152,
    n56153, n56154, n56155, n56156, n56157, n56158,
    n56159, n56160, n56161, n56162, n56163, n56164,
    n56165, n56166, n56167, n56168, n56169, n56170,
    n56171, n56172, n56173, n56174, n56175, n56176,
    n56177, n56178, n56179, n56180, n56181, n56182,
    n56183, n56184, n56185, n56186, n56187, n56188,
    n56189, n56190, n56191, n56192, n56193, n56194,
    n56195, n56196, n56197, n56198, n56199, n56200,
    n56201, n56202, n56203, n56204, n56205, n56206,
    n56207, n56208, n56209, n56210, n56211, n56212,
    n56213, n56214, n56215, n56216, n56217, n56218,
    n56219, n56220, n56221, n56222, n56223, n56224,
    n56225, n56226, n56227, n56228, n56229, n56230,
    n56231, n56232, n56233, n56234, n56235, n56236,
    n56237, n56238, n56239, n56240, n56241, n56242,
    n56243, n56244, n56245, n56246, n56247, n56248,
    n56249, n56250, n56251, n56252, n56253, n56254,
    n56255, n56256, n56257, n56258, n56259, n56260,
    n56261, n56262, n56263, n56264, n56265, n56266,
    n56267, n56268, n56269, n56270, n56271, n56272,
    n56273, n56274, n56275, n56276, n56277, n56278,
    n56279, n56280, n56281, n56282, n56283, n56284,
    n56285, n56286, n56287, n56288, n56289, n56290,
    n56291, n56292, n56293, n56294, n56295, n56296,
    n56297, n56298, n56299, n56300, n56301, n56302,
    n56303, n56304, n56305, n56306, n56307, n56308,
    n56309, n56310, n56311, n56312, n56313, n56314,
    n56315, n56316, n56317, n56318, n56319, n56320,
    n56321, n56322, n56323, n56324, n56325, n56326,
    n56327, n56328, n56329, n56330, n56331, n56332,
    n56333, n56334, n56335, n56336, n56337, n56338,
    n56339, n56340, n56341, n56342, n56343, n56344,
    n56345, n56346, n56347, n56348, n56349, n56350,
    n56351, n56352, n56353, n56354, n56355, n56356,
    n56357, n56358, n56359, n56360, n56361, n56362,
    n56363, n56364, n56365, n56366, n56367, n56368,
    n56369, n56370, n56371, n56372, n56373, n56374,
    n56375, n56376, n56377, n56378, n56379, n56380,
    n56381, n56382, n56383, n56384, n56385, n56386,
    n56387, n56388, n56389, n56390, n56391, n56392,
    n56393, n56394, n56395, n56396, n56397, n56398,
    n56399, n56400, n56401, n56402, n56403, n56404,
    n56405, n56406, n56407, n56408, n56409, n56410,
    n56411, n56412, n56413, n56414, n56415, n56416,
    n56417, n56418, n56419, n56420, n56421, n56422,
    n56423, n56424, n56425, n56426, n56427, n56428,
    n56429, n56430, n56431, n56432, n56433, n56434,
    n56435, n56436, n56437, n56438, n56439, n56440,
    n56441, n56442, n56443, n56444, n56445, n56446,
    n56447, n56448, n56449, n56450, n56451, n56452,
    n56453, n56454, n56455, n56456, n56457, n56458,
    n56459, n56460, n56461, n56462, n56463, n56464,
    n56465, n56466, n56467, n56468, n56469, n56470,
    n56471, n56472, n56473, n56474, n56475, n56476,
    n56477, n56478, n56479, n56480, n56481, n56482,
    n56483, n56484, n56485, n56486, n56487, n56488,
    n56489, n56490, n56491, n56492, n56493, n56494,
    n56495, n56496, n56497, n56498, n56499, n56500,
    n56501, n56502, n56503, n56504, n56505, n56506,
    n56507, n56508, n56509, n56510, n56511, n56512,
    n56513, n56514, n56515, n56516, n56517, n56518,
    n56519, n56520, n56521, n56522, n56523, n56524,
    n56525, n56526, n56527, n56528, n56529, n56530,
    n56531, n56532, n56533, n56534, n56535, n56536,
    n56537, n56538, n56539, n56540, n56541, n56542,
    n56543, n56544, n56545, n56546, n56547, n56548,
    n56549, n56550, n56551, n56552, n56553, n56554,
    n56555, n56556, n56557, n56558, n56559, n56560,
    n56561, n56562, n56563, n56564, n56565, n56566,
    n56567, n56568, n56569, n56570, n56571, n56572,
    n56573, n56574, n56575, n56576, n56577, n56578,
    n56579, n56580, n56581, n56582, n56583, n56584,
    n56585, n56586, n56587, n56588, n56589, n56590,
    n56591, n56592, n56593, n56594, n56595, n56596,
    n56597, n56598, n56599, n56600, n56601, n56602,
    n56603, n56604, n56605, n56606, n56607, n56608,
    n56609, n56610, n56611, n56612, n56613, n56614,
    n56615, n56616, n56617, n56618, n56619, n56620,
    n56621, n56622, n56623, n56624, n56625, n56626,
    n56627, n56628, n56629, n56630, n56631, n56632,
    n56633, n56634, n56635, n56636, n56637, n56638,
    n56639, n56640, n56641, n56642, n56643, n56644,
    n56645, n56646, n56647, n56648, n56649, n56650,
    n56651, n56652, n56653, n56654, n56655, n56656,
    n56657, n56658, n56659, n56660, n56661, n56662,
    n56663, n56664, n56665, n56666, n56667, n56668,
    n56669, n56670, n56671, n56672, n56673, n56674,
    n56675, n56676, n56677, n56678, n56679, n56680,
    n56681, n56682, n56683, n56684, n56685, n56686,
    n56687, n56688, n56689, n56690, n56691, n56692,
    n56693, n56694, n56695, n56696, n56697, n56698,
    n56699, n56700, n56701, n56702, n56703, n56704,
    n56705, n56706, n56707, n56708, n56709, n56710,
    n56711, n56712, n56713, n56714, n56715, n56716,
    n56717, n56718, n56719, n56720, n56721, n56722,
    n56723, n56724, n56725, n56726, n56727, n56728,
    n56729, n56730, n56731, n56732, n56733, n56734,
    n56735, n56736, n56737, n56738, n56739, n56740,
    n56741, n56742, n56743, n56744, n56745, n56746,
    n56747, n56748, n56749, n56750, n56751, n56752,
    n56753, n56754, n56755, n56756, n56757, n56758,
    n56759, n56760, n56761, n56762, n56763, n56764,
    n56765, n56766, n56767, n56768, n56769, n56770,
    n56771, n56772, n56773, n56774, n56775, n56776,
    n56777, n56778, n56779, n56780, n56781, n56782,
    n56783, n56784, n56785, n56786, n56787, n56788,
    n56789, n56790, n56791, n56792, n56793, n56794,
    n56795, n56796, n56797, n56798, n56799, n56800,
    n56801, n56802, n56803, n56804, n56805, n56806,
    n56807, n56808, n56809, n56810, n56811, n56812,
    n56813, n56814, n56815, n56816, n56817, n56818,
    n56819, n56820, n56821, n56822, n56823, n56824,
    n56825, n56826, n56827, n56828, n56829, n56830,
    n56831, n56832, n56833, n56834, n56835, n56836,
    n56837, n56838, n56839, n56840, n56841, n56842,
    n56843, n56844, n56845, n56846, n56847, n56848,
    n56849, n56850, n56851, n56852, n56853, n56854,
    n56855, n56856, n56857, n56858, n56859, n56860,
    n56861, n56862, n56863, n56864, n56865, n56866,
    n56867, n56868, n56869, n56870, n56871, n56872,
    n56873, n56874, n56875, n56876, n56877, n56878,
    n56879, n56880, n56881, n56882, n56883, n56884,
    n56885, n56886, n56887, n56888, n56889, n56890,
    n56891, n56892, n56893, n56894, n56895, n56896,
    n56897, n56898, n56899, n56900, n56901, n56902,
    n56903, n56904, n56905, n56906, n56907, n56908,
    n56909, n56910, n56911, n56912, n56913, n56914,
    n56915, n56916, n56917, n56918, n56919, n56920,
    n56921, n56922, n56923, n56924, n56925, n56926,
    n56927, n56928, n56929, n56930, n56931, n56932,
    n56933, n56934, n56935, n56936, n56937, n56938,
    n56939, n56940, n56941, n56942, n56943, n56944,
    n56945, n56946, n56947, n56948, n56949, n56950,
    n56951, n56952, n56953, n56954, n56955, n56956,
    n56957, n56958, n56959, n56960, n56961, n56962,
    n56963, n56964, n56965, n56966, n56967, n56968,
    n56969, n56970, n56971, n56972, n56973, n56974,
    n56975, n56976, n56977, n56978, n56979, n56980,
    n56981, n56982, n56983, n56984, n56985, n56986,
    n56987, n56988, n56989, n56990, n56991, n56992,
    n56993, n56994, n56995, n56996, n56997, n56998,
    n56999, n57000, n57001, n57002, n57003, n57004,
    n57005, n57006, n57007, n57008, n57009, n57010,
    n57011, n57012, n57013, n57014, n57015, n57016,
    n57017, n57018, n57019, n57020, n57021, n57022,
    n57023, n57024, n57025, n57026, n57027, n57028,
    n57029, n57030, n57031, n57032, n57033, n57034,
    n57035, n57036, n57037, n57038, n57039, n57040,
    n57041, n57042, n57043, n57044, n57045, n57046,
    n57047, n57048, n57049, n57050, n57051, n57052,
    n57053, n57054, n57055, n57056, n57057, n57058,
    n57059, n57060, n57061, n57062, n57063, n57064,
    n57065, n57066, n57067, n57068, n57069, n57070,
    n57071, n57072, n57073, n57074, n57075, n57076,
    n57077, n57078, n57079, n57080, n57081, n57082,
    n57083, n57084, n57085, n57086, n57087, n57088,
    n57089, n57090, n57091, n57092, n57093, n57094,
    n57095, n57096, n57097, n57098, n57099, n57100,
    n57101, n57102, n57103, n57104, n57105, n57106,
    n57107, n57108, n57109, n57110, n57111, n57112,
    n57113, n57114, n57115, n57116, n57117, n57118,
    n57119, n57120, n57121, n57122, n57123, n57124,
    n57125, n57126, n57127, n57128, n57129, n57130,
    n57131, n57132, n57133, n57134, n57135, n57136,
    n57137, n57138, n57139, n57140, n57141, n57142,
    n57143, n57144, n57145, n57146, n57147, n57148,
    n57149, n57150, n57151, n57152, n57153, n57154,
    n57155, n57156, n57157, n57158, n57159, n57160,
    n57161, n57162, n57163, n57164, n57165, n57166,
    n57167, n57168, n57169, n57170, n57171, n57172,
    n57173, n57174, n57175, n57176, n57177, n57178,
    n57179, n57180, n57181, n57182, n57183, n57184,
    n57185, n57186, n57187, n57188, n57189, n57190,
    n57191, n57192, n57193, n57194, n57195, n57196,
    n57197, n57198, n57199, n57200, n57201, n57202,
    n57203, n57204, n57205, n57206, n57207, n57208,
    n57209, n57210, n57211, n57212, n57213, n57214,
    n57215, n57216, n57217, n57218, n57219, n57220,
    n57221, n57222, n57223, n57224, n57225, n57226,
    n57227, n57228, n57229, n57230, n57231, n57232,
    n57233, n57234, n57235, n57236, n57237, n57238,
    n57239, n57240, n57241, n57242, n57243, n57244,
    n57245, n57246, n57247, n57248, n57249, n57250,
    n57251, n57252, n57253, n57254, n57255, n57256,
    n57257, n57258, n57259, n57260, n57261, n57262,
    n57263, n57264, n57265, n57266, n57267, n57268,
    n57269, n57270, n57271, n57272, n57273, n57274,
    n57275, n57276, n57277, n57278, n57279, n57280,
    n57281, n57282, n57283, n57284, n57285, n57286,
    n57287, n57288, n57289, n57290, n57291, n57292,
    n57293, n57294, n57295, n57296, n57297, n57298,
    n57299, n57300, n57301, n57302, n57303, n57304,
    n57305, n57306, n57307, n57308, n57309, n57310,
    n57311, n57312, n57313, n57314, n57315, n57316,
    n57317, n57318, n57319, n57320, n57321, n57322,
    n57323, n57324, n57325, n57326, n57327, n57328,
    n57329, n57330, n57331, n57332, n57333, n57334,
    n57335, n57336, n57337, n57338, n57339, n57340,
    n57341, n57342, n57343, n57344, n57345, n57346,
    n57347, n57348, n57349, n57350, n57351, n57352,
    n57353, n57354, n57355, n57356, n57357, n57358,
    n57359, n57360, n57361, n57362, n57363, n57364,
    n57365, n57366, n57367, n57368, n57369, n57370,
    n57371, n57372, n57373, n57374, n57375, n57376,
    n57377, n57378, n57379, n57380, n57381, n57382,
    n57383, n57384, n57385, n57386, n57387, n57388,
    n57389, n57390, n57391, n57392, n57393, n57394,
    n57395, n57396, n57397, n57398, n57399, n57400,
    n57401, n57402, n57403, n57404, n57405, n57406,
    n57407, n57408, n57409, n57410, n57411, n57412,
    n57413, n57414, n57415, n57416, n57417, n57418,
    n57419, n57420, n57421, n57422, n57423, n57424,
    n57425, n57426, n57427, n57428, n57429, n57430,
    n57431, n57432, n57433, n57434, n57435, n57437,
    n57438, n57439, n57440, n57441, n57442, n57443,
    n57444, n57445, n57446, n57447, n57448, n57449,
    n57450, n57451, n57452, n57453, n57454, n57455,
    n57456, n57457, n57458, n57459, n57460, n57461,
    n57462, n57463, n57464, n57465, n57466, n57467,
    n57468, n57469, n57470, n57471, n57472, n57473,
    n57474, n57475, n57476, n57477, n57478, n57479,
    n57480, n57481, n57482, n57483, n57484, n57485,
    n57486, n57487, n57488, n57489, n57490, n57491,
    n57492, n57493, n57494, n57495, n57496, n57497,
    n57498, n57499, n57500, n57501, n57502, n57503,
    n57504, n57505, n57506, n57507, n57508, n57509,
    n57510, n57511, n57512, n57513, n57514, n57515,
    n57516, n57517, n57518, n57519, n57520, n57521,
    n57522, n57523, n57524, n57525, n57526, n57527,
    n57528, n57529, n57530, n57531, n57532, n57533,
    n57534, n57535, n57536, n57537, n57538, n57539,
    n57540, n57541, n57542, n57543, n57544, n57545,
    n57546, n57547, n57548, n57549, n57550, n57551,
    n57552, n57553, n57554, n57555, n57556, n57557,
    n57558, n57559, n57560, n57561, n57562, n57563,
    n57564, n57565, n57566, n57567, n57568, n57569,
    n57570, n57571, n57572, n57573, n57574, n57575,
    n57576, n57577, n57578, n57579, n57580, n57581,
    n57582, n57583, n57584, n57585, n57586, n57587,
    n57588, n57589, n57590, n57591, n57592, n57593,
    n57594, n57595, n57596, n57597, n57598, n57599,
    n57600, n57601, n57602, n57603, n57604, n57605,
    n57606, n57607, n57608, n57609, n57610, n57611,
    n57612, n57613, n57614, n57615, n57616, n57617,
    n57619, n57620, n57621, n57622, n57623, n57624,
    n57625, n57626, n57627, n57628, n57629, n57630,
    n57631, n57632, n57633, n57634, n57635, n57636,
    n57637, n57638, n57639, n57640, n57641, n57642,
    n57643, n57644, n57645, n57646, n57647, n57648,
    n57649, n57650, n57651, n57652, n57653, n57654,
    n57655, n57656, n57657, n57658, n57659, n57660,
    n57661, n57662, n57663, n57664, n57665, n57666,
    n57667, n57668, n57670, n57671, n57672, n57673,
    n57674, n57675, n57676, n57677, n57678, n57679,
    n57680, n57681, n57682, n57683, n57684, n57685,
    n57686, n57687, n57688, n57689, n57690, n57691,
    n57692, n57693, n57694, n57695, n57696, n57697,
    n57698, n57699, n57700, n57701, n57702, n57703,
    n57704, n57705, n57706, n57707, n57708, n57709,
    n57710, n57711, n57712, n57713, n57714, n57715,
    n57716, n57717, n57718, n57719, n57720, n57721,
    n57722, n57723, n57724, n57725, n57726, n57727,
    n57728, n57729, n57730, n57731, n57732, n57733,
    n57734, n57735, n57736, n57737, n57738, n57739,
    n57740, n57741, n57742, n57743, n57744, n57745,
    n57746, n57747, n57748, n57749, n57750, n57751,
    n57752, n57753, n57754, n57755, n57756, n57757,
    n57758, n57759, n57760, n57761, n57762, n57763,
    n57764, n57765, n57766, n57767, n57768, n57769,
    n57770, n57771, n57772, n57773, n57774, n57775,
    n57776, n57777, n57778, n57779, n57780, n57781,
    n57782, n57783, n57785, n57786, n57787, n57788,
    n57789, n57790, n57791, n57792, n57793, n57794,
    n57795, n57796, n57797, n57798, n57799, n57800,
    n57801, n57802, n57803, n57804, n57805, n57806,
    n57807, n57808, n57809, n57810, n57811, n57812,
    n57813, n57814, n57815, n57816, n57817, n57818,
    n57819, n57820, n57821, n57822, n57823, n57824,
    n57825, n57826, n57827, n57828, n57829, n57830,
    n57831, n57832, n57833, n57834, n57835, n57836,
    n57837, n57838, n57839, n57840, n57841, n57842,
    n57843, n57844, n57845, n57846, n57847, n57848,
    n57849, n57850, n57851, n57852, n57853, n57854,
    n57855, n57856, n57857, n57858, n57859, n57860,
    n57861, n57862, n57863, n57864, n57865, n57866,
    n57867, n57868, n57869, n57870, n57871, n57872,
    n57873, n57874, n57875, n57876, n57877, n57878,
    n57879, n57880, n57881, n57882, n57883, n57884,
    n57885, n57886, n57887, n57888, n57889, n57890,
    n57891, n57892, n57893, n57894, n57895, n57896,
    n57897, n57898, n57899, n57900, n57901, n57902,
    n57903, n57904, n57905, n57906, n57907, n57908,
    n57909, n57910, n57911, n57912, n57913, n57914,
    n57915, n57916, n57917, n57918, n57919, n57920,
    n57921, n57922, n57923, n57924, n57925, n57926,
    n57927, n57928, n57929, n57930, n57931, n57932,
    n57933, n57934, n57935, n57936, n57937, n57938,
    n57939, n57940, n57941, n57942, n57943, n57944,
    n57945, n57946, n57947, n57948, n57949, n57951,
    n57952, n57953, n57954, n57955, n57956, n57957,
    n57958, n57959, n57960, n57961, n57962, n57963,
    n57964, n57965, n57966, n57967, n57968, n57969,
    n57970, n57971, n57972, n57973, n57974, n57975,
    n57976, n57977, n57978, n57979, n57980, n57981,
    n57982, n57983, n57984, n57985, n57986, n57987,
    n57988, n57989, n57990, n57991, n57992, n57993,
    n57994, n57995, n57996, n57997, n57998, n57999,
    n58000, n58001, n58002, n58003, n58004, n58005,
    n58006, n58007, n58008, n58009, n58010, n58011,
    n58012, n58013, n58014, n58015, n58016, n58018,
    n58019, n58020, n58021, n58022, n58023, n58024,
    n58025, n58026, n58027, n58028, n58029, n58030,
    n58031, n58032, n58033, n58034, n58035, n58036,
    n58037, n58038, n58039, n58040, n58041, n58042,
    n58043, n58044, n58045, n58046, n58047, n58048,
    n58049, n58050, n58051, n58052, n58053, n58054,
    n58055, n58056, n58057, n58058, n58059, n58060,
    n58061, n58062, n58063, n58064, n58065, n58066,
    n58067, n58068, n58069, n58070, n58071, n58072,
    n58073, n58074, n58075, n58076, n58077, n58078,
    n58079, n58080, n58081, n58082, n58083, n58084,
    n58085, n58086, n58087, n58088, n58089, n58090,
    n58091, n58092, n58093, n58094, n58095, n58096,
    n58097, n58098, n58099, n58100, n58101, n58102,
    n58103, n58104, n58105, n58106, n58107, n58108,
    n58109, n58110, n58111, n58112, n58113, n58114,
    n58115, n58116, n58117, n58118, n58119, n58120,
    n58121, n58122, n58124, n58125, n58126, n58127,
    n58128, n58129, n58130, n58131, n58132, n58133,
    n58134, n58135, n58136, n58137, n58138, n58139,
    n58140, n58141, n58142, n58143, n58144, n58145,
    n58146, n58147, n58148, n58149, n58150, n58151,
    n58152, n58153, n58154, n58155, n58156, n58157,
    n58158, n58159, n58160, n58161, n58162, n58163,
    n58164, n58165, n58167, n58168, n58169, n58170,
    n58171, n58172, n58173, n58174, n58175, n58176,
    n58177, n58178, n58179, n58180, n58181, n58182,
    n58183, n58184, n58185, n58186, n58187, n58188,
    n58189, n58190, n58191, n58192, n58193, n58194,
    n58195, n58196, n58197, n58198, n58199, n58200,
    n58201, n58202, n58203, n58204, n58205, n58206,
    n58207, n58208, n58209, n58210, n58211, n58212,
    n58213, n58214, n58215, n58216, n58217, n58218,
    n58219, n58220, n58221, n58222, n58223, n58224,
    n58225, n58226, n58227, n58228, n58229, n58230,
    n58231, n58232, n58233, n58234, n58235, n58236,
    n58237, n58238, n58239, n58240, n58241, n58242,
    n58243, n58244, n58245, n58246, n58247, n58248,
    n58249, n58250, n58251, n58252, n58253, n58254,
    n58255, n58256, n58257, n58258, n58259, n58260,
    n58261, n58262, n58263, n58264, n58265, n58266,
    n58267, n58268, n58269, n58270, n58271, n58272,
    n58273, n58274, n58275, n58276, n58277, n58278,
    n58279, n58280, n58281, n58282, n58283, n58284,
    n58285, n58286, n58287, n58288, n58289, n58290,
    n58291, n58292, n58293, n58294, n58295, n58296,
    n58297, n58298, n58299, n58300, n58301, n58302,
    n58303, n58304, n58305, n58306, n58307, n58308,
    n58309, n58310, n58311, n58312, n58313, n58314,
    n58315, n58316, n58317, n58318, n58319, n58320,
    n58321, n58322, n58323, n58324, n58325, n58326,
    n58327, n58328, n58329, n58330, n58331, n58332,
    n58333, n58334, n58335, n58336, n58337, n58338,
    n58339, n58340, n58341, n58342, n58343, n58344,
    n58345, n58346, n58347, n58348, n58349, n58350,
    n58351, n58352, n58353, n58354, n58355, n58356,
    n58357, n58358, n58359, n58360, n58361, n58362,
    n58363, n58364, n58365, n58366, n58367, n58368,
    n58369, n58370, n58371, n58372, n58373, n58374,
    n58375, n58376, n58377, n58378, n58379, n58380,
    n58381, n58382, n58383, n58384, n58385, n58386,
    n58387, n58388, n58389, n58390, n58391, n58392,
    n58393, n58394, n58395, n58396, n58397, n58398,
    n58399, n58400, n58401, n58402, n58403, n58404,
    n58405, n58406, n58407, n58408, n58409, n58410,
    n58411, n58412, n58413, n58414, n58415, n58416,
    n58417, n58418, n58419, n58420, n58422, n58423,
    n58424, n58425, n58426, n58427, n58428, n58429,
    n58430, n58431, n58432, n58433, n58434, n58435,
    n58436, n58437, n58438, n58439, n58440, n58441,
    n58442, n58443, n58444, n58445, n58446, n58447,
    n58448, n58449, n58450, n58451, n58452, n58453,
    n58454, n58455, n58456, n58457, n58458, n58459,
    n58460, n58461, n58462, n58463, n58465, n58466,
    n58467, n58468, n58469, n58470, n58471, n58472,
    n58473, n58474, n58475, n58476, n58477, n58478,
    n58479, n58480, n58481, n58482, n58483, n58484,
    n58485, n58486, n58487, n58488, n58489, n58490,
    n58491, n58492, n58493, n58494, n58495, n58496,
    n58497, n58498, n58499, n58500, n58501, n58502,
    n58503, n58504, n58505, n58506, n58507, n58508,
    n58509, n58510, n58511, n58513, n58514, n58516,
    n58518, n58519, n58520, n58521, n58522, n58523,
    n58524, n58525, n58526, n58527, n58528, n58529,
    n58530, n58531, n58532, n58533, n58534, n58535,
    n58536, n58537, n58538, n58539, n58540, n58542,
    n58543, n58544, n58545, n58546, n58547, n58548,
    n58549, n58550, n58551, n58552, n58553, n58554,
    n58555, n58556, n58557, n58558, n58560, n58561,
    n58562, n58563, n58564, n58565, n58566, n58567,
    n58569, n58570, n58571, n58572, n58573, n58574,
    n58575, n58576, n58577, n58578, n58579, n58580,
    n58581, n58582, n58583, n58584, n58585, n58586,
    n58587, n58588, n58589, n58590, n58591, n58592,
    n58593, n58594, n58595, n58596, n58597, n58598,
    n58599, n58600, n58601, n58602, n58603, n58604,
    n58605, n58606, n58607, n58608, n58609, n58610,
    n58611, n58612, n58613, n58614, n58615, n58616,
    n58617, n58618, n58619, n58620, n58621, n58622,
    n58623, n58624, n58625, n58626, n58627, n58628,
    n58629, n58630, n58631, n58632, n58633, n58634,
    n58635, n58636, n58637, n58638, n58639, n58640,
    n58641, n58642, n58643, n58644, n58645, n58646,
    n58647, n58649, n58650, n58651, n58652, n58653,
    n58654, n58655, n58656, n58657, n58658, n58659,
    n58660, n58661, n58662, n58663, n58664, n58665,
    n58666, n58667, n58669, n58670, n58671, n58672,
    n58673, n58674, n58675, n58676, n58677, n58678,
    n58679, n58680, n58681, n58682, n58683, n58684,
    n58685, n58686, n58687, n58688, n58689, n58690,
    n58691, n58692, n58693, n58694, n58695, n58696,
    n58697, n58698, n58699, n58700, n58701, n58702,
    n58703, n58704, n58705, n58706, n58707, n58708,
    n58709, n58710, n58711, n58712, n58713, n58714,
    n58715, n58716, n58717, n58718, n58719, n58720,
    n58721, n58722, n58723, n58724, n58725, n58726,
    n58727, n58728, n58729, n58730, n58731, n58732,
    n58733, n58734, n58735, n58736, n58737, n58738,
    n58739, n58740, n58741, n58742, n58743, n58744,
    n58745, n58746, n58747, n58748, n58749, n58750,
    n58751, n58752, n58753, n58754, n58755, n58756,
    n58758, n58760, n58762, n58763, n58764, n58766,
    n58768, n58770, n58772, n58774, n58776, n58778,
    n58779, n58780, n58781, n58782, n58783, n58784,
    n58785, n58786, n58787, n58788, n58789, n58790,
    n58791, n58792, n58793, n58794, n58795, n58796,
    n58797, n58798, n58799, n58800, n58801, n58802,
    n58803, n58804, n58805, n58806, n58807, n58808,
    n58809, n58810, n58811, n58812, n58813, n58814,
    n58815, n58816, n58817, n58818, n58819, n58820,
    n58821, n58822, n58823, n58824, n58825, n58826,
    n58827, n58828, n58829, n58830, n58831, n58832,
    n58833, n58834, n58835, n58836, n58837, n58838,
    n58839, n58840, n58841, n58842, n58843, n58844,
    n58845, n58846, n58847, n58848, n58849, n58850,
    n58851, n58852, n58853, n58854, n58855, n58856,
    n58857, n58858, n58859, n58860, n58861, n58862,
    n58863, n58864, n58865, n58866, n58867, n58868,
    n58869, n58870, n58871, n58872, n58873, n58874,
    n58875, n58876, n58877, n58878, n58879, n58880,
    n58881, n58882, n58883, n58884, n58885, n58886,
    n58887, n58888, n58889, n58890, n58891, n58892,
    n58893, n58894, n58895, n58896, n58897, n58898,
    n58899, n58900, n58901, n58902, n58903, n58904,
    n58905, n58906, n58907, n58909, n58910, n58911,
    n58912, n58913, n58914, n58915, n58916, n58917,
    n58918, n58919, n58920, n58921, n58922, n58923,
    n58924, n58925, n58926, n58927, n58928, n58929,
    n58930, n58931, n58932, n58933, n58934, n58935,
    n58936, n58937, n58938, n58939, n58940, n58941,
    n58942, n58943, n58944, n58945, n58946, n58947,
    n58948, n58949, n58950, n58951, n58952, n58953,
    n58954, n58955, n58956, n58957, n58958, n58959,
    n58960, n58961, n58962, n58963, n58964, n58965,
    n58966, n58967, n58968, n58969, n58970, n58971,
    n58972, n58973, n58974, n58975, n58976, n58977,
    n58978, n58979, n58980, n58981, n58982, n58983,
    n58984, n58985, n58986, n58987, n58988, n58989,
    n58990, n58991, n58992, n58993, n58994, n58995,
    n58996, n58997, n58998, n58999, n59000, n59001,
    n59002, n59003, n59004, n59005, n59006, n59007,
    n59008, n59009, n59010, n59011, n59012, n59013,
    n59014, n59015, n59016, n59017, n59018, n59019,
    n59020, n59021, n59022, n59023, n59024, n59025,
    n59026, n59027, n59028, n59029, n59030, n59031,
    n59032, n59033, n59034, n59035, n59036, n59037,
    n59038, n59039, n59040, n59041, n59042, n59043,
    n59044, n59045, n59046, n59047, n59048, n59049,
    n59050, n59051, n59052, n59053, n59054, n59055,
    n59056, n59057, n59058, n59059, n59060, n59061,
    n59062, n59063, n59064, n59066, n59067, n59068,
    n59069, n59070, n59071, n59072, n59073, n59074,
    n59075, n59076, n59077, n59079, n59080, n59081,
    n59082, n59083, n59084, n59085, n59086, n59087,
    n59088, n59089, n59090, n59092, n59093, n59094,
    n59095, n59096, n59097, n59098, n59099, n59100,
    n59101, n59102, n59103, n59104, n59105, n59106,
    n59107, n59108, n59109, n59110, n59111, n59112,
    n59113, n59114, n59115, n59116, n59117, n59118,
    n59119, n59120, n59121, n59122, n59123, n59124,
    n59125, n59126, n59127, n59128, n59129, n59130,
    n59131, n59132, n59133, n59134, n59135, n59136,
    n59137, n59138, n59139, n59140, n59141, n59142,
    n59143, n59144, n59145, n59146, n59147, n59148,
    n59149, n59150, n59151, n59152, n59153, n59154,
    n59155, n59156, n59157, n59158, n59159, n59160,
    n59161, n59162, n59163, n59164, n59165, n59166,
    n59167, n59168, n59169, n59170, n59171, n59172,
    n59173, n59174, n59175, n59176, n59177, n59178,
    n59179, n59180, n59181, n59182, n59183, n59184,
    n59185, n59186, n59187, n59188, n59189, n59190,
    n59191, n59192, n59193, n59194, n59195, n59196,
    n59197, n59198, n59199, n59200, n59201, n59202,
    n59203, n59204, n59205, n59206, n59207, n59208,
    n59209, n59210, n59211, n59212, n59213, n59214,
    n59215, n59216, n59217, n59218, n59219, n59220,
    n59221, n59222, n59223, n59224, n59225, n59226,
    n59227, n59228, n59229, n59230, n59231, n59232,
    n59233, n59234, n59235, n59236, n59237, n59238,
    n59239, n59240, n59241, n59242, n59243, n59244,
    n59245, n59246, n59247, n59248, n59249, n59250,
    n59251, n59252, n59253, n59254, n59255, n59256,
    n59257, n59258, n59259, n59260, n59261, n59262,
    n59263, n59264, n59265, n59266, n59267, n59268,
    n59269, n59270, n59271, n59272, n59273, n59274,
    n59275, n59276, n59277, n59278, n59279, n59280,
    n59281, n59282, n59283, n59284, n59285, n59286,
    n59287, n59288, n59289, n59290, n59291, n59292,
    n59293, n59294, n59295, n59296, n59297, n59298,
    n59299, n59300, n59301, n59302, n59303, n59304,
    n59305, n59306, n59307, n59308, n59309, n59310,
    n59311, n59312, n59313, n59314, n59315, n59316,
    n59317, n59318, n59319, n59320, n59321, n59322,
    n59323, n59324, n59325, n59326, n59327, n59328,
    n59329, n59330, n59331, n59332, n59333, n59334,
    n59335, n59336, n59337, n59338, n59339, n59340,
    n59341, n59342, n59343, n59344, n59345, n59346,
    n59347, n59348, n59349, n59350, n59351, n59352,
    n59353, n59354, n59355, n59356, n59357, n59358,
    n59359, n59360, n59361, n59362, n59363, n59364,
    n59365, n59366, n59367, n59368, n59369, n59370,
    n59371, n59372, n59373, n59374, n59375, n59376,
    n59377, n59378, n59379, n59380, n59381, n59382,
    n59383, n59384, n59385, n59386, n59387, n59388,
    n59389, n59390, n59391, n59392, n59393, n59394,
    n59395, n59396, n59397, n59398, n59399, n59400,
    n59401, n59402, n59403, n59404, n59405, n59406,
    n59407, n59408, n59409, n59410, n59411, n59412,
    n59413, n59414, n59415, n59416, n59417, n59418,
    n59419, n59420, n59421, n59422, n59423, n59424,
    n59425, n59426, n59427, n59428, n59429, n59430,
    n59431, n59432, n59433, n59434, n59435, n59436,
    n59437, n59438, n59439, n59440, n59441, n59442,
    n59443, n59444, n59445, n59446, n59447, n59448,
    n59449, n59450, n59451, n59452, n59453, n59454,
    n59455, n59456, n59457, n59458, n59459, n59460,
    n59461, n59462, n59463, n59464, n59465, n59466,
    n59467, n59468, n59469, n59470, n59471, n59472,
    n59473, n59474, n59475, n59476, n59477, n59478,
    n59479, n59480, n59481, n59482, n59483, n59484,
    n59485, n59486, n59487, n59488, n59489, n59490,
    n59491, n59492, n59493, n59494, n59495, n59496,
    n59497, n59498, n59499, n59500, n59501, n59502,
    n59503, n59504, n59505, n59506, n59507, n59508,
    n59509, n59510, n59511, n59512, n59513, n59514,
    n59515, n59516, n59517, n59518, n59519, n59520,
    n59521, n59522, n59523, n59524, n59525, n59526,
    n59527, n59528, n59529, n59530, n59531, n59532,
    n59533, n59534, n59535, n59536, n59537, n59538,
    n59539, n59540, n59541, n59542, n59543, n59544,
    n59545, n59546, n59547, n59548, n59549, n59550,
    n59551, n59552, n59553, n59554, n59555, n59556,
    n59557, n59558, n59559, n59560, n59561, n59562,
    n59563, n59564, n59565, n59566, n59567, n59568,
    n59569, n59570, n59571, n59572, n59573, n59574,
    n59575, n59576, n59577, n59578, n59579, n59580,
    n59581, n59582, n59583, n59584, n59585, n59586,
    n59587, n59588, n59589, n59590, n59591, n59592,
    n59593, n59594, n59595, n59596, n59597, n59598,
    n59599, n59600, n59601, n59602, n59603, n59604,
    n59605, n59606, n59607, n59608, n59609, n59610,
    n59611, n59612, n59613, n59614, n59615, n59616,
    n59617, n59618, n59619, n59620, n59621, n59622,
    n59623, n59624, n59625, n59626, n59627, n59628,
    n59629, n59630, n59631, n59632, n59633, n59634,
    n59635, n59636, n59637, n59638, n59639, n59640,
    n59641, n59642, n59643, n59644, n59645, n59646,
    n59647, n59648, n59649, n59650, n59651, n59652,
    n59653, n59654, n59655, n59656, n59657, n59658,
    n59659, n59660, n59661, n59662, n59663, n59664,
    n59665, n59666, n59667, n59668, n59669, n59670,
    n59671, n59672, n59673, n59674, n59675, n59676,
    n59677, n59678, n59679, n59680, n59681, n59682,
    n59683, n59684, n59685, n59686, n59687, n59688,
    n59689, n59690, n59691, n59692, n59693, n59694,
    n59695, n59696, n59697, n59698, n59699, n59700,
    n59701, n59702, n59703, n59704, n59705, n59706,
    n59707, n59708, n59709, n59710, n59711, n59712,
    n59713, n59714, n59715, n59716, n59717, n59718,
    n59719, n59720, n59721, n59722, n59723, n59724,
    n59725, n59726, n59727, n59728, n59729, n59730,
    n59731, n59732, n59733, n59734, n59735, n59736,
    n59737, n59738, n59739, n59740, n59741, n59742,
    n59743, n59744, n59745, n59746, n59747, n59748,
    n59749, n59750, n59751, n59752, n59753, n59754,
    n59755, n59756, n59757, n59758, n59759, n59760,
    n59761, n59762, n59763, n59764, n59765, n59766,
    n59767, n59768, n59769, n59770, n59771, n59772,
    n59773, n59774, n59775, n59776, n59777, n59778,
    n59779, n59780, n59781, n59782, n59783, n59784,
    n59785, n59786, n59787, n59788, n59789, n59790,
    n59791, n59792, n59793, n59794, n59795, n59796,
    n59797, n59798, n59799, n59800, n59801, n59802,
    n59803, n59804, n59805, n59806, n59807, n59808,
    n59809, n59810, n59811, n59812, n59813, n59814,
    n59815, n59816, n59817, n59818, n59819, n59820,
    n59821, n59822, n59823, n59824, n59825, n59826,
    n59827, n59828, n59829, n59830, n59831, n59832,
    n59833, n59834, n59835, n59836, n59837, n59838,
    n59839, n59840, n59841, n59842, n59843, n59844,
    n59845, n59846, n59847, n59848, n59849, n59850,
    n59851, n59852, n59853, n59854, n59855, n59856,
    n59857, n59858, n59859, n59860, n59861, n59862,
    n59863, n59864, n59865, n59866, n59867, n59868,
    n59869, n59870, n59871, n59872, n59873, n59874,
    n59875, n59876, n59877, n59878, n59879, n59880,
    n59881, n59882, n59883, n59884, n59885, n59886,
    n59887, n59888, n59889, n59890, n59891, n59892,
    n59893, n59894, n59895, n59896, n59897, n59898,
    n59899, n59900, n59901, n59902, n59903, n59904,
    n59905, n59906, n59907, n59908, n59909, n59910,
    n59911, n59912, n59913, n59914, n59915, n59916,
    n59917, n59918, n59919, n59920, n59921, n59922,
    n59923, n59924, n59925, n59926, n59927, n59928,
    n59929, n59930, n59931, n59932, n59933, n59934,
    n59935, n59936, n59937, n59938, n59939, n59940,
    n59941, n59942, n59943, n59944, n59945, n59946,
    n59947, n59948, n59949, n59950, n59951, n59952,
    n59953, n59954, n59955, n59956, n59957, n59958,
    n59959, n59960, n59961, n59962, n59963, n59964,
    n59965, n59966, n59967, n59968, n59969, n59970,
    n59971, n59972, n59973, n59974, n59975, n59976,
    n59977, n59978, n59979, n59980, n59981, n59982,
    n59983, n59984, n59985, n59986, n59987, n59988,
    n59989, n59990, n59991, n59992, n59993, n59994,
    n59995, n59996, n59997, n59998, n59999, n60000,
    n60001, n60002, n60003, n60004, n60005, n60006,
    n60007, n60008, n60009, n60010, n60011, n60012,
    n60013, n60014, n60015, n60016, n60017, n60018,
    n60019, n60020, n60021, n60022, n60023, n60024,
    n60025, n60026, n60027, n60028, n60029, n60030,
    n60031, n60032, n60033, n60034, n60035, n60036,
    n60037, n60038, n60039, n60040, n60041, n60042,
    n60043, n60044, n60045, n60046, n60047, n60048,
    n60049, n60050, n60051, n60052, n60053, n60054,
    n60055, n60056, n60057, n60058, n60059, n60060,
    n60061, n60062, n60063, n60064, n60065, n60066,
    n60067, n60068, n60069, n60070, n60071, n60072,
    n60073, n60074, n60075, n60076, n60077, n60078,
    n60079, n60080, n60081, n60082, n60083, n60084,
    n60085, n60086, n60087, n60088, n60089, n60090,
    n60091, n60092, n60093, n60094, n60095, n60096,
    n60097, n60098, n60099, n60100, n60101, n60102,
    n60103, n60104, n60105, n60106, n60107, n60108,
    n60109, n60110, n60111, n60112, n60113, n60114,
    n60115, n60116, n60117, n60118, n60119, n60120,
    n60121, n60122, n60123, n60124, n60125, n60126,
    n60127, n60128, n60129, n60130, n60131, n60132,
    n60133, n60134, n60135, n60136, n60137, n60138,
    n60139, n60140, n60141, n60142, n60143, n60144,
    n60145, n60146, n60147, n60148, n60149, n60150,
    n60151, n60152, n60153, n60154, n60155, n60156,
    n60157, n60158, n60159, n60160, n60161, n60162,
    n60163, n60164, n60165, n60166, n60167, n60168,
    n60169, n60170, n60171, n60172, n60173, n60174,
    n60175, n60176, n60177, n60178, n60179, n60180,
    n60181, n60182, n60183, n60184, n60185, n60186,
    n60187, n60188, n60189, n60190, n60192, n60193,
    n60195, n60196, n60197, n60198, n60199, n60200,
    n60201, n60202, n60203, n60204, n60205, n60206,
    n60207, n60208, n60209, n60210, n60211, n60212,
    n60213, n60214, n60215, n60216, n60217, n60218,
    n60219, n60220, n60221, n60222, n60223, n60224,
    n60225, n60226, n60227, n60228, n60229, n60230,
    n60231, n60232, n60233, n60234, n60235, n60236,
    n60237, n60238, n60239, n60240, n60241, n60242,
    n60243, n60244, n60245, n60246, n60248, n60249,
    n60250, n60251, n60252, n60253, n60254, n60255,
    n60256, n60257, n60258, n60259, n60260, n60261,
    n60262, n60263, n60264, n60265, n60266, n60267,
    n60268, n60269, n60270, n60271, n60272, n60273,
    n60274, n60275, n60276, n60277, n60278, n60279,
    n60280, n60281, n60282, n60283, n60284, n60285,
    n60286, n60287, n60288, n60289, n60290, n60291,
    n60292, n60293, n60294, n60295, n60296, n60297,
    n60298, n60299, n60300, n60301, n60302, n60303,
    n60304, n60305, n60307, n60308, n60309, n60310,
    n60311, n60312, n60313, n60314, n60315, n60316,
    n60317, n60318, n60319, n60320, n60321, n60322,
    n60323, n60324, n60325, n60326, n60327, n60328,
    n60329, n60330, n60331, n60332, n60333, n60334,
    n60335, n60336, n60337, n60338, n60339, n60340,
    n60341, n60342, n60343, n60344, n60345, n60346,
    n60347, n60348, n60349, n60350, n60351, n60352,
    n60353, n60354, n60355, n60356, n60357, n60358,
    n60359, n60360, n60361, n60362, n60363, n60364,
    n60365, n60366, n60367, n60368, n60369, n60370,
    n60371, n60372, n60373, n60374, n60376, n60377,
    n60378, n60379, n60380, n60381, n60382, n60383,
    n60384, n60385, n60386, n60387, n60388, n60389,
    n60390, n60391, n60392, n60393, n60394, n60395,
    n60396, n60397, n60398, n60399, n60400, n60401,
    n60402, n60403, n60404, n60405, n60406, n60407,
    n60408, n60409, n60410, n60411, n60412, n60413,
    n60414, n60415, n60416, n60417, n60418, n60419,
    n60420, n60421, n60422, n60423, n60424, n60425,
    n60426, n60427, n60428, n60429, n60430, n60431,
    n60432, n60433, n60434, n60435, n60436, n60437,
    n60438, n60439, n60440, n60441, n60442, n60443,
    n60444, n60445, n60446, n60447, n60448, n60449,
    n60450, n60451, n60452, n60453, n60454, n60455,
    n60456, n60457, n60458, n60459, n60460, n60461,
    n60462, n60463, n60464, n60465, n60466, n60467,
    n60468, n60469, n60470, n60471, n60472, n60473,
    n60474, n60475, n60476, n60477, n60478, n60479,
    n60480, n60481, n60482, n60483, n60484, n60485,
    n60486, n60487, n60488, n60489, n60490, n60491,
    n60492, n60493, n60494, n60495, n60496, n60497,
    n60498, n60499, n60500, n60501, n60502, n60503,
    n60504, n60505, n60506, n60507, n60508, n60509,
    n60510, n60511, n60512, n60513, n60514, n60515,
    n60516, n60517, n60518, n60519, n60520, n60521,
    n60522, n60523, n60524, n60525, n60526, n60527,
    n60528, n60529, n60530, n60531, n60532, n60533,
    n60534, n60535, n60536, n60537, n60538, n60539,
    n60540, n60541, n60542, n60543, n60544, n60545,
    n60546, n60547, n60548, n60549, n60550, n60551,
    n60552, n60553, n60554, n60555, n60556, n60557,
    n60558, n60559, n60560, n60561, n60562, n60563,
    n60564, n60565, n60566, n60567, n60568, n60569,
    n60570, n60571, n60572, n60573, n60574, n60575,
    n60576, n60577, n60578, n60579, n60580, n60581,
    n60582, n60583, n60584, n60585, n60586, n60587,
    n60588, n60589, n60590, n60591, n60592, n60593,
    n60594, n60595, n60596, n60597, n60598, n60599,
    n60600, n60601, n60602, n60603, n60604, n60605,
    n60606, n60607, n60608, n60609, n60610, n60611,
    n60612, n60613, n60614, n60615, n60616, n60617,
    n60619, n60620, n60621, n60622, n60623, n60624,
    n60625, n60626, n60627, n60628, n60629, n60630,
    n60631, n60632, n60633, n60634, n60635, n60636,
    n60637, n60638, n60639, n60640, n60641, n60642,
    n60643, n60644, n60645, n60646, n60647, n60648,
    n60649, n60650, n60651, n60652, n60653, n60654,
    n60655, n60656, n60657, n60658, n60659, n60660,
    n60661, n60662, n60663, n60664, n60665, n60666,
    n60667, n60668, n60669, n60670, n60671, n60672,
    n60673, n60674, n60675, n60676, n60677, n60678,
    n60679, n60680, n60681, n60682, n60683, n60684,
    n60685, n60686, n60687, n60688, n60689, n60690,
    n60691, n60692, n60693, n60694, n60695, n60696,
    n60697, n60698, n60699, n60700, n60701, n60702,
    n60703, n60704, n60705, n60706, n60707, n60708,
    n60709, n60710, n60711, n60712, n60713, n60714,
    n60715, n60716, n60717, n60718, n60719, n60720,
    n60721, n60722, n60723, n60724, n60725, n60726,
    n60727, n60728, n60729, n60730, n60731, n60732,
    n60733, n60734, n60735, n60736, n60737, n60738,
    n60739, n60740, n60741, n60742, n60743, n60744,
    n60745, n60746, n60747, n60748, n60749, n60750,
    n60751, n60752, n60753, n60754, n60755, n60756,
    n60757, n60758, n60759, n60760, n60761, n60762,
    n60763, n60764, n60765, n60766, n60767, n60768,
    n60769, n60770, n60771, n60772, n60773, n60774,
    n60775, n60776, n60777, n60778, n60779, n60780,
    n60781, n60782, n60783, n60784, n60785, n60786,
    n60787, n60788, n60789, n60790, n60791, n60792,
    n60793, n60794, n60795, n60796, n60797, n60798,
    n60799, n60800, n60801, n60802, n60803, n60804,
    n60805, n60806, n60807, n60808, n60809, n60810,
    n60811, n60812, n60813, n60814, n60815, n60816,
    n60817, n60818, n60819, n60820, n60821, n60822,
    n60823, n60824, n60825, n60826, n60827, n60828,
    n60829, n60830, n60831, n60832, n60833, n60834,
    n60835, n60836, n60837, n60838, n60839, n60840,
    n60841, n60842, n60843, n60844, n60845, n60846,
    n60847, n60848, n60849, n60850, n60851, n60852,
    n60853, n60854, n60855, n60856, n60857, n60858,
    n60859, n60860, n60861, n60862, n60863, n60864,
    n60865, n60866, n60867, n60868, n60869, n60870,
    n60871, n60872, n60873, n60874, n60875, n60876,
    n60877, n60878, n60879, n60880, n60881, n60882,
    n60883, n60884, n60885, n60886, n60887, n60888,
    n60889, n60890, n60891, n60892, n60893, n60894,
    n60895, n60896, n60897, n60898, n60899, n60900,
    n60901, n60902, n60903, n60904, n60905, n60906,
    n60907, n60908, n60909, n60910, n60911, n60912,
    n60913, n60914, n60915, n60916, n60917, n60918,
    n60919, n60920, n60921, n60922, n60923, n60924,
    n60925, n60926, n60927, n60928, n60929, n60930,
    n60931, n60932, n60933, n60934, n60935, n60936,
    n60937, n60938, n60939, n60940, n60941, n60942,
    n60943, n60944, n60945, n60946, n60947, n60948,
    n60949, n60950, n60951, n60952, n60953, n60954,
    n60955, n60956, n60957, n60958, n60959, n60960,
    n60961, n60962, n60963, n60964, n60965, n60966,
    n60968, n60969, n60970, n60971, n60972, n60973,
    n60974, n60975, n60976, n60977, n60978, n60979,
    n60980, n60981, n60982, n60983, n60984, n60985,
    n60986, n60987, n60988, n60989, n60990, n60991,
    n60992, n60993, n60994, n60995, n60996, n60997,
    n60998, n60999, n61000, n61001, n61002, n61003,
    n61004, n61005, n61006, n61007, n61008, n61009,
    n61010, n61011, n61012, n61013, n61014, n61015,
    n61017, n61018, n61019, n61020, n61021, n61022,
    n61023, n61024, n61025, n61026, n61027, n61028,
    n61029, n61030, n61031, n61032, n61033, n61034,
    n61035, n61036, n61037, n61038, n61039, n61040,
    n61041, n61042, n61043, n61044, n61045, n61046,
    n61047, n61048, n61049, n61050, n61051, n61052,
    n61053, n61054, n61055, n61056, n61057, n61058,
    n61059, n61060, n61061, n61062, n61063, n61064,
    n61066, n61067, n61068, n61069, n61070, n61071,
    n61072, n61073, n61074, n61075, n61076, n61077,
    n61078, n61079, n61080, n61081, n61082, n61083,
    n61084, n61085, n61086, n61087, n61088, n61089,
    n61090, n61091, n61092, n61093, n61094, n61095,
    n61096, n61097, n61098, n61099, n61100, n61101,
    n61102, n61103, n61104, n61105, n61106, n61107,
    n61108, n61109, n61110, n61111, n61112, n61113,
    n61115, n61116, n61117, n61118, n61119, n61120,
    n61121, n61122, n61123, n61124, n61125, n61126,
    n61127, n61128, n61129, n61130, n61131, n61132,
    n61133, n61134, n61135, n61136, n61137, n61138,
    n61139, n61140, n61141, n61142, n61143, n61144,
    n61145, n61146, n61147, n61148, n61149, n61150,
    n61151, n61152, n61153, n61154, n61155, n61156,
    n61157, n61158, n61159, n61160, n61161, n61162,
    n61163, n61164, n61165, n61166, n61167, n61168,
    n61169, n61170, n61171, n61172, n61173, n61174,
    n61175, n61176, n61177, n61178, n61179, n61180,
    n61181, n61182, n61183, n61184, n61185, n61186,
    n61187, n61188, n61189, n61190, n61191, n61192,
    n61193, n61194, n61195, n61196, n61197, n61198,
    n61199, n61200, n61201, n61202, n61203, n61204,
    n61205, n61206, n61207, n61208, n61209, n61210,
    n61211, n61212, n61213, n61214, n61215, n61216,
    n61217, n61218, n61219, n61220, n61221, n61222,
    n61223, n61224, n61225, n61226, n61227, n61228,
    n61229, n61230, n61231, n61232, n61233, n61234,
    n61235, n61236, n61237, n61238, n61239, n61240,
    n61241, n61242, n61243, n61244, n61245, n61246,
    n61247, n61248, n61249, n61250, n61251, n61252,
    n61253, n61254, n61255, n61256, n61257, n61258,
    n61259, n61260, n61261, n61262, n61263, n61264,
    n61265, n61266, n61267, n61268, n61269, n61270,
    n61271, n61272, n61273, n61274, n61275, n61276,
    n61277, n61278, n61279, n61280, n61281, n61282,
    n61283, n61284, n61285, n61286, n61287, n61288,
    n61289, n61290, n61291, n61292, n61293, n61294,
    n61295, n61296, n61297, n61298, n61299, n61300,
    n61301, n61302, n61303, n61304, n61305, n61306,
    n61307, n61308, n61309, n61310, n61311, n61312,
    n61313, n61314, n61315, n61316, n61317, n61318,
    n61319, n61320, n61321, n61322, n61323, n61324,
    n61325, n61326, n61327, n61328, n61329, n61330,
    n61331, n61332, n61333, n61334, n61335, n61336,
    n61337, n61338, n61339, n61340, n61341, n61342,
    n61343, n61344, n61345, n61346, n61347, n61348,
    n61349, n61350, n61351, n61352, n61353, n61354,
    n61355, n61356, n61357, n61358, n61359, n61360,
    n61361, n61362, n61363, n61364, n61365, n61366,
    n61367, n61368, n61369, n61370, n61371, n61372,
    n61373, n61374, n61375, n61376, n61377, n61378,
    n61379, n61380, n61381, n61382, n61383, n61384,
    n61385, n61386, n61387, n61388, n61389, n61390,
    n61391, n61392, n61393, n61394, n61395, n61396,
    n61397, n61398, n61399, n61400, n61401, n61402,
    n61403, n61404, n61405, n61406, n61407, n61408,
    n61409, n61410, n61411, n61412, n61413, n61414,
    n61415, n61416, n61417, n61418, n61419, n61420,
    n61421, n61422, n61423, n61424, n61425, n61426,
    n61427, n61428, n61429, n61430, n61431, n61432,
    n61433, n61434, n61435, n61436, n61437, n61438,
    n61439, n61440, n61441, n61442, n61443, n61444,
    n61445, n61446, n61447, n61448, n61449, n61450,
    n61451, n61452, n61453, n61454, n61455, n61456,
    n61457, n61458, n61459, n61460, n61461, n61462,
    n61463, n61464, n61465, n61466, n61467, n61468,
    n61469, n61470, n61471, n61472, n61473, n61474,
    n61475, n61476, n61477, n61478, n61479, n61480,
    n61481, n61482, n61483, n61484, n61485, n61486,
    n61487, n61488, n61490, n61491, n61492, n61493,
    n61494, n61495, n61496, n61497, n61498, n61499,
    n61500, n61501, n61502, n61503, n61504, n61505,
    n61506, n61507, n61508, n61509, n61510, n61511,
    n61512, n61513, n61514, n61515, n61516, n61517,
    n61518, n61519, n61520, n61521, n61522, n61523,
    n61524, n61525, n61526, n61527, n61528, n61529,
    n61530, n61531, n61532, n61533, n61534, n61535,
    n61536, n61537, n61538, n61539, n61540, n61541,
    n61542, n61543, n61544, n61545, n61546, n61547,
    n61548, n61549, n61550, n61551, n61552, n61553,
    n61554, n61555, n61556, n61557, n61558, n61559,
    n61560, n61561, n61562, n61563, n61564, n61565,
    n61566, n61567, n61568, n61570, n61571, n61572,
    n61573, n61574, n61575, n61576, n61577, n61578,
    n61579, n61580, n61581, n61582, n61583, n61584,
    n61585, n61586, n61587, n61588, n61589, n61590,
    n61591, n61592, n61593, n61594, n61595, n61596,
    n61597, n61598, n61599, n61600, n61601, n61602,
    n61604, n61605, n61606, n61607, n61608, n61609,
    n61610, n61611, n61612, n61613, n61615, n61616,
    n61617, n61618, n61619, n61620, n61621, n61622,
    n61623, n61624, n61626, n61627, n61629, n61630,
    n61631, n61632, n61633, n61634, n61635, n61637,
    n61638, n61640, n61641, n61642, n61643, n61644,
    n61645, n61646, n61647, n61648, n61649, n61650,
    n61651, n61652, n61653, n61654, n61655, n61656,
    n61657, n61658, n61659, n61660, n61661, n61662,
    n61663, n61664, n61665, n61666, n61667, n61668,
    n61669, n61670, n61671, n61672, n61673, n61674,
    n61675, n61676, n61677, n61678, n61679, n61680,
    n61681, n61682, n61683, n61684, n61685, n61686,
    n61687, n61688, n61689, n61690, n61691, n61692,
    n61693, n61694, n61695, n61696, n61697, n61698,
    n61699, n61700, n61701, n61702, n61703, n61704,
    n61705, n61706, n61707, n61708, n61709, n61710,
    n61711, n61712, n61713, n61714, n61715, n61716,
    n61717, n61718, n61719, n61720, n61721, n61722,
    n61723, n61724, n61725, n61726, n61727, n61728,
    n61729, n61730, n61731, n61732, n61733, n61734,
    n61735, n61736, n61737, n61738, n61739, n61740,
    n61741, n61742, n61743, n61744, n61745, n61746,
    n61747, n61748, n61749, n61750, n61751, n61752,
    n61753, n61754, n61755, n61756, n61757, n61758,
    n61759, n61760, n61761, n61762, n61763, n61765,
    n61766, n61767, n61768, n61769, n61770, n61771,
    n61772, n61773, n61774, n61775, n61776, n61777,
    n61778, n61779, n61780, n61781, n61782, n61783,
    n61784, n61785, n61786, n61787, n61788, n61789,
    n61790, n61791, n61792, n61793, n61794, n61795,
    n61796, n61797, n61798, n61799, n61800, n61801,
    n61802, n61804, n61805, n61807, n61808, n61809,
    n61810, n61811, n61812, n61813, n61814, n61815,
    n61816, n61817, n61818, n61819, n61821, n61822,
    n61823, n61824, n61825, n61826, n61827, n61828,
    n61829, n61830, n61831, n61832, n61833, n61834,
    n61835, n61837, n61838, n61839, n61840, n61841,
    n61842, n61843, n61844, n61845, n61846, n61847,
    n61848, n61849, n61850, n61851, n61852, n61853,
    n61854, n61855, n61856, n61857, n61858, n61860,
    n61861, n61862, n61863, n61864, n61865, n61866,
    n61867, n61868, n61869, n61870, n61871, n61872,
    n61873, n61874, n61875, n61876, n61877, n61878,
    n61879, n61880, n61881, n61882, n61883, n61884,
    n61885, n61886, n61887, n61888, n61889, n61890,
    n61891, n61892, n61893, n61894, n61895, n61896,
    n61897, n61898, n61899, n61900, n61901, n61902,
    n61903, n61904, n61905, n61906, n61907, n61908,
    n61909, n61911, n61912, n61913, n61914, n61915,
    n61916, n61917, n61918, n61920, n61921, n61922,
    n61923, n61924, n61925, n61926, n61927, n61928,
    n61929, n61930, n61932, n61933, n61934, n61935,
    n61936, n61937, n61938, n61939, n61941, n61942,
    n61943, n61944, n61945, n61947, n61948, n61949,
    n61950, n61951, n61952, n61954, n61955, n61956,
    n61957, n61958, n61959, n61960, n61961, n61962,
    n61963, n61964, n61965, n61966, n61967, n61968,
    n61969, n61970, n61971, n61972, n61973, n61974,
    n61975, n61976, n61977, n61978, n61979, n61980,
    n61981, n61982, n61983, n61984, n61985, n61986,
    n61987, n61988, n61989, n61990, n61991, n61992,
    n61993, n61994, n61995, n61996, n61997, n61998,
    n61999, n62000, n62001, n62002, n62003, n62004,
    n62005, n62006, n62007, n62008, n62009, n62010,
    n62011, n62012, n62013, n62014, n62015, n62016,
    n62017, n62018, n62019, n62020, n62021, n62022,
    n62023, n62024, n62025, n62026, n62027, n62028,
    n62029, n62030, n62031, n62032, n62033, n62034,
    n62035, n62036, n62037, n62038, n62039, n62040,
    n62041, n62042, n62043, n62044, n62045, n62046,
    n62047, n62048, n62049, n62050, n62051, n62052,
    n62053, n62054, n62055, n62056, n62057, n62058,
    n62059, n62060, n62061, n62062, n62063, n62064,
    n62065, n62066, n62067, n62068, n62069, n62070,
    n62071, n62072, n62073, n62074, n62075, n62076,
    n62077, n62078, n62079, n62080, n62081, n62082,
    n62083, n62084, n62085, n62086, n62087, n62088,
    n62089, n62090, n62091, n62092, n62093, n62094,
    n62095, n62096, n62097, n62098, n62099, n62100,
    n62101, n62102, n62103, n62104, n62105, n62106,
    n62107, n62108, n62109, n62110, n62111, n62112,
    n62113, n62114, n62115, n62116, n62117, n62118,
    n62119, n62120, n62121, n62122, n62123, n62124,
    n62125, n62126, n62127, n62128, n62129, n62130,
    n62131, n62132, n62133, n62134, n62135, n62136,
    n62137, n62138, n62139, n62140, n62141, n62142,
    n62143, n62144, n62145, n62146, n62147, n62148,
    n62149, n62150, n62151, n62152, n62153, n62154,
    n62155, n62156, n62157, n62158, n62159, n62160,
    n62161, n62162, n62163, n62164, n62165, n62166,
    n62167, n62168, n62169, n62170, n62171, n62172,
    n62173, n62174, n62175, n62176, n62177, n62178,
    n62179, n62180, n62181, n62182, n62183, n62184,
    n62185, n62186, n62187, n62188, n62189, n62190,
    n62191, n62192, n62193, n62194, n62195, n62196,
    n62197, n62198, n62199, n62200, n62201, n62202,
    n62203, n62204, n62205, n62206, n62207, n62208,
    n62209, n62210, n62211, n62212, n62213, n62214,
    n62215, n62216, n62217, n62218, n62219, n62220,
    n62221, n62222, n62223, n62224, n62225, n62226,
    n62227, n62228, n62229, n62230, n62231, n62232,
    n62233, n62234, n62235, n62236, n62237, n62238,
    n62239, n62240, n62241, n62242, n62243, n62244,
    n62245, n62246, n62247, n62248, n62249, n62250,
    n62251, n62252, n62253, n62254, n62255, n62256,
    n62257, n62258, n62259, n62260, n62261, n62262,
    n62263, n62264, n62265, n62266, n62267, n62268,
    n62270, n62271, n62272, n62273, n62274, n62275,
    n62276, n62277, n62278, n62279, n62280, n62281,
    n62282, n62283, n62284, n62285, n62286, n62287,
    n62288, n62289, n62290, n62291, n62292, n62293,
    n62294, n62295, n62296, n62297, n62298, n62299,
    n62300, n62301, n62302, n62303, n62304, n62305,
    n62306, n62307, n62308, n62309, n62310, n62311,
    n62313, n62314, n62315, n62316, n62317, n62318,
    n62331, n62332, n62333, n62334, n62335, n62336,
    n62337, n62338, n62339, n62340, n62341, n62342,
    n62343, n62344, n62345, n62346, n62347, n62348,
    n62349, n62350, n62351, n62352, n62353, n62354,
    n62355, n62356, n62357, n62358, n62359, n62360,
    n62361, n62362, n62363, n62364, n62365, n62366,
    n62367, n62368, n62369, n62370, n62371, n62372,
    n62373, n62374, n62375, n62376, n62377, n62378,
    n62379, n62380, n62381, n62382, n62383, n62384,
    n62385, n62386, n62387, n62388, n62389, n62390,
    n62391, n62392, n62393, n62394, n62395, n62396,
    n62397, n62398, n62399, n62400, n62401, n62402,
    n62403, n62404, n62405, n62406, n62407, n62408,
    n62409, n62410, n62411, n62412, n62413, n62414,
    n62415, n62416, n62417, n62418, n62419, n62420,
    n62421, n62422, n62423, n62424, n62425, n62426,
    n62427, n62428, n62429, n62430, n62431, n62432,
    n62433, n62434, n62435, n62436, n62437, n62438,
    n62439, n62440, n62441, n62442, n62443, n62444,
    n62445, n62446, n62447, n62448, n62449, n62450,
    n62451, n62452, n62453, n62454, n62455, n62456,
    n62457, n62458, n62459, n62460, n62461, n62462,
    n62463, n62464, n62465, n62466, n62467, n62468,
    n62469, n62470, n62471, n62472, n62473, n62474,
    n62475, n62476, n62477, n62478, n62479, n62480,
    n62481, n62482, n62483, n62484, n62485, n62486,
    n62487, n62488, n62489, n62490, n62491, n62492,
    n62493, n62494, n62495, n62496, n62497, n62498,
    n62499, n62500, n62501, n62502, n62503, n62504,
    n62505, n62506, n62507, n62508, n62509, n62510,
    n62511, n62512, n62513, n62514, n62515, n62516,
    n62517, n62518, n62519, n62520, n62521, n62522,
    n62523, n62524, n62525, n62526, n62527, n62528,
    n62529, n62530, n62531, n62532, n62533, n62534,
    n62535, n62536, n62537, n62538, n62539, n62540,
    n62541, n62542, n62543, n62544, n62545, n62546,
    n62547, n62548, n62549, n62550, n62551, n62552,
    n62553, n62554, n62555, n62556, n62557, n62558,
    n62559, n62560, n62561, n62562, n62563, n62564,
    n62565, n62566, n62567, n62568, n62569, n62570,
    n62571, n62572, n62573, n62574, n62575, n62576,
    n62577, n62578, n62579, n62580, n62581, n62582,
    n62583, n62584, n62585, n62586, n62587, n62588,
    n62589, n62590, n62591, n62592, n62593, n62594,
    n62595, n62596, n62597, n62598, n62599, n62600,
    n62601, n62602, n62603, n62604, n62605, n62606,
    n62607, n62608, n62609, n62610, n62611, n62612,
    n62613, n62614, n62615, n62616, n62617, n62618,
    n62619, n62620, n62621, n62622, n62623, n62624,
    n62625, n62626, n62627, n62628, n62629, n62630,
    n62631, n62632, n62633, n62634, n62635, n62636,
    n62637, n62638, n62639, n62640, n62641, n62642,
    n62643, n62644, n62645, n62646, n62647, n62648,
    n62649, n62650, n62651, n62652, n62653, n62654,
    n62655, n62656, n62657, n62658, n62659, n62660,
    n62661, n62662, n62663, n62664, n62665, n62666,
    n62667, n62668, n62669, n62670, n62671, n62672,
    n62673, n62674, n62675, n62676, n62677, n62678,
    n62679, n62680, n62681, n62682, n62683, n62684,
    n62685, n62686, n62687, n62688, n62689, n62690,
    n62691, n62692, n62693, n62694, n62695, n62696,
    n62697, n62698, n62699, n62700, n62701, n62702,
    n62703, n62704, n62705, n62706, n62707, n62708,
    n62709, n62710, n62711, n62712, n62713, n62714,
    n62715, n62716, n62717, n62718, n62719, n62720,
    n62721, n62722, n62723, n62724, n62725, n62726,
    n62727, n62728, n62729, n62730, n62731, n62732,
    n62733, n62734, n62735, n62736, n62737, n62738,
    n62739, n62740, n62741, n62742, n62743, n62744,
    n62745, n62746, n62747, n62748, n62749, n62750,
    n62751, n62752, n62753, n62754, n62755, n62756,
    n62757, n62758, n62759, n62760, n62761, n62762,
    n62763, n62764, n62765, n62766, n62767, n62768,
    n62769, n62770, n62771, n62772, n62773, n62774,
    n62775, n62776, n62777, n62778, n62779, n62780,
    n62781, n62782, n62783, n62784, n62785, n62786,
    n62787, n62788, n62789, n62790, n62791, n62792,
    n62793, n62794, n62795, n62796, n62797, n62798,
    n62799, n62800, n62801, n62802, n62803, n62804,
    n62805, n62806, n62807, n62808, n62809, n62810,
    n62811, n62812, n62813, n62814, n62815, n62816,
    n62817, n62818, n62819, n62820, n62821, n62822,
    n62823, n62824, n62825, n62826, n62827, n62828,
    n62829, n62830, n62831, n62832, n62833, n62834,
    n62835, n62836, n62837, n62838, n62839, n62840,
    n62841, n62842, n62843, n62844, n62845, n62846,
    n62847, n62848, n62849, n62850, n62851, n62852,
    n62853, n62854, n62855, n62856, n62857, n62858,
    n62859, n62860, n62861, n62862, n62863, n62864,
    n62865, n62866, n62867, n62868, n62869, n62870,
    n62871, n62872, n62873, n62874, n62875, n62876,
    n62877, n62878, n62879, n62880, n62881, n62882,
    n62883, n62884, n62885, n62886, n62887, n62888,
    n62889, n62890, n62891, n62892, n62893, n62894,
    n62895, n62896, n62897, n62898, n62899, n62900,
    n62901, n62902, n62903, n62904, n62905, n62906,
    n62907, n62908, n62909, n62910, n62911, n62912,
    n62913, n62914, n62915, n62916, n62917, n62918,
    n62919, n62920, n62921, n62922, n62923, n62924,
    n62925, n62926, n62927, n62928, n62929, n62930,
    n62931, n62932, n62933, n62934, n62935, n62936,
    n62937, n62938, n62939, n62940, n62941, n62942,
    n62943, n62944, n62945, n62946, n62947, n62948,
    n62949, n62950, n62951, n62952, n62953, n62954,
    n62955, n62956, n62957, n62958, n62959, n62960,
    n62961, n62962, n62963, n62964, n62965, n62966,
    n62967, n62968, n62969, n62970, n62971, n62972,
    n62973, n62974, n62975, n62976, n62977, n62978,
    n62979, n62980, n62981, n62982, n62983, n62984,
    n62985, n62986, n62987, n62988, n62989, n62990,
    n62991, n62992, n62993, n62994, n62995, n62996,
    n62997, n62998, n62999, n63000, n63001, n63002,
    n63003, n63004, n63005, n63006, n63007, n63008,
    n63009, n63010, n63011, n63012, n63013, n63014,
    n63015, n63016, n63017, n63018, n63019, n63020,
    n63021, n63022, n63023, n63024, n63025, n63026,
    n63027, n63028, n63029, n63030, n63031, n63032,
    n63033, n63034, n63035, n63036, n63037, n63038,
    n63039, n63040, n63041, n63042, n63043, n63044,
    n63045, n63046, n63047, n63048, n63049, n63050,
    n63051, n63052, n63053, n63054, n63055, n63056,
    n63057, n63058, n63059, n63060, n63061, n63062,
    n63063, n63064, n63065, n63066, n63067, n63068,
    n63069, n63070, n63071, n63072, n63073, n63074,
    n63075, n63076, n63077, n63078, n63079, n63080,
    n63081, n63082, n63083, n63084, n63085, n63086,
    n63087, n63088, n63089, n63090, n63091, n63092,
    n63093, n63094, n63095, n63096, n63097, n63098,
    n63099, n63100, n63101, n63102, n63103, n63104,
    n63105, n63106, n63107, n63108, n63109, n63110,
    n63111, n63112, n63113, n63114, n63115, n63116,
    n63117, n63118, n63119, n63120, n63121, n63122,
    n63123, n63124, n63125, n63126, n63127, n63128,
    n63129, n63130, n63131, n63132, n63133, n63134,
    n63135, n63136, n63137, n63138, n63139, n63140,
    n63141, n63142, n63143, n63144, n63145, n63146,
    n63147, n63148, n63149, n63150, n63151, n63152,
    n63153, n63154, n63155, n63156, n63157, n63158,
    n63159, n63160, n63161, n63162, n63163, n63164,
    n63165, n63166, n63167, n63168, n63169, n63170,
    n63171, n63172, n63173, n63174, n63175, n63176,
    n63177, n63178, n63179, n63180, n63181, n63182,
    n63183, n63184, n63185, n63186, n63187, n63188,
    n63189, n63190, n63191, n63192, n63193, n63194,
    n63195, n63196, n63197, n63198, n63199, n63200,
    n63201, n63202, n63203, n63204, n63205, n63206,
    n63207, n63208, n63209, n63210, n63211, n63212,
    n63213, n63214, n63215, n63216, n63217, n63218,
    n63219, n63220, n63221, n63222, n63223, n63224,
    n63225, n63226, n63227, n63228, n63229, n63230,
    n63231, n63232, n63233, n63234, n63235, n63236,
    n63237, n63238, n63239, n63240, n63241, n63242,
    n63243, n63244, n63245, n63246, n63247, n63248,
    n63249, n63250, n63251, n63252, n63253, n63254,
    n63255, n63256, n63257, n63258, n63259, n63260,
    n63261, n63262, n63263, n63264, n63265, n63266,
    n63267, n63268, n63269, n63270, n63271, n63272,
    n63273, n63274, n63275, n63276, n63277, n63278,
    n63279, n63280, n63281, n63282, n63283, n63284,
    n63285, n63286, n63287, n63288, n63289, n63290,
    n63291, n63292, n63293, n63294, n63295, n63296,
    n63297, n63298, n63299, n63300, n63301, n63302,
    n63303, n63304, n63305, n63306, n63307, n63308,
    n63309, n63310, n63311, n63312, n63313, n63314,
    n63315, n63316, n63317, n63318, n63319, n63320,
    n63321, n63322, n63323, n63324, n63325, n63326,
    n63327, n63328, n63329, n63330, n63331, n63332,
    n63333, n63334, n63335, n63336, n63337, n63338,
    n63339, n63340, n63341, n63342, n63343, n63344,
    n63345, n63346, n63347, n63348, n63349, n63350,
    n63351, n63352, n63353, n63354, n63355, n63356,
    n63357, n63358, n63359, n63360, n63361, n63362,
    n63363, n63364, n63365, n63366, n63367, n63368,
    n63369, n63370, n63371, n63372, n63373, n63374,
    n63375, n63376, n63377, n63378, n63379, n63380,
    n63381, n63382, n63383, n63384, n63385, n63386,
    n63387, n63388, n63389, n63390, n63391, n63392,
    n63393, n63394, n63395, n63396, n63397, n63398,
    n63399, n63400, n63401, n63402, n63403, n63404,
    n63405, n63406, n63407, n63408, n63409, n63410,
    n63411, n63412, n63413, n63414, n63415, n63416,
    n63417, n63418, n63419, n63420, n63421, n63422,
    n63423, n63424, n63425, n63426, n63427, n63428,
    n63429, n63430, n63431, n63432, n63433, n63434,
    n63435, n63436, n63437, n63438, n63439, n63440,
    n63441, n63442, n63443, n63444, n63445, n63446,
    n63447, n63448, n63449, n63450, n63451, n63452,
    n63453, n63454, n63455, n63456, n63457, n63458,
    n63459, n63460, n63461, n63462, n63463, n63464,
    n63465, n63466, n63467, n63468, n63469, n63470,
    n63471, n63472, n63473, n63474, n63475, n63476,
    n63477, n63478, n63479, n63480, n63481, n63482,
    n63483, n63484, n63485, n63486, n63487, n63488,
    n63489, n63490, n63491, n63492, n63493, n63494,
    n63495, n63496, n63497, n63498, n63499, n63500,
    n63501, n63502, n63503, n63504, n63505, n63506,
    n63507, n63508, n63509, n63510, n63511, n63512,
    n63513, n63514, n63515, n63516, n63517, n63518,
    n63519, n63520, n63521, n63522, n63523, n63524,
    n63525, n63526, n63527, n63528, n63529, n63530,
    n63531, n63532, n63533, n63534, n63535, n63536,
    n63537, n63538, n63539, n63540, n63541, n63542,
    n63543, n63544, n63545, n63546, n63547, n63548,
    n63549, n63550, n63551, n63552, n63553, n63554,
    n63555, n63556, n63557, n63558, n63559, n63560,
    n63561, n63562, n63563, n63564, n63565, n63566,
    n63567, n63568, n63569, n63570, n63571, n63572,
    n63573, n63574, n63575, n63576, n63577, n63578,
    n63579, n63580, n63581, n63582, n63583, n63584,
    n63585, n63586, n63587, n63588, n63589, n63590,
    n63591, n63592, n63593, n63594, n63595, n63596,
    n63597, n63598, n63599, n63600, n63601, n63602,
    n63603, n63604, n63605, n63606, n63607, n63608,
    n63609, n63610, n63611, n63612, n63613, n63614,
    n63615, n63616, n63617, n63618, n63619, n63620,
    n63621, n63622, n63623, n63624, n63625, n63626,
    n63627, n63628, n63629, n63630, n63631, n63632,
    n63633, n63634, n63635, n63636, n63637, n63638,
    n63639, n63640, n63641, n63642, n63643, n63644,
    n63645, n63646, n63647, n63648, n63649, n63650,
    n63651, n63652, n63653, n63654, n63655, n63656,
    n63657, n63658, n63659, n63660, n63661, n63662,
    n63663, n63664, n63665, n63666, n63667, n63668,
    n63669, n63670, n63671, n63672, n63673, n63674,
    n63675, n63676, n63677, n63678, n63679, n63680,
    n63681, n63682, n63683, n63684, n63685, n63686,
    n63687, n63688, n63689, n63690, n63691, n63692,
    n63693, n63694, n63695, n63696, n63697, n63698,
    n63699, n63700, n63701, n63702, n63703, n63704,
    n63705, n63706, n63707, n63708, n63709, n63710,
    n63711, n63712, n63713, n63714, n63715, n63716,
    n63717, n63718, n63719, n63720, n63721, n63722,
    n63723, n63724, n63725, n63726, n63727, n63728,
    n63729, n63730, n63731, n63732, n63733, n63734,
    n63735, n63736, n63737, n63738, n63739, n63740,
    n63741, n63742, n63743, n63744, n63745, n63746,
    n63747, n63748, n63749, n63750, n63751, n63752,
    n63753, n63754, n63755, n63756, n63757, n63758,
    n63759, n63760, n63761, n63762, n63763, n63764,
    n63765, n63766, n63767, n63768, n63769, n63770,
    n63771, n63772, n63773, n63774, n63775, n63776,
    n63777, n63778, n63779, n63780, n63781, n63782,
    n63783, n63784, n63785, n63786, n63787, n63788,
    n63789, n63790, n63791, n63792, n63793, n63794,
    n63795, n63796, n63797, n63798, n63799, n63800,
    n63801, n63802, n63803, n63804, n63805, n63806,
    n63807, n63808, n63809, n63811, n63812, n63813,
    n63814, n63815, n63816, n63817, n63818, n63819,
    n63820, n63821, n63822, n63823, n63824, n63825,
    n63826, n63827, n63828, n63829, n63830, n63831,
    n63833, n63834, n63835, n63836, n63837, n63838,
    n63839, n63840, n63841, n63842, n63843, n63844,
    n63845, n63846, n63847, n63848, n63849, n63850,
    n63851, n63852, n63853, n63854, n63855, n63856,
    n63857, n63858, n63859, n63860, n63861, n63862,
    n63863, n63864, n63865, n63866, n63867, n63868,
    n63869, n63870, n63871, n63872, n63873, n63874,
    n63875, n63876, n63877, n63879, n63880, n63881,
    n63882, n63883, n63885, n63886, n63887, n63888,
    n63889, n63890, n63891, n63892, n63893, n63894,
    n63895, n63896, n63897, n63898, n63899, n63900,
    n63901, n63902, n63903, n63904, n63905, n63906,
    n63907, n63908, n63909, n63910, n63911, n63912,
    n63913, n63914, n63915, n63916, n63917, n63918,
    n63919, n63920, n63921, n63922, n63923, n63924,
    n63925, n63926, n63927, n63928, n63929, n63930,
    n63931, n63932, n63933, n63934, n63935, n63936,
    n63937, n63938, n63939, n63940, n63941, n63942,
    n63943, n63944, n63945, n63946, n63947, n63948,
    n63949, n63950, n63951, n63952, n63953, n63954,
    n63955, n63956, n63957, n63958, n63959, n63960,
    n63961, n63962, n63963, n63964, n63965, n63966,
    n63967, n63968, n63969, n63970, n63971, n63972,
    n63973, n63974, n63975, n63976, n63977, n63978,
    n63979, n63980, n63981, n63982, n63983, n63984,
    n63985, n63986, n63987, n63988, n63989, n63991,
    n63992, n63993, n63994, n63995, n63996, n63997,
    n63998, n63999, n64000, n64001, n64002, n64003,
    n64004, n64005, n64006, n64007, n64008, n64009,
    n64010, n64011, n64012, n64013, n64014, n64015,
    n64016, n64017, n64018, n64019, n64020, n64021,
    n64022, n64023, n64024, n64025, n64026, n64027,
    n64028, n64029, n64030, n64031, n64032, n64033,
    n64034, n64035, n64036, n64037, n64038, n64039,
    n64040, n64041, n64042, n64043, n64044, n64045,
    n64046, n64047, n64048, n64049, n64050, n64051,
    n64052, n64053, n64054, n64055, n64056, n64057,
    n64058, n64059, n64060, n64061, n64062, n64063,
    n64064, n64065, n64066, n64067, n64068, n64069,
    n64070, n64071, n64072, n64073, n64074, n64075,
    n64076, n64077, n64078, n64079, n64080, n64081,
    n64082, n64083, n64084, n64085, n64086, n64087,
    n64088, n64089, n64090, n64091, n64092, n64093,
    n64094, n64095, n64096, n64097, n64098, n64099,
    n64100, n64101, n64102, n64103, n64104, n64105,
    n64106, n64107, n64108, n64109, n64110, n64111,
    n64112, n64113, n64114, n64115, n64116, n64117,
    n64118, n64119, n64120, n64121, n64122, n64123,
    n64124, n64125, n64126, n64127, n64128, n64129,
    n64130, n64131, n64132, n64133, n64134, n64135,
    n64136, n64137, n64138, n64139, n64140, n64141,
    n64142, n64143, n64144, n64145, n64146, n64147,
    n64148, n64149, n64150, n64151, n64152, n64153,
    n64154, n64155, n64156, n64157, n64158, n64159,
    n64160, n64161, n64162, n64163, n64164, n64165,
    n64166, n64167, n64168, n64169, n64170, n64171,
    n64172, n64173, n64174, n64175, n64176, n64177,
    n64178, n64179, n64180, n64181, n64182, n64183,
    n64184, n64185, n64186, n64187, n64188, n64189,
    n64190, n64191, n64192, n64193, n64194, n64195,
    n64196, n64197, n64198, n64199, n64200, n64201,
    n64202, n64203, n64204, n64205, n64206, n64207,
    n64208, n64209, n64210, n64211, n64212, n64213,
    n64214, n64215, n64216, n64217, n64218, n64219,
    n64220, n64221, n64222, n64223, n64224, n64225,
    n64226, n64227, n64228, n64229, n64230, n64231,
    n64232, n64233, n64234, n64235, n64236, n64237,
    n64238, n64239, n64240, n64241, n64242, n64243,
    n64244, n64245, n64246, n64247, n64248, n64249,
    n64250, n64251, n64252, n64253, n64254, n64255,
    n64256, n64257, n64258, n64259, n64260, n64261,
    n64262, n64263, n64264, n64265, n64266, n64267,
    n64268, n64269, n64270, n64271, n64272, n64273,
    n64274, n64275, n64276, n64277, n64278, n64279,
    n64280, n64281, n64282, n64283, n64284, n64285,
    n64286, n64287, n64288, n64289, n64290, n64291,
    n64292, n64293, n64294, n64295, n64296, n64297,
    n64298, n64299, n64300, n64301, n64302, n64303,
    n64304, n64305, n64306, n64307, n64308, n64309,
    n64310, n64311, n64312, n64313, n64314, n64315,
    n64316, n64317, n64319, n64320, n64321, n64322,
    n64323, n64324, n64325, n64326, n64327, n64328,
    n64329, n64330, n64331, n64332, n64333, n64334,
    n64335, n64336, n64337, n64338, n64339, n64340,
    n64341, n64342, n64343, n64344, n64345, n64346,
    n64347, n64348, n64349, n64350, n64351, n64352,
    n64353, n64354, n64355, n64356, n64357, n64358,
    n64359, n64360, n64361, n64362, n64363, n64364,
    n64365, n64366, n64367, n64368, n64369, n64370,
    n64371, n64372, n64373, n64374, n64375, n64376,
    n64377, n64378, n64379, n64380, n64381, n64382,
    n64383, n64384, n64385, n64386, n64387, n64388,
    n64389, n64390, n64391, n64392, n64393, n64394,
    n64395, n64396, n64397, n64398, n64399, n64400,
    n64401, n64402, n64403, n64404, n64405, n64406,
    n64407, n64408, n64409, n64410, n64411, n64412,
    n64413, n64414, n64415, n64416, n64417, n64418,
    n64419, n64420, n64421, n64422, n64423, n64424,
    n64425, n64426, n64427, n64428, n64429, n64430,
    n64431, n64432, n64433, n64434, n64435, n64436,
    n64437, n64438, n64439, n64440, n64441, n64442,
    n64443, n64444, n64445, n64446, n64447, n64448,
    n64449, n64450, n64451, n64452, n64453, n64454,
    n64455, n64456, n64457, n64458, n64459, n64460,
    n64461, n64462, n64463, n64464, n64465, n64466,
    n64467, n64468, n64469, n64470, n64471, n64472,
    n64473, n64474, n64475, n64476, n64477, n64478,
    n64479, n64480, n64481, n64482, n64483, n64484,
    n64485, n64486, n64487, n64488, n64489, n64490,
    n64491, n64492, n64493, n64494, n64495, n64496,
    n64497, n64498, n64499, n64500, n64501, n64502,
    n64503, n64504, n64505, n64506, n64507, n64508,
    n64509, n64510, n64511, n64512, n64513, n64514,
    n64515, n64516, n64517, n64518, n64519, n64520,
    n64521, n64522, n64523, n64524, n64525, n64526,
    n64527, n64528, n64529, n64530, n64531, n64532,
    n64533, n64534, n64535, n64536, n64537, n64538,
    n64539, n64540, n64541, n64542, n64543, n64544,
    n64545, n64546, n64547, n64548, n64549, n64550,
    n64551, n64552, n64553, n64554, n64555, n64556,
    n64557, n64558, n64559, n64560, n64561, n64562,
    n64563, n64564, n64565, n64566, n64567, n64568,
    n64569, n64570, n64571, n64572, n64573, n64574,
    n64575, n64576, n64577, n64578, n64579, n64580,
    n64581, n64582, n64583, n64585, n64586, n64587,
    n64588, n64589, n64590, n64591, n64592, n64593,
    n64594, n64595, n64596, n64597, n64598, n64599,
    n64600, n64601, n64602, n64603, n64604, n64605,
    n64606, n64607, n64608, n64609, n64610, n64611,
    n64612, n64613, n64614, n64615, n64616, n64617,
    n64618, n64619, n64620, n64621, n64622, n64623,
    n64624, n64625, n64626, n64627, n64628, n64629,
    n64630, n64631, n64632, n64633, n64634, n64635,
    n64636, n64637, n64638, n64639, n64640, n64641,
    n64642, n64643, n64644, n64645, n64646, n64647,
    n64648, n64649, n64650, n64651, n64652, n64653,
    n64654, n64655, n64656, n64657, n64658, n64659,
    n64660, n64661, n64662, n64663, n64664, n64665,
    n64666, n64667, n64668, n64669, n64670, n64671,
    n64672, n64673, n64674, n64675, n64676, n64677,
    n64678, n64679, n64680, n64681, n64682, n64683,
    n64684, n64685, n64686, n64688, n64689, n64690,
    n64691, n64692, n64693, n64694, n64695, n64696,
    n64697, n64698, n64699, n64700, n64701, n64702,
    n64703, n64704, n64705, n64706, n64707, n64708,
    n64709, n64710, n64711, n64713, n64714, n64715,
    n64716, n64717, n64718, n64719, n64720, n64721,
    n64722, n64723, n64724, n64725, n64726, n64727,
    n64728, n64729, n64730, n64731, n64732, n64733,
    n64734, n64735, n64736, n64737, n64738, n64739,
    n64740, n64741, n64742, n64743, n64744, n64745,
    n64746, n64747, n64748, n64749, n64750, n64751,
    n64752, n64753, n64754, n64755, n64756, n64757,
    n64758, n64759, n64760, n64761, n64762, n64763,
    n64764, n64765, n64766, n64767, n64768, n64769,
    n64770, n64771, n64772, n64773, n64774, n64775,
    n64776, n64777, n64778, n64779, n64780, n64781,
    n64782, n64783, n64784, n64785, n64786, n64787,
    n64788, n64789, n64790, n64791, n64792, n64793,
    n64794, n64795, n64796, n64797, n64798, n64799,
    n64800, n64801, n64802, n64803, n64804, n64805,
    n64806, n64807, n64808, n64809, n64810, n64811,
    n64812, n64813, n64814, n64815, n64816, n64817,
    n64818, n64819, n64820, n64821, n64822, n64823,
    n64824, n64825, n64826, n64827, n64828, n64829,
    n64830, n64831, n64832, n64833, n64834, n64835,
    n64836, n64837, n64838, n64839, n64840, n64841,
    n64842, n64843, n64844, n64845, n64846, n64847,
    n64848, n64849, n64850, n64851, n64852, n64853,
    n64854, n64855, n64856, n64857, n64858, n64860,
    n64861, n64862, n64863, n64864, n64865, n64866,
    n64867, n64868, n64869, n64870, n64871, n64872,
    n64873, n64874, n64875, n64876, n64877, n64878,
    n64879, n64880, n64881, n64882, n64883, n64884,
    n64885, n64886, n64887, n64888, n64889, n64890,
    n64891, n64892, n64893, n64894, n64895, n64896,
    n64897, n64898, n64899, n64900, n64901, n64902,
    n64903, n64905, n64906, n64907, n64908, n64909,
    n64910, n64911, n64912, n64914, n64915, n64916,
    n64917, n64918, n64919, n64920, n64921, n64922,
    n64923, n64924, n64925, n64926, n64927, n64928,
    n64930, n64931, n64932, n64933, n64934, n64935,
    n64936, n64937, n64939, n64940, n64941, n64942,
    n64943, n64944, n64945, n64946, n64947, n64948,
    n64949, n64950, n64951, n64952, n64953, n64954,
    n64955, n64956, n64957, n64958, n64959, n64960,
    n64961, n64962, n64963, n64964, n64965, n64966,
    n64967, n64968, n64969, n64970, n64971, n64973,
    n64974, n64975, n64976, n64977, n64978, n64979,
    n64980, n64981, n64982, n64983, n64984, n64985,
    n64986, n64987, n64988, n64989, n64990, n64991,
    n64992, n64994, n64995, n64996, n64997, n65000,
    n65001, n65002, n65003, n65004, n65005, n65006,
    n65007, n65008, n65009, n65010, n65011, n65012,
    n65013, n65014, n65015, n65016, n65017, n65018,
    n65019, n65020, n65021, n65022, n65023, n65024,
    n65025, n65026, n65027, n65028, n65029, n65030,
    n65031, n65032, n65033, n65034, n65035, n65036,
    n65037, n65038, n65039, n65040, n65041, n65042,
    n65043, n65044, n65046, n65047, n65048, n65049,
    n65050, n65051, n65052, n65053, n65055, n65058,
    n65059, n65060, n65062, n65063, n65065, n65066,
    n65068, n65070, n65071, n65072, n65074, n65075,
    n65076, n65077, n65078, n65079, n65081, n65082,
    n65083, n65084, n65086, n65087, n65088, n65089,
    n65090, n65091, n65092, n65093, n65094, n65095,
    n65096, n65097, n65098, n65099, n65100, n65101,
    n65102, n65103, n65104, n65105, n65106, n65107,
    n65108, n65109, n65110, n65111, n65112, n65113,
    n65114, n65115, n65116, n65117, n65118, n65119,
    n65120, n65121, n65122, n65123, n65124, n65125,
    n65126, n65127, n65128, n65129, n65130, n65131,
    n65132, n65133, n65134, n65135, n65136, n65137,
    n65138, n65139, n65140, n65141, n65142, n65143,
    n65144, n65145, n65146, n65147, n65148, n65149,
    n65150, n65151, n65152, n65153, n65154, n65155,
    n65156, n65157, n65158, n65159, n65160, n65161,
    n65162, n65163, n65164, n65165, n65166, n65167,
    n65168, n65169, n65170, n65171, n65172, n65173,
    n65174, n65175, n65176, n65177, n65178, n65179,
    n65180, n65181, n65182, n65183, n65184, n65185,
    n65186, n65187, n65188, n65189, n65190, n65191,
    n65192, n65193, n65194, n65195, n65196, n65197,
    n65198, n65199, n65200, n65201, n65202, n65203,
    n65204, n65205, n65206, n65207, n65208, n65209,
    n65210, n65211, n65212, n65213, n65214, n65215,
    n65216, n65217, n65218, n65219, n65220, n65221,
    n65222, n65223, n65224, n65225, n65226, n65227,
    n65228, n65229, n65230, n65231, n65232, n65233,
    n65234, n65235, n65236, n65237, n65238, n65239,
    n65240, n65241, n65242, n65243, n65244, n65245,
    n65246, n65247, n65248, n65249, n65250, n65251,
    n65252, n65253, n65254, n65255, n65256, n65257,
    n65258, n65259, n65260, n65261, n65262, n65263,
    n65264, n65265, n65266, n65267, n65268, n65269,
    n65270, n65271, n65272, n65273, n65274, n65275,
    n65276, n65277, n65278, n65279, n65280, n65281,
    n65282, n65283, n65284, n65285, n65286, n65287,
    n65288, n65289, n65290, n65291, n65292, n65293,
    n65294, n65295, n65296, n65297, n65298, n65299,
    n65300, n65301, n65302, n65303, n65304, n65305,
    n65306, n65307, n65308, n65309, n65310, n65311,
    n65312, n65313, n65314, n65315, n65316, n65317,
    n65318, n65319, n65320, n65321, n65322, n65323,
    n65324, n65325, n65326, n65327, n65328, n65329,
    n65330, n65331, n65332, n65333, n65334, n65335,
    n65336, n65337, n65338, n65339, n65340, n65341,
    n65342, n65343, n65344, n65345, n65346, n65347,
    n65348, n65349, n65350, n65351, n65352, n65353,
    n65354, n65355, n65356, n65357, n65358, n65359,
    n65360, n65361, n65362, n65363, n65364, n65365,
    n65366, n65367, n65368, n65369, n65370, n65371,
    n65372, n65373, n65374, n65375, n65376, n65377,
    n65378, n65379, n65380, n65381, n65382, n65383,
    n65384, n65385, n65386, n65387, n65388, n65389,
    n65390, n65391, n65392, n65393, n65394, n65395,
    n65396, n65397, n65398, n65399, n65400, n65401,
    n65402, n65403, n65404, n65405, n65406, n65407,
    n65408, n65409, n65410, n65411, n65412, n65413,
    n65414, n65415, n65416, n65417, n65418, n65419,
    n65420, n65421, n65422, n65423, n65424, n65425,
    n65426, n65427, n65428, n65429, n65430, n65431,
    n65432, n65433, n65434, n65435, n65436, n65437,
    n65438, n65439, n65440, n65441, n65442, n65443,
    n65444, n65445, n65446, n65447, n65448, n65449,
    n65450, n65451, n65452, n65453, n65454, n65455,
    n65456, n65457, n65458, n65459, n65460, n65461,
    n65462, n65463, n65464, n65465, n65466, n65467,
    n65468, n65469, n65470, n65471, n65472, n65473,
    n65474, n65475, n65476, n65477, n65478, n65479,
    n65480, n65481, n65482, n65483, n65484, n65485,
    n65486, n65487, n65488, n65489, n65490, n65491,
    n65492, n65493, n65494, n65495, n65496, n65497,
    n65498, n65499, n65500, n65501, n65502, n65503,
    n65504, n65505, n65506, n65507, n65508, n65509,
    n65510, n65511, n65512, n65513, n65514, n65515,
    n65516, n65517, n65518, n65519, n65520, n65521,
    n65522, n65523, n65524, n65525, n65526, n65527,
    n65528, n65529, n65530, n65531, n65532, n65533,
    n65534, n65535, n65536, n65537, n65538, n65539,
    n65540, n65541, n65542, n65543, n65544, n65545,
    n65546, n65547, n65548, n65549, n65550, n65551,
    n65552, n65553, n65554, n65555, n65556, n65557,
    n65558, n65559, n65560, n65561, n65562, n65563,
    n65564, n65565, n65566, n65567, n65568, n65569,
    n65570, n65571, n65572, n65573, n65574, n65575,
    n65576, n65577, n65578, n65579, n65580, n65581,
    n65582, n65583, n65584, n65585, n65586, n65587,
    n65588, n65589, n65590, n65591, n65592, n65593,
    n65594, n65595, n65596, n65597, n65598, n65599,
    n65600, n65601, n65602, n65603, n65604, n65605,
    n65606, n65607, n65608, n65609, n65610, n65611,
    n65612, n65613, n65614, n65615, n65616, n65617,
    n65618, n65619, n65620, n65621, n65622, n65623,
    n65624, n65625, n65626, n65627, n65628, n65629,
    n65630, n65631, n65632, n65633, n65634, n65635,
    n65636, n65637, n65638, n65639, n65640, n65641,
    n65642, n65643, n65644, n65645, n65646, n65647,
    n65648, n65649, n65650, n65651, n65652, n65653,
    n65654, n65655, n65656, n65657, n65658, n65659,
    n65660, n65661, n65662, n65663, n65664, n65665,
    n65666, n65667, n65668, n65669, n65670, n65671,
    n65672, n65673, n65674, n65675, n65676, n65677,
    n65678, n65679, n65680, n65681, n65682, n65683,
    n65684, n65685, n65686, n65687, n65688, n65689,
    n65690, n65691, n65692, n65693, n65694, n65695,
    n65696, n65697, n65698, n65699, n65700, n65701,
    n65702, n65703, n65704, n65705, n65706, n65707,
    n65708, n65709, n65710, n65711, n65712, n65713,
    n65714, n65715, n65719, n65720, n65721, n65722,
    n65723, n65724, n65725, n65727, n65729, n65730,
    n65731, n65732, n65733, n65735, n65736, n65737,
    n65738, n65739, n65741, n65742, n65744, n65745,
    n65747, n65748, n65750, n65751, n65752, n65753,
    n65754, n65755, n65756, n65757, n65758, n65759,
    n65760, n65761, n65762, n65763, n65764, n65765,
    n65766, n65767, n65768, n65769, n65770, n65771,
    n65772, n65773, n65774, n65775, n65776, n65777,
    n65778, n65779, n65780, n65781, n65782, n65783,
    n65784, n65785, n65786, n65787, n65788, n65789,
    n65790, n65791, n65792, n65793, n65794, n65795,
    n65796, n65797, n65798, n65799, n65800, n65801,
    n65802, n65803, n65804, n65883, n65884, n65885,
    n65886, n65887, n65888, n65889, n65890, n65891,
    n65892, n65893, n65894, n65895, n65896, n65897,
    n65898, n65899, n65900, n65901, n65902, n65903,
    n65904, n65905, n65906, n65907, n65908, n65909,
    n65910, n65911, n65912, n65913, n65914, n65915,
    n65916, n65917, n65918, n65934, n65935, n65936,
    n65937, n65938, n65939, n65940, n65941, n65942,
    n65943, n65944, n65945, n65946, n65947, n65948,
    n65949, n65950, n65951, n65952, n65953, n65954,
    n65955, n65957, n65958, n65959, n65960, n65961,
    n65962, n65963, n65964, n65965, n65966, n65975,
    n65976, n65978, n65984, n65985, n65986, n65987,
    n65988, n65989, n65990, n65991, n65992, n65993,
    n65994, n65996, n65997, n65998, n65999, n66000,
    n66001, n66002, n66035, n66036, n66037, n66038,
    n66039, n66040, n66041;
  assign po166 = 1'b1;
  assign n2437 = ~pi426 & ~pi430;
  assign n2438 = pi426 & pi430;
  assign n2439 = pi426 & ~pi430;
  assign n2440 = ~pi426 & pi430;
  assign n2441 = ~n2439 & ~n2440;
  assign n2442 = ~n2437 & ~n2438;
  assign n2443 = pi427 & ~pi428;
  assign n2444 = ~pi427 & pi428;
  assign n2445 = ~pi427 & ~pi428;
  assign n2446 = pi427 & pi428;
  assign n2447 = ~n2445 & ~n2446;
  assign n2448 = ~n2443 & ~n2444;
  assign n2449 = pi417 & ~pi464;
  assign n2450 = ~pi417 & pi464;
  assign n2451 = ~n2449 & ~n2450;
  assign n2452 = pi437 & ~pi453;
  assign n2453 = ~pi437 & pi453;
  assign n2454 = ~pi437 & ~pi453;
  assign n2455 = pi437 & pi453;
  assign n2456 = ~n2454 & ~n2455;
  assign n2457 = ~n2452 & ~n2453;
  assign n2458 = pi418 & n62333;
  assign n2459 = ~pi418 & ~n62333;
  assign n2460 = ~n2458 & ~n2459;
  assign n2461 = n2451 & n2460;
  assign n2462 = ~n2451 & ~n2460;
  assign n2463 = ~pi417 & ~pi418;
  assign n2464 = pi417 & pi418;
  assign n2465 = pi417 & ~pi418;
  assign n2466 = ~pi417 & pi418;
  assign n2467 = ~n2465 & ~n2466;
  assign n2468 = ~n2463 & ~n2464;
  assign n2469 = pi464 & n62333;
  assign n2470 = ~pi464 & ~n62333;
  assign n2471 = ~n2469 & ~n2470;
  assign n2472 = n62334 & n2471;
  assign n2473 = ~n62334 & ~n2471;
  assign n2474 = ~n2472 & ~n2473;
  assign n2475 = pi464 & n62334;
  assign n2476 = ~pi464 & ~n62334;
  assign n2477 = ~n2475 & ~n2476;
  assign n2478 = ~n62333 & n2477;
  assign n2479 = n62333 & ~n2477;
  assign n2480 = ~n2478 & ~n2479;
  assign n2481 = pi437 & ~n62334;
  assign n2482 = ~pi437 & n62334;
  assign n2483 = ~n2481 & ~n2482;
  assign n2484 = pi453 & ~pi464;
  assign n2485 = ~pi453 & pi464;
  assign n2486 = ~n2484 & ~n2485;
  assign n2487 = n2483 & n2486;
  assign n2488 = ~n2483 & ~n2486;
  assign n2489 = ~n2487 & ~n2488;
  assign n2490 = ~n2461 & ~n2462;
  assign n2491 = pi415 & ~pi431;
  assign n2492 = ~pi415 & pi431;
  assign n2493 = ~pi415 & ~pi431;
  assign n2494 = pi415 & pi431;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = ~n2491 & ~n2492;
  assign n2497 = pi416 & ~pi438;
  assign n2498 = ~pi416 & pi438;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = ~n62336 & n2499;
  assign n2501 = n62336 & ~n2499;
  assign n2502 = n62336 & n2499;
  assign n2503 = ~n62336 & ~n2499;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = ~n2500 & ~n2501;
  assign n2506 = n62335 & n62337;
  assign n2507 = ~n62335 & ~n62337;
  assign n2508 = pi1197 & ~n2507;
  assign n2509 = pi1197 & ~n2506;
  assign n2510 = ~n2507 & n2509;
  assign n2511 = ~n2506 & n2508;
  assign n2512 = ~pi421 & ~pi454;
  assign n2513 = pi421 & pi454;
  assign n2514 = pi421 & ~pi454;
  assign n2515 = ~pi421 & pi454;
  assign n2516 = ~n2514 & ~n2515;
  assign n2517 = ~n2512 & ~n2513;
  assign n2518 = pi432 & ~pi459;
  assign n2519 = ~pi432 & pi459;
  assign n2520 = ~n2518 & ~n2519;
  assign n2521 = n62339 & ~n2520;
  assign n2522 = ~n62339 & n2520;
  assign n2523 = ~n2521 & ~n2522;
  assign n2524 = pi419 & ~pi420;
  assign n2525 = ~pi419 & pi420;
  assign n2526 = ~pi419 & ~pi420;
  assign n2527 = pi419 & pi420;
  assign n2528 = ~n2526 & ~n2527;
  assign n2529 = ~n2524 & ~n2525;
  assign n2530 = pi423 & ~pi424;
  assign n2531 = ~pi423 & pi424;
  assign n2532 = ~pi423 & ~pi424;
  assign n2533 = pi423 & pi424;
  assign n2534 = ~n2532 & ~n2533;
  assign n2535 = ~n2530 & ~n2531;
  assign n2536 = n62340 & n62341;
  assign n2537 = ~n62340 & ~n62341;
  assign n2538 = ~n2536 & ~n2537;
  assign n2539 = n2523 & n2538;
  assign n2540 = ~n2523 & ~n2538;
  assign n2541 = n2520 & ~n62341;
  assign n2542 = ~n2520 & n62341;
  assign n2543 = ~n2541 & ~n2542;
  assign n2544 = ~n62339 & ~n2543;
  assign n2545 = n62339 & n2543;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = ~n62340 & n2546;
  assign n2548 = n62340 & ~n2546;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = pi459 & ~n62340;
  assign n2551 = ~pi459 & n62340;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = pi432 & n62341;
  assign n2554 = ~pi432 & ~n62341;
  assign n2555 = ~n2553 & ~n2554;
  assign n2556 = ~n2552 & n2555;
  assign n2557 = n2552 & ~n2555;
  assign n2558 = ~n2556 & ~n2557;
  assign n2559 = n62339 & n2558;
  assign n2560 = ~n62339 & ~n2558;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = pi432 & ~n62339;
  assign n2563 = ~pi432 & n62339;
  assign n2564 = ~n2562 & ~n2563;
  assign n2565 = ~n62341 & ~n2564;
  assign n2566 = n62341 & n2564;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = n2552 & n2567;
  assign n2569 = ~n2552 & ~n2567;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = ~n2539 & ~n2540;
  assign n2572 = pi425 & n62342;
  assign n2573 = ~pi425 & ~n62342;
  assign n2574 = pi1198 & ~n2573;
  assign n2575 = pi1198 & ~n2572;
  assign n2576 = ~n2573 & n2575;
  assign n2577 = ~n2572 & n2574;
  assign n2578 = ~n62338 & ~n62343;
  assign n2579 = ~pi54 & ~pi92;
  assign n2580 = ~pi74 & n2579;
  assign n2581 = ~pi122 & pi829;
  assign n2582 = pi950 & pi1092;
  assign n2583 = ~pi824 & ~pi829;
  assign n2584 = n2582 & ~n2583;
  assign n2585 = ~pi35 & ~pi70;
  assign n2586 = ~pi58 & ~pi90;
  assign n2587 = ~pi63 & ~pi107;
  assign n2588 = ~pi83 & ~pi103;
  assign n2589 = ~pi61 & ~pi76;
  assign n2590 = ~pi85 & ~pi106;
  assign n2591 = n2589 & n2590;
  assign n2592 = ~pi48 & n2591;
  assign n2593 = ~pi89 & n2592;
  assign n2594 = ~pi49 & n2593;
  assign n2595 = ~pi104 & n2594;
  assign n2596 = ~pi45 & n2595;
  assign n2597 = ~pi68 & ~pi84;
  assign n2598 = ~pi82 & ~pi111;
  assign n2599 = ~pi36 & n2598;
  assign n2600 = n2597 & n2599;
  assign n2601 = ~pi66 & ~pi73;
  assign n2602 = n2600 & n2601;
  assign n2603 = n2596 & n2600;
  assign n2604 = n2601 & n2603;
  assign n2605 = n2596 & n2602;
  assign n2606 = ~pi67 & ~pi69;
  assign n2607 = ~pi67 & n62344;
  assign n2608 = ~pi69 & n2607;
  assign n2609 = n62344 & n2606;
  assign n2610 = n2588 & n62345;
  assign n2611 = ~pi88 & ~pi98;
  assign n2612 = ~pi77 & n2611;
  assign n2613 = ~pi50 & n2612;
  assign n2614 = ~pi81 & ~pi102;
  assign n2615 = ~pi64 & ~pi65;
  assign n2616 = ~pi64 & ~pi81;
  assign n2617 = ~pi65 & ~pi102;
  assign n2618 = n2616 & n2617;
  assign n2619 = n2614 & n2615;
  assign n2620 = ~pi65 & ~pi71;
  assign n2621 = ~pi102 & n2616;
  assign n2622 = n2620 & n2621;
  assign n2623 = ~pi71 & n62346;
  assign n2624 = n2613 & n62347;
  assign n2625 = n2610 & n2620;
  assign n2626 = ~pi102 & n2613;
  assign n2627 = n2616 & n2626;
  assign n2628 = n2625 & n2627;
  assign n2629 = n2610 & n2624;
  assign n2630 = n2587 & n2625;
  assign n2631 = n2627 & n2630;
  assign n2632 = ~pi64 & n2630;
  assign n2633 = ~pi81 & n2632;
  assign n2634 = n2626 & n2633;
  assign n2635 = n2587 & n62348;
  assign n2636 = ~pi47 & ~pi91;
  assign n2637 = ~pi53 & ~pi60;
  assign n2638 = ~pi86 & n2637;
  assign n2639 = ~pi97 & ~pi108;
  assign n2640 = ~pi94 & n2639;
  assign n2641 = ~pi109 & ~pi110;
  assign n2642 = ~pi46 & n2641;
  assign n2643 = ~pi46 & n2639;
  assign n2644 = ~pi46 & n2640;
  assign n2645 = ~pi94 & n2643;
  assign n2646 = n2641 & n62350;
  assign n2647 = n2641 & n2643;
  assign n2648 = ~pi94 & n2647;
  assign n2649 = n2640 & n2642;
  assign n2650 = ~pi46 & n2638;
  assign n2651 = n2640 & n2650;
  assign n2652 = n2638 & n62350;
  assign n2653 = n2641 & n62352;
  assign n2654 = n2638 & n62351;
  assign n2655 = ~pi47 & n62353;
  assign n2656 = ~pi91 & n2655;
  assign n2657 = n2636 & n62353;
  assign n2658 = n62349 & n62354;
  assign n2659 = n2586 & n2658;
  assign n2660 = ~pi841 & n2659;
  assign n2661 = pi93 & ~n2660;
  assign n2662 = n2585 & ~n2661;
  assign n2663 = ~pi58 & ~pi91;
  assign n2664 = ~pi47 & n2663;
  assign n2665 = n2641 & n2664;
  assign n2666 = n62351 & n2664;
  assign n2667 = n62350 & n2665;
  assign n2668 = n62352 & n2665;
  assign n2669 = n2638 & n62355;
  assign n2670 = n2627 & n62356;
  assign n2671 = n62349 & n62352;
  assign n2672 = n2665 & n2671;
  assign n2673 = n2630 & n2670;
  assign n2674 = ~pi841 & n62357;
  assign n2675 = pi90 & n2674;
  assign n2676 = ~pi93 & ~n2675;
  assign n2677 = n2662 & ~n2676;
  assign n2678 = ~pi51 & ~n2677;
  assign n2679 = ~pi102 & n2633;
  assign n2680 = n2614 & n2632;
  assign n2681 = ~pi88 & pi98;
  assign n2682 = ~pi86 & ~pi94;
  assign n2683 = ~pi50 & n2637;
  assign n2684 = ~pi77 & n2683;
  assign n2685 = n2682 & n2684;
  assign n2686 = n2681 & n2685;
  assign n2687 = ~pi50 & ~pi77;
  assign n2688 = ~pi94 & n2687;
  assign n2689 = n62358 & n2688;
  assign n2690 = n2638 & n2681;
  assign n2691 = n2689 & n2690;
  assign n2692 = n62358 & n2686;
  assign n2693 = ~pi97 & ~n62359;
  assign n2694 = ~pi90 & ~pi93;
  assign n2695 = ~pi35 & n2694;
  assign n2696 = ~pi70 & n2695;
  assign n2697 = n2636 & n2641;
  assign n2698 = ~pi109 & n2643;
  assign n2699 = ~pi110 & n2636;
  assign n2700 = n2698 & n2699;
  assign n2701 = n2636 & n2647;
  assign n2702 = n2636 & n2639;
  assign n2703 = n2642 & n2702;
  assign n2704 = n2643 & n2697;
  assign n2705 = ~pi58 & n62360;
  assign n2706 = n2643 & n2665;
  assign n2707 = n2696 & n62361;
  assign n2708 = ~n2693 & n62361;
  assign n2709 = n2696 & n2708;
  assign n2710 = ~pi90 & n62361;
  assign n2711 = n62359 & n2710;
  assign n2712 = n2662 & n2711;
  assign n2713 = ~n2693 & n2707;
  assign n2714 = n2678 & ~n62362;
  assign n2715 = ~pi93 & n2586;
  assign n2716 = n62354 & n2715;
  assign n2717 = ~pi93 & n2659;
  assign n2718 = n62349 & n2716;
  assign n2719 = ~pi35 & ~pi93;
  assign n2720 = n2586 & n2719;
  assign n2721 = n2659 & n2719;
  assign n2722 = n2658 & n2720;
  assign n2723 = ~pi70 & n62364;
  assign n2724 = n2585 & n62363;
  assign n2725 = pi51 & ~n62365;
  assign n2726 = ~pi40 & ~pi72;
  assign n2727 = ~pi32 & ~pi95;
  assign n2728 = n2726 & n2727;
  assign n2729 = ~pi72 & ~pi96;
  assign n2730 = ~pi40 & n2729;
  assign n2731 = n2727 & n2730;
  assign n2732 = ~pi96 & n2728;
  assign n2733 = ~pi96 & ~n2725;
  assign n2734 = n2728 & n2733;
  assign n2735 = ~n2725 & n62366;
  assign n2736 = ~n2714 & ~n2725;
  assign n2737 = n62366 & n2736;
  assign n2738 = ~n2714 & n62367;
  assign n2739 = n2584 & n62368;
  assign n2740 = ~n2581 & n2739;
  assign n2741 = ~pi96 & ~n2736;
  assign n2742 = n2581 & n2582;
  assign n2743 = ~pi51 & n2585;
  assign n2744 = ~pi93 & n2660;
  assign n2745 = ~pi841 & n62363;
  assign n2746 = n2743 & n62369;
  assign n2747 = pi96 & ~n2746;
  assign n2748 = n2726 & ~n2747;
  assign n2749 = n2727 & n2748;
  assign n2750 = ~pi32 & ~pi40;
  assign n2751 = ~pi95 & n2750;
  assign n2752 = ~n2747 & n2751;
  assign n2753 = ~pi72 & n2752;
  assign n2754 = n2728 & ~n2747;
  assign n2755 = ~pi72 & n2742;
  assign n2756 = n2752 & n2755;
  assign n2757 = n2742 & n62370;
  assign n2758 = ~n2741 & n2752;
  assign n2759 = n2755 & n2758;
  assign n2760 = ~n2741 & n62371;
  assign n2761 = ~n2740 & ~n62372;
  assign n2762 = ~pi1093 & ~n2761;
  assign n2763 = ~pi87 & ~n2762;
  assign n2764 = ~pi38 & ~pi39;
  assign n2765 = ~pi75 & ~pi100;
  assign n2766 = ~pi38 & ~pi100;
  assign n2767 = ~pi100 & n2764;
  assign n2768 = ~pi39 & n2766;
  assign n2769 = ~pi75 & n62373;
  assign n2770 = n2764 & n2765;
  assign n2771 = ~pi70 & ~pi96;
  assign n2772 = ~pi51 & ~pi72;
  assign n2773 = ~pi51 & ~pi70;
  assign n2774 = n2729 & n2773;
  assign n2775 = n2771 & n2772;
  assign n2776 = n2730 & n2773;
  assign n2777 = ~pi40 & n62375;
  assign n2778 = n2727 & n62376;
  assign n2779 = ~pi70 & n62366;
  assign n2780 = n2728 & n2771;
  assign n2781 = ~pi51 & n62378;
  assign n2782 = n2751 & n62375;
  assign n2783 = n2715 & n2743;
  assign n2784 = n62366 & n2783;
  assign n2785 = n2720 & n62377;
  assign n2786 = n62364 & n62377;
  assign n2787 = ~pi51 & ~pi96;
  assign n2788 = ~pi51 & n62366;
  assign n2789 = n2728 & n2787;
  assign n2790 = n62365 & n62381;
  assign n2791 = n2729 & n2743;
  assign n2792 = ~pi35 & n62375;
  assign n2793 = n62364 & n62375;
  assign n2794 = n62363 & n62382;
  assign n2795 = n2750 & n62383;
  assign n2796 = ~pi95 & n2795;
  assign n2797 = n2658 & n62379;
  assign po740 = ~pi1093 & n2584;
  assign n2799 = n62380 & po740;
  assign n2800 = pi87 & ~n2799;
  assign n2801 = n62374 & ~n2800;
  assign n2802 = ~n2763 & n2801;
  assign n2803 = ~pi567 & ~n2802;
  assign n2804 = n2580 & ~n2803;
  assign n2805 = ~pi39 & ~pi87;
  assign n2806 = n2766 & n2805;
  assign n2807 = ~pi144 & ~pi174;
  assign n2808 = ~pi189 & n2807;
  assign n2809 = ~pi299 & ~n2808;
  assign n2810 = ~pi152 & ~pi161;
  assign n2811 = ~pi166 & n2810;
  assign n2812 = pi299 & ~n2811;
  assign n2813 = ~n2809 & ~n2812;
  assign n2814 = ~pi332 & ~pi468;
  assign n2815 = pi232 & n2814;
  assign n2816 = n2813 & n2815;
  assign n2817 = n2806 & ~n2816;
  assign n2818 = ~pi24 & n62364;
  assign n2819 = n62377 & n2818;
  assign n2820 = ~pi24 & n62380;
  assign n2821 = pi252 & n62380;
  assign n2822 = ~pi24 & n2821;
  assign n2823 = pi252 & n62384;
  assign n2824 = ~pi833 & pi957;
  assign n2825 = ~pi41 & ~pi99;
  assign n2826 = ~pi101 & n2825;
  assign n2827 = ~pi113 & ~pi116;
  assign n2828 = ~pi52 & n2827;
  assign n2829 = ~pi114 & ~pi115;
  assign n2830 = ~pi42 & ~pi43;
  assign n2831 = ~pi42 & ~pi114;
  assign n2832 = ~pi42 & n2829;
  assign n2833 = ~pi115 & n2831;
  assign n2834 = ~pi43 & n62386;
  assign n2835 = ~pi114 & n2830;
  assign n2836 = ~pi115 & n2835;
  assign n2837 = n2829 & n2830;
  assign n2838 = ~pi52 & n2830;
  assign n2839 = n2827 & n2829;
  assign n2840 = n2838 & n2839;
  assign n2841 = n2828 & n62387;
  assign n2842 = n2826 & n62388;
  assign n2843 = ~pi44 & n2842;
  assign n2844 = ~n2824 & ~n2843;
  assign n2845 = pi1091 & n2844;
  assign n2846 = n2742 & n2845;
  assign n2847 = n62385 & n2846;
  assign n2848 = pi1093 & n2847;
  assign n2849 = n2817 & n2848;
  assign n2850 = pi75 & ~n2849;
  assign n2851 = pi1093 & ~n2824;
  assign n2852 = pi824 & n2582;
  assign n2853 = ~n2678 & n62367;
  assign n2854 = n2852 & n2853;
  assign n2855 = ~pi829 & n2854;
  assign n2856 = n62349 & n2655;
  assign n2857 = pi91 & n2856;
  assign n2858 = ~pi24 & n2857;
  assign n2859 = n2611 & n62358;
  assign n2860 = n2612 & n62358;
  assign n2861 = n2683 & n2860;
  assign n2862 = n2682 & n2861;
  assign n2863 = n2685 & n2859;
  assign n2864 = ~pi91 & pi97;
  assign n2865 = ~pi108 & n2864;
  assign n2866 = ~pi47 & ~pi110;
  assign n2867 = ~pi46 & ~pi109;
  assign n2868 = n2866 & n2867;
  assign n2869 = n2865 & n2868;
  assign n2870 = ~pi47 & n2641;
  assign n2871 = ~pi46 & pi97;
  assign n2872 = ~pi108 & n2871;
  assign n2873 = n2870 & n2872;
  assign n2874 = n62389 & n2873;
  assign n2875 = ~pi91 & n2874;
  assign n2876 = n62389 & n2869;
  assign n2877 = ~n2858 & ~n62390;
  assign n2878 = n2586 & n2662;
  assign n2879 = ~n2877 & n2878;
  assign n2880 = n2678 & ~n2879;
  assign n2881 = ~n2725 & ~n2880;
  assign n2882 = ~pi96 & ~n2881;
  assign n2883 = pi829 & n2582;
  assign n2884 = ~pi72 & pi950;
  assign n2885 = n2752 & n2884;
  assign n2886 = pi950 & n62370;
  assign n2887 = pi829 & pi1092;
  assign n2888 = n62391 & n2887;
  assign n2889 = n62370 & n2883;
  assign n2890 = ~n2882 & n62392;
  assign n2891 = ~n2855 & ~n2890;
  assign n2892 = ~pi122 & ~n2891;
  assign n2893 = pi122 & n2584;
  assign n2894 = n2853 & n2893;
  assign n2895 = ~n2892 & ~n2894;
  assign n2896 = n2851 & ~n2895;
  assign n2897 = pi1091 & ~n2896;
  assign n2898 = ~n2762 & n2897;
  assign n2899 = ~pi1091 & ~n2762;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = ~pi39 & ~n2900;
  assign n2902 = pi603 & ~pi642;
  assign n2903 = ~pi614 & ~pi616;
  assign n2904 = n2902 & n2903;
  assign n2905 = ~pi662 & pi680;
  assign n2906 = ~pi661 & n2905;
  assign n2907 = ~pi681 & n2906;
  assign n2908 = ~n2904 & ~n2907;
  assign n2909 = ~n2814 & ~n2908;
  assign n2910 = ~pi960 & ~pi963;
  assign n2911 = ~pi970 & ~pi972;
  assign n2912 = ~pi975 & ~pi978;
  assign n2913 = n2911 & n2912;
  assign n2914 = n2910 & n2913;
  assign n2915 = ~pi907 & ~pi947;
  assign n2916 = ~pi907 & n2914;
  assign n2917 = ~pi947 & n2916;
  assign n2918 = n2914 & n2915;
  assign n2919 = n2814 & ~n62393;
  assign n2920 = ~n2909 & ~n2919;
  assign n2921 = pi829 & pi950;
  assign n2922 = ~n2824 & n2921;
  assign n2923 = pi1092 & pi1093;
  assign n2924 = pi1091 & pi1093;
  assign n2925 = pi1092 & n2924;
  assign n2926 = pi1091 & n2923;
  assign n2927 = ~n2824 & n2924;
  assign n2928 = n2883 & n2927;
  assign n2929 = pi1091 & ~n2824;
  assign n2930 = n2921 & n2923;
  assign n2931 = n2929 & n2930;
  assign n2932 = n2922 & n62394;
  assign n2933 = ~pi287 & n62380;
  assign n2934 = pi835 & pi984;
  assign n2935 = ~pi252 & ~pi1001;
  assign n2936 = ~pi979 & ~n2935;
  assign n2937 = ~n2934 & n2936;
  assign n2938 = pi835 & n2937;
  assign n2939 = n2933 & n2938;
  assign n2940 = n2921 & n2939;
  assign n2941 = pi1092 & n2940;
  assign n2942 = n2883 & n2939;
  assign n2943 = n2927 & n62396;
  assign n2944 = ~n2824 & n2940;
  assign n2945 = n2922 & n2939;
  assign n2946 = n2923 & n62398;
  assign n2947 = n2851 & n62396;
  assign n2948 = pi1091 & n62399;
  assign n2949 = n62395 & n2939;
  assign n2950 = n2909 & n62397;
  assign n2951 = n62393 & ~n2950;
  assign n2952 = ~n2814 & ~n2904;
  assign n2953 = ~n2907 & n2952;
  assign n2954 = n62397 & ~n2953;
  assign n2955 = ~n62393 & ~n2954;
  assign n2956 = ~n2951 & ~n2955;
  assign n2957 = ~n2920 & n62397;
  assign n2958 = ~pi216 & pi221;
  assign n2959 = ~pi215 & pi299;
  assign n2960 = ~pi215 & pi221;
  assign n2961 = pi299 & n2960;
  assign n2962 = ~pi216 & n2961;
  assign n2963 = n2958 & n2959;
  assign n2964 = n62400 & n62401;
  assign n2965 = ~pi969 & ~pi971;
  assign n2966 = ~pi974 & ~pi977;
  assign n2967 = n2965 & n2966;
  assign n2968 = ~pi587 & ~pi602;
  assign n2969 = ~pi961 & ~pi967;
  assign n2970 = n2968 & n2969;
  assign n2971 = n2967 & n2970;
  assign n2972 = n2814 & ~n2971;
  assign n2973 = ~n2909 & ~n2972;
  assign n2974 = ~n2950 & n2971;
  assign n2975 = ~n2954 & ~n2971;
  assign n2976 = ~n2974 & ~n2975;
  assign n2977 = n62397 & ~n2973;
  assign n2978 = pi222 & ~pi224;
  assign n2979 = ~pi223 & ~pi299;
  assign n2980 = pi222 & ~pi223;
  assign n2981 = ~pi299 & n2980;
  assign n2982 = pi222 & n2979;
  assign n2983 = ~pi224 & n62403;
  assign n2984 = n2978 & n2979;
  assign n2985 = n62402 & n62404;
  assign n2986 = pi39 & ~n2985;
  assign n2987 = pi39 & ~n2964;
  assign n2988 = ~n2985 & n2987;
  assign n2989 = ~n2964 & n2986;
  assign n2990 = ~pi38 & ~n62405;
  assign n2991 = ~n2901 & n2990;
  assign n2992 = ~pi100 & ~n2991;
  assign n2993 = pi1093 & n2742;
  assign n2994 = n2844 & n2993;
  assign n2995 = n62380 & n2994;
  assign n2996 = pi1091 & n2995;
  assign n2997 = pi228 & ~n2816;
  assign n2998 = n2764 & n2997;
  assign n2999 = pi228 & n2996;
  assign n3000 = n2764 & ~n2816;
  assign n3001 = n2999 & n3000;
  assign n3002 = n2996 & n2998;
  assign n3003 = pi100 & ~n62406;
  assign n3004 = ~pi87 & ~n3003;
  assign n3005 = ~n2992 & n3004;
  assign n3006 = ~pi1091 & ~n2799;
  assign n3007 = pi1093 & n2824;
  assign n3008 = n2584 & ~n3007;
  assign n3009 = n62380 & n3008;
  assign n3010 = pi1091 & ~n3009;
  assign n3011 = pi87 & ~pi100;
  assign n3012 = pi87 & n62373;
  assign n3013 = n2764 & n3011;
  assign n3014 = ~n3010 & n62407;
  assign n3015 = ~n3006 & n62407;
  assign n3016 = ~n3010 & n3015;
  assign n3017 = ~n3006 & n3014;
  assign n3018 = ~pi75 & ~n62408;
  assign n3019 = ~n3005 & n3018;
  assign n3020 = ~n2850 & ~n3019;
  assign n3021 = pi567 & ~n3020;
  assign n3022 = n2804 & ~n3021;
  assign n3023 = ~pi592 & ~n3022;
  assign n3024 = n62385 & n2994;
  assign n3025 = pi1091 & ~n3024;
  assign n3026 = n2817 & ~n3025;
  assign n3027 = ~pi98 & n2852;
  assign n3028 = ~pi122 & pi1093;
  assign n3029 = n3027 & n3028;
  assign n3030 = ~pi1091 & ~n3029;
  assign n3031 = n3026 & ~n3030;
  assign n3032 = ~pi1091 & pi1093;
  assign n3033 = ~pi122 & n3027;
  assign n3034 = ~pi1091 & n3029;
  assign n3035 = n2852 & n3028;
  assign n3036 = ~pi1091 & n3035;
  assign n3037 = ~pi98 & n3036;
  assign n3038 = n3032 & n3033;
  assign n3039 = ~n2817 & n62409;
  assign n3040 = pi75 & ~n3039;
  assign n3041 = ~n3031 & n3040;
  assign n3042 = ~pi39 & ~n2898;
  assign n3043 = pi122 & n2854;
  assign n3044 = ~n3033 & ~n3043;
  assign n3045 = pi1093 & ~n3044;
  assign n3046 = n2899 & ~n3045;
  assign n3047 = n3042 & ~n3046;
  assign n3048 = pi1091 & ~n62399;
  assign n3049 = ~n3030 & ~n3048;
  assign n3050 = pi1091 & n2953;
  assign n3051 = ~n2953 & n3049;
  assign n3052 = n2953 & n62409;
  assign n3053 = ~n3051 & ~n3052;
  assign n3054 = n3049 & ~n3050;
  assign n3055 = ~n62393 & n62410;
  assign n3056 = ~pi216 & n2960;
  assign n3057 = pi1091 & ~n2909;
  assign n3058 = ~n2909 & ~n62409;
  assign n3059 = n2909 & ~n3049;
  assign n3060 = ~n3058 & ~n3059;
  assign n3061 = n2909 & n3049;
  assign n3062 = ~n2909 & n62409;
  assign n3063 = ~n3061 & ~n3062;
  assign n3064 = n3049 & ~n3057;
  assign n3065 = n62393 & ~n62411;
  assign n3066 = n3056 & ~n3065;
  assign n3067 = ~n3055 & n3056;
  assign n3068 = ~n3065 & n3067;
  assign n3069 = ~n3055 & n3066;
  assign n3070 = n3036 & ~n3056;
  assign n3071 = ~pi98 & n3070;
  assign n3072 = n62409 & ~n3056;
  assign n3073 = pi299 & ~n62413;
  assign n3074 = ~n62412 & n3073;
  assign n3075 = n2971 & ~n62411;
  assign n3076 = ~pi223 & n2978;
  assign n3077 = ~n2971 & n62410;
  assign n3078 = n3076 & ~n3077;
  assign n3079 = ~n3075 & n3076;
  assign n3080 = ~n3077 & n3079;
  assign n3081 = ~n3075 & n3078;
  assign n3082 = n3036 & ~n3076;
  assign n3083 = ~pi98 & n3082;
  assign n3084 = n62409 & ~n3076;
  assign n3085 = ~pi299 & ~n62415;
  assign n3086 = ~n62414 & n3085;
  assign n3087 = pi39 & ~n3086;
  assign n3088 = pi39 & ~n3074;
  assign n3089 = ~n3086 & n3088;
  assign n3090 = ~n3074 & n3087;
  assign n3091 = ~n3047 & ~n62416;
  assign n3092 = ~pi38 & ~n3091;
  assign n3093 = pi38 & n3036;
  assign n3094 = ~pi98 & n3093;
  assign n3095 = pi38 & n62409;
  assign n3096 = ~pi100 & ~n62417;
  assign n3097 = ~n3092 & n3096;
  assign n3098 = n2997 & ~n62409;
  assign n3099 = pi1091 & ~n2995;
  assign n3100 = ~n3030 & ~n3099;
  assign n3101 = n2997 & ~n3100;
  assign n3102 = ~n2996 & n3098;
  assign n3103 = ~n2997 & ~n62409;
  assign n3104 = n2764 & ~n3103;
  assign n3105 = ~n62418 & n3104;
  assign n3106 = ~n2764 & n62409;
  assign n3107 = pi100 & ~n3106;
  assign n3108 = ~n3105 & n3107;
  assign n3109 = n3003 & ~n62409;
  assign n3110 = ~pi87 & ~n62419;
  assign n3111 = ~n3097 & n3110;
  assign n3112 = pi824 & pi950;
  assign n3113 = pi950 & n62380;
  assign n3114 = pi824 & n3113;
  assign n3115 = n62380 & n3112;
  assign n3116 = pi1092 & n62420;
  assign n3117 = n62380 & n2852;
  assign n3118 = pi122 & n62421;
  assign n3119 = ~n3033 & ~n3118;
  assign n3120 = pi1093 & ~n3119;
  assign n3121 = n3006 & ~n3120;
  assign n3122 = n62373 & ~n3010;
  assign n3123 = ~n3121 & n3122;
  assign n3124 = ~n62409 & ~n3123;
  assign n3125 = pi87 & ~n3124;
  assign n3126 = ~pi75 & ~n3125;
  assign n3127 = ~n3111 & n3126;
  assign n3128 = ~n3041 & ~n3127;
  assign n3129 = pi567 & ~n3128;
  assign n3130 = n2804 & ~n3129;
  assign n3131 = pi567 & ~n2580;
  assign n3132 = pi567 & n62409;
  assign n3133 = ~n2580 & n3132;
  assign n3134 = n62409 & n3131;
  assign n3135 = ~n3130 & ~n62422;
  assign n3136 = pi592 & n3135;
  assign n3137 = ~n3023 & ~n3136;
  assign n3138 = ~n2578 & ~n3137;
  assign n3139 = pi443 & ~pi592;
  assign n3140 = n3135 & ~n3139;
  assign n3141 = pi434 & ~pi446;
  assign n3142 = ~pi434 & pi446;
  assign n3143 = ~pi434 & ~pi446;
  assign n3144 = pi434 & pi446;
  assign n3145 = ~n3143 & ~n3144;
  assign n3146 = ~n3141 & ~n3142;
  assign n3147 = ~pi414 & ~pi435;
  assign n3148 = pi414 & pi435;
  assign n3149 = pi414 & ~pi435;
  assign n3150 = ~pi414 & pi435;
  assign n3151 = ~n3149 & ~n3150;
  assign n3152 = ~n3147 & ~n3148;
  assign n3153 = ~pi422 & ~pi429;
  assign n3154 = pi422 & pi429;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = ~n62424 & ~n3155;
  assign n3157 = n62424 & n3155;
  assign n3158 = ~n3156 & ~n3157;
  assign n3159 = ~n62423 & n3158;
  assign n3160 = n62423 & ~n3158;
  assign n3161 = n62423 & ~n3155;
  assign n3162 = ~n62423 & n3155;
  assign n3163 = ~n3161 & ~n3162;
  assign n3164 = n62424 & n3163;
  assign n3165 = ~n62424 & ~n3163;
  assign n3166 = ~n3164 & ~n3165;
  assign n3167 = pi414 & ~pi422;
  assign n3168 = ~pi414 & pi422;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = ~n62423 & n3169;
  assign n3171 = n62423 & ~n3169;
  assign n3172 = ~n3170 & ~n3171;
  assign n3173 = pi429 & ~n3172;
  assign n3174 = ~pi429 & n3172;
  assign n3175 = ~n3173 & ~n3174;
  assign n3176 = pi435 & n3175;
  assign n3177 = ~pi435 & ~n3175;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = ~pi429 & ~pi435;
  assign n3180 = pi429 & pi435;
  assign n3181 = ~n3179 & ~n3180;
  assign n3182 = n3172 & n3181;
  assign n3183 = ~n3172 & ~n3181;
  assign n3184 = ~n3182 & ~n3183;
  assign n3185 = ~n3159 & ~n3160;
  assign n3186 = pi436 & ~pi444;
  assign n3187 = ~pi436 & pi444;
  assign n3188 = ~n3186 & ~n3187;
  assign n3189 = n62425 & n3188;
  assign n3190 = ~n62425 & ~n3188;
  assign n3191 = n62425 & ~n3188;
  assign n3192 = ~n62425 & n3188;
  assign n3193 = ~n3191 & ~n3192;
  assign n3194 = ~n3189 & ~n3190;
  assign n3195 = ~n3022 & n3139;
  assign n3196 = ~n62426 & ~n3195;
  assign n3197 = ~n3140 & n3196;
  assign n3198 = ~pi443 & ~pi592;
  assign n3199 = n3135 & ~n3198;
  assign n3200 = ~n3022 & n3198;
  assign n3201 = n62426 & ~n3200;
  assign n3202 = ~n3199 & n3201;
  assign n3203 = ~n3197 & ~n3202;
  assign n3204 = pi1196 & ~n3203;
  assign n3205 = ~pi1196 & ~n3135;
  assign n3206 = n2578 & ~n3205;
  assign n3207 = ~pi1196 & n3135;
  assign n3208 = pi1196 & ~n3202;
  assign n3209 = pi1196 & ~n3197;
  assign n3210 = ~n3202 & n3209;
  assign n3211 = ~n3197 & n3208;
  assign n3212 = ~n3207 & ~n62427;
  assign n3213 = n2578 & ~n3212;
  assign n3214 = ~n3204 & n3206;
  assign n3215 = ~n3138 & ~n62428;
  assign n3216 = ~n62332 & ~n3215;
  assign n3217 = n62332 & ~n3137;
  assign n3218 = ~n62332 & n3215;
  assign n3219 = n62332 & n3137;
  assign n3220 = ~n3218 & ~n3219;
  assign n3221 = pi428 & n3215;
  assign n3222 = ~pi428 & n3137;
  assign n3223 = pi427 & ~n3222;
  assign n3224 = ~n3221 & n3223;
  assign n3225 = ~pi428 & n3215;
  assign n3226 = pi428 & n3137;
  assign n3227 = ~pi427 & ~n3226;
  assign n3228 = ~n3225 & n3227;
  assign n3229 = ~n3224 & ~n3228;
  assign n3230 = ~n3216 & ~n3217;
  assign n3231 = n62331 & ~n62429;
  assign n3232 = ~n62332 & n3137;
  assign n3233 = n62332 & n3215;
  assign n3234 = n62332 & ~n3215;
  assign n3235 = ~n62332 & ~n3137;
  assign n3236 = ~n3234 & ~n3235;
  assign n3237 = ~n3232 & ~n3233;
  assign n3238 = ~n62331 & n62430;
  assign n3239 = pi430 & n62429;
  assign n3240 = ~pi430 & ~n62430;
  assign n3241 = ~pi430 & n62430;
  assign n3242 = pi430 & ~n62429;
  assign n3243 = ~n3241 & ~n3242;
  assign n3244 = ~n3239 & ~n3240;
  assign n3245 = pi426 & ~n62431;
  assign n3246 = ~pi430 & n62429;
  assign n3247 = pi430 & ~n62430;
  assign n3248 = pi430 & n62430;
  assign n3249 = ~pi430 & ~n62429;
  assign n3250 = ~n3248 & ~n3249;
  assign n3251 = ~n3246 & ~n3247;
  assign n3252 = ~pi426 & ~n3247;
  assign n3253 = ~n3246 & n3252;
  assign n3254 = ~pi426 & ~n62432;
  assign n3255 = ~n3245 & ~n62433;
  assign n3256 = ~pi426 & n62432;
  assign n3257 = pi426 & n62431;
  assign n3258 = ~n3256 & ~n3257;
  assign n3259 = ~n3231 & ~n3238;
  assign n3260 = pi445 & n62434;
  assign n3261 = pi433 & ~pi451;
  assign n3262 = ~pi433 & pi451;
  assign n3263 = ~pi433 & ~pi451;
  assign n3264 = pi433 & pi451;
  assign n3265 = ~n3263 & ~n3264;
  assign n3266 = ~n3261 & ~n3262;
  assign n3267 = pi449 & ~n62435;
  assign n3268 = ~pi449 & n62435;
  assign n3269 = ~n3267 & ~n3268;
  assign n3270 = pi448 & n3269;
  assign n3271 = ~pi448 & ~n3269;
  assign n3272 = pi448 & ~n3269;
  assign n3273 = ~pi448 & n3269;
  assign n3274 = ~n3272 & ~n3273;
  assign n3275 = ~n3270 & ~n3271;
  assign n3276 = n62331 & n62430;
  assign n3277 = ~n62331 & ~n62429;
  assign n3278 = pi426 & ~n62432;
  assign n3279 = ~pi426 & ~n62431;
  assign n3280 = ~n3278 & ~n3279;
  assign n3281 = ~pi426 & n62431;
  assign n3282 = pi426 & n62432;
  assign n3283 = ~n3281 & ~n3282;
  assign n3284 = ~n3276 & ~n3277;
  assign n3285 = ~pi445 & n62437;
  assign n3286 = n62436 & ~n3285;
  assign n3287 = ~n3260 & n3286;
  assign n3288 = pi445 & n62437;
  assign n3289 = ~pi445 & n62434;
  assign n3290 = ~n62436 & ~n3289;
  assign n3291 = ~n62436 & ~n3288;
  assign n3292 = ~n3289 & n3291;
  assign n3293 = ~n3288 & n3290;
  assign n3294 = pi1199 & ~n62438;
  assign n3295 = ~n3288 & ~n3289;
  assign n3296 = pi448 & n3295;
  assign n3297 = ~n3260 & ~n3285;
  assign n3298 = ~pi448 & n3297;
  assign n3299 = ~n3269 & ~n3298;
  assign n3300 = ~n3269 & ~n3296;
  assign n3301 = ~n3298 & n3300;
  assign n3302 = ~n3296 & n3299;
  assign n3303 = ~pi448 & n3295;
  assign n3304 = pi448 & n3297;
  assign n3305 = n3269 & ~n3304;
  assign n3306 = n3269 & ~n3303;
  assign n3307 = ~n3304 & n3306;
  assign n3308 = ~n3303 & n3305;
  assign n3309 = ~n62439 & ~n62440;
  assign n3310 = pi1199 & ~n3309;
  assign n3311 = ~n3287 & n3294;
  assign n3312 = ~pi590 & ~pi591;
  assign n3313 = ~pi1199 & ~n3215;
  assign n3314 = n3312 & ~n3313;
  assign n3315 = ~n62441 & n3314;
  assign n3316 = ~pi285 & ~pi286;
  assign n3317 = ~pi289 & n3316;
  assign n3318 = ~pi288 & n3317;
  assign n3319 = ~n3135 & ~n3312;
  assign n3320 = ~n3318 & ~n3319;
  assign n3321 = ~n3315 & n3320;
  assign n3322 = pi824 & pi1093;
  assign n3323 = pi1093 & n2852;
  assign n3324 = n2582 & n3322;
  assign n3325 = pi1093 & n2854;
  assign n3326 = n2853 & n62442;
  assign n3327 = n2990 & n62443;
  assign n3328 = ~n2897 & n3327;
  assign n3329 = n2992 & ~n3328;
  assign n3330 = ~n3003 & ~n3329;
  assign n3331 = ~pi87 & ~n3330;
  assign n3332 = n3032 & ~n62421;
  assign n3333 = ~n3009 & ~n3032;
  assign n3334 = n62373 & ~n3333;
  assign n3335 = ~n3332 & n3334;
  assign n3336 = pi87 & ~n3335;
  assign n3337 = ~n3331 & ~n3336;
  assign n3338 = ~pi75 & ~n3337;
  assign n3339 = ~n2850 & ~n3338;
  assign n3340 = pi567 & ~n3339;
  assign n3341 = n2804 & ~n3340;
  assign n3342 = pi592 & ~n3341;
  assign n3343 = ~n3023 & ~n3342;
  assign n3344 = ~n2578 & n3343;
  assign n3345 = ~pi443 & ~n3341;
  assign n3346 = ~n3195 & ~n3345;
  assign n3347 = ~n62426 & ~n3346;
  assign n3348 = pi443 & ~n3341;
  assign n3349 = ~n3200 & ~n3348;
  assign n3350 = n62426 & ~n3349;
  assign n3351 = ~n3342 & ~n3350;
  assign n3352 = ~n3347 & n3351;
  assign n3353 = ~n3139 & ~n3341;
  assign n3354 = ~n3195 & ~n3353;
  assign n3355 = ~pi444 & ~n3354;
  assign n3356 = ~n3198 & ~n3341;
  assign n3357 = ~n3200 & ~n3356;
  assign n3358 = pi444 & ~n3357;
  assign n3359 = ~n3355 & ~n3358;
  assign n3360 = ~pi436 & ~n3359;
  assign n3361 = ~pi444 & ~n3357;
  assign n3362 = pi444 & ~n3354;
  assign n3363 = ~n3361 & ~n3362;
  assign n3364 = pi436 & ~n3363;
  assign n3365 = ~n62425 & ~n3364;
  assign n3366 = ~n62425 & ~n3360;
  assign n3367 = ~n3364 & n3366;
  assign n3368 = ~n3360 & n3365;
  assign n3369 = ~pi436 & ~n3363;
  assign n3370 = pi436 & ~n3359;
  assign n3371 = n62425 & ~n3370;
  assign n3372 = n62425 & ~n3369;
  assign n3373 = ~n3370 & n3372;
  assign n3374 = ~n3369 & n3371;
  assign n3375 = pi1196 & ~n62445;
  assign n3376 = ~n62444 & n3375;
  assign n3377 = pi1196 & ~n62444;
  assign n3378 = ~n62445 & n3377;
  assign n3379 = pi1196 & ~n3352;
  assign n3380 = ~pi1196 & ~n3341;
  assign n3381 = n2578 & ~n3380;
  assign n3382 = ~n62446 & n3381;
  assign n3383 = ~n62446 & ~n3380;
  assign n3384 = n2578 & ~n3383;
  assign n3385 = ~n2578 & ~n3343;
  assign n3386 = ~n3384 & ~n3385;
  assign n3387 = ~n3344 & ~n3382;
  assign n3388 = pi428 & n62447;
  assign n3389 = ~pi428 & n3343;
  assign n3390 = pi427 & ~n3389;
  assign n3391 = ~n3388 & n3390;
  assign n3392 = ~pi428 & n62447;
  assign n3393 = pi428 & n3343;
  assign n3394 = ~pi427 & ~n3393;
  assign n3395 = ~n3392 & n3394;
  assign n3396 = pi428 & ~n3343;
  assign n3397 = ~pi428 & ~n62447;
  assign n3398 = ~n3396 & ~n3397;
  assign n3399 = ~n3392 & ~n3393;
  assign n3400 = ~pi427 & n62448;
  assign n3401 = ~n3388 & ~n3389;
  assign n3402 = pi427 & ~n3401;
  assign n3403 = ~n3400 & ~n3402;
  assign n3404 = ~n3391 & ~n3395;
  assign n3405 = n62331 & n62449;
  assign n3406 = pi445 & ~pi448;
  assign n3407 = ~pi445 & pi448;
  assign n3408 = ~pi445 & ~pi448;
  assign n3409 = pi445 & pi448;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = ~n3406 & ~n3407;
  assign n3412 = n3269 & ~n62450;
  assign n3413 = ~n3269 & n62450;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = ~n62332 & n3343;
  assign n3416 = n62332 & n62447;
  assign n3417 = ~pi427 & ~n3401;
  assign n3418 = pi427 & n62448;
  assign n3419 = ~n3417 & ~n3418;
  assign n3420 = ~n3415 & ~n3416;
  assign n3421 = ~n62331 & n62451;
  assign n3422 = ~n3414 & ~n3421;
  assign n3423 = ~n3405 & n3422;
  assign n3424 = ~n62331 & n62449;
  assign n3425 = n62331 & n62451;
  assign n3426 = n3414 & ~n3425;
  assign n3427 = ~n3424 & n3426;
  assign n3428 = pi1199 & ~n3427;
  assign n3429 = pi430 & ~n62449;
  assign n3430 = ~pi430 & ~n62451;
  assign n3431 = ~n3429 & ~n3430;
  assign n3432 = pi426 & ~n3431;
  assign n3433 = pi430 & ~n62451;
  assign n3434 = ~pi430 & ~n62449;
  assign n3435 = ~n3433 & ~n3434;
  assign n3436 = ~pi426 & ~n3435;
  assign n3437 = ~n3432 & ~n3436;
  assign n3438 = pi445 & ~n3437;
  assign n3439 = pi426 & ~n3435;
  assign n3440 = ~pi426 & ~n3431;
  assign n3441 = ~n3439 & ~n3440;
  assign n3442 = ~pi445 & ~n3441;
  assign n3443 = ~n3438 & ~n3442;
  assign n3444 = ~pi445 & n3441;
  assign n3445 = pi445 & n3437;
  assign n3446 = n62436 & ~n3445;
  assign n3447 = ~n3444 & n3446;
  assign n3448 = n62436 & ~n3443;
  assign n3449 = pi445 & ~n3441;
  assign n3450 = ~pi445 & ~n3437;
  assign n3451 = ~n3449 & ~n3450;
  assign n3452 = ~pi445 & n3437;
  assign n3453 = pi445 & n3441;
  assign n3454 = ~n62436 & ~n3453;
  assign n3455 = ~n3452 & n3454;
  assign n3456 = ~n62436 & ~n3451;
  assign n3457 = pi1199 & ~n62453;
  assign n3458 = ~n62452 & n3457;
  assign n3459 = pi1199 & ~n62452;
  assign n3460 = ~n62453 & n3459;
  assign n3461 = ~n3423 & n3428;
  assign n3462 = ~pi1199 & ~n62447;
  assign n3463 = n3312 & ~n3462;
  assign n3464 = ~n62454 & n3463;
  assign n3465 = ~n3312 & n3341;
  assign n3466 = n3318 & ~n3465;
  assign n3467 = ~n3464 & n3466;
  assign n3468 = ~n3321 & ~n3467;
  assign n3469 = pi588 & ~n3468;
  assign n3470 = ~pi56 & ~pi62;
  assign n3471 = ~pi55 & n3470;
  assign n3472 = ~pi57 & ~pi59;
  assign n3473 = n3470 & n3472;
  assign n3474 = ~pi55 & n3473;
  assign n3475 = ~pi59 & n3471;
  assign n3476 = ~pi57 & n3475;
  assign n3477 = n3471 & n3472;
  assign n3478 = ~pi351 & pi1199;
  assign n3479 = pi323 & ~pi450;
  assign n3480 = ~pi323 & pi450;
  assign n3481 = ~n3479 & ~n3480;
  assign n3482 = pi345 & ~pi346;
  assign n3483 = ~pi345 & pi346;
  assign n3484 = ~pi345 & ~pi346;
  assign n3485 = pi345 & pi346;
  assign n3486 = ~n3484 & ~n3485;
  assign n3487 = ~n3482 & ~n3483;
  assign n3488 = pi358 & n62456;
  assign n3489 = ~pi358 & ~n62456;
  assign n3490 = ~n3488 & ~n3489;
  assign n3491 = n3481 & n3490;
  assign n3492 = ~n3481 & ~n3490;
  assign n3493 = pi450 & n62456;
  assign n3494 = ~pi450 & ~n62456;
  assign n3495 = ~n3493 & ~n3494;
  assign n3496 = pi323 & ~pi358;
  assign n3497 = ~pi323 & pi358;
  assign n3498 = ~n3496 & ~n3497;
  assign n3499 = n3495 & n3498;
  assign n3500 = ~n3495 & ~n3498;
  assign n3501 = ~n3499 & ~n3500;
  assign n3502 = pi323 & n62456;
  assign n3503 = ~pi323 & ~n62456;
  assign n3504 = ~n3502 & ~n3503;
  assign n3505 = pi358 & ~n3504;
  assign n3506 = ~pi358 & n3504;
  assign n3507 = ~n3505 & ~n3506;
  assign n3508 = pi450 & n3507;
  assign n3509 = ~pi450 & ~n3507;
  assign n3510 = ~n3508 & ~n3509;
  assign n3511 = pi358 & ~pi450;
  assign n3512 = ~pi358 & pi450;
  assign n3513 = ~n3511 & ~n3512;
  assign n3514 = n3504 & ~n3513;
  assign n3515 = ~n3504 & n3513;
  assign n3516 = ~n3514 & ~n3515;
  assign n3517 = ~n3491 & ~n3492;
  assign n3518 = ~pi327 & ~pi362;
  assign n3519 = pi327 & pi362;
  assign n3520 = pi327 & ~pi362;
  assign n3521 = ~pi327 & pi362;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = ~n3518 & ~n3519;
  assign n3524 = pi343 & ~pi344;
  assign n3525 = ~pi343 & pi344;
  assign n3526 = ~n3524 & ~n3525;
  assign n3527 = ~n62458 & n3526;
  assign n3528 = n62458 & ~n3526;
  assign n3529 = pi343 & n62458;
  assign n3530 = ~pi343 & ~n62458;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = pi344 & n3531;
  assign n3533 = ~pi344 & ~n3531;
  assign n3534 = ~n3532 & ~n3533;
  assign n3535 = ~n62458 & ~n3526;
  assign n3536 = n62458 & n3526;
  assign n3537 = ~n3535 & ~n3536;
  assign n3538 = ~n3527 & ~n3528;
  assign n3539 = ~n62457 & ~n62459;
  assign n3540 = n62457 & n62459;
  assign n3541 = pi1197 & ~n3540;
  assign n3542 = pi1197 & ~n3539;
  assign n3543 = ~n3540 & n3542;
  assign n3544 = ~n3539 & n3541;
  assign n3545 = pi342 & ~pi361;
  assign n3546 = ~pi342 & pi361;
  assign n3547 = ~n3545 & ~n3546;
  assign n3548 = pi320 & ~pi460;
  assign n3549 = ~pi320 & pi460;
  assign n3550 = ~pi320 & ~pi460;
  assign n3551 = pi320 & pi460;
  assign n3552 = ~n3550 & ~n3551;
  assign n3553 = ~n3548 & ~n3549;
  assign n3554 = pi441 & n62461;
  assign n3555 = ~pi441 & ~n62461;
  assign n3556 = ~n3554 & ~n3555;
  assign n3557 = n3547 & n3556;
  assign n3558 = ~n3547 & ~n3556;
  assign n3559 = pi342 & n62461;
  assign n3560 = ~pi342 & ~n62461;
  assign n3561 = ~n3559 & ~n3560;
  assign n3562 = pi361 & ~pi441;
  assign n3563 = ~pi361 & pi441;
  assign n3564 = ~n3562 & ~n3563;
  assign n3565 = n3561 & n3564;
  assign n3566 = ~n3561 & ~n3564;
  assign n3567 = ~n3565 & ~n3566;
  assign n3568 = ~n3557 & ~n3558;
  assign n3569 = ~pi355 & ~pi458;
  assign n3570 = pi355 & pi458;
  assign n3571 = pi355 & ~pi458;
  assign n3572 = ~pi355 & pi458;
  assign n3573 = ~n3571 & ~n3572;
  assign n3574 = ~n3569 & ~n3570;
  assign n3575 = ~pi452 & ~pi455;
  assign n3576 = pi452 & pi455;
  assign n3577 = pi452 & ~pi455;
  assign n3578 = ~pi452 & pi455;
  assign n3579 = ~n3577 & ~n3578;
  assign n3580 = ~n3575 & ~n3576;
  assign n3581 = ~n62463 & n62464;
  assign n3582 = n62463 & ~n62464;
  assign n3583 = ~n3581 & ~n3582;
  assign n3584 = n62462 & n3583;
  assign n3585 = ~n62462 & ~n3583;
  assign n3586 = n62462 & n62463;
  assign n3587 = ~n62462 & ~n62463;
  assign n3588 = pi458 & n62462;
  assign n3589 = ~pi458 & ~n62462;
  assign n3590 = ~n3588 & ~n3589;
  assign n3591 = pi355 & ~n3590;
  assign n3592 = ~pi355 & n3590;
  assign n3593 = ~n3591 & ~n3592;
  assign n3594 = pi355 & ~n62462;
  assign n3595 = ~pi355 & n62462;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = pi458 & n3596;
  assign n3598 = ~pi458 & ~n3596;
  assign n3599 = ~n3597 & ~n3598;
  assign n3600 = ~n3586 & ~n3587;
  assign n3601 = ~n62464 & n62465;
  assign n3602 = n62464 & ~n62465;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = n62464 & n62465;
  assign n3605 = ~n62464 & ~n62465;
  assign n3606 = ~n3604 & ~n3605;
  assign n3607 = pi355 & n62464;
  assign n3608 = ~pi355 & ~n62464;
  assign n3609 = ~n3607 & ~n3608;
  assign n3610 = n3590 & n3609;
  assign n3611 = ~n3590 & ~n3609;
  assign n3612 = ~n3610 & ~n3611;
  assign n3613 = ~n3584 & ~n3585;
  assign n3614 = pi1196 & n62466;
  assign n3615 = ~n62460 & ~n3614;
  assign n3616 = ~n3137 & ~n3615;
  assign n3617 = pi316 & ~pi349;
  assign n3618 = ~pi316 & pi349;
  assign n3619 = ~pi316 & ~pi349;
  assign n3620 = pi316 & pi349;
  assign n3621 = ~n3619 & ~n3620;
  assign n3622 = ~n3617 & ~n3618;
  assign n3623 = ~pi315 & ~pi359;
  assign n3624 = pi315 & pi359;
  assign n3625 = pi315 & ~pi359;
  assign n3626 = ~pi315 & pi359;
  assign n3627 = ~n3625 & ~n3626;
  assign n3628 = ~n3623 & ~n3624;
  assign n3629 = pi321 & ~pi347;
  assign n3630 = ~pi321 & pi347;
  assign n3631 = ~pi321 & ~pi347;
  assign n3632 = pi321 & pi347;
  assign n3633 = ~n3631 & ~n3632;
  assign n3634 = ~n3629 & ~n3630;
  assign n3635 = pi322 & ~pi348;
  assign n3636 = ~pi322 & pi348;
  assign n3637 = ~n3635 & ~n3636;
  assign n3638 = ~n62469 & n3637;
  assign n3639 = n62469 & ~n3637;
  assign n3640 = ~n3638 & ~n3639;
  assign n3641 = ~n62468 & ~n3640;
  assign n3642 = n62468 & n3640;
  assign n3643 = ~n3641 & ~n3642;
  assign n3644 = ~n62467 & n3643;
  assign n3645 = n62467 & ~n3643;
  assign n3646 = ~n62467 & n3637;
  assign n3647 = n62467 & ~n3637;
  assign n3648 = ~n3646 & ~n3647;
  assign n3649 = ~n62469 & ~n3648;
  assign n3650 = n62469 & n3648;
  assign n3651 = pi348 & n62469;
  assign n3652 = ~pi348 & ~n62469;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = pi322 & n62467;
  assign n3655 = ~pi322 & ~n62467;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = n3653 & ~n3656;
  assign n3658 = ~n3653 & n3656;
  assign n3659 = ~n3657 & ~n3658;
  assign n3660 = ~n3649 & ~n3650;
  assign n3661 = n62468 & n62470;
  assign n3662 = ~n62468 & ~n62470;
  assign n3663 = ~n3661 & ~n3662;
  assign n3664 = n62468 & ~n62470;
  assign n3665 = ~n62468 & n62470;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = pi348 & ~n62467;
  assign n3668 = ~pi348 & n62467;
  assign n3669 = ~n3667 & ~n3668;
  assign n3670 = pi322 & n62468;
  assign n3671 = ~pi322 & ~n62468;
  assign n3672 = ~n3670 & ~n3671;
  assign n3673 = n3669 & ~n3672;
  assign n3674 = ~n3669 & n3672;
  assign n3675 = ~n3673 & ~n3674;
  assign n3676 = ~n62469 & n3675;
  assign n3677 = n62469 & ~n3675;
  assign n3678 = ~n3676 & ~n3677;
  assign n3679 = ~n3644 & ~n3645;
  assign n3680 = pi350 & n62471;
  assign n3681 = ~pi350 & ~n62471;
  assign n3682 = pi350 & ~n62471;
  assign n3683 = ~pi350 & n62471;
  assign n3684 = ~n3682 & ~n3683;
  assign n3685 = ~n3680 & ~n3681;
  assign n3686 = ~pi592 & pi1198;
  assign n3687 = ~n3680 & n3686;
  assign n3688 = ~n3681 & n3687;
  assign n3689 = ~n62472 & n3686;
  assign n3690 = n3022 & n62473;
  assign n3691 = n3615 & ~n3690;
  assign n3692 = ~n3135 & ~n62473;
  assign n3693 = n3691 & ~n3692;
  assign n3694 = pi1198 & n3614;
  assign n3695 = ~n62460 & ~n3694;
  assign n3696 = ~n3137 & ~n3695;
  assign n3697 = pi350 & ~pi592;
  assign n3698 = ~n3022 & n3697;
  assign n3699 = ~n62471 & ~n3698;
  assign n3700 = n3135 & ~n3697;
  assign n3701 = n3699 & ~n3700;
  assign n3702 = ~pi350 & ~pi592;
  assign n3703 = ~n3022 & n3702;
  assign n3704 = n62471 & ~n3703;
  assign n3705 = n3135 & ~n3702;
  assign n3706 = n3704 & ~n3705;
  assign n3707 = pi1198 & ~n3614;
  assign n3708 = ~n3706 & n3707;
  assign n3709 = ~n3701 & n3708;
  assign n3710 = pi1196 & n62465;
  assign n3711 = n3137 & n3710;
  assign n3712 = ~n3135 & ~n62465;
  assign n3713 = n62464 & ~n3712;
  assign n3714 = ~n3711 & n3713;
  assign n3715 = pi1196 & ~n62465;
  assign n3716 = n3137 & n3715;
  assign n3717 = ~n3135 & n62465;
  assign n3718 = ~n62464 & ~n3717;
  assign n3719 = ~n3716 & n3718;
  assign n3720 = ~n3714 & ~n3719;
  assign n3721 = ~pi1198 & ~n3205;
  assign n3722 = ~n3720 & n3721;
  assign n3723 = ~n3709 & ~n3722;
  assign n3724 = ~n62460 & ~n3723;
  assign n3725 = ~n3696 & ~n3724;
  assign n3726 = ~n3137 & n62460;
  assign n3727 = pi455 & ~n3137;
  assign n3728 = ~pi455 & n3135;
  assign n3729 = ~n3727 & ~n3728;
  assign n3730 = ~pi452 & ~n3729;
  assign n3731 = ~pi455 & ~n3137;
  assign n3732 = pi455 & n3135;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = pi452 & ~n3733;
  assign n3735 = ~n62465 & ~n3734;
  assign n3736 = ~n62465 & ~n3730;
  assign n3737 = ~n3734 & n3736;
  assign n3738 = ~n3730 & n3735;
  assign n3739 = ~pi452 & ~n3733;
  assign n3740 = pi452 & ~n3729;
  assign n3741 = n62465 & ~n3740;
  assign n3742 = n62465 & ~n3739;
  assign n3743 = ~n3740 & n3742;
  assign n3744 = ~n3739 & n3741;
  assign n3745 = pi1196 & ~n62476;
  assign n3746 = pi1196 & ~n62475;
  assign n3747 = ~n62476 & n3746;
  assign n3748 = ~n62475 & n3745;
  assign n3749 = ~pi1198 & ~n3207;
  assign n3750 = ~n62477 & n3749;
  assign n3751 = ~n3614 & ~n3706;
  assign n3752 = ~n3614 & ~n3701;
  assign n3753 = ~n3706 & n3752;
  assign n3754 = ~n3701 & n3751;
  assign n3755 = ~n3137 & n3614;
  assign n3756 = pi1198 & ~n3755;
  assign n3757 = ~n62478 & n3756;
  assign n3758 = ~n62460 & ~n3757;
  assign n3759 = ~n3750 & n3758;
  assign n3760 = ~n3726 & ~n3759;
  assign n3761 = ~n3616 & ~n3693;
  assign n3762 = ~n3478 & ~n62474;
  assign n3763 = pi1199 & ~n3137;
  assign n3764 = ~pi351 & n3763;
  assign n3765 = ~n3762 & ~n3764;
  assign n3766 = ~pi461 & ~n3765;
  assign n3767 = pi351 & pi1199;
  assign n3768 = ~n62474 & ~n3767;
  assign n3769 = pi351 & n3763;
  assign n3770 = ~n3768 & ~n3769;
  assign n3771 = pi461 & ~n3770;
  assign n3772 = ~n3766 & ~n3771;
  assign n3773 = ~pi357 & ~n3772;
  assign n3774 = ~pi461 & ~n3770;
  assign n3775 = pi461 & ~n3765;
  assign n3776 = ~n3774 & ~n3775;
  assign n3777 = pi357 & ~n3776;
  assign n3778 = ~n3773 & ~n3777;
  assign n3779 = pi356 & n3778;
  assign n3780 = pi360 & ~pi462;
  assign n3781 = ~pi360 & pi462;
  assign n3782 = ~pi360 & ~pi462;
  assign n3783 = pi360 & pi462;
  assign n3784 = ~n3782 & ~n3783;
  assign n3785 = ~n3780 & ~n3781;
  assign n3786 = pi352 & ~pi353;
  assign n3787 = ~pi352 & pi353;
  assign n3788 = ~n3786 & ~n3787;
  assign n3789 = ~n62479 & n3788;
  assign n3790 = n62479 & ~n3788;
  assign n3791 = n62479 & n3788;
  assign n3792 = ~n62479 & ~n3788;
  assign n3793 = ~n3791 & ~n3792;
  assign n3794 = ~n3789 & ~n3790;
  assign n3795 = pi354 & ~n62480;
  assign n3796 = ~pi354 & n62480;
  assign n3797 = pi354 & n62480;
  assign n3798 = ~pi354 & ~n62480;
  assign n3799 = ~n3797 & ~n3798;
  assign n3800 = ~n3795 & ~n3796;
  assign n3801 = ~pi357 & ~n3776;
  assign n3802 = pi357 & ~n3772;
  assign n3803 = ~n3801 & ~n3802;
  assign n3804 = ~pi356 & n3803;
  assign n3805 = n62481 & ~n3804;
  assign n3806 = ~pi356 & ~n3803;
  assign n3807 = pi356 & ~n3778;
  assign n3808 = ~n3806 & ~n3807;
  assign n3809 = n62481 & ~n3808;
  assign n3810 = ~n3779 & n3805;
  assign n3811 = pi356 & n3803;
  assign n3812 = ~pi356 & n3778;
  assign n3813 = ~n62481 & ~n3812;
  assign n3814 = ~pi356 & ~n3778;
  assign n3815 = pi356 & ~n3803;
  assign n3816 = ~n3814 & ~n3815;
  assign n3817 = ~n62481 & ~n3816;
  assign n3818 = ~n3811 & n3813;
  assign n3819 = pi590 & ~n62483;
  assign n3820 = ~n62482 & n3819;
  assign n3821 = pi592 & ~n3022;
  assign n3822 = ~pi592 & n3135;
  assign n3823 = ~n3821 & ~n3822;
  assign n3824 = pi1198 & ~n3823;
  assign n3825 = pi338 & ~pi388;
  assign n3826 = ~pi338 & pi388;
  assign n3827 = ~pi338 & ~pi388;
  assign n3828 = pi338 & pi388;
  assign n3829 = ~n3827 & ~n3828;
  assign n3830 = ~n3825 & ~n3826;
  assign n3831 = pi337 & n62484;
  assign n3832 = ~pi337 & ~n62484;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = pi363 & ~pi372;
  assign n3835 = ~pi363 & pi372;
  assign n3836 = ~pi363 & ~pi372;
  assign n3837 = pi363 & pi372;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = ~n3834 & ~n3835;
  assign n3840 = ~pi339 & ~pi386;
  assign n3841 = pi339 & pi386;
  assign n3842 = pi339 & ~pi386;
  assign n3843 = ~pi339 & pi386;
  assign n3844 = ~n3842 & ~n3843;
  assign n3845 = ~n3840 & ~n3841;
  assign n3846 = ~pi380 & ~pi387;
  assign n3847 = pi380 & pi387;
  assign n3848 = pi380 & ~pi387;
  assign n3849 = ~pi380 & pi387;
  assign n3850 = ~n3848 & ~n3849;
  assign n3851 = ~n3846 & ~n3847;
  assign n3852 = ~n62486 & n62487;
  assign n3853 = n62486 & ~n62487;
  assign n3854 = ~n3852 & ~n3853;
  assign n3855 = ~n62485 & n3854;
  assign n3856 = n62485 & ~n3854;
  assign n3857 = ~n62485 & n62487;
  assign n3858 = n62485 & ~n62487;
  assign n3859 = ~n3857 & ~n3858;
  assign n3860 = n62486 & n3859;
  assign n3861 = ~n62486 & ~n3859;
  assign n3862 = ~n3860 & ~n3861;
  assign n3863 = ~n3855 & ~n3856;
  assign n3864 = n3833 & ~n62488;
  assign n3865 = ~n3833 & n62488;
  assign n3866 = pi1196 & ~n3865;
  assign n3867 = pi386 & ~n62485;
  assign n3868 = ~pi386 & n62485;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = pi337 & ~pi339;
  assign n3871 = ~pi337 & pi339;
  assign n3872 = ~n3870 & ~n3871;
  assign n3873 = ~n62484 & n3872;
  assign n3874 = n62484 & ~n3872;
  assign n3875 = ~n3873 & ~n3874;
  assign n3876 = n3869 & ~n3875;
  assign n3877 = ~n3869 & n3875;
  assign n3878 = ~n3876 & ~n3877;
  assign n3879 = n62487 & n3878;
  assign n3880 = ~n62487 & ~n3878;
  assign n3881 = pi387 & n3872;
  assign n3882 = ~pi387 & ~n3872;
  assign n3883 = ~n3881 & ~n3882;
  assign n3884 = pi380 & ~n3883;
  assign n3885 = ~pi380 & n3883;
  assign n3886 = ~n3884 & ~n3885;
  assign n3887 = ~n62484 & ~n3886;
  assign n3888 = n62484 & n3886;
  assign n3889 = ~n3887 & ~n3888;
  assign n3890 = n3869 & n3889;
  assign n3891 = ~n3869 & ~n3889;
  assign n3892 = ~n3890 & ~n3891;
  assign n3893 = ~n3879 & ~n3880;
  assign n3894 = pi1196 & ~n62489;
  assign n3895 = ~n3864 & n3866;
  assign n3896 = ~pi368 & ~pi389;
  assign n3897 = pi368 & pi389;
  assign n3898 = pi368 & ~pi389;
  assign n3899 = ~pi368 & pi389;
  assign n3900 = ~n3898 & ~n3899;
  assign n3901 = ~n3896 & ~n3897;
  assign n3902 = pi336 & ~pi383;
  assign n3903 = ~pi336 & pi383;
  assign n3904 = ~pi336 & ~pi383;
  assign n3905 = pi336 & pi383;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = ~n3902 & ~n3903;
  assign n3908 = pi364 & ~pi366;
  assign n3909 = ~pi364 & pi366;
  assign n3910 = ~n3908 & ~n3909;
  assign n3911 = ~n62492 & n3910;
  assign n3912 = n62492 & ~n3910;
  assign n3913 = n62492 & n3910;
  assign n3914 = ~n62492 & ~n3910;
  assign n3915 = ~n3913 & ~n3914;
  assign n3916 = ~n3911 & ~n3912;
  assign n3917 = pi365 & ~pi447;
  assign n3918 = ~pi365 & pi447;
  assign n3919 = ~pi365 & ~pi447;
  assign n3920 = pi365 & pi447;
  assign n3921 = ~n3919 & ~n3920;
  assign n3922 = ~n3917 & ~n3918;
  assign n3923 = pi367 & n62494;
  assign n3924 = ~pi367 & ~n62494;
  assign n3925 = pi367 & ~n62494;
  assign n3926 = ~pi367 & n62494;
  assign n3927 = ~n3925 & ~n3926;
  assign n3928 = ~n3923 & ~n3924;
  assign n3929 = ~n62493 & ~n62495;
  assign n3930 = n62493 & n62495;
  assign n3931 = ~n62493 & ~n62494;
  assign n3932 = n62493 & n62494;
  assign n3933 = ~n3931 & ~n3932;
  assign n3934 = pi367 & ~n3933;
  assign n3935 = ~pi367 & n3933;
  assign n3936 = ~n3934 & ~n3935;
  assign n3937 = ~n3929 & ~n3930;
  assign n3938 = n62491 & ~n62496;
  assign n3939 = ~n62491 & n62496;
  assign n3940 = pi1197 & ~n3939;
  assign n3941 = n62491 & ~n62495;
  assign n3942 = ~n62491 & n62495;
  assign n3943 = ~n3941 & ~n3942;
  assign n3944 = ~n62493 & n3943;
  assign n3945 = n62493 & ~n3943;
  assign n3946 = ~n62491 & n3933;
  assign n3947 = n62491 & ~n3933;
  assign n3948 = ~n3946 & ~n3947;
  assign n3949 = pi367 & ~n3948;
  assign n3950 = ~pi367 & n3948;
  assign n3951 = ~n3949 & ~n3950;
  assign n3952 = ~n3944 & ~n3945;
  assign n3953 = pi1197 & n62497;
  assign n3954 = pi1197 & ~n3938;
  assign n3955 = ~n3939 & n3954;
  assign n3956 = ~n3938 & n3940;
  assign n3957 = ~n62490 & ~n62498;
  assign n3958 = pi379 & ~pi382;
  assign n3959 = ~pi379 & pi382;
  assign n3960 = ~pi379 & ~pi382;
  assign n3961 = pi379 & pi382;
  assign n3962 = ~n3960 & ~n3961;
  assign n3963 = ~n3958 & ~n3959;
  assign n3964 = pi377 & n62499;
  assign n3965 = ~pi377 & ~n62499;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = ~pi317 & ~pi385;
  assign n3968 = pi317 & pi385;
  assign n3969 = pi317 & ~pi385;
  assign n3970 = ~pi317 & pi385;
  assign n3971 = ~n3969 & ~n3970;
  assign n3972 = ~n3967 & ~n3968;
  assign n3973 = pi376 & ~pi439;
  assign n3974 = ~pi376 & pi439;
  assign n3975 = ~pi376 & ~pi439;
  assign n3976 = pi376 & pi439;
  assign n3977 = ~n3975 & ~n3976;
  assign n3978 = ~n3973 & ~n3974;
  assign n3979 = ~n62500 & ~n62501;
  assign n3980 = n62500 & n62501;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = pi378 & ~pi381;
  assign n3983 = ~pi378 & pi381;
  assign n3984 = ~n3982 & ~n3983;
  assign n3985 = n3981 & ~n3984;
  assign n3986 = ~n3981 & n3984;
  assign n3987 = pi381 & ~n62501;
  assign n3988 = ~pi381 & n62501;
  assign n3989 = ~n3987 & ~n3988;
  assign n3990 = pi378 & n62500;
  assign n3991 = ~pi378 & ~n62500;
  assign n3992 = ~n3990 & ~n3991;
  assign n3993 = n3989 & ~n3992;
  assign n3994 = ~n3989 & n3992;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = ~n3985 & ~n3986;
  assign n3997 = n3966 & n62502;
  assign n3998 = ~n3966 & ~n62502;
  assign n3999 = ~n62499 & n62502;
  assign n4000 = n62499 & ~n62502;
  assign n4001 = ~n62501 & n3984;
  assign n4002 = n62501 & ~n3984;
  assign n4003 = ~n4001 & ~n4002;
  assign n4004 = ~n62499 & ~n4003;
  assign n4005 = n62499 & n4003;
  assign n4006 = pi381 & n62499;
  assign n4007 = ~pi381 & ~n62499;
  assign n4008 = ~n4006 & ~n4007;
  assign n4009 = pi378 & n62501;
  assign n4010 = ~pi378 & ~n62501;
  assign n4011 = ~n4009 & ~n4010;
  assign n4012 = n4008 & ~n4011;
  assign n4013 = ~n4008 & n4011;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = ~n4004 & ~n4005;
  assign n4016 = n62500 & n62503;
  assign n4017 = ~n62500 & ~n62503;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = n62500 & ~n62503;
  assign n4020 = ~n62500 & n62503;
  assign n4021 = ~n4019 & ~n4020;
  assign n4022 = ~n3999 & ~n4000;
  assign n4023 = pi377 & ~n62504;
  assign n4024 = ~pi377 & n62504;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = ~pi377 & ~n62504;
  assign n4027 = pi377 & n62504;
  assign n4028 = ~n4026 & ~n4027;
  assign n4029 = ~n3997 & ~n3998;
  assign n4030 = pi1199 & ~n62505;
  assign n4031 = n3957 & ~n4030;
  assign n4032 = pi592 & ~n4031;
  assign n4033 = ~n3022 & n4032;
  assign n4034 = n3135 & ~n4032;
  assign n4035 = n3823 & ~n3957;
  assign n4036 = ~pi377 & pi592;
  assign n4037 = ~n3022 & n4036;
  assign n4038 = n62504 & ~n4037;
  assign n4039 = n3135 & ~n4036;
  assign n4040 = n4038 & ~n4039;
  assign n4041 = pi377 & pi592;
  assign n4042 = ~n3022 & n4041;
  assign n4043 = ~n62504 & ~n4042;
  assign n4044 = n3135 & ~n4041;
  assign n4045 = n4043 & ~n4044;
  assign n4046 = ~n4040 & ~n4045;
  assign n4047 = pi1199 & ~n4046;
  assign n4048 = ~pi1199 & ~n3135;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = n3957 & ~n4049;
  assign n4051 = ~n4035 & ~n4050;
  assign n4052 = ~n3135 & n3957;
  assign n4053 = ~pi1199 & ~n4052;
  assign n4054 = ~n4035 & n4053;
  assign n4055 = n3957 & ~n4046;
  assign n4056 = pi1199 & ~n4035;
  assign n4057 = ~n4055 & n4056;
  assign n4058 = ~n4054 & ~n4057;
  assign n4059 = ~n4033 & ~n4034;
  assign n4060 = ~pi1198 & n62506;
  assign n4061 = ~pi1198 & ~n62506;
  assign n4062 = pi1198 & n3823;
  assign n4063 = ~n4061 & ~n4062;
  assign n4064 = ~n3824 & ~n4060;
  assign n4065 = ~pi374 & ~n62507;
  assign n4066 = pi374 & ~n62506;
  assign n4067 = ~pi369 & ~n4066;
  assign n4068 = ~pi374 & n62507;
  assign n4069 = pi374 & n62506;
  assign n4070 = ~n4065 & ~n4066;
  assign n4071 = ~n4068 & ~n4069;
  assign n4072 = ~pi369 & n62508;
  assign n4073 = ~n4065 & n4067;
  assign n4074 = pi374 & ~n62507;
  assign n4075 = ~pi374 & ~n62506;
  assign n4076 = pi369 & ~n4075;
  assign n4077 = ~pi374 & n62506;
  assign n4078 = pi374 & n62507;
  assign n4079 = ~n4074 & ~n4075;
  assign n4080 = ~n4077 & ~n4078;
  assign n4081 = pi369 & n62510;
  assign n4082 = ~n4074 & n4076;
  assign n4083 = ~pi369 & ~n62508;
  assign n4084 = pi369 & ~n62510;
  assign n4085 = ~n4083 & ~n4084;
  assign n4086 = ~n62509 & ~n62511;
  assign n4087 = pi384 & ~pi442;
  assign n4088 = ~pi384 & pi442;
  assign n4089 = ~pi384 & ~pi442;
  assign n4090 = pi384 & pi442;
  assign n4091 = ~n4089 & ~n4090;
  assign n4092 = ~n4087 & ~n4088;
  assign n4093 = pi375 & ~pi440;
  assign n4094 = ~pi375 & pi440;
  assign n4095 = ~n4093 & ~n4094;
  assign n4096 = ~n62513 & n4095;
  assign n4097 = n62513 & ~n4095;
  assign n4098 = pi440 & n62513;
  assign n4099 = ~pi440 & ~n62513;
  assign n4100 = ~n4098 & ~n4099;
  assign n4101 = pi375 & ~n4100;
  assign n4102 = ~pi375 & n4100;
  assign n4103 = ~n4101 & ~n4102;
  assign n4104 = pi375 & n4100;
  assign n4105 = ~pi375 & ~n4100;
  assign n4106 = ~n4104 & ~n4105;
  assign n4107 = ~n4096 & ~n4097;
  assign n4108 = pi371 & ~pi373;
  assign n4109 = ~pi371 & pi373;
  assign n4110 = ~n4108 & ~n4109;
  assign n4111 = ~n62514 & n4110;
  assign n4112 = n62514 & ~n4110;
  assign n4113 = pi373 & n62514;
  assign n4114 = ~pi373 & ~n62514;
  assign n4115 = pi373 & ~pi375;
  assign n4116 = ~pi373 & pi375;
  assign n4117 = ~n4115 & ~n4116;
  assign n4118 = n4100 & n4117;
  assign n4119 = ~n4100 & ~n4117;
  assign n4120 = ~n4118 & ~n4119;
  assign n4121 = pi373 & ~n4100;
  assign n4122 = ~pi373 & n4100;
  assign n4123 = ~n4121 & ~n4122;
  assign n4124 = pi375 & n4123;
  assign n4125 = ~pi375 & ~n4123;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = ~n4113 & ~n4114;
  assign n4128 = pi371 & n62515;
  assign n4129 = ~pi371 & ~n62515;
  assign n4130 = ~n4128 & ~n4129;
  assign n4131 = ~n4111 & ~n4112;
  assign n4132 = pi370 & ~n62516;
  assign n4133 = ~pi370 & n62516;
  assign n4134 = pi370 & ~pi371;
  assign n4135 = ~pi370 & pi371;
  assign n4136 = ~pi370 & ~pi371;
  assign n4137 = pi370 & pi371;
  assign n4138 = ~n4136 & ~n4137;
  assign n4139 = ~n4134 & ~n4135;
  assign n4140 = ~n62515 & ~n62517;
  assign n4141 = n62515 & n62517;
  assign n4142 = ~n4140 & ~n4141;
  assign n4143 = n62515 & ~n62517;
  assign n4144 = ~n62515 & n62517;
  assign n4145 = ~n4143 & ~n4144;
  assign n4146 = pi370 & n62516;
  assign n4147 = ~pi370 & ~n62516;
  assign n4148 = ~n4146 & ~n4147;
  assign n4149 = ~n4132 & ~n4133;
  assign n4150 = n62512 & ~n62518;
  assign n4151 = pi369 & ~pi374;
  assign n4152 = ~pi369 & pi374;
  assign n4153 = ~pi369 & ~pi374;
  assign n4154 = pi369 & pi374;
  assign n4155 = ~n4153 & ~n4154;
  assign n4156 = ~n4151 & ~n4152;
  assign n4157 = ~n62507 & n62519;
  assign n4158 = ~n62506 & ~n62519;
  assign n4159 = n62518 & ~n4158;
  assign n4160 = ~n4157 & n4159;
  assign n4161 = ~pi590 & ~n4160;
  assign n4162 = ~n4150 & n4161;
  assign n4163 = ~pi591 & ~n4162;
  assign n4164 = ~n3820 & n4163;
  assign n4165 = pi335 & ~pi393;
  assign n4166 = ~pi335 & pi393;
  assign n4167 = ~n4165 & ~n4166;
  assign n4168 = pi407 & ~pi463;
  assign n4169 = ~pi407 & pi463;
  assign n4170 = ~pi407 & ~pi463;
  assign n4171 = pi407 & pi463;
  assign n4172 = ~n4170 & ~n4171;
  assign n4173 = ~n4168 & ~n4169;
  assign n4174 = ~pi334 & ~pi413;
  assign n4175 = pi334 & pi413;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = ~n62520 & ~n4176;
  assign n4178 = n62520 & n4176;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180 = n4167 & n4179;
  assign n4181 = ~n4167 & ~n4179;
  assign n4182 = pi335 & ~pi413;
  assign n4183 = ~pi335 & pi413;
  assign n4184 = ~n4182 & ~n4183;
  assign n4185 = ~n62520 & n4184;
  assign n4186 = n62520 & ~n4184;
  assign n4187 = n62520 & n4184;
  assign n4188 = ~n62520 & ~n4184;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = ~n4185 & ~n4186;
  assign n4191 = pi334 & n62521;
  assign n4192 = ~pi334 & ~n62521;
  assign n4193 = pi334 & ~n62521;
  assign n4194 = ~pi334 & n62521;
  assign n4195 = ~n4193 & ~n4194;
  assign n4196 = ~n4191 & ~n4192;
  assign n4197 = pi393 & n62522;
  assign n4198 = ~pi393 & ~n62522;
  assign n4199 = ~n4197 & ~n4198;
  assign n4200 = pi393 & ~n62522;
  assign n4201 = ~pi393 & n62522;
  assign n4202 = ~n4200 & ~n4201;
  assign n4203 = ~n4180 & ~n4181;
  assign n4204 = ~pi392 & n62523;
  assign n4205 = pi392 & ~n62523;
  assign n4206 = ~n4204 & ~n4205;
  assign n4207 = pi391 & ~n4206;
  assign n4208 = ~pi391 & n4206;
  assign n4209 = ~n4207 & ~n4208;
  assign n4210 = ~pi333 & pi1197;
  assign n4211 = ~n3137 & n4210;
  assign n4212 = pi319 & ~pi324;
  assign n4213 = ~pi319 & pi324;
  assign n4214 = ~pi319 & ~pi324;
  assign n4215 = pi319 & pi324;
  assign n4216 = ~n4214 & ~n4215;
  assign n4217 = ~n4212 & ~n4213;
  assign n4218 = pi456 & n62524;
  assign n4219 = ~pi456 & ~n62524;
  assign n4220 = ~n4218 & ~n4219;
  assign n4221 = pi411 & ~n4220;
  assign n4222 = ~pi411 & n4220;
  assign n4223 = ~n4221 & ~n4222;
  assign n4224 = pi390 & ~pi410;
  assign n4225 = ~pi390 & pi410;
  assign n4226 = ~pi390 & ~pi410;
  assign n4227 = pi390 & pi410;
  assign n4228 = ~n4226 & ~n4227;
  assign n4229 = ~n4224 & ~n4225;
  assign n4230 = pi412 & ~n62525;
  assign n4231 = ~pi412 & n62525;
  assign n4232 = ~n4230 & ~n4231;
  assign n4233 = pi397 & ~pi404;
  assign n4234 = ~pi397 & pi404;
  assign n4235 = ~pi397 & ~pi404;
  assign n4236 = pi397 & pi404;
  assign n4237 = ~n4235 & ~n4236;
  assign n4238 = ~n4233 & ~n4234;
  assign n4239 = n4232 & n62526;
  assign n4240 = ~n4232 & ~n62526;
  assign n4241 = pi397 & ~pi412;
  assign n4242 = ~pi397 & pi412;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = pi404 & n4243;
  assign n4245 = ~pi404 & ~n4243;
  assign n4246 = pi412 & n62526;
  assign n4247 = ~pi412 & ~n62526;
  assign n4248 = ~n4246 & ~n4247;
  assign n4249 = ~n4244 & ~n4245;
  assign n4250 = n62525 & n62527;
  assign n4251 = ~n62525 & ~n62527;
  assign n4252 = ~n4250 & ~n4251;
  assign n4253 = ~n4239 & ~n4240;
  assign n4254 = n4223 & ~n62528;
  assign n4255 = ~n4223 & n62528;
  assign n4256 = pi411 & n62526;
  assign n4257 = ~pi411 & ~n62526;
  assign n4258 = ~n4256 & ~n4257;
  assign n4259 = n62525 & n4258;
  assign n4260 = ~n62525 & ~n4258;
  assign n4261 = pi411 & n62525;
  assign n4262 = ~pi411 & ~n62525;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264 = n62526 & ~n4263;
  assign n4265 = ~n62526 & n4263;
  assign n4266 = ~n4264 & ~n4265;
  assign n4267 = ~n62525 & n4258;
  assign n4268 = n62525 & ~n4258;
  assign n4269 = ~n4267 & ~n4268;
  assign n4270 = ~n4259 & ~n4260;
  assign n4271 = pi412 & ~n4220;
  assign n4272 = ~pi412 & n4220;
  assign n4273 = ~n4271 & ~n4272;
  assign n4274 = n62529 & n4273;
  assign n4275 = ~n62529 & ~n4273;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = ~n4220 & ~n62527;
  assign n4278 = n4220 & n62527;
  assign n4279 = ~n4277 & ~n4278;
  assign n4280 = ~n62525 & n4279;
  assign n4281 = n62525 & ~n4279;
  assign n4282 = n4220 & n62528;
  assign n4283 = ~n4220 & ~n62528;
  assign n4284 = ~n4282 & ~n4283;
  assign n4285 = ~n4280 & ~n4281;
  assign n4286 = pi411 & ~n62531;
  assign n4287 = ~pi411 & n62531;
  assign n4288 = ~n4286 & ~n4287;
  assign n4289 = ~n4254 & ~n4255;
  assign n4290 = n2899 & n62530;
  assign n4291 = n3047 & ~n4290;
  assign n4292 = ~pi403 & ~pi405;
  assign n4293 = pi403 & pi405;
  assign n4294 = pi403 & ~pi405;
  assign n4295 = ~pi403 & pi405;
  assign n4296 = ~n4294 & ~n4295;
  assign n4297 = ~n4292 & ~n4293;
  assign n4298 = pi406 & n62532;
  assign n4299 = ~pi406 & ~n62532;
  assign n4300 = ~n4298 & ~n4299;
  assign n4301 = pi318 & ~pi409;
  assign n4302 = ~pi318 & pi409;
  assign n4303 = ~pi318 & ~pi409;
  assign n4304 = pi318 & pi409;
  assign n4305 = ~n4303 & ~n4304;
  assign n4306 = ~n4301 & ~n4302;
  assign n4307 = n4300 & n62533;
  assign n4308 = ~n4300 & ~n62533;
  assign n4309 = ~n4307 & ~n4308;
  assign n4310 = ~pi401 & ~pi402;
  assign n4311 = pi401 & pi402;
  assign n4312 = pi401 & ~pi402;
  assign n4313 = ~pi401 & pi402;
  assign n4314 = ~n4312 & ~n4313;
  assign n4315 = ~n4310 & ~n4311;
  assign n4316 = pi325 & ~pi326;
  assign n4317 = ~pi325 & pi326;
  assign n4318 = ~n4316 & ~n4317;
  assign n4319 = ~n62534 & ~n4318;
  assign n4320 = n62534 & n4318;
  assign n4321 = ~n4319 & ~n4320;
  assign n4322 = n4309 & n4321;
  assign n4323 = ~n4309 & ~n4321;
  assign n4324 = pi325 & n62533;
  assign n4325 = ~pi325 & ~n62533;
  assign n4326 = ~n4324 & ~n4325;
  assign n4327 = pi326 & ~n4326;
  assign n4328 = ~pi326 & n4326;
  assign n4329 = ~n4327 & ~n4328;
  assign n4330 = n4300 & n62534;
  assign n4331 = ~n4300 & ~n62534;
  assign n4332 = ~n4330 & ~n4331;
  assign n4333 = n4329 & n4332;
  assign n4334 = ~n4329 & ~n4332;
  assign n4335 = ~n4333 & ~n4334;
  assign n4336 = pi326 & ~pi406;
  assign n4337 = ~pi326 & pi406;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = n62534 & n4338;
  assign n4340 = ~n62534 & ~n4338;
  assign n4341 = ~n4339 & ~n4340;
  assign n4342 = ~n62532 & ~n4341;
  assign n4343 = n62532 & n4341;
  assign n4344 = ~n4342 & ~n4343;
  assign n4345 = n4326 & n4344;
  assign n4346 = ~n4326 & ~n4344;
  assign n4347 = ~n4345 & ~n4346;
  assign n4348 = pi406 & n62534;
  assign n4349 = ~pi406 & ~n62534;
  assign n4350 = ~n4348 & ~n4349;
  assign n4351 = ~n62532 & n4318;
  assign n4352 = n62532 & ~n4318;
  assign n4353 = ~n4351 & ~n4352;
  assign n4354 = n4350 & ~n4353;
  assign n4355 = ~n4350 & n4353;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = ~n62533 & n4356;
  assign n4358 = n62533 & ~n4356;
  assign n4359 = ~n4357 & ~n4358;
  assign n4360 = ~n4322 & ~n4323;
  assign n4361 = n2854 & n62535;
  assign n4362 = pi122 & ~n4361;
  assign n4363 = n3027 & n62535;
  assign n4364 = ~pi122 & ~n4363;
  assign n4365 = pi1093 & ~n4364;
  assign n4366 = n3045 & n62535;
  assign n4367 = ~n4362 & n4365;
  assign n4368 = n2899 & ~n62536;
  assign n4369 = n4291 & ~n4368;
  assign n4370 = pi1093 & ~n2909;
  assign n4371 = n2971 & n4370;
  assign n4372 = n2953 & ~n2971;
  assign n4373 = n3076 & ~n4372;
  assign n4374 = ~n4371 & n4373;
  assign n4375 = ~n2975 & n3076;
  assign n4376 = ~n2974 & n4375;
  assign n4377 = n62402 & n3076;
  assign n4378 = n62397 & n4374;
  assign n4379 = ~pi299 & ~n62537;
  assign n4380 = n62393 & n4370;
  assign n4381 = ~n62393 & n2953;
  assign n4382 = n3056 & ~n4381;
  assign n4383 = ~n4380 & n4382;
  assign n4384 = ~n2955 & n3056;
  assign n4385 = ~n2951 & n4384;
  assign n4386 = n62400 & n3056;
  assign n4387 = n62397 & n4383;
  assign n4388 = pi299 & ~n62538;
  assign n4389 = ~n2964 & ~n2985;
  assign n4390 = ~n4379 & ~n4388;
  assign n4391 = n3029 & ~n62530;
  assign n4392 = ~pi1091 & n4391;
  assign n4393 = n62409 & ~n62530;
  assign n4394 = n3028 & n4363;
  assign n4395 = n3029 & n62535;
  assign n4396 = ~pi1091 & n62541;
  assign n4397 = n62409 & n62535;
  assign n4398 = ~n62530 & n62542;
  assign n4399 = n62535 & n62540;
  assign n4400 = n62539 & ~n62543;
  assign n4401 = ~n3076 & n62540;
  assign n4402 = ~pi299 & ~n4401;
  assign n4403 = ~n3076 & n62542;
  assign n4404 = ~pi299 & ~n4403;
  assign n4405 = ~n4402 & ~n4404;
  assign n4406 = ~n2950 & ~n62543;
  assign n4407 = n2971 & n4406;
  assign n4408 = ~n2954 & ~n62543;
  assign n4409 = ~n2971 & n4408;
  assign n4410 = n3076 & ~n4409;
  assign n4411 = n3076 & ~n4407;
  assign n4412 = ~n4409 & n4411;
  assign n4413 = ~n4407 & n4410;
  assign n4414 = ~n4405 & ~n62544;
  assign n4415 = n4379 & ~n62543;
  assign n4416 = ~n3056 & n62540;
  assign n4417 = pi299 & ~n4416;
  assign n4418 = ~n3056 & n62542;
  assign n4419 = pi299 & ~n4418;
  assign n4420 = ~n3056 & n62543;
  assign n4421 = pi299 & ~n4420;
  assign n4422 = ~n4417 & ~n4419;
  assign n4423 = ~n62400 & ~n62543;
  assign n4424 = n62393 & n4406;
  assign n4425 = ~n62393 & n4408;
  assign n4426 = n3056 & ~n4425;
  assign n4427 = ~n4424 & n4426;
  assign n4428 = n3056 & ~n4424;
  assign n4429 = ~n4425 & n4428;
  assign n4430 = n3056 & ~n4423;
  assign n4431 = n62546 & ~n62547;
  assign n4432 = pi39 & ~n4431;
  assign n4433 = ~n62545 & n4432;
  assign n4434 = pi39 & ~n62545;
  assign n4435 = ~n4431 & n4434;
  assign n4436 = pi39 & ~n4400;
  assign n4437 = ~n4369 & ~n62548;
  assign n4438 = ~pi38 & ~n4437;
  assign n4439 = pi38 & n62540;
  assign n4440 = ~pi100 & ~n4439;
  assign n4441 = pi38 & n62542;
  assign n4442 = ~pi100 & ~n4441;
  assign n4443 = ~n4440 & ~n4442;
  assign n4444 = ~n4438 & ~n4443;
  assign n4445 = ~pi1091 & ~n62543;
  assign n4446 = ~n2998 & ~n62543;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = n2995 & n4447;
  assign n4449 = pi100 & ~n62543;
  assign n4450 = ~n2995 & ~n62543;
  assign n4451 = n4447 & ~n4450;
  assign n4452 = pi100 & ~n4451;
  assign n4453 = n2809 & n2996;
  assign n4454 = ~n2812 & n2814;
  assign n4455 = ~n2809 & ~n4454;
  assign n4456 = ~n4445 & n4455;
  assign n4457 = ~n3099 & n4456;
  assign n4458 = ~n4453 & ~n4457;
  assign n4459 = pi228 & ~n4458;
  assign n4460 = pi228 & n4455;
  assign n4461 = n62543 & ~n4460;
  assign n4462 = pi232 & ~n4461;
  assign n4463 = ~n4459 & n4462;
  assign n4464 = ~pi232 & ~n62543;
  assign n4465 = ~n2999 & n4464;
  assign n4466 = n2764 & ~n4465;
  assign n4467 = ~n4463 & n4466;
  assign n4468 = ~n2764 & n62543;
  assign n4469 = pi100 & ~n4468;
  assign n4470 = ~n4467 & n4469;
  assign n4471 = ~n4448 & n4449;
  assign n4472 = ~n4444 & ~n62549;
  assign n4473 = ~pi87 & ~n4472;
  assign n4474 = ~n62373 & n62540;
  assign n4475 = pi87 & ~n4474;
  assign n4476 = ~n62373 & n62542;
  assign n4477 = pi87 & ~n4476;
  assign n4478 = ~n4475 & ~n4477;
  assign n4479 = n3006 & n62530;
  assign n4480 = n3006 & ~n62535;
  assign n4481 = n3123 & ~n4480;
  assign n4482 = ~n4479 & n4481;
  assign n4483 = ~n4478 & ~n4482;
  assign n4484 = ~n4473 & ~n4483;
  assign n4485 = ~pi75 & ~n4484;
  assign n4486 = ~n2817 & n62540;
  assign n4487 = pi75 & ~n4486;
  assign n4488 = ~n2817 & n62542;
  assign n4489 = pi75 & ~n4488;
  assign n4490 = ~n4487 & ~n4489;
  assign n4491 = n3026 & ~n4445;
  assign n4492 = ~n4490 & ~n4491;
  assign n4493 = ~n4485 & ~n4492;
  assign n4494 = ~pi592 & pi1196;
  assign n4495 = pi567 & n62540;
  assign n4496 = ~n2580 & n4495;
  assign n4497 = n3131 & n62540;
  assign n4498 = n4363 & n62550;
  assign n4499 = n4494 & ~n4498;
  assign n4500 = ~n4493 & n4499;
  assign n4501 = n4477 & ~n4481;
  assign n4502 = n3003 & ~n62542;
  assign n4503 = n3042 & ~n4368;
  assign n4504 = n62539 & ~n62542;
  assign n4505 = ~n2954 & ~n62542;
  assign n4506 = ~n2971 & n4505;
  assign n4507 = ~n2950 & ~n62542;
  assign n4508 = n2971 & n4507;
  assign n4509 = n3076 & ~n4508;
  assign n4510 = n3076 & ~n4506;
  assign n4511 = ~n4508 & n4510;
  assign n4512 = ~n4506 & n4509;
  assign n4513 = n4404 & ~n62551;
  assign n4514 = ~n62393 & n4505;
  assign n4515 = n62393 & n4507;
  assign n4516 = n3056 & ~n4515;
  assign n4517 = n3056 & ~n4514;
  assign n4518 = ~n4515 & n4517;
  assign n4519 = ~n4514 & n4516;
  assign n4520 = n4419 & ~n62552;
  assign n4521 = pi39 & ~n4520;
  assign n4522 = ~n4513 & n4521;
  assign n4523 = pi39 & ~n4513;
  assign n4524 = ~n4520 & n4523;
  assign n4525 = pi39 & ~n4504;
  assign n4526 = ~n4503 & ~n62553;
  assign n4527 = ~pi38 & ~n4526;
  assign n4528 = n4442 & ~n4527;
  assign n4529 = ~n4502 & ~n4528;
  assign n4530 = ~pi87 & ~n4529;
  assign n4531 = ~n4501 & ~n4530;
  assign n4532 = ~pi75 & ~n4531;
  assign n4533 = ~pi1091 & ~n62541;
  assign n4534 = n3026 & ~n4533;
  assign n4535 = n4489 & ~n4534;
  assign n4536 = ~n4532 & ~n4535;
  assign n4537 = ~pi592 & ~pi1196;
  assign n4538 = pi567 & n62542;
  assign n4539 = ~n2580 & n4538;
  assign n4540 = n62422 & n62535;
  assign n4541 = n4537 & ~n62554;
  assign n4542 = ~n4536 & n4541;
  assign n4543 = ~n4500 & ~n4542;
  assign n4544 = pi567 & ~n4543;
  assign n4545 = ~n4499 & ~n4541;
  assign n4546 = ~n2804 & ~n4545;
  assign n4547 = pi1199 & ~n4546;
  assign n4548 = ~n4544 & n4547;
  assign n4549 = pi328 & ~pi408;
  assign n4550 = ~pi328 & pi408;
  assign n4551 = ~n4549 & ~n4550;
  assign n4552 = pi398 & ~pi399;
  assign n4553 = ~pi398 & pi399;
  assign n4554 = ~pi398 & ~pi399;
  assign n4555 = pi398 & pi399;
  assign n4556 = ~n4554 & ~n4555;
  assign n4557 = ~n4552 & ~n4553;
  assign n4558 = pi394 & ~n62555;
  assign n4559 = ~pi394 & n62555;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = pi329 & ~pi395;
  assign n4562 = ~pi329 & pi395;
  assign n4563 = ~pi329 & ~pi395;
  assign n4564 = pi329 & pi395;
  assign n4565 = ~n4563 & ~n4564;
  assign n4566 = ~n4561 & ~n4562;
  assign n4567 = pi396 & ~pi400;
  assign n4568 = ~pi396 & pi400;
  assign n4569 = ~n4567 & ~n4568;
  assign n4570 = ~n62556 & n4569;
  assign n4571 = n62556 & ~n4569;
  assign n4572 = ~n4570 & ~n4571;
  assign n4573 = n4560 & ~n4572;
  assign n4574 = ~n4560 & n4572;
  assign n4575 = pi396 & n62556;
  assign n4576 = ~pi396 & ~n62556;
  assign n4577 = ~n4575 & ~n4576;
  assign n4578 = pi394 & ~pi400;
  assign n4579 = ~pi394 & pi400;
  assign n4580 = ~n4578 & ~n4579;
  assign n4581 = n62555 & n4580;
  assign n4582 = ~n62555 & ~n4580;
  assign n4583 = ~n4581 & ~n4582;
  assign n4584 = n4577 & ~n4583;
  assign n4585 = ~n4577 & n4583;
  assign n4586 = ~n4584 & ~n4585;
  assign n4587 = ~n4573 & ~n4574;
  assign n4588 = n4551 & n62557;
  assign n4589 = ~n4551 & ~n62557;
  assign n4590 = pi400 & n62555;
  assign n4591 = ~pi400 & ~n62555;
  assign n4592 = ~n4590 & ~n4591;
  assign n4593 = pi394 & ~n4551;
  assign n4594 = ~pi394 & n4551;
  assign n4595 = ~n4593 & ~n4594;
  assign n4596 = n4592 & ~n4595;
  assign n4597 = ~n4592 & n4595;
  assign n4598 = ~n4596 & ~n4597;
  assign n4599 = n4577 & n4598;
  assign n4600 = ~n4577 & ~n4598;
  assign n4601 = ~n4599 & ~n4600;
  assign n4602 = ~pi394 & ~pi396;
  assign n4603 = pi394 & pi396;
  assign n4604 = ~n4602 & ~n4603;
  assign n4605 = n4551 & ~n4604;
  assign n4606 = ~n4551 & n4604;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = pi395 & ~n62555;
  assign n4609 = ~pi395 & n62555;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = pi329 & ~n4610;
  assign n4612 = ~pi329 & n4610;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 = pi400 & ~n4613;
  assign n4615 = ~pi400 & n4613;
  assign n4616 = ~n4614 & ~n4615;
  assign n4617 = n4607 & n4616;
  assign n4618 = ~n4607 & ~n4616;
  assign n4619 = ~n4617 & ~n4618;
  assign n4620 = ~n4588 & ~n4589;
  assign n4621 = pi1198 & ~n62558;
  assign n4622 = ~n2954 & ~n62540;
  assign n4623 = ~n2971 & n4622;
  assign n4624 = ~n2950 & ~n62540;
  assign n4625 = n2971 & n4624;
  assign n4626 = n3076 & ~n4625;
  assign n4627 = n3076 & ~n4623;
  assign n4628 = ~n4625 & n4627;
  assign n4629 = ~n4623 & n4626;
  assign n4630 = n4402 & ~n62559;
  assign n4631 = n4379 & ~n62540;
  assign n4632 = pi299 & ~n62540;
  assign n4633 = ~n62393 & n4622;
  assign n4634 = n62393 & n4624;
  assign n4635 = n3056 & ~n4634;
  assign n4636 = n3056 & ~n4633;
  assign n4637 = ~n4634 & n4636;
  assign n4638 = ~n4633 & n4635;
  assign n4639 = n4417 & ~n62561;
  assign n4640 = ~n62538 & n4632;
  assign n4641 = pi39 & ~n62562;
  assign n4642 = n62539 & ~n62540;
  assign n4643 = pi39 & ~n4642;
  assign n4644 = pi39 & ~n62560;
  assign n4645 = ~n62562 & n4644;
  assign n4646 = ~n62560 & n4641;
  assign n4647 = ~n4291 & ~n62563;
  assign n4648 = ~pi38 & ~n4647;
  assign n4649 = n4440 & ~n4648;
  assign n4650 = n3003 & ~n62540;
  assign n4651 = ~n4649 & ~n4650;
  assign n4652 = ~pi87 & ~n4651;
  assign n4653 = n3123 & ~n4479;
  assign n4654 = n4475 & ~n4653;
  assign n4655 = ~n4652 & ~n4654;
  assign n4656 = ~pi75 & ~n4655;
  assign n4657 = ~pi1091 & ~n4391;
  assign n4658 = n3026 & ~n4657;
  assign n4659 = n4487 & ~n4658;
  assign n4660 = ~n4656 & ~n4659;
  assign n4661 = pi567 & ~n4660;
  assign n4662 = n2804 & ~n4661;
  assign n4663 = n4494 & ~n62550;
  assign n4664 = ~n4662 & n4663;
  assign n4665 = ~pi1199 & ~n3207;
  assign n4666 = ~n4664 & n4665;
  assign n4667 = ~n4621 & ~n4666;
  assign n4668 = ~n4548 & n4667;
  assign n4669 = n3023 & n4621;
  assign n4670 = ~n3136 & ~n4669;
  assign n4671 = ~n4668 & n4670;
  assign n4672 = ~n4210 & ~n4671;
  assign n4673 = ~pi1197 & ~n4671;
  assign n4674 = pi1197 & ~n3137;
  assign n4675 = ~n4673 & ~n4674;
  assign n4676 = ~pi333 & ~n4675;
  assign n4677 = pi333 & ~n4671;
  assign n4678 = ~n4676 & ~n4677;
  assign n4679 = ~n4211 & ~n4672;
  assign n4680 = n4209 & ~n62564;
  assign n4681 = pi333 & pi1197;
  assign n4682 = ~n3137 & n4681;
  assign n4683 = ~n4671 & ~n4681;
  assign n4684 = n4671 & ~n4681;
  assign n4685 = n3137 & n4681;
  assign n4686 = ~n4684 & ~n4685;
  assign n4687 = ~pi333 & ~n4671;
  assign n4688 = pi333 & ~n4675;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = ~n4682 & ~n4683;
  assign n4691 = ~n4209 & n62565;
  assign n4692 = ~pi590 & ~n4691;
  assign n4693 = ~n4680 & n4692;
  assign n4694 = pi590 & ~n3135;
  assign n4695 = pi591 & ~n4694;
  assign n4696 = ~n4693 & n4695;
  assign n4697 = ~n3318 & ~n4696;
  assign n4698 = ~pi370 & n62512;
  assign n4699 = ~pi369 & n62510;
  assign n4700 = pi369 & n62508;
  assign n4701 = pi369 & ~n62508;
  assign n4702 = ~pi369 & ~n62510;
  assign n4703 = ~n4701 & ~n4702;
  assign n4704 = ~n4699 & ~n4700;
  assign n4705 = pi370 & n62566;
  assign n4706 = pi370 & ~n62566;
  assign n4707 = ~pi370 & ~n62512;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = ~n4698 & ~n4705;
  assign n4710 = ~pi371 & n62567;
  assign n4711 = ~pi370 & n62566;
  assign n4712 = pi370 & n62512;
  assign n4713 = pi370 & ~n62512;
  assign n4714 = ~pi370 & ~n62566;
  assign n4715 = ~n4713 & ~n4714;
  assign n4716 = ~n4711 & ~n4712;
  assign n4717 = pi371 & n62568;
  assign n4718 = ~n4710 & ~n4717;
  assign n4719 = pi371 & ~n62568;
  assign n4720 = ~pi371 & ~n62567;
  assign n4721 = ~n62515 & ~n4720;
  assign n4722 = ~n4719 & n4721;
  assign n4723 = ~n62515 & ~n4718;
  assign n4724 = ~pi371 & n62568;
  assign n4725 = pi371 & n62567;
  assign n4726 = ~n4724 & ~n4725;
  assign n4727 = pi371 & ~n62567;
  assign n4728 = ~pi371 & ~n62568;
  assign n4729 = n62515 & ~n4728;
  assign n4730 = ~n4727 & n4729;
  assign n4731 = n62515 & ~n4726;
  assign n4732 = ~pi591 & ~n62570;
  assign n4733 = ~pi591 & ~n62569;
  assign n4734 = ~n62570 & n4733;
  assign n4735 = ~n62515 & ~n4710;
  assign n4736 = ~n4717 & n4735;
  assign n4737 = n62515 & ~n4724;
  assign n4738 = ~n4725 & n4737;
  assign n4739 = ~n4736 & ~n4738;
  assign n4740 = ~pi591 & ~n4739;
  assign n4741 = ~n62569 & n4732;
  assign n4742 = ~pi391 & ~n62564;
  assign n4743 = pi391 & n62565;
  assign n4744 = pi391 & ~n62565;
  assign n4745 = ~pi391 & n62564;
  assign n4746 = ~n4744 & ~n4745;
  assign n4747 = ~n4742 & ~n4743;
  assign n4748 = ~pi392 & n62572;
  assign n4749 = ~pi391 & n62565;
  assign n4750 = pi391 & ~n62564;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = pi392 & ~n4751;
  assign n4753 = ~n4748 & ~n4752;
  assign n4754 = pi392 & n4751;
  assign n4755 = ~pi392 & ~n62572;
  assign n4756 = n62523 & ~n4755;
  assign n4757 = ~n4754 & n4756;
  assign n4758 = n62523 & ~n4754;
  assign n4759 = ~n4755 & n4758;
  assign n4760 = n62523 & ~n4753;
  assign n4761 = ~pi392 & ~n4751;
  assign n4762 = pi392 & n62572;
  assign n4763 = ~n4761 & ~n4762;
  assign n4764 = pi392 & ~n62572;
  assign n4765 = ~pi392 & n4751;
  assign n4766 = ~n62523 & ~n4765;
  assign n4767 = ~n4764 & n4766;
  assign n4768 = ~n62523 & ~n4763;
  assign n4769 = pi591 & ~n62574;
  assign n4770 = pi591 & ~n62573;
  assign n4771 = ~n62574 & n4770;
  assign n4772 = ~n62573 & n4769;
  assign n4773 = ~pi590 & ~n62575;
  assign n4774 = ~n62571 & n4773;
  assign n4775 = ~pi591 & ~n62482;
  assign n4776 = ~pi591 & ~n62483;
  assign n4777 = ~n62482 & n4776;
  assign n4778 = ~n62483 & n4775;
  assign n4779 = pi591 & ~n3135;
  assign n4780 = pi590 & ~n4779;
  assign n4781 = ~n62576 & n4780;
  assign n4782 = ~n3318 & ~n4781;
  assign n4783 = ~n4774 & n4782;
  assign n4784 = ~n3318 & ~n4774;
  assign n4785 = ~n4781 & n4784;
  assign n4786 = ~n4164 & n4697;
  assign n4787 = ~n3341 & ~n4032;
  assign n4788 = ~n3341 & ~n4041;
  assign n4789 = n4043 & ~n4788;
  assign n4790 = ~n3341 & ~n4036;
  assign n4791 = n4038 & ~n4790;
  assign n4792 = ~n4789 & ~n4791;
  assign n4793 = n3957 & ~n4792;
  assign n4794 = ~pi592 & ~n3341;
  assign n4795 = ~n3821 & ~n4794;
  assign n4796 = ~n3957 & n4795;
  assign n4797 = ~n4793 & ~n4796;
  assign n4798 = pi1199 & n4797;
  assign n4799 = n3341 & ~n62498;
  assign n4800 = n62498 & n4795;
  assign n4801 = ~n4799 & ~n4800;
  assign n4802 = n62489 & ~n4801;
  assign n4803 = ~pi1196 & ~n62498;
  assign n4804 = n4795 & ~n4803;
  assign n4805 = ~pi1196 & n4799;
  assign n4806 = ~n4804 & ~n4805;
  assign n4807 = ~n62489 & ~n4806;
  assign n4808 = ~pi1199 & ~n4807;
  assign n4809 = ~pi1199 & ~n4802;
  assign n4810 = ~n4807 & n4809;
  assign n4811 = ~n4802 & n4808;
  assign n4812 = ~n4798 & ~n62578;
  assign n4813 = ~n4033 & ~n4787;
  assign n4814 = ~n62519 & n62579;
  assign n4815 = ~pi1198 & ~n62579;
  assign n4816 = pi1198 & ~n4795;
  assign n4817 = ~pi1198 & n62578;
  assign n4818 = ~pi1198 & pi1199;
  assign n4819 = n4797 & n4818;
  assign n4820 = ~n4816 & ~n4819;
  assign n4821 = ~n4817 & n4820;
  assign n4822 = ~n4815 & ~n4816;
  assign n4823 = n62519 & n62580;
  assign n4824 = ~pi374 & ~n62579;
  assign n4825 = pi374 & ~n62580;
  assign n4826 = ~n4824 & ~n4825;
  assign n4827 = ~pi369 & ~n4826;
  assign n4828 = ~pi374 & ~n62580;
  assign n4829 = pi374 & ~n62579;
  assign n4830 = ~n4828 & ~n4829;
  assign n4831 = pi369 & ~n4830;
  assign n4832 = ~n4827 & ~n4831;
  assign n4833 = ~n4814 & ~n4823;
  assign n4834 = n62517 & n62581;
  assign n4835 = n62519 & n62579;
  assign n4836 = ~n62519 & n62580;
  assign n4837 = pi369 & ~n4826;
  assign n4838 = ~pi369 & ~n4830;
  assign n4839 = ~n4837 & ~n4838;
  assign n4840 = ~n4835 & ~n4836;
  assign n4841 = ~n62517 & n62582;
  assign n4842 = ~n62517 & ~n62582;
  assign n4843 = n62517 & ~n62581;
  assign n4844 = ~n4842 & ~n4843;
  assign n4845 = ~pi370 & ~n62582;
  assign n4846 = pi370 & ~n62581;
  assign n4847 = ~n4845 & ~n4846;
  assign n4848 = pi370 & n62581;
  assign n4849 = ~pi370 & n62582;
  assign n4850 = ~pi371 & ~n4849;
  assign n4851 = ~n4848 & n4850;
  assign n4852 = ~pi371 & ~n4847;
  assign n4853 = ~pi370 & ~n62581;
  assign n4854 = pi370 & ~n62582;
  assign n4855 = ~n4853 & ~n4854;
  assign n4856 = pi370 & n62582;
  assign n4857 = ~pi370 & n62581;
  assign n4858 = pi371 & ~n4857;
  assign n4859 = ~n4856 & n4858;
  assign n4860 = pi371 & ~n4855;
  assign n4861 = ~n62584 & ~n62585;
  assign n4862 = ~n4834 & ~n4841;
  assign n4863 = pi373 & ~n62583;
  assign n4864 = ~n62517 & n62581;
  assign n4865 = n62517 & n62582;
  assign n4866 = ~pi371 & ~n4855;
  assign n4867 = pi371 & ~n4847;
  assign n4868 = ~n4866 & ~n4867;
  assign n4869 = ~n4864 & ~n4865;
  assign n4870 = ~pi373 & ~n62586;
  assign n4871 = n62514 & ~n4870;
  assign n4872 = n62514 & ~n4863;
  assign n4873 = ~n4870 & n4872;
  assign n4874 = ~n4863 & n4871;
  assign n4875 = pi373 & ~n62586;
  assign n4876 = ~pi373 & ~n62583;
  assign n4877 = ~n62514 & ~n4876;
  assign n4878 = ~n4875 & n4877;
  assign n4879 = ~pi590 & ~n4878;
  assign n4880 = ~n62587 & n4879;
  assign n4881 = ~n3343 & ~n3615;
  assign n4882 = n3341 & ~n62473;
  assign n4883 = n3691 & ~n4882;
  assign n4884 = n3343 & n62464;
  assign n4885 = n3341 & ~n62464;
  assign n4886 = ~pi455 & n3343;
  assign n4887 = pi455 & n3341;
  assign n4888 = ~pi452 & ~n4887;
  assign n4889 = ~pi455 & ~n3343;
  assign n4890 = pi455 & ~n3341;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = ~pi452 & ~n4891;
  assign n4893 = ~n4886 & n4888;
  assign n4894 = pi455 & n3343;
  assign n4895 = ~pi455 & n3341;
  assign n4896 = pi452 & ~n4895;
  assign n4897 = pi455 & ~n3343;
  assign n4898 = ~pi455 & ~n3341;
  assign n4899 = ~n4897 & ~n4898;
  assign n4900 = pi452 & ~n4899;
  assign n4901 = ~n4894 & n4896;
  assign n4902 = ~n62588 & ~n62589;
  assign n4903 = ~n4884 & ~n4885;
  assign n4904 = ~pi355 & ~n62590;
  assign n4905 = n3341 & n62464;
  assign n4906 = n3343 & ~n62464;
  assign n4907 = ~pi452 & ~n4899;
  assign n4908 = pi452 & ~n4891;
  assign n4909 = ~n4907 & ~n4908;
  assign n4910 = ~n3343 & ~n62464;
  assign n4911 = ~n3341 & n62464;
  assign n4912 = ~n4910 & ~n4911;
  assign n4913 = ~n4905 & ~n4906;
  assign n4914 = pi355 & ~n62591;
  assign n4915 = pi355 & n62591;
  assign n4916 = ~pi355 & n62590;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = ~n4904 & ~n4914;
  assign n4919 = pi458 & n62592;
  assign n4920 = ~pi355 & ~n62591;
  assign n4921 = pi355 & ~n62590;
  assign n4922 = ~pi355 & n62591;
  assign n4923 = pi355 & n62590;
  assign n4924 = ~n4922 & ~n4923;
  assign n4925 = ~n4920 & ~n4921;
  assign n4926 = ~pi458 & n62593;
  assign n4927 = n62462 & ~n4926;
  assign n4928 = n62462 & ~n4919;
  assign n4929 = ~n4926 & n4928;
  assign n4930 = ~n4919 & n4927;
  assign n4931 = pi458 & n62593;
  assign n4932 = ~pi458 & n62592;
  assign n4933 = ~n62462 & ~n4932;
  assign n4934 = ~n62462 & ~n4931;
  assign n4935 = ~n4932 & n4934;
  assign n4936 = ~n4931 & n4933;
  assign n4937 = pi1196 & ~n62595;
  assign n4938 = pi1196 & ~n62594;
  assign n4939 = ~n62595 & n4938;
  assign n4940 = ~n62594 & n4937;
  assign n4941 = ~pi1198 & ~n3380;
  assign n4942 = ~n62596 & n4941;
  assign n4943 = ~n3341 & ~n3702;
  assign n4944 = n3704 & ~n4943;
  assign n4945 = ~n3341 & ~n3697;
  assign n4946 = n3699 & ~n4945;
  assign n4947 = ~n3614 & ~n4946;
  assign n4948 = ~n3614 & ~n4944;
  assign n4949 = ~n4946 & n4948;
  assign n4950 = ~n4944 & n4947;
  assign n4951 = ~n3343 & n3614;
  assign n4952 = pi1198 & ~n4951;
  assign n4953 = ~n62597 & n4952;
  assign n4954 = ~n62460 & ~n4953;
  assign n4955 = ~n4942 & n4954;
  assign n4956 = ~n3343 & n62460;
  assign n4957 = ~n4955 & ~n4956;
  assign n4958 = ~n4942 & ~n4953;
  assign n4959 = ~n62460 & ~n4958;
  assign n4960 = n3343 & n62460;
  assign n4961 = ~n4959 & ~n4960;
  assign n4962 = ~n4881 & ~n4883;
  assign n4963 = ~n3478 & ~n62598;
  assign n4964 = pi1199 & ~n3343;
  assign n4965 = ~pi351 & n4964;
  assign n4966 = ~n4963 & ~n4965;
  assign n4967 = pi461 & ~n4966;
  assign n4968 = pi356 & ~pi357;
  assign n4969 = ~pi356 & pi357;
  assign n4970 = ~pi356 & ~pi357;
  assign n4971 = pi356 & pi357;
  assign n4972 = ~n4970 & ~n4971;
  assign n4973 = ~n4968 & ~n4969;
  assign n4974 = ~n62481 & ~n62599;
  assign n4975 = n62481 & n62599;
  assign n4976 = pi356 & ~n62481;
  assign n4977 = ~pi356 & n62481;
  assign n4978 = ~n4976 & ~n4977;
  assign n4979 = pi357 & ~n4978;
  assign n4980 = ~pi357 & n4978;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = ~n4974 & ~n4975;
  assign n4983 = ~n3767 & ~n62598;
  assign n4984 = pi351 & n4964;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = ~pi461 & ~n4985;
  assign n4987 = n62600 & ~n4986;
  assign n4988 = ~n4967 & n4987;
  assign n4989 = pi461 & ~n4985;
  assign n4990 = ~pi461 & ~n4966;
  assign n4991 = ~n62600 & ~n4990;
  assign n4992 = ~n4989 & n4991;
  assign n4993 = pi590 & ~n4992;
  assign n4994 = ~n4988 & n4993;
  assign n4995 = ~n4880 & ~n4994;
  assign n4996 = ~pi591 & ~n4995;
  assign n4997 = n3343 & n4621;
  assign n4998 = ~pi75 & ~pi592;
  assign n4999 = ~n3339 & ~n4998;
  assign n5000 = ~pi1196 & ~n3338;
  assign n5001 = n3328 & ~n62530;
  assign n5002 = n2992 & ~n5001;
  assign n5003 = n3004 & ~n5002;
  assign n5004 = n62421 & ~n62530;
  assign n5005 = n3032 & ~n5004;
  assign n5006 = pi87 & n3334;
  assign n5007 = n62407 & ~n3333;
  assign n5008 = ~n5005 & n62601;
  assign n5009 = n4998 & ~n5008;
  assign n5010 = ~n5003 & n5009;
  assign n5011 = pi1196 & ~n5010;
  assign n5012 = ~pi1199 & ~n5011;
  assign n5013 = pi1196 & n4998;
  assign n5014 = ~n5008 & n5013;
  assign n5015 = ~n5003 & n5014;
  assign n5016 = ~pi1196 & n3338;
  assign n5017 = ~n5015 & ~n5016;
  assign n5018 = ~pi1199 & ~n5017;
  assign n5019 = ~n5000 & n5012;
  assign n5020 = pi1196 & n62530;
  assign n5021 = ~pi75 & n5020;
  assign n5022 = n62535 & ~n5021;
  assign n5023 = n3328 & n5022;
  assign n5024 = n2992 & ~n5023;
  assign n5025 = n3004 & ~n5024;
  assign n5026 = n62535 & ~n5020;
  assign n5027 = n62421 & n5026;
  assign n5028 = n3032 & ~n5027;
  assign n5029 = n62421 & n62535;
  assign n5030 = n3032 & ~n5029;
  assign n5031 = n62601 & ~n5030;
  assign n5032 = pi1196 & n5005;
  assign n5033 = n5031 & ~n5032;
  assign n5034 = n62601 & ~n5028;
  assign n5035 = pi1199 & n4998;
  assign n5036 = ~n5005 & n5031;
  assign n5037 = ~pi1196 & n5031;
  assign n5038 = n5035 & ~n5037;
  assign n5039 = ~n5036 & n5038;
  assign n5040 = n5035 & ~n5036;
  assign n5041 = ~n5037 & n5040;
  assign n5042 = ~n62603 & n5035;
  assign n5043 = ~n5025 & n62604;
  assign n5044 = ~n62602 & ~n5043;
  assign n5045 = ~n4999 & ~n5043;
  assign n5046 = ~n62602 & n5045;
  assign n5047 = ~n4999 & n5044;
  assign n5048 = pi567 & ~n62605;
  assign n5049 = n2804 & ~n4621;
  assign n5050 = ~n5048 & n5049;
  assign n5051 = ~n4997 & ~n5050;
  assign n5052 = ~n4210 & n5051;
  assign n5053 = pi1197 & ~n3343;
  assign n5054 = ~pi333 & n5053;
  assign n5055 = ~pi1197 & n5051;
  assign n5056 = ~n5053 & ~n5055;
  assign n5057 = ~pi333 & ~n5056;
  assign n5058 = pi333 & n5051;
  assign n5059 = ~n5057 & ~n5058;
  assign n5060 = pi333 & ~n5051;
  assign n5061 = ~pi333 & n5056;
  assign n5062 = ~n5060 & ~n5061;
  assign n5063 = ~n5052 & ~n5054;
  assign n5064 = n62523 & n62606;
  assign n5065 = ~pi391 & ~pi392;
  assign n5066 = pi391 & pi392;
  assign n5067 = ~n5065 & ~n5066;
  assign n5068 = ~n4681 & n5051;
  assign n5069 = pi333 & n5053;
  assign n5070 = pi333 & ~n5056;
  assign n5071 = ~pi333 & n5051;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = ~n5068 & ~n5069;
  assign n5074 = ~n62523 & n62607;
  assign n5075 = ~n5067 & ~n5074;
  assign n5076 = ~n5064 & n5075;
  assign n5077 = n62523 & n62607;
  assign n5078 = ~n62523 & n62606;
  assign n5079 = n5067 & ~n5078;
  assign n5080 = ~n5077 & n5079;
  assign n5081 = ~pi590 & ~n5080;
  assign n5082 = ~n5076 & n5081;
  assign n5083 = pi590 & n3341;
  assign n5084 = pi591 & ~n5083;
  assign n5085 = ~n5082 & n5084;
  assign n5086 = n3318 & ~n5085;
  assign n5087 = ~n4989 & ~n4990;
  assign n5088 = ~pi357 & ~n5087;
  assign n5089 = ~n4967 & ~n4986;
  assign n5090 = pi357 & ~n5089;
  assign n5091 = ~n5088 & ~n5090;
  assign n5092 = n4978 & ~n5091;
  assign n5093 = ~pi357 & ~n5089;
  assign n5094 = pi357 & ~n5087;
  assign n5095 = ~n5093 & ~n5094;
  assign n5096 = ~n4978 & ~n5095;
  assign n5097 = ~pi591 & ~n5096;
  assign n5098 = ~pi356 & ~n5091;
  assign n5099 = pi356 & ~n5095;
  assign n5100 = ~n5098 & ~n5099;
  assign n5101 = pi356 & n5095;
  assign n5102 = ~pi356 & n5091;
  assign n5103 = ~n62481 & ~n5102;
  assign n5104 = ~n5101 & n5103;
  assign n5105 = ~n62481 & ~n5100;
  assign n5106 = ~pi356 & ~n5095;
  assign n5107 = pi356 & ~n5091;
  assign n5108 = ~n5106 & ~n5107;
  assign n5109 = pi356 & n5091;
  assign n5110 = ~pi356 & n5095;
  assign n5111 = n62481 & ~n5110;
  assign n5112 = ~n5109 & n5111;
  assign n5113 = n62481 & ~n5108;
  assign n5114 = ~pi591 & ~n62609;
  assign n5115 = ~n62608 & n5114;
  assign n5116 = ~pi591 & ~n62608;
  assign n5117 = ~n62609 & n5116;
  assign n5118 = ~n5092 & n5097;
  assign n5119 = pi591 & n3341;
  assign n5120 = pi590 & ~n5119;
  assign n5121 = ~n62610 & n5120;
  assign n5122 = pi373 & n62586;
  assign n5123 = ~pi373 & n62583;
  assign n5124 = ~n5122 & ~n5123;
  assign n5125 = ~n4875 & ~n4876;
  assign n5126 = ~pi375 & ~n62611;
  assign n5127 = ~pi373 & n62586;
  assign n5128 = pi373 & n62583;
  assign n5129 = ~n5127 & ~n5128;
  assign n5130 = ~n4863 & ~n4870;
  assign n5131 = pi375 & ~n62612;
  assign n5132 = n4100 & ~n5131;
  assign n5133 = n4100 & ~n5126;
  assign n5134 = ~n5131 & n5133;
  assign n5135 = ~n5126 & n5132;
  assign n5136 = pi375 & ~n62611;
  assign n5137 = ~pi375 & ~n62612;
  assign n5138 = ~n4100 & ~n5137;
  assign n5139 = ~n4100 & ~n5136;
  assign n5140 = ~n5137 & n5139;
  assign n5141 = ~n5136 & n5138;
  assign n5142 = ~pi591 & ~n62614;
  assign n5143 = ~pi591 & ~n62613;
  assign n5144 = ~n62614 & n5143;
  assign n5145 = ~n62613 & n5142;
  assign n5146 = pi391 & ~n62607;
  assign n5147 = ~pi391 & ~n62606;
  assign n5148 = ~n5146 & ~n5147;
  assign n5149 = ~pi392 & ~n5148;
  assign n5150 = ~pi391 & ~n62607;
  assign n5151 = pi391 & ~n62606;
  assign n5152 = ~n5150 & ~n5151;
  assign n5153 = pi392 & ~n5152;
  assign n5154 = ~n5149 & ~n5153;
  assign n5155 = ~pi393 & ~n5154;
  assign n5156 = ~pi392 & ~n5152;
  assign n5157 = pi392 & ~n5148;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = pi393 & ~n5158;
  assign n5160 = ~n5155 & ~n5159;
  assign n5161 = ~pi334 & n5160;
  assign n5162 = ~pi393 & ~n5158;
  assign n5163 = pi393 & ~n5154;
  assign n5164 = ~n5162 & ~n5163;
  assign n5165 = pi334 & n5164;
  assign n5166 = ~n62521 & ~n5165;
  assign n5167 = ~n62521 & ~n5161;
  assign n5168 = ~n5165 & n5167;
  assign n5169 = ~n5161 & n5166;
  assign n5170 = ~pi334 & n5164;
  assign n5171 = pi334 & n5160;
  assign n5172 = n62521 & ~n5171;
  assign n5173 = n62521 & ~n5170;
  assign n5174 = ~n5171 & n5173;
  assign n5175 = ~n5170 & n5172;
  assign n5176 = pi591 & ~n62617;
  assign n5177 = pi591 & ~n62616;
  assign n5178 = ~n62617 & n5177;
  assign n5179 = ~n62616 & n5176;
  assign n5180 = ~pi590 & ~n62618;
  assign n5181 = ~n62616 & ~n62617;
  assign n5182 = pi591 & ~n5181;
  assign n5183 = ~pi591 & ~n4878;
  assign n5184 = ~n62587 & n5183;
  assign n5185 = ~n5182 & ~n5184;
  assign n5186 = ~pi590 & ~n5185;
  assign n5187 = ~n62615 & n5180;
  assign n5188 = n3318 & ~n62619;
  assign n5189 = ~n5121 & n5188;
  assign n5190 = ~n4996 & n5086;
  assign n5191 = ~pi588 & ~n62620;
  assign n5192 = ~pi588 & ~n62577;
  assign n5193 = ~n62620 & n5192;
  assign n5194 = ~n62577 & n5191;
  assign n5195 = n62455 & ~n62621;
  assign n5196 = ~n3469 & n62455;
  assign n5197 = ~n62621 & n5196;
  assign n5198 = ~n3469 & n5195;
  assign n5199 = ~pi333 & ~n4209;
  assign n5200 = pi333 & n4209;
  assign n5201 = pi1197 & ~n5200;
  assign n5202 = pi1197 & ~n5199;
  assign n5203 = ~n5200 & n5202;
  assign n5204 = ~n5199 & n5201;
  assign n5205 = ~n4621 & ~n62623;
  assign n5206 = n62558 & n4681;
  assign n5207 = ~n4209 & n5206;
  assign n5208 = pi1199 & ~n62535;
  assign n5209 = n3132 & ~n5020;
  assign n5210 = ~n5208 & n5209;
  assign n5211 = ~n5207 & ~n5210;
  assign n5212 = n5205 & ~n5211;
  assign n5213 = pi592 & n3132;
  assign n5214 = pi591 & ~n5213;
  assign n5215 = ~n5205 & ~n5213;
  assign n5216 = pi1199 & ~n5213;
  assign n5217 = ~pi592 & ~n5020;
  assign n5218 = ~pi592 & n4538;
  assign n5219 = ~n5020 & n5218;
  assign n5220 = n4538 & n5217;
  assign n5221 = n5216 & ~n62624;
  assign n5222 = n4494 & n4495;
  assign n5223 = n3132 & ~n4494;
  assign n5224 = ~pi1199 & ~n5223;
  assign n5225 = ~n5222 & n5224;
  assign n5226 = ~n5221 & ~n5225;
  assign n5227 = ~n5207 & ~n5226;
  assign n5228 = pi1197 & ~n5213;
  assign n5229 = ~pi1197 & ~n5226;
  assign n5230 = ~n5228 & ~n5229;
  assign n5231 = pi333 & ~n5230;
  assign n5232 = pi1198 & ~n5213;
  assign n5233 = n5226 & ~n5232;
  assign n5234 = ~n62558 & ~n5233;
  assign n5235 = ~pi333 & ~n5226;
  assign n5236 = ~n5234 & ~n5235;
  assign n5237 = ~n5231 & n5236;
  assign n5238 = ~pi391 & ~n5237;
  assign n5239 = ~pi333 & ~n5230;
  assign n5240 = n5226 & ~n5234;
  assign n5241 = ~n5239 & n5240;
  assign n5242 = pi391 & ~n5241;
  assign n5243 = ~n5238 & ~n5242;
  assign n5244 = ~pi392 & ~n5243;
  assign n5245 = ~pi391 & ~n5241;
  assign n5246 = pi391 & ~n5237;
  assign n5247 = ~n5245 & ~n5246;
  assign n5248 = pi392 & ~n5247;
  assign n5249 = ~n5244 & ~n5248;
  assign n5250 = ~pi393 & ~n5249;
  assign n5251 = ~pi392 & ~n5247;
  assign n5252 = pi392 & ~n5243;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = pi393 & ~n5253;
  assign n5255 = ~n62522 & ~n5254;
  assign n5256 = ~n62522 & ~n5250;
  assign n5257 = ~n5254 & n5256;
  assign n5258 = ~n5250 & n5255;
  assign n5259 = ~pi393 & ~n5253;
  assign n5260 = pi393 & ~n5249;
  assign n5261 = n62522 & ~n5260;
  assign n5262 = n62522 & ~n5259;
  assign n5263 = ~n5260 & n5262;
  assign n5264 = ~n5259 & n5261;
  assign n5265 = ~n62625 & ~n62626;
  assign n5266 = ~n62523 & ~n5244;
  assign n5267 = ~n5248 & n5266;
  assign n5268 = n62523 & ~n5251;
  assign n5269 = ~n5252 & n5268;
  assign n5270 = ~n5267 & ~n5269;
  assign n5271 = ~n5215 & ~n5227;
  assign n5272 = pi591 & n62627;
  assign n5273 = ~n5212 & n5214;
  assign n5274 = pi592 & ~n3957;
  assign n5275 = n3957 & n62505;
  assign n5276 = pi592 & ~n5275;
  assign n5277 = n3132 & ~n5276;
  assign n5278 = pi1199 & ~n5277;
  assign n5279 = ~n5274 & ~n5278;
  assign n5280 = ~n62518 & n62519;
  assign n5281 = n62518 & ~n62519;
  assign n5282 = pi1198 & ~n5281;
  assign n5283 = ~n5280 & n5282;
  assign n5284 = n5213 & ~n5283;
  assign n5285 = ~pi592 & n3132;
  assign n5286 = n5213 & n5279;
  assign n5287 = ~pi1198 & n5286;
  assign n5288 = ~pi370 & ~n62519;
  assign n5289 = pi370 & n62519;
  assign n5290 = ~n5288 & ~n5289;
  assign n5291 = ~pi371 & ~n5290;
  assign n5292 = pi371 & n5290;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~pi373 & ~n5293;
  assign n5295 = pi373 & n5293;
  assign n5296 = ~n5294 & ~n5295;
  assign n5297 = pi375 & ~n5296;
  assign n5298 = ~pi375 & n5296;
  assign n5299 = ~n5297 & ~n5298;
  assign n5300 = ~n4100 & ~n5299;
  assign n5301 = n4100 & n5299;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = n5286 & n5302;
  assign n5304 = ~n5285 & ~n5303;
  assign n5305 = ~n5285 & ~n5287;
  assign n5306 = ~n5303 & n5305;
  assign n5307 = ~n5287 & n5304;
  assign n5308 = ~n5285 & ~n62629;
  assign n5309 = n5279 & n5284;
  assign n5310 = ~pi591 & ~n5285;
  assign n5311 = ~n62630 & n5310;
  assign n5312 = ~n62628 & ~n5311;
  assign n5313 = ~pi590 & ~n5312;
  assign n5314 = ~pi592 & n62466;
  assign n5315 = n3132 & ~n5314;
  assign n5316 = n3132 & ~n3561;
  assign n5317 = ~n5314 & n5316;
  assign n5318 = pi361 & ~pi458;
  assign n5319 = ~pi361 & pi458;
  assign n5320 = ~n5318 & ~n5319;
  assign n5321 = n3609 & n5320;
  assign n5322 = ~n3609 & ~n5320;
  assign n5323 = pi355 & ~pi361;
  assign n5324 = ~pi355 & pi361;
  assign n5325 = ~n5323 & ~n5324;
  assign n5326 = pi458 & ~n62464;
  assign n5327 = ~pi458 & n62464;
  assign n5328 = ~n5326 & ~n5327;
  assign n5329 = n5325 & n5328;
  assign n5330 = ~n5325 & ~n5328;
  assign n5331 = ~n5329 & ~n5330;
  assign n5332 = ~n5321 & ~n5322;
  assign n5333 = ~pi441 & ~n62631;
  assign n5334 = pi441 & n62631;
  assign n5335 = ~pi592 & ~n5334;
  assign n5336 = ~pi592 & ~n5333;
  assign n5337 = ~n5334 & n5336;
  assign n5338 = ~n5333 & n5335;
  assign n5339 = n3132 & n3561;
  assign n5340 = ~n62632 & n5339;
  assign n5341 = pi1196 & ~n5340;
  assign n5342 = ~n5317 & n5341;
  assign n5343 = pi1196 & ~n5315;
  assign n5344 = ~pi1198 & ~n62633;
  assign n5345 = ~n3614 & n62472;
  assign n5346 = pi1198 & n5285;
  assign n5347 = n62472 & n5285;
  assign n5348 = n3707 & n5347;
  assign n5349 = n5345 & n5346;
  assign n5350 = ~n5344 & ~n62634;
  assign n5351 = ~n62460 & ~n5350;
  assign n5352 = ~pi592 & ~n5351;
  assign n5353 = n3132 & ~n5352;
  assign n5354 = ~n3478 & ~n5353;
  assign n5355 = ~pi351 & n5216;
  assign n5356 = pi461 & ~n62599;
  assign n5357 = ~pi461 & n62599;
  assign n5358 = ~n5356 & ~n5357;
  assign n5359 = n62481 & n5358;
  assign n5360 = ~n62481 & ~n5358;
  assign n5361 = pi461 & ~n62481;
  assign n5362 = ~pi461 & n62481;
  assign n5363 = ~n5361 & ~n5362;
  assign n5364 = n62599 & n5363;
  assign n5365 = ~n62599 & ~n5363;
  assign n5366 = ~n5364 & ~n5365;
  assign n5367 = ~n5359 & ~n5360;
  assign n5368 = ~n5355 & n62635;
  assign n5369 = ~n5354 & n5368;
  assign n5370 = ~n3767 & ~n5353;
  assign n5371 = pi351 & n5216;
  assign n5372 = ~n62635 & ~n5371;
  assign n5373 = ~n5370 & n5372;
  assign n5374 = ~n5370 & ~n5371;
  assign n5375 = ~pi461 & ~n5374;
  assign n5376 = ~n5354 & ~n5355;
  assign n5377 = pi461 & ~n5376;
  assign n5378 = ~n5375 & ~n5377;
  assign n5379 = ~pi357 & ~n5378;
  assign n5380 = ~pi461 & ~n5376;
  assign n5381 = pi461 & ~n5374;
  assign n5382 = ~n5380 & ~n5381;
  assign n5383 = pi357 & ~n5382;
  assign n5384 = ~n5379 & ~n5383;
  assign n5385 = ~pi356 & ~n5384;
  assign n5386 = ~pi357 & ~n5382;
  assign n5387 = pi357 & ~n5378;
  assign n5388 = ~n5386 & ~n5387;
  assign n5389 = pi356 & ~n5388;
  assign n5390 = n62481 & ~n5389;
  assign n5391 = n62481 & ~n5385;
  assign n5392 = ~n5389 & n5391;
  assign n5393 = ~n5385 & n5390;
  assign n5394 = ~pi356 & ~n5388;
  assign n5395 = pi356 & ~n5384;
  assign n5396 = ~n62481 & ~n5395;
  assign n5397 = ~n62481 & ~n5394;
  assign n5398 = ~n5395 & n5397;
  assign n5399 = ~n5394 & n5396;
  assign n5400 = ~n62636 & ~n62637;
  assign n5401 = ~n5369 & ~n5373;
  assign n5402 = ~pi591 & ~n62638;
  assign n5403 = pi591 & n3132;
  assign n5404 = pi590 & ~n5403;
  assign n5405 = ~n5402 & n5404;
  assign n5406 = pi461 & n5374;
  assign n5407 = ~pi461 & n5376;
  assign n5408 = ~n62600 & ~n5407;
  assign n5409 = ~n5406 & n5408;
  assign n5410 = pi461 & n5376;
  assign n5411 = ~pi461 & n5374;
  assign n5412 = n62600 & ~n5411;
  assign n5413 = ~n5410 & n5412;
  assign n5414 = pi590 & ~n5413;
  assign n5415 = ~n5409 & n5414;
  assign n5416 = pi590 & ~n62638;
  assign n5417 = ~pi590 & ~n62629;
  assign n5418 = ~pi591 & ~n5417;
  assign n5419 = ~n62639 & n5418;
  assign n5420 = ~pi590 & ~n62627;
  assign n5421 = pi590 & n3132;
  assign n5422 = pi591 & ~n5421;
  assign n5423 = ~n5420 & n5422;
  assign n5424 = ~n5419 & ~n5423;
  assign n5425 = ~n5313 & ~n5405;
  assign n5426 = ~pi588 & ~n62640;
  assign n5427 = ~n3318 & ~n62455;
  assign n5428 = pi436 & ~pi443;
  assign n5429 = ~pi436 & pi443;
  assign n5430 = ~pi436 & ~pi443;
  assign n5431 = pi436 & pi443;
  assign n5432 = ~n5430 & ~n5431;
  assign n5433 = ~n5428 & ~n5429;
  assign n5434 = ~pi444 & ~n62641;
  assign n5435 = pi444 & n62641;
  assign n5436 = ~n5434 & ~n5435;
  assign n5437 = n62425 & n5436;
  assign n5438 = ~n62425 & ~n5436;
  assign n5439 = n4494 & ~n5438;
  assign n5440 = n4494 & ~n5437;
  assign n5441 = ~n5438 & n5440;
  assign n5442 = ~n5437 & n5439;
  assign n5443 = n2578 & ~n62642;
  assign n5444 = n62331 & n3269;
  assign n5445 = ~n62331 & ~n3269;
  assign n5446 = pi426 & n3269;
  assign n5447 = ~pi426 & ~n3269;
  assign n5448 = pi426 & ~n3269;
  assign n5449 = ~pi426 & n3269;
  assign n5450 = ~n5448 & ~n5449;
  assign n5451 = ~n5446 & ~n5447;
  assign n5452 = pi430 & ~n62643;
  assign n5453 = ~pi430 & n62643;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = ~n5444 & ~n5445;
  assign n5456 = n62332 & ~n62450;
  assign n5457 = ~n62332 & n62450;
  assign n5458 = pi445 & n62332;
  assign n5459 = ~pi445 & ~n62332;
  assign n5460 = ~n5458 & ~n5459;
  assign n5461 = pi448 & ~n5460;
  assign n5462 = ~pi448 & n5460;
  assign n5463 = ~n5461 & ~n5462;
  assign n5464 = ~n5456 & ~n5457;
  assign n5465 = n62644 & n62645;
  assign n5466 = ~n62644 & ~n62645;
  assign n5467 = pi1199 & ~n5466;
  assign n5468 = n62450 & n62644;
  assign n5469 = ~n62450 & ~n62644;
  assign n5470 = ~n5468 & ~n5469;
  assign n5471 = n62332 & ~n5470;
  assign n5472 = ~n62332 & n5470;
  assign n5473 = pi1199 & ~n5472;
  assign n5474 = ~n5471 & n5473;
  assign n5475 = ~n5465 & n5467;
  assign n5476 = n3312 & n5285;
  assign n5477 = ~n62646 & n5476;
  assign n5478 = n5443 & n5476;
  assign n5479 = ~n62646 & n5478;
  assign n5480 = n5443 & n5477;
  assign n5481 = ~pi592 & n3312;
  assign n5482 = n3132 & ~n5481;
  assign n5483 = pi588 & ~n5482;
  assign n5484 = n5285 & n5443;
  assign n5485 = n62331 & n62645;
  assign n5486 = ~n62331 & ~n62645;
  assign n5487 = pi430 & n62332;
  assign n5488 = ~pi430 & ~n62332;
  assign n5489 = ~n5487 & ~n5488;
  assign n5490 = ~pi426 & ~n5489;
  assign n5491 = pi426 & n5489;
  assign n5492 = ~n5490 & ~n5491;
  assign n5493 = ~pi445 & ~n5492;
  assign n5494 = pi445 & n5492;
  assign n5495 = ~n5493 & ~n5494;
  assign n5496 = ~pi448 & ~n5495;
  assign n5497 = pi448 & n5495;
  assign n5498 = ~n5496 & ~n5497;
  assign n5499 = ~n5485 & ~n5486;
  assign n5500 = n5484 & ~n62648;
  assign n5501 = ~n5213 & ~n5500;
  assign n5502 = n3269 & ~n5501;
  assign n5503 = n5484 & n62648;
  assign n5504 = ~n5213 & ~n5503;
  assign n5505 = ~n3269 & ~n5504;
  assign n5506 = pi1199 & ~n5505;
  assign n5507 = pi1199 & ~n5502;
  assign n5508 = ~n5505 & n5507;
  assign n5509 = ~n5502 & n5506;
  assign n5510 = ~pi1199 & ~n5213;
  assign n5511 = ~n5484 & n5510;
  assign n5512 = n3312 & ~n5511;
  assign n5513 = ~n62649 & n5512;
  assign n5514 = n3132 & ~n3312;
  assign n5515 = pi588 & ~n5514;
  assign n5516 = ~n5513 & n5515;
  assign n5517 = ~n62647 & n5483;
  assign n5518 = n5427 & ~n62650;
  assign n5519 = ~n5426 & n5518;
  assign n5520 = ~pi217 & ~n5519;
  assign n5521 = ~n62622 & n5520;
  assign n5522 = n3318 & ~n3341;
  assign n5523 = n3135 & ~n3318;
  assign n5524 = n62455 & ~n5523;
  assign n5525 = ~n5522 & n5524;
  assign n5526 = n3132 & n5427;
  assign n5527 = pi217 & ~n5526;
  assign n5528 = ~n5525 & n5527;
  assign n5529 = ~pi1161 & ~pi1162;
  assign n5530 = ~pi1163 & n5529;
  assign n5531 = ~n5528 & n5530;
  assign n5532 = ~n5521 & n5531;
  assign n5533 = pi1161 & ~pi1163;
  assign n5534 = n2923 & n5533;
  assign n5535 = ~pi31 & pi1162;
  assign n5536 = n5534 & n5535;
  assign n5537 = ~n5532 & ~n5536;
  assign n5538 = pi98 & pi1092;
  assign n5539 = pi1093 & n5538;
  assign n5540 = ~pi567 & n2923;
  assign n5541 = ~n5539 & ~n5540;
  assign n5542 = pi591 & ~n5541;
  assign n5543 = pi590 & ~n5542;
  assign n5544 = n5345 & n5541;
  assign n5545 = pi592 & ~n5541;
  assign n5546 = ~pi88 & n2638;
  assign n5547 = ~pi58 & n2699;
  assign n5548 = ~pi110 & n2664;
  assign n5549 = n2698 & n5546;
  assign n5550 = n62651 & n5549;
  assign n5551 = n62361 & n5546;
  assign n5552 = n2689 & n62652;
  assign n5553 = n2696 & n5552;
  assign n5554 = n62381 & n3112;
  assign n5555 = n5553 & n5554;
  assign n5556 = ~pi98 & ~n5555;
  assign n5557 = pi1092 & ~n5556;
  assign n5558 = pi1091 & n5539;
  assign n5559 = n62373 & ~n5558;
  assign n5560 = pi87 & n5559;
  assign n5561 = n62407 & ~n5558;
  assign n5562 = ~n5557 & n62653;
  assign n5563 = n62407 & ~n5557;
  assign n5564 = pi51 & n5553;
  assign n5565 = pi90 & pi93;
  assign n5566 = ~pi841 & ~n2694;
  assign n5567 = ~n5565 & n5566;
  assign n5568 = n2743 & n5567;
  assign n5569 = n5552 & n5568;
  assign n5570 = ~n5564 & ~n5569;
  assign n5571 = n62366 & n3112;
  assign n5572 = ~n5570 & n5571;
  assign n5573 = ~pi98 & ~n5572;
  assign n5574 = pi1092 & ~n5573;
  assign n5575 = ~pi87 & n5559;
  assign n5576 = n2806 & ~n5558;
  assign n5577 = ~n5574 & n62655;
  assign n5578 = n2806 & ~n5574;
  assign n5579 = ~n62654 & ~n62656;
  assign n5580 = pi122 & ~n5579;
  assign n5581 = ~n3036 & ~n5539;
  assign n5582 = ~pi122 & n5581;
  assign n5583 = n3032 & ~n5582;
  assign n5584 = n62373 & ~n5583;
  assign n5585 = ~n5580 & ~n5584;
  assign n5586 = ~pi75 & ~n5558;
  assign n5587 = n5559 & ~n5583;
  assign n5588 = ~n5580 & ~n5587;
  assign n5589 = ~pi75 & ~n5588;
  assign n5590 = ~n5585 & n5586;
  assign n5591 = ~n62374 & n5581;
  assign n5592 = pi567 & n2580;
  assign n5593 = ~n5591 & n5592;
  assign n5594 = ~n62657 & n5593;
  assign n5595 = ~n2580 & ~n5581;
  assign n5596 = ~n5540 & ~n5595;
  assign n5597 = ~n5594 & n5596;
  assign n5598 = ~pi592 & ~n5597;
  assign n5599 = ~n5545 & ~n5598;
  assign n5600 = ~n5345 & n5599;
  assign n5601 = ~n5544 & ~n5600;
  assign n5602 = pi1198 & ~n5601;
  assign n5603 = ~pi1196 & ~n5541;
  assign n5604 = ~pi1198 & ~n5603;
  assign n5605 = n62464 & n5541;
  assign n5606 = ~n62464 & n5599;
  assign n5607 = ~n5605 & ~n5606;
  assign n5608 = pi355 & ~n5607;
  assign n5609 = pi455 & ~n5541;
  assign n5610 = ~pi455 & ~n5599;
  assign n5611 = ~n5609 & ~n5610;
  assign n5612 = ~pi452 & ~n5611;
  assign n5613 = ~pi455 & ~n5541;
  assign n5614 = pi455 & ~n5599;
  assign n5615 = ~n5613 & ~n5614;
  assign n5616 = pi452 & ~n5615;
  assign n5617 = ~n5612 & ~n5616;
  assign n5618 = ~pi355 & n5617;
  assign n5619 = ~n5608 & ~n5618;
  assign n5620 = ~pi458 & n5619;
  assign n5621 = ~pi355 & ~n5607;
  assign n5622 = pi355 & n5617;
  assign n5623 = ~n5621 & ~n5622;
  assign n5624 = pi458 & n5623;
  assign n5625 = ~n62462 & ~n5624;
  assign n5626 = ~n62462 & ~n5620;
  assign n5627 = ~n5624 & n5626;
  assign n5628 = ~n5620 & n5625;
  assign n5629 = pi458 & n5619;
  assign n5630 = ~pi458 & n5623;
  assign n5631 = n62462 & ~n5630;
  assign n5632 = n62462 & ~n5629;
  assign n5633 = ~n5630 & n5632;
  assign n5634 = ~n5629 & n5631;
  assign n5635 = pi1196 & ~n62659;
  assign n5636 = pi1196 & ~n62658;
  assign n5637 = ~n62659 & n5636;
  assign n5638 = ~n62658 & n5635;
  assign n5639 = n5604 & ~n62660;
  assign n5640 = ~n5602 & ~n5639;
  assign n5641 = ~n62460 & ~n5640;
  assign n5642 = n62460 & n5599;
  assign n5643 = ~n5641 & ~n5642;
  assign n5644 = ~n3478 & n5643;
  assign n5645 = pi1199 & ~n5599;
  assign n5646 = ~pi351 & n5645;
  assign n5647 = n62635 & ~n5646;
  assign n5648 = ~n5644 & n5647;
  assign n5649 = ~n3767 & n5643;
  assign n5650 = pi351 & n5645;
  assign n5651 = ~n62635 & ~n5650;
  assign n5652 = ~n5649 & n5651;
  assign n5653 = ~pi591 & ~n5652;
  assign n5654 = ~n5644 & ~n5646;
  assign n5655 = ~pi461 & ~n5654;
  assign n5656 = ~n5649 & ~n5650;
  assign n5657 = pi461 & ~n5656;
  assign n5658 = ~n5655 & ~n5657;
  assign n5659 = ~pi357 & ~n5658;
  assign n5660 = ~pi461 & ~n5656;
  assign n5661 = pi461 & ~n5654;
  assign n5662 = ~n5660 & ~n5661;
  assign n5663 = pi357 & ~n5662;
  assign n5664 = ~n5659 & ~n5663;
  assign n5665 = pi357 & n5662;
  assign n5666 = ~pi357 & n5658;
  assign n5667 = ~pi356 & ~n5666;
  assign n5668 = ~n5665 & n5667;
  assign n5669 = ~pi356 & ~n5664;
  assign n5670 = ~pi357 & ~n5662;
  assign n5671 = pi357 & ~n5658;
  assign n5672 = ~n5670 & ~n5671;
  assign n5673 = pi357 & n5658;
  assign n5674 = ~pi357 & n5662;
  assign n5675 = pi356 & ~n5674;
  assign n5676 = ~n5673 & n5675;
  assign n5677 = pi356 & ~n5672;
  assign n5678 = ~n62661 & ~n62662;
  assign n5679 = ~pi354 & ~n5678;
  assign n5680 = ~n62599 & n5662;
  assign n5681 = n62599 & n5658;
  assign n5682 = ~pi356 & ~n5672;
  assign n5683 = pi356 & ~n5664;
  assign n5684 = ~n5682 & ~n5683;
  assign n5685 = ~n5680 & ~n5681;
  assign n5686 = pi354 & ~n62663;
  assign n5687 = ~n62480 & ~n5686;
  assign n5688 = ~n62480 & ~n5679;
  assign n5689 = ~n5686 & n5688;
  assign n5690 = ~n5679 & n5687;
  assign n5691 = pi354 & ~n5678;
  assign n5692 = ~pi354 & ~n62663;
  assign n5693 = n62480 & ~n5692;
  assign n5694 = n62480 & ~n5691;
  assign n5695 = ~n5692 & n5694;
  assign n5696 = ~n5691 & n5693;
  assign n5697 = ~pi591 & ~n62665;
  assign n5698 = ~n62664 & n5697;
  assign n5699 = ~pi591 & ~n62664;
  assign n5700 = ~n62665 & n5699;
  assign n5701 = ~n5648 & n5653;
  assign n5702 = n5543 & ~n62666;
  assign n5703 = ~pi592 & ~n5541;
  assign n5704 = pi592 & ~n5597;
  assign n5705 = ~n5703 & ~n5704;
  assign n5706 = ~pi367 & ~n5705;
  assign n5707 = pi367 & ~n5541;
  assign n5708 = ~n5706 & ~n5707;
  assign n5709 = ~n62491 & ~n5708;
  assign n5710 = pi367 & ~n5705;
  assign n5711 = ~pi367 & ~n5541;
  assign n5712 = ~n5710 & ~n5711;
  assign n5713 = n62491 & ~n5712;
  assign n5714 = ~n5709 & ~n5713;
  assign n5715 = ~n62494 & ~n5714;
  assign n5716 = n62491 & ~n5708;
  assign n5717 = ~n62491 & ~n5712;
  assign n5718 = n62491 & n5708;
  assign n5719 = ~n62491 & n5712;
  assign n5720 = ~n5718 & ~n5719;
  assign n5721 = ~n5716 & ~n5717;
  assign n5722 = n62494 & n62667;
  assign n5723 = n62493 & ~n5722;
  assign n5724 = n62493 & ~n5715;
  assign n5725 = ~n5722 & n5724;
  assign n5726 = ~n5715 & n5723;
  assign n5727 = n62494 & ~n5714;
  assign n5728 = ~n62494 & n62667;
  assign n5729 = ~n62493 & ~n5728;
  assign n5730 = ~n62493 & ~n5727;
  assign n5731 = ~n5728 & n5730;
  assign n5732 = ~n5727 & n5729;
  assign n5733 = pi1197 & ~n62669;
  assign n5734 = pi1197 & ~n62668;
  assign n5735 = ~n62669 & n5734;
  assign n5736 = ~n62668 & n5733;
  assign n5737 = ~pi1197 & ~n5541;
  assign n5738 = ~n62490 & ~n5737;
  assign n5739 = ~n62670 & n5738;
  assign n5740 = n62490 & n5705;
  assign n5741 = ~pi1199 & ~n5740;
  assign n5742 = ~n5739 & n5741;
  assign n5743 = ~pi1198 & n5742;
  assign n5744 = pi1198 & ~n5705;
  assign n5745 = ~n5275 & n5705;
  assign n5746 = n5275 & n5541;
  assign n5747 = ~n5745 & ~n5746;
  assign n5748 = n4818 & n5747;
  assign n5749 = ~n5744 & ~n5748;
  assign n5750 = pi1199 & ~n5746;
  assign n5751 = pi1199 & n5747;
  assign n5752 = ~n5745 & n5750;
  assign n5753 = ~n5742 & ~n62671;
  assign n5754 = ~pi1198 & ~n5753;
  assign n5755 = ~n5744 & ~n5754;
  assign n5756 = ~n5743 & n5749;
  assign n5757 = pi374 & ~n62672;
  assign n5758 = ~pi369 & n62518;
  assign n5759 = pi369 & ~n62518;
  assign n5760 = ~n5758 & ~n5759;
  assign n5761 = ~pi374 & ~n5753;
  assign n5762 = ~n5760 & ~n5761;
  assign n5763 = ~n5757 & n5762;
  assign n5764 = ~pi374 & ~n62672;
  assign n5765 = pi374 & ~n5753;
  assign n5766 = n5760 & ~n5765;
  assign n5767 = ~n5764 & n5766;
  assign n5768 = ~pi591 & ~n5767;
  assign n5769 = ~pi591 & ~n5763;
  assign n5770 = ~n5767 & n5769;
  assign n5771 = ~n5757 & ~n5761;
  assign n5772 = ~pi369 & ~n5771;
  assign n5773 = ~n5764 & ~n5765;
  assign n5774 = pi369 & ~n5773;
  assign n5775 = n62518 & ~n5774;
  assign n5776 = n62518 & ~n5772;
  assign n5777 = ~n5774 & n5776;
  assign n5778 = ~n5772 & n5775;
  assign n5779 = pi369 & ~n5771;
  assign n5780 = ~pi369 & ~n5773;
  assign n5781 = ~n62518 & ~n5780;
  assign n5782 = ~n62518 & ~n5779;
  assign n5783 = ~n5780 & n5782;
  assign n5784 = ~n5779 & n5781;
  assign n5785 = ~pi591 & ~n62675;
  assign n5786 = ~n62674 & n5785;
  assign n5787 = ~pi591 & ~n62674;
  assign n5788 = ~n62675 & n5787;
  assign n5789 = ~n5763 & n5768;
  assign n5790 = n2580 & ~n5540;
  assign n5791 = ~pi122 & n2852;
  assign n5792 = ~n5538 & ~n5791;
  assign n5793 = ~n3032 & ~n5558;
  assign n5794 = n2852 & ~n62535;
  assign n5795 = ~pi122 & ~n5538;
  assign n5796 = ~n5794 & n5795;
  assign n5797 = ~n5793 & ~n5796;
  assign n5798 = ~n5792 & n5797;
  assign n5799 = pi567 & n5798;
  assign n5800 = ~n5540 & ~n5799;
  assign n5801 = ~n62530 & ~n5538;
  assign n5802 = ~n2852 & ~n5538;
  assign n5803 = ~n5801 & ~n5802;
  assign n5804 = n2852 & n62529;
  assign n5805 = ~n5538 & ~n5804;
  assign n5806 = pi412 & ~n5805;
  assign n5807 = n62526 & n4263;
  assign n5808 = ~n62526 & ~n4263;
  assign n5809 = n2852 & ~n5808;
  assign n5810 = ~n5807 & n5809;
  assign n5811 = n2852 & ~n62529;
  assign n5812 = ~n5538 & ~n62676;
  assign n5813 = ~pi412 & ~n5812;
  assign n5814 = ~n4220 & ~n5813;
  assign n5815 = ~n4220 & ~n5806;
  assign n5816 = ~n5813 & n5815;
  assign n5817 = ~n5806 & n5814;
  assign n5818 = ~pi412 & ~n5805;
  assign n5819 = pi412 & ~n5812;
  assign n5820 = n4220 & ~n5819;
  assign n5821 = n4220 & ~n5818;
  assign n5822 = ~n5819 & n5821;
  assign n5823 = ~n5818 & n5820;
  assign n5824 = ~pi122 & ~n62678;
  assign n5825 = ~n62677 & n5824;
  assign n5826 = ~pi122 & ~n62677;
  assign n5827 = ~n62678 & n5826;
  assign n5828 = ~pi122 & n5803;
  assign n5829 = ~n5538 & ~n62679;
  assign n5830 = n3032 & ~n5829;
  assign n5831 = ~n5558 & ~n5830;
  assign n5832 = pi567 & ~n5831;
  assign n5833 = n5800 & ~n5832;
  assign n5834 = ~n5790 & ~n5833;
  assign n5835 = n62373 & ~n5797;
  assign n5836 = ~n5830 & n5835;
  assign n5837 = ~n62535 & n5574;
  assign n5838 = n62535 & n5538;
  assign n5839 = ~n5837 & ~n5838;
  assign n5840 = n62655 & n5839;
  assign n5841 = n62530 & ~n5574;
  assign n5842 = ~n62530 & n5538;
  assign n5843 = n62530 & n5574;
  assign n5844 = ~n5842 & ~n5843;
  assign n5845 = ~pi411 & n5538;
  assign n5846 = ~n62531 & ~n5845;
  assign n5847 = pi411 & n5574;
  assign n5848 = n5846 & ~n5847;
  assign n5849 = n62531 & ~n5538;
  assign n5850 = ~n4287 & ~n5849;
  assign n5851 = ~pi411 & n5574;
  assign n5852 = ~n5850 & ~n5851;
  assign n5853 = ~n5848 & ~n5852;
  assign n5854 = ~n5801 & ~n5841;
  assign n5855 = pi411 & ~n62530;
  assign n5856 = n62531 & ~n5851;
  assign n5857 = ~n5848 & ~n5856;
  assign n5858 = ~n62680 & ~n5855;
  assign n5859 = n5840 & ~n62681;
  assign n5860 = n62530 & ~n5557;
  assign n5861 = pi411 & n5557;
  assign n5862 = n5846 & ~n5861;
  assign n5863 = ~pi411 & n5557;
  assign n5864 = ~n5850 & ~n5863;
  assign n5865 = ~n5862 & ~n5864;
  assign n5866 = ~n5801 & ~n5860;
  assign n5867 = ~n62535 & n5557;
  assign n5868 = n62653 & ~n5867;
  assign n5869 = n62407 & ~n62682;
  assign n5870 = ~n5867 & n5869;
  assign n5871 = ~n62682 & n5868;
  assign n5872 = ~n5859 & ~n62683;
  assign n5873 = ~pi122 & n5794;
  assign n5874 = ~n62679 & ~n5873;
  assign n5875 = ~n5872 & n5874;
  assign n5876 = ~n5836 & ~n5875;
  assign n5877 = ~pi75 & ~n5876;
  assign n5878 = ~n62374 & ~n5798;
  assign n5879 = ~n5830 & n5878;
  assign n5880 = n5592 & ~n5879;
  assign n5881 = ~n5877 & n5880;
  assign n5882 = ~n5834 & ~n5881;
  assign n5883 = n4494 & ~n5882;
  assign n5884 = ~n5790 & ~n5800;
  assign n5885 = ~n5838 & ~n5867;
  assign n5886 = n62653 & n5885;
  assign n5887 = ~n5840 & ~n5886;
  assign n5888 = pi122 & ~n5887;
  assign n5889 = ~n5835 & ~n5888;
  assign n5890 = ~pi75 & ~n5889;
  assign n5891 = n5592 & ~n5878;
  assign n5892 = ~n5890 & n5891;
  assign n5893 = ~n5884 & ~n5892;
  assign n5894 = n4537 & ~n5893;
  assign n5895 = pi1199 & ~n5894;
  assign n5896 = ~n5883 & n5895;
  assign n5897 = ~pi1199 & ~n5603;
  assign n5898 = ~n5540 & ~n5832;
  assign n5899 = ~n5790 & ~n5898;
  assign n5900 = n62655 & n62680;
  assign n5901 = ~n5869 & ~n5900;
  assign n5902 = ~n62679 & ~n5901;
  assign n5903 = ~pi122 & ~n62679;
  assign n5904 = ~pi122 & ~n5803;
  assign n5905 = ~n5793 & ~n62684;
  assign n5906 = n3032 & ~n62684;
  assign n5907 = n5559 & ~n5906;
  assign n5908 = n62373 & ~n5905;
  assign n5909 = ~n5902 & ~n62685;
  assign n5910 = ~pi75 & ~n5909;
  assign n5911 = ~n62374 & n5831;
  assign n5912 = n5592 & ~n5911;
  assign n5913 = pi122 & ~n62680;
  assign n5914 = ~n62679 & ~n5913;
  assign n5915 = n3032 & ~n5914;
  assign n5916 = n62655 & ~n5915;
  assign n5917 = pi122 & n62682;
  assign n5918 = ~n62679 & ~n5917;
  assign n5919 = n3032 & ~n5918;
  assign n5920 = n62653 & ~n5919;
  assign n5921 = ~n62373 & n5831;
  assign n5922 = ~n5920 & ~n5921;
  assign n5923 = ~n5916 & n5922;
  assign n5924 = ~pi75 & ~n5923;
  assign n5925 = pi75 & n5831;
  assign n5926 = n5592 & ~n5925;
  assign n5927 = ~n5924 & n5926;
  assign n5928 = ~n5910 & n5912;
  assign n5929 = ~n5899 & ~n62686;
  assign n5930 = n4494 & ~n5929;
  assign n5931 = n5897 & ~n5930;
  assign n5932 = n5205 & ~n5931;
  assign n5933 = ~n5896 & n5932;
  assign n5934 = ~n5205 & n5598;
  assign n5935 = ~n5545 & ~n5934;
  assign n5936 = ~n5933 & n5935;
  assign n5937 = ~pi1197 & ~n4621;
  assign n5938 = n5599 & ~n5937;
  assign n5939 = ~n5896 & ~n5931;
  assign n5940 = ~n5603 & ~n5930;
  assign n5941 = ~pi1199 & ~n5940;
  assign n5942 = ~n5883 & ~n5894;
  assign n5943 = pi1199 & ~n5942;
  assign n5944 = ~n5545 & ~n5943;
  assign n5945 = ~n5941 & n5944;
  assign n5946 = ~n5545 & ~n5939;
  assign n5947 = n5937 & n62687;
  assign n5948 = ~n5938 & ~n5947;
  assign n5949 = pi333 & ~n5948;
  assign n5950 = n4621 & ~n5599;
  assign n5951 = ~n4621 & ~n62687;
  assign n5952 = ~n5950 & ~n5951;
  assign n5953 = ~pi333 & n5952;
  assign n5954 = ~pi333 & ~n5952;
  assign n5955 = pi333 & n5948;
  assign n5956 = ~n5954 & ~n5955;
  assign n5957 = ~n5949 & ~n5953;
  assign n5958 = pi391 & n62688;
  assign n5959 = pi333 & ~n5952;
  assign n5960 = ~pi333 & n5948;
  assign n5961 = ~n5959 & ~n5960;
  assign n5962 = ~pi391 & n5961;
  assign n5963 = ~pi391 & ~n5961;
  assign n5964 = pi391 & ~n62688;
  assign n5965 = ~n5963 & ~n5964;
  assign n5966 = ~n5958 & ~n5962;
  assign n5967 = pi392 & ~n62689;
  assign n5968 = ~pi391 & ~n62688;
  assign n5969 = pi391 & ~n5961;
  assign n5970 = ~n5968 & ~n5969;
  assign n5971 = ~pi392 & ~n5970;
  assign n5972 = ~n62523 & ~n5971;
  assign n5973 = ~n5967 & n5972;
  assign n5974 = ~pi392 & ~n62689;
  assign n5975 = pi392 & ~n5970;
  assign n5976 = n62523 & ~n5975;
  assign n5977 = ~n5974 & n5976;
  assign n5978 = pi591 & ~n5977;
  assign n5979 = ~n5973 & n5978;
  assign n5980 = ~pi392 & n62689;
  assign n5981 = pi392 & n5970;
  assign n5982 = ~n5974 & ~n5975;
  assign n5983 = ~n5980 & ~n5981;
  assign n5984 = pi393 & n62691;
  assign n5985 = pi392 & n62689;
  assign n5986 = ~pi392 & n5970;
  assign n5987 = ~n5985 & ~n5986;
  assign n5988 = ~pi393 & ~n5987;
  assign n5989 = ~n5984 & ~n5988;
  assign n5990 = pi393 & ~n62691;
  assign n5991 = ~pi393 & n5987;
  assign n5992 = ~n62522 & ~n5991;
  assign n5993 = ~n5990 & n5992;
  assign n5994 = ~n62522 & ~n5989;
  assign n5995 = pi393 & ~n5987;
  assign n5996 = ~pi393 & n62691;
  assign n5997 = ~n5995 & ~n5996;
  assign n5998 = ~pi393 & ~n62691;
  assign n5999 = pi393 & n5987;
  assign n6000 = n62522 & ~n5999;
  assign n6001 = ~n5998 & n6000;
  assign n6002 = n62522 & ~n5997;
  assign n6003 = pi591 & ~n62693;
  assign n6004 = ~n62692 & n6003;
  assign n6005 = pi591 & ~n62692;
  assign n6006 = ~n62693 & n6005;
  assign n6007 = pi591 & ~n5936;
  assign n6008 = ~pi590 & ~n62690;
  assign n6009 = ~n62673 & n6008;
  assign n6010 = ~pi588 & ~n6009;
  assign n6011 = ~n5702 & n6010;
  assign n6012 = ~n3312 & n5541;
  assign n6013 = pi588 & ~n6012;
  assign n6014 = ~n2578 & n5599;
  assign n6015 = n2578 & ~n5603;
  assign n6016 = pi443 & ~n5541;
  assign n6017 = n62426 & ~n6016;
  assign n6018 = ~pi443 & ~n5599;
  assign n6019 = n6017 & ~n6018;
  assign n6020 = ~pi443 & ~n5541;
  assign n6021 = ~n62426 & ~n6020;
  assign n6022 = pi443 & ~n5599;
  assign n6023 = n6021 & ~n6022;
  assign n6024 = pi1196 & ~n6023;
  assign n6025 = ~n6020 & ~n6022;
  assign n6026 = n3188 & n6025;
  assign n6027 = ~n6016 & ~n6018;
  assign n6028 = ~n3188 & n6027;
  assign n6029 = ~n6026 & ~n6028;
  assign n6030 = ~pi435 & ~n6029;
  assign n6031 = n3188 & n6027;
  assign n6032 = ~n3188 & n6025;
  assign n6033 = ~pi444 & n6027;
  assign n6034 = pi444 & n6025;
  assign n6035 = ~pi436 & ~n6034;
  assign n6036 = ~pi436 & ~n6033;
  assign n6037 = ~n6034 & n6036;
  assign n6038 = ~n6033 & n6035;
  assign n6039 = ~pi444 & n6025;
  assign n6040 = pi444 & n6027;
  assign n6041 = pi436 & ~n6040;
  assign n6042 = pi436 & ~n6039;
  assign n6043 = ~n6040 & n6042;
  assign n6044 = ~n6039 & n6041;
  assign n6045 = ~n62694 & ~n62695;
  assign n6046 = ~n6031 & ~n6032;
  assign n6047 = pi435 & n62696;
  assign n6048 = ~n6030 & ~n6047;
  assign n6049 = ~pi429 & n6048;
  assign n6050 = pi435 & ~n6029;
  assign n6051 = ~pi435 & n62696;
  assign n6052 = ~n6050 & ~n6051;
  assign n6053 = pi429 & n6052;
  assign n6054 = ~n3172 & ~n6053;
  assign n6055 = ~n3172 & ~n6049;
  assign n6056 = ~n6053 & n6055;
  assign n6057 = ~n6049 & n6054;
  assign n6058 = ~pi429 & n6052;
  assign n6059 = pi429 & n6048;
  assign n6060 = n3172 & ~n6059;
  assign n6061 = n3172 & ~n6058;
  assign n6062 = ~n6059 & n6061;
  assign n6063 = ~n6058 & n6060;
  assign n6064 = pi1196 & ~n62698;
  assign n6065 = ~n62697 & n6064;
  assign n6066 = pi1196 & ~n62697;
  assign n6067 = ~n62698 & n6066;
  assign n6068 = ~n6019 & n6024;
  assign n6069 = n6015 & ~n62699;
  assign n6070 = ~n6014 & ~n6069;
  assign n6071 = pi428 & ~n6070;
  assign n6072 = ~pi428 & n5599;
  assign n6073 = ~n6071 & ~n6072;
  assign n6074 = ~pi427 & ~n6073;
  assign n6075 = ~pi428 & ~n6070;
  assign n6076 = pi428 & n5599;
  assign n6077 = pi428 & ~n5599;
  assign n6078 = ~pi428 & n6070;
  assign n6079 = ~n6077 & ~n6078;
  assign n6080 = ~n6075 & ~n6076;
  assign n6081 = pi427 & n62700;
  assign n6082 = ~n6074 & ~n6081;
  assign n6083 = pi430 & n6082;
  assign n6084 = ~n62450 & ~n62643;
  assign n6085 = n62450 & n62643;
  assign n6086 = ~n6084 & ~n6085;
  assign n6087 = ~pi427 & n62700;
  assign n6088 = pi427 & ~n6073;
  assign n6089 = ~n6087 & ~n6088;
  assign n6090 = ~pi430 & n6089;
  assign n6091 = ~n6086 & ~n6090;
  assign n6092 = ~n6083 & ~n6086;
  assign n6093 = ~n6090 & n6092;
  assign n6094 = ~n6083 & n6091;
  assign n6095 = ~pi430 & n6082;
  assign n6096 = pi430 & n6089;
  assign n6097 = n6086 & ~n6096;
  assign n6098 = ~n6095 & n6097;
  assign n6099 = pi1199 & ~n6098;
  assign n6100 = pi430 & ~n6082;
  assign n6101 = ~pi430 & ~n6089;
  assign n6102 = ~n6100 & ~n6101;
  assign n6103 = pi426 & ~n6102;
  assign n6104 = pi430 & ~n6089;
  assign n6105 = ~pi430 & ~n6082;
  assign n6106 = ~n6104 & ~n6105;
  assign n6107 = ~pi426 & ~n6106;
  assign n6108 = ~n6103 & ~n6107;
  assign n6109 = pi445 & ~n6108;
  assign n6110 = pi426 & ~n6106;
  assign n6111 = ~pi426 & ~n6102;
  assign n6112 = ~n6110 & ~n6111;
  assign n6113 = ~pi445 & ~n6112;
  assign n6114 = ~n6109 & ~n6113;
  assign n6115 = ~pi448 & n6114;
  assign n6116 = pi445 & ~n6112;
  assign n6117 = ~pi445 & ~n6108;
  assign n6118 = ~n6116 & ~n6117;
  assign n6119 = pi448 & n6118;
  assign n6120 = n3269 & ~n6119;
  assign n6121 = n3269 & ~n6115;
  assign n6122 = ~n6119 & n6121;
  assign n6123 = ~n6115 & n6120;
  assign n6124 = pi448 & n6114;
  assign n6125 = ~pi448 & n6118;
  assign n6126 = ~n3269 & ~n6125;
  assign n6127 = ~n3269 & ~n6124;
  assign n6128 = ~n6125 & n6127;
  assign n6129 = ~n6124 & n6126;
  assign n6130 = pi1199 & ~n62703;
  assign n6131 = ~n62702 & n6130;
  assign n6132 = pi1199 & ~n62702;
  assign n6133 = ~n62703 & n6132;
  assign n6134 = ~n62701 & n6099;
  assign n6135 = ~pi1199 & n6070;
  assign n6136 = n3312 & ~n6135;
  assign n6137 = ~n62704 & n6136;
  assign n6138 = n6013 & ~n6137;
  assign n6139 = ~n3318 & ~n6138;
  assign n6140 = ~n3318 & ~n6011;
  assign n6141 = ~n6138 & n6140;
  assign n6142 = ~n6011 & n6139;
  assign n6143 = ~n2580 & n5541;
  assign n6144 = n62407 & ~n5793;
  assign n6145 = n5557 & n6144;
  assign n6146 = n2806 & ~n5793;
  assign n6147 = n5574 & n6146;
  assign n6148 = ~n6145 & ~n6147;
  assign n6149 = ~pi75 & ~n6148;
  assign n6150 = ~n62374 & n5539;
  assign n6151 = pi75 & n5539;
  assign n6152 = ~n62373 & n5539;
  assign n6153 = ~n6145 & ~n6152;
  assign n6154 = ~n6147 & n6153;
  assign n6155 = ~pi75 & ~n6154;
  assign n6156 = ~n6151 & ~n6155;
  assign n6157 = ~n6149 & ~n6150;
  assign n6158 = pi567 & ~n62706;
  assign n6159 = n5790 & ~n6158;
  assign n6160 = ~n6143 & ~n6159;
  assign n6161 = ~pi592 & n6160;
  assign n6162 = ~n5545 & ~n6161;
  assign n6163 = ~n5345 & n6162;
  assign n6164 = ~n5544 & ~n6163;
  assign n6165 = pi1198 & ~n6164;
  assign n6166 = ~n62464 & n6162;
  assign n6167 = ~n5605 & ~n6166;
  assign n6168 = ~pi355 & ~n6167;
  assign n6169 = ~pi455 & ~n6162;
  assign n6170 = ~n5609 & ~n6169;
  assign n6171 = ~pi452 & ~n6170;
  assign n6172 = pi455 & ~n6162;
  assign n6173 = ~n5613 & ~n6172;
  assign n6174 = pi452 & ~n6173;
  assign n6175 = ~n6171 & ~n6174;
  assign n6176 = pi355 & n6175;
  assign n6177 = ~n6168 & ~n6176;
  assign n6178 = ~pi458 & n6177;
  assign n6179 = pi355 & ~n6167;
  assign n6180 = ~pi355 & n6175;
  assign n6181 = ~n6179 & ~n6180;
  assign n6182 = pi458 & n6181;
  assign n6183 = n62462 & ~n6182;
  assign n6184 = n62462 & ~n6178;
  assign n6185 = ~n6182 & n6184;
  assign n6186 = ~n6178 & n6183;
  assign n6187 = ~pi458 & n6181;
  assign n6188 = pi458 & n6177;
  assign n6189 = ~n62462 & ~n6188;
  assign n6190 = ~n62462 & ~n6187;
  assign n6191 = ~n6188 & n6190;
  assign n6192 = ~n6187 & n6189;
  assign n6193 = pi1196 & ~n62708;
  assign n6194 = pi1196 & ~n62707;
  assign n6195 = ~n62708 & n6194;
  assign n6196 = ~n62707 & n6193;
  assign n6197 = n5604 & ~n62709;
  assign n6198 = ~n6165 & ~n6197;
  assign n6199 = ~n62460 & ~n6198;
  assign n6200 = n62460 & n6162;
  assign n6201 = ~n6199 & ~n6200;
  assign n6202 = ~n3767 & n6201;
  assign n6203 = pi1199 & ~n6162;
  assign n6204 = pi351 & n6203;
  assign n6205 = ~n62635 & ~n6204;
  assign n6206 = ~n6202 & n6205;
  assign n6207 = ~n3478 & n6201;
  assign n6208 = ~pi351 & n6203;
  assign n6209 = n62635 & ~n6208;
  assign n6210 = ~n6207 & n6209;
  assign n6211 = ~pi591 & ~n6210;
  assign n6212 = ~pi591 & ~n6206;
  assign n6213 = ~n6210 & n6212;
  assign n6214 = ~n6207 & ~n6208;
  assign n6215 = ~pi461 & ~n6214;
  assign n6216 = ~n6202 & ~n6204;
  assign n6217 = pi461 & ~n6216;
  assign n6218 = ~n6215 & ~n6217;
  assign n6219 = ~pi357 & ~n6218;
  assign n6220 = ~pi461 & ~n6216;
  assign n6221 = pi461 & ~n6214;
  assign n6222 = ~n6220 & ~n6221;
  assign n6223 = pi357 & ~n6222;
  assign n6224 = ~n6219 & ~n6223;
  assign n6225 = pi357 & n6222;
  assign n6226 = ~pi357 & n6218;
  assign n6227 = ~pi356 & ~n6226;
  assign n6228 = ~n6225 & n6227;
  assign n6229 = ~pi356 & ~n6224;
  assign n6230 = ~pi357 & ~n6222;
  assign n6231 = pi357 & ~n6218;
  assign n6232 = ~n6230 & ~n6231;
  assign n6233 = pi357 & n6218;
  assign n6234 = ~pi357 & n6222;
  assign n6235 = pi356 & ~n6234;
  assign n6236 = ~n6233 & n6235;
  assign n6237 = pi356 & ~n6232;
  assign n6238 = ~n62711 & ~n62712;
  assign n6239 = ~pi354 & ~n6238;
  assign n6240 = ~n62599 & n6222;
  assign n6241 = n62599 & n6218;
  assign n6242 = ~pi356 & ~n6232;
  assign n6243 = pi356 & ~n6224;
  assign n6244 = ~n6242 & ~n6243;
  assign n6245 = ~n6240 & ~n6241;
  assign n6246 = pi354 & ~n62713;
  assign n6247 = ~n62480 & ~n6246;
  assign n6248 = ~n62480 & ~n6239;
  assign n6249 = ~n6246 & n6248;
  assign n6250 = ~n6239 & n6247;
  assign n6251 = pi354 & ~n6238;
  assign n6252 = ~pi354 & ~n62713;
  assign n6253 = n62480 & ~n6252;
  assign n6254 = n62480 & ~n6251;
  assign n6255 = ~n6252 & n6254;
  assign n6256 = ~n6251 & n6253;
  assign n6257 = ~pi591 & ~n62715;
  assign n6258 = ~n62714 & n6257;
  assign n6259 = ~pi591 & ~n62714;
  assign n6260 = ~n62715 & n6259;
  assign n6261 = ~n6206 & n6211;
  assign n6262 = n5543 & ~n62710;
  assign n6263 = pi592 & n6160;
  assign n6264 = ~n5703 & ~n6263;
  assign n6265 = pi1198 & ~n6264;
  assign n6266 = n62518 & ~n6265;
  assign n6267 = n62519 & ~n6266;
  assign n6268 = ~n62519 & n6265;
  assign n6269 = ~n62518 & ~n6265;
  assign n6270 = ~n62519 & ~n6269;
  assign n6271 = pi1198 & ~n6270;
  assign n6272 = n5282 & ~n6268;
  assign n6273 = n4031 & ~n5541;
  assign n6274 = ~n4031 & ~n6264;
  assign n6275 = ~n5275 & n6264;
  assign n6276 = n5750 & ~n6275;
  assign n6277 = n62497 & n6264;
  assign n6278 = ~n62497 & n5541;
  assign n6279 = pi1197 & ~n6278;
  assign n6280 = ~n6277 & n6279;
  assign n6281 = n5738 & ~n6280;
  assign n6282 = n62490 & n6264;
  assign n6283 = ~pi1199 & ~n6282;
  assign n6284 = ~n6281 & n6283;
  assign n6285 = ~n6276 & ~n6284;
  assign n6286 = ~n6273 & ~n6274;
  assign n6287 = n62518 & n62717;
  assign n6288 = ~n62716 & ~n6287;
  assign n6289 = ~n6267 & ~n6288;
  assign n6290 = ~n62518 & ~n6268;
  assign n6291 = ~pi1198 & ~n62717;
  assign n6292 = ~n6265 & ~n6291;
  assign n6293 = ~pi374 & ~n6292;
  assign n6294 = pi374 & ~n62717;
  assign n6295 = ~n6293 & ~n6294;
  assign n6296 = ~pi369 & ~n6295;
  assign n6297 = ~pi374 & ~n62717;
  assign n6298 = pi374 & ~n6292;
  assign n6299 = ~n6297 & ~n6298;
  assign n6300 = pi369 & ~n6299;
  assign n6301 = ~n62518 & ~n6300;
  assign n6302 = ~n6296 & n6301;
  assign n6303 = ~n62518 & ~n6296;
  assign n6304 = ~n6300 & n6303;
  assign n6305 = n62717 & n6290;
  assign n6306 = ~n62518 & n62717;
  assign n6307 = n6267 & ~n6306;
  assign n6308 = ~n62518 & n6270;
  assign n6309 = n62717 & ~n6308;
  assign n6310 = ~n62716 & ~n6309;
  assign n6311 = ~n6307 & ~n6310;
  assign n6312 = ~n6289 & ~n62718;
  assign n6313 = ~pi591 & n62719;
  assign n6314 = ~n5545 & ~n5603;
  assign n6315 = ~pi1199 & n6314;
  assign n6316 = ~n5545 & n5897;
  assign n6317 = n4494 & ~n6143;
  assign n6318 = ~n62680 & n6146;
  assign n6319 = n62682 & n6144;
  assign n6320 = ~n6318 & ~n6319;
  assign n6321 = ~pi75 & ~n6320;
  assign n6322 = ~n6152 & ~n6319;
  assign n6323 = ~n6318 & n6322;
  assign n6324 = ~pi75 & ~n6323;
  assign n6325 = ~n6151 & ~n6324;
  assign n6326 = ~n6150 & ~n6321;
  assign n6327 = pi567 & ~n62721;
  assign n6328 = n5790 & ~n6327;
  assign n6329 = n6317 & ~n6328;
  assign n6330 = n62720 & ~n6329;
  assign n6331 = ~n5839 & n6147;
  assign n6332 = ~n62535 & n6145;
  assign n6333 = ~n6152 & ~n6332;
  assign n6334 = ~n6331 & n6333;
  assign n6335 = ~n6331 & ~n6332;
  assign n6336 = n6323 & n6335;
  assign n6337 = n6320 & n6334;
  assign n6338 = n6317 & ~n62722;
  assign n6339 = ~n5885 & n6145;
  assign n6340 = ~n6152 & ~n6339;
  assign n6341 = ~n6331 & n6340;
  assign n6342 = n4537 & ~n6143;
  assign n6343 = ~n6341 & n6342;
  assign n6344 = ~n6338 & ~n6343;
  assign n6345 = ~pi75 & pi567;
  assign n6346 = ~n6344 & n6345;
  assign n6347 = n4998 & n5790;
  assign n6348 = ~n5541 & ~n6347;
  assign n6349 = pi1199 & ~n6348;
  assign n6350 = ~n6346 & n6349;
  assign n6351 = n5205 & ~n6350;
  assign n6352 = ~n6330 & n6351;
  assign n6353 = ~n5205 & ~n6162;
  assign n6354 = pi591 & ~n6353;
  assign n6355 = ~n6352 & n6354;
  assign n6356 = ~n6313 & ~n6355;
  assign n6357 = ~n5937 & ~n6162;
  assign n6358 = ~n4621 & ~n6350;
  assign n6359 = ~n6330 & n6358;
  assign n6360 = ~pi1197 & n6359;
  assign n6361 = ~n6357 & ~n6360;
  assign n6362 = ~pi333 & ~n6361;
  assign n6363 = n4621 & ~n6162;
  assign n6364 = ~n6359 & ~n6363;
  assign n6365 = pi333 & ~n6364;
  assign n6366 = ~n6362 & ~n6365;
  assign n6367 = ~pi391 & ~n6366;
  assign n6368 = pi333 & ~n6361;
  assign n6369 = ~pi333 & ~n6364;
  assign n6370 = ~n6368 & ~n6369;
  assign n6371 = pi391 & ~n6370;
  assign n6372 = ~n6367 & ~n6371;
  assign n6373 = pi392 & ~n6372;
  assign n6374 = ~pi391 & ~n6370;
  assign n6375 = pi391 & ~n6366;
  assign n6376 = ~n6374 & ~n6375;
  assign n6377 = ~pi392 & ~n6376;
  assign n6378 = ~n62523 & ~n6377;
  assign n6379 = ~n6373 & n6378;
  assign n6380 = ~pi392 & ~n6372;
  assign n6381 = pi392 & ~n6376;
  assign n6382 = n62523 & ~n6381;
  assign n6383 = ~n6380 & n6382;
  assign n6384 = pi591 & ~n6383;
  assign n6385 = ~n6380 & ~n6381;
  assign n6386 = ~pi393 & ~n6385;
  assign n6387 = ~n6373 & ~n6377;
  assign n6388 = pi393 & ~n6387;
  assign n6389 = n62522 & ~n6388;
  assign n6390 = n62522 & ~n6386;
  assign n6391 = ~n6388 & n6390;
  assign n6392 = ~n6386 & n6389;
  assign n6393 = ~pi393 & ~n6387;
  assign n6394 = pi393 & ~n6385;
  assign n6395 = ~n62522 & ~n6394;
  assign n6396 = ~n62522 & ~n6393;
  assign n6397 = ~n6394 & n6396;
  assign n6398 = ~n6393 & n6395;
  assign n6399 = pi591 & ~n62724;
  assign n6400 = ~n62723 & n6399;
  assign n6401 = pi591 & ~n62723;
  assign n6402 = ~n62724 & n6401;
  assign n6403 = ~n6379 & n6384;
  assign n6404 = ~pi369 & ~n6299;
  assign n6405 = pi369 & ~n6295;
  assign n6406 = n62518 & ~n6405;
  assign n6407 = n62518 & ~n6404;
  assign n6408 = ~n6405 & n6407;
  assign n6409 = ~n6404 & n6406;
  assign n6410 = ~pi591 & ~n62718;
  assign n6411 = ~n62726 & n6410;
  assign n6412 = ~pi591 & ~n62726;
  assign n6413 = ~n62718 & n6412;
  assign n6414 = ~pi591 & ~n62719;
  assign n6415 = ~pi590 & ~n62727;
  assign n6416 = ~n62725 & n6415;
  assign n6417 = ~pi590 & ~n6356;
  assign n6418 = ~pi588 & ~n62728;
  assign n6419 = ~n6262 & n6418;
  assign n6420 = ~n2578 & n6162;
  assign n6421 = ~pi443 & ~n6162;
  assign n6422 = n6017 & ~n6421;
  assign n6423 = pi443 & ~n6162;
  assign n6424 = n6021 & ~n6423;
  assign n6425 = pi1196 & ~n6424;
  assign n6426 = ~n6020 & ~n6423;
  assign n6427 = n3188 & n6426;
  assign n6428 = ~n6016 & ~n6421;
  assign n6429 = ~n3188 & n6428;
  assign n6430 = ~n6427 & ~n6429;
  assign n6431 = ~pi435 & ~n6430;
  assign n6432 = n3188 & n6428;
  assign n6433 = ~n3188 & n6426;
  assign n6434 = ~pi444 & n6428;
  assign n6435 = pi444 & n6426;
  assign n6436 = ~pi436 & ~n6435;
  assign n6437 = ~pi436 & ~n6434;
  assign n6438 = ~n6435 & n6437;
  assign n6439 = ~n6434 & n6436;
  assign n6440 = ~pi444 & n6426;
  assign n6441 = pi444 & n6428;
  assign n6442 = pi436 & ~n6441;
  assign n6443 = pi436 & ~n6440;
  assign n6444 = ~n6441 & n6443;
  assign n6445 = ~n6440 & n6442;
  assign n6446 = ~n62729 & ~n62730;
  assign n6447 = ~n6432 & ~n6433;
  assign n6448 = pi435 & n62731;
  assign n6449 = ~n6431 & ~n6448;
  assign n6450 = ~pi429 & n6449;
  assign n6451 = pi435 & ~n6430;
  assign n6452 = ~pi435 & n62731;
  assign n6453 = ~n6451 & ~n6452;
  assign n6454 = pi429 & n6453;
  assign n6455 = ~n3172 & ~n6454;
  assign n6456 = ~n3172 & ~n6450;
  assign n6457 = ~n6454 & n6456;
  assign n6458 = ~n6450 & n6455;
  assign n6459 = ~pi429 & n6453;
  assign n6460 = pi429 & n6449;
  assign n6461 = n3172 & ~n6460;
  assign n6462 = n3172 & ~n6459;
  assign n6463 = ~n6460 & n6462;
  assign n6464 = ~n6459 & n6461;
  assign n6465 = pi1196 & ~n62733;
  assign n6466 = ~n62732 & n6465;
  assign n6467 = pi1196 & ~n62732;
  assign n6468 = ~n62733 & n6467;
  assign n6469 = ~n6422 & n6425;
  assign n6470 = n6015 & ~n62734;
  assign n6471 = ~n6420 & ~n6470;
  assign n6472 = pi428 & ~n6471;
  assign n6473 = ~pi428 & n6162;
  assign n6474 = ~n6472 & ~n6473;
  assign n6475 = ~pi427 & ~n6474;
  assign n6476 = ~pi428 & ~n6471;
  assign n6477 = pi428 & n6162;
  assign n6478 = pi428 & ~n6162;
  assign n6479 = ~pi428 & n6471;
  assign n6480 = ~n6478 & ~n6479;
  assign n6481 = ~n6476 & ~n6477;
  assign n6482 = pi427 & n62735;
  assign n6483 = ~n6475 & ~n6482;
  assign n6484 = pi430 & n6483;
  assign n6485 = ~pi427 & n62735;
  assign n6486 = pi427 & ~n6474;
  assign n6487 = ~n6485 & ~n6486;
  assign n6488 = ~pi430 & n6487;
  assign n6489 = ~n6086 & ~n6488;
  assign n6490 = ~n6086 & ~n6484;
  assign n6491 = ~n6488 & n6490;
  assign n6492 = ~n6484 & n6489;
  assign n6493 = ~pi430 & n6483;
  assign n6494 = pi430 & n6487;
  assign n6495 = n6086 & ~n6494;
  assign n6496 = ~n6493 & n6495;
  assign n6497 = pi1199 & ~n6496;
  assign n6498 = pi430 & ~n6483;
  assign n6499 = ~pi430 & ~n6487;
  assign n6500 = ~n6498 & ~n6499;
  assign n6501 = pi426 & ~n6500;
  assign n6502 = pi430 & ~n6487;
  assign n6503 = ~pi430 & ~n6483;
  assign n6504 = ~n6502 & ~n6503;
  assign n6505 = ~pi426 & ~n6504;
  assign n6506 = ~n6501 & ~n6505;
  assign n6507 = pi445 & ~n6506;
  assign n6508 = pi426 & ~n6504;
  assign n6509 = ~pi426 & ~n6500;
  assign n6510 = ~n6508 & ~n6509;
  assign n6511 = ~pi445 & ~n6510;
  assign n6512 = ~n6507 & ~n6511;
  assign n6513 = pi448 & n6512;
  assign n6514 = pi445 & ~n6510;
  assign n6515 = ~pi445 & ~n6506;
  assign n6516 = ~n6514 & ~n6515;
  assign n6517 = ~pi448 & n6516;
  assign n6518 = ~n3269 & ~n6517;
  assign n6519 = ~n3269 & ~n6513;
  assign n6520 = ~n6517 & n6519;
  assign n6521 = ~n6513 & n6518;
  assign n6522 = pi448 & n6516;
  assign n6523 = ~pi448 & n6512;
  assign n6524 = n3269 & ~n6523;
  assign n6525 = n3269 & ~n6522;
  assign n6526 = ~n6523 & n6525;
  assign n6527 = ~n6522 & n6524;
  assign n6528 = pi1199 & ~n62738;
  assign n6529 = ~n62737 & n6528;
  assign n6530 = pi1199 & ~n62737;
  assign n6531 = ~n62738 & n6530;
  assign n6532 = ~n62736 & n6497;
  assign n6533 = ~pi1199 & n6471;
  assign n6534 = n3312 & ~n6533;
  assign n6535 = ~n62739 & n6534;
  assign n6536 = n6013 & ~n6535;
  assign n6537 = n3318 & ~n6536;
  assign n6538 = n3318 & ~n6419;
  assign n6539 = ~n6536 & n6538;
  assign n6540 = ~n6419 & n6537;
  assign n6541 = ~pi80 & n62455;
  assign n6542 = ~n62740 & n6541;
  assign n6543 = ~n62705 & n6541;
  assign n6544 = ~n62740 & n6543;
  assign n6545 = ~n62705 & n6542;
  assign n6546 = ~pi1196 & n5800;
  assign n6547 = ~pi592 & ~n6546;
  assign n6548 = ~n5833 & n6547;
  assign n6549 = pi1199 & ~n5545;
  assign n6550 = ~n6548 & n6549;
  assign n6551 = n4494 & ~n5898;
  assign n6552 = n62720 & ~n6551;
  assign n6553 = n5205 & ~n6552;
  assign n6554 = ~n5800 & ~n62720;
  assign n6555 = pi1196 & ~n5898;
  assign n6556 = ~n6554 & ~n6555;
  assign n6557 = ~pi592 & ~n6556;
  assign n6558 = ~pi1199 & n5603;
  assign n6559 = ~n5545 & ~n6558;
  assign n6560 = n6314 & ~n6551;
  assign n6561 = ~pi1199 & ~n6560;
  assign n6562 = n4494 & ~n5833;
  assign n6563 = n4537 & ~n5800;
  assign n6564 = ~n5545 & ~n6563;
  assign n6565 = ~n6562 & n6564;
  assign n6566 = pi1199 & ~n6565;
  assign n6567 = ~n6561 & ~n6566;
  assign n6568 = ~n6557 & n6559;
  assign n6569 = n5205 & ~n62742;
  assign n6570 = ~n6550 & n6553;
  assign n6571 = ~n5285 & n5541;
  assign n6572 = ~n5205 & ~n6571;
  assign n6573 = pi591 & ~n6572;
  assign n6574 = ~n62743 & n6573;
  assign n6575 = n5279 & ~n5283;
  assign n6576 = n3132 & ~n3686;
  assign n6577 = n3132 & ~n5279;
  assign n6578 = ~pi1198 & ~n6577;
  assign n6579 = ~n5232 & ~n62630;
  assign n6580 = ~n6578 & n6579;
  assign n6581 = ~n5232 & ~n6578;
  assign n6582 = ~n62630 & n6581;
  assign n6583 = ~n6575 & n6576;
  assign n6584 = ~pi591 & n5541;
  assign n6585 = ~n62744 & n6584;
  assign n6586 = ~n6574 & ~n6585;
  assign n6587 = ~n5937 & ~n6571;
  assign n6588 = n5937 & ~n62742;
  assign n6589 = ~n6587 & ~n6588;
  assign n6590 = pi333 & ~n6589;
  assign n6591 = n4621 & ~n6571;
  assign n6592 = ~n4621 & ~n62742;
  assign n6593 = ~n6591 & ~n6592;
  assign n6594 = ~pi333 & ~n6593;
  assign n6595 = ~n6590 & ~n6594;
  assign n6596 = pi391 & ~n6595;
  assign n6597 = ~pi333 & ~n6589;
  assign n6598 = pi333 & ~n6593;
  assign n6599 = ~n6597 & ~n6598;
  assign n6600 = ~pi391 & ~n6599;
  assign n6601 = ~n4206 & ~n6600;
  assign n6602 = ~n4206 & ~n6596;
  assign n6603 = ~n6600 & n6602;
  assign n6604 = ~n6596 & n6601;
  assign n6605 = pi391 & ~n6599;
  assign n6606 = ~pi391 & ~n6595;
  assign n6607 = n4206 & ~n6606;
  assign n6608 = n4206 & ~n6605;
  assign n6609 = ~n6606 & n6608;
  assign n6610 = ~n6605 & n6607;
  assign n6611 = pi591 & ~n62746;
  assign n6612 = pi591 & ~n62745;
  assign n6613 = ~n62746 & n6612;
  assign n6614 = ~n62745 & n6611;
  assign n6615 = n5541 & ~n62744;
  assign n6616 = ~pi591 & ~n6615;
  assign n6617 = ~pi590 & ~n6616;
  assign n6618 = ~n62747 & n6617;
  assign n6619 = ~pi590 & ~n6586;
  assign n6620 = n3767 & ~n62635;
  assign n6621 = n3478 & n62635;
  assign n6622 = ~n5213 & n5541;
  assign n6623 = ~n6621 & n6622;
  assign n6624 = ~n6620 & n6623;
  assign n6625 = n5351 & n6624;
  assign n6626 = ~pi591 & ~n6571;
  assign n6627 = n5351 & n6622;
  assign n6628 = ~n3478 & n6627;
  assign n6629 = ~n6571 & ~n6628;
  assign n6630 = pi461 & ~n6629;
  assign n6631 = ~n3767 & n6627;
  assign n6632 = ~n6571 & ~n6631;
  assign n6633 = ~pi461 & ~n6632;
  assign n6634 = ~n6630 & ~n6633;
  assign n6635 = ~n62599 & n6634;
  assign n6636 = pi461 & ~n6632;
  assign n6637 = ~pi461 & ~n6629;
  assign n6638 = ~n6636 & ~n6637;
  assign n6639 = n62599 & n6638;
  assign n6640 = pi357 & ~n6634;
  assign n6641 = ~pi357 & ~n6638;
  assign n6642 = ~n6640 & ~n6641;
  assign n6643 = pi356 & ~n6642;
  assign n6644 = pi357 & ~n6638;
  assign n6645 = ~pi357 & ~n6634;
  assign n6646 = ~n6644 & ~n6645;
  assign n6647 = ~pi356 & ~n6646;
  assign n6648 = ~n6643 & ~n6647;
  assign n6649 = ~n6635 & ~n6639;
  assign n6650 = pi354 & n62749;
  assign n6651 = n62599 & ~n6634;
  assign n6652 = ~n62599 & ~n6638;
  assign n6653 = pi357 & n6638;
  assign n6654 = ~pi357 & n6634;
  assign n6655 = pi356 & ~n6654;
  assign n6656 = ~n6653 & n6655;
  assign n6657 = pi356 & ~n6646;
  assign n6658 = pi357 & n6634;
  assign n6659 = ~pi357 & n6638;
  assign n6660 = ~pi356 & ~n6659;
  assign n6661 = ~n6658 & n6660;
  assign n6662 = ~pi356 & ~n6642;
  assign n6663 = ~n62750 & ~n62751;
  assign n6664 = ~n6651 & ~n6652;
  assign n6665 = ~pi354 & n62752;
  assign n6666 = ~n62480 & ~n6665;
  assign n6667 = ~n62480 & ~n6650;
  assign n6668 = ~n6665 & n6667;
  assign n6669 = ~n6650 & n6666;
  assign n6670 = pi354 & n62752;
  assign n6671 = ~pi354 & n62749;
  assign n6672 = n62480 & ~n6671;
  assign n6673 = n62480 & ~n6670;
  assign n6674 = ~n6671 & n6673;
  assign n6675 = ~n6670 & n6672;
  assign n6676 = ~pi591 & ~n62754;
  assign n6677 = ~n62753 & n6676;
  assign n6678 = ~pi591 & ~n62753;
  assign n6679 = ~n62754 & n6678;
  assign n6680 = ~n6625 & n6626;
  assign n6681 = n5543 & ~n62755;
  assign n6682 = ~pi588 & ~n6681;
  assign n6683 = ~pi588 & ~n62748;
  assign n6684 = ~n6681 & n6683;
  assign n6685 = ~n62748 & n6682;
  assign n6686 = pi592 & ~n2578;
  assign n6687 = n3132 & ~n5443;
  assign n6688 = ~n6686 & n6687;
  assign n6689 = n5541 & ~n6688;
  assign n6690 = ~n62332 & ~n6689;
  assign n6691 = n62332 & ~n6571;
  assign n6692 = ~n62332 & n6689;
  assign n6693 = n62332 & n6571;
  assign n6694 = ~n6692 & ~n6693;
  assign n6695 = ~pi428 & n6689;
  assign n6696 = pi428 & n6571;
  assign n6697 = ~pi427 & ~n6696;
  assign n6698 = ~pi428 & ~n6689;
  assign n6699 = pi428 & ~n6571;
  assign n6700 = ~n6698 & ~n6699;
  assign n6701 = ~pi427 & ~n6700;
  assign n6702 = ~n6695 & n6697;
  assign n6703 = pi428 & n6689;
  assign n6704 = ~pi428 & n6571;
  assign n6705 = pi427 & ~n6704;
  assign n6706 = pi428 & ~n6689;
  assign n6707 = ~pi428 & ~n6571;
  assign n6708 = ~n6706 & ~n6707;
  assign n6709 = pi427 & ~n6708;
  assign n6710 = ~n6703 & n6705;
  assign n6711 = ~n62758 & ~n62759;
  assign n6712 = ~n6690 & ~n6691;
  assign n6713 = n62331 & n62757;
  assign n6714 = ~n62332 & n6571;
  assign n6715 = n62332 & n6689;
  assign n6716 = n62332 & ~n6689;
  assign n6717 = ~n62332 & ~n6571;
  assign n6718 = ~n6716 & ~n6717;
  assign n6719 = ~pi427 & ~n6708;
  assign n6720 = pi427 & ~n6700;
  assign n6721 = ~n6719 & ~n6720;
  assign n6722 = ~n6714 & ~n6715;
  assign n6723 = ~n62331 & ~n62760;
  assign n6724 = ~n3414 & ~n6723;
  assign n6725 = ~n6713 & n6724;
  assign n6726 = n62331 & ~n62760;
  assign n6727 = ~n62331 & n62757;
  assign n6728 = n3414 & ~n6727;
  assign n6729 = ~n6726 & n6728;
  assign n6730 = pi1199 & ~n6729;
  assign n6731 = ~pi430 & ~n62760;
  assign n6732 = pi430 & n62757;
  assign n6733 = ~pi430 & n62760;
  assign n6734 = pi430 & ~n62757;
  assign n6735 = ~n6733 & ~n6734;
  assign n6736 = ~n6731 & ~n6732;
  assign n6737 = ~pi426 & n62761;
  assign n6738 = ~pi430 & n62757;
  assign n6739 = pi430 & ~n62760;
  assign n6740 = ~n6738 & ~n6739;
  assign n6741 = pi426 & ~n6740;
  assign n6742 = ~n6737 & ~n6741;
  assign n6743 = ~pi445 & ~n6742;
  assign n6744 = ~pi426 & ~n6740;
  assign n6745 = pi426 & n62761;
  assign n6746 = ~n6744 & ~n6745;
  assign n6747 = pi445 & ~n6746;
  assign n6748 = n62436 & ~n6747;
  assign n6749 = ~n6743 & n6748;
  assign n6750 = ~pi445 & ~n6746;
  assign n6751 = pi445 & ~n6742;
  assign n6752 = ~n62436 & ~n6751;
  assign n6753 = ~n6750 & n6752;
  assign n6754 = pi1199 & ~n6753;
  assign n6755 = ~n6749 & n6754;
  assign n6756 = ~n6743 & ~n6747;
  assign n6757 = ~pi448 & ~n6756;
  assign n6758 = ~n6750 & ~n6751;
  assign n6759 = pi448 & ~n6758;
  assign n6760 = ~n3269 & ~n6759;
  assign n6761 = ~n3269 & ~n6757;
  assign n6762 = ~n6759 & n6761;
  assign n6763 = ~n6757 & n6760;
  assign n6764 = pi448 & ~n6756;
  assign n6765 = ~pi448 & ~n6758;
  assign n6766 = n3269 & ~n6765;
  assign n6767 = n3269 & ~n6764;
  assign n6768 = ~n6765 & n6767;
  assign n6769 = ~n6764 & n6766;
  assign n6770 = pi1199 & ~n62764;
  assign n6771 = ~n62763 & n6770;
  assign n6772 = pi1199 & ~n62763;
  assign n6773 = ~n62764 & n6772;
  assign n6774 = ~n6725 & n6730;
  assign n6775 = ~pi1199 & ~n6689;
  assign n6776 = n3312 & ~n6775;
  assign n6777 = ~n62762 & n6776;
  assign n6778 = n6013 & ~n6777;
  assign n6779 = ~n3318 & ~n6778;
  assign n6780 = ~n62756 & n6779;
  assign n6781 = n3318 & n5541;
  assign n6782 = ~pi80 & ~n62455;
  assign n6783 = ~n6781 & n6782;
  assign n6784 = ~n6780 & n6783;
  assign n6785 = ~pi217 & ~n6784;
  assign n6786 = ~n62741 & n6785;
  assign n6787 = ~pi80 & ~n5541;
  assign n6788 = pi217 & ~n6787;
  assign n6789 = n5530 & ~n6788;
  assign po238 = ~n6786 & n6789;
  assign n6791 = ~pi87 & ~pi100;
  assign n6792 = ~pi54 & ~pi74;
  assign n6793 = ~pi75 & ~pi92;
  assign n6794 = n6792 & n6793;
  assign n6795 = ~pi75 & ~pi87;
  assign n6796 = ~pi92 & n6795;
  assign n6797 = n6792 & n6796;
  assign n6798 = ~pi100 & n6797;
  assign n6799 = n6791 & n6794;
  assign n6800 = pi140 & ~n62765;
  assign n6801 = pi40 & ~n62383;
  assign n6802 = n2727 & ~n6801;
  assign n6803 = n2687 & n5546;
  assign n6804 = ~pi66 & ~pi84;
  assign n6805 = n2616 & n6804;
  assign n6806 = ~pi36 & ~pi67;
  assign n6807 = ~pi103 & n6806;
  assign n6808 = n6805 & n6807;
  assign n6809 = ~pi68 & ~pi73;
  assign n6810 = ~pi69 & ~pi83;
  assign n6811 = n2620 & n6810;
  assign n6812 = n6809 & n6811;
  assign n6813 = n6808 & n6812;
  assign n6814 = pi45 & n2587;
  assign n6815 = pi45 & n2598;
  assign n6816 = n2587 & n6815;
  assign n6817 = n2598 & n6814;
  assign n6818 = n6813 & n62766;
  assign n6819 = n2595 & n6818;
  assign n6820 = ~pi102 & ~n6819;
  assign n6821 = pi102 & ~n2633;
  assign n6822 = ~pi98 & ~n6821;
  assign n6823 = ~n6820 & n6822;
  assign n6824 = n6803 & n6823;
  assign n6825 = ~pi96 & n2696;
  assign n6826 = n2695 & n2771;
  assign n6827 = n2772 & n62767;
  assign n6828 = ~pi93 & n62382;
  assign n6829 = ~pi35 & ~pi51;
  assign n6830 = ~pi96 & n2743;
  assign n6831 = n2771 & n6829;
  assign n6832 = ~pi72 & ~pi93;
  assign n6833 = n62770 & n6832;
  assign n6834 = n2719 & n62375;
  assign n6835 = ~pi90 & n62769;
  assign n6836 = n2694 & n62382;
  assign n6837 = n62355 & n62768;
  assign n6838 = n6824 & n6837;
  assign n6839 = ~pi40 & ~n6838;
  assign n6840 = n6802 & ~n6839;
  assign n6841 = ~pi252 & ~n6840;
  assign n6842 = pi35 & ~n62369;
  assign n6843 = n62375 & ~n6842;
  assign n6844 = ~pi40 & n6843;
  assign n6845 = pi47 & n62349;
  assign n6846 = n62353 & n6845;
  assign n6847 = pi47 & ~n6846;
  assign n6848 = n2663 & ~n6847;
  assign n6849 = ~pi91 & ~n6847;
  assign n6850 = n2715 & n6849;
  assign n6851 = n2694 & n6848;
  assign n6852 = n62351 & n6824;
  assign n6853 = ~pi47 & ~n6852;
  assign n6854 = ~pi97 & n62389;
  assign n6855 = pi108 & ~pi110;
  assign n6856 = pi108 & n2642;
  assign n6857 = n2867 & n6855;
  assign n6858 = n6854 & n62772;
  assign n6859 = pi314 & n6858;
  assign n6860 = n6853 & ~n6859;
  assign n6861 = n62771 & ~n6860;
  assign n6862 = ~pi35 & ~n6861;
  assign n6863 = n6844 & ~n6862;
  assign n6864 = pi40 & n62383;
  assign n6865 = pi252 & ~n6864;
  assign n6866 = ~n6863 & n6865;
  assign n6867 = ~n6841 & ~n6866;
  assign n6868 = n2727 & n6867;
  assign n6869 = pi1092 & ~n3112;
  assign n6870 = pi1092 & n6868;
  assign n6871 = ~n3112 & n6870;
  assign n6872 = n6868 & n6869;
  assign n6873 = ~pi98 & n62358;
  assign n6874 = pi88 & ~n6873;
  assign n6875 = n2687 & ~n6874;
  assign n6876 = ~pi88 & ~n6823;
  assign n6877 = n6875 & ~n6876;
  assign n6878 = n62353 & n6877;
  assign n6879 = ~pi47 & ~n6859;
  assign n6880 = ~pi47 & ~n6878;
  assign n6881 = ~n6859 & n6880;
  assign n6882 = ~n6878 & n6879;
  assign n6883 = n62771 & ~n62774;
  assign n6884 = ~pi35 & ~n6883;
  assign n6885 = pi252 & n6843;
  assign n6886 = ~n6884 & n6885;
  assign n6887 = n2638 & n6837;
  assign n6888 = n62356 & n62768;
  assign n6889 = ~pi252 & n62775;
  assign n6890 = n6877 & n6889;
  assign n6891 = ~pi40 & ~n6890;
  assign n6892 = ~n6886 & n6891;
  assign n6893 = n2852 & n6802;
  assign n6894 = ~n6892 & n6893;
  assign n6895 = ~n62773 & ~n6894;
  assign n6896 = pi1093 & ~n6895;
  assign n6897 = ~n2824 & ~n6896;
  assign po1106 = n2824 & n62394;
  assign n6899 = n2824 & n2924;
  assign n6900 = n6870 & n6899;
  assign n6901 = n6868 & po1106;
  assign n6902 = ~n2929 & ~n62776;
  assign n6903 = ~n6897 & ~n6902;
  assign n6904 = ~pi1091 & n6896;
  assign n6905 = ~n6903 & ~n6904;
  assign n6906 = ~pi210 & n6905;
  assign n6907 = ~n6801 & ~n6892;
  assign n6908 = ~pi32 & ~n6907;
  assign n6909 = n2730 & n2746;
  assign n6910 = pi32 & ~n6909;
  assign n6911 = ~pi95 & ~n6910;
  assign n6912 = ~pi95 & n2582;
  assign n6913 = ~n6910 & n6912;
  assign n6914 = pi824 & n6913;
  assign n6915 = n2852 & n6911;
  assign n6916 = ~n6908 & n6913;
  assign n6917 = pi824 & n6916;
  assign n6918 = ~n6908 & n62777;
  assign n6919 = ~n62773 & ~n62778;
  assign n6920 = ~pi32 & ~n6867;
  assign n6921 = ~pi824 & n2582;
  assign n6922 = ~pi824 & n6913;
  assign n6923 = n6911 & n6921;
  assign n6924 = ~n6920 & n62779;
  assign n6925 = n6913 & ~n6920;
  assign n6926 = ~pi824 & pi829;
  assign n6927 = n6925 & n6926;
  assign n6928 = pi829 & n6924;
  assign n6929 = n6919 & ~n62780;
  assign n6930 = pi1093 & ~n6929;
  assign n6931 = ~n2824 & ~n6930;
  assign n6932 = ~n6902 & ~n6931;
  assign n6933 = n3032 & ~n6919;
  assign n6934 = ~n6932 & ~n6933;
  assign n6935 = pi210 & n6934;
  assign n6936 = ~n6906 & ~n6935;
  assign n6937 = pi299 & ~n6936;
  assign n6938 = ~pi198 & n6905;
  assign n6939 = pi198 & n6934;
  assign n6940 = ~n6938 & ~n6939;
  assign n6941 = ~pi299 & ~n6940;
  assign n6942 = ~pi299 & n6940;
  assign n6943 = pi299 & n6936;
  assign n6944 = ~n6942 & ~n6943;
  assign n6945 = ~n6937 & ~n6941;
  assign n6946 = ~pi39 & ~n62781;
  assign n6947 = n2933 & ~n2937;
  assign n6948 = ~pi120 & ~n6947;
  assign n6949 = pi120 & ~n62380;
  assign n6950 = ~n6948 & ~n6949;
  assign n6951 = n2923 & n6950;
  assign n6952 = ~n2814 & n6951;
  assign n6953 = n2923 & n6947;
  assign n6954 = ~pi120 & ~n6953;
  assign n6955 = n62380 & n2923;
  assign n6956 = ~pi287 & n2937;
  assign n6957 = pi835 & pi950;
  assign n6958 = n6956 & n6957;
  assign n6959 = ~n2583 & ~n2824;
  assign n6960 = n6958 & n6959;
  assign n6961 = n6955 & ~n6960;
  assign n6962 = pi120 & ~n6961;
  assign n6963 = pi1091 & ~n6962;
  assign n6964 = ~n6954 & n6963;
  assign n6965 = pi120 & ~n6955;
  assign n6966 = ~pi1091 & ~n6965;
  assign n6967 = pi120 & pi824;
  assign n6968 = n6958 & n6967;
  assign n6969 = n6966 & ~n6968;
  assign n6970 = ~n6954 & n6969;
  assign n6971 = ~n6964 & ~n6970;
  assign n6972 = n2814 & ~n6971;
  assign n6973 = ~n6952 & ~n6972;
  assign n6974 = ~n2904 & n6973;
  assign n6975 = n2904 & n6971;
  assign n6976 = ~n2902 & ~n6951;
  assign n6977 = n2814 & ~n6951;
  assign n6978 = ~n2814 & n6971;
  assign n6979 = ~n6977 & ~n6978;
  assign n6980 = n2902 & ~n6979;
  assign n6981 = ~n6976 & ~n6980;
  assign n6982 = ~pi614 & ~n6981;
  assign n6983 = ~pi616 & n6982;
  assign n6984 = n2903 & ~n6981;
  assign n6985 = ~n6973 & ~n62782;
  assign n6986 = ~n6974 & ~n6975;
  assign n6987 = pi681 & ~n62783;
  assign n6988 = pi616 & ~n6951;
  assign n6989 = pi614 & ~n6951;
  assign n6990 = ~n6982 & ~n6989;
  assign n6991 = ~pi616 & ~n6990;
  assign n6992 = ~n6988 & ~n6991;
  assign n6993 = ~n2905 & ~n6992;
  assign n6994 = n2905 & n6971;
  assign n6995 = ~n2814 & ~n6994;
  assign n6996 = ~n6993 & n6995;
  assign n6997 = ~n6972 & ~n6996;
  assign n6998 = ~pi661 & ~n6997;
  assign n6999 = pi661 & n62783;
  assign n7000 = ~pi681 & ~n6999;
  assign n7001 = ~n6998 & n7000;
  assign n7002 = ~n6987 & ~n7001;
  assign n7003 = ~n2971 & ~n7002;
  assign n7004 = n2907 & n6979;
  assign n7005 = ~n2907 & n6992;
  assign n7006 = pi681 & ~n6992;
  assign n7007 = ~pi661 & ~pi681;
  assign n7008 = ~pi662 & n7007;
  assign n7009 = ~pi616 & ~n7008;
  assign n7010 = n6990 & n7009;
  assign n7011 = ~pi680 & n6991;
  assign n7012 = pi680 & ~n6979;
  assign n7013 = ~pi616 & n7008;
  assign n7014 = ~n7012 & n7013;
  assign n7015 = ~n7011 & n7014;
  assign n7016 = ~n7010 & ~n7015;
  assign n7017 = ~pi680 & ~n6951;
  assign n7018 = pi616 & n7008;
  assign n7019 = ~n7017 & n7018;
  assign n7020 = ~n7012 & n7019;
  assign n7021 = pi616 & n6951;
  assign n7022 = ~n7008 & n7021;
  assign n7023 = ~n7020 & ~n7022;
  assign n7024 = ~pi681 & n7023;
  assign n7025 = n7016 & n7024;
  assign n7026 = ~n7006 & ~n7025;
  assign n7027 = ~n7004 & ~n7005;
  assign n7028 = n2971 & ~n62784;
  assign n7029 = ~n2971 & n7002;
  assign n7030 = n2971 & n62784;
  assign n7031 = ~n7029 & ~n7030;
  assign n7032 = ~n7003 & ~n7028;
  assign n7033 = pi223 & n62785;
  assign n7034 = ~pi222 & ~pi224;
  assign n7035 = n2824 & n6953;
  assign n7036 = ~pi824 & ~n6947;
  assign n7037 = ~pi984 & ~n2582;
  assign n7038 = pi835 & ~n7037;
  assign n7039 = n2936 & ~n7038;
  assign n7040 = n2933 & ~n7039;
  assign n7041 = pi1092 & n7040;
  assign n7042 = ~n6921 & ~n7041;
  assign n7043 = ~n7036 & ~n7042;
  assign n7044 = ~pi829 & ~n7043;
  assign n7045 = pi829 & ~n7041;
  assign n7046 = n2851 & ~n7045;
  assign n7047 = ~n7044 & n7046;
  assign n7048 = ~n7035 & ~n7047;
  assign n7049 = pi1091 & ~n7048;
  assign n7050 = ~pi120 & ~n7049;
  assign n7051 = ~n6965 & ~n7050;
  assign n7052 = pi1093 & n7043;
  assign n7053 = ~pi120 & ~n7052;
  assign n7054 = n6966 & ~n7053;
  assign n7055 = ~n7051 & ~n7054;
  assign n7056 = n2814 & ~n7055;
  assign n7057 = ~n6952 & ~n7056;
  assign n7058 = ~n2904 & n7057;
  assign n7059 = n2904 & n7055;
  assign n7060 = n2904 & ~n7055;
  assign n7061 = ~n2904 & ~n7057;
  assign n7062 = ~n7060 & ~n7061;
  assign n7063 = ~n7058 & ~n7059;
  assign n7064 = ~n2907 & n62786;
  assign n7065 = n2907 & n7055;
  assign n7066 = ~n2906 & ~n62786;
  assign n7067 = n2906 & ~n7055;
  assign n7068 = ~pi681 & ~n7067;
  assign n7069 = ~n7066 & n7068;
  assign n7070 = pi681 & n62786;
  assign n7071 = ~n7069 & ~n7070;
  assign n7072 = ~n7064 & ~n7065;
  assign n7073 = ~n2971 & n62787;
  assign n7074 = ~pi603 & ~n6951;
  assign n7075 = ~n2814 & n7055;
  assign n7076 = ~n6977 & ~n7075;
  assign n7077 = pi603 & ~n7076;
  assign n7078 = ~n7074 & ~n7077;
  assign n7079 = ~pi642 & ~n7078;
  assign n7080 = ~n6976 & ~n7079;
  assign n7081 = ~pi614 & ~n7080;
  assign n7082 = ~n6989 & ~n7081;
  assign n7083 = ~pi616 & ~n7082;
  assign n7084 = ~n6988 & ~n7083;
  assign n7085 = pi681 & ~n7084;
  assign n7086 = ~pi616 & ~n7080;
  assign n7087 = ~pi614 & ~n2907;
  assign n7088 = ~n6988 & n7087;
  assign n7089 = ~n6988 & ~n7086;
  assign n7090 = n7087 & n7089;
  assign n7091 = ~n7086 & n7088;
  assign n7092 = ~pi614 & n2907;
  assign n7093 = n7076 & n7092;
  assign n7094 = ~n62788 & ~n7093;
  assign n7095 = pi680 & ~n7076;
  assign n7096 = pi614 & n7008;
  assign n7097 = ~n7017 & n7096;
  assign n7098 = ~n7095 & n7097;
  assign n7099 = pi614 & n6951;
  assign n7100 = ~n7008 & n7099;
  assign n7101 = ~n7098 & ~n7100;
  assign n7102 = ~pi681 & n7101;
  assign n7103 = n7094 & n7102;
  assign n7104 = ~n7085 & ~n7103;
  assign n7105 = n2971 & n7104;
  assign n7106 = n2971 & ~n7104;
  assign n7107 = ~n2971 & ~n62787;
  assign n7108 = ~n7106 & ~n7107;
  assign n7109 = ~n7073 & ~n7105;
  assign n7110 = ~n7034 & n62789;
  assign n7111 = n6950 & n7034;
  assign n7112 = n6955 & n7111;
  assign n7113 = n6951 & n7034;
  assign n7114 = ~pi223 & ~n62790;
  assign n7115 = ~n7110 & n7114;
  assign n7116 = ~n7033 & ~n7115;
  assign n7117 = ~pi299 & ~n7116;
  assign n7118 = ~pi216 & ~pi221;
  assign n7119 = n2914 & ~n7104;
  assign n7120 = ~n2914 & ~n62787;
  assign n7121 = n2915 & ~n7120;
  assign n7122 = ~n7119 & n7121;
  assign n7123 = ~n7118 & n7122;
  assign n7124 = ~n2915 & n62787;
  assign n7125 = ~n7118 & n7124;
  assign n7126 = n6951 & n7118;
  assign n7127 = ~pi215 & ~n7126;
  assign n7128 = ~n6951 & n7118;
  assign n7129 = ~n7118 & ~n7124;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = ~pi215 & ~n7130;
  assign n7132 = ~n7125 & n7127;
  assign n7133 = ~n7123 & n62791;
  assign n7134 = ~n2915 & n7002;
  assign n7135 = ~n2914 & ~n7002;
  assign n7136 = n2914 & ~n62784;
  assign n7137 = n2915 & ~n7136;
  assign n7138 = ~n7135 & n7137;
  assign n7139 = ~n7134 & ~n7138;
  assign n7140 = pi215 & n7139;
  assign n7141 = ~n7133 & ~n7140;
  assign n7142 = pi299 & ~n7141;
  assign n7143 = ~n7117 & ~n7142;
  assign n7144 = pi39 & n7143;
  assign n7145 = ~pi39 & n62781;
  assign n7146 = pi39 & ~n7143;
  assign n7147 = ~n7145 & ~n7146;
  assign n7148 = ~n6946 & ~n7144;
  assign n7149 = pi761 & n62792;
  assign n7150 = pi621 & n6903;
  assign n7151 = ~pi198 & ~n7150;
  assign n7152 = pi621 & n6932;
  assign n7153 = pi198 & ~n7152;
  assign n7154 = ~n7151 & ~n7153;
  assign n7155 = pi621 & ~n6904;
  assign n7156 = ~n6905 & ~n7155;
  assign n7157 = ~pi198 & n7156;
  assign n7158 = pi621 & ~n6933;
  assign n7159 = ~n6934 & ~n7158;
  assign n7160 = pi198 & n7159;
  assign n7161 = ~n7157 & ~n7160;
  assign n7162 = ~pi603 & ~n7161;
  assign n7163 = ~n7154 & ~n7162;
  assign n7164 = ~pi299 & ~n7163;
  assign n7165 = ~pi210 & ~n7150;
  assign n7166 = pi210 & ~n7152;
  assign n7167 = ~n7165 & ~n7166;
  assign n7168 = pi603 & ~n7167;
  assign n7169 = n6936 & ~n7168;
  assign n7170 = pi299 & n7169;
  assign n7171 = pi299 & ~n7169;
  assign n7172 = ~pi299 & n7163;
  assign n7173 = ~n7171 & ~n7172;
  assign n7174 = ~n7164 & ~n7170;
  assign n7175 = ~pi39 & n62793;
  assign n7176 = pi621 & pi1091;
  assign n7177 = n6951 & n7176;
  assign n7178 = n2814 & ~n7177;
  assign n7179 = n7051 & n7176;
  assign n7180 = ~n2814 & ~n7179;
  assign n7181 = ~n7178 & ~n7180;
  assign n7182 = pi603 & ~n7181;
  assign n7183 = n7076 & ~n7182;
  assign n7184 = n2907 & ~n7183;
  assign n7185 = ~pi614 & ~pi642;
  assign n7186 = ~pi616 & n7185;
  assign n7187 = pi603 & ~n7176;
  assign n7188 = n6951 & ~n7187;
  assign n7189 = ~n7186 & n7188;
  assign n7190 = ~n7074 & n7186;
  assign n7191 = ~n7182 & n7190;
  assign n7192 = ~n7189 & ~n7191;
  assign n7193 = ~n2907 & n7192;
  assign n7194 = ~n7184 & ~n7193;
  assign n7195 = n62393 & ~n7194;
  assign n7196 = pi621 & ~n7054;
  assign n7197 = ~n7055 & ~n7196;
  assign n7198 = ~pi603 & n7197;
  assign n7199 = ~n7179 & ~n7198;
  assign n7200 = n62787 & ~n7199;
  assign n7201 = ~n62393 & ~n7200;
  assign n7202 = ~n7118 & ~n7201;
  assign n7203 = ~n62393 & n7200;
  assign n7204 = n62393 & n7194;
  assign n7205 = ~n7203 & ~n7204;
  assign n7206 = ~n7118 & ~n7205;
  assign n7207 = ~n7118 & ~n7195;
  assign n7208 = ~n7201 & n7207;
  assign n7209 = ~n7195 & n7202;
  assign n7210 = n7118 & n7188;
  assign n7211 = n7126 & ~n7187;
  assign n7212 = ~pi215 & ~n62795;
  assign n7213 = ~n62794 & n7212;
  assign n7214 = pi621 & n6964;
  assign n7215 = ~n2814 & ~n7214;
  assign n7216 = ~n7178 & ~n7215;
  assign n7217 = pi603 & ~n7216;
  assign n7218 = n7004 & ~n7217;
  assign n7219 = n7190 & ~n7217;
  assign n7220 = ~n7189 & ~n7219;
  assign n7221 = ~n2907 & ~n7220;
  assign n7222 = ~n7218 & ~n7221;
  assign n7223 = n62393 & ~n7222;
  assign n7224 = n2923 & ~n7187;
  assign n7225 = ~n6973 & n7224;
  assign n7226 = n2904 & ~n6964;
  assign n7227 = n7225 & ~n7226;
  assign n7228 = ~n2907 & ~n7227;
  assign n7229 = ~n6971 & n7224;
  assign n7230 = pi680 & ~n7229;
  assign n7231 = n7008 & n7230;
  assign n7232 = n2907 & ~n7229;
  assign n7233 = ~n7228 & ~n62796;
  assign n7234 = ~n62393 & n7233;
  assign n7235 = pi215 & ~n7234;
  assign n7236 = ~n7223 & n7235;
  assign n7237 = ~n62794 & ~n62795;
  assign n7238 = ~pi215 & ~n7237;
  assign n7239 = n62393 & n7222;
  assign n7240 = ~n62393 & ~n7233;
  assign n7241 = pi215 & ~n7240;
  assign n7242 = ~n7239 & n7241;
  assign n7243 = ~n7238 & ~n7242;
  assign n7244 = ~n7213 & ~n7236;
  assign n7245 = pi299 & ~n62797;
  assign n7246 = n2971 & ~n7194;
  assign n7247 = ~n2971 & ~n7200;
  assign n7248 = ~n7034 & ~n7247;
  assign n7249 = n2971 & n7194;
  assign n7250 = ~n2971 & n7200;
  assign n7251 = ~n7249 & ~n7250;
  assign n7252 = ~n7034 & ~n7251;
  assign n7253 = ~n7034 & ~n7246;
  assign n7254 = ~n7247 & n7253;
  assign n7255 = ~n7246 & n7248;
  assign n7256 = n7034 & n7188;
  assign n7257 = n62790 & ~n7187;
  assign n7258 = ~pi223 & ~n62799;
  assign n7259 = ~n62798 & n7258;
  assign n7260 = n2971 & ~n7222;
  assign n7261 = ~n2971 & n7233;
  assign n7262 = pi223 & ~n7261;
  assign n7263 = ~n7260 & n7262;
  assign n7264 = ~n62798 & ~n62799;
  assign n7265 = ~pi223 & ~n7264;
  assign n7266 = n2971 & n7222;
  assign n7267 = ~n2971 & ~n7233;
  assign n7268 = pi223 & ~n7267;
  assign n7269 = ~n7266 & n7268;
  assign n7270 = ~n7265 & ~n7269;
  assign n7271 = ~n7259 & ~n7263;
  assign n7272 = ~pi299 & ~n62800;
  assign n7273 = pi299 & n62797;
  assign n7274 = ~pi299 & n62800;
  assign n7275 = ~n7273 & ~n7274;
  assign n7276 = ~n7245 & ~n7272;
  assign n7277 = pi39 & n62801;
  assign n7278 = ~pi39 & ~n62793;
  assign n7279 = pi39 & ~n62801;
  assign n7280 = ~n7278 & ~n7279;
  assign n7281 = ~n7175 & ~n7277;
  assign n7282 = ~pi761 & n62802;
  assign n7283 = ~pi140 & ~n7282;
  assign n7284 = ~n7149 & n7283;
  assign n7285 = pi603 & ~n7161;
  assign n7286 = ~pi299 & ~n7285;
  assign n7287 = ~pi210 & ~n7156;
  assign n7288 = pi210 & ~n7159;
  assign n7289 = ~n7287 & ~n7288;
  assign n7290 = pi603 & n7289;
  assign n7291 = pi299 & ~n7290;
  assign n7292 = ~n7286 & ~n7291;
  assign n7293 = ~pi39 & ~n7292;
  assign n7294 = n62787 & n7187;
  assign n7295 = ~n62393 & ~n7294;
  assign n7296 = n7076 & n7187;
  assign n7297 = n2907 & ~n7296;
  assign n7298 = n6951 & n7187;
  assign n7299 = ~n7186 & n7298;
  assign n7300 = n7186 & n7296;
  assign n7301 = n7186 & ~n7296;
  assign n7302 = ~n7186 & ~n7298;
  assign n7303 = ~n7301 & ~n7302;
  assign n7304 = ~n7299 & ~n7300;
  assign n7305 = ~n2907 & ~n62803;
  assign n7306 = n2907 & n7296;
  assign n7307 = ~n2907 & n62803;
  assign n7308 = ~n7306 & ~n7307;
  assign n7309 = ~n7297 & ~n7305;
  assign n7310 = n62393 & n62804;
  assign n7311 = ~n7118 & ~n7310;
  assign n7312 = ~n7118 & ~n7295;
  assign n7313 = ~n7310 & n7312;
  assign n7314 = ~n7295 & n7311;
  assign n7315 = n6950 & n7118;
  assign n7316 = n2923 & n7187;
  assign n7317 = n7126 & n7187;
  assign n7318 = n7118 & n7298;
  assign n7319 = n7315 & n7316;
  assign n7320 = ~pi215 & ~n62806;
  assign n7321 = ~n62805 & n7320;
  assign n7322 = ~n6978 & n7298;
  assign n7323 = ~n6973 & n7298;
  assign n7324 = n6978 & n7186;
  assign n7325 = n7323 & ~n7324;
  assign n7326 = ~n2907 & n7325;
  assign n7327 = ~n7322 & ~n7326;
  assign n7328 = ~n62393 & n6973;
  assign n7329 = ~n7327 & ~n7328;
  assign n7330 = pi215 & ~n7329;
  assign n7331 = pi299 & ~n7330;
  assign n7332 = ~n7321 & n7331;
  assign n7333 = n7034 & n7298;
  assign n7334 = n62790 & n7187;
  assign n7335 = n7111 & n7316;
  assign n7336 = ~pi223 & ~n62807;
  assign n7337 = n2971 & n62804;
  assign n7338 = ~n2971 & ~n7294;
  assign n7339 = ~n7034 & ~n7338;
  assign n7340 = ~n7034 & ~n7337;
  assign n7341 = ~n7338 & n7340;
  assign n7342 = ~n7337 & n7339;
  assign n7343 = n7336 & ~n62808;
  assign n7344 = ~n2971 & n6973;
  assign n7345 = ~n7327 & ~n7344;
  assign n7346 = pi223 & ~n7345;
  assign n7347 = ~pi299 & ~n7346;
  assign n7348 = ~n7343 & n7347;
  assign n7349 = ~n7332 & ~n7348;
  assign n7350 = pi39 & n7349;
  assign n7351 = ~n7293 & ~n7350;
  assign n7352 = pi140 & ~pi761;
  assign n7353 = n7351 & n7352;
  assign n7354 = ~n7284 & ~n7353;
  assign n7355 = ~pi38 & ~n7354;
  assign n7356 = ~pi39 & n62380;
  assign n7357 = n2923 & n7356;
  assign n7358 = ~pi140 & ~n7357;
  assign n7359 = n7316 & n7356;
  assign n7360 = ~pi761 & n7359;
  assign n7361 = ~n7358 & ~n7360;
  assign n7362 = pi38 & ~n7361;
  assign n7363 = ~n7355 & ~n7362;
  assign n7364 = pi738 & ~n7363;
  assign n7365 = pi680 & ~n7008;
  assign n7366 = pi665 & pi1091;
  assign n7367 = ~n7187 & ~n7366;
  assign n7368 = n6951 & ~n7367;
  assign n7369 = pi616 & ~n7368;
  assign n7370 = pi614 & ~n7368;
  assign n7371 = pi642 & ~n7368;
  assign n7372 = n7078 & ~n7367;
  assign n7373 = ~pi642 & ~n7372;
  assign n7374 = ~n7371 & ~n7373;
  assign n7375 = ~pi614 & ~n7374;
  assign n7376 = ~n7370 & ~n7375;
  assign n7377 = ~pi616 & ~n7376;
  assign n7378 = ~n7369 & ~n7377;
  assign n7379 = n7365 & ~n7378;
  assign n7380 = ~pi680 & ~n7084;
  assign n7381 = n6951 & n7366;
  assign n7382 = n2814 & ~n7381;
  assign n7383 = n7051 & n7366;
  assign n7384 = ~n2814 & ~n7383;
  assign n7385 = ~n7382 & ~n7384;
  assign n7386 = ~pi603 & ~n7385;
  assign n7387 = pi603 & ~pi665;
  assign n7388 = n7176 & n7387;
  assign n7389 = ~n7077 & ~n7388;
  assign n7390 = ~n7386 & n7389;
  assign n7391 = n2907 & ~n7390;
  assign n7392 = ~n7380 & ~n7391;
  assign n7393 = ~n7379 & n7392;
  assign n7394 = n2971 & n7393;
  assign n7395 = ~n62786 & ~n7367;
  assign n7396 = n7365 & ~n7395;
  assign n7397 = ~pi680 & n62786;
  assign n7398 = pi603 & n7197;
  assign n7399 = pi603 & ~pi621;
  assign n7400 = n7383 & ~n7399;
  assign n7401 = n2907 & ~n7400;
  assign n7402 = ~n7398 & n7401;
  assign n7403 = ~n7397 & ~n7402;
  assign n7404 = ~n7396 & n7403;
  assign n7405 = ~n2971 & n7404;
  assign n7406 = ~n7034 & ~n7405;
  assign n7407 = ~n7394 & n7406;
  assign n7408 = pi680 & n7367;
  assign n7409 = n6951 & ~n7408;
  assign n7410 = n7034 & ~n7409;
  assign n7411 = ~pi223 & ~n7410;
  assign n7412 = n2971 & ~n7393;
  assign n7413 = ~n2971 & ~n7404;
  assign n7414 = ~n7034 & ~n7413;
  assign n7415 = ~n7394 & ~n7405;
  assign n7416 = ~n7034 & ~n7415;
  assign n7417 = ~n7412 & n7414;
  assign n7418 = n7034 & ~n7408;
  assign n7419 = n7034 & n7409;
  assign n7420 = n6951 & n7418;
  assign n7421 = ~n62809 & ~n62810;
  assign n7422 = ~pi223 & ~n7421;
  assign n7423 = ~n7407 & n7411;
  assign n7424 = pi665 & n6964;
  assign n7425 = ~n6971 & n7298;
  assign n7426 = ~n7424 & ~n7425;
  assign n7427 = n6952 & n7366;
  assign n7428 = ~pi603 & n7427;
  assign n7429 = n7426 & ~n7428;
  assign n7430 = ~n2814 & ~n7424;
  assign n7431 = ~n7382 & ~n7430;
  assign n7432 = ~pi642 & ~n7431;
  assign n7433 = ~pi642 & ~n7322;
  assign n7434 = ~n7431 & n7433;
  assign n7435 = ~n7322 & n7432;
  assign n7436 = n7429 & n62812;
  assign n7437 = ~n7371 & ~n7436;
  assign n7438 = ~pi614 & ~n7437;
  assign n7439 = ~n7370 & ~n7438;
  assign n7440 = ~pi616 & ~n7439;
  assign n7441 = ~n7369 & ~n7440;
  assign n7442 = n7365 & ~n7441;
  assign n7443 = ~pi680 & ~n6992;
  assign n7444 = n2907 & ~n7431;
  assign n7445 = ~n7322 & n7444;
  assign n7446 = ~n7443 & ~n7445;
  assign n7447 = ~n7442 & n7446;
  assign n7448 = n2971 & ~n7447;
  assign n7449 = ~n7424 & ~n7427;
  assign n7450 = ~n7323 & n7449;
  assign n7451 = ~n7186 & n7450;
  assign n7452 = n7186 & n7429;
  assign n7453 = ~n7451 & ~n7452;
  assign n7454 = n7365 & ~n7453;
  assign n7455 = ~pi680 & ~n62783;
  assign n7456 = n2907 & n7426;
  assign n7457 = ~n7455 & ~n7456;
  assign n7458 = ~n7454 & ~n7456;
  assign n7459 = ~n7455 & n7458;
  assign n7460 = ~n7454 & n7457;
  assign n7461 = ~n2971 & ~n62813;
  assign n7462 = pi223 & ~n7461;
  assign n7463 = ~n7448 & n7462;
  assign n7464 = ~pi223 & ~n62810;
  assign n7465 = ~n62809 & n7464;
  assign n7466 = n2971 & n7447;
  assign n7467 = ~n2971 & n62813;
  assign n7468 = pi223 & ~n7467;
  assign n7469 = ~n7466 & n7468;
  assign n7470 = ~n7465 & ~n7469;
  assign n7471 = ~n62811 & ~n7463;
  assign n7472 = ~pi299 & n62814;
  assign n7473 = n62393 & n7393;
  assign n7474 = ~n62393 & n7404;
  assign n7475 = ~n7118 & ~n7474;
  assign n7476 = n62393 & ~n7393;
  assign n7477 = ~n62393 & ~n7404;
  assign n7478 = ~n7473 & ~n7474;
  assign n7479 = ~n7476 & ~n7477;
  assign n7480 = ~n7118 & n62815;
  assign n7481 = ~n7473 & n7475;
  assign n7482 = n7118 & ~n7409;
  assign n7483 = ~pi215 & ~n7482;
  assign n7484 = n7118 & n7409;
  assign n7485 = n7126 & ~n7408;
  assign n7486 = ~n7118 & ~n7477;
  assign n7487 = ~n7118 & ~n62815;
  assign n7488 = ~n7476 & n7486;
  assign n7489 = ~n62817 & ~n62818;
  assign n7490 = ~pi215 & ~n7489;
  assign n7491 = ~n62816 & n7483;
  assign n7492 = n62393 & ~n7447;
  assign n7493 = ~n62393 & ~n62813;
  assign n7494 = pi215 & ~n7493;
  assign n7495 = ~n7492 & n7494;
  assign n7496 = ~pi215 & ~n62817;
  assign n7497 = ~n62818 & n7496;
  assign n7498 = n62393 & n7447;
  assign n7499 = ~n62393 & n62813;
  assign n7500 = pi215 & ~n7499;
  assign n7501 = ~n7498 & n7500;
  assign n7502 = ~n7497 & ~n7501;
  assign n7503 = ~n62819 & ~n7495;
  assign n7504 = pi299 & n62820;
  assign n7505 = ~pi299 & ~n62814;
  assign n7506 = pi299 & ~n62820;
  assign n7507 = ~n7505 & ~n7506;
  assign n7508 = ~n7472 & ~n7504;
  assign n7509 = ~pi140 & ~n62821;
  assign n7510 = ~pi665 & n7051;
  assign n7511 = pi665 & ~n7054;
  assign n7512 = ~n7055 & ~n7511;
  assign n7513 = ~n7054 & ~n7510;
  assign n7514 = ~pi603 & n7057;
  assign n7515 = n2814 & n7179;
  assign n7516 = n6952 & n7176;
  assign n7517 = pi603 & ~n7516;
  assign n7518 = n2814 & n7051;
  assign n7519 = ~n6952 & ~n7518;
  assign n7520 = pi603 & n7519;
  assign n7521 = ~n7187 & ~n7520;
  assign n7522 = ~n7515 & n7517;
  assign n7523 = ~n7514 & n62823;
  assign n7524 = n62822 & n7523;
  assign n7525 = pi616 & ~n7524;
  assign n7526 = ~n7185 & n7524;
  assign n7527 = ~n7057 & n62822;
  assign n7528 = ~pi603 & ~n7527;
  assign n7529 = ~pi665 & n7179;
  assign n7530 = n7176 & n7510;
  assign n7531 = pi603 & ~n62824;
  assign n7532 = ~n7528 & ~n7531;
  assign n7533 = n7185 & n7532;
  assign n7534 = ~pi616 & ~n7533;
  assign n7535 = ~n7524 & n7534;
  assign n7536 = ~n7526 & n7534;
  assign n7537 = ~n7525 & ~n62825;
  assign n7538 = ~n7008 & ~n7537;
  assign n7539 = n2907 & n62822;
  assign n7540 = ~n7531 & n7539;
  assign n7541 = ~n7365 & ~n7540;
  assign n7542 = ~n7538 & ~n7541;
  assign n7543 = ~n62393 & ~n7542;
  assign n7544 = n6951 & ~n7366;
  assign n7545 = ~n7187 & n7544;
  assign n7546 = n7188 & ~n7366;
  assign n7547 = pi616 & ~n62826;
  assign n7548 = n7365 & ~n7547;
  assign n7549 = pi603 & pi665;
  assign n7550 = ~pi603 & ~n7544;
  assign n7551 = ~n7549 & ~n7550;
  assign n7552 = ~n7182 & n7551;
  assign n7553 = n7185 & n7552;
  assign n7554 = ~n7185 & n62826;
  assign n7555 = ~pi616 & ~n7554;
  assign n7556 = ~n7553 & n7555;
  assign n7557 = n7548 & ~n7556;
  assign n7558 = n7076 & n7391;
  assign n7559 = ~n7557 & ~n7558;
  assign n7560 = n62393 & n7559;
  assign n7561 = ~n7118 & ~n7560;
  assign n7562 = ~n7543 & n7561;
  assign n7563 = pi680 & ~n7366;
  assign n7564 = n2923 & n7563;
  assign n7565 = ~n7187 & n7564;
  assign n7566 = n7126 & n7563;
  assign n7567 = pi680 & n7544;
  assign n7568 = n6951 & n7563;
  assign n7569 = n7118 & n62828;
  assign n7570 = n7315 & n7564;
  assign n7571 = ~n7187 & n62827;
  assign n7572 = n7126 & n7408;
  assign n7573 = n7315 & n7565;
  assign n7574 = ~pi215 & ~n62829;
  assign n7575 = ~n7562 & n7574;
  assign n7576 = ~n7220 & ~n7366;
  assign n7577 = ~pi616 & ~n7576;
  assign n7578 = n7548 & ~n7577;
  assign n7579 = ~n7217 & n7551;
  assign n7580 = n7218 & n7551;
  assign n7581 = n7004 & n7579;
  assign n7582 = ~n7578 & ~n62830;
  assign n7583 = n62393 & ~n7582;
  assign n7584 = n7225 & n7551;
  assign n7585 = n7186 & n7217;
  assign n7586 = ~pi642 & ~n7579;
  assign n7587 = n2903 & n7586;
  assign n7588 = n7584 & ~n7587;
  assign n7589 = ~pi614 & n7586;
  assign n7590 = n7584 & ~n7589;
  assign n7591 = pi614 & ~pi616;
  assign n7592 = ~n7584 & n7591;
  assign n7593 = n7584 & ~n7586;
  assign n7594 = n2903 & ~n7593;
  assign n7595 = ~n7592 & ~n7594;
  assign n7596 = ~pi616 & ~n7590;
  assign n7597 = pi616 & ~n7584;
  assign n7598 = n62832 & ~n7597;
  assign n7599 = n7584 & ~n7585;
  assign n7600 = ~n7008 & ~n62831;
  assign n7601 = ~n6971 & n7408;
  assign n7602 = ~n7365 & ~n7601;
  assign n7603 = ~n7600 & ~n7602;
  assign n7604 = ~n62393 & n7603;
  assign n7605 = pi215 & ~n7604;
  assign n7606 = pi215 & ~n7583;
  assign n7607 = ~n7604 & n7606;
  assign n7608 = ~n7583 & n7605;
  assign n7609 = ~n7575 & ~n62833;
  assign n7610 = pi299 & ~n7609;
  assign n7611 = ~n2971 & n7542;
  assign n7612 = n2971 & ~n7559;
  assign n7613 = ~n7034 & ~n7612;
  assign n7614 = ~n7611 & n7613;
  assign n7615 = ~n7187 & ~n7563;
  assign n7616 = ~n7316 & ~n7565;
  assign n7617 = n6951 & ~n7616;
  assign n7618 = n6951 & ~n7615;
  assign n7619 = n7034 & ~n62834;
  assign n7620 = ~pi223 & ~n7619;
  assign n7621 = ~n62807 & n7620;
  assign n7622 = n7336 & ~n7619;
  assign n7623 = ~n7614 & n62835;
  assign n7624 = n2971 & n7582;
  assign n7625 = ~n2971 & ~n7603;
  assign n7626 = pi223 & ~n7625;
  assign n7627 = pi223 & ~n7624;
  assign n7628 = ~n7625 & n7627;
  assign n7629 = ~n7624 & n7626;
  assign n7630 = ~pi299 & ~n62836;
  assign n7631 = ~n7623 & n7630;
  assign n7632 = ~n7610 & ~n7631;
  assign n7633 = pi140 & n7632;
  assign n7634 = pi761 & ~n7633;
  assign n7635 = ~n7509 & n7634;
  assign n7636 = ~n7398 & ~n7532;
  assign n7637 = n7186 & ~n7636;
  assign n7638 = ~n7057 & n7187;
  assign n7639 = ~n7527 & ~n7638;
  assign n7640 = ~n7186 & ~n7639;
  assign n7641 = n7365 & ~n7640;
  assign n7642 = ~n7186 & n7639;
  assign n7643 = n7186 & ~n7532;
  assign n7644 = ~n7398 & n7643;
  assign n7645 = ~n7642 & ~n7644;
  assign n7646 = n7365 & ~n7645;
  assign n7647 = ~n7637 & n7641;
  assign n7648 = ~n7365 & ~n7539;
  assign n7649 = ~n7294 & n7648;
  assign n7650 = ~n62837 & ~n7649;
  assign n7651 = ~n62393 & ~n7650;
  assign n7652 = n7366 & ~n7399;
  assign n7653 = n6951 & ~n7652;
  assign n7654 = ~n7186 & n7653;
  assign n7655 = n7365 & ~n7654;
  assign n7656 = ~n7296 & ~n7552;
  assign n7657 = n7186 & ~n7656;
  assign n7658 = n7655 & ~n7657;
  assign n7659 = n7076 & n62822;
  assign n7660 = n2907 & ~n7659;
  assign n7661 = ~n7296 & n7660;
  assign n7662 = n7297 & ~n7659;
  assign n7663 = ~pi680 & ~n62803;
  assign n7664 = ~n62838 & ~n7663;
  assign n7665 = ~n7658 & n7664;
  assign n7666 = n62393 & ~n7665;
  assign n7667 = ~n7118 & ~n7666;
  assign n7668 = ~n62393 & n7650;
  assign n7669 = n62393 & n7665;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~n7118 & ~n7670;
  assign n7672 = ~n7651 & n7667;
  assign n7673 = n7126 & ~n7615;
  assign n7674 = n7118 & n62834;
  assign n7675 = ~pi215 & ~n62840;
  assign n7676 = ~n62839 & n7675;
  assign n7677 = ~n2904 & n7544;
  assign n7678 = ~n6978 & n7544;
  assign n7679 = ~n7677 & ~n7678;
  assign n7680 = ~n7322 & n7679;
  assign n7681 = n7186 & ~n7680;
  assign n7682 = n7655 & ~n7681;
  assign n7683 = n7008 & ~n7678;
  assign n7684 = pi680 & ~n7683;
  assign n7685 = n7327 & ~n7684;
  assign n7686 = ~n7682 & ~n7685;
  assign n7687 = n62393 & n7686;
  assign n7688 = ~n7326 & ~n7425;
  assign n7689 = ~n7679 & n7684;
  assign n7690 = ~n6973 & n7544;
  assign n7691 = n7689 & n7690;
  assign n7692 = n7688 & ~n7691;
  assign n7693 = ~n62393 & ~n7692;
  assign n7694 = pi215 & ~n7693;
  assign n7695 = ~n7687 & n7694;
  assign n7696 = ~n7676 & ~n7695;
  assign n7697 = pi299 & ~n7696;
  assign n7698 = ~n2971 & n7650;
  assign n7699 = n2971 & n7665;
  assign n7700 = ~n7034 & ~n7699;
  assign n7701 = ~n7698 & n7700;
  assign n7702 = n7620 & ~n7701;
  assign n7703 = n2971 & ~n7686;
  assign n7704 = ~n2971 & n7692;
  assign n7705 = pi223 & ~n7704;
  assign n7706 = ~n7703 & n7705;
  assign n7707 = ~pi299 & ~n7706;
  assign n7708 = ~n7702 & n7707;
  assign n7709 = ~n7697 & ~n7708;
  assign n7710 = pi140 & n7709;
  assign n7711 = n7191 & n7366;
  assign n7712 = n7381 & ~n7399;
  assign n7713 = ~n7186 & n7712;
  assign n7714 = n7365 & ~n7713;
  assign n7715 = ~n7711 & n7714;
  assign n7716 = ~pi680 & n7192;
  assign n7717 = n7385 & n7652;
  assign n7718 = n2907 & ~n7717;
  assign n7719 = ~n7716 & ~n7718;
  assign n7720 = ~n7715 & ~n7718;
  assign n7721 = ~n7716 & n7720;
  assign n7722 = ~n7715 & n7719;
  assign n7723 = n2971 & ~n62841;
  assign n7724 = ~n62786 & ~n7187;
  assign n7725 = ~pi680 & ~n7724;
  assign n7726 = ~n2952 & n7383;
  assign n7727 = ~n2904 & n7381;
  assign n7728 = ~n2814 & n7727;
  assign n7729 = ~n2904 & n7427;
  assign n7730 = n2952 & n7381;
  assign n7731 = ~n7726 & ~n62842;
  assign n7732 = n7652 & ~n7731;
  assign n7733 = n7365 & ~n7732;
  assign n7734 = ~n7401 & ~n7733;
  assign n7735 = ~n7725 & n7734;
  assign n7736 = ~n2971 & ~n7735;
  assign n7737 = ~n7034 & ~n7736;
  assign n7738 = ~n2971 & n7735;
  assign n7739 = n2971 & n62841;
  assign n7740 = ~n7723 & ~n7736;
  assign n7741 = ~n7738 & ~n7739;
  assign n7742 = ~n7034 & n62843;
  assign n7743 = ~n7723 & n7737;
  assign n7744 = n6955 & n7615;
  assign n7745 = ~n6948 & n7744;
  assign n7746 = n7034 & n7745;
  assign n7747 = ~pi223 & ~n7746;
  assign n7748 = ~n62844 & n7747;
  assign n7749 = ~n7220 & ~n7449;
  assign n7750 = n7365 & ~n7749;
  assign n7751 = ~pi680 & ~n7227;
  assign n7752 = pi680 & ~n7424;
  assign n7753 = ~n7399 & ~n7752;
  assign n7754 = n2907 & ~n7753;
  assign n7755 = ~n7751 & ~n7754;
  assign n7756 = ~n7750 & n7755;
  assign n7757 = ~n2971 & n7756;
  assign n7758 = n7221 & ~n7563;
  assign n7759 = n2907 & ~n7399;
  assign n7760 = n7431 & n7759;
  assign n7761 = ~n7758 & ~n7760;
  assign n7762 = n2971 & ~n7761;
  assign n7763 = pi223 & ~n7762;
  assign n7764 = pi223 & ~n7757;
  assign n7765 = ~n7762 & n7764;
  assign n7766 = ~n7757 & n7763;
  assign n7767 = ~n7034 & ~n62843;
  assign n7768 = n7034 & ~n7745;
  assign n7769 = ~pi223 & ~n7768;
  assign n7770 = ~n7767 & n7769;
  assign n7771 = ~n2971 & ~n7756;
  assign n7772 = n2971 & n7761;
  assign n7773 = pi223 & ~n7772;
  assign n7774 = ~n7771 & n7773;
  assign n7775 = ~n7770 & ~n7774;
  assign n7776 = ~n7748 & ~n62845;
  assign n7777 = ~pi299 & n62846;
  assign n7778 = n62393 & ~n62841;
  assign n7779 = ~n62393 & ~n7735;
  assign n7780 = ~n7118 & ~n7779;
  assign n7781 = ~n62393 & n7735;
  assign n7782 = n62393 & n62841;
  assign n7783 = ~n7778 & ~n7779;
  assign n7784 = ~n7781 & ~n7782;
  assign n7785 = ~n7118 & n62847;
  assign n7786 = ~n7778 & n7780;
  assign n7787 = n7118 & n7745;
  assign n7788 = ~pi215 & ~n7787;
  assign n7789 = ~n62848 & n7788;
  assign n7790 = ~n62393 & n7756;
  assign n7791 = n62393 & ~n7761;
  assign n7792 = pi215 & ~n7791;
  assign n7793 = pi215 & ~n7790;
  assign n7794 = ~n7791 & n7793;
  assign n7795 = ~n7790 & n7792;
  assign n7796 = ~n7118 & ~n62847;
  assign n7797 = n7118 & ~n7745;
  assign n7798 = ~pi215 & ~n7797;
  assign n7799 = ~n7796 & n7798;
  assign n7800 = ~n62393 & ~n7756;
  assign n7801 = n62393 & n7761;
  assign n7802 = pi215 & ~n7801;
  assign n7803 = ~n7800 & n7802;
  assign n7804 = ~n7799 & ~n7803;
  assign n7805 = ~n7789 & ~n62849;
  assign n7806 = pi299 & n62850;
  assign n7807 = ~pi299 & ~n62846;
  assign n7808 = pi299 & ~n62850;
  assign n7809 = ~n7807 & ~n7808;
  assign n7810 = ~n7777 & ~n7806;
  assign n7811 = ~pi140 & n62851;
  assign n7812 = ~pi761 & ~n7811;
  assign n7813 = ~n7710 & n7812;
  assign n7814 = ~n7635 & ~n7813;
  assign n7815 = pi39 & ~n7814;
  assign n7816 = pi665 & n6932;
  assign n7817 = pi198 & ~n7816;
  assign n7818 = pi665 & n6903;
  assign n7819 = ~pi198 & ~n7818;
  assign n7820 = ~n7817 & ~n7819;
  assign n7821 = pi680 & ~n7820;
  assign n7822 = n6940 & ~n7821;
  assign n7823 = ~pi299 & ~n7822;
  assign n7824 = ~pi210 & ~n7818;
  assign n7825 = pi210 & ~n7816;
  assign n7826 = ~n7824 & ~n7825;
  assign n7827 = pi680 & ~n7826;
  assign n7828 = n6936 & ~n7827;
  assign n7829 = pi299 & ~n7828;
  assign n7830 = ~n7823 & ~n7829;
  assign n7831 = pi680 & n7292;
  assign n7832 = ~n7830 & ~n7831;
  assign n7833 = ~pi140 & ~n7832;
  assign n7834 = pi665 & ~n6904;
  assign n7835 = ~n6905 & ~n7834;
  assign n7836 = ~pi198 & ~n7835;
  assign n7837 = pi665 & ~n6933;
  assign n7838 = ~n6934 & ~n7837;
  assign n7839 = pi198 & ~n7838;
  assign n7840 = ~n7836 & ~n7839;
  assign n7841 = ~pi603 & ~n7840;
  assign n7842 = pi603 & ~n7154;
  assign n7843 = ~n7549 & ~n7842;
  assign n7844 = ~n7841 & n7843;
  assign n7845 = pi680 & n7844;
  assign n7846 = ~pi299 & ~n7845;
  assign n7847 = pi210 & ~n7838;
  assign n7848 = ~pi210 & ~n7835;
  assign n7849 = ~n7847 & ~n7848;
  assign n7850 = ~pi603 & ~n7849;
  assign n7851 = ~n7168 & ~n7549;
  assign n7852 = ~n7850 & n7851;
  assign n7853 = pi680 & n7852;
  assign n7854 = pi299 & ~n7853;
  assign n7855 = ~n7846 & ~n7854;
  assign n7856 = pi140 & ~n7855;
  assign n7857 = pi761 & ~n7856;
  assign n7858 = pi761 & ~n7833;
  assign n7859 = ~n7856 & n7858;
  assign n7860 = ~n7833 & n7857;
  assign n7861 = n62793 & n7830;
  assign n7862 = ~pi140 & n7861;
  assign n7863 = pi680 & n7840;
  assign n7864 = ~pi299 & ~n7863;
  assign n7865 = pi680 & n7849;
  assign n7866 = pi299 & ~n7865;
  assign n7867 = ~n7864 & ~n7866;
  assign n7868 = ~n7292 & ~n7867;
  assign n7869 = pi140 & ~n7867;
  assign n7870 = ~n7292 & n7869;
  assign n7871 = pi140 & n7868;
  assign n7872 = ~pi761 & ~n62853;
  assign n7873 = ~n7862 & n7872;
  assign n7874 = ~pi39 & ~n7873;
  assign n7875 = pi140 & n7855;
  assign n7876 = ~pi140 & n7832;
  assign n7877 = pi761 & ~n7876;
  assign n7878 = ~n7875 & n7877;
  assign n7879 = ~pi140 & ~n7861;
  assign n7880 = pi140 & ~n7868;
  assign n7881 = ~pi761 & ~n7880;
  assign n7882 = ~n7862 & ~n62853;
  assign n7883 = ~pi761 & ~n7882;
  assign n7884 = ~n7879 & n7881;
  assign n7885 = ~n7878 & ~n62854;
  assign n7886 = ~pi39 & ~n7885;
  assign n7887 = ~n62852 & n7874;
  assign n7888 = ~pi38 & ~n62855;
  assign n7889 = ~n7815 & n7888;
  assign n7890 = pi761 & n7187;
  assign n7891 = n7357 & ~n7615;
  assign n7892 = n6955 & ~n7615;
  assign n7893 = ~pi39 & n7892;
  assign n7894 = n7356 & ~n7616;
  assign n7895 = ~n7890 & n62856;
  assign n7896 = ~n7358 & ~n7895;
  assign n7897 = ~pi761 & n7892;
  assign n7898 = ~pi140 & ~n6955;
  assign n7899 = n6955 & n7408;
  assign n7900 = n62380 & n7565;
  assign n7901 = pi761 & n62857;
  assign n7902 = ~pi39 & ~n7901;
  assign n7903 = ~n7898 & n7902;
  assign n7904 = ~pi140 & ~n7744;
  assign n7905 = pi140 & ~n7616;
  assign n7906 = n62380 & n7905;
  assign n7907 = ~pi761 & ~n7906;
  assign n7908 = ~n7904 & n7907;
  assign n7909 = pi761 & ~n62857;
  assign n7910 = pi761 & ~n7898;
  assign n7911 = ~n62857 & n7910;
  assign n7912 = ~n7898 & n7909;
  assign n7913 = ~n7908 & ~n62858;
  assign n7914 = ~pi39 & ~n7913;
  assign n7915 = ~n7897 & n7903;
  assign n7916 = pi39 & pi140;
  assign n7917 = pi38 & ~n7916;
  assign n7918 = ~n62859 & n7917;
  assign n7919 = pi38 & ~n7896;
  assign n7920 = ~n7889 & ~n62860;
  assign n7921 = ~pi738 & ~n7920;
  assign n7922 = n62765 & ~n7921;
  assign n7923 = n62765 & ~n7364;
  assign n7924 = ~n7921 & n7923;
  assign n7925 = ~n7364 & n7922;
  assign n7926 = ~n6800 & ~n62861;
  assign n7927 = ~pi778 & ~n7926;
  assign n7928 = pi625 & n7926;
  assign n7929 = n62765 & n7363;
  assign n7930 = ~n6800 & ~n7929;
  assign n7931 = ~pi625 & n7930;
  assign n7932 = pi1153 & ~n7931;
  assign n7933 = ~n7928 & n7932;
  assign n7934 = n2904 & n7385;
  assign n7935 = pi680 & ~n7727;
  assign n7936 = ~n7934 & n7935;
  assign n7937 = ~n7380 & ~n7936;
  assign n7938 = ~n7008 & n7937;
  assign n7939 = pi680 & ~n7385;
  assign n7940 = n7008 & ~n7939;
  assign n7941 = ~n7380 & n7940;
  assign n7942 = ~n7938 & ~n7941;
  assign n7943 = n62393 & n7942;
  assign n7944 = ~n7008 & ~n7731;
  assign n7945 = n7008 & n7383;
  assign n7946 = pi680 & ~n7945;
  assign n7947 = ~n7944 & n7946;
  assign n7948 = ~n7397 & ~n7947;
  assign n7949 = ~n62393 & ~n7948;
  assign n7950 = ~n7118 & ~n7949;
  assign n7951 = ~n7943 & n7950;
  assign n7952 = n2923 & ~n7563;
  assign n7953 = n7126 & ~n7563;
  assign n7954 = n7315 & n7952;
  assign n7955 = ~pi215 & ~n62862;
  assign n7956 = ~n7951 & n7955;
  assign n7957 = ~n7431 & n7935;
  assign n7958 = ~n7444 & ~n7957;
  assign n7959 = ~n7443 & ~n7957;
  assign n7960 = ~n7444 & n7959;
  assign n7961 = ~n7443 & n7958;
  assign n7962 = n62393 & n62863;
  assign n7963 = ~n62842 & n7752;
  assign n7964 = ~n7455 & ~n7963;
  assign n7965 = n7958 & n7964;
  assign n7966 = ~n62393 & n7965;
  assign n7967 = pi215 & ~n7966;
  assign n7968 = pi215 & ~n7962;
  assign n7969 = ~n7966 & n7968;
  assign n7970 = ~n7962 & n7967;
  assign n7971 = ~n7951 & ~n62862;
  assign n7972 = ~pi215 & ~n7971;
  assign n7973 = n62393 & ~n62863;
  assign n7974 = ~n62393 & ~n7965;
  assign n7975 = pi215 & ~n7974;
  assign n7976 = ~n7973 & n7975;
  assign n7977 = ~n7972 & ~n7976;
  assign n7978 = ~n7956 & ~n62864;
  assign n7979 = pi299 & ~n62865;
  assign n7980 = n2971 & n7942;
  assign n7981 = ~n2971 & ~n7948;
  assign n7982 = ~n7034 & ~n7981;
  assign n7983 = ~n7980 & n7982;
  assign n7984 = n62790 & ~n7563;
  assign n7985 = n7111 & n7952;
  assign n7986 = ~pi223 & ~n62866;
  assign n7987 = ~n7983 & n7986;
  assign n7988 = n2971 & n62863;
  assign n7989 = ~n2971 & n7965;
  assign n7990 = pi223 & ~n7989;
  assign n7991 = pi223 & ~n7988;
  assign n7992 = ~n7989 & n7991;
  assign n7993 = ~n7988 & n7990;
  assign n7994 = ~n7983 & ~n62866;
  assign n7995 = ~pi223 & ~n7994;
  assign n7996 = n2971 & ~n62863;
  assign n7997 = ~n2971 & ~n7965;
  assign n7998 = pi223 & ~n7997;
  assign n7999 = ~n7996 & n7998;
  assign n8000 = ~n7995 & ~n7999;
  assign n8001 = ~n7987 & ~n62867;
  assign n8002 = ~pi299 & ~n62868;
  assign n8003 = ~pi299 & n62868;
  assign n8004 = pi299 & n62865;
  assign n8005 = ~n8003 & ~n8004;
  assign n8006 = ~n7979 & ~n8002;
  assign n8007 = pi39 & n62869;
  assign n8008 = ~pi39 & n7830;
  assign n8009 = ~n8007 & ~n8008;
  assign n8010 = ~pi140 & n8009;
  assign n8011 = ~pi39 & n7867;
  assign n8012 = n62790 & n7563;
  assign n8013 = ~n62786 & n7563;
  assign n8014 = ~n7008 & n8013;
  assign n8015 = ~n7539 & ~n8014;
  assign n8016 = ~n2971 & n8015;
  assign n8017 = n2904 & n7659;
  assign n8018 = ~n7677 & ~n8017;
  assign n8019 = ~n7008 & n8018;
  assign n8020 = n7008 & ~n7659;
  assign n8021 = pi680 & ~n8020;
  assign n8022 = ~n8019 & n8021;
  assign n8023 = n2971 & ~n8022;
  assign n8024 = ~n7034 & ~n8023;
  assign n8025 = ~n7034 & ~n8016;
  assign n8026 = ~n8023 & n8025;
  assign n8027 = ~n8016 & n8024;
  assign n8028 = ~n8012 & ~n62870;
  assign n8029 = ~pi223 & ~n8028;
  assign n8030 = pi680 & ~n7679;
  assign n8031 = ~n7344 & n8030;
  assign n8032 = pi223 & ~n7683;
  assign n8033 = n8031 & n8032;
  assign n8034 = ~n8029 & ~n8033;
  assign n8035 = ~pi299 & ~n8034;
  assign n8036 = ~n62393 & ~n8015;
  assign n8037 = n62393 & n8022;
  assign n8038 = ~n7118 & ~n8037;
  assign n8039 = ~n8036 & n8038;
  assign n8040 = n7118 & ~n62828;
  assign n8041 = ~pi215 & ~n8040;
  assign n8042 = ~n62393 & n8015;
  assign n8043 = n62393 & ~n8022;
  assign n8044 = ~n7118 & ~n8043;
  assign n8045 = ~n7118 & ~n8042;
  assign n8046 = ~n8043 & n8045;
  assign n8047 = ~n8042 & n8044;
  assign n8048 = ~n62827 & ~n62871;
  assign n8049 = ~pi215 & ~n8048;
  assign n8050 = ~n8039 & n8041;
  assign n8051 = pi215 & ~n7328;
  assign n8052 = ~n7328 & n8030;
  assign n8053 = pi215 & ~n7683;
  assign n8054 = n8052 & n8053;
  assign n8055 = n7689 & n8051;
  assign n8056 = ~n62872 & ~n62873;
  assign n8057 = pi299 & ~n8056;
  assign n8058 = ~n8035 & ~n8057;
  assign n8059 = pi39 & ~n8058;
  assign n8060 = ~pi39 & ~n7867;
  assign n8061 = pi39 & n8058;
  assign n8062 = ~n8060 & ~n8061;
  assign n8063 = ~n8011 & ~n8059;
  assign n8064 = pi140 & n62874;
  assign n8065 = ~pi38 & ~n8064;
  assign n8066 = ~pi140 & ~n62869;
  assign n8067 = pi140 & ~n8058;
  assign n8068 = pi39 & ~n8067;
  assign n8069 = ~n7916 & ~n8007;
  assign n8070 = ~n8067 & ~n8069;
  assign n8071 = ~n8066 & n8068;
  assign n8072 = pi140 & n7867;
  assign n8073 = ~pi140 & ~n7830;
  assign n8074 = ~pi39 & ~n8073;
  assign n8075 = ~pi140 & n7830;
  assign n8076 = ~n7869 & ~n8075;
  assign n8077 = ~pi39 & ~n8076;
  assign n8078 = ~pi39 & ~n8072;
  assign n8079 = ~n8073 & n8078;
  assign n8080 = ~n8072 & n8074;
  assign n8081 = ~n62875 & ~n62876;
  assign n8082 = ~pi38 & ~n8081;
  assign n8083 = ~n8010 & n8065;
  assign n8084 = n7356 & n7564;
  assign n8085 = pi38 & ~n8084;
  assign n8086 = ~n7358 & n8085;
  assign n8087 = ~pi738 & ~n8086;
  assign n8088 = ~n62877 & n8087;
  assign n8089 = pi38 & ~n7357;
  assign n8090 = ~pi38 & ~n62792;
  assign n8091 = ~n8089 & ~n8090;
  assign n8092 = ~pi140 & pi738;
  assign n8093 = ~n8091 & n8092;
  assign n8094 = n62765 & ~n8093;
  assign n8095 = ~n8088 & n8094;
  assign n8096 = ~n6800 & ~n8095;
  assign n8097 = ~pi625 & n8096;
  assign n8098 = n62765 & n8091;
  assign n8099 = pi625 & ~n8098;
  assign n8100 = ~pi140 & ~n8098;
  assign n8101 = pi625 & n8100;
  assign n8102 = ~pi140 & n8099;
  assign n8103 = ~pi1153 & ~n62878;
  assign n8104 = ~n8097 & n8103;
  assign n8105 = pi608 & ~n8104;
  assign n8106 = ~n7933 & n8105;
  assign n8107 = ~pi625 & n7926;
  assign n8108 = pi625 & n7930;
  assign n8109 = ~pi1153 & ~n8108;
  assign n8110 = ~n8107 & n8109;
  assign n8111 = pi625 & n8096;
  assign n8112 = ~pi625 & n8100;
  assign n8113 = pi1153 & ~n8112;
  assign n8114 = ~n8111 & n8113;
  assign n8115 = ~pi608 & ~n8114;
  assign n8116 = ~n8110 & n8115;
  assign n8117 = pi778 & ~n8116;
  assign n8118 = ~n8106 & n8117;
  assign n8119 = ~n8106 & ~n8116;
  assign n8120 = pi778 & ~n8119;
  assign n8121 = ~pi778 & n7926;
  assign n8122 = ~n8120 & ~n8121;
  assign n8123 = ~n7927 & ~n8118;
  assign n8124 = ~pi609 & ~n62879;
  assign n8125 = ~pi778 & ~n8096;
  assign n8126 = ~n8104 & ~n8114;
  assign n8127 = pi778 & ~n8126;
  assign n8128 = ~n8125 & ~n8127;
  assign n8129 = pi609 & n8128;
  assign n8130 = ~pi1155 & ~n8129;
  assign n8131 = ~n8124 & n8130;
  assign n8132 = pi608 & ~pi1153;
  assign n8133 = ~pi608 & pi1153;
  assign n8134 = ~n8132 & ~n8133;
  assign n8135 = pi778 & ~n8134;
  assign n8136 = pi609 & ~n8135;
  assign n8137 = ~n8100 & ~n8136;
  assign n8138 = ~n7930 & ~n8135;
  assign n8139 = pi609 & n8138;
  assign n8140 = ~n8137 & ~n8139;
  assign n8141 = pi1155 & ~n8140;
  assign n8142 = ~pi660 & ~n8141;
  assign n8143 = ~n8131 & n8142;
  assign n8144 = pi609 & ~n62879;
  assign n8145 = ~pi609 & n8128;
  assign n8146 = pi1155 & ~n8145;
  assign n8147 = ~n8144 & n8146;
  assign n8148 = ~pi609 & ~n8135;
  assign n8149 = ~n8100 & ~n8148;
  assign n8150 = ~pi609 & n8138;
  assign n8151 = ~n8149 & ~n8150;
  assign n8152 = ~pi1155 & ~n8151;
  assign n8153 = pi660 & ~n8152;
  assign n8154 = ~n8147 & n8153;
  assign n8155 = ~n8143 & ~n8154;
  assign n8156 = pi785 & ~n8155;
  assign n8157 = ~pi785 & ~n62879;
  assign n8158 = ~n8156 & ~n8157;
  assign n8159 = ~pi618 & ~n8158;
  assign n8160 = pi660 & ~pi1155;
  assign n8161 = ~pi660 & pi1155;
  assign n8162 = ~n8160 & ~n8161;
  assign n8163 = ~pi660 & ~pi1155;
  assign n8164 = pi660 & pi1155;
  assign n8165 = pi785 & ~n8164;
  assign n8166 = ~n8163 & n8165;
  assign n8167 = pi785 & ~n8163;
  assign n8168 = ~n8164 & n8167;
  assign n8169 = pi785 & ~n8162;
  assign n8170 = ~n8128 & ~n62880;
  assign n8171 = ~n8100 & n62880;
  assign n8172 = n8128 & ~n62880;
  assign n8173 = n8100 & n62880;
  assign n8174 = ~n8172 & ~n8173;
  assign n8175 = ~n8170 & ~n8171;
  assign n8176 = pi618 & ~n62881;
  assign n8177 = ~pi1154 & ~n8176;
  assign n8178 = ~n8159 & n8177;
  assign n8179 = ~n8100 & n8135;
  assign n8180 = ~n8138 & ~n8179;
  assign n8181 = ~pi785 & ~n8180;
  assign n8182 = ~n8141 & ~n8152;
  assign n8183 = pi785 & ~n8182;
  assign n8184 = ~n8181 & ~n8183;
  assign n8185 = pi618 & n8184;
  assign n8186 = ~pi618 & n8100;
  assign n8187 = pi1154 & ~n8186;
  assign n8188 = ~n8185 & n8187;
  assign n8189 = ~pi627 & ~n8188;
  assign n8190 = ~n8178 & n8189;
  assign n8191 = pi618 & ~n8158;
  assign n8192 = ~pi618 & ~n62881;
  assign n8193 = pi1154 & ~n8192;
  assign n8194 = ~n8191 & n8193;
  assign n8195 = ~pi618 & n8184;
  assign n8196 = pi618 & n8100;
  assign n8197 = ~pi1154 & ~n8196;
  assign n8198 = ~n8195 & n8197;
  assign n8199 = pi627 & ~n8198;
  assign n8200 = ~n8194 & n8199;
  assign n8201 = ~n8190 & ~n8200;
  assign n8202 = pi781 & ~n8201;
  assign n8203 = ~pi781 & ~n8158;
  assign n8204 = ~n8202 & ~n8203;
  assign n8205 = ~pi619 & ~n8204;
  assign n8206 = pi627 & ~pi1154;
  assign n8207 = ~pi627 & pi1154;
  assign n8208 = ~n8206 & ~n8207;
  assign n8209 = ~pi627 & ~pi1154;
  assign n8210 = pi627 & pi1154;
  assign n8211 = pi781 & ~n8210;
  assign n8212 = ~n8209 & n8211;
  assign n8213 = pi781 & ~n8209;
  assign n8214 = ~n8210 & n8213;
  assign n8215 = pi781 & ~n8208;
  assign n8216 = ~n62881 & ~n62882;
  assign n8217 = n8100 & n62882;
  assign n8218 = n62881 & ~n62882;
  assign n8219 = ~n8100 & n62882;
  assign n8220 = ~n8218 & ~n8219;
  assign n8221 = ~n8216 & ~n8217;
  assign n8222 = pi619 & n62883;
  assign n8223 = ~pi1159 & ~n8222;
  assign n8224 = ~n8205 & n8223;
  assign n8225 = ~pi781 & ~n8184;
  assign n8226 = ~n8188 & ~n8198;
  assign n8227 = pi781 & ~n8226;
  assign n8228 = ~n8225 & ~n8227;
  assign n8229 = pi619 & n8228;
  assign n8230 = ~pi619 & n8100;
  assign n8231 = pi1159 & ~n8230;
  assign n8232 = ~n8229 & n8231;
  assign n8233 = ~pi648 & ~n8232;
  assign n8234 = ~n8224 & n8233;
  assign n8235 = pi619 & ~n8204;
  assign n8236 = ~pi619 & n62883;
  assign n8237 = pi1159 & ~n8236;
  assign n8238 = ~n8235 & n8237;
  assign n8239 = ~pi619 & n8228;
  assign n8240 = pi619 & n8100;
  assign n8241 = ~pi1159 & ~n8240;
  assign n8242 = ~n8239 & n8241;
  assign n8243 = pi648 & ~n8242;
  assign n8244 = ~n8238 & n8243;
  assign n8245 = ~n8234 & ~n8244;
  assign n8246 = pi789 & ~n8245;
  assign n8247 = ~pi789 & ~n8204;
  assign n8248 = ~n8246 & ~n8247;
  assign n8249 = ~pi788 & n8248;
  assign n8250 = ~pi626 & n8248;
  assign n8251 = ~pi648 & ~pi1159;
  assign n8252 = pi648 & pi1159;
  assign n8253 = ~pi648 & pi1159;
  assign n8254 = pi648 & ~pi1159;
  assign n8255 = ~n8253 & ~n8254;
  assign n8256 = ~n8251 & ~n8252;
  assign n8257 = pi789 & ~n62884;
  assign n8258 = ~n62883 & ~n8257;
  assign n8259 = ~n8100 & n8257;
  assign n8260 = n62883 & ~n8257;
  assign n8261 = n8100 & n8257;
  assign n8262 = ~n8260 & ~n8261;
  assign n8263 = ~n8258 & ~n8259;
  assign n8264 = pi626 & n62885;
  assign n8265 = ~pi641 & ~n8264;
  assign n8266 = ~n8250 & n8265;
  assign n8267 = ~pi641 & ~pi1158;
  assign n8268 = ~pi789 & ~n8228;
  assign n8269 = ~n8232 & ~n8242;
  assign n8270 = pi789 & ~n8269;
  assign n8271 = ~n8268 & ~n8270;
  assign n8272 = ~pi626 & n8271;
  assign n8273 = pi626 & n8100;
  assign n8274 = ~pi1158 & ~n8273;
  assign n8275 = ~n8272 & n8274;
  assign n8276 = ~n8267 & ~n8275;
  assign n8277 = ~n8266 & ~n8276;
  assign n8278 = pi626 & n8248;
  assign n8279 = ~pi626 & n62885;
  assign n8280 = pi641 & ~n8279;
  assign n8281 = ~n8278 & n8280;
  assign n8282 = pi641 & pi1158;
  assign n8283 = pi626 & n8271;
  assign n8284 = ~pi626 & n8100;
  assign n8285 = pi1158 & ~n8284;
  assign n8286 = ~n8283 & n8285;
  assign n8287 = ~n8282 & ~n8286;
  assign n8288 = ~n8281 & ~n8287;
  assign n8289 = ~n8277 & ~n8288;
  assign n8290 = pi788 & ~n8289;
  assign n8291 = ~n8249 & ~n8290;
  assign n8292 = ~pi628 & n8291;
  assign n8293 = ~n8275 & ~n8286;
  assign n8294 = pi788 & ~n8293;
  assign n8295 = ~pi788 & ~n8271;
  assign n8296 = ~n8294 & ~n8295;
  assign n8297 = pi628 & n8296;
  assign n8298 = ~pi1156 & ~n8297;
  assign n8299 = ~n8292 & n8298;
  assign n8300 = ~pi641 & pi1158;
  assign n8301 = pi641 & ~pi1158;
  assign n8302 = ~n8300 & ~n8301;
  assign n8303 = pi788 & ~n8302;
  assign n8304 = ~n62885 & ~n8303;
  assign n8305 = n8100 & n8303;
  assign n8306 = n62885 & ~n8303;
  assign n8307 = ~n8100 & n8303;
  assign n8308 = ~n8306 & ~n8307;
  assign n8309 = ~n8304 & ~n8305;
  assign n8310 = pi628 & n62886;
  assign n8311 = ~pi628 & n8100;
  assign n8312 = pi1156 & ~n8311;
  assign n8313 = ~n8310 & n8312;
  assign n8314 = ~pi629 & ~n8313;
  assign n8315 = ~n8299 & n8314;
  assign n8316 = pi628 & n8291;
  assign n8317 = ~pi628 & n8296;
  assign n8318 = pi1156 & ~n8317;
  assign n8319 = ~n8316 & n8318;
  assign n8320 = ~pi628 & n62886;
  assign n8321 = pi628 & n8100;
  assign n8322 = ~pi1156 & ~n8321;
  assign n8323 = ~n8320 & n8322;
  assign n8324 = pi629 & ~n8323;
  assign n8325 = ~n8319 & n8324;
  assign n8326 = ~n8315 & ~n8325;
  assign n8327 = pi792 & ~n8326;
  assign n8328 = ~pi792 & n8291;
  assign n8329 = ~n8327 & ~n8328;
  assign n8330 = ~pi647 & ~n8329;
  assign n8331 = ~pi629 & pi1156;
  assign n8332 = pi629 & ~pi1156;
  assign n8333 = ~n8331 & ~n8332;
  assign n8334 = pi792 & ~n8333;
  assign n8335 = n8296 & ~n8334;
  assign n8336 = n8100 & n8334;
  assign n8337 = ~n8335 & ~n8336;
  assign n8338 = pi647 & ~n8337;
  assign n8339 = ~pi1157 & ~n8338;
  assign n8340 = ~n8330 & n8339;
  assign n8341 = ~pi792 & ~n62886;
  assign n8342 = ~n8313 & ~n8323;
  assign n8343 = pi792 & ~n8342;
  assign n8344 = ~n8341 & ~n8343;
  assign n8345 = pi647 & n8344;
  assign n8346 = ~pi647 & n8100;
  assign n8347 = pi1157 & ~n8346;
  assign n8348 = ~n8345 & n8347;
  assign n8349 = ~pi630 & ~n8348;
  assign n8350 = ~n8340 & n8349;
  assign n8351 = pi647 & ~n8329;
  assign n8352 = ~pi647 & ~n8337;
  assign n8353 = pi1157 & ~n8352;
  assign n8354 = ~n8351 & n8353;
  assign n8355 = ~pi647 & n8344;
  assign n8356 = pi647 & n8100;
  assign n8357 = ~pi1157 & ~n8356;
  assign n8358 = ~n8355 & n8357;
  assign n8359 = pi630 & ~n8358;
  assign n8360 = ~n8354 & n8359;
  assign n8361 = ~n8350 & ~n8360;
  assign n8362 = pi787 & ~n8361;
  assign n8363 = ~pi787 & ~n8329;
  assign n8364 = ~n8362 & ~n8363;
  assign n8365 = ~pi644 & ~n8364;
  assign n8366 = ~pi787 & ~n8344;
  assign n8367 = ~n8348 & ~n8358;
  assign n8368 = pi787 & ~n8367;
  assign n8369 = ~n8366 & ~n8368;
  assign n8370 = pi644 & n8369;
  assign n8371 = ~pi715 & ~n8370;
  assign n8372 = ~n8365 & n8371;
  assign n8373 = ~pi630 & pi1157;
  assign n8374 = pi630 & ~pi1157;
  assign n8375 = ~n8373 & ~n8374;
  assign n8376 = pi787 & ~n8375;
  assign n8377 = n8337 & ~n8376;
  assign n8378 = ~n8100 & n8376;
  assign n8379 = ~n8337 & ~n8376;
  assign n8380 = n8100 & n8376;
  assign n8381 = ~n8379 & ~n8380;
  assign n8382 = ~n8377 & ~n8378;
  assign n8383 = ~pi644 & ~n62887;
  assign n8384 = pi644 & n8100;
  assign n8385 = pi715 & ~n8384;
  assign n8386 = ~n8383 & n8385;
  assign n8387 = ~pi1160 & ~n8386;
  assign n8388 = ~n8372 & n8387;
  assign n8389 = pi644 & ~n8364;
  assign n8390 = ~pi644 & n8369;
  assign n8391 = pi715 & ~n8390;
  assign n8392 = ~n8389 & n8391;
  assign n8393 = pi644 & ~n62887;
  assign n8394 = ~pi644 & n8100;
  assign n8395 = ~pi715 & ~n8394;
  assign n8396 = ~n8393 & n8395;
  assign n8397 = pi1160 & ~n8396;
  assign n8398 = ~n8392 & n8397;
  assign n8399 = pi790 & ~n8398;
  assign n8400 = pi790 & ~n8388;
  assign n8401 = ~n8398 & n8400;
  assign n8402 = ~n8388 & n8399;
  assign n8403 = ~pi790 & n8364;
  assign n8404 = n62455 & ~n8403;
  assign n8405 = ~n62888 & n8404;
  assign n8406 = ~pi140 & ~n62455;
  assign n8407 = ~pi832 & ~n8406;
  assign n8408 = ~n8405 & n8407;
  assign n8409 = pi630 & ~pi647;
  assign n8410 = pi1157 & n8409;
  assign n8411 = ~pi630 & pi647;
  assign n8412 = ~pi1157 & n8411;
  assign n8413 = ~n8410 & ~n8412;
  assign n8414 = ~pi140 & ~n2923;
  assign n8415 = n8334 & ~n8414;
  assign n8416 = ~pi626 & pi1158;
  assign n8417 = pi626 & ~pi1158;
  assign n8418 = ~n8416 & ~n8417;
  assign n8419 = n8414 & ~n8418;
  assign n8420 = n2923 & n8135;
  assign n8421 = ~pi761 & n7316;
  assign n8422 = ~n8414 & ~n8421;
  assign n8423 = ~n8420 & ~n8422;
  assign n8424 = ~pi785 & ~n8423;
  assign n8425 = n2923 & ~n8136;
  assign n8426 = ~n8422 & ~n8425;
  assign n8427 = pi1155 & ~n8426;
  assign n8428 = pi609 & n2923;
  assign n8429 = n8423 & ~n8428;
  assign n8430 = ~pi1155 & ~n8429;
  assign n8431 = ~n8427 & ~n8430;
  assign n8432 = pi785 & ~n8431;
  assign n8433 = ~n8424 & ~n8432;
  assign n8434 = ~pi781 & ~n8433;
  assign n8435 = ~pi618 & n2923;
  assign n8436 = n8433 & ~n8435;
  assign n8437 = pi1154 & ~n8436;
  assign n8438 = pi618 & n2923;
  assign n8439 = n8433 & ~n8438;
  assign n8440 = ~pi1154 & ~n8439;
  assign n8441 = ~n8437 & ~n8440;
  assign n8442 = pi781 & ~n8441;
  assign n8443 = ~n8434 & ~n8442;
  assign n8444 = ~pi789 & ~n8443;
  assign n8445 = pi619 & n8443;
  assign n8446 = ~pi619 & n8414;
  assign n8447 = pi1159 & ~n8446;
  assign n8448 = ~n8445 & n8447;
  assign n8449 = ~pi619 & n8443;
  assign n8450 = pi619 & n8414;
  assign n8451 = ~pi1159 & ~n8450;
  assign n8452 = ~n8449 & n8451;
  assign n8453 = ~n8448 & ~n8452;
  assign n8454 = pi789 & ~n8453;
  assign n8455 = ~n8444 & ~n8454;
  assign n8456 = n8418 & n8455;
  assign n8457 = pi626 & n8455;
  assign n8458 = ~pi626 & n8414;
  assign n8459 = pi1158 & ~n8458;
  assign n8460 = ~n8457 & n8459;
  assign n8461 = ~pi626 & n8455;
  assign n8462 = pi626 & n8414;
  assign n8463 = ~pi1158 & ~n8462;
  assign n8464 = ~n8461 & n8463;
  assign n8465 = ~n8460 & ~n8464;
  assign n8466 = ~n8419 & ~n8456;
  assign n8467 = pi788 & n62889;
  assign n8468 = ~pi788 & n8455;
  assign n8469 = ~pi788 & ~n8455;
  assign n8470 = pi788 & ~n62889;
  assign n8471 = ~n8469 & ~n8470;
  assign n8472 = ~n8467 & ~n8468;
  assign n8473 = ~n8334 & ~n62890;
  assign n8474 = ~n8334 & n62890;
  assign n8475 = n8334 & n8414;
  assign n8476 = ~n8474 & ~n8475;
  assign n8477 = ~n8415 & ~n8473;
  assign n8478 = ~n8413 & n62891;
  assign n8479 = ~pi738 & n7564;
  assign n8480 = ~n8414 & ~n8479;
  assign n8481 = ~pi778 & n8480;
  assign n8482 = ~pi625 & n8479;
  assign n8483 = ~n8480 & ~n8482;
  assign n8484 = pi1153 & ~n8483;
  assign n8485 = ~pi1153 & ~n8414;
  assign n8486 = ~n8482 & n8485;
  assign n8487 = ~n8484 & ~n8486;
  assign n8488 = pi778 & ~n8487;
  assign n8489 = ~n8481 & ~n8488;
  assign n8490 = n2923 & n62880;
  assign n8491 = n8489 & ~n8490;
  assign n8492 = n2923 & n62882;
  assign n8493 = n8491 & ~n8492;
  assign n8494 = n2923 & n8257;
  assign n8495 = n8493 & ~n8494;
  assign n8496 = n2923 & n8303;
  assign n8497 = n8495 & ~n8496;
  assign n8498 = ~pi628 & pi1156;
  assign n8499 = pi628 & ~pi1156;
  assign n8500 = ~n8498 & ~n8499;
  assign n8501 = ~pi628 & ~pi1156;
  assign n8502 = pi628 & pi1156;
  assign n8503 = pi792 & ~n8502;
  assign n8504 = ~n8501 & n8503;
  assign n8505 = pi792 & ~n8501;
  assign n8506 = ~n8502 & n8505;
  assign n8507 = pi792 & ~n8500;
  assign n8508 = n2923 & n62892;
  assign n8509 = n8497 & ~n8508;
  assign n8510 = pi647 & ~n8509;
  assign n8511 = ~pi647 & ~n8414;
  assign n8512 = ~n8510 & ~n8511;
  assign n8513 = n8373 & ~n8512;
  assign n8514 = ~pi647 & n8509;
  assign n8515 = pi647 & n8414;
  assign n8516 = ~pi1157 & ~n8515;
  assign n8517 = ~n8514 & n8516;
  assign n8518 = pi630 & n8517;
  assign n8519 = ~n8513 & ~n8518;
  assign n8520 = ~n8478 & n8519;
  assign n8521 = pi787 & ~n8520;
  assign n8522 = ~pi626 & pi641;
  assign n8523 = pi626 & ~pi641;
  assign n8524 = ~n8522 & ~n8523;
  assign n8525 = ~n8418 & ~n8524;
  assign n8526 = n8495 & n8525;
  assign n8527 = ~n8302 & n62889;
  assign n8528 = ~n8526 & ~n8527;
  assign n8529 = pi788 & ~n8528;
  assign n8530 = ~n7187 & ~n8480;
  assign n8531 = pi625 & n8530;
  assign n8532 = n8422 & ~n8530;
  assign n8533 = ~n8531 & ~n8532;
  assign n8534 = n8485 & ~n8533;
  assign n8535 = ~pi608 & ~n8484;
  assign n8536 = ~n8534 & n8535;
  assign n8537 = pi1153 & n8422;
  assign n8538 = ~n8531 & n8537;
  assign n8539 = pi608 & ~n8486;
  assign n8540 = ~n8538 & n8539;
  assign n8541 = ~n8536 & ~n8540;
  assign n8542 = pi778 & ~n8541;
  assign n8543 = ~pi778 & ~n8532;
  assign n8544 = ~n8542 & ~n8543;
  assign n8545 = ~pi609 & ~n8544;
  assign n8546 = pi609 & n8489;
  assign n8547 = ~pi1155 & ~n8546;
  assign n8548 = ~n8545 & n8547;
  assign n8549 = ~pi660 & ~n8427;
  assign n8550 = ~n8548 & n8549;
  assign n8551 = pi609 & ~n8544;
  assign n8552 = ~pi609 & n8489;
  assign n8553 = pi1155 & ~n8552;
  assign n8554 = ~n8551 & n8553;
  assign n8555 = pi660 & ~n8430;
  assign n8556 = ~n8554 & n8555;
  assign n8557 = ~n8550 & ~n8556;
  assign n8558 = pi785 & ~n8557;
  assign n8559 = ~pi785 & ~n8544;
  assign n8560 = ~n8558 & ~n8559;
  assign n8561 = ~pi618 & ~n8560;
  assign n8562 = pi618 & n8491;
  assign n8563 = ~pi1154 & ~n8562;
  assign n8564 = ~n8561 & n8563;
  assign n8565 = ~pi627 & ~n8437;
  assign n8566 = ~n8564 & n8565;
  assign n8567 = pi618 & ~n8560;
  assign n8568 = ~pi618 & n8491;
  assign n8569 = pi1154 & ~n8568;
  assign n8570 = ~n8567 & n8569;
  assign n8571 = pi627 & ~n8440;
  assign n8572 = ~n8570 & n8571;
  assign n8573 = ~n8566 & ~n8572;
  assign n8574 = pi781 & ~n8573;
  assign n8575 = ~pi781 & ~n8560;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = pi619 & ~n8576;
  assign n8578 = ~pi619 & n8493;
  assign n8579 = pi1159 & ~n8578;
  assign n8580 = ~n8577 & n8579;
  assign n8581 = pi648 & ~n8452;
  assign n8582 = ~n8580 & n8581;
  assign n8583 = ~pi619 & ~n8576;
  assign n8584 = pi619 & n8493;
  assign n8585 = ~pi1159 & ~n8584;
  assign n8586 = ~n8583 & n8585;
  assign n8587 = ~pi648 & ~n8448;
  assign n8588 = ~n8586 & n8587;
  assign n8589 = pi789 & ~n8588;
  assign n8590 = pi789 & ~n8582;
  assign n8591 = ~n8588 & n8590;
  assign n8592 = ~n8582 & n8589;
  assign n8593 = ~pi789 & n8576;
  assign n8594 = n8418 & n8524;
  assign n8595 = pi788 & ~n8418;
  assign n8596 = ~n8303 & ~n8595;
  assign n8597 = pi788 & ~n8594;
  assign n8598 = ~n8593 & n62894;
  assign n8599 = ~n62893 & n8598;
  assign n8600 = ~n8529 & ~n8599;
  assign n8601 = ~pi628 & n8600;
  assign n8602 = pi628 & ~n62890;
  assign n8603 = ~pi1156 & ~n8602;
  assign n8604 = ~n8601 & n8603;
  assign n8605 = ~pi628 & n2923;
  assign n8606 = pi1156 & ~n8605;
  assign n8607 = n8497 & n8606;
  assign n8608 = ~pi629 & ~n8607;
  assign n8609 = ~n8604 & n8608;
  assign n8610 = pi628 & n8600;
  assign n8611 = ~pi628 & ~n62890;
  assign n8612 = pi1156 & ~n8611;
  assign n8613 = ~n8610 & n8612;
  assign n8614 = pi628 & n2923;
  assign n8615 = ~pi1156 & ~n8614;
  assign n8616 = n8497 & n8615;
  assign n8617 = pi629 & ~n8616;
  assign n8618 = ~n8613 & n8617;
  assign n8619 = pi792 & ~n8618;
  assign n8620 = pi792 & ~n8609;
  assign n8621 = ~n8618 & n8620;
  assign n8622 = ~pi628 & ~n8600;
  assign n8623 = pi628 & n62890;
  assign n8624 = ~pi1156 & ~n8623;
  assign n8625 = ~n8622 & n8624;
  assign n8626 = n8497 & ~n8605;
  assign n8627 = pi1156 & ~n8626;
  assign n8628 = ~pi629 & ~n8627;
  assign n8629 = ~n8625 & n8628;
  assign n8630 = pi628 & ~n8600;
  assign n8631 = ~pi628 & n62890;
  assign n8632 = pi1156 & ~n8631;
  assign n8633 = ~n8630 & n8632;
  assign n8634 = n8497 & ~n8614;
  assign n8635 = ~pi1156 & ~n8634;
  assign n8636 = pi629 & ~n8635;
  assign n8637 = ~n8633 & n8636;
  assign n8638 = ~n8629 & ~n8637;
  assign n8639 = pi792 & ~n8638;
  assign n8640 = ~n8609 & n8619;
  assign n8641 = ~pi792 & ~n8600;
  assign n8642 = ~pi647 & pi1157;
  assign n8643 = pi647 & ~pi1157;
  assign n8644 = ~n8642 & ~n8643;
  assign n8645 = ~pi630 & ~pi647;
  assign n8646 = ~pi1157 & n8645;
  assign n8647 = pi630 & pi647;
  assign n8648 = pi1157 & n8647;
  assign n8649 = ~n8646 & ~n8648;
  assign n8650 = n8375 & n8644;
  assign n8651 = pi787 & n62896;
  assign n8652 = ~n8641 & ~n8651;
  assign n8653 = ~n62895 & n8652;
  assign n8654 = ~n62895 & ~n8641;
  assign n8655 = ~pi647 & ~n8654;
  assign n8656 = pi647 & ~n62891;
  assign n8657 = ~pi1157 & ~n8656;
  assign n8658 = ~n8655 & n8657;
  assign n8659 = pi647 & n8509;
  assign n8660 = ~pi647 & n8414;
  assign n8661 = pi1157 & ~n8660;
  assign n8662 = pi1157 & ~n8512;
  assign n8663 = ~n8659 & n8661;
  assign n8664 = ~pi630 & ~n62897;
  assign n8665 = ~n8658 & n8664;
  assign n8666 = pi647 & ~n8654;
  assign n8667 = ~pi647 & ~n62891;
  assign n8668 = pi1157 & ~n8667;
  assign n8669 = ~n8666 & n8668;
  assign n8670 = pi630 & ~n8517;
  assign n8671 = ~n8669 & n8670;
  assign n8672 = ~n8665 & ~n8671;
  assign n8673 = pi787 & ~n8672;
  assign n8674 = ~pi787 & ~n8654;
  assign n8675 = ~n8673 & ~n8674;
  assign n8676 = ~n8521 & ~n8653;
  assign n8677 = pi644 & ~n62898;
  assign n8678 = ~pi787 & ~n8509;
  assign n8679 = ~n8517 & ~n62897;
  assign n8680 = pi787 & ~n8679;
  assign n8681 = ~n8678 & ~n8680;
  assign n8682 = ~pi644 & n8681;
  assign n8683 = pi715 & ~n8682;
  assign n8684 = ~n8677 & n8683;
  assign n8685 = ~n8334 & ~n8376;
  assign n8686 = ~n8414 & ~n8685;
  assign n8687 = ~n8376 & n8473;
  assign n8688 = n8376 & ~n8414;
  assign n8689 = ~n8376 & n62891;
  assign n8690 = ~n8688 & ~n8689;
  assign n8691 = ~n8686 & ~n8687;
  assign n8692 = pi644 & n62899;
  assign n8693 = ~pi644 & n8414;
  assign n8694 = ~pi715 & ~n8693;
  assign n8695 = ~n8692 & n8694;
  assign n8696 = pi1160 & ~n8695;
  assign n8697 = ~n8684 & n8696;
  assign n8698 = ~pi644 & ~n62898;
  assign n8699 = pi644 & n8681;
  assign n8700 = ~pi715 & ~n8699;
  assign n8701 = ~n8698 & n8700;
  assign n8702 = ~pi644 & n62899;
  assign n8703 = pi644 & n8414;
  assign n8704 = pi715 & ~n8703;
  assign n8705 = ~n8702 & n8704;
  assign n8706 = ~pi1160 & ~n8705;
  assign n8707 = ~n8701 & n8706;
  assign n8708 = ~n8697 & ~n8707;
  assign n8709 = pi790 & ~n8708;
  assign n8710 = ~pi790 & ~n62898;
  assign n8711 = pi832 & ~n8710;
  assign n8712 = ~n8709 & n8711;
  assign po297 = ~n8408 & ~n8712;
  assign n8714 = pi141 & ~n62765;
  assign n8715 = ~pi141 & ~n7357;
  assign n8716 = pi749 & n7359;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = pi38 & ~n8717;
  assign n8719 = ~pi749 & n7143;
  assign n8720 = pi141 & n7349;
  assign n8721 = ~n8719 & ~n8720;
  assign n8722 = pi39 & ~n8721;
  assign n8723 = ~pi141 & n62802;
  assign n8724 = pi141 & n7293;
  assign n8725 = pi749 & ~n8724;
  assign n8726 = ~n8723 & n8725;
  assign n8727 = ~pi141 & ~pi749;
  assign n8728 = ~n6946 & n8727;
  assign n8729 = ~n8726 & ~n8728;
  assign n8730 = ~pi38 & ~n8729;
  assign n8731 = ~n8722 & n8730;
  assign n8732 = ~n8718 & ~n8731;
  assign n8733 = ~pi706 & ~n8732;
  assign n8734 = ~pi141 & ~n62821;
  assign n8735 = pi141 & n7632;
  assign n8736 = ~pi749 & ~n8735;
  assign n8737 = ~n8734 & n8736;
  assign n8738 = pi141 & n7709;
  assign n8739 = ~pi141 & n62851;
  assign n8740 = pi749 & ~n8739;
  assign n8741 = ~n8738 & n8740;
  assign n8742 = pi39 & ~n8741;
  assign n8743 = ~n8737 & n8742;
  assign n8744 = ~pi141 & n7832;
  assign n8745 = pi141 & n7855;
  assign n8746 = ~pi749 & ~n8745;
  assign n8747 = ~pi749 & ~n8744;
  assign n8748 = ~n8745 & n8747;
  assign n8749 = ~n8744 & n8746;
  assign n8750 = ~pi141 & ~n7861;
  assign n8751 = pi141 & ~n7868;
  assign n8752 = pi749 & ~n8751;
  assign n8753 = ~n8750 & n8752;
  assign n8754 = ~pi39 & ~n8753;
  assign n8755 = ~n62900 & n8754;
  assign n8756 = ~pi38 & ~n8755;
  assign n8757 = ~pi39 & ~n7832;
  assign n8758 = pi39 & n62821;
  assign n8759 = ~n8757 & ~n8758;
  assign n8760 = ~pi141 & n8759;
  assign n8761 = pi39 & ~n7632;
  assign n8762 = ~pi39 & ~n7855;
  assign n8763 = ~n8761 & ~n8762;
  assign n8764 = pi141 & n8763;
  assign n8765 = ~pi749 & ~n8764;
  assign n8766 = ~n8760 & n8765;
  assign n8767 = pi39 & ~n8739;
  assign n8768 = ~n8738 & n8767;
  assign n8769 = ~pi39 & ~n8751;
  assign n8770 = ~n8750 & n8769;
  assign n8771 = ~n8768 & ~n8770;
  assign n8772 = pi39 & ~n7709;
  assign n8773 = ~n7292 & n8060;
  assign n8774 = n7293 & ~n7867;
  assign n8775 = ~n8772 & ~n62901;
  assign n8776 = pi141 & n8775;
  assign n8777 = pi39 & n62851;
  assign n8778 = ~pi39 & ~n7861;
  assign n8779 = ~n8777 & ~n8778;
  assign n8780 = ~pi141 & ~n8779;
  assign n8781 = pi749 & ~n8780;
  assign n8782 = ~n8776 & n8781;
  assign n8783 = pi749 & ~n8771;
  assign n8784 = ~n8766 & ~n62902;
  assign n8785 = ~pi38 & ~n8784;
  assign n8786 = ~n8743 & n8756;
  assign n8787 = ~n7187 & n7357;
  assign n8788 = n7224 & n7356;
  assign n8789 = n7563 & n62904;
  assign n8790 = ~n7187 & n8084;
  assign n8791 = ~pi39 & n62857;
  assign n8792 = n7356 & n7565;
  assign n8793 = pi38 & ~n62905;
  assign n8794 = n8717 & n8793;
  assign n8795 = pi706 & ~n8794;
  assign n8796 = ~n62903 & n8795;
  assign n8797 = n62765 & ~n8796;
  assign n8798 = n62765 & ~n8733;
  assign n8799 = ~n8796 & n8798;
  assign n8800 = ~n8733 & n8797;
  assign n8801 = ~n8714 & ~n62906;
  assign n8802 = ~pi778 & ~n8801;
  assign n8803 = ~pi625 & n8801;
  assign n8804 = n62765 & n8732;
  assign n8805 = ~n8714 & ~n8804;
  assign n8806 = pi625 & n8805;
  assign n8807 = ~pi1153 & ~n8806;
  assign n8808 = ~n8803 & n8807;
  assign n8809 = ~pi141 & n8009;
  assign n8810 = pi141 & n62874;
  assign n8811 = ~pi38 & ~n8810;
  assign n8812 = ~n8809 & n8811;
  assign n8813 = n8085 & ~n8715;
  assign n8814 = pi706 & ~n8813;
  assign n8815 = ~n8812 & n8814;
  assign n8816 = ~pi141 & ~pi706;
  assign n8817 = ~n8091 & n8816;
  assign n8818 = n62765 & ~n8817;
  assign n8819 = ~n8815 & n8818;
  assign n8820 = ~n8714 & ~n8819;
  assign n8821 = pi625 & n8820;
  assign n8822 = ~pi141 & ~n8098;
  assign n8823 = ~pi625 & n8822;
  assign n8824 = pi1153 & ~n8823;
  assign n8825 = ~n8821 & n8824;
  assign n8826 = ~pi608 & ~n8825;
  assign n8827 = ~n8808 & n8826;
  assign n8828 = pi625 & n8801;
  assign n8829 = ~pi625 & n8805;
  assign n8830 = pi1153 & ~n8829;
  assign n8831 = ~n8828 & n8830;
  assign n8832 = ~pi625 & n8820;
  assign n8833 = pi625 & n8822;
  assign n8834 = ~pi1153 & ~n8833;
  assign n8835 = ~n8832 & n8834;
  assign n8836 = pi608 & ~n8835;
  assign n8837 = ~n8831 & n8836;
  assign n8838 = pi778 & ~n8837;
  assign n8839 = pi778 & ~n8827;
  assign n8840 = ~n8837 & n8839;
  assign n8841 = ~n8827 & n8838;
  assign n8842 = ~n8827 & ~n8837;
  assign n8843 = pi778 & ~n8842;
  assign n8844 = ~pi778 & n8801;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = ~n8802 & ~n62907;
  assign n8847 = ~pi609 & ~n62908;
  assign n8848 = ~pi778 & ~n8820;
  assign n8849 = ~n8825 & ~n8835;
  assign n8850 = pi778 & ~n8849;
  assign n8851 = ~n8848 & ~n8850;
  assign n8852 = pi609 & n8851;
  assign n8853 = ~pi1155 & ~n8852;
  assign n8854 = ~n8847 & n8853;
  assign n8855 = ~n8136 & ~n8822;
  assign n8856 = ~n8135 & ~n8805;
  assign n8857 = pi609 & n8856;
  assign n8858 = ~n8855 & ~n8857;
  assign n8859 = pi1155 & ~n8858;
  assign n8860 = ~pi660 & ~n8859;
  assign n8861 = ~n8854 & n8860;
  assign n8862 = pi609 & ~n62908;
  assign n8863 = ~pi609 & n8851;
  assign n8864 = pi1155 & ~n8863;
  assign n8865 = ~n8862 & n8864;
  assign n8866 = ~n8148 & ~n8822;
  assign n8867 = ~pi609 & n8856;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = ~pi1155 & ~n8868;
  assign n8870 = pi660 & ~n8869;
  assign n8871 = ~n8865 & n8870;
  assign n8872 = ~n8861 & ~n8871;
  assign n8873 = pi785 & ~n8872;
  assign n8874 = ~pi785 & ~n62908;
  assign n8875 = ~n8873 & ~n8874;
  assign n8876 = ~pi618 & ~n8875;
  assign n8877 = ~n62880 & ~n8851;
  assign n8878 = n62880 & ~n8822;
  assign n8879 = ~n62880 & n8851;
  assign n8880 = n62880 & n8822;
  assign n8881 = ~n8879 & ~n8880;
  assign n8882 = ~n8877 & ~n8878;
  assign n8883 = pi618 & ~n62909;
  assign n8884 = ~pi1154 & ~n8883;
  assign n8885 = ~n8876 & n8884;
  assign n8886 = n8135 & ~n8822;
  assign n8887 = ~n8856 & ~n8886;
  assign n8888 = ~pi785 & ~n8887;
  assign n8889 = ~n8859 & ~n8869;
  assign n8890 = pi785 & ~n8889;
  assign n8891 = ~n8888 & ~n8890;
  assign n8892 = pi618 & n8891;
  assign n8893 = ~pi618 & n8822;
  assign n8894 = pi1154 & ~n8893;
  assign n8895 = ~n8892 & n8894;
  assign n8896 = ~pi627 & ~n8895;
  assign n8897 = ~n8885 & n8896;
  assign n8898 = pi618 & ~n8875;
  assign n8899 = ~pi618 & ~n62909;
  assign n8900 = pi1154 & ~n8899;
  assign n8901 = ~n8898 & n8900;
  assign n8902 = ~pi618 & n8891;
  assign n8903 = pi618 & n8822;
  assign n8904 = ~pi1154 & ~n8903;
  assign n8905 = ~n8902 & n8904;
  assign n8906 = pi627 & ~n8905;
  assign n8907 = ~n8901 & n8906;
  assign n8908 = ~n8897 & ~n8907;
  assign n8909 = pi781 & ~n8908;
  assign n8910 = ~pi781 & ~n8875;
  assign n8911 = ~n8909 & ~n8910;
  assign n8912 = ~pi619 & ~n8911;
  assign n8913 = ~n62882 & ~n62909;
  assign n8914 = n62882 & n8822;
  assign n8915 = n62882 & ~n8822;
  assign n8916 = ~n62882 & n62909;
  assign n8917 = ~n8915 & ~n8916;
  assign n8918 = ~n8913 & ~n8914;
  assign n8919 = pi619 & n62910;
  assign n8920 = ~pi1159 & ~n8919;
  assign n8921 = ~n8912 & n8920;
  assign n8922 = ~pi781 & ~n8891;
  assign n8923 = ~n8895 & ~n8905;
  assign n8924 = pi781 & ~n8923;
  assign n8925 = ~n8922 & ~n8924;
  assign n8926 = pi619 & n8925;
  assign n8927 = ~pi619 & n8822;
  assign n8928 = pi1159 & ~n8927;
  assign n8929 = ~n8926 & n8928;
  assign n8930 = ~pi648 & ~n8929;
  assign n8931 = ~n8921 & n8930;
  assign n8932 = pi619 & ~n8911;
  assign n8933 = ~pi619 & n62910;
  assign n8934 = pi1159 & ~n8933;
  assign n8935 = ~n8932 & n8934;
  assign n8936 = ~pi619 & n8925;
  assign n8937 = pi619 & n8822;
  assign n8938 = ~pi1159 & ~n8937;
  assign n8939 = ~n8936 & n8938;
  assign n8940 = pi648 & ~n8939;
  assign n8941 = ~n8935 & n8940;
  assign n8942 = ~n8931 & ~n8941;
  assign n8943 = pi789 & ~n8942;
  assign n8944 = ~pi789 & ~n8911;
  assign n8945 = ~n8943 & ~n8944;
  assign n8946 = ~pi788 & n8945;
  assign n8947 = ~pi626 & n8945;
  assign n8948 = n8257 & ~n8822;
  assign n8949 = ~n8257 & ~n62910;
  assign n8950 = ~n8257 & n62910;
  assign n8951 = n8257 & n8822;
  assign n8952 = ~n8950 & ~n8951;
  assign n8953 = ~n8948 & ~n8949;
  assign n8954 = pi626 & n62911;
  assign n8955 = ~pi641 & ~n8954;
  assign n8956 = ~n8947 & n8955;
  assign n8957 = ~pi789 & ~n8925;
  assign n8958 = ~n8929 & ~n8939;
  assign n8959 = pi789 & ~n8958;
  assign n8960 = ~n8957 & ~n8959;
  assign n8961 = ~pi626 & n8960;
  assign n8962 = pi626 & n8822;
  assign n8963 = ~pi1158 & ~n8962;
  assign n8964 = ~n8961 & n8963;
  assign n8965 = ~n8267 & ~n8964;
  assign n8966 = ~n8956 & ~n8965;
  assign n8967 = pi626 & n8945;
  assign n8968 = ~pi626 & n62911;
  assign n8969 = pi641 & ~n8968;
  assign n8970 = ~n8967 & n8969;
  assign n8971 = pi626 & n8960;
  assign n8972 = ~pi626 & n8822;
  assign n8973 = pi1158 & ~n8972;
  assign n8974 = ~n8971 & n8973;
  assign n8975 = ~n8282 & ~n8974;
  assign n8976 = ~n8970 & ~n8975;
  assign n8977 = ~n8966 & ~n8976;
  assign n8978 = pi788 & ~n8977;
  assign n8979 = ~n8946 & ~n8978;
  assign n8980 = ~pi628 & n8979;
  assign n8981 = ~n8964 & ~n8974;
  assign n8982 = pi788 & ~n8981;
  assign n8983 = ~pi788 & ~n8960;
  assign n8984 = ~n8982 & ~n8983;
  assign n8985 = pi628 & n8984;
  assign n8986 = ~pi1156 & ~n8985;
  assign n8987 = ~n8980 & n8986;
  assign n8988 = ~n8303 & ~n62911;
  assign n8989 = n8303 & n8822;
  assign n8990 = n8303 & ~n8822;
  assign n8991 = ~n8303 & n62911;
  assign n8992 = ~n8990 & ~n8991;
  assign n8993 = ~n8988 & ~n8989;
  assign n8994 = pi628 & n62912;
  assign n8995 = ~pi628 & n8822;
  assign n8996 = pi1156 & ~n8995;
  assign n8997 = ~n8994 & n8996;
  assign n8998 = ~pi629 & ~n8997;
  assign n8999 = ~n8987 & n8998;
  assign n9000 = pi628 & n8979;
  assign n9001 = ~pi628 & n8984;
  assign n9002 = pi1156 & ~n9001;
  assign n9003 = ~n9000 & n9002;
  assign n9004 = ~pi628 & n62912;
  assign n9005 = pi628 & n8822;
  assign n9006 = ~pi1156 & ~n9005;
  assign n9007 = ~n9004 & n9006;
  assign n9008 = pi629 & ~n9007;
  assign n9009 = ~n9003 & n9008;
  assign n9010 = ~n8999 & ~n9009;
  assign n9011 = pi792 & ~n9010;
  assign n9012 = ~pi792 & n8979;
  assign n9013 = ~n9011 & ~n9012;
  assign n9014 = ~pi647 & ~n9013;
  assign n9015 = ~n8334 & n8984;
  assign n9016 = n8334 & n8822;
  assign n9017 = ~n9015 & ~n9016;
  assign n9018 = pi647 & ~n9017;
  assign n9019 = ~pi1157 & ~n9018;
  assign n9020 = ~n9014 & n9019;
  assign n9021 = ~pi792 & ~n62912;
  assign n9022 = ~n8997 & ~n9007;
  assign n9023 = pi792 & ~n9022;
  assign n9024 = ~n9021 & ~n9023;
  assign n9025 = pi647 & n9024;
  assign n9026 = ~pi647 & n8822;
  assign n9027 = pi1157 & ~n9026;
  assign n9028 = ~n9025 & n9027;
  assign n9029 = ~pi630 & ~n9028;
  assign n9030 = ~n9020 & n9029;
  assign n9031 = pi647 & ~n9013;
  assign n9032 = ~pi647 & ~n9017;
  assign n9033 = pi1157 & ~n9032;
  assign n9034 = ~n9031 & n9033;
  assign n9035 = ~pi647 & n9024;
  assign n9036 = pi647 & n8822;
  assign n9037 = ~pi1157 & ~n9036;
  assign n9038 = ~n9035 & n9037;
  assign n9039 = pi630 & ~n9038;
  assign n9040 = ~n9034 & n9039;
  assign n9041 = ~n9030 & ~n9040;
  assign n9042 = pi787 & ~n9041;
  assign n9043 = ~pi787 & ~n9013;
  assign n9044 = ~n9042 & ~n9043;
  assign n9045 = ~pi644 & ~n9044;
  assign n9046 = ~pi787 & ~n9024;
  assign n9047 = ~n9028 & ~n9038;
  assign n9048 = pi787 & ~n9047;
  assign n9049 = ~n9046 & ~n9048;
  assign n9050 = pi644 & n9049;
  assign n9051 = ~pi715 & ~n9050;
  assign n9052 = ~n9045 & n9051;
  assign n9053 = n8376 & ~n8822;
  assign n9054 = ~n8376 & n9017;
  assign n9055 = ~n8376 & ~n9017;
  assign n9056 = n8376 & n8822;
  assign n9057 = ~n9055 & ~n9056;
  assign n9058 = ~n9053 & ~n9054;
  assign n9059 = ~pi644 & ~n62913;
  assign n9060 = pi644 & n8822;
  assign n9061 = pi715 & ~n9060;
  assign n9062 = ~n9059 & n9061;
  assign n9063 = ~pi1160 & ~n9062;
  assign n9064 = ~n9052 & n9063;
  assign n9065 = pi644 & ~n9044;
  assign n9066 = ~pi644 & n9049;
  assign n9067 = pi715 & ~n9066;
  assign n9068 = ~n9065 & n9067;
  assign n9069 = pi644 & ~n62913;
  assign n9070 = ~pi644 & n8822;
  assign n9071 = ~pi715 & ~n9070;
  assign n9072 = ~n9069 & n9071;
  assign n9073 = pi1160 & ~n9072;
  assign n9074 = ~n9068 & n9073;
  assign n9075 = pi790 & ~n9074;
  assign n9076 = pi790 & ~n9064;
  assign n9077 = ~n9074 & n9076;
  assign n9078 = ~n9064 & n9075;
  assign n9079 = ~pi790 & n9044;
  assign n9080 = n62455 & ~n9079;
  assign n9081 = ~n62914 & n9080;
  assign n9082 = ~pi141 & ~n62455;
  assign n9083 = ~pi832 & ~n9082;
  assign n9084 = ~n9081 & n9083;
  assign n9085 = ~pi141 & ~n2923;
  assign n9086 = n8334 & ~n9085;
  assign n9087 = ~n8418 & n9085;
  assign n9088 = pi749 & n7316;
  assign n9089 = ~n9085 & ~n9088;
  assign n9090 = ~n8420 & ~n9089;
  assign n9091 = ~pi785 & ~n9090;
  assign n9092 = ~n8425 & ~n9089;
  assign n9093 = pi1155 & ~n9092;
  assign n9094 = ~n8428 & n9090;
  assign n9095 = ~pi1155 & ~n9094;
  assign n9096 = ~n9093 & ~n9095;
  assign n9097 = pi785 & ~n9096;
  assign n9098 = ~n9091 & ~n9097;
  assign n9099 = ~pi781 & ~n9098;
  assign n9100 = ~n8435 & n9098;
  assign n9101 = pi1154 & ~n9100;
  assign n9102 = ~n8438 & n9098;
  assign n9103 = ~pi1154 & ~n9102;
  assign n9104 = ~n9101 & ~n9103;
  assign n9105 = pi781 & ~n9104;
  assign n9106 = ~n9099 & ~n9105;
  assign n9107 = ~pi789 & ~n9106;
  assign n9108 = pi619 & n9106;
  assign n9109 = ~pi619 & n9085;
  assign n9110 = pi1159 & ~n9109;
  assign n9111 = ~n9108 & n9110;
  assign n9112 = ~pi619 & n9106;
  assign n9113 = pi619 & n9085;
  assign n9114 = ~pi1159 & ~n9113;
  assign n9115 = ~n9112 & n9114;
  assign n9116 = ~n9111 & ~n9115;
  assign n9117 = pi789 & ~n9116;
  assign n9118 = ~n9107 & ~n9117;
  assign n9119 = n8418 & n9118;
  assign n9120 = pi626 & n9118;
  assign n9121 = ~pi626 & n9085;
  assign n9122 = pi1158 & ~n9121;
  assign n9123 = ~n9120 & n9122;
  assign n9124 = ~pi626 & n9118;
  assign n9125 = pi626 & n9085;
  assign n9126 = ~pi1158 & ~n9125;
  assign n9127 = ~n9124 & n9126;
  assign n9128 = ~n9123 & ~n9127;
  assign n9129 = ~n9087 & ~n9119;
  assign n9130 = pi788 & n62915;
  assign n9131 = ~pi788 & n9118;
  assign n9132 = ~pi788 & ~n9118;
  assign n9133 = pi788 & ~n62915;
  assign n9134 = ~n9132 & ~n9133;
  assign n9135 = ~n9130 & ~n9131;
  assign n9136 = ~n8334 & ~n62916;
  assign n9137 = ~n8334 & n62916;
  assign n9138 = n8334 & n9085;
  assign n9139 = ~n9137 & ~n9138;
  assign n9140 = ~n9086 & ~n9136;
  assign n9141 = ~n8413 & n62917;
  assign n9142 = pi706 & n7564;
  assign n9143 = ~n9085 & ~n9142;
  assign n9144 = ~pi778 & n9143;
  assign n9145 = ~pi625 & n9142;
  assign n9146 = ~n9143 & ~n9145;
  assign n9147 = pi1153 & ~n9146;
  assign n9148 = ~pi1153 & ~n9085;
  assign n9149 = ~n9145 & n9148;
  assign n9150 = ~n9147 & ~n9149;
  assign n9151 = pi778 & ~n9150;
  assign n9152 = ~n9144 & ~n9151;
  assign n9153 = ~n8490 & n9152;
  assign n9154 = ~n8492 & n9153;
  assign n9155 = ~n8494 & n9154;
  assign n9156 = ~n8496 & n9155;
  assign n9157 = ~n8508 & n9156;
  assign n9158 = pi647 & ~n9157;
  assign n9159 = ~pi647 & ~n9085;
  assign n9160 = ~n9158 & ~n9159;
  assign n9161 = n8373 & ~n9160;
  assign n9162 = ~pi647 & n9157;
  assign n9163 = pi647 & n9085;
  assign n9164 = ~pi1157 & ~n9163;
  assign n9165 = ~n9162 & n9164;
  assign n9166 = pi630 & n9165;
  assign n9167 = ~n9161 & ~n9166;
  assign n9168 = ~n9141 & n9167;
  assign n9169 = pi787 & ~n9168;
  assign n9170 = n8525 & n9155;
  assign n9171 = ~n8302 & n62915;
  assign n9172 = ~n9170 & ~n9171;
  assign n9173 = pi788 & ~n9172;
  assign n9174 = ~n7187 & ~n9143;
  assign n9175 = pi625 & n9174;
  assign n9176 = n9089 & ~n9174;
  assign n9177 = ~n9175 & ~n9176;
  assign n9178 = n9148 & ~n9177;
  assign n9179 = ~pi608 & ~n9147;
  assign n9180 = ~n9178 & n9179;
  assign n9181 = pi1153 & n9089;
  assign n9182 = ~n9175 & n9181;
  assign n9183 = pi608 & ~n9149;
  assign n9184 = ~n9182 & n9183;
  assign n9185 = ~n9180 & ~n9184;
  assign n9186 = pi778 & ~n9185;
  assign n9187 = ~pi778 & ~n9176;
  assign n9188 = ~n9186 & ~n9187;
  assign n9189 = ~pi609 & ~n9188;
  assign n9190 = pi609 & n9152;
  assign n9191 = ~pi1155 & ~n9190;
  assign n9192 = ~n9189 & n9191;
  assign n9193 = ~pi660 & ~n9093;
  assign n9194 = ~n9192 & n9193;
  assign n9195 = pi609 & ~n9188;
  assign n9196 = ~pi609 & n9152;
  assign n9197 = pi1155 & ~n9196;
  assign n9198 = ~n9195 & n9197;
  assign n9199 = pi660 & ~n9095;
  assign n9200 = ~n9198 & n9199;
  assign n9201 = ~n9194 & ~n9200;
  assign n9202 = pi785 & ~n9201;
  assign n9203 = ~pi785 & ~n9188;
  assign n9204 = ~n9202 & ~n9203;
  assign n9205 = ~pi618 & ~n9204;
  assign n9206 = pi618 & n9153;
  assign n9207 = ~pi1154 & ~n9206;
  assign n9208 = ~n9205 & n9207;
  assign n9209 = ~pi627 & ~n9101;
  assign n9210 = ~n9208 & n9209;
  assign n9211 = pi618 & ~n9204;
  assign n9212 = ~pi618 & n9153;
  assign n9213 = pi1154 & ~n9212;
  assign n9214 = ~n9211 & n9213;
  assign n9215 = pi627 & ~n9103;
  assign n9216 = ~n9214 & n9215;
  assign n9217 = ~n9210 & ~n9216;
  assign n9218 = pi781 & ~n9217;
  assign n9219 = ~pi781 & ~n9204;
  assign n9220 = ~n9218 & ~n9219;
  assign n9221 = pi619 & ~n9220;
  assign n9222 = ~pi619 & n9154;
  assign n9223 = pi1159 & ~n9222;
  assign n9224 = ~n9221 & n9223;
  assign n9225 = pi648 & ~n9115;
  assign n9226 = ~n9224 & n9225;
  assign n9227 = ~pi619 & ~n9220;
  assign n9228 = pi619 & n9154;
  assign n9229 = ~pi1159 & ~n9228;
  assign n9230 = ~n9227 & n9229;
  assign n9231 = ~pi648 & ~n9111;
  assign n9232 = ~n9230 & n9231;
  assign n9233 = pi789 & ~n9232;
  assign n9234 = pi789 & ~n9226;
  assign n9235 = ~n9232 & n9234;
  assign n9236 = ~n9226 & n9233;
  assign n9237 = ~pi789 & n9220;
  assign n9238 = n62894 & ~n9237;
  assign n9239 = ~n62918 & n9238;
  assign n9240 = ~n9173 & ~n9239;
  assign n9241 = ~pi628 & n9240;
  assign n9242 = pi628 & ~n62916;
  assign n9243 = ~pi1156 & ~n9242;
  assign n9244 = ~n9241 & n9243;
  assign n9245 = n8606 & n9156;
  assign n9246 = ~pi629 & ~n9245;
  assign n9247 = ~n9244 & n9246;
  assign n9248 = pi628 & n9240;
  assign n9249 = ~pi628 & ~n62916;
  assign n9250 = pi1156 & ~n9249;
  assign n9251 = ~n9248 & n9250;
  assign n9252 = n8615 & n9156;
  assign n9253 = pi629 & ~n9252;
  assign n9254 = ~n9251 & n9253;
  assign n9255 = pi792 & ~n9254;
  assign n9256 = ~pi628 & ~n9240;
  assign n9257 = pi628 & n62916;
  assign n9258 = ~pi1156 & ~n9257;
  assign n9259 = ~n9256 & n9258;
  assign n9260 = ~n8605 & n9156;
  assign n9261 = pi1156 & ~n9260;
  assign n9262 = ~pi629 & ~n9261;
  assign n9263 = ~n9259 & n9262;
  assign n9264 = pi628 & ~n9240;
  assign n9265 = ~pi628 & n62916;
  assign n9266 = pi1156 & ~n9265;
  assign n9267 = ~n9264 & n9266;
  assign n9268 = ~n8614 & n9156;
  assign n9269 = ~pi1156 & ~n9268;
  assign n9270 = pi629 & ~n9269;
  assign n9271 = ~n9267 & n9270;
  assign n9272 = ~n9263 & ~n9271;
  assign n9273 = pi792 & ~n9272;
  assign n9274 = ~n9247 & n9255;
  assign n9275 = ~pi792 & ~n9240;
  assign n9276 = ~n8651 & ~n9275;
  assign n9277 = ~n62919 & n9276;
  assign n9278 = ~n62919 & ~n9275;
  assign n9279 = ~pi647 & ~n9278;
  assign n9280 = pi647 & ~n62917;
  assign n9281 = ~pi1157 & ~n9280;
  assign n9282 = ~n9279 & n9281;
  assign n9283 = pi647 & n9157;
  assign n9284 = ~pi647 & n9085;
  assign n9285 = pi1157 & ~n9284;
  assign n9286 = pi1157 & ~n9160;
  assign n9287 = ~n9283 & n9285;
  assign n9288 = ~pi630 & ~n62920;
  assign n9289 = ~n9282 & n9288;
  assign n9290 = pi647 & ~n9278;
  assign n9291 = ~pi647 & ~n62917;
  assign n9292 = pi1157 & ~n9291;
  assign n9293 = ~n9290 & n9292;
  assign n9294 = pi630 & ~n9165;
  assign n9295 = ~n9293 & n9294;
  assign n9296 = ~n9289 & ~n9295;
  assign n9297 = pi787 & ~n9296;
  assign n9298 = ~pi787 & ~n9278;
  assign n9299 = ~n9297 & ~n9298;
  assign n9300 = ~n9169 & ~n9277;
  assign n9301 = pi644 & ~n62921;
  assign n9302 = ~pi787 & ~n9157;
  assign n9303 = ~n9165 & ~n62920;
  assign n9304 = pi787 & ~n9303;
  assign n9305 = ~n9302 & ~n9304;
  assign n9306 = ~pi644 & n9305;
  assign n9307 = pi715 & ~n9306;
  assign n9308 = ~n9301 & n9307;
  assign n9309 = ~n8685 & ~n9085;
  assign n9310 = ~n8376 & n9136;
  assign n9311 = n8376 & ~n9085;
  assign n9312 = ~n8376 & n62917;
  assign n9313 = ~n9311 & ~n9312;
  assign n9314 = ~n9309 & ~n9310;
  assign n9315 = pi644 & n62922;
  assign n9316 = ~pi644 & n9085;
  assign n9317 = ~pi715 & ~n9316;
  assign n9318 = ~n9315 & n9317;
  assign n9319 = pi1160 & ~n9318;
  assign n9320 = ~n9308 & n9319;
  assign n9321 = ~pi644 & ~n62921;
  assign n9322 = pi644 & n9305;
  assign n9323 = ~pi715 & ~n9322;
  assign n9324 = ~n9321 & n9323;
  assign n9325 = ~pi644 & n62922;
  assign n9326 = pi644 & n9085;
  assign n9327 = pi715 & ~n9326;
  assign n9328 = ~n9325 & n9327;
  assign n9329 = ~pi1160 & ~n9328;
  assign n9330 = ~n9324 & n9329;
  assign n9331 = ~n9320 & ~n9330;
  assign n9332 = pi790 & ~n9331;
  assign n9333 = ~pi790 & ~n62921;
  assign n9334 = pi832 & ~n9333;
  assign n9335 = ~n9332 & n9334;
  assign po298 = ~n9084 & ~n9335;
  assign n9337 = pi142 & ~n62765;
  assign n9338 = ~pi142 & ~n7665;
  assign n9339 = pi142 & n62841;
  assign n9340 = pi743 & ~n9339;
  assign n9341 = pi743 & ~n9338;
  assign n9342 = ~n9339 & n9341;
  assign n9343 = ~n9338 & n9340;
  assign n9344 = pi142 & n7393;
  assign n9345 = ~pi142 & n7559;
  assign n9346 = ~pi743 & ~n9345;
  assign n9347 = ~n9344 & n9346;
  assign n9348 = pi142 & ~n62841;
  assign n9349 = ~pi142 & n7665;
  assign n9350 = pi743 & ~n9349;
  assign n9351 = ~n9348 & n9350;
  assign n9352 = pi142 & ~n7393;
  assign n9353 = ~pi142 & ~n7559;
  assign n9354 = ~pi743 & ~n9353;
  assign n9355 = ~n9352 & n9354;
  assign n9356 = ~n9351 & ~n9355;
  assign n9357 = ~n62923 & ~n9347;
  assign n9358 = pi735 & n62924;
  assign n9359 = pi142 & n7194;
  assign n9360 = ~pi142 & n62804;
  assign n9361 = pi743 & ~n9360;
  assign n9362 = ~n9359 & n9361;
  assign n9363 = pi142 & ~n7104;
  assign n9364 = ~pi743 & n9363;
  assign n9365 = ~n9359 & ~n9360;
  assign n9366 = pi743 & ~n9365;
  assign n9367 = ~pi743 & ~n9363;
  assign n9368 = ~n9366 & ~n9367;
  assign n9369 = ~n9362 & ~n9364;
  assign n9370 = ~pi735 & n62925;
  assign n9371 = pi735 & ~n62924;
  assign n9372 = ~pi735 & ~n62925;
  assign n9373 = ~n9371 & ~n9372;
  assign n9374 = ~n9358 & ~n9370;
  assign n9375 = n62393 & n62926;
  assign n9376 = ~pi142 & ~n7650;
  assign n9377 = pi142 & n7735;
  assign n9378 = pi743 & ~n9377;
  assign n9379 = ~n9376 & n9378;
  assign n9380 = ~pi142 & ~n7542;
  assign n9381 = pi142 & n7404;
  assign n9382 = ~pi743 & ~n9381;
  assign n9383 = ~n9380 & n9382;
  assign n9384 = ~pi142 & n7650;
  assign n9385 = pi142 & ~n7735;
  assign n9386 = pi743 & ~n9385;
  assign n9387 = ~n9384 & n9386;
  assign n9388 = ~pi142 & n7542;
  assign n9389 = pi142 & ~n7404;
  assign n9390 = ~pi743 & ~n9389;
  assign n9391 = ~n9388 & n9390;
  assign n9392 = ~n9387 & ~n9391;
  assign n9393 = ~n9379 & ~n9383;
  assign n9394 = pi735 & n62927;
  assign n9395 = pi142 & ~n62787;
  assign n9396 = ~pi743 & ~n9395;
  assign n9397 = pi142 & ~n7200;
  assign n9398 = pi743 & ~n7294;
  assign n9399 = ~n9397 & n9398;
  assign n9400 = ~n9396 & ~n9399;
  assign n9401 = ~pi735 & n9400;
  assign n9402 = pi735 & ~n62927;
  assign n9403 = ~pi735 & ~n9400;
  assign n9404 = ~n9402 & ~n9403;
  assign n9405 = ~n9394 & ~n9401;
  assign n9406 = ~n62393 & n62928;
  assign n9407 = ~n7118 & ~n9406;
  assign n9408 = ~n9375 & n9407;
  assign n9409 = pi743 & n7316;
  assign n9410 = pi743 & n7298;
  assign n9411 = n6950 & n9409;
  assign n9412 = ~pi735 & n62929;
  assign n9413 = pi142 & ~n6951;
  assign n9414 = pi142 & ~n6955;
  assign n9415 = n62380 & n9409;
  assign n9416 = ~n9414 & ~n9415;
  assign n9417 = ~n62857 & n9416;
  assign n9418 = pi735 & ~n6948;
  assign n9419 = ~n9417 & n9418;
  assign n9420 = ~n9413 & ~n9419;
  assign n9421 = ~n62929 & ~n9413;
  assign n9422 = ~pi735 & n9421;
  assign n9423 = ~n6948 & ~n9417;
  assign n9424 = pi735 & ~n9423;
  assign n9425 = ~n9413 & n9424;
  assign n9426 = ~n9422 & ~n9425;
  assign n9427 = ~n9412 & n9420;
  assign n9428 = n7118 & ~n62930;
  assign n9429 = ~pi215 & ~n9428;
  assign n9430 = ~n9408 & n9429;
  assign n9431 = pi142 & n7756;
  assign n9432 = ~pi142 & n7692;
  assign n9433 = pi743 & ~n9432;
  assign n9434 = ~n9431 & n9433;
  assign n9435 = pi142 & n62813;
  assign n9436 = ~pi142 & ~n7603;
  assign n9437 = ~pi743 & ~n9436;
  assign n9438 = ~pi743 & ~n9435;
  assign n9439 = ~n9436 & n9438;
  assign n9440 = ~n9435 & n9437;
  assign n9441 = pi142 & ~n7756;
  assign n9442 = ~pi142 & ~n7692;
  assign n9443 = pi743 & ~n9442;
  assign n9444 = ~n9441 & n9443;
  assign n9445 = pi142 & ~n62813;
  assign n9446 = ~pi142 & n7603;
  assign n9447 = ~pi743 & ~n9446;
  assign n9448 = ~n9445 & n9447;
  assign n9449 = ~n9444 & ~n9448;
  assign n9450 = ~n9434 & ~n62931;
  assign n9451 = pi735 & n62932;
  assign n9452 = pi142 & ~n7002;
  assign n9453 = ~pi743 & ~n9452;
  assign n9454 = pi142 & ~n7233;
  assign n9455 = pi743 & n7688;
  assign n9456 = ~n9454 & n9455;
  assign n9457 = ~n9453 & ~n9456;
  assign n9458 = ~pi735 & n9457;
  assign n9459 = pi735 & ~n62932;
  assign n9460 = ~pi735 & ~n9457;
  assign n9461 = ~n9459 & ~n9460;
  assign n9462 = ~n9451 & ~n9458;
  assign n9463 = ~n62393 & ~n62933;
  assign n9464 = ~pi142 & ~n7686;
  assign n9465 = pi142 & ~n7761;
  assign n9466 = pi743 & ~n9465;
  assign n9467 = pi743 & ~n9464;
  assign n9468 = ~n9465 & n9467;
  assign n9469 = ~n9464 & n9466;
  assign n9470 = pi142 & n7447;
  assign n9471 = ~pi142 & n7582;
  assign n9472 = ~pi743 & ~n9471;
  assign n9473 = ~n9470 & n9472;
  assign n9474 = pi142 & n7761;
  assign n9475 = ~pi142 & n7686;
  assign n9476 = pi743 & ~n9475;
  assign n9477 = ~n9474 & n9476;
  assign n9478 = pi142 & ~n7447;
  assign n9479 = ~pi142 & ~n7582;
  assign n9480 = ~pi743 & ~n9479;
  assign n9481 = ~n9478 & n9480;
  assign n9482 = ~n9477 & ~n9481;
  assign n9483 = ~n62934 & ~n9473;
  assign n9484 = pi735 & n62935;
  assign n9485 = pi142 & n7222;
  assign n9486 = n7327 & ~n9485;
  assign n9487 = pi743 & ~n9486;
  assign n9488 = pi142 & ~n62784;
  assign n9489 = ~pi743 & n9488;
  assign n9490 = ~pi743 & ~n9488;
  assign n9491 = pi743 & n7327;
  assign n9492 = ~n9485 & n9491;
  assign n9493 = ~n9490 & ~n9492;
  assign n9494 = ~n9487 & ~n9489;
  assign n9495 = ~pi735 & n62936;
  assign n9496 = pi735 & ~n62935;
  assign n9497 = ~pi735 & ~n62936;
  assign n9498 = ~n9496 & ~n9497;
  assign n9499 = ~n9484 & ~n9495;
  assign n9500 = n62393 & ~n62937;
  assign n9501 = pi215 & ~n9500;
  assign n9502 = ~n9463 & n9501;
  assign n9503 = ~n9430 & ~n9502;
  assign n9504 = pi299 & ~n9503;
  assign n9505 = n2971 & n62926;
  assign n9506 = ~n2971 & n62928;
  assign n9507 = ~n7034 & ~n9506;
  assign n9508 = ~n9505 & n9507;
  assign n9509 = n7034 & ~n62930;
  assign n9510 = ~pi223 & ~n9509;
  assign n9511 = ~n9508 & n9510;
  assign n9512 = ~n2971 & ~n62933;
  assign n9513 = n2971 & ~n62937;
  assign n9514 = pi223 & ~n9513;
  assign n9515 = ~n9512 & n9514;
  assign n9516 = ~n9511 & ~n9515;
  assign n9517 = ~pi299 & ~n9516;
  assign n9518 = pi39 & ~n9517;
  assign n9519 = pi39 & ~n9504;
  assign n9520 = ~n9517 & n9519;
  assign n9521 = ~n9504 & n9518;
  assign n9522 = pi142 & n7169;
  assign n9523 = ~n7827 & n9522;
  assign n9524 = ~pi142 & ~n7290;
  assign n9525 = ~n7865 & n9524;
  assign n9526 = pi299 & ~n9525;
  assign n9527 = ~n9523 & n9526;
  assign n9528 = pi142 & ~n7163;
  assign n9529 = n7822 & n9528;
  assign n9530 = ~pi142 & ~n7285;
  assign n9531 = ~n7863 & n9530;
  assign n9532 = ~pi299 & ~n9531;
  assign n9533 = ~n9529 & n9532;
  assign n9534 = pi743 & ~n9533;
  assign n9535 = ~n9527 & n9534;
  assign n9536 = ~pi142 & n7853;
  assign n9537 = pi142 & ~n7828;
  assign n9538 = ~n7290 & n9537;
  assign n9539 = pi299 & ~n9538;
  assign n9540 = ~n9536 & n9539;
  assign n9541 = ~pi142 & n7845;
  assign n9542 = pi142 & ~n7822;
  assign n9543 = ~n7285 & n9542;
  assign n9544 = ~pi299 & ~n9543;
  assign n9545 = ~n9541 & n9544;
  assign n9546 = ~n9540 & ~n9545;
  assign n9547 = ~pi743 & ~n9546;
  assign n9548 = pi735 & ~n9547;
  assign n9549 = ~n9529 & ~n9531;
  assign n9550 = pi743 & ~n9549;
  assign n9551 = ~pi743 & ~n9543;
  assign n9552 = ~n9541 & n9551;
  assign n9553 = ~pi299 & ~n9552;
  assign n9554 = ~n9550 & n9553;
  assign n9555 = ~n9523 & ~n9525;
  assign n9556 = pi743 & ~n9555;
  assign n9557 = ~pi743 & ~n9538;
  assign n9558 = ~n9536 & n9557;
  assign n9559 = pi299 & ~n9558;
  assign n9560 = pi299 & ~n9556;
  assign n9561 = ~n9558 & n9560;
  assign n9562 = ~n9556 & n9559;
  assign n9563 = ~n9554 & ~n62939;
  assign n9564 = pi735 & ~n9563;
  assign n9565 = ~n9535 & n9548;
  assign n9566 = pi142 & ~n6936;
  assign n9567 = ~pi743 & ~n9566;
  assign n9568 = pi743 & ~n9524;
  assign n9569 = ~n9566 & ~n9568;
  assign n9570 = ~n9524 & ~n9567;
  assign n9571 = ~n9522 & ~n62941;
  assign n9572 = pi299 & ~n9571;
  assign n9573 = pi743 & ~n9530;
  assign n9574 = ~n9528 & n9573;
  assign n9575 = pi142 & ~pi743;
  assign n9576 = ~n6940 & n9575;
  assign n9577 = ~pi299 & ~n9576;
  assign n9578 = ~n9574 & n9577;
  assign n9579 = ~n9572 & ~n9578;
  assign n9580 = ~pi735 & n9579;
  assign n9581 = ~pi39 & ~n9580;
  assign n9582 = ~n62940 & n9581;
  assign n9583 = ~n62938 & ~n9582;
  assign n9584 = ~pi38 & ~n9583;
  assign n9585 = pi39 & pi142;
  assign n9586 = pi38 & ~n9585;
  assign n9587 = pi735 & n7565;
  assign n9588 = pi735 & n7564;
  assign n9589 = pi735 & n7563;
  assign n9590 = n6955 & n9589;
  assign n9591 = n62380 & n9588;
  assign n9592 = ~n7187 & n62942;
  assign n9593 = pi735 & n62857;
  assign n9594 = n62380 & n9587;
  assign n9595 = n9416 & ~n62943;
  assign n9596 = ~pi39 & ~n9595;
  assign n9597 = n9586 & ~n9596;
  assign n9598 = n62765 & ~n9597;
  assign n9599 = ~n9584 & n9598;
  assign n9600 = ~n9337 & ~n9599;
  assign n9601 = pi625 & n9600;
  assign n9602 = ~n62393 & n9457;
  assign n9603 = n62393 & n62936;
  assign n9604 = pi215 & ~n9603;
  assign n9605 = ~n9602 & n9604;
  assign n9606 = n62393 & ~n62925;
  assign n9607 = ~n62393 & ~n9400;
  assign n9608 = ~n7118 & ~n9607;
  assign n9609 = n62393 & n62925;
  assign n9610 = ~n62393 & n9400;
  assign n9611 = ~n9609 & ~n9610;
  assign n9612 = ~n7118 & ~n9611;
  assign n9613 = ~n9606 & n9608;
  assign n9614 = n7118 & ~n9421;
  assign n9615 = ~pi215 & ~n9614;
  assign n9616 = ~n62944 & n9615;
  assign n9617 = ~n9605 & ~n9616;
  assign n9618 = pi299 & ~n9617;
  assign n9619 = n2971 & n62925;
  assign n9620 = ~n2971 & n9400;
  assign n9621 = ~n7034 & ~n9620;
  assign n9622 = ~n9619 & n9621;
  assign n9623 = n7034 & n9421;
  assign n9624 = ~pi223 & ~n9623;
  assign n9625 = ~n9622 & n9624;
  assign n9626 = ~n2971 & ~n9457;
  assign n9627 = n2971 & ~n62936;
  assign n9628 = pi223 & ~n9627;
  assign n9629 = ~n9626 & n9628;
  assign n9630 = ~pi299 & ~n9629;
  assign n9631 = ~n9625 & n9630;
  assign n9632 = pi39 & ~n9631;
  assign n9633 = ~n9618 & n9632;
  assign n9634 = ~pi39 & n9579;
  assign n9635 = ~pi38 & ~n9634;
  assign n9636 = ~n9633 & n9635;
  assign n9637 = ~pi39 & ~n9416;
  assign n9638 = n9586 & ~n9637;
  assign n9639 = n62765 & ~n9638;
  assign n9640 = ~n9636 & n9639;
  assign n9641 = ~n9337 & ~n9640;
  assign n9642 = ~pi625 & n9641;
  assign n9643 = pi1153 & ~n9642;
  assign n9644 = ~n9601 & n9643;
  assign n9645 = pi142 & ~n7942;
  assign n9646 = ~pi142 & ~n8022;
  assign n9647 = pi735 & ~n9646;
  assign n9648 = ~n9645 & n9647;
  assign n9649 = ~pi735 & n9363;
  assign n9650 = ~n9645 & ~n9646;
  assign n9651 = pi735 & ~n9650;
  assign n9652 = ~pi735 & ~n9363;
  assign n9653 = ~n9651 & ~n9652;
  assign n9654 = ~n9648 & ~n9649;
  assign n9655 = n2971 & n62945;
  assign n9656 = ~pi142 & n8015;
  assign n9657 = pi142 & n7948;
  assign n9658 = pi735 & ~n9657;
  assign n9659 = ~n9656 & n9658;
  assign n9660 = ~pi735 & n9395;
  assign n9661 = ~n9656 & ~n9657;
  assign n9662 = pi735 & ~n9661;
  assign n9663 = ~pi735 & ~n9395;
  assign n9664 = ~n9662 & ~n9663;
  assign n9665 = ~n9659 & ~n9660;
  assign n9666 = ~n2971 & n62946;
  assign n9667 = ~n7034 & ~n9666;
  assign n9668 = ~n9655 & n9667;
  assign n9669 = n6951 & n9589;
  assign n9670 = n6950 & n9588;
  assign n9671 = ~n9413 & ~n62947;
  assign n9672 = n7034 & n9671;
  assign n9673 = ~pi223 & ~n9672;
  assign n9674 = ~n9668 & n9673;
  assign n9675 = ~pi735 & ~n9452;
  assign n9676 = pi142 & ~n7965;
  assign n9677 = ~pi142 & n7689;
  assign n9678 = n7690 & n9677;
  assign n9679 = pi735 & ~n9678;
  assign n9680 = ~n9676 & n9679;
  assign n9681 = ~n9676 & ~n9678;
  assign n9682 = pi735 & ~n9681;
  assign n9683 = ~pi735 & n9452;
  assign n9684 = ~n9682 & ~n9683;
  assign n9685 = ~n9675 & ~n9680;
  assign n9686 = ~n2971 & n62948;
  assign n9687 = ~pi735 & ~n9488;
  assign n9688 = pi142 & ~n62863;
  assign n9689 = pi735 & ~n9677;
  assign n9690 = ~n9688 & n9689;
  assign n9691 = ~n9687 & ~n9690;
  assign n9692 = n2971 & ~n9691;
  assign n9693 = pi223 & ~n9692;
  assign n9694 = ~n9686 & n9693;
  assign n9695 = ~pi299 & ~n9694;
  assign n9696 = ~n9674 & n9695;
  assign n9697 = n62393 & n62945;
  assign n9698 = ~n62393 & n62946;
  assign n9699 = ~n7118 & ~n9698;
  assign n9700 = ~n9697 & n9699;
  assign n9701 = n7118 & n9671;
  assign n9702 = ~pi215 & ~n9701;
  assign n9703 = ~n9700 & n9702;
  assign n9704 = ~n62393 & n62948;
  assign n9705 = n62393 & ~n9691;
  assign n9706 = pi215 & ~n9705;
  assign n9707 = ~n9704 & n9706;
  assign n9708 = pi299 & ~n9707;
  assign n9709 = ~n9703 & n9708;
  assign n9710 = pi39 & ~n9709;
  assign n9711 = pi39 & ~n9696;
  assign n9712 = ~n9709 & n9711;
  assign n9713 = ~n9696 & n9710;
  assign n9714 = ~pi142 & ~n7867;
  assign n9715 = pi142 & n7830;
  assign n9716 = pi735 & ~n9715;
  assign n9717 = pi735 & ~n9714;
  assign n9718 = ~n9715 & n9717;
  assign n9719 = ~n9714 & n9716;
  assign n9720 = pi142 & ~pi735;
  assign n9721 = n62781 & n9720;
  assign n9722 = ~n62950 & ~n9721;
  assign n9723 = ~pi39 & ~n9722;
  assign n9724 = ~pi38 & ~n9723;
  assign n9725 = ~n62949 & n9724;
  assign n9726 = ~n9414 & ~n62942;
  assign n9727 = ~pi39 & ~n9726;
  assign n9728 = n9586 & ~n9727;
  assign n9729 = n62765 & ~n9728;
  assign n9730 = ~n9725 & n9729;
  assign n9731 = ~n9337 & ~n9730;
  assign n9732 = ~pi625 & n9731;
  assign n9733 = n62765 & ~n8089;
  assign n9734 = pi142 & ~n9733;
  assign n9735 = ~pi38 & ~pi87;
  assign n9736 = ~pi100 & n9735;
  assign n9737 = ~pi38 & n6791;
  assign n9738 = n6793 & n62951;
  assign n9739 = n6792 & n9738;
  assign n9740 = ~pi38 & n62765;
  assign n9741 = n6794 & n62951;
  assign n9742 = ~n62393 & ~n9452;
  assign n9743 = n62393 & ~n9488;
  assign n9744 = pi39 & pi215;
  assign n9745 = pi299 & n9744;
  assign n9746 = ~n9743 & n9745;
  assign n9747 = ~n9742 & n9746;
  assign n9748 = ~n62393 & n62787;
  assign n9749 = n62393 & n7104;
  assign n9750 = ~n62393 & ~n62787;
  assign n9751 = n2915 & n7119;
  assign n9752 = ~n9750 & ~n9751;
  assign n9753 = ~n7122 & ~n7124;
  assign n9754 = ~n9748 & ~n9749;
  assign n9755 = ~n7118 & n62953;
  assign n9756 = n2959 & ~n7126;
  assign n9757 = ~n9755 & n9756;
  assign n9758 = pi39 & ~n9757;
  assign n9759 = ~n7117 & n9758;
  assign n9760 = pi142 & ~n6946;
  assign n9761 = ~n9759 & n9760;
  assign n9762 = pi39 & ~n7117;
  assign n9763 = n9760 & ~n9762;
  assign n9764 = pi215 & ~n9743;
  assign n9765 = ~n9742 & n9764;
  assign n9766 = n62393 & n9363;
  assign n9767 = ~n62393 & n9395;
  assign n9768 = ~n7118 & ~n9767;
  assign n9769 = ~n62393 & ~n9395;
  assign n9770 = n62393 & ~n9363;
  assign n9771 = ~n9769 & ~n9770;
  assign n9772 = ~n7118 & ~n9771;
  assign n9773 = ~n9766 & n9768;
  assign n9774 = n7118 & ~n9413;
  assign n9775 = ~pi215 & ~n9774;
  assign n9776 = ~n62954 & n9775;
  assign n9777 = ~n9765 & ~n9776;
  assign n9778 = pi39 & pi299;
  assign n9779 = ~n9777 & n9778;
  assign n9780 = ~n9763 & ~n9779;
  assign n9781 = ~n9747 & ~n9761;
  assign n9782 = n62952 & ~n62955;
  assign n9783 = ~n9734 & ~n9782;
  assign n9784 = pi625 & n9783;
  assign n9785 = ~pi1153 & ~n9784;
  assign n9786 = ~n9732 & n9785;
  assign n9787 = pi608 & ~n9786;
  assign n9788 = ~n9644 & n9787;
  assign n9789 = ~pi625 & n9600;
  assign n9790 = pi625 & n9641;
  assign n9791 = ~pi1153 & ~n9790;
  assign n9792 = ~n9789 & n9791;
  assign n9793 = pi625 & n9731;
  assign n9794 = ~pi625 & n9783;
  assign n9795 = pi1153 & ~n9794;
  assign n9796 = ~n9793 & n9795;
  assign n9797 = ~pi608 & ~n9796;
  assign n9798 = ~n9792 & n9797;
  assign n9799 = ~n9788 & ~n9798;
  assign n9800 = pi778 & ~n9799;
  assign n9801 = ~pi778 & n9600;
  assign n9802 = ~n9800 & ~n9801;
  assign n9803 = ~pi609 & ~n9802;
  assign n9804 = ~pi778 & ~n9731;
  assign n9805 = ~n9786 & ~n9796;
  assign n9806 = pi778 & ~n9805;
  assign n9807 = ~n9804 & ~n9806;
  assign n9808 = pi609 & n9807;
  assign n9809 = ~pi1155 & ~n9808;
  assign n9810 = ~n9803 & n9809;
  assign n9811 = ~n8136 & ~n9783;
  assign n9812 = ~n8135 & ~n9641;
  assign n9813 = pi609 & n9812;
  assign n9814 = ~n9811 & ~n9813;
  assign n9815 = pi1155 & ~n9814;
  assign n9816 = ~pi660 & ~n9815;
  assign n9817 = ~n9810 & n9816;
  assign n9818 = pi609 & ~n9802;
  assign n9819 = ~pi609 & n9807;
  assign n9820 = pi1155 & ~n9819;
  assign n9821 = ~n9818 & n9820;
  assign n9822 = ~n8148 & ~n9783;
  assign n9823 = ~pi609 & n9812;
  assign n9824 = ~n9822 & ~n9823;
  assign n9825 = ~pi1155 & ~n9824;
  assign n9826 = pi660 & ~n9825;
  assign n9827 = ~n9821 & n9826;
  assign n9828 = ~n9817 & ~n9827;
  assign n9829 = pi785 & ~n9828;
  assign n9830 = ~pi785 & ~n9802;
  assign n9831 = ~n9829 & ~n9830;
  assign n9832 = ~pi618 & ~n9831;
  assign n9833 = ~n62880 & n9807;
  assign n9834 = n62880 & n9783;
  assign n9835 = ~n62880 & ~n9807;
  assign n9836 = n62880 & ~n9783;
  assign n9837 = ~n9835 & ~n9836;
  assign n9838 = ~n9833 & ~n9834;
  assign n9839 = pi618 & n62956;
  assign n9840 = ~pi1154 & ~n9839;
  assign n9841 = ~n9832 & n9840;
  assign n9842 = n8135 & ~n9783;
  assign n9843 = ~n9812 & ~n9842;
  assign n9844 = ~pi785 & ~n9843;
  assign n9845 = ~n9815 & ~n9825;
  assign n9846 = pi785 & ~n9845;
  assign n9847 = ~n9844 & ~n9846;
  assign n9848 = pi618 & n9847;
  assign n9849 = ~pi618 & n9783;
  assign n9850 = pi1154 & ~n9849;
  assign n9851 = ~n9848 & n9850;
  assign n9852 = ~pi627 & ~n9851;
  assign n9853 = ~n9841 & n9852;
  assign n9854 = pi618 & ~n9831;
  assign n9855 = ~pi618 & n62956;
  assign n9856 = pi1154 & ~n9855;
  assign n9857 = ~n9854 & n9856;
  assign n9858 = ~pi618 & n9847;
  assign n9859 = pi618 & n9783;
  assign n9860 = ~pi1154 & ~n9859;
  assign n9861 = ~n9858 & n9860;
  assign n9862 = pi627 & ~n9861;
  assign n9863 = ~n9857 & n9862;
  assign n9864 = ~n9853 & ~n9863;
  assign n9865 = pi781 & ~n9864;
  assign n9866 = ~pi781 & ~n9831;
  assign n9867 = ~n9865 & ~n9866;
  assign n9868 = ~pi619 & ~n9867;
  assign n9869 = n62882 & ~n9783;
  assign n9870 = ~n62882 & ~n62956;
  assign n9871 = ~n62882 & n62956;
  assign n9872 = n62882 & n9783;
  assign n9873 = ~n9871 & ~n9872;
  assign n9874 = ~n9869 & ~n9870;
  assign n9875 = pi619 & ~n62957;
  assign n9876 = ~pi1159 & ~n9875;
  assign n9877 = ~n9868 & n9876;
  assign n9878 = ~pi781 & ~n9847;
  assign n9879 = ~n9851 & ~n9861;
  assign n9880 = pi781 & ~n9879;
  assign n9881 = ~n9878 & ~n9880;
  assign n9882 = pi619 & n9881;
  assign n9883 = ~pi619 & n9783;
  assign n9884 = pi1159 & ~n9883;
  assign n9885 = ~n9882 & n9884;
  assign n9886 = ~pi648 & ~n9885;
  assign n9887 = ~n9877 & n9886;
  assign n9888 = pi619 & ~n9867;
  assign n9889 = ~pi619 & ~n62957;
  assign n9890 = pi1159 & ~n9889;
  assign n9891 = ~n9888 & n9890;
  assign n9892 = ~pi619 & n9881;
  assign n9893 = pi619 & n9783;
  assign n9894 = ~pi1159 & ~n9893;
  assign n9895 = ~n9892 & n9894;
  assign n9896 = pi648 & ~n9895;
  assign n9897 = ~n9891 & n9896;
  assign n9898 = ~n9887 & ~n9897;
  assign n9899 = pi789 & ~n9898;
  assign n9900 = ~pi789 & ~n9867;
  assign n9901 = ~n9899 & ~n9900;
  assign n9902 = ~pi788 & n9901;
  assign n9903 = ~pi626 & n9901;
  assign n9904 = ~n8257 & ~n62957;
  assign n9905 = n8257 & n9783;
  assign n9906 = n8257 & ~n9783;
  assign n9907 = ~n8257 & n62957;
  assign n9908 = ~n9906 & ~n9907;
  assign n9909 = ~n9904 & ~n9905;
  assign n9910 = pi626 & ~n62958;
  assign n9911 = ~pi641 & ~n9910;
  assign n9912 = ~n9903 & n9911;
  assign n9913 = ~pi789 & ~n9881;
  assign n9914 = ~n9885 & ~n9895;
  assign n9915 = pi789 & ~n9914;
  assign n9916 = ~n9913 & ~n9915;
  assign n9917 = ~pi626 & n9916;
  assign n9918 = pi626 & n9783;
  assign n9919 = ~pi1158 & ~n9918;
  assign n9920 = ~n9917 & n9919;
  assign n9921 = ~n8267 & ~n9920;
  assign n9922 = ~n9912 & ~n9921;
  assign n9923 = pi626 & n9901;
  assign n9924 = ~pi626 & ~n62958;
  assign n9925 = pi641 & ~n9924;
  assign n9926 = ~n9923 & n9925;
  assign n9927 = pi626 & n9916;
  assign n9928 = ~pi626 & n9783;
  assign n9929 = pi1158 & ~n9928;
  assign n9930 = ~n9927 & n9929;
  assign n9931 = ~n8282 & ~n9930;
  assign n9932 = ~n9926 & ~n9931;
  assign n9933 = ~n9922 & ~n9932;
  assign n9934 = pi788 & ~n9933;
  assign n9935 = ~n9902 & ~n9934;
  assign n9936 = ~pi628 & n9935;
  assign n9937 = ~n9920 & ~n9930;
  assign n9938 = pi788 & ~n9937;
  assign n9939 = ~pi788 & ~n9916;
  assign n9940 = ~n9938 & ~n9939;
  assign n9941 = pi628 & n9940;
  assign n9942 = ~pi1156 & ~n9941;
  assign n9943 = ~n9936 & n9942;
  assign n9944 = ~n8303 & n62958;
  assign n9945 = n8303 & n9783;
  assign n9946 = ~n8303 & ~n62958;
  assign n9947 = n8303 & ~n9783;
  assign n9948 = ~n9946 & ~n9947;
  assign n9949 = ~n9944 & ~n9945;
  assign n9950 = pi628 & n62959;
  assign n9951 = ~pi628 & n9783;
  assign n9952 = pi1156 & ~n9951;
  assign n9953 = ~n9950 & n9952;
  assign n9954 = ~pi629 & ~n9953;
  assign n9955 = ~n9943 & n9954;
  assign n9956 = pi628 & n9935;
  assign n9957 = ~pi628 & n9940;
  assign n9958 = pi1156 & ~n9957;
  assign n9959 = ~n9956 & n9958;
  assign n9960 = ~pi628 & n62959;
  assign n9961 = pi628 & n9783;
  assign n9962 = ~pi1156 & ~n9961;
  assign n9963 = ~n9960 & n9962;
  assign n9964 = pi629 & ~n9963;
  assign n9965 = ~n9959 & n9964;
  assign n9966 = ~n9955 & ~n9965;
  assign n9967 = pi792 & ~n9966;
  assign n9968 = ~pi792 & n9935;
  assign n9969 = ~n9967 & ~n9968;
  assign n9970 = ~pi647 & ~n9969;
  assign n9971 = ~n8334 & n9940;
  assign n9972 = n8334 & n9783;
  assign n9973 = ~n8334 & ~n9940;
  assign n9974 = n8334 & ~n9783;
  assign n9975 = ~n9973 & ~n9974;
  assign n9976 = ~n9971 & ~n9972;
  assign n9977 = pi647 & n62960;
  assign n9978 = ~pi1157 & ~n9977;
  assign n9979 = ~n9970 & n9978;
  assign n9980 = ~pi792 & ~n62959;
  assign n9981 = ~n9953 & ~n9963;
  assign n9982 = pi792 & ~n9981;
  assign n9983 = ~n9980 & ~n9982;
  assign n9984 = pi647 & n9983;
  assign n9985 = ~pi647 & n9783;
  assign n9986 = pi1157 & ~n9985;
  assign n9987 = ~n9984 & n9986;
  assign n9988 = ~pi630 & ~n9987;
  assign n9989 = ~n9979 & n9988;
  assign n9990 = pi647 & ~n9969;
  assign n9991 = ~pi647 & n62960;
  assign n9992 = pi1157 & ~n9991;
  assign n9993 = ~n9990 & n9992;
  assign n9994 = ~pi647 & n9983;
  assign n9995 = pi647 & n9783;
  assign n9996 = ~pi1157 & ~n9995;
  assign n9997 = ~n9994 & n9996;
  assign n9998 = pi630 & ~n9997;
  assign n9999 = ~n9993 & n9998;
  assign n10000 = ~n9989 & ~n9999;
  assign n10001 = pi787 & ~n10000;
  assign n10002 = ~pi787 & ~n9969;
  assign n10003 = ~n10001 & ~n10002;
  assign n10004 = ~pi644 & ~n10003;
  assign n10005 = ~pi787 & ~n9983;
  assign n10006 = ~n9987 & ~n9997;
  assign n10007 = pi787 & ~n10006;
  assign n10008 = ~n10005 & ~n10007;
  assign n10009 = pi644 & n10008;
  assign n10010 = ~pi715 & ~n10009;
  assign n10011 = ~n10004 & n10010;
  assign n10012 = n8376 & ~n9783;
  assign n10013 = ~n8376 & ~n62960;
  assign n10014 = ~n8376 & n62960;
  assign n10015 = n8376 & n9783;
  assign n10016 = ~n10014 & ~n10015;
  assign n10017 = ~n10012 & ~n10013;
  assign n10018 = ~pi644 & ~n62961;
  assign n10019 = pi644 & n9783;
  assign n10020 = pi715 & ~n10019;
  assign n10021 = ~n10018 & n10020;
  assign n10022 = ~pi1160 & ~n10021;
  assign n10023 = ~n10011 & n10022;
  assign n10024 = pi644 & ~n10003;
  assign n10025 = ~pi644 & n10008;
  assign n10026 = pi715 & ~n10025;
  assign n10027 = ~n10024 & n10026;
  assign n10028 = pi644 & ~n62961;
  assign n10029 = ~pi644 & n9783;
  assign n10030 = ~pi715 & ~n10029;
  assign n10031 = ~n10028 & n10030;
  assign n10032 = pi1160 & ~n10031;
  assign n10033 = ~n10027 & n10032;
  assign n10034 = pi790 & ~n10033;
  assign n10035 = pi790 & ~n10023;
  assign n10036 = ~n10033 & n10035;
  assign n10037 = ~n10023 & n10034;
  assign n10038 = ~pi790 & n10003;
  assign n10039 = n3475 & ~n10038;
  assign n10040 = ~n62962 & n10039;
  assign n10041 = ~pi142 & ~n3475;
  assign n10042 = ~pi57 & ~n10041;
  assign n10043 = ~n10040 & n10042;
  assign n10044 = pi57 & pi142;
  assign n10045 = ~pi832 & ~n10044;
  assign n10046 = ~n10043 & n10045;
  assign n10047 = pi142 & ~n2923;
  assign n10048 = ~n8418 & n10047;
  assign n10049 = ~n8135 & n9409;
  assign n10050 = pi609 & n10049;
  assign n10051 = pi1155 & ~n10047;
  assign n10052 = ~n10050 & n10051;
  assign n10053 = ~pi609 & n10049;
  assign n10054 = ~pi1155 & ~n10047;
  assign n10055 = ~n10053 & n10054;
  assign n10056 = ~n10052 & ~n10055;
  assign n10057 = pi785 & ~n10056;
  assign n10058 = ~pi785 & ~n10047;
  assign n10059 = ~n10049 & n10058;
  assign n10060 = ~n10057 & ~n10059;
  assign n10061 = ~pi781 & ~n10060;
  assign n10062 = pi618 & n10060;
  assign n10063 = ~pi618 & n10047;
  assign n10064 = pi1154 & ~n10063;
  assign n10065 = ~n10062 & n10064;
  assign n10066 = ~pi618 & n10060;
  assign n10067 = pi618 & n10047;
  assign n10068 = ~pi1154 & ~n10067;
  assign n10069 = ~n10066 & n10068;
  assign n10070 = ~n10065 & ~n10069;
  assign n10071 = pi781 & ~n10070;
  assign n10072 = ~n10061 & ~n10071;
  assign n10073 = ~pi789 & ~n10072;
  assign n10074 = pi619 & n10072;
  assign n10075 = ~pi619 & n10047;
  assign n10076 = pi1159 & ~n10075;
  assign n10077 = ~n10074 & n10076;
  assign n10078 = ~pi619 & n10072;
  assign n10079 = pi619 & n10047;
  assign n10080 = ~pi1159 & ~n10079;
  assign n10081 = ~n10078 & n10080;
  assign n10082 = ~n10077 & ~n10081;
  assign n10083 = pi789 & ~n10082;
  assign n10084 = ~n10073 & ~n10083;
  assign n10085 = n8418 & n10084;
  assign n10086 = pi626 & n10084;
  assign n10087 = ~pi626 & n10047;
  assign n10088 = pi1158 & ~n10087;
  assign n10089 = ~n10086 & n10088;
  assign n10090 = ~pi626 & n10084;
  assign n10091 = pi626 & n10047;
  assign n10092 = ~pi1158 & ~n10091;
  assign n10093 = ~n10090 & n10092;
  assign n10094 = ~n10089 & ~n10093;
  assign n10095 = ~n10048 & ~n10085;
  assign n10096 = ~n8302 & n62963;
  assign n10097 = pi625 & pi1153;
  assign n10098 = ~pi625 & ~pi1153;
  assign n10099 = pi778 & ~n10098;
  assign n10100 = ~pi625 & pi1153;
  assign n10101 = pi625 & ~pi1153;
  assign n10102 = ~n10100 & ~n10101;
  assign n10103 = pi778 & ~n10102;
  assign n10104 = ~n10097 & n10099;
  assign n10105 = n9588 & ~n62964;
  assign n10106 = ~n62880 & ~n62882;
  assign n10107 = n10105 & n10106;
  assign n10108 = ~n10047 & ~n10105;
  assign n10109 = ~n62880 & ~n10108;
  assign n10110 = ~n62882 & n10109;
  assign n10111 = n10106 & ~n10108;
  assign n10112 = ~n10047 & ~n62965;
  assign n10113 = ~n10047 & ~n10107;
  assign n10114 = n8257 & ~n10047;
  assign n10115 = n8525 & ~n10114;
  assign n10116 = ~n62966 & n10115;
  assign n10117 = ~n10096 & ~n10116;
  assign n10118 = pi788 & ~n10117;
  assign n10119 = pi625 & n9587;
  assign n10120 = ~n9409 & ~n10047;
  assign n10121 = ~n9587 & n10120;
  assign n10122 = ~n10119 & ~n10121;
  assign n10123 = ~pi1153 & ~n10122;
  assign n10124 = pi625 & n9588;
  assign n10125 = pi1153 & ~n10047;
  assign n10126 = ~n10124 & n10125;
  assign n10127 = ~pi608 & ~n10126;
  assign n10128 = ~n10123 & n10127;
  assign n10129 = ~n9409 & ~n10119;
  assign n10130 = pi1153 & ~n10129;
  assign n10131 = n9588 & n10098;
  assign n10132 = ~n10047 & ~n10131;
  assign n10133 = ~n10130 & n10132;
  assign n10134 = pi608 & ~n10133;
  assign n10135 = ~n10128 & ~n10134;
  assign n10136 = pi778 & ~n10135;
  assign n10137 = ~pi778 & ~n10121;
  assign n10138 = ~n10136 & ~n10137;
  assign n10139 = ~pi609 & ~n10138;
  assign n10140 = pi609 & ~n10108;
  assign n10141 = ~pi1155 & ~n10140;
  assign n10142 = ~n10139 & n10141;
  assign n10143 = ~pi660 & ~n10052;
  assign n10144 = ~n10142 & n10143;
  assign n10145 = pi609 & ~n10138;
  assign n10146 = ~pi609 & ~n10108;
  assign n10147 = pi1155 & ~n10146;
  assign n10148 = ~n10145 & n10147;
  assign n10149 = pi660 & ~n10055;
  assign n10150 = ~n10148 & n10149;
  assign n10151 = ~n10144 & ~n10150;
  assign n10152 = pi785 & ~n10151;
  assign n10153 = ~pi785 & ~n10138;
  assign n10154 = ~n10152 & ~n10153;
  assign n10155 = ~pi618 & ~n10154;
  assign n10156 = n62880 & ~n10047;
  assign n10157 = ~n62880 & n10105;
  assign n10158 = ~n10047 & ~n10157;
  assign n10159 = ~n10047 & ~n10109;
  assign n10160 = ~n10108 & ~n10156;
  assign n10161 = pi618 & ~n62967;
  assign n10162 = ~pi1154 & ~n10161;
  assign n10163 = ~n10155 & n10162;
  assign n10164 = ~pi627 & ~n10065;
  assign n10165 = ~n10163 & n10164;
  assign n10166 = pi618 & ~n10154;
  assign n10167 = ~pi618 & ~n62967;
  assign n10168 = pi1154 & ~n10167;
  assign n10169 = ~n10166 & n10168;
  assign n10170 = pi627 & ~n10069;
  assign n10171 = ~n10169 & n10170;
  assign n10172 = ~n10165 & ~n10171;
  assign n10173 = pi781 & ~n10172;
  assign n10174 = ~pi781 & ~n10154;
  assign n10175 = ~n10173 & ~n10174;
  assign n10176 = pi619 & ~n10175;
  assign n10177 = ~pi619 & ~n62966;
  assign n10178 = pi1159 & ~n10177;
  assign n10179 = ~n10176 & n10178;
  assign n10180 = pi648 & ~n10081;
  assign n10181 = ~n10179 & n10180;
  assign n10182 = ~pi619 & ~n10175;
  assign n10183 = pi619 & ~n62966;
  assign n10184 = ~pi1159 & ~n10183;
  assign n10185 = ~n10182 & n10184;
  assign n10186 = ~pi648 & ~n10077;
  assign n10187 = ~n10185 & n10186;
  assign n10188 = pi789 & ~n10187;
  assign n10189 = pi789 & ~n10181;
  assign n10190 = ~n10187 & n10189;
  assign n10191 = ~n10181 & n10188;
  assign n10192 = ~pi789 & n10175;
  assign n10193 = n62894 & ~n10192;
  assign n10194 = ~n62968 & n10193;
  assign n10195 = ~n10118 & ~n10194;
  assign n10196 = ~pi628 & n10195;
  assign n10197 = pi788 & n62963;
  assign n10198 = ~pi788 & n10084;
  assign n10199 = ~pi788 & ~n10084;
  assign n10200 = pi788 & ~n62963;
  assign n10201 = ~n10199 & ~n10200;
  assign n10202 = ~n10197 & ~n10198;
  assign n10203 = pi628 & ~n62969;
  assign n10204 = ~pi1156 & ~n10203;
  assign n10205 = ~n10196 & n10204;
  assign n10206 = ~n8257 & ~n8303;
  assign n10207 = n10106 & n10206;
  assign n10208 = n62965 & n10206;
  assign n10209 = ~n10108 & n10207;
  assign n10210 = pi628 & n62970;
  assign n10211 = ~n10047 & ~n10210;
  assign n10212 = pi1156 & ~n10211;
  assign n10213 = ~pi629 & ~n10212;
  assign n10214 = ~n10205 & n10213;
  assign n10215 = pi628 & n10195;
  assign n10216 = ~pi628 & ~n62969;
  assign n10217 = pi1156 & ~n10216;
  assign n10218 = ~n10215 & n10217;
  assign n10219 = ~pi628 & n62970;
  assign n10220 = ~n10047 & ~n10219;
  assign n10221 = ~pi1156 & ~n10220;
  assign n10222 = pi629 & ~n10221;
  assign n10223 = ~n10218 & n10222;
  assign n10224 = ~pi628 & ~n10195;
  assign n10225 = pi628 & n62969;
  assign n10226 = ~pi1156 & ~n10225;
  assign n10227 = ~n10224 & n10226;
  assign n10228 = pi1156 & ~n10047;
  assign n10229 = ~n10210 & n10228;
  assign n10230 = ~pi629 & ~n10229;
  assign n10231 = ~n10227 & n10230;
  assign n10232 = pi628 & ~n10195;
  assign n10233 = ~pi628 & n62969;
  assign n10234 = pi1156 & ~n10233;
  assign n10235 = ~n10232 & n10234;
  assign n10236 = ~pi1156 & ~n10047;
  assign n10237 = ~n10219 & n10236;
  assign n10238 = pi629 & ~n10237;
  assign n10239 = ~n10235 & n10238;
  assign n10240 = ~n10231 & ~n10239;
  assign n10241 = ~n10214 & ~n10223;
  assign n10242 = pi792 & n62971;
  assign n10243 = ~pi792 & n10195;
  assign n10244 = pi792 & ~n62971;
  assign n10245 = ~pi792 & ~n10195;
  assign n10246 = ~n10244 & ~n10245;
  assign n10247 = ~n10242 & ~n10243;
  assign n10248 = ~pi647 & ~n62972;
  assign n10249 = ~n8334 & n62969;
  assign n10250 = n8334 & n10047;
  assign n10251 = n8334 & ~n10047;
  assign n10252 = ~n8334 & ~n62969;
  assign n10253 = ~n10251 & ~n10252;
  assign n10254 = ~n10249 & ~n10250;
  assign n10255 = pi647 & n62973;
  assign n10256 = ~pi1157 & ~n10255;
  assign n10257 = ~n10248 & n10256;
  assign n10258 = ~n62892 & n62970;
  assign n10259 = pi647 & n10258;
  assign n10260 = pi1157 & ~n10047;
  assign n10261 = ~n10259 & n10260;
  assign n10262 = ~pi630 & ~n10261;
  assign n10263 = ~n10257 & n10262;
  assign n10264 = pi647 & ~n62972;
  assign n10265 = ~pi647 & n62973;
  assign n10266 = pi1157 & ~n10265;
  assign n10267 = ~n10264 & n10266;
  assign n10268 = ~pi647 & n10258;
  assign n10269 = ~pi1157 & ~n10047;
  assign n10270 = ~n10268 & n10269;
  assign n10271 = pi630 & ~n10270;
  assign n10272 = ~n10267 & n10271;
  assign n10273 = ~pi647 & n62972;
  assign n10274 = pi647 & ~n62973;
  assign n10275 = ~pi1157 & ~n10274;
  assign n10276 = ~n10273 & n10275;
  assign n10277 = ~n10047 & ~n10259;
  assign n10278 = pi1157 & ~n10277;
  assign n10279 = ~pi630 & ~n10278;
  assign n10280 = ~n10276 & n10279;
  assign n10281 = pi647 & n62972;
  assign n10282 = ~pi647 & ~n62973;
  assign n10283 = pi1157 & ~n10282;
  assign n10284 = ~n10281 & n10283;
  assign n10285 = ~n10047 & ~n10268;
  assign n10286 = ~pi1157 & ~n10285;
  assign n10287 = pi630 & ~n10286;
  assign n10288 = ~n10284 & n10287;
  assign n10289 = ~n10280 & ~n10288;
  assign n10290 = ~n10263 & ~n10272;
  assign n10291 = pi787 & n62974;
  assign n10292 = ~pi787 & ~n62972;
  assign n10293 = pi787 & ~n62974;
  assign n10294 = ~pi787 & n62972;
  assign n10295 = ~n10293 & ~n10294;
  assign n10296 = ~n10291 & ~n10292;
  assign n10297 = pi644 & n62975;
  assign n10298 = pi787 & ~n8644;
  assign n10299 = n10258 & ~n10298;
  assign n10300 = ~n10047 & ~n10299;
  assign n10301 = ~pi644 & ~n10300;
  assign n10302 = pi715 & ~n10301;
  assign n10303 = ~n10297 & n10302;
  assign n10304 = n8376 & ~n10047;
  assign n10305 = ~n8376 & ~n62973;
  assign n10306 = ~n8376 & n62973;
  assign n10307 = n8376 & n10047;
  assign n10308 = ~n10306 & ~n10307;
  assign n10309 = ~n10304 & ~n10305;
  assign n10310 = pi644 & ~n62976;
  assign n10311 = ~pi644 & n10047;
  assign n10312 = ~pi715 & ~n10311;
  assign n10313 = ~n10310 & n10312;
  assign n10314 = pi1160 & ~n10313;
  assign n10315 = ~n10303 & n10314;
  assign n10316 = ~pi644 & n62975;
  assign n10317 = pi644 & ~n10300;
  assign n10318 = ~pi715 & ~n10317;
  assign n10319 = ~n10316 & n10318;
  assign n10320 = ~pi644 & ~n62976;
  assign n10321 = pi644 & n10047;
  assign n10322 = pi715 & ~n10321;
  assign n10323 = ~n10320 & n10322;
  assign n10324 = ~pi1160 & ~n10323;
  assign n10325 = ~n10319 & n10324;
  assign n10326 = ~n10315 & ~n10325;
  assign n10327 = pi790 & ~n10326;
  assign n10328 = ~pi790 & n62975;
  assign n10329 = pi832 & ~n10328;
  assign n10330 = ~n10327 & n10329;
  assign po299 = ~n10046 & ~n10330;
  assign n10332 = pi143 & ~n62765;
  assign n10333 = ~pi143 & ~n8091;
  assign n10334 = pi774 & ~n10333;
  assign n10335 = pi38 & ~pi39;
  assign n10336 = n7316 & n10335;
  assign n10337 = pi38 & n7359;
  assign n10338 = n62380 & n10336;
  assign n10339 = ~pi38 & n7351;
  assign n10340 = pi143 & ~n10339;
  assign n10341 = ~pi38 & ~n62802;
  assign n10342 = pi38 & ~n62904;
  assign n10343 = ~n10341 & ~n10342;
  assign n10344 = ~pi143 & ~pi774;
  assign n10345 = n10343 & n10344;
  assign n10346 = ~n10340 & ~n10345;
  assign n10347 = ~n62977 & ~n10346;
  assign n10348 = ~n10334 & ~n10347;
  assign n10349 = ~pi687 & n10348;
  assign n10350 = n7357 & ~n7408;
  assign n10351 = pi38 & n10350;
  assign n10352 = ~pi38 & ~n8759;
  assign n10353 = ~n10351 & ~n10352;
  assign n10354 = ~pi143 & n10353;
  assign n10355 = ~pi38 & n8763;
  assign n10356 = pi143 & n10355;
  assign n10357 = pi38 & n62905;
  assign n10358 = pi774 & ~n10357;
  assign n10359 = ~n10356 & n10358;
  assign n10360 = ~n10354 & n10359;
  assign n10361 = ~pi38 & ~n8775;
  assign n10362 = pi38 & ~n62856;
  assign n10363 = ~n10361 & ~n10362;
  assign n10364 = pi143 & n10363;
  assign n10365 = ~pi38 & n8778;
  assign n10366 = ~pi39 & n7744;
  assign n10367 = pi38 & ~n10366;
  assign n10368 = ~n8777 & ~n10367;
  assign n10369 = ~pi38 & ~n8778;
  assign n10370 = pi38 & n7615;
  assign n10371 = n7357 & n10370;
  assign n10372 = n7744 & n10335;
  assign n10373 = ~n10365 & ~n10367;
  assign n10374 = ~n10369 & ~n62978;
  assign n10375 = ~n8777 & n62979;
  assign n10376 = ~pi38 & n8779;
  assign n10377 = ~n62978 & ~n10376;
  assign n10378 = ~n10365 & n10368;
  assign n10379 = ~pi143 & ~n62980;
  assign n10380 = ~pi774 & ~n10379;
  assign n10381 = ~n10364 & n10380;
  assign n10382 = pi687 & ~n10381;
  assign n10383 = ~n10360 & n10382;
  assign n10384 = n62765 & ~n10383;
  assign n10385 = n62765 & ~n10349;
  assign n10386 = ~n10383 & n10385;
  assign n10387 = ~n10349 & n10384;
  assign n10388 = ~n10332 & ~n62981;
  assign n10389 = ~pi625 & n10388;
  assign n10390 = n62765 & ~n10348;
  assign n10391 = ~n10332 & ~n10390;
  assign n10392 = pi625 & n10391;
  assign n10393 = ~pi1153 & ~n10392;
  assign n10394 = ~n10389 & n10393;
  assign n10395 = ~pi143 & n8009;
  assign n10396 = pi143 & n62874;
  assign n10397 = ~pi38 & ~n10396;
  assign n10398 = ~n10395 & n10397;
  assign n10399 = ~pi143 & ~n7357;
  assign n10400 = n8085 & ~n10399;
  assign n10401 = pi687 & ~n10400;
  assign n10402 = ~n10398 & n10401;
  assign n10403 = ~pi687 & n10333;
  assign n10404 = n62765 & ~n10403;
  assign n10405 = n62765 & ~n10402;
  assign n10406 = ~n10403 & n10405;
  assign n10407 = ~n10402 & n10404;
  assign n10408 = ~n10332 & ~n62982;
  assign n10409 = pi625 & n10408;
  assign n10410 = ~pi143 & ~n8098;
  assign n10411 = ~pi625 & n10410;
  assign n10412 = pi1153 & ~n10411;
  assign n10413 = ~n10409 & n10412;
  assign n10414 = ~pi608 & ~n10413;
  assign n10415 = ~n10394 & n10414;
  assign n10416 = pi625 & n10388;
  assign n10417 = ~pi625 & n10391;
  assign n10418 = pi1153 & ~n10417;
  assign n10419 = ~n10416 & n10418;
  assign n10420 = ~pi625 & n10408;
  assign n10421 = pi625 & n10410;
  assign n10422 = ~pi1153 & ~n10421;
  assign n10423 = ~n10420 & n10422;
  assign n10424 = pi608 & ~n10423;
  assign n10425 = ~n10419 & n10424;
  assign n10426 = ~n10415 & ~n10425;
  assign n10427 = pi778 & ~n10426;
  assign n10428 = ~pi778 & n10388;
  assign n10429 = ~pi778 & ~n10388;
  assign n10430 = pi778 & ~n10425;
  assign n10431 = ~n10415 & n10430;
  assign n10432 = ~n10429 & ~n10431;
  assign n10433 = ~n10427 & ~n10428;
  assign n10434 = ~pi609 & n62983;
  assign n10435 = ~pi778 & ~n10408;
  assign n10436 = ~n10413 & ~n10423;
  assign n10437 = pi778 & ~n10436;
  assign n10438 = ~n10435 & ~n10437;
  assign n10439 = pi609 & n10438;
  assign n10440 = ~pi1155 & ~n10439;
  assign n10441 = ~n10434 & n10440;
  assign n10442 = ~n8136 & ~n10410;
  assign n10443 = ~n8135 & ~n10391;
  assign n10444 = pi609 & n10443;
  assign n10445 = ~n10442 & ~n10444;
  assign n10446 = pi1155 & ~n10445;
  assign n10447 = ~pi660 & ~n10446;
  assign n10448 = ~n10441 & n10447;
  assign n10449 = pi609 & n62983;
  assign n10450 = ~pi609 & n10438;
  assign n10451 = pi1155 & ~n10450;
  assign n10452 = ~n10449 & n10451;
  assign n10453 = ~n8148 & ~n10410;
  assign n10454 = ~pi609 & n10443;
  assign n10455 = ~n10453 & ~n10454;
  assign n10456 = ~pi1155 & ~n10455;
  assign n10457 = pi660 & ~n10456;
  assign n10458 = ~n10452 & n10457;
  assign n10459 = ~n10448 & ~n10458;
  assign n10460 = pi785 & ~n10459;
  assign n10461 = ~pi785 & n62983;
  assign n10462 = ~n10460 & ~n10461;
  assign n10463 = ~pi618 & ~n10462;
  assign n10464 = ~n62880 & ~n10438;
  assign n10465 = n62880 & ~n10410;
  assign n10466 = ~n62880 & n10438;
  assign n10467 = n62880 & n10410;
  assign n10468 = ~n10466 & ~n10467;
  assign n10469 = ~n10464 & ~n10465;
  assign n10470 = pi618 & ~n62984;
  assign n10471 = ~pi1154 & ~n10470;
  assign n10472 = ~n10463 & n10471;
  assign n10473 = n8135 & ~n10410;
  assign n10474 = ~n10443 & ~n10473;
  assign n10475 = ~pi785 & ~n10474;
  assign n10476 = ~n10446 & ~n10456;
  assign n10477 = pi785 & ~n10476;
  assign n10478 = ~n10475 & ~n10477;
  assign n10479 = pi618 & n10478;
  assign n10480 = ~pi618 & n10410;
  assign n10481 = pi1154 & ~n10480;
  assign n10482 = ~n10479 & n10481;
  assign n10483 = ~pi627 & ~n10482;
  assign n10484 = ~n10472 & n10483;
  assign n10485 = pi618 & ~n10462;
  assign n10486 = ~pi618 & ~n62984;
  assign n10487 = pi1154 & ~n10486;
  assign n10488 = ~n10485 & n10487;
  assign n10489 = ~pi618 & n10478;
  assign n10490 = pi618 & n10410;
  assign n10491 = ~pi1154 & ~n10490;
  assign n10492 = ~n10489 & n10491;
  assign n10493 = pi627 & ~n10492;
  assign n10494 = ~n10488 & n10493;
  assign n10495 = ~n10484 & ~n10494;
  assign n10496 = pi781 & ~n10495;
  assign n10497 = ~pi781 & ~n10462;
  assign n10498 = ~n10496 & ~n10497;
  assign n10499 = ~pi619 & ~n10498;
  assign n10500 = ~n62882 & ~n62984;
  assign n10501 = n62882 & n10410;
  assign n10502 = n62882 & ~n10410;
  assign n10503 = ~n62882 & n62984;
  assign n10504 = ~n10502 & ~n10503;
  assign n10505 = ~n10500 & ~n10501;
  assign n10506 = pi619 & n62985;
  assign n10507 = ~pi1159 & ~n10506;
  assign n10508 = ~n10499 & n10507;
  assign n10509 = ~pi781 & ~n10478;
  assign n10510 = ~n10482 & ~n10492;
  assign n10511 = pi781 & ~n10510;
  assign n10512 = ~n10509 & ~n10511;
  assign n10513 = pi619 & n10512;
  assign n10514 = ~pi619 & n10410;
  assign n10515 = pi1159 & ~n10514;
  assign n10516 = ~n10513 & n10515;
  assign n10517 = ~pi648 & ~n10516;
  assign n10518 = ~n10508 & n10517;
  assign n10519 = pi619 & ~n10498;
  assign n10520 = ~pi619 & n62985;
  assign n10521 = pi1159 & ~n10520;
  assign n10522 = ~n10519 & n10521;
  assign n10523 = ~pi619 & n10512;
  assign n10524 = pi619 & n10410;
  assign n10525 = ~pi1159 & ~n10524;
  assign n10526 = ~n10523 & n10525;
  assign n10527 = pi648 & ~n10526;
  assign n10528 = ~n10522 & n10527;
  assign n10529 = ~n10518 & ~n10528;
  assign n10530 = pi789 & ~n10529;
  assign n10531 = ~pi789 & ~n10498;
  assign n10532 = ~n10530 & ~n10531;
  assign n10533 = ~pi788 & n10532;
  assign n10534 = ~pi626 & n10532;
  assign n10535 = n8257 & ~n10410;
  assign n10536 = ~n8257 & ~n62985;
  assign n10537 = ~n8257 & n62985;
  assign n10538 = n8257 & n10410;
  assign n10539 = ~n10537 & ~n10538;
  assign n10540 = ~n10535 & ~n10536;
  assign n10541 = pi626 & n62986;
  assign n10542 = ~pi641 & ~n10541;
  assign n10543 = ~n10534 & n10542;
  assign n10544 = ~pi789 & ~n10512;
  assign n10545 = ~n10516 & ~n10526;
  assign n10546 = pi789 & ~n10545;
  assign n10547 = ~n10544 & ~n10546;
  assign n10548 = ~pi626 & n10547;
  assign n10549 = pi626 & n10410;
  assign n10550 = ~pi1158 & ~n10549;
  assign n10551 = ~n10548 & n10550;
  assign n10552 = ~n8267 & ~n10551;
  assign n10553 = ~n10543 & ~n10552;
  assign n10554 = pi626 & n10532;
  assign n10555 = ~pi626 & n62986;
  assign n10556 = pi641 & ~n10555;
  assign n10557 = ~n10554 & n10556;
  assign n10558 = pi626 & n10547;
  assign n10559 = ~pi626 & n10410;
  assign n10560 = pi1158 & ~n10559;
  assign n10561 = ~n10558 & n10560;
  assign n10562 = ~n8282 & ~n10561;
  assign n10563 = ~n10557 & ~n10562;
  assign n10564 = ~n10553 & ~n10563;
  assign n10565 = pi788 & ~n10564;
  assign n10566 = ~n10533 & ~n10565;
  assign n10567 = ~pi628 & n10566;
  assign n10568 = ~n10551 & ~n10561;
  assign n10569 = pi788 & ~n10568;
  assign n10570 = ~pi788 & ~n10547;
  assign n10571 = ~n10569 & ~n10570;
  assign n10572 = pi628 & n10571;
  assign n10573 = ~pi1156 & ~n10572;
  assign n10574 = ~n10567 & n10573;
  assign n10575 = ~n8303 & ~n62986;
  assign n10576 = n8303 & n10410;
  assign n10577 = n8303 & ~n10410;
  assign n10578 = ~n8303 & n62986;
  assign n10579 = ~n10577 & ~n10578;
  assign n10580 = ~n10575 & ~n10576;
  assign n10581 = pi628 & n62987;
  assign n10582 = ~pi628 & n10410;
  assign n10583 = pi1156 & ~n10582;
  assign n10584 = ~n10581 & n10583;
  assign n10585 = ~pi629 & ~n10584;
  assign n10586 = ~n10574 & n10585;
  assign n10587 = pi628 & n10566;
  assign n10588 = ~pi628 & n10571;
  assign n10589 = pi1156 & ~n10588;
  assign n10590 = ~n10587 & n10589;
  assign n10591 = ~pi628 & n62987;
  assign n10592 = pi628 & n10410;
  assign n10593 = ~pi1156 & ~n10592;
  assign n10594 = ~n10591 & n10593;
  assign n10595 = pi629 & ~n10594;
  assign n10596 = ~n10590 & n10595;
  assign n10597 = ~n10586 & ~n10596;
  assign n10598 = pi792 & ~n10597;
  assign n10599 = ~pi792 & n10566;
  assign n10600 = ~n10598 & ~n10599;
  assign n10601 = ~pi647 & ~n10600;
  assign n10602 = ~n8334 & n10571;
  assign n10603 = n8334 & n10410;
  assign n10604 = ~n10602 & ~n10603;
  assign n10605 = pi647 & ~n10604;
  assign n10606 = ~pi1157 & ~n10605;
  assign n10607 = ~n10601 & n10606;
  assign n10608 = ~pi792 & ~n62987;
  assign n10609 = ~n10584 & ~n10594;
  assign n10610 = pi792 & ~n10609;
  assign n10611 = ~n10608 & ~n10610;
  assign n10612 = pi647 & n10611;
  assign n10613 = ~pi647 & n10410;
  assign n10614 = pi1157 & ~n10613;
  assign n10615 = ~n10612 & n10614;
  assign n10616 = ~pi630 & ~n10615;
  assign n10617 = ~n10607 & n10616;
  assign n10618 = pi647 & ~n10600;
  assign n10619 = ~pi647 & ~n10604;
  assign n10620 = pi1157 & ~n10619;
  assign n10621 = ~n10618 & n10620;
  assign n10622 = ~pi647 & n10611;
  assign n10623 = pi647 & n10410;
  assign n10624 = ~pi1157 & ~n10623;
  assign n10625 = ~n10622 & n10624;
  assign n10626 = pi630 & ~n10625;
  assign n10627 = ~n10621 & n10626;
  assign n10628 = ~n10617 & ~n10627;
  assign n10629 = pi787 & ~n10628;
  assign n10630 = ~pi787 & ~n10600;
  assign n10631 = ~n10629 & ~n10630;
  assign n10632 = ~pi644 & ~n10631;
  assign n10633 = ~pi787 & ~n10611;
  assign n10634 = ~n10615 & ~n10625;
  assign n10635 = pi787 & ~n10634;
  assign n10636 = ~n10633 & ~n10635;
  assign n10637 = pi644 & n10636;
  assign n10638 = ~pi715 & ~n10637;
  assign n10639 = ~n10632 & n10638;
  assign n10640 = n8376 & ~n10410;
  assign n10641 = ~n8376 & n10604;
  assign n10642 = ~n8376 & ~n10604;
  assign n10643 = n8376 & n10410;
  assign n10644 = ~n10642 & ~n10643;
  assign n10645 = ~n10640 & ~n10641;
  assign n10646 = ~pi644 & ~n62988;
  assign n10647 = pi644 & n10410;
  assign n10648 = pi715 & ~n10647;
  assign n10649 = ~n10646 & n10648;
  assign n10650 = ~pi1160 & ~n10649;
  assign n10651 = ~n10639 & n10650;
  assign n10652 = pi644 & ~n10631;
  assign n10653 = ~pi644 & n10636;
  assign n10654 = pi715 & ~n10653;
  assign n10655 = ~n10652 & n10654;
  assign n10656 = pi644 & ~n62988;
  assign n10657 = ~pi644 & n10410;
  assign n10658 = ~pi715 & ~n10657;
  assign n10659 = ~n10656 & n10658;
  assign n10660 = pi1160 & ~n10659;
  assign n10661 = ~n10655 & n10660;
  assign n10662 = pi790 & ~n10661;
  assign n10663 = pi790 & ~n10651;
  assign n10664 = ~n10661 & n10663;
  assign n10665 = ~n10651 & n10662;
  assign n10666 = ~pi790 & n10631;
  assign n10667 = n62455 & ~n10666;
  assign n10668 = ~n62989 & n10667;
  assign n10669 = ~pi143 & ~n62455;
  assign n10670 = ~pi832 & ~n10669;
  assign n10671 = ~n10668 & n10670;
  assign n10672 = ~pi143 & ~n2923;
  assign n10673 = n8334 & ~n10672;
  assign n10674 = ~n8418 & n10672;
  assign n10675 = ~pi774 & n7316;
  assign n10676 = ~n10672 & ~n10675;
  assign n10677 = ~n8420 & ~n10676;
  assign n10678 = ~pi785 & ~n10677;
  assign n10679 = ~n8425 & ~n10676;
  assign n10680 = pi1155 & ~n10679;
  assign n10681 = ~n8428 & n10677;
  assign n10682 = ~pi1155 & ~n10681;
  assign n10683 = ~n10680 & ~n10682;
  assign n10684 = pi785 & ~n10683;
  assign n10685 = ~n10678 & ~n10684;
  assign n10686 = ~pi781 & ~n10685;
  assign n10687 = ~n8435 & n10685;
  assign n10688 = pi1154 & ~n10687;
  assign n10689 = ~n8438 & n10685;
  assign n10690 = ~pi1154 & ~n10689;
  assign n10691 = ~n10688 & ~n10690;
  assign n10692 = pi781 & ~n10691;
  assign n10693 = ~n10686 & ~n10692;
  assign n10694 = ~pi789 & ~n10693;
  assign n10695 = pi619 & n10693;
  assign n10696 = ~pi619 & n10672;
  assign n10697 = pi1159 & ~n10696;
  assign n10698 = ~n10695 & n10697;
  assign n10699 = ~pi619 & n10693;
  assign n10700 = pi619 & n10672;
  assign n10701 = ~pi1159 & ~n10700;
  assign n10702 = ~n10699 & n10701;
  assign n10703 = ~n10698 & ~n10702;
  assign n10704 = pi789 & ~n10703;
  assign n10705 = ~n10694 & ~n10704;
  assign n10706 = n8418 & n10705;
  assign n10707 = pi626 & n10705;
  assign n10708 = ~pi626 & n10672;
  assign n10709 = pi1158 & ~n10708;
  assign n10710 = ~n10707 & n10709;
  assign n10711 = ~pi626 & n10705;
  assign n10712 = pi626 & n10672;
  assign n10713 = ~pi1158 & ~n10712;
  assign n10714 = ~n10711 & n10713;
  assign n10715 = ~n10710 & ~n10714;
  assign n10716 = ~n10674 & ~n10706;
  assign n10717 = pi788 & n62990;
  assign n10718 = ~pi788 & n10705;
  assign n10719 = ~pi788 & ~n10705;
  assign n10720 = pi788 & ~n62990;
  assign n10721 = ~n10719 & ~n10720;
  assign n10722 = ~n10717 & ~n10718;
  assign n10723 = ~n8334 & ~n62991;
  assign n10724 = ~n8334 & n62991;
  assign n10725 = n8334 & n10672;
  assign n10726 = ~n10724 & ~n10725;
  assign n10727 = ~n10673 & ~n10723;
  assign n10728 = ~n8413 & n62992;
  assign n10729 = pi687 & n7564;
  assign n10730 = ~n10672 & ~n10729;
  assign n10731 = ~pi778 & n10730;
  assign n10732 = ~pi625 & n10729;
  assign n10733 = ~n10730 & ~n10732;
  assign n10734 = pi1153 & ~n10733;
  assign n10735 = ~pi1153 & ~n10672;
  assign n10736 = ~n10732 & n10735;
  assign n10737 = ~n10734 & ~n10736;
  assign n10738 = pi778 & ~n10737;
  assign n10739 = ~n10731 & ~n10738;
  assign n10740 = ~n8490 & n10739;
  assign n10741 = ~n8492 & n10740;
  assign n10742 = ~n8494 & n10741;
  assign n10743 = ~n8496 & n10742;
  assign n10744 = ~n8508 & n10743;
  assign n10745 = pi647 & ~n10744;
  assign n10746 = ~pi647 & ~n10672;
  assign n10747 = ~n10745 & ~n10746;
  assign n10748 = n8373 & ~n10747;
  assign n10749 = ~pi647 & n10744;
  assign n10750 = pi647 & n10672;
  assign n10751 = ~pi1157 & ~n10750;
  assign n10752 = ~n10749 & n10751;
  assign n10753 = pi630 & n10752;
  assign n10754 = ~n10748 & ~n10753;
  assign n10755 = ~n10728 & n10754;
  assign n10756 = pi787 & ~n10755;
  assign n10757 = n8525 & n10742;
  assign n10758 = ~n8302 & n62990;
  assign n10759 = ~n10757 & ~n10758;
  assign n10760 = pi788 & ~n10759;
  assign n10761 = ~n7187 & ~n10730;
  assign n10762 = pi625 & n10761;
  assign n10763 = n10676 & ~n10761;
  assign n10764 = ~n10762 & ~n10763;
  assign n10765 = n10735 & ~n10764;
  assign n10766 = ~pi608 & ~n10734;
  assign n10767 = ~n10765 & n10766;
  assign n10768 = pi1153 & n10676;
  assign n10769 = ~n10762 & n10768;
  assign n10770 = pi608 & ~n10736;
  assign n10771 = ~n10769 & n10770;
  assign n10772 = ~n10767 & ~n10771;
  assign n10773 = pi778 & ~n10772;
  assign n10774 = ~pi778 & ~n10763;
  assign n10775 = ~n10773 & ~n10774;
  assign n10776 = ~pi609 & ~n10775;
  assign n10777 = pi609 & n10739;
  assign n10778 = ~pi1155 & ~n10777;
  assign n10779 = ~n10776 & n10778;
  assign n10780 = ~pi660 & ~n10680;
  assign n10781 = ~n10779 & n10780;
  assign n10782 = pi609 & ~n10775;
  assign n10783 = ~pi609 & n10739;
  assign n10784 = pi1155 & ~n10783;
  assign n10785 = ~n10782 & n10784;
  assign n10786 = pi660 & ~n10682;
  assign n10787 = ~n10785 & n10786;
  assign n10788 = ~n10781 & ~n10787;
  assign n10789 = pi785 & ~n10788;
  assign n10790 = ~pi785 & ~n10775;
  assign n10791 = ~n10789 & ~n10790;
  assign n10792 = ~pi618 & ~n10791;
  assign n10793 = pi618 & n10740;
  assign n10794 = ~pi1154 & ~n10793;
  assign n10795 = ~n10792 & n10794;
  assign n10796 = ~pi627 & ~n10688;
  assign n10797 = ~n10795 & n10796;
  assign n10798 = pi618 & ~n10791;
  assign n10799 = ~pi618 & n10740;
  assign n10800 = pi1154 & ~n10799;
  assign n10801 = ~n10798 & n10800;
  assign n10802 = pi627 & ~n10690;
  assign n10803 = ~n10801 & n10802;
  assign n10804 = ~n10797 & ~n10803;
  assign n10805 = pi781 & ~n10804;
  assign n10806 = ~pi781 & ~n10791;
  assign n10807 = ~n10805 & ~n10806;
  assign n10808 = pi619 & ~n10807;
  assign n10809 = ~pi619 & n10741;
  assign n10810 = pi1159 & ~n10809;
  assign n10811 = ~n10808 & n10810;
  assign n10812 = pi648 & ~n10702;
  assign n10813 = ~n10811 & n10812;
  assign n10814 = ~pi619 & ~n10807;
  assign n10815 = pi619 & n10741;
  assign n10816 = ~pi1159 & ~n10815;
  assign n10817 = ~n10814 & n10816;
  assign n10818 = ~pi648 & ~n10698;
  assign n10819 = ~n10817 & n10818;
  assign n10820 = pi789 & ~n10819;
  assign n10821 = pi789 & ~n10813;
  assign n10822 = ~n10819 & n10821;
  assign n10823 = ~n10813 & n10820;
  assign n10824 = ~pi789 & n10807;
  assign n10825 = n62894 & ~n10824;
  assign n10826 = ~n62993 & n10825;
  assign n10827 = ~n10760 & ~n10826;
  assign n10828 = ~pi628 & n10827;
  assign n10829 = pi628 & ~n62991;
  assign n10830 = ~pi1156 & ~n10829;
  assign n10831 = ~n10828 & n10830;
  assign n10832 = n8606 & n10743;
  assign n10833 = ~pi629 & ~n10832;
  assign n10834 = ~n10831 & n10833;
  assign n10835 = pi628 & n10827;
  assign n10836 = ~pi628 & ~n62991;
  assign n10837 = pi1156 & ~n10836;
  assign n10838 = ~n10835 & n10837;
  assign n10839 = n8615 & n10743;
  assign n10840 = pi629 & ~n10839;
  assign n10841 = ~n10838 & n10840;
  assign n10842 = pi792 & ~n10841;
  assign n10843 = ~pi628 & ~n10827;
  assign n10844 = pi628 & n62991;
  assign n10845 = ~pi1156 & ~n10844;
  assign n10846 = ~n10843 & n10845;
  assign n10847 = ~n8605 & n10743;
  assign n10848 = pi1156 & ~n10847;
  assign n10849 = ~pi629 & ~n10848;
  assign n10850 = ~n10846 & n10849;
  assign n10851 = pi628 & ~n10827;
  assign n10852 = ~pi628 & n62991;
  assign n10853 = pi1156 & ~n10852;
  assign n10854 = ~n10851 & n10853;
  assign n10855 = ~n8614 & n10743;
  assign n10856 = ~pi1156 & ~n10855;
  assign n10857 = pi629 & ~n10856;
  assign n10858 = ~n10854 & n10857;
  assign n10859 = ~n10850 & ~n10858;
  assign n10860 = pi792 & ~n10859;
  assign n10861 = ~n10834 & n10842;
  assign n10862 = ~pi792 & ~n10827;
  assign n10863 = ~n8651 & ~n10862;
  assign n10864 = ~n62994 & n10863;
  assign n10865 = ~n62994 & ~n10862;
  assign n10866 = ~pi647 & ~n10865;
  assign n10867 = pi647 & ~n62992;
  assign n10868 = ~pi1157 & ~n10867;
  assign n10869 = ~n10866 & n10868;
  assign n10870 = pi647 & n10744;
  assign n10871 = ~pi647 & n10672;
  assign n10872 = pi1157 & ~n10871;
  assign n10873 = pi1157 & ~n10747;
  assign n10874 = ~n10870 & n10872;
  assign n10875 = ~pi630 & ~n62995;
  assign n10876 = ~n10869 & n10875;
  assign n10877 = pi647 & ~n10865;
  assign n10878 = ~pi647 & ~n62992;
  assign n10879 = pi1157 & ~n10878;
  assign n10880 = ~n10877 & n10879;
  assign n10881 = pi630 & ~n10752;
  assign n10882 = ~n10880 & n10881;
  assign n10883 = ~n10876 & ~n10882;
  assign n10884 = pi787 & ~n10883;
  assign n10885 = ~pi787 & ~n10865;
  assign n10886 = ~n10884 & ~n10885;
  assign n10887 = ~n10756 & ~n10864;
  assign n10888 = pi644 & ~n62996;
  assign n10889 = ~pi787 & ~n10744;
  assign n10890 = ~n10752 & ~n62995;
  assign n10891 = pi787 & ~n10890;
  assign n10892 = ~n10889 & ~n10891;
  assign n10893 = ~pi644 & n10892;
  assign n10894 = pi715 & ~n10893;
  assign n10895 = ~n10888 & n10894;
  assign n10896 = ~n8685 & ~n10672;
  assign n10897 = ~n8376 & n10723;
  assign n10898 = n8376 & ~n10672;
  assign n10899 = ~n8376 & n62992;
  assign n10900 = ~n10898 & ~n10899;
  assign n10901 = ~n10896 & ~n10897;
  assign n10902 = pi644 & n62997;
  assign n10903 = ~pi644 & n10672;
  assign n10904 = ~pi715 & ~n10903;
  assign n10905 = ~n10902 & n10904;
  assign n10906 = pi1160 & ~n10905;
  assign n10907 = ~n10895 & n10906;
  assign n10908 = ~pi644 & ~n62996;
  assign n10909 = pi644 & n10892;
  assign n10910 = ~pi715 & ~n10909;
  assign n10911 = ~n10908 & n10910;
  assign n10912 = ~pi644 & n62997;
  assign n10913 = pi644 & n10672;
  assign n10914 = pi715 & ~n10913;
  assign n10915 = ~n10912 & n10914;
  assign n10916 = ~pi1160 & ~n10915;
  assign n10917 = ~n10911 & n10916;
  assign n10918 = ~n10907 & ~n10917;
  assign n10919 = pi790 & ~n10918;
  assign n10920 = ~pi790 & ~n62996;
  assign n10921 = pi832 & ~n10920;
  assign n10922 = ~n10919 & n10921;
  assign po300 = ~n10671 & ~n10922;
  assign n10924 = pi144 & ~n62765;
  assign n10925 = ~pi758 & ~n7143;
  assign n10926 = pi758 & ~n62801;
  assign n10927 = ~n10925 & ~n10926;
  assign n10928 = pi39 & ~n10927;
  assign n10929 = pi758 & n62793;
  assign n10930 = ~pi758 & ~n62781;
  assign n10931 = ~pi39 & ~n10930;
  assign n10932 = ~n10929 & n10931;
  assign n10933 = ~n10928 & ~n10932;
  assign n10934 = pi144 & ~n10933;
  assign n10935 = ~pi144 & pi758;
  assign n10936 = n7351 & n10935;
  assign n10937 = ~n10934 & ~n10936;
  assign n10938 = ~pi38 & ~n10937;
  assign n10939 = pi758 & n7187;
  assign n10940 = n7357 & ~n10939;
  assign n10941 = ~pi144 & ~n7357;
  assign n10942 = pi38 & ~n10941;
  assign n10943 = pi38 & ~n10940;
  assign n10944 = ~n10941 & n10943;
  assign n10945 = ~n10940 & n10942;
  assign n10946 = ~n10938 & ~n62998;
  assign n10947 = ~pi736 & n10946;
  assign n10948 = pi144 & n62821;
  assign n10949 = ~pi144 & ~n7632;
  assign n10950 = ~pi758 & ~n10949;
  assign n10951 = ~n10948 & n10950;
  assign n10952 = ~pi144 & ~n7709;
  assign n10953 = pi144 & ~n62851;
  assign n10954 = pi758 & ~n10953;
  assign n10955 = ~n10952 & n10954;
  assign n10956 = pi39 & ~n10955;
  assign n10957 = ~n10951 & n10956;
  assign n10958 = ~pi144 & ~n7855;
  assign n10959 = pi144 & ~n7832;
  assign n10960 = ~pi758 & ~n10959;
  assign n10961 = ~pi758 & ~n10958;
  assign n10962 = ~n10959 & n10961;
  assign n10963 = ~n10958 & n10960;
  assign n10964 = pi144 & n7861;
  assign n10965 = ~pi144 & n7868;
  assign n10966 = pi758 & ~n10965;
  assign n10967 = ~n10964 & n10966;
  assign n10968 = ~pi39 & ~n10967;
  assign n10969 = pi144 & ~n7861;
  assign n10970 = ~pi144 & ~n7868;
  assign n10971 = pi758 & ~n10970;
  assign n10972 = ~n10969 & n10971;
  assign n10973 = pi144 & n7832;
  assign n10974 = ~pi144 & n7855;
  assign n10975 = ~pi758 & ~n10974;
  assign n10976 = ~n10973 & n10975;
  assign n10977 = ~n10972 & ~n10976;
  assign n10978 = ~pi39 & ~n10977;
  assign n10979 = ~n62999 & n10968;
  assign n10980 = ~pi38 & ~n63000;
  assign n10981 = ~n10957 & n10980;
  assign n10982 = pi736 & ~n10357;
  assign n10983 = ~n62998 & n10982;
  assign n10984 = ~n10981 & n10983;
  assign n10985 = n62765 & ~n10984;
  assign n10986 = ~n10947 & n10985;
  assign n10987 = ~n10924 & ~n10986;
  assign n10988 = ~pi625 & n10987;
  assign n10989 = n62765 & ~n10946;
  assign n10990 = ~n10924 & ~n10989;
  assign n10991 = pi625 & n10990;
  assign n10992 = ~pi1153 & ~n10991;
  assign n10993 = ~n10988 & n10992;
  assign n10994 = pi736 & n62765;
  assign n10995 = n7357 & ~n7563;
  assign n10996 = n7356 & n7952;
  assign n10997 = pi38 & ~n63001;
  assign n10998 = ~n10941 & n10997;
  assign n10999 = pi144 & ~n8009;
  assign n11000 = ~pi144 & ~n62874;
  assign n11001 = ~pi38 & ~n11000;
  assign n11002 = ~n10999 & n11001;
  assign n11003 = ~n10998 & ~n11002;
  assign n11004 = n10994 & ~n11003;
  assign n11005 = pi144 & ~n8098;
  assign n11006 = ~n10994 & n11005;
  assign n11007 = ~n10994 & ~n11005;
  assign n11008 = n10994 & ~n10998;
  assign n11009 = ~n11002 & n11008;
  assign n11010 = ~n11007 & ~n11009;
  assign n11011 = ~n11004 & ~n11006;
  assign n11012 = pi625 & ~n63002;
  assign n11013 = ~pi625 & ~n11005;
  assign n11014 = pi1153 & ~n11013;
  assign n11015 = ~n11012 & n11014;
  assign n11016 = ~pi608 & ~n11015;
  assign n11017 = ~n10993 & n11016;
  assign n11018 = pi625 & n10987;
  assign n11019 = ~pi625 & n10990;
  assign n11020 = pi1153 & ~n11019;
  assign n11021 = ~n11018 & n11020;
  assign n11022 = ~pi625 & ~n63002;
  assign n11023 = pi625 & ~n11005;
  assign n11024 = ~pi1153 & ~n11023;
  assign n11025 = ~n11022 & n11024;
  assign n11026 = pi608 & ~n11025;
  assign n11027 = ~n11021 & n11026;
  assign n11028 = ~n11017 & ~n11027;
  assign n11029 = pi778 & ~n11028;
  assign n11030 = ~pi778 & n10987;
  assign n11031 = ~n11029 & ~n11030;
  assign n11032 = ~pi609 & ~n11031;
  assign n11033 = ~pi778 & n63002;
  assign n11034 = ~n11015 & ~n11025;
  assign n11035 = pi778 & ~n11034;
  assign n11036 = ~n11033 & ~n11035;
  assign n11037 = pi609 & n11036;
  assign n11038 = ~pi1155 & ~n11037;
  assign n11039 = ~n11032 & n11038;
  assign n11040 = ~n8135 & ~n10990;
  assign n11041 = n8135 & n11005;
  assign n11042 = n8135 & ~n11005;
  assign n11043 = ~n8135 & n10990;
  assign n11044 = ~n11042 & ~n11043;
  assign n11045 = ~n11040 & ~n11041;
  assign n11046 = pi609 & ~n63003;
  assign n11047 = ~pi609 & ~n11005;
  assign n11048 = pi1155 & ~n11047;
  assign n11049 = ~n11046 & n11048;
  assign n11050 = ~pi660 & ~n11049;
  assign n11051 = ~n11039 & n11050;
  assign n11052 = pi609 & ~n11031;
  assign n11053 = ~pi609 & n11036;
  assign n11054 = pi1155 & ~n11053;
  assign n11055 = ~n11052 & n11054;
  assign n11056 = ~pi609 & ~n63003;
  assign n11057 = pi609 & ~n11005;
  assign n11058 = ~pi1155 & ~n11057;
  assign n11059 = ~n11056 & n11058;
  assign n11060 = pi660 & ~n11059;
  assign n11061 = ~n11055 & n11060;
  assign n11062 = ~n11051 & ~n11061;
  assign n11063 = pi785 & ~n11062;
  assign n11064 = ~pi785 & ~n11031;
  assign n11065 = ~n11063 & ~n11064;
  assign n11066 = ~pi618 & ~n11065;
  assign n11067 = n62880 & ~n11005;
  assign n11068 = ~n62880 & n11036;
  assign n11069 = ~n62880 & ~n11036;
  assign n11070 = n62880 & n11005;
  assign n11071 = ~n11069 & ~n11070;
  assign n11072 = ~n11067 & ~n11068;
  assign n11073 = pi618 & n63004;
  assign n11074 = ~pi1154 & ~n11073;
  assign n11075 = ~n11066 & n11074;
  assign n11076 = ~pi785 & n63003;
  assign n11077 = ~n11049 & ~n11059;
  assign n11078 = pi785 & ~n11077;
  assign n11079 = ~n11076 & ~n11078;
  assign n11080 = pi618 & n11079;
  assign n11081 = ~pi618 & ~n11005;
  assign n11082 = pi1154 & ~n11081;
  assign n11083 = ~n11080 & n11082;
  assign n11084 = ~pi627 & ~n11083;
  assign n11085 = ~n11075 & n11084;
  assign n11086 = pi618 & ~n11065;
  assign n11087 = ~pi618 & n63004;
  assign n11088 = pi1154 & ~n11087;
  assign n11089 = ~n11086 & n11088;
  assign n11090 = ~pi618 & n11079;
  assign n11091 = pi618 & ~n11005;
  assign n11092 = ~pi1154 & ~n11091;
  assign n11093 = ~n11090 & n11092;
  assign n11094 = pi627 & ~n11093;
  assign n11095 = ~n11089 & n11094;
  assign n11096 = ~n11085 & ~n11095;
  assign n11097 = pi781 & ~n11096;
  assign n11098 = ~pi781 & ~n11065;
  assign n11099 = ~n11097 & ~n11098;
  assign n11100 = ~pi619 & ~n11099;
  assign n11101 = ~n62882 & ~n63004;
  assign n11102 = n62882 & n11005;
  assign n11103 = n62882 & ~n11005;
  assign n11104 = ~n62882 & n63004;
  assign n11105 = ~n11103 & ~n11104;
  assign n11106 = ~n11101 & ~n11102;
  assign n11107 = pi619 & ~n63005;
  assign n11108 = ~pi1159 & ~n11107;
  assign n11109 = ~n11100 & n11108;
  assign n11110 = ~pi781 & ~n11079;
  assign n11111 = ~n11083 & ~n11093;
  assign n11112 = pi781 & ~n11111;
  assign n11113 = ~n11110 & ~n11112;
  assign n11114 = pi619 & n11113;
  assign n11115 = ~pi619 & ~n11005;
  assign n11116 = pi1159 & ~n11115;
  assign n11117 = ~n11114 & n11116;
  assign n11118 = ~pi648 & ~n11117;
  assign n11119 = ~n11109 & n11118;
  assign n11120 = pi619 & ~n11099;
  assign n11121 = ~pi619 & ~n63005;
  assign n11122 = pi1159 & ~n11121;
  assign n11123 = ~n11120 & n11122;
  assign n11124 = ~pi619 & n11113;
  assign n11125 = pi619 & ~n11005;
  assign n11126 = ~pi1159 & ~n11125;
  assign n11127 = ~n11124 & n11126;
  assign n11128 = pi648 & ~n11127;
  assign n11129 = ~n11123 & n11128;
  assign n11130 = ~n11119 & ~n11129;
  assign n11131 = pi789 & ~n11130;
  assign n11132 = ~pi789 & ~n11099;
  assign n11133 = ~n11131 & ~n11132;
  assign n11134 = ~pi788 & n11133;
  assign n11135 = ~pi626 & n11133;
  assign n11136 = n8257 & ~n11005;
  assign n11137 = ~n8257 & ~n63005;
  assign n11138 = ~n8257 & n63005;
  assign n11139 = n8257 & n11005;
  assign n11140 = ~n11138 & ~n11139;
  assign n11141 = ~n11136 & ~n11137;
  assign n11142 = pi626 & ~n63006;
  assign n11143 = ~pi641 & ~n11142;
  assign n11144 = ~n11135 & n11143;
  assign n11145 = ~pi789 & ~n11113;
  assign n11146 = ~n11117 & ~n11127;
  assign n11147 = pi789 & ~n11146;
  assign n11148 = ~n11145 & ~n11147;
  assign n11149 = ~pi626 & n11148;
  assign n11150 = pi626 & ~n11005;
  assign n11151 = ~pi1158 & ~n11150;
  assign n11152 = ~n11149 & n11151;
  assign n11153 = ~n8267 & ~n11152;
  assign n11154 = ~n11144 & ~n11153;
  assign n11155 = pi626 & n11133;
  assign n11156 = ~pi626 & ~n63006;
  assign n11157 = pi641 & ~n11156;
  assign n11158 = ~n11155 & n11157;
  assign n11159 = pi626 & n11148;
  assign n11160 = ~pi626 & ~n11005;
  assign n11161 = pi1158 & ~n11160;
  assign n11162 = ~n11159 & n11161;
  assign n11163 = ~n8282 & ~n11162;
  assign n11164 = ~n11158 & ~n11163;
  assign n11165 = ~n11154 & ~n11164;
  assign n11166 = pi788 & ~n11165;
  assign n11167 = ~n11134 & ~n11166;
  assign n11168 = ~pi628 & n11167;
  assign n11169 = ~n11152 & ~n11162;
  assign n11170 = pi788 & ~n11169;
  assign n11171 = ~pi788 & ~n11148;
  assign n11172 = ~n11170 & ~n11171;
  assign n11173 = pi628 & n11172;
  assign n11174 = ~pi1156 & ~n11173;
  assign n11175 = ~n11168 & n11174;
  assign n11176 = ~n8303 & ~n63006;
  assign n11177 = n8303 & n11005;
  assign n11178 = n8303 & ~n11005;
  assign n11179 = ~n8303 & n63006;
  assign n11180 = ~n11178 & ~n11179;
  assign n11181 = ~n11176 & ~n11177;
  assign n11182 = pi628 & ~n63007;
  assign n11183 = ~pi628 & ~n11005;
  assign n11184 = pi1156 & ~n11183;
  assign n11185 = ~n11182 & n11184;
  assign n11186 = ~pi629 & ~n11185;
  assign n11187 = ~n11175 & n11186;
  assign n11188 = pi628 & n11167;
  assign n11189 = ~pi628 & n11172;
  assign n11190 = pi1156 & ~n11189;
  assign n11191 = ~n11188 & n11190;
  assign n11192 = ~pi628 & ~n63007;
  assign n11193 = pi628 & ~n11005;
  assign n11194 = ~pi1156 & ~n11193;
  assign n11195 = ~n11192 & n11194;
  assign n11196 = pi629 & ~n11195;
  assign n11197 = ~n11191 & n11196;
  assign n11198 = ~n11187 & ~n11197;
  assign n11199 = pi792 & ~n11198;
  assign n11200 = ~pi792 & n11167;
  assign n11201 = ~n11199 & ~n11200;
  assign n11202 = ~pi647 & ~n11201;
  assign n11203 = ~n8334 & ~n11172;
  assign n11204 = n8334 & n11005;
  assign n11205 = ~n11203 & ~n11204;
  assign n11206 = pi647 & n11205;
  assign n11207 = ~pi1157 & ~n11206;
  assign n11208 = ~n11202 & n11207;
  assign n11209 = ~pi792 & n63007;
  assign n11210 = ~n11185 & ~n11195;
  assign n11211 = pi792 & ~n11210;
  assign n11212 = ~n11209 & ~n11211;
  assign n11213 = pi647 & n11212;
  assign n11214 = ~pi647 & ~n11005;
  assign n11215 = pi1157 & ~n11214;
  assign n11216 = ~n11213 & n11215;
  assign n11217 = ~pi630 & ~n11216;
  assign n11218 = ~n11208 & n11217;
  assign n11219 = pi647 & ~n11201;
  assign n11220 = ~pi647 & n11205;
  assign n11221 = pi1157 & ~n11220;
  assign n11222 = ~n11219 & n11221;
  assign n11223 = ~pi647 & n11212;
  assign n11224 = pi647 & ~n11005;
  assign n11225 = ~pi1157 & ~n11224;
  assign n11226 = ~n11223 & n11225;
  assign n11227 = pi630 & ~n11226;
  assign n11228 = ~n11222 & n11227;
  assign n11229 = ~n11218 & ~n11228;
  assign n11230 = pi787 & ~n11229;
  assign n11231 = ~pi787 & ~n11201;
  assign n11232 = ~n11230 & ~n11231;
  assign n11233 = ~pi644 & ~n11232;
  assign n11234 = ~pi787 & ~n11212;
  assign n11235 = ~n11216 & ~n11226;
  assign n11236 = pi787 & ~n11235;
  assign n11237 = ~n11234 & ~n11236;
  assign n11238 = pi644 & n11237;
  assign n11239 = ~pi715 & ~n11238;
  assign n11240 = ~n11233 & n11239;
  assign n11241 = n8376 & ~n11005;
  assign n11242 = ~n8376 & n11205;
  assign n11243 = ~n8376 & ~n11205;
  assign n11244 = n8376 & n11005;
  assign n11245 = ~n11243 & ~n11244;
  assign n11246 = ~n11241 & ~n11242;
  assign n11247 = ~pi644 & n63008;
  assign n11248 = pi644 & ~n11005;
  assign n11249 = pi715 & ~n11248;
  assign n11250 = ~n11247 & n11249;
  assign n11251 = ~pi1160 & ~n11250;
  assign n11252 = ~n11240 & n11251;
  assign n11253 = pi644 & ~n11232;
  assign n11254 = ~pi644 & n11237;
  assign n11255 = pi715 & ~n11254;
  assign n11256 = ~n11253 & n11255;
  assign n11257 = pi644 & n63008;
  assign n11258 = ~pi644 & ~n11005;
  assign n11259 = ~pi715 & ~n11258;
  assign n11260 = ~n11257 & n11259;
  assign n11261 = pi1160 & ~n11260;
  assign n11262 = ~n11256 & n11261;
  assign n11263 = pi790 & ~n11262;
  assign n11264 = pi790 & ~n11252;
  assign n11265 = ~n11262 & n11264;
  assign n11266 = ~n11252 & n11263;
  assign n11267 = ~pi790 & n11232;
  assign n11268 = n3475 & ~n11267;
  assign n11269 = ~n63009 & n11268;
  assign n11270 = ~pi144 & ~n3475;
  assign n11271 = ~pi57 & ~n11270;
  assign n11272 = ~n11269 & n11271;
  assign n11273 = pi57 & pi144;
  assign n11274 = ~pi832 & ~n11273;
  assign n11275 = ~n11272 & n11274;
  assign n11276 = pi144 & ~n2923;
  assign n11277 = pi736 & n7564;
  assign n11278 = ~n11276 & ~n11277;
  assign n11279 = ~pi778 & n11278;
  assign n11280 = pi625 & n11277;
  assign n11281 = ~n11278 & ~n11280;
  assign n11282 = ~pi1153 & ~n11281;
  assign n11283 = pi1153 & ~n11276;
  assign n11284 = ~n11280 & n11283;
  assign n11285 = ~n11282 & ~n11284;
  assign n11286 = pi778 & ~n11285;
  assign n11287 = ~n11279 & ~n11286;
  assign n11288 = ~n62880 & n11287;
  assign n11289 = ~n62882 & n11288;
  assign n11290 = ~n8257 & n11289;
  assign n11291 = ~n8303 & n11290;
  assign n11292 = n10207 & n11287;
  assign n11293 = ~pi628 & n63010;
  assign n11294 = pi629 & ~n11293;
  assign n11295 = pi609 & pi1155;
  assign n11296 = ~pi609 & ~pi1155;
  assign n11297 = pi785 & ~n11296;
  assign n11298 = pi785 & ~n11295;
  assign n11299 = ~n11296 & n11298;
  assign n11300 = ~n11295 & n11297;
  assign n11301 = pi758 & n7316;
  assign n11302 = ~n63011 & n11301;
  assign n11303 = ~pi619 & pi1159;
  assign n11304 = pi619 & ~pi1159;
  assign n11305 = ~n11303 & ~n11304;
  assign n11306 = pi789 & ~n11305;
  assign n11307 = pi618 & pi1154;
  assign n11308 = ~pi618 & ~pi1154;
  assign n11309 = pi781 & ~n11308;
  assign n11310 = pi781 & ~n11307;
  assign n11311 = ~n11308 & n11310;
  assign n11312 = ~n11307 & n11309;
  assign n11313 = ~n8135 & ~n63012;
  assign n11314 = ~n8135 & ~n11306;
  assign n11315 = ~n63012 & n11314;
  assign n11316 = ~n11306 & n11313;
  assign n11317 = n11302 & n63013;
  assign n11318 = ~n8595 & n11317;
  assign n11319 = pi628 & ~n11318;
  assign n11320 = ~n11294 & ~n11319;
  assign n11321 = ~pi1156 & ~n11320;
  assign n11322 = pi628 & n63010;
  assign n11323 = ~pi628 & ~n11318;
  assign n11324 = pi629 & ~n11323;
  assign n11325 = pi1156 & ~n11324;
  assign n11326 = ~n11322 & n11325;
  assign n11327 = ~n11321 & ~n11326;
  assign n11328 = pi792 & ~n11276;
  assign n11329 = ~n11276 & ~n11327;
  assign n11330 = pi792 & n11329;
  assign n11331 = ~n11327 & n11328;
  assign n11332 = pi736 & n7565;
  assign n11333 = ~n7187 & n11277;
  assign n11334 = ~n7187 & n11280;
  assign n11335 = pi625 & n63015;
  assign n11336 = ~n11276 & ~n11301;
  assign n11337 = ~n63015 & n11336;
  assign n11338 = ~n63016 & ~n11337;
  assign n11339 = ~pi1153 & ~n11338;
  assign n11340 = ~pi608 & ~n11284;
  assign n11341 = ~n11339 & n11340;
  assign n11342 = pi1153 & n11336;
  assign n11343 = n11283 & ~n11301;
  assign n11344 = ~n63016 & n63017;
  assign n11345 = pi608 & ~n11282;
  assign n11346 = ~n11344 & n11345;
  assign n11347 = ~n11341 & ~n11346;
  assign n11348 = pi778 & ~n11347;
  assign n11349 = ~pi778 & ~n11337;
  assign n11350 = ~n11348 & ~n11349;
  assign n11351 = ~pi609 & ~n11350;
  assign n11352 = pi609 & n11287;
  assign n11353 = ~pi1155 & ~n11352;
  assign n11354 = ~n11351 & n11353;
  assign n11355 = n8136 & n11301;
  assign n11356 = pi1155 & ~n11276;
  assign n11357 = ~n11355 & n11356;
  assign n11358 = ~pi660 & ~n11357;
  assign n11359 = ~n11354 & n11358;
  assign n11360 = pi609 & ~n11350;
  assign n11361 = ~pi609 & n11287;
  assign n11362 = pi1155 & ~n11361;
  assign n11363 = ~n11360 & n11362;
  assign n11364 = n8148 & n11301;
  assign n11365 = ~pi1155 & ~n11276;
  assign n11366 = ~n11364 & n11365;
  assign n11367 = pi660 & ~n11366;
  assign n11368 = ~n11363 & n11367;
  assign n11369 = ~n11359 & ~n11368;
  assign n11370 = pi785 & ~n11369;
  assign n11371 = ~pi785 & ~n11350;
  assign n11372 = ~pi618 & n8209;
  assign n11373 = pi627 & n11307;
  assign n11374 = pi618 & n8210;
  assign n11375 = pi781 & ~n63018;
  assign n11376 = ~n11372 & n11375;
  assign n11377 = ~n11371 & ~n11376;
  assign n11378 = ~n11370 & n11377;
  assign n11379 = pi618 & n8209;
  assign n11380 = ~pi618 & pi627;
  assign n11381 = pi1154 & n11380;
  assign n11382 = ~pi618 & n8210;
  assign n11383 = ~n11379 & ~n63019;
  assign n11384 = ~n11288 & ~n11383;
  assign n11385 = ~n8208 & ~n11302;
  assign n11386 = pi618 & ~n8135;
  assign n11387 = n8207 & ~n11386;
  assign n11388 = ~pi618 & ~n8135;
  assign n11389 = n8206 & ~n11388;
  assign n11390 = ~n11387 & ~n11389;
  assign n11391 = ~n11385 & n11390;
  assign n11392 = ~n11384 & n11391;
  assign n11393 = pi781 & ~n11276;
  assign n11394 = ~n11392 & n11393;
  assign n11395 = ~n11370 & ~n11371;
  assign n11396 = ~pi618 & ~n11395;
  assign n11397 = ~n11276 & ~n11288;
  assign n11398 = pi618 & ~n11397;
  assign n11399 = ~pi1154 & ~n11398;
  assign n11400 = ~n11396 & n11399;
  assign n11401 = n11302 & n11386;
  assign n11402 = pi1154 & ~n11276;
  assign n11403 = ~n11401 & n11402;
  assign n11404 = ~pi627 & ~n11403;
  assign n11405 = ~n11400 & n11404;
  assign n11406 = pi618 & ~n11395;
  assign n11407 = ~pi618 & ~n11397;
  assign n11408 = pi1154 & ~n11407;
  assign n11409 = ~n11406 & n11408;
  assign n11410 = n11302 & n11388;
  assign n11411 = ~pi1154 & ~n11276;
  assign n11412 = ~n11410 & n11411;
  assign n11413 = pi627 & ~n11412;
  assign n11414 = ~n11409 & n11413;
  assign n11415 = ~n11405 & ~n11414;
  assign n11416 = pi781 & ~n11415;
  assign n11417 = ~pi781 & ~n11395;
  assign n11418 = ~n11416 & ~n11417;
  assign n11419 = ~n11378 & ~n11394;
  assign n11420 = ~pi619 & ~pi648;
  assign n11421 = ~pi1159 & n11420;
  assign n11422 = pi619 & pi648;
  assign n11423 = pi1159 & n11422;
  assign n11424 = n62884 & n11305;
  assign n11425 = pi619 & ~pi648;
  assign n11426 = ~pi648 & n11304;
  assign n11427 = ~pi1159 & n11425;
  assign n11428 = ~pi619 & pi648;
  assign n11429 = pi648 & n11303;
  assign n11430 = pi1159 & n11428;
  assign n11431 = ~n63022 & ~n63023;
  assign n11432 = n62884 & n11431;
  assign n11433 = ~n11421 & ~n11423;
  assign n11434 = pi789 & ~n63021;
  assign n11435 = n63020 & ~n11434;
  assign n11436 = n11302 & n11313;
  assign n11437 = n11302 & ~n63012;
  assign n11438 = ~pi619 & ~n8135;
  assign n11439 = n11437 & n11438;
  assign n11440 = ~pi619 & n11436;
  assign n11441 = pi648 & ~n63024;
  assign n11442 = pi619 & ~n11289;
  assign n11443 = ~n11441 & ~n11442;
  assign n11444 = ~pi1159 & ~n11443;
  assign n11445 = ~pi619 & ~n11289;
  assign n11446 = pi648 & ~n11445;
  assign n11447 = pi619 & ~n8135;
  assign n11448 = n11437 & n11447;
  assign n11449 = pi619 & n11436;
  assign n11450 = pi1159 & ~n63025;
  assign n11451 = ~n11446 & n11450;
  assign n11452 = ~n11444 & ~n11451;
  assign n11453 = pi789 & ~n11276;
  assign n11454 = ~n11452 & n11453;
  assign n11455 = n62894 & ~n11454;
  assign n11456 = ~pi619 & ~n63020;
  assign n11457 = ~n11276 & ~n11289;
  assign n11458 = pi619 & ~n11457;
  assign n11459 = ~pi1159 & ~n11458;
  assign n11460 = ~n11456 & n11459;
  assign n11461 = pi1159 & ~n11276;
  assign n11462 = ~n63025 & n11461;
  assign n11463 = ~pi648 & ~n11462;
  assign n11464 = ~n11460 & n11463;
  assign n11465 = pi619 & ~n63020;
  assign n11466 = ~pi619 & ~n11457;
  assign n11467 = pi1159 & ~n11466;
  assign n11468 = ~n11465 & n11467;
  assign n11469 = ~pi1159 & ~n11276;
  assign n11470 = ~n63024 & n11469;
  assign n11471 = pi648 & ~n11470;
  assign n11472 = ~n11468 & n11471;
  assign n11473 = pi789 & ~n11472;
  assign n11474 = pi789 & ~n11464;
  assign n11475 = ~n11472 & n11474;
  assign n11476 = ~n11464 & n11473;
  assign n11477 = ~pi789 & n63020;
  assign n11478 = n62894 & ~n11477;
  assign n11479 = ~n63026 & n11478;
  assign n11480 = ~n11435 & n11455;
  assign n11481 = n8333 & n8500;
  assign n11482 = ~pi628 & ~pi629;
  assign n11483 = ~pi1156 & n11482;
  assign n11484 = ~pi629 & n8501;
  assign n11485 = pi628 & pi629;
  assign n11486 = pi1156 & n11485;
  assign n11487 = pi629 & n8502;
  assign n11488 = pi792 & ~n63029;
  assign n11489 = ~n63028 & n11488;
  assign n11490 = pi792 & ~n63028;
  assign n11491 = ~n63029 & n11490;
  assign n11492 = pi792 & ~n11481;
  assign n11493 = n8257 & ~n11276;
  assign n11494 = ~n11457 & ~n11493;
  assign n11495 = ~n11276 & ~n11290;
  assign n11496 = n8417 & n63031;
  assign n11497 = pi626 & n11317;
  assign n11498 = ~n11276 & ~n11497;
  assign n11499 = pi1158 & ~n11498;
  assign n11500 = ~pi641 & ~n11499;
  assign n11501 = ~n11496 & n11500;
  assign n11502 = n8416 & n63031;
  assign n11503 = ~pi626 & n11317;
  assign n11504 = ~n11276 & ~n11503;
  assign n11505 = ~pi1158 & ~n11504;
  assign n11506 = pi641 & ~n11505;
  assign n11507 = ~n11502 & n11506;
  assign n11508 = pi788 & ~n11507;
  assign n11509 = pi788 & ~n11501;
  assign n11510 = ~n11507 & n11509;
  assign n11511 = ~n11501 & n11508;
  assign n11512 = ~n63030 & ~n63032;
  assign n11513 = ~n63027 & n11512;
  assign n11514 = ~n63014 & ~n11513;
  assign n11515 = ~n63027 & ~n63032;
  assign n11516 = ~n63014 & ~n11515;
  assign n11517 = ~n11329 & n63030;
  assign n11518 = ~n8651 & ~n11517;
  assign n11519 = ~n11516 & n11518;
  assign n11520 = ~n8651 & ~n11514;
  assign n11521 = ~n62892 & n63010;
  assign n11522 = ~pi630 & ~n11521;
  assign n11523 = pi647 & ~n11522;
  assign n11524 = ~n8334 & n11318;
  assign n11525 = pi630 & n11524;
  assign n11526 = pi1157 & ~n11525;
  assign n11527 = ~n11523 & n11526;
  assign n11528 = pi630 & ~n11521;
  assign n11529 = ~pi647 & ~n11528;
  assign n11530 = ~pi630 & n11524;
  assign n11531 = ~pi1157 & ~n11530;
  assign n11532 = pi647 & ~n11530;
  assign n11533 = ~n11528 & ~n11532;
  assign n11534 = ~pi1157 & ~n11533;
  assign n11535 = ~n11529 & n11531;
  assign n11536 = ~n11527 & ~n63034;
  assign n11537 = pi787 & ~n11276;
  assign n11538 = ~n11536 & n11537;
  assign n11539 = ~pi715 & ~pi1160;
  assign n11540 = ~pi644 & ~n11539;
  assign n11541 = pi715 & pi1160;
  assign n11542 = pi644 & ~n11541;
  assign n11543 = ~pi644 & n11539;
  assign n11544 = pi644 & n11541;
  assign n11545 = ~n11543 & ~n11544;
  assign n11546 = ~n11540 & ~n11542;
  assign n11547 = pi790 & n63035;
  assign n11548 = ~n11538 & ~n11547;
  assign n11549 = ~n63033 & n11548;
  assign n11550 = ~pi644 & ~n11541;
  assign n11551 = pi644 & ~n11539;
  assign n11552 = pi644 & n11539;
  assign n11553 = ~pi644 & n11541;
  assign n11554 = ~n11552 & ~n11553;
  assign n11555 = ~n11550 & ~n11551;
  assign n11556 = ~n10298 & ~n63036;
  assign n11557 = n11521 & n11556;
  assign n11558 = ~n8595 & n8685;
  assign n11559 = ~n8376 & n11524;
  assign n11560 = n11317 & n11558;
  assign n11561 = ~pi1160 & n63037;
  assign n11562 = ~n11276 & ~n11561;
  assign n11563 = n11540 & ~n11562;
  assign n11564 = pi1160 & n63037;
  assign n11565 = ~n11276 & ~n11564;
  assign n11566 = n11542 & ~n11565;
  assign n11567 = ~n11563 & ~n11566;
  assign n11568 = ~n11557 & n11567;
  assign n11569 = pi790 & ~n11568;
  assign n11570 = pi832 & ~n11569;
  assign n11571 = ~n63033 & ~n11538;
  assign n11572 = pi644 & n11571;
  assign n11573 = ~n10298 & n11521;
  assign n11574 = ~n11276 & ~n11573;
  assign n11575 = ~pi644 & ~n11574;
  assign n11576 = pi715 & ~n11575;
  assign n11577 = ~n11572 & n11576;
  assign n11578 = pi644 & n63037;
  assign n11579 = ~pi715 & ~n11276;
  assign n11580 = ~n11578 & n11579;
  assign n11581 = pi1160 & ~n11580;
  assign n11582 = ~n11577 & n11581;
  assign n11583 = ~pi644 & n11571;
  assign n11584 = pi644 & ~n11574;
  assign n11585 = ~pi715 & ~n11584;
  assign n11586 = ~n11583 & n11585;
  assign n11587 = ~pi644 & n63037;
  assign n11588 = pi715 & ~n11276;
  assign n11589 = ~n11587 & n11588;
  assign n11590 = ~pi1160 & ~n11589;
  assign n11591 = ~n11586 & n11590;
  assign n11592 = ~n11582 & ~n11591;
  assign n11593 = pi790 & ~n11592;
  assign n11594 = ~pi790 & n11571;
  assign n11595 = pi832 & ~n11594;
  assign n11596 = ~n11593 & n11595;
  assign n11597 = ~n11549 & n11570;
  assign po301 = ~n11275 & ~n63038;
  assign n11599 = ~pi145 & ~n8098;
  assign n11600 = n8257 & ~n11599;
  assign n11601 = ~pi698 & n62765;
  assign n11602 = n11599 & ~n11601;
  assign n11603 = pi145 & n62874;
  assign n11604 = ~pi38 & ~n11603;
  assign n11605 = n62765 & ~n11604;
  assign n11606 = ~pi145 & n8009;
  assign n11607 = ~n11605 & ~n11606;
  assign n11608 = ~pi145 & ~n7357;
  assign n11609 = n8085 & ~n11608;
  assign n11610 = ~pi698 & ~n11609;
  assign n11611 = ~n11607 & n11610;
  assign n11612 = ~n11602 & ~n11611;
  assign n11613 = ~pi778 & n11612;
  assign n11614 = pi625 & ~n11612;
  assign n11615 = ~pi625 & n11599;
  assign n11616 = pi1153 & ~n11615;
  assign n11617 = ~n11614 & n11616;
  assign n11618 = ~pi625 & ~n11612;
  assign n11619 = pi625 & n11599;
  assign n11620 = ~pi1153 & ~n11619;
  assign n11621 = ~n11618 & n11620;
  assign n11622 = ~n11617 & ~n11621;
  assign n11623 = pi778 & ~n11622;
  assign n11624 = ~n11613 & ~n11623;
  assign n11625 = ~n62880 & ~n11624;
  assign n11626 = n62880 & ~n11599;
  assign n11627 = ~n62880 & n11624;
  assign n11628 = n62880 & n11599;
  assign n11629 = ~n11627 & ~n11628;
  assign n11630 = ~n11625 & ~n11626;
  assign n11631 = ~n62882 & ~n63039;
  assign n11632 = n62882 & n11599;
  assign n11633 = n62882 & ~n11599;
  assign n11634 = ~n62882 & n63039;
  assign n11635 = ~n11633 & ~n11634;
  assign n11636 = ~n11631 & ~n11632;
  assign n11637 = ~n8257 & ~n63040;
  assign n11638 = ~n8257 & n63040;
  assign n11639 = n8257 & n11599;
  assign n11640 = ~n11638 & ~n11639;
  assign n11641 = ~n11600 & ~n11637;
  assign n11642 = ~n8303 & ~n63041;
  assign n11643 = n8303 & n11599;
  assign n11644 = ~n11642 & ~n11643;
  assign n11645 = ~pi792 & n11644;
  assign n11646 = pi628 & ~n11644;
  assign n11647 = ~pi628 & n11599;
  assign n11648 = pi1156 & ~n11647;
  assign n11649 = ~n11646 & n11648;
  assign n11650 = ~pi628 & ~n11644;
  assign n11651 = pi628 & n11599;
  assign n11652 = ~pi1156 & ~n11651;
  assign n11653 = ~n11650 & n11652;
  assign n11654 = ~n11649 & ~n11653;
  assign n11655 = pi792 & ~n11654;
  assign n11656 = ~n11645 & ~n11655;
  assign n11657 = pi647 & n11656;
  assign n11658 = ~pi647 & n11599;
  assign n11659 = pi1157 & ~n11658;
  assign n11660 = pi647 & ~n11656;
  assign n11661 = ~pi647 & ~n11599;
  assign n11662 = ~n11660 & ~n11661;
  assign n11663 = pi1157 & ~n11662;
  assign n11664 = ~n11657 & n11659;
  assign n11665 = ~pi647 & n11656;
  assign n11666 = pi647 & n11599;
  assign n11667 = ~pi1157 & ~n11666;
  assign n11668 = ~n11665 & n11667;
  assign n11669 = ~pi647 & ~n11656;
  assign n11670 = pi647 & ~n11599;
  assign n11671 = ~n11669 & ~n11670;
  assign n11672 = ~pi1157 & n11671;
  assign n11673 = pi1157 & n11662;
  assign n11674 = ~n11672 & ~n11673;
  assign n11675 = ~n63042 & ~n11668;
  assign n11676 = pi787 & n63043;
  assign n11677 = ~pi787 & ~n11656;
  assign n11678 = pi787 & ~n63043;
  assign n11679 = ~pi787 & n11656;
  assign n11680 = ~n11678 & ~n11679;
  assign n11681 = ~n11676 & ~n11677;
  assign n11682 = ~pi644 & ~n63044;
  assign n11683 = pi715 & ~n11682;
  assign n11684 = pi145 & ~n62765;
  assign n11685 = ~pi767 & n7359;
  assign n11686 = ~n11608 & ~n11685;
  assign n11687 = pi38 & ~n11686;
  assign n11688 = ~pi145 & n62802;
  assign n11689 = pi145 & ~n7351;
  assign n11690 = ~pi767 & ~n11689;
  assign n11691 = ~n11688 & n11690;
  assign n11692 = ~pi145 & pi767;
  assign n11693 = ~n62792 & n11692;
  assign n11694 = pi767 & ~n62792;
  assign n11695 = ~pi767 & ~n11688;
  assign n11696 = ~n11694 & ~n11695;
  assign n11697 = ~pi145 & ~n11696;
  assign n11698 = n7351 & n11695;
  assign n11699 = ~n11697 & ~n11698;
  assign n11700 = ~pi145 & ~n62792;
  assign n11701 = pi767 & ~n11700;
  assign n11702 = ~pi145 & ~pi767;
  assign n11703 = n62802 & n11702;
  assign n11704 = ~n11689 & ~n11703;
  assign n11705 = ~n11701 & n11704;
  assign n11706 = ~n11691 & ~n11693;
  assign n11707 = ~pi38 & ~n63045;
  assign n11708 = ~pi38 & n63045;
  assign n11709 = pi38 & ~n11608;
  assign n11710 = ~n11685 & n11709;
  assign n11711 = ~n11708 & ~n11710;
  assign n11712 = ~n11687 & ~n11707;
  assign n11713 = n62765 & ~n63046;
  assign n11714 = ~n11684 & ~n11713;
  assign n11715 = ~n8135 & ~n11714;
  assign n11716 = n8135 & ~n11599;
  assign n11717 = ~n11715 & ~n11716;
  assign n11718 = ~pi785 & ~n11717;
  assign n11719 = ~n8136 & ~n11599;
  assign n11720 = pi609 & n11715;
  assign n11721 = ~n11719 & ~n11720;
  assign n11722 = pi1155 & ~n11721;
  assign n11723 = ~n8148 & ~n11599;
  assign n11724 = ~pi609 & n11715;
  assign n11725 = ~n11723 & ~n11724;
  assign n11726 = ~pi1155 & ~n11725;
  assign n11727 = ~n11722 & ~n11726;
  assign n11728 = pi785 & ~n11727;
  assign n11729 = ~n11718 & ~n11728;
  assign n11730 = ~pi781 & ~n11729;
  assign n11731 = pi618 & n11729;
  assign n11732 = ~pi618 & n11599;
  assign n11733 = pi1154 & ~n11732;
  assign n11734 = ~n11731 & n11733;
  assign n11735 = ~pi618 & n11729;
  assign n11736 = pi618 & n11599;
  assign n11737 = ~pi1154 & ~n11736;
  assign n11738 = ~n11735 & n11737;
  assign n11739 = ~n11734 & ~n11738;
  assign n11740 = pi781 & ~n11739;
  assign n11741 = ~n11730 & ~n11740;
  assign n11742 = ~pi619 & ~n11741;
  assign n11743 = pi619 & ~n11599;
  assign n11744 = ~pi1159 & ~n11743;
  assign n11745 = ~n11742 & n11744;
  assign n11746 = pi619 & ~n11741;
  assign n11747 = ~pi619 & ~n11599;
  assign n11748 = pi1159 & ~n11747;
  assign n11749 = ~n11746 & n11748;
  assign n11750 = pi619 & n11741;
  assign n11751 = ~pi619 & n11599;
  assign n11752 = pi1159 & ~n11751;
  assign n11753 = ~n11750 & n11752;
  assign n11754 = ~pi619 & n11741;
  assign n11755 = pi619 & n11599;
  assign n11756 = ~pi1159 & ~n11755;
  assign n11757 = ~n11754 & n11756;
  assign n11758 = ~n11753 & ~n11757;
  assign n11759 = ~n11745 & ~n11749;
  assign n11760 = pi789 & n63047;
  assign n11761 = ~pi789 & n11741;
  assign n11762 = ~pi789 & ~n11741;
  assign n11763 = pi789 & ~n63047;
  assign n11764 = ~n11762 & ~n11763;
  assign n11765 = ~n11760 & ~n11761;
  assign n11766 = n8418 & n63048;
  assign n11767 = ~n8418 & n11599;
  assign n11768 = pi626 & n63048;
  assign n11769 = ~pi626 & n11599;
  assign n11770 = pi1158 & ~n11769;
  assign n11771 = ~n11768 & n11770;
  assign n11772 = ~pi626 & n63048;
  assign n11773 = pi626 & n11599;
  assign n11774 = ~pi1158 & ~n11773;
  assign n11775 = ~n11772 & n11774;
  assign n11776 = ~n11771 & ~n11775;
  assign n11777 = ~n11766 & ~n11767;
  assign n11778 = pi788 & n63049;
  assign n11779 = ~pi788 & n63048;
  assign n11780 = ~pi788 & ~n63048;
  assign n11781 = pi788 & ~n63049;
  assign n11782 = ~n11780 & ~n11781;
  assign n11783 = ~n11778 & ~n11779;
  assign n11784 = ~n8334 & n63050;
  assign n11785 = n8334 & n11599;
  assign n11786 = ~n11784 & ~n11785;
  assign n11787 = ~n8376 & ~n11786;
  assign n11788 = n8376 & n11599;
  assign n11789 = n8376 & ~n11599;
  assign n11790 = ~n8376 & n11786;
  assign n11791 = ~n11789 & ~n11790;
  assign n11792 = ~n11787 & ~n11788;
  assign n11793 = pi644 & n63051;
  assign n11794 = ~pi644 & n11599;
  assign n11795 = ~pi715 & ~n11794;
  assign n11796 = ~n11793 & n11795;
  assign n11797 = pi1160 & ~n11796;
  assign n11798 = ~n11683 & n11797;
  assign n11799 = pi628 & ~pi629;
  assign n11800 = ~pi1156 & ~n11799;
  assign n11801 = ~pi628 & pi629;
  assign n11802 = pi1156 & ~n11801;
  assign n11803 = pi1156 & n11801;
  assign n11804 = ~pi1156 & n11799;
  assign n11805 = ~n11803 & ~n11804;
  assign n11806 = ~n11800 & ~n11802;
  assign n11807 = ~n63050 & ~n63052;
  assign n11808 = ~pi629 & n11649;
  assign n11809 = pi629 & n11653;
  assign n11810 = ~n11808 & ~n11809;
  assign n11811 = ~n11807 & n11810;
  assign n11812 = pi792 & ~n11811;
  assign n11813 = n8525 & ~n63041;
  assign n11814 = ~n8302 & n63049;
  assign n11815 = ~n11813 & ~n11814;
  assign n11816 = pi788 & ~n11815;
  assign n11817 = pi698 & n63046;
  assign n11818 = ~pi145 & ~n62821;
  assign n11819 = pi145 & n7632;
  assign n11820 = pi767 & ~n11819;
  assign n11821 = ~n11818 & n11820;
  assign n11822 = pi145 & n7709;
  assign n11823 = ~pi145 & n62851;
  assign n11824 = ~pi767 & ~n11823;
  assign n11825 = ~n11822 & n11824;
  assign n11826 = pi39 & ~n11825;
  assign n11827 = ~n11821 & n11826;
  assign n11828 = pi145 & n7855;
  assign n11829 = ~pi145 & n7832;
  assign n11830 = pi767 & ~n11829;
  assign n11831 = ~n11828 & n11830;
  assign n11832 = ~pi145 & ~n7861;
  assign n11833 = pi145 & ~n7868;
  assign n11834 = ~pi767 & ~n11833;
  assign n11835 = ~n11832 & n11834;
  assign n11836 = ~pi39 & ~n11835;
  assign n11837 = pi145 & ~n7855;
  assign n11838 = ~pi145 & ~n7832;
  assign n11839 = pi767 & ~n11838;
  assign n11840 = pi767 & ~n11837;
  assign n11841 = ~n11838 & n11840;
  assign n11842 = ~n11837 & n11839;
  assign n11843 = ~pi145 & n7861;
  assign n11844 = pi145 & n7868;
  assign n11845 = ~pi767 & ~n11844;
  assign n11846 = ~n11843 & n11845;
  assign n11847 = ~n63053 & ~n11846;
  assign n11848 = ~pi39 & ~n11847;
  assign n11849 = ~n11831 & n11836;
  assign n11850 = ~pi38 & ~n63054;
  assign n11851 = ~n11827 & n11850;
  assign n11852 = ~pi767 & ~n7744;
  assign n11853 = n10350 & ~n11852;
  assign n11854 = ~pi145 & ~n11853;
  assign n11855 = ~pi767 & n7316;
  assign n11856 = ~n7565 & ~n11855;
  assign n11857 = pi145 & ~n11856;
  assign n11858 = n7356 & n11857;
  assign n11859 = pi38 & ~n11858;
  assign n11860 = ~n11854 & n11859;
  assign n11861 = ~pi698 & ~n11860;
  assign n11862 = ~n11851 & n11861;
  assign n11863 = n62765 & ~n11862;
  assign n11864 = ~n11817 & n11863;
  assign n11865 = ~n11684 & ~n11864;
  assign n11866 = ~pi625 & n11865;
  assign n11867 = pi625 & n11714;
  assign n11868 = ~pi1153 & ~n11867;
  assign n11869 = ~n11866 & n11868;
  assign n11870 = ~pi608 & ~n11617;
  assign n11871 = ~n11869 & n11870;
  assign n11872 = pi625 & n11865;
  assign n11873 = ~pi625 & n11714;
  assign n11874 = pi1153 & ~n11873;
  assign n11875 = ~n11872 & n11874;
  assign n11876 = pi608 & ~n11621;
  assign n11877 = ~n11875 & n11876;
  assign n11878 = ~n11871 & ~n11877;
  assign n11879 = pi778 & ~n11878;
  assign n11880 = ~pi778 & n11865;
  assign n11881 = ~n11879 & ~n11880;
  assign n11882 = ~pi609 & ~n11881;
  assign n11883 = pi609 & n11624;
  assign n11884 = ~pi1155 & ~n11883;
  assign n11885 = ~n11882 & n11884;
  assign n11886 = ~pi660 & ~n11722;
  assign n11887 = ~n11885 & n11886;
  assign n11888 = pi609 & ~n11881;
  assign n11889 = ~pi609 & n11624;
  assign n11890 = pi1155 & ~n11889;
  assign n11891 = ~n11888 & n11890;
  assign n11892 = pi660 & ~n11726;
  assign n11893 = ~n11891 & n11892;
  assign n11894 = ~n11887 & ~n11893;
  assign n11895 = pi785 & ~n11894;
  assign n11896 = ~pi785 & ~n11881;
  assign n11897 = ~n11895 & ~n11896;
  assign n11898 = pi618 & ~n11897;
  assign n11899 = ~pi618 & ~n63039;
  assign n11900 = pi1154 & ~n11899;
  assign n11901 = ~n11898 & n11900;
  assign n11902 = pi627 & ~n11738;
  assign n11903 = ~n11901 & n11902;
  assign n11904 = ~pi618 & ~n11897;
  assign n11905 = pi618 & ~n63039;
  assign n11906 = ~pi1154 & ~n11905;
  assign n11907 = ~n11904 & n11906;
  assign n11908 = ~pi627 & ~n11734;
  assign n11909 = ~n11907 & n11908;
  assign n11910 = pi781 & ~n11909;
  assign n11911 = ~n11903 & n11910;
  assign n11912 = ~n11431 & ~n63040;
  assign n11913 = ~n62884 & ~n63047;
  assign n11914 = ~n11912 & ~n11913;
  assign n11915 = pi789 & ~n11914;
  assign n11916 = ~pi781 & n11897;
  assign n11917 = ~n11915 & ~n11916;
  assign n11918 = ~n11911 & n11917;
  assign n11919 = n11434 & n11914;
  assign n11920 = ~n11918 & ~n11919;
  assign n11921 = ~n11903 & ~n11909;
  assign n11922 = pi781 & ~n11921;
  assign n11923 = ~pi781 & ~n11897;
  assign n11924 = ~n11922 & ~n11923;
  assign n11925 = ~pi619 & ~n11924;
  assign n11926 = pi619 & n63040;
  assign n11927 = ~pi1159 & ~n11926;
  assign n11928 = ~n11925 & n11927;
  assign n11929 = ~pi648 & ~n11753;
  assign n11930 = ~n11928 & n11929;
  assign n11931 = pi619 & ~n11924;
  assign n11932 = ~pi619 & n63040;
  assign n11933 = pi1159 & ~n11932;
  assign n11934 = ~n11931 & n11933;
  assign n11935 = pi648 & ~n11757;
  assign n11936 = ~n11934 & n11935;
  assign n11937 = pi789 & ~n11936;
  assign n11938 = pi789 & ~n11930;
  assign n11939 = ~n11936 & n11938;
  assign n11940 = ~n11930 & n11937;
  assign n11941 = ~pi789 & n11924;
  assign n11942 = n62894 & ~n11941;
  assign n11943 = ~n63055 & n11942;
  assign n11944 = n62894 & ~n11920;
  assign n11945 = ~n63030 & ~n63056;
  assign n11946 = ~n63030 & ~n11816;
  assign n11947 = ~n63056 & n11946;
  assign n11948 = ~n11816 & n11945;
  assign n11949 = ~n11812 & ~n63057;
  assign n11950 = ~n8651 & ~n11949;
  assign n11951 = ~n8413 & n11786;
  assign n11952 = n8373 & ~n11662;
  assign n11953 = ~pi630 & n63042;
  assign n11954 = n8374 & ~n11671;
  assign n11955 = pi630 & n11668;
  assign n11956 = ~n63058 & ~n63059;
  assign n11957 = ~n11951 & n11956;
  assign n11958 = pi787 & ~n11957;
  assign n11959 = ~n11950 & ~n11958;
  assign n11960 = ~pi644 & n11959;
  assign n11961 = pi644 & ~n63044;
  assign n11962 = ~pi715 & ~n11961;
  assign n11963 = ~n11960 & n11962;
  assign n11964 = ~pi644 & n63051;
  assign n11965 = pi644 & n11599;
  assign n11966 = pi715 & ~n11965;
  assign n11967 = ~n11964 & n11966;
  assign n11968 = ~pi1160 & ~n11967;
  assign n11969 = ~n11963 & n11968;
  assign n11970 = ~n11798 & ~n11969;
  assign n11971 = pi790 & ~n11970;
  assign n11972 = pi644 & n11797;
  assign n11973 = pi790 & ~n11972;
  assign n11974 = n11959 & ~n11973;
  assign n11975 = ~n11971 & ~n11974;
  assign n11976 = n62455 & ~n11975;
  assign n11977 = ~pi145 & ~n62455;
  assign n11978 = ~pi832 & ~n11977;
  assign n11979 = ~n11976 & n11978;
  assign n11980 = ~pi145 & ~n2923;
  assign n11981 = ~n11855 & ~n11980;
  assign n11982 = ~n8420 & ~n11981;
  assign n11983 = ~pi785 & ~n11982;
  assign n11984 = ~n8425 & ~n11981;
  assign n11985 = pi1155 & ~n11984;
  assign n11986 = ~n8428 & n11982;
  assign n11987 = ~pi1155 & ~n11986;
  assign n11988 = ~n11985 & ~n11987;
  assign n11989 = pi785 & ~n11988;
  assign n11990 = ~n11983 & ~n11989;
  assign n11991 = ~pi781 & ~n11990;
  assign n11992 = ~n8435 & n11990;
  assign n11993 = pi1154 & ~n11992;
  assign n11994 = ~n8438 & n11990;
  assign n11995 = ~pi1154 & ~n11994;
  assign n11996 = ~n11993 & ~n11995;
  assign n11997 = pi781 & ~n11996;
  assign n11998 = ~n11991 & ~n11997;
  assign n11999 = ~pi619 & ~n11998;
  assign n12000 = pi619 & ~n11980;
  assign n12001 = ~pi1159 & ~n12000;
  assign n12002 = ~n11999 & n12001;
  assign n12003 = pi619 & ~n11998;
  assign n12004 = ~pi619 & ~n11980;
  assign n12005 = pi1159 & ~n12004;
  assign n12006 = ~n12003 & n12005;
  assign n12007 = pi619 & n11998;
  assign n12008 = ~pi619 & n11980;
  assign n12009 = pi1159 & ~n12008;
  assign n12010 = ~n12007 & n12009;
  assign n12011 = ~pi619 & n11998;
  assign n12012 = pi619 & n11980;
  assign n12013 = ~pi1159 & ~n12012;
  assign n12014 = ~n12011 & n12013;
  assign n12015 = ~n12010 & ~n12014;
  assign n12016 = ~n12002 & ~n12006;
  assign n12017 = pi789 & n63060;
  assign n12018 = ~pi789 & n11998;
  assign n12019 = ~pi789 & ~n11998;
  assign n12020 = pi789 & ~n63060;
  assign n12021 = ~n12019 & ~n12020;
  assign n12022 = ~n12017 & ~n12018;
  assign n12023 = n8418 & n63061;
  assign n12024 = ~n8418 & n11980;
  assign n12025 = pi626 & n63061;
  assign n12026 = ~pi626 & n11980;
  assign n12027 = pi1158 & ~n12026;
  assign n12028 = ~n12025 & n12027;
  assign n12029 = ~pi626 & n63061;
  assign n12030 = pi626 & n11980;
  assign n12031 = ~pi1158 & ~n12030;
  assign n12032 = ~n12029 & n12031;
  assign n12033 = ~n12028 & ~n12032;
  assign n12034 = ~n12023 & ~n12024;
  assign n12035 = pi788 & n63062;
  assign n12036 = ~pi788 & n63061;
  assign n12037 = ~pi788 & ~n63061;
  assign n12038 = pi788 & ~n63062;
  assign n12039 = ~n12037 & ~n12038;
  assign n12040 = ~n12035 & ~n12036;
  assign n12041 = ~n8334 & n63063;
  assign n12042 = n8334 & n11980;
  assign n12043 = ~n8413 & ~n12042;
  assign n12044 = ~n12041 & ~n12042;
  assign n12045 = ~n8413 & n12044;
  assign n12046 = ~n12041 & n12043;
  assign n12047 = ~pi698 & n7564;
  assign n12048 = ~n11980 & ~n12047;
  assign n12049 = ~pi778 & n12048;
  assign n12050 = ~pi625 & n12047;
  assign n12051 = ~n12048 & ~n12050;
  assign n12052 = pi1153 & ~n12051;
  assign n12053 = ~pi1153 & ~n11980;
  assign n12054 = ~n12050 & n12053;
  assign n12055 = ~n12052 & ~n12054;
  assign n12056 = pi778 & ~n12055;
  assign n12057 = ~n12049 & ~n12056;
  assign n12058 = ~n8490 & n12057;
  assign n12059 = ~n8492 & n12058;
  assign n12060 = ~n8494 & n12059;
  assign n12061 = ~n8496 & n12060;
  assign n12062 = ~n8508 & n12061;
  assign n12063 = pi647 & ~n12062;
  assign n12064 = ~pi647 & ~n11980;
  assign n12065 = ~n12063 & ~n12064;
  assign n12066 = n8373 & ~n12065;
  assign n12067 = ~pi647 & n12062;
  assign n12068 = pi647 & n11980;
  assign n12069 = ~pi1157 & ~n12068;
  assign n12070 = ~n12067 & n12069;
  assign n12071 = pi630 & n12070;
  assign n12072 = ~n12066 & ~n12071;
  assign n12073 = ~n63064 & n12072;
  assign n12074 = pi787 & ~n12073;
  assign n12075 = n8525 & n12060;
  assign n12076 = ~n8302 & n63062;
  assign n12077 = ~n12075 & ~n12076;
  assign n12078 = pi788 & ~n12077;
  assign n12079 = ~n7187 & ~n12048;
  assign n12080 = pi625 & n12079;
  assign n12081 = n11981 & ~n12079;
  assign n12082 = ~n12080 & ~n12081;
  assign n12083 = n12053 & ~n12082;
  assign n12084 = ~pi608 & ~n12052;
  assign n12085 = ~n12083 & n12084;
  assign n12086 = pi1153 & n11981;
  assign n12087 = ~n12080 & n12086;
  assign n12088 = pi608 & ~n12054;
  assign n12089 = ~n12087 & n12088;
  assign n12090 = ~n12085 & ~n12089;
  assign n12091 = pi778 & ~n12090;
  assign n12092 = ~pi778 & ~n12081;
  assign n12093 = ~n12091 & ~n12092;
  assign n12094 = ~pi609 & ~n12093;
  assign n12095 = pi609 & n12057;
  assign n12096 = ~pi1155 & ~n12095;
  assign n12097 = ~n12094 & n12096;
  assign n12098 = ~pi660 & ~n11985;
  assign n12099 = ~n12097 & n12098;
  assign n12100 = pi609 & ~n12093;
  assign n12101 = ~pi609 & n12057;
  assign n12102 = pi1155 & ~n12101;
  assign n12103 = ~n12100 & n12102;
  assign n12104 = pi660 & ~n11987;
  assign n12105 = ~n12103 & n12104;
  assign n12106 = ~n12099 & ~n12105;
  assign n12107 = pi785 & ~n12106;
  assign n12108 = ~pi785 & ~n12093;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = pi618 & ~n12109;
  assign n12111 = ~pi618 & n12058;
  assign n12112 = pi1154 & ~n12111;
  assign n12113 = ~n12110 & n12112;
  assign n12114 = pi627 & ~n11995;
  assign n12115 = ~n12113 & n12114;
  assign n12116 = ~pi618 & ~n12109;
  assign n12117 = pi618 & n12058;
  assign n12118 = ~pi1154 & ~n12117;
  assign n12119 = ~n12116 & n12118;
  assign n12120 = ~pi627 & ~n11993;
  assign n12121 = ~n12119 & n12120;
  assign n12122 = pi781 & ~n12121;
  assign n12123 = ~n12115 & n12122;
  assign n12124 = ~n11431 & ~n12059;
  assign n12125 = ~n62884 & ~n63060;
  assign n12126 = ~n12124 & ~n12125;
  assign n12127 = pi789 & ~n12126;
  assign n12128 = ~pi781 & n12109;
  assign n12129 = ~n12127 & ~n12128;
  assign n12130 = ~n12123 & n12129;
  assign n12131 = n11434 & n12126;
  assign n12132 = ~n12130 & ~n12131;
  assign n12133 = ~n12115 & ~n12121;
  assign n12134 = pi781 & ~n12133;
  assign n12135 = ~pi781 & ~n12109;
  assign n12136 = ~n12134 & ~n12135;
  assign n12137 = ~pi619 & ~n12136;
  assign n12138 = pi619 & n12059;
  assign n12139 = ~pi1159 & ~n12138;
  assign n12140 = ~n12137 & n12139;
  assign n12141 = ~pi648 & ~n12010;
  assign n12142 = ~n12140 & n12141;
  assign n12143 = pi619 & ~n12136;
  assign n12144 = ~pi619 & n12059;
  assign n12145 = pi1159 & ~n12144;
  assign n12146 = ~n12143 & n12145;
  assign n12147 = pi648 & ~n12014;
  assign n12148 = ~n12146 & n12147;
  assign n12149 = pi789 & ~n12148;
  assign n12150 = pi789 & ~n12142;
  assign n12151 = ~n12148 & n12150;
  assign n12152 = ~n12142 & n12149;
  assign n12153 = ~pi789 & n12136;
  assign n12154 = n62894 & ~n12153;
  assign n12155 = ~n63065 & n12154;
  assign n12156 = n62894 & ~n12132;
  assign n12157 = ~n12078 & ~n63066;
  assign n12158 = ~n63030 & ~n12157;
  assign n12159 = n8498 & n63063;
  assign n12160 = n8615 & n12061;
  assign n12161 = pi629 & ~n12160;
  assign n12162 = ~n12159 & n12161;
  assign n12163 = n8499 & n63063;
  assign n12164 = n8606 & n12061;
  assign n12165 = ~pi629 & ~n12164;
  assign n12166 = ~n12163 & n12165;
  assign n12167 = pi792 & ~n12166;
  assign n12168 = pi792 & ~n12162;
  assign n12169 = ~n12166 & n12168;
  assign n12170 = ~n12163 & ~n12164;
  assign n12171 = ~pi629 & ~n12170;
  assign n12172 = ~n12159 & ~n12160;
  assign n12173 = pi629 & ~n12172;
  assign n12174 = ~n12171 & ~n12173;
  assign n12175 = pi792 & ~n12174;
  assign n12176 = ~n12162 & n12167;
  assign n12177 = ~n8651 & ~n63067;
  assign n12178 = ~n12158 & n12177;
  assign n12179 = ~n12074 & ~n12178;
  assign n12180 = pi644 & n12179;
  assign n12181 = ~pi787 & ~n12062;
  assign n12182 = pi1157 & ~n12065;
  assign n12183 = ~n12070 & ~n12182;
  assign n12184 = pi787 & ~n12183;
  assign n12185 = ~n12181 & ~n12184;
  assign n12186 = ~pi644 & n12185;
  assign n12187 = pi715 & ~n12186;
  assign n12188 = ~n12180 & n12187;
  assign n12189 = ~n8685 & n11980;
  assign n12190 = ~n8376 & n12041;
  assign n12191 = ~n8376 & ~n12044;
  assign n12192 = n8376 & n11980;
  assign n12193 = ~n12191 & ~n12192;
  assign n12194 = ~n12189 & ~n12190;
  assign n12195 = pi644 & ~n63068;
  assign n12196 = ~pi644 & n11980;
  assign n12197 = ~pi715 & ~n12196;
  assign n12198 = ~n12195 & n12197;
  assign n12199 = pi1160 & ~n12198;
  assign n12200 = ~n12188 & n12199;
  assign n12201 = ~pi644 & n12179;
  assign n12202 = pi644 & n12185;
  assign n12203 = ~pi715 & ~n12202;
  assign n12204 = ~n12201 & n12203;
  assign n12205 = ~pi644 & ~n63068;
  assign n12206 = pi644 & n11980;
  assign n12207 = pi715 & ~n12206;
  assign n12208 = ~n12205 & n12207;
  assign n12209 = ~pi1160 & ~n12208;
  assign n12210 = ~n12204 & n12209;
  assign n12211 = ~n12200 & ~n12210;
  assign n12212 = pi790 & ~n12211;
  assign n12213 = ~pi790 & n12179;
  assign n12214 = pi832 & ~n12213;
  assign n12215 = ~n12212 & n12214;
  assign po302 = ~n11979 & ~n12215;
  assign n12217 = ~pi173 & ~n8098;
  assign n12218 = n8257 & ~n12217;
  assign n12219 = ~pi723 & n62765;
  assign n12220 = n12217 & ~n12219;
  assign n12221 = pi173 & n62874;
  assign n12222 = ~pi38 & ~n12221;
  assign n12223 = n62765 & ~n12222;
  assign n12224 = ~pi173 & n8009;
  assign n12225 = ~n12223 & ~n12224;
  assign n12226 = ~pi173 & ~n7357;
  assign n12227 = n8085 & ~n12226;
  assign n12228 = ~pi723 & ~n12227;
  assign n12229 = ~n12225 & n12228;
  assign n12230 = ~n12220 & ~n12229;
  assign n12231 = ~pi778 & n12230;
  assign n12232 = pi625 & ~n12230;
  assign n12233 = ~pi625 & n12217;
  assign n12234 = pi1153 & ~n12233;
  assign n12235 = ~n12232 & n12234;
  assign n12236 = ~pi625 & ~n12230;
  assign n12237 = pi625 & n12217;
  assign n12238 = ~pi1153 & ~n12237;
  assign n12239 = ~n12236 & n12238;
  assign n12240 = ~n12235 & ~n12239;
  assign n12241 = pi778 & ~n12240;
  assign n12242 = ~n12231 & ~n12241;
  assign n12243 = ~n62880 & ~n12242;
  assign n12244 = n62880 & ~n12217;
  assign n12245 = ~n62880 & n12242;
  assign n12246 = n62880 & n12217;
  assign n12247 = ~n12245 & ~n12246;
  assign n12248 = ~n12243 & ~n12244;
  assign n12249 = ~n62882 & ~n63069;
  assign n12250 = n62882 & n12217;
  assign n12251 = n62882 & ~n12217;
  assign n12252 = ~n62882 & n63069;
  assign n12253 = ~n12251 & ~n12252;
  assign n12254 = ~n12249 & ~n12250;
  assign n12255 = ~n8257 & ~n63070;
  assign n12256 = ~n8257 & n63070;
  assign n12257 = n8257 & n12217;
  assign n12258 = ~n12256 & ~n12257;
  assign n12259 = ~n12218 & ~n12255;
  assign n12260 = ~n8303 & ~n63071;
  assign n12261 = n8303 & n12217;
  assign n12262 = ~n12260 & ~n12261;
  assign n12263 = ~pi792 & n12262;
  assign n12264 = pi628 & ~n12262;
  assign n12265 = ~pi628 & n12217;
  assign n12266 = pi1156 & ~n12265;
  assign n12267 = ~n12264 & n12266;
  assign n12268 = ~pi628 & ~n12262;
  assign n12269 = pi628 & n12217;
  assign n12270 = ~pi1156 & ~n12269;
  assign n12271 = ~n12268 & n12270;
  assign n12272 = ~n12267 & ~n12271;
  assign n12273 = pi792 & ~n12272;
  assign n12274 = ~n12263 & ~n12273;
  assign n12275 = pi647 & n12274;
  assign n12276 = ~pi647 & n12217;
  assign n12277 = pi1157 & ~n12276;
  assign n12278 = pi647 & ~n12274;
  assign n12279 = ~pi647 & ~n12217;
  assign n12280 = ~n12278 & ~n12279;
  assign n12281 = pi1157 & ~n12280;
  assign n12282 = ~n12275 & n12277;
  assign n12283 = ~pi647 & n12274;
  assign n12284 = pi647 & n12217;
  assign n12285 = ~pi1157 & ~n12284;
  assign n12286 = ~n12283 & n12285;
  assign n12287 = ~pi647 & ~n12274;
  assign n12288 = pi647 & ~n12217;
  assign n12289 = ~n12287 & ~n12288;
  assign n12290 = ~pi1157 & n12289;
  assign n12291 = pi1157 & n12280;
  assign n12292 = ~n12290 & ~n12291;
  assign n12293 = ~n63072 & ~n12286;
  assign n12294 = pi787 & n63073;
  assign n12295 = ~pi787 & ~n12274;
  assign n12296 = pi787 & ~n63073;
  assign n12297 = ~pi787 & n12274;
  assign n12298 = ~n12296 & ~n12297;
  assign n12299 = ~n12294 & ~n12295;
  assign n12300 = ~pi644 & ~n63074;
  assign n12301 = pi715 & ~n12300;
  assign n12302 = pi173 & ~n62765;
  assign n12303 = ~pi745 & n7359;
  assign n12304 = ~n12226 & ~n12303;
  assign n12305 = pi38 & ~n12304;
  assign n12306 = ~pi173 & n62802;
  assign n12307 = pi173 & ~n7351;
  assign n12308 = ~pi745 & ~n12307;
  assign n12309 = ~n12306 & n12308;
  assign n12310 = ~pi173 & pi745;
  assign n12311 = ~n62792 & n12310;
  assign n12312 = pi745 & ~n62792;
  assign n12313 = ~pi745 & ~n12306;
  assign n12314 = ~n12312 & ~n12313;
  assign n12315 = ~pi173 & ~n12314;
  assign n12316 = n7351 & n12313;
  assign n12317 = ~n12315 & ~n12316;
  assign n12318 = ~pi173 & ~n62792;
  assign n12319 = pi745 & ~n12318;
  assign n12320 = ~pi173 & ~pi745;
  assign n12321 = n62802 & n12320;
  assign n12322 = ~n12307 & ~n12321;
  assign n12323 = ~n12319 & n12322;
  assign n12324 = ~n12309 & ~n12311;
  assign n12325 = ~pi38 & ~n63075;
  assign n12326 = ~pi38 & n63075;
  assign n12327 = pi38 & ~n12226;
  assign n12328 = ~n12303 & n12327;
  assign n12329 = ~n12326 & ~n12328;
  assign n12330 = ~n12305 & ~n12325;
  assign n12331 = n62765 & ~n63076;
  assign n12332 = ~n12302 & ~n12331;
  assign n12333 = ~n8135 & ~n12332;
  assign n12334 = n8135 & ~n12217;
  assign n12335 = ~n12333 & ~n12334;
  assign n12336 = ~pi785 & ~n12335;
  assign n12337 = ~n8136 & ~n12217;
  assign n12338 = pi609 & n12333;
  assign n12339 = ~n12337 & ~n12338;
  assign n12340 = pi1155 & ~n12339;
  assign n12341 = ~n8148 & ~n12217;
  assign n12342 = ~pi609 & n12333;
  assign n12343 = ~n12341 & ~n12342;
  assign n12344 = ~pi1155 & ~n12343;
  assign n12345 = ~n12340 & ~n12344;
  assign n12346 = pi785 & ~n12345;
  assign n12347 = ~n12336 & ~n12346;
  assign n12348 = ~pi781 & ~n12347;
  assign n12349 = pi618 & n12347;
  assign n12350 = ~pi618 & n12217;
  assign n12351 = pi1154 & ~n12350;
  assign n12352 = ~n12349 & n12351;
  assign n12353 = ~pi618 & n12347;
  assign n12354 = pi618 & n12217;
  assign n12355 = ~pi1154 & ~n12354;
  assign n12356 = ~n12353 & n12355;
  assign n12357 = ~n12352 & ~n12356;
  assign n12358 = pi781 & ~n12357;
  assign n12359 = ~n12348 & ~n12358;
  assign n12360 = ~pi619 & ~n12359;
  assign n12361 = pi619 & ~n12217;
  assign n12362 = ~pi1159 & ~n12361;
  assign n12363 = ~n12360 & n12362;
  assign n12364 = pi619 & ~n12359;
  assign n12365 = ~pi619 & ~n12217;
  assign n12366 = pi1159 & ~n12365;
  assign n12367 = ~n12364 & n12366;
  assign n12368 = pi619 & n12359;
  assign n12369 = ~pi619 & n12217;
  assign n12370 = pi1159 & ~n12369;
  assign n12371 = ~n12368 & n12370;
  assign n12372 = ~pi619 & n12359;
  assign n12373 = pi619 & n12217;
  assign n12374 = ~pi1159 & ~n12373;
  assign n12375 = ~n12372 & n12374;
  assign n12376 = ~n12371 & ~n12375;
  assign n12377 = ~n12363 & ~n12367;
  assign n12378 = pi789 & n63077;
  assign n12379 = ~pi789 & n12359;
  assign n12380 = ~pi789 & ~n12359;
  assign n12381 = pi789 & ~n63077;
  assign n12382 = ~n12380 & ~n12381;
  assign n12383 = ~n12378 & ~n12379;
  assign n12384 = n8418 & n63078;
  assign n12385 = ~n8418 & n12217;
  assign n12386 = pi626 & n63078;
  assign n12387 = ~pi626 & n12217;
  assign n12388 = pi1158 & ~n12387;
  assign n12389 = ~n12386 & n12388;
  assign n12390 = ~pi626 & n63078;
  assign n12391 = pi626 & n12217;
  assign n12392 = ~pi1158 & ~n12391;
  assign n12393 = ~n12390 & n12392;
  assign n12394 = ~n12389 & ~n12393;
  assign n12395 = ~n12384 & ~n12385;
  assign n12396 = pi788 & n63079;
  assign n12397 = ~pi788 & n63078;
  assign n12398 = ~pi788 & ~n63078;
  assign n12399 = pi788 & ~n63079;
  assign n12400 = ~n12398 & ~n12399;
  assign n12401 = ~n12396 & ~n12397;
  assign n12402 = ~n8334 & n63080;
  assign n12403 = n8334 & n12217;
  assign n12404 = ~n12402 & ~n12403;
  assign n12405 = ~n8376 & ~n12404;
  assign n12406 = n8376 & n12217;
  assign n12407 = n8376 & ~n12217;
  assign n12408 = ~n8376 & n12404;
  assign n12409 = ~n12407 & ~n12408;
  assign n12410 = ~n12405 & ~n12406;
  assign n12411 = pi644 & n63081;
  assign n12412 = ~pi644 & n12217;
  assign n12413 = ~pi715 & ~n12412;
  assign n12414 = ~n12411 & n12413;
  assign n12415 = pi1160 & ~n12414;
  assign n12416 = ~n12301 & n12415;
  assign n12417 = ~n63052 & ~n63080;
  assign n12418 = ~pi629 & n12267;
  assign n12419 = pi629 & n12271;
  assign n12420 = ~n12418 & ~n12419;
  assign n12421 = ~n12417 & n12420;
  assign n12422 = pi792 & ~n12421;
  assign n12423 = n8525 & ~n63071;
  assign n12424 = ~n8302 & n63079;
  assign n12425 = ~n12423 & ~n12424;
  assign n12426 = pi788 & ~n12425;
  assign n12427 = pi723 & n63076;
  assign n12428 = ~pi173 & ~n62821;
  assign n12429 = pi173 & n7632;
  assign n12430 = pi745 & ~n12429;
  assign n12431 = ~n12428 & n12430;
  assign n12432 = pi173 & n7709;
  assign n12433 = ~pi173 & n62851;
  assign n12434 = ~pi745 & ~n12433;
  assign n12435 = ~n12432 & n12434;
  assign n12436 = pi39 & ~n12435;
  assign n12437 = ~n12431 & n12436;
  assign n12438 = pi173 & n7855;
  assign n12439 = ~pi173 & n7832;
  assign n12440 = pi745 & ~n12439;
  assign n12441 = ~n12438 & n12440;
  assign n12442 = ~pi173 & ~n7861;
  assign n12443 = pi173 & ~n7868;
  assign n12444 = ~pi745 & ~n12443;
  assign n12445 = ~n12442 & n12444;
  assign n12446 = ~pi39 & ~n12445;
  assign n12447 = pi173 & ~n7855;
  assign n12448 = ~pi173 & ~n7832;
  assign n12449 = pi745 & ~n12448;
  assign n12450 = pi745 & ~n12447;
  assign n12451 = ~n12448 & n12450;
  assign n12452 = ~n12447 & n12449;
  assign n12453 = ~pi173 & n7861;
  assign n12454 = pi173 & n7868;
  assign n12455 = ~pi745 & ~n12454;
  assign n12456 = ~n12453 & n12455;
  assign n12457 = ~n63082 & ~n12456;
  assign n12458 = ~pi39 & ~n12457;
  assign n12459 = ~n12441 & n12446;
  assign n12460 = ~pi38 & ~n63083;
  assign n12461 = ~n12437 & n12460;
  assign n12462 = ~pi745 & ~n7744;
  assign n12463 = n10350 & ~n12462;
  assign n12464 = ~pi173 & ~n12463;
  assign n12465 = ~pi745 & n7316;
  assign n12466 = ~n7565 & ~n12465;
  assign n12467 = pi173 & ~n12466;
  assign n12468 = n7356 & n12467;
  assign n12469 = pi38 & ~n12468;
  assign n12470 = ~n12464 & n12469;
  assign n12471 = ~pi723 & ~n12470;
  assign n12472 = ~n12461 & n12471;
  assign n12473 = n62765 & ~n12472;
  assign n12474 = ~n12427 & n12473;
  assign n12475 = ~n12302 & ~n12474;
  assign n12476 = ~pi625 & n12475;
  assign n12477 = pi625 & n12332;
  assign n12478 = ~pi1153 & ~n12477;
  assign n12479 = ~n12476 & n12478;
  assign n12480 = ~pi608 & ~n12235;
  assign n12481 = ~n12479 & n12480;
  assign n12482 = pi625 & n12475;
  assign n12483 = ~pi625 & n12332;
  assign n12484 = pi1153 & ~n12483;
  assign n12485 = ~n12482 & n12484;
  assign n12486 = pi608 & ~n12239;
  assign n12487 = ~n12485 & n12486;
  assign n12488 = ~n12481 & ~n12487;
  assign n12489 = pi778 & ~n12488;
  assign n12490 = ~pi778 & n12475;
  assign n12491 = ~n12489 & ~n12490;
  assign n12492 = ~pi609 & ~n12491;
  assign n12493 = pi609 & n12242;
  assign n12494 = ~pi1155 & ~n12493;
  assign n12495 = ~n12492 & n12494;
  assign n12496 = ~pi660 & ~n12340;
  assign n12497 = ~n12495 & n12496;
  assign n12498 = pi609 & ~n12491;
  assign n12499 = ~pi609 & n12242;
  assign n12500 = pi1155 & ~n12499;
  assign n12501 = ~n12498 & n12500;
  assign n12502 = pi660 & ~n12344;
  assign n12503 = ~n12501 & n12502;
  assign n12504 = ~n12497 & ~n12503;
  assign n12505 = pi785 & ~n12504;
  assign n12506 = ~pi785 & ~n12491;
  assign n12507 = ~n12505 & ~n12506;
  assign n12508 = pi618 & ~n12507;
  assign n12509 = ~pi618 & ~n63069;
  assign n12510 = pi1154 & ~n12509;
  assign n12511 = ~n12508 & n12510;
  assign n12512 = pi627 & ~n12356;
  assign n12513 = ~n12511 & n12512;
  assign n12514 = ~pi618 & ~n12507;
  assign n12515 = pi618 & ~n63069;
  assign n12516 = ~pi1154 & ~n12515;
  assign n12517 = ~n12514 & n12516;
  assign n12518 = ~pi627 & ~n12352;
  assign n12519 = ~n12517 & n12518;
  assign n12520 = pi781 & ~n12519;
  assign n12521 = ~n12513 & n12520;
  assign n12522 = ~n11431 & ~n63070;
  assign n12523 = ~n62884 & ~n63077;
  assign n12524 = ~n12522 & ~n12523;
  assign n12525 = pi789 & ~n12524;
  assign n12526 = ~pi781 & n12507;
  assign n12527 = ~n12525 & ~n12526;
  assign n12528 = ~n12521 & n12527;
  assign n12529 = n11434 & n12524;
  assign n12530 = ~n12528 & ~n12529;
  assign n12531 = ~n12513 & ~n12519;
  assign n12532 = pi781 & ~n12531;
  assign n12533 = ~pi781 & ~n12507;
  assign n12534 = ~n12532 & ~n12533;
  assign n12535 = ~pi619 & ~n12534;
  assign n12536 = pi619 & n63070;
  assign n12537 = ~pi1159 & ~n12536;
  assign n12538 = ~n12535 & n12537;
  assign n12539 = ~pi648 & ~n12371;
  assign n12540 = ~n12538 & n12539;
  assign n12541 = pi619 & ~n12534;
  assign n12542 = ~pi619 & n63070;
  assign n12543 = pi1159 & ~n12542;
  assign n12544 = ~n12541 & n12543;
  assign n12545 = pi648 & ~n12375;
  assign n12546 = ~n12544 & n12545;
  assign n12547 = pi789 & ~n12546;
  assign n12548 = pi789 & ~n12540;
  assign n12549 = ~n12546 & n12548;
  assign n12550 = ~n12540 & n12547;
  assign n12551 = ~pi789 & n12534;
  assign n12552 = n62894 & ~n12551;
  assign n12553 = ~n63084 & n12552;
  assign n12554 = n62894 & ~n12530;
  assign n12555 = ~n63030 & ~n63085;
  assign n12556 = ~n63030 & ~n12426;
  assign n12557 = ~n63085 & n12556;
  assign n12558 = ~n12426 & n12555;
  assign n12559 = ~n12422 & ~n63086;
  assign n12560 = ~n8651 & ~n12559;
  assign n12561 = ~n8413 & n12404;
  assign n12562 = n8373 & ~n12280;
  assign n12563 = ~pi630 & n63072;
  assign n12564 = n8374 & ~n12289;
  assign n12565 = pi630 & n12286;
  assign n12566 = ~n63087 & ~n63088;
  assign n12567 = ~n12561 & n12566;
  assign n12568 = pi787 & ~n12567;
  assign n12569 = ~n12560 & ~n12568;
  assign n12570 = ~pi644 & n12569;
  assign n12571 = pi644 & ~n63074;
  assign n12572 = ~pi715 & ~n12571;
  assign n12573 = ~n12570 & n12572;
  assign n12574 = ~pi644 & n63081;
  assign n12575 = pi644 & n12217;
  assign n12576 = pi715 & ~n12575;
  assign n12577 = ~n12574 & n12576;
  assign n12578 = ~pi1160 & ~n12577;
  assign n12579 = ~n12573 & n12578;
  assign n12580 = ~n12416 & ~n12579;
  assign n12581 = pi790 & ~n12580;
  assign n12582 = pi644 & n12415;
  assign n12583 = pi790 & ~n12582;
  assign n12584 = n12569 & ~n12583;
  assign n12585 = ~n12581 & ~n12584;
  assign n12586 = n62455 & ~n12585;
  assign n12587 = ~pi173 & ~n62455;
  assign n12588 = ~pi832 & ~n12587;
  assign n12589 = ~n12586 & n12588;
  assign n12590 = ~pi173 & ~n2923;
  assign n12591 = ~n8418 & n12590;
  assign n12592 = ~n12465 & ~n12590;
  assign n12593 = ~n8420 & ~n12592;
  assign n12594 = ~pi785 & ~n12593;
  assign n12595 = n8148 & n12465;
  assign n12596 = n12593 & ~n12595;
  assign n12597 = pi1155 & ~n12596;
  assign n12598 = ~pi1155 & ~n12590;
  assign n12599 = ~n12595 & n12598;
  assign n12600 = ~n12597 & ~n12599;
  assign n12601 = pi785 & ~n12600;
  assign n12602 = ~n12594 & ~n12601;
  assign n12603 = ~pi781 & ~n12602;
  assign n12604 = ~n8435 & n12602;
  assign n12605 = pi1154 & ~n12604;
  assign n12606 = ~n8438 & n12602;
  assign n12607 = ~pi1154 & ~n12606;
  assign n12608 = ~n12605 & ~n12607;
  assign n12609 = pi781 & ~n12608;
  assign n12610 = ~n12603 & ~n12609;
  assign n12611 = ~pi789 & ~n12610;
  assign n12612 = ~pi619 & n2923;
  assign n12613 = n12610 & ~n12612;
  assign n12614 = pi1159 & ~n12613;
  assign n12615 = pi619 & n2923;
  assign n12616 = n12610 & ~n12615;
  assign n12617 = ~pi1159 & ~n12616;
  assign n12618 = ~n12614 & ~n12617;
  assign n12619 = pi789 & ~n12618;
  assign n12620 = ~n12611 & ~n12619;
  assign n12621 = n8418 & n12620;
  assign n12622 = pi626 & n12620;
  assign n12623 = ~pi626 & n12590;
  assign n12624 = pi1158 & ~n12623;
  assign n12625 = ~n12622 & n12624;
  assign n12626 = ~pi626 & n12620;
  assign n12627 = pi626 & n12590;
  assign n12628 = ~pi1158 & ~n12627;
  assign n12629 = ~n12626 & n12628;
  assign n12630 = ~n12625 & ~n12629;
  assign n12631 = ~n12591 & ~n12621;
  assign n12632 = pi788 & n63089;
  assign n12633 = ~pi788 & n12620;
  assign n12634 = ~pi788 & ~n12620;
  assign n12635 = pi788 & ~n63089;
  assign n12636 = ~n12634 & ~n12635;
  assign n12637 = ~n12632 & ~n12633;
  assign n12638 = ~n8334 & n63090;
  assign n12639 = n8334 & n12590;
  assign n12640 = ~n8413 & ~n12639;
  assign n12641 = ~n12638 & ~n12639;
  assign n12642 = ~n8413 & n12641;
  assign n12643 = ~n12638 & n12640;
  assign n12644 = ~pi723 & n7564;
  assign n12645 = ~n12590 & ~n12644;
  assign n12646 = ~pi778 & ~n12645;
  assign n12647 = ~pi625 & n12644;
  assign n12648 = ~n12645 & ~n12647;
  assign n12649 = pi1153 & ~n12648;
  assign n12650 = ~pi1153 & ~n12590;
  assign n12651 = ~n12647 & n12650;
  assign n12652 = pi778 & ~n12651;
  assign n12653 = ~n12649 & n12652;
  assign n12654 = ~n12646 & ~n12653;
  assign n12655 = ~n8490 & ~n12654;
  assign n12656 = ~n8492 & n12655;
  assign n12657 = ~n8494 & n12656;
  assign n12658 = ~n8496 & n12657;
  assign n12659 = ~n8508 & n12658;
  assign n12660 = pi647 & ~n12659;
  assign n12661 = ~pi647 & ~n12590;
  assign n12662 = ~n12660 & ~n12661;
  assign n12663 = n8373 & ~n12662;
  assign n12664 = ~pi647 & n12659;
  assign n12665 = pi647 & n12590;
  assign n12666 = ~pi1157 & ~n12665;
  assign n12667 = ~n12664 & n12666;
  assign n12668 = pi630 & n12667;
  assign n12669 = ~n12663 & ~n12668;
  assign n12670 = ~n63091 & n12669;
  assign n12671 = pi787 & ~n12670;
  assign n12672 = n8525 & n12657;
  assign n12673 = ~n8302 & n63089;
  assign n12674 = ~n12672 & ~n12673;
  assign n12675 = pi788 & ~n12674;
  assign n12676 = ~n7187 & ~n12645;
  assign n12677 = pi625 & n12676;
  assign n12678 = n12592 & ~n12676;
  assign n12679 = ~n12677 & ~n12678;
  assign n12680 = n12650 & ~n12679;
  assign n12681 = ~pi608 & ~n12649;
  assign n12682 = ~n12680 & n12681;
  assign n12683 = pi1153 & n12592;
  assign n12684 = ~n12677 & n12683;
  assign n12685 = pi608 & ~n12651;
  assign n12686 = ~n12684 & n12685;
  assign n12687 = ~n12682 & ~n12686;
  assign n12688 = pi778 & ~n12687;
  assign n12689 = ~pi778 & ~n12678;
  assign n12690 = ~n12688 & ~n12689;
  assign n12691 = ~pi609 & ~n12690;
  assign n12692 = pi609 & ~n12654;
  assign n12693 = ~pi1155 & ~n12692;
  assign n12694 = ~n12691 & n12693;
  assign n12695 = ~pi660 & ~n12597;
  assign n12696 = ~n12694 & n12695;
  assign n12697 = pi609 & ~n12690;
  assign n12698 = ~pi609 & ~n12654;
  assign n12699 = pi1155 & ~n12698;
  assign n12700 = ~n12697 & n12699;
  assign n12701 = pi660 & ~n12599;
  assign n12702 = ~n12700 & n12701;
  assign n12703 = ~n12696 & ~n12702;
  assign n12704 = pi785 & ~n12703;
  assign n12705 = ~pi785 & ~n12690;
  assign n12706 = ~n12704 & ~n12705;
  assign n12707 = ~pi618 & ~n12706;
  assign n12708 = pi618 & n12655;
  assign n12709 = ~pi1154 & ~n12708;
  assign n12710 = ~n12707 & n12709;
  assign n12711 = ~pi627 & ~n12605;
  assign n12712 = ~n12710 & n12711;
  assign n12713 = pi618 & ~n12706;
  assign n12714 = ~pi618 & n12655;
  assign n12715 = pi1154 & ~n12714;
  assign n12716 = ~n12713 & n12715;
  assign n12717 = pi627 & ~n12607;
  assign n12718 = ~n12716 & n12717;
  assign n12719 = ~n12712 & ~n12718;
  assign n12720 = pi781 & ~n12719;
  assign n12721 = ~pi781 & ~n12706;
  assign n12722 = ~n12720 & ~n12721;
  assign n12723 = pi619 & ~n12722;
  assign n12724 = ~pi619 & n12656;
  assign n12725 = pi1159 & ~n12724;
  assign n12726 = ~n12723 & n12725;
  assign n12727 = pi648 & ~n12617;
  assign n12728 = ~n12726 & n12727;
  assign n12729 = ~pi619 & ~n12722;
  assign n12730 = pi619 & n12656;
  assign n12731 = ~pi1159 & ~n12730;
  assign n12732 = ~n12729 & n12731;
  assign n12733 = ~pi648 & ~n12614;
  assign n12734 = ~n12732 & n12733;
  assign n12735 = pi789 & ~n12734;
  assign n12736 = pi789 & ~n12728;
  assign n12737 = ~n12734 & n12736;
  assign n12738 = ~n12728 & n12735;
  assign n12739 = ~pi789 & n12722;
  assign n12740 = n62894 & ~n12739;
  assign n12741 = ~n63092 & n12740;
  assign n12742 = ~n12675 & ~n12741;
  assign n12743 = ~n63030 & ~n12742;
  assign n12744 = n8498 & n63090;
  assign n12745 = n8615 & n12658;
  assign n12746 = pi629 & ~n12745;
  assign n12747 = ~n12744 & n12746;
  assign n12748 = n8499 & n63090;
  assign n12749 = n8606 & n12658;
  assign n12750 = ~pi629 & ~n12749;
  assign n12751 = ~n12748 & n12750;
  assign n12752 = pi792 & ~n12751;
  assign n12753 = pi792 & ~n12747;
  assign n12754 = ~n12751 & n12753;
  assign n12755 = ~n12748 & ~n12749;
  assign n12756 = ~pi629 & ~n12755;
  assign n12757 = ~n12744 & ~n12745;
  assign n12758 = pi629 & ~n12757;
  assign n12759 = ~n12756 & ~n12758;
  assign n12760 = pi792 & ~n12759;
  assign n12761 = ~n12747 & n12752;
  assign n12762 = ~n8651 & ~n63093;
  assign n12763 = ~n12743 & n12762;
  assign n12764 = ~n12671 & ~n12763;
  assign n12765 = pi644 & n12764;
  assign n12766 = ~pi787 & ~n12659;
  assign n12767 = pi1157 & ~n12662;
  assign n12768 = ~n12667 & ~n12767;
  assign n12769 = pi787 & ~n12768;
  assign n12770 = ~n12766 & ~n12769;
  assign n12771 = ~pi644 & n12770;
  assign n12772 = pi715 & ~n12771;
  assign n12773 = ~n12765 & n12772;
  assign n12774 = ~n8685 & n12590;
  assign n12775 = ~n8376 & n12638;
  assign n12776 = ~n8376 & ~n12641;
  assign n12777 = n8376 & n12590;
  assign n12778 = ~n12776 & ~n12777;
  assign n12779 = ~n12774 & ~n12775;
  assign n12780 = pi644 & ~n63094;
  assign n12781 = ~pi644 & n12590;
  assign n12782 = ~pi715 & ~n12781;
  assign n12783 = ~n12780 & n12782;
  assign n12784 = pi1160 & ~n12783;
  assign n12785 = ~n12773 & n12784;
  assign n12786 = ~pi644 & n12764;
  assign n12787 = pi644 & n12770;
  assign n12788 = ~pi715 & ~n12787;
  assign n12789 = ~n12786 & n12788;
  assign n12790 = ~pi644 & ~n63094;
  assign n12791 = pi644 & n12590;
  assign n12792 = pi715 & ~n12791;
  assign n12793 = ~n12790 & n12792;
  assign n12794 = ~pi1160 & ~n12793;
  assign n12795 = ~n12789 & n12794;
  assign n12796 = ~n12785 & ~n12795;
  assign n12797 = pi790 & ~n12796;
  assign n12798 = ~pi790 & n12764;
  assign n12799 = pi832 & ~n12798;
  assign n12800 = ~n12797 & n12799;
  assign po330 = ~n12589 & ~n12800;
  assign n12802 = pi174 & ~n8098;
  assign n12803 = ~n8685 & n12802;
  assign n12804 = pi174 & ~n62765;
  assign n12805 = ~pi759 & ~n7143;
  assign n12806 = pi759 & ~n62801;
  assign n12807 = ~n12805 & ~n12806;
  assign n12808 = pi39 & ~n12807;
  assign n12809 = pi759 & n62793;
  assign n12810 = ~pi759 & ~n62781;
  assign n12811 = ~pi39 & ~n12810;
  assign n12812 = ~n12809 & n12811;
  assign n12813 = ~n12808 & ~n12812;
  assign n12814 = pi174 & ~n12813;
  assign n12815 = ~pi174 & pi759;
  assign n12816 = n7351 & n12815;
  assign n12817 = ~n12814 & ~n12816;
  assign n12818 = ~pi38 & ~n12817;
  assign n12819 = pi759 & n7187;
  assign n12820 = n7357 & ~n12819;
  assign n12821 = ~pi174 & ~n7357;
  assign n12822 = pi38 & ~n12821;
  assign n12823 = pi38 & ~n12820;
  assign n12824 = ~n12821 & n12823;
  assign n12825 = ~n12820 & n12822;
  assign n12826 = ~n12818 & ~n63095;
  assign n12827 = n62765 & ~n12826;
  assign n12828 = ~n12804 & ~n12827;
  assign n12829 = ~n8135 & ~n12828;
  assign n12830 = n8135 & n12802;
  assign n12831 = n8135 & ~n12802;
  assign n12832 = ~n8135 & n12828;
  assign n12833 = ~n12831 & ~n12832;
  assign n12834 = ~n12829 & ~n12830;
  assign n12835 = ~pi785 & n63096;
  assign n12836 = pi609 & ~n63096;
  assign n12837 = ~pi609 & ~n12802;
  assign n12838 = pi1155 & ~n12837;
  assign n12839 = ~n12836 & n12838;
  assign n12840 = ~pi609 & ~n63096;
  assign n12841 = pi609 & ~n12802;
  assign n12842 = ~pi1155 & ~n12841;
  assign n12843 = ~n12840 & n12842;
  assign n12844 = ~n12839 & ~n12843;
  assign n12845 = pi785 & ~n12844;
  assign n12846 = ~n12835 & ~n12845;
  assign n12847 = ~pi781 & ~n12846;
  assign n12848 = pi618 & n12846;
  assign n12849 = ~pi618 & ~n12802;
  assign n12850 = pi1154 & ~n12849;
  assign n12851 = ~n12848 & n12850;
  assign n12852 = ~pi618 & n12846;
  assign n12853 = pi618 & ~n12802;
  assign n12854 = ~pi1154 & ~n12853;
  assign n12855 = ~n12852 & n12854;
  assign n12856 = ~n12851 & ~n12855;
  assign n12857 = pi781 & ~n12856;
  assign n12858 = ~n12847 & ~n12857;
  assign n12859 = ~n11306 & n12858;
  assign n12860 = n11306 & ~n12802;
  assign n12861 = ~pi789 & ~n12858;
  assign n12862 = pi619 & n12858;
  assign n12863 = ~pi619 & ~n12802;
  assign n12864 = pi1159 & ~n12863;
  assign n12865 = ~n12862 & n12864;
  assign n12866 = ~pi619 & n12858;
  assign n12867 = pi619 & ~n12802;
  assign n12868 = ~pi1159 & ~n12867;
  assign n12869 = ~n12866 & n12868;
  assign n12870 = ~n12865 & ~n12869;
  assign n12871 = pi789 & ~n12870;
  assign n12872 = ~n12861 & ~n12871;
  assign n12873 = ~n12859 & ~n12860;
  assign n12874 = ~n8595 & ~n63097;
  assign n12875 = n8595 & n12802;
  assign n12876 = ~n12874 & ~n12875;
  assign n12877 = ~n8334 & ~n12876;
  assign n12878 = ~n8376 & n12877;
  assign n12879 = n8334 & n12802;
  assign n12880 = ~n12877 & ~n12879;
  assign n12881 = ~n8376 & ~n12880;
  assign n12882 = n8376 & n12802;
  assign n12883 = ~n12881 & ~n12882;
  assign n12884 = n8376 & ~n12802;
  assign n12885 = ~n8376 & n12880;
  assign n12886 = ~n12884 & ~n12885;
  assign n12887 = ~n12803 & ~n12878;
  assign n12888 = pi644 & n63098;
  assign n12889 = ~pi644 & ~n12802;
  assign n12890 = ~pi715 & ~n12889;
  assign n12891 = ~n12888 & n12890;
  assign n12892 = pi1160 & ~n12891;
  assign n12893 = n8257 & ~n12802;
  assign n12894 = n62880 & ~n12802;
  assign n12895 = pi696 & n62765;
  assign n12896 = n10997 & ~n12821;
  assign n12897 = pi174 & ~n8009;
  assign n12898 = ~pi174 & ~n62874;
  assign n12899 = ~pi38 & ~n12898;
  assign n12900 = ~n12897 & n12899;
  assign n12901 = ~n12896 & ~n12900;
  assign n12902 = n12895 & ~n12901;
  assign n12903 = n12802 & ~n12895;
  assign n12904 = ~n12802 & ~n12895;
  assign n12905 = n12895 & ~n12896;
  assign n12906 = ~n12900 & n12905;
  assign n12907 = ~n12904 & ~n12906;
  assign n12908 = ~n12902 & ~n12903;
  assign n12909 = ~pi778 & n63099;
  assign n12910 = pi625 & ~n63099;
  assign n12911 = ~pi625 & ~n12802;
  assign n12912 = pi1153 & ~n12911;
  assign n12913 = ~n12910 & n12912;
  assign n12914 = ~pi625 & ~n63099;
  assign n12915 = pi625 & ~n12802;
  assign n12916 = ~pi1153 & ~n12915;
  assign n12917 = ~n12914 & n12916;
  assign n12918 = ~n12913 & ~n12917;
  assign n12919 = pi778 & ~n12918;
  assign n12920 = ~n12909 & ~n12919;
  assign n12921 = ~n62880 & n12920;
  assign n12922 = ~n62880 & ~n12920;
  assign n12923 = n62880 & n12802;
  assign n12924 = ~n12922 & ~n12923;
  assign n12925 = ~n12894 & ~n12921;
  assign n12926 = ~n62882 & ~n63100;
  assign n12927 = n62882 & n12802;
  assign n12928 = n62882 & ~n12802;
  assign n12929 = ~n62882 & n63100;
  assign n12930 = ~n12928 & ~n12929;
  assign n12931 = ~n12926 & ~n12927;
  assign n12932 = ~n8257 & ~n63101;
  assign n12933 = ~n8257 & n63101;
  assign n12934 = n8257 & n12802;
  assign n12935 = ~n12933 & ~n12934;
  assign n12936 = ~n12893 & ~n12932;
  assign n12937 = ~n8303 & ~n63102;
  assign n12938 = n8303 & n12802;
  assign n12939 = n8303 & ~n12802;
  assign n12940 = ~n8303 & n63102;
  assign n12941 = ~n12939 & ~n12940;
  assign n12942 = ~n12937 & ~n12938;
  assign n12943 = ~pi792 & n63103;
  assign n12944 = pi628 & ~n63103;
  assign n12945 = ~pi628 & ~n12802;
  assign n12946 = pi1156 & ~n12945;
  assign n12947 = ~n12944 & n12946;
  assign n12948 = ~pi628 & ~n63103;
  assign n12949 = pi628 & ~n12802;
  assign n12950 = ~pi1156 & ~n12949;
  assign n12951 = ~n12948 & n12950;
  assign n12952 = ~n12947 & ~n12951;
  assign n12953 = pi792 & ~n12952;
  assign n12954 = ~n12943 & ~n12953;
  assign n12955 = ~pi787 & ~n12954;
  assign n12956 = pi647 & n12954;
  assign n12957 = ~pi647 & ~n12802;
  assign n12958 = pi1157 & ~n12957;
  assign n12959 = pi647 & ~n12954;
  assign n12960 = ~pi647 & n12802;
  assign n12961 = ~n12959 & ~n12960;
  assign n12962 = pi1157 & ~n12961;
  assign n12963 = ~n12956 & n12958;
  assign n12964 = ~pi647 & n12954;
  assign n12965 = pi647 & ~n12802;
  assign n12966 = ~pi1157 & ~n12965;
  assign n12967 = ~n12964 & n12966;
  assign n12968 = ~n63104 & ~n12967;
  assign n12969 = pi787 & ~n12968;
  assign n12970 = ~n12955 & ~n12969;
  assign n12971 = ~pi644 & n12970;
  assign n12972 = pi715 & ~n12971;
  assign n12973 = n8373 & ~n12961;
  assign n12974 = pi630 & n12967;
  assign n12975 = ~n8413 & ~n12880;
  assign n12976 = ~n12974 & ~n12975;
  assign n12977 = ~n12973 & n12976;
  assign n12978 = pi787 & ~n12977;
  assign n12979 = ~n8302 & ~n8524;
  assign n12980 = n63097 & n12979;
  assign n12981 = ~pi641 & ~n63102;
  assign n12982 = pi641 & n12802;
  assign n12983 = n8417 & ~n12982;
  assign n12984 = ~n12981 & n12983;
  assign n12985 = pi641 & ~n63102;
  assign n12986 = ~pi641 & n12802;
  assign n12987 = n8416 & ~n12986;
  assign n12988 = ~n12985 & n12987;
  assign n12989 = ~n12984 & ~n12988;
  assign n12990 = ~n12980 & n12989;
  assign n12991 = pi788 & ~n12990;
  assign n12992 = ~pi696 & n12818;
  assign n12993 = pi174 & ~n62821;
  assign n12994 = ~pi174 & n7632;
  assign n12995 = ~pi759 & ~n12994;
  assign n12996 = ~n12993 & n12995;
  assign n12997 = ~pi174 & n7709;
  assign n12998 = pi174 & n62851;
  assign n12999 = pi759 & ~n12998;
  assign n13000 = ~n12997 & n12999;
  assign n13001 = pi39 & ~n13000;
  assign n13002 = ~n12996 & n13001;
  assign n13003 = pi174 & ~n7832;
  assign n13004 = ~pi174 & ~n7855;
  assign n13005 = ~pi759 & ~n13004;
  assign n13006 = ~pi759 & ~n13003;
  assign n13007 = ~n13004 & n13006;
  assign n13008 = ~n13003 & n13005;
  assign n13009 = pi174 & n7861;
  assign n13010 = ~pi174 & n7868;
  assign n13011 = pi759 & ~n13010;
  assign n13012 = ~n13009 & n13011;
  assign n13013 = ~n63105 & ~n13012;
  assign n13014 = ~pi39 & ~n13013;
  assign n13015 = ~pi38 & ~n13014;
  assign n13016 = ~n13002 & n13015;
  assign n13017 = pi696 & ~n8793;
  assign n13018 = pi174 & n62821;
  assign n13019 = ~pi174 & ~n7632;
  assign n13020 = ~pi759 & ~n13019;
  assign n13021 = ~n13018 & n13020;
  assign n13022 = ~pi174 & ~n7709;
  assign n13023 = pi174 & ~n62851;
  assign n13024 = pi759 & ~n13023;
  assign n13025 = ~n13022 & n13024;
  assign n13026 = pi39 & ~n13025;
  assign n13027 = ~n13021 & n13026;
  assign n13028 = ~pi39 & ~n13012;
  assign n13029 = ~n63105 & n13028;
  assign n13030 = ~pi38 & ~n13029;
  assign n13031 = ~n13027 & n13030;
  assign n13032 = ~n10357 & ~n13031;
  assign n13033 = pi696 & ~n13032;
  assign n13034 = ~n13016 & n13017;
  assign n13035 = ~n63095 & ~n63106;
  assign n13036 = ~n12992 & n13035;
  assign n13037 = ~pi696 & n12826;
  assign n13038 = pi696 & ~n10357;
  assign n13039 = ~n63095 & n13038;
  assign n13040 = ~n13031 & n13039;
  assign n13041 = n62765 & ~n13040;
  assign n13042 = ~n13037 & n13041;
  assign n13043 = n62765 & ~n13036;
  assign n13044 = ~n12804 & ~n63107;
  assign n13045 = pi625 & n13044;
  assign n13046 = ~pi625 & n12828;
  assign n13047 = pi1153 & ~n13046;
  assign n13048 = ~n13045 & n13047;
  assign n13049 = pi608 & ~n12917;
  assign n13050 = ~n13048 & n13049;
  assign n13051 = ~pi625 & n13044;
  assign n13052 = pi625 & n12828;
  assign n13053 = ~pi1153 & ~n13052;
  assign n13054 = ~n13051 & n13053;
  assign n13055 = ~pi608 & ~n12913;
  assign n13056 = ~n13054 & n13055;
  assign n13057 = ~n13050 & ~n13056;
  assign n13058 = pi778 & ~n13057;
  assign n13059 = ~pi778 & n13044;
  assign n13060 = ~n13058 & ~n13059;
  assign n13061 = ~pi609 & ~n13060;
  assign n13062 = pi609 & n12920;
  assign n13063 = ~pi1155 & ~n13062;
  assign n13064 = ~n13061 & n13063;
  assign n13065 = ~pi660 & ~n12839;
  assign n13066 = ~n13064 & n13065;
  assign n13067 = pi609 & ~n13060;
  assign n13068 = ~pi609 & n12920;
  assign n13069 = pi1155 & ~n13068;
  assign n13070 = ~n13067 & n13069;
  assign n13071 = pi660 & ~n12843;
  assign n13072 = ~n13070 & n13071;
  assign n13073 = ~n13066 & ~n13072;
  assign n13074 = pi785 & ~n13073;
  assign n13075 = ~pi785 & ~n13060;
  assign n13076 = ~n13074 & ~n13075;
  assign n13077 = ~pi618 & ~n13076;
  assign n13078 = pi618 & n63100;
  assign n13079 = ~pi1154 & ~n13078;
  assign n13080 = ~n13077 & n13079;
  assign n13081 = ~pi627 & ~n12851;
  assign n13082 = ~n13080 & n13081;
  assign n13083 = pi618 & ~n13076;
  assign n13084 = ~pi618 & n63100;
  assign n13085 = pi1154 & ~n13084;
  assign n13086 = ~n13083 & n13085;
  assign n13087 = pi627 & ~n12855;
  assign n13088 = ~n13086 & n13087;
  assign n13089 = ~n13082 & ~n13088;
  assign n13090 = pi781 & ~n13089;
  assign n13091 = ~pi781 & ~n13076;
  assign n13092 = ~n11434 & ~n13091;
  assign n13093 = ~n13090 & n13092;
  assign n13094 = n8253 & ~n12863;
  assign n13095 = ~n12862 & n13094;
  assign n13096 = n8254 & ~n12867;
  assign n13097 = ~n12866 & n13096;
  assign n13098 = ~n11431 & n63101;
  assign n13099 = ~n13097 & ~n13098;
  assign n13100 = ~n13095 & n13099;
  assign n13101 = pi789 & ~n13100;
  assign n13102 = n62894 & ~n13101;
  assign n13103 = ~n13090 & ~n13091;
  assign n13104 = ~pi619 & ~n13103;
  assign n13105 = pi619 & ~n63101;
  assign n13106 = ~pi1159 & ~n13105;
  assign n13107 = ~n13104 & n13106;
  assign n13108 = ~pi648 & ~n12865;
  assign n13109 = ~n13107 & n13108;
  assign n13110 = pi619 & ~n13103;
  assign n13111 = ~pi619 & ~n63101;
  assign n13112 = pi1159 & ~n13111;
  assign n13113 = ~n13110 & n13112;
  assign n13114 = pi648 & ~n12869;
  assign n13115 = ~n13113 & n13114;
  assign n13116 = pi789 & ~n13115;
  assign n13117 = ~n13109 & n13116;
  assign n13118 = ~pi789 & n13103;
  assign n13119 = n62894 & ~n13118;
  assign n13120 = ~n13117 & n13119;
  assign n13121 = ~n13093 & n13102;
  assign n13122 = ~n13109 & ~n13115;
  assign n13123 = pi789 & ~n13122;
  assign n13124 = ~pi789 & ~n13103;
  assign n13125 = ~n13123 & ~n13124;
  assign n13126 = ~pi788 & n13125;
  assign n13127 = ~pi626 & n13125;
  assign n13128 = pi626 & ~n63102;
  assign n13129 = ~pi641 & ~n13128;
  assign n13130 = ~n13127 & n13129;
  assign n13131 = ~pi626 & ~n63097;
  assign n13132 = pi626 & n12802;
  assign n13133 = pi641 & ~n13132;
  assign n13134 = ~n13131 & n13133;
  assign n13135 = ~pi1158 & ~n13134;
  assign n13136 = ~n13130 & n13135;
  assign n13137 = pi626 & n13125;
  assign n13138 = ~pi626 & ~n63102;
  assign n13139 = pi641 & ~n13138;
  assign n13140 = ~n13137 & n13139;
  assign n13141 = pi626 & ~n63097;
  assign n13142 = ~pi626 & n12802;
  assign n13143 = ~pi641 & ~n13142;
  assign n13144 = ~n13141 & n13143;
  assign n13145 = pi1158 & ~n13144;
  assign n13146 = ~n13140 & n13145;
  assign n13147 = ~n13136 & ~n13146;
  assign n13148 = pi788 & ~n13147;
  assign n13149 = ~n13126 & ~n13148;
  assign n13150 = ~n12991 & ~n63108;
  assign n13151 = ~pi628 & n63109;
  assign n13152 = pi628 & n12876;
  assign n13153 = ~pi1156 & ~n13152;
  assign n13154 = ~n13151 & n13153;
  assign n13155 = ~pi629 & ~n12947;
  assign n13156 = ~n13154 & n13155;
  assign n13157 = pi628 & n63109;
  assign n13158 = ~pi628 & n12876;
  assign n13159 = pi1156 & ~n13158;
  assign n13160 = ~n13157 & n13159;
  assign n13161 = pi629 & ~n12951;
  assign n13162 = ~n13160 & n13161;
  assign n13163 = ~n13156 & ~n13162;
  assign n13164 = pi792 & ~n13163;
  assign n13165 = ~pi792 & n63109;
  assign n13166 = ~n8651 & ~n13165;
  assign n13167 = ~n13164 & n13166;
  assign n13168 = ~n13164 & ~n13165;
  assign n13169 = ~pi647 & ~n13168;
  assign n13170 = pi647 & n12880;
  assign n13171 = ~pi1157 & ~n13170;
  assign n13172 = ~n13169 & n13171;
  assign n13173 = ~pi630 & ~n63104;
  assign n13174 = ~n13172 & n13173;
  assign n13175 = pi647 & ~n13168;
  assign n13176 = ~pi647 & n12880;
  assign n13177 = pi1157 & ~n13176;
  assign n13178 = ~n13175 & n13177;
  assign n13179 = pi630 & ~n12967;
  assign n13180 = ~n13178 & n13179;
  assign n13181 = ~n13174 & ~n13180;
  assign n13182 = pi787 & ~n13181;
  assign n13183 = ~pi787 & ~n13168;
  assign n13184 = ~n13182 & ~n13183;
  assign n13185 = ~n12978 & ~n13167;
  assign n13186 = pi644 & ~n63110;
  assign n13187 = n12972 & ~n13186;
  assign n13188 = n12892 & ~n13187;
  assign n13189 = ~pi644 & ~n63110;
  assign n13190 = pi644 & n12970;
  assign n13191 = ~pi715 & ~n13190;
  assign n13192 = ~n13189 & n13191;
  assign n13193 = ~pi644 & n63098;
  assign n13194 = pi644 & ~n12802;
  assign n13195 = pi715 & ~n13194;
  assign n13196 = ~n13193 & n13195;
  assign n13197 = ~pi1160 & ~n13196;
  assign n13198 = ~n13192 & n13197;
  assign n13199 = pi790 & ~n13198;
  assign n13200 = pi790 & ~n13188;
  assign n13201 = ~n13198 & n13200;
  assign n13202 = ~n13188 & n13199;
  assign n13203 = ~pi790 & n63110;
  assign n13204 = n3475 & ~n13203;
  assign n13205 = n12892 & ~n12972;
  assign n13206 = ~n13198 & ~n13205;
  assign n13207 = pi790 & ~n13206;
  assign n13208 = pi644 & n12892;
  assign n13209 = pi790 & ~n13208;
  assign n13210 = ~n63110 & ~n13209;
  assign n13211 = ~n13207 & ~n13210;
  assign n13212 = n3475 & ~n13211;
  assign n13213 = ~n63111 & n13204;
  assign n13214 = ~pi174 & ~n3475;
  assign n13215 = ~pi57 & ~n13214;
  assign n13216 = ~n63112 & n13215;
  assign n13217 = pi57 & pi174;
  assign n13218 = ~pi832 & ~n13217;
  assign n13219 = ~n13216 & n13218;
  assign n13220 = pi696 & n7564;
  assign n13221 = pi696 & n7565;
  assign n13222 = ~n7187 & n13220;
  assign n13223 = pi625 & n13220;
  assign n13224 = ~n7187 & n13223;
  assign n13225 = pi625 & n63113;
  assign n13226 = pi174 & ~n2923;
  assign n13227 = pi759 & n7316;
  assign n13228 = ~n13226 & ~n13227;
  assign n13229 = ~n63113 & n13228;
  assign n13230 = ~n63114 & ~n13229;
  assign n13231 = ~pi1153 & ~n13230;
  assign n13232 = pi1153 & ~n13226;
  assign n13233 = ~n13223 & n13232;
  assign n13234 = ~pi608 & ~n13233;
  assign n13235 = ~n13231 & n13234;
  assign n13236 = pi1153 & n13228;
  assign n13237 = ~n13227 & n13232;
  assign n13238 = ~n63114 & n63115;
  assign n13239 = ~n13220 & ~n13226;
  assign n13240 = ~n13223 & ~n13239;
  assign n13241 = ~pi1153 & ~n13240;
  assign n13242 = pi608 & ~n13241;
  assign n13243 = pi608 & ~n13238;
  assign n13244 = ~n13241 & n13243;
  assign n13245 = ~n13238 & n13242;
  assign n13246 = ~n13235 & ~n63116;
  assign n13247 = pi778 & ~n13246;
  assign n13248 = ~pi778 & ~n13229;
  assign n13249 = ~n13247 & ~n13248;
  assign n13250 = ~pi609 & ~n13249;
  assign n13251 = ~pi778 & n13239;
  assign n13252 = ~n13233 & ~n13241;
  assign n13253 = pi778 & ~n13252;
  assign n13254 = ~n13251 & ~n13253;
  assign n13255 = pi609 & n13254;
  assign n13256 = ~pi1155 & ~n13255;
  assign n13257 = ~n13250 & n13256;
  assign n13258 = n8136 & n13227;
  assign n13259 = pi1155 & ~n13226;
  assign n13260 = ~n13258 & n13259;
  assign n13261 = ~pi660 & ~n13260;
  assign n13262 = ~n13257 & n13261;
  assign n13263 = pi609 & ~n13249;
  assign n13264 = ~pi609 & n13254;
  assign n13265 = pi1155 & ~n13264;
  assign n13266 = ~n13263 & n13265;
  assign n13267 = n8148 & n13227;
  assign n13268 = ~pi1155 & ~n13226;
  assign n13269 = ~n13267 & n13268;
  assign n13270 = pi660 & ~n13269;
  assign n13271 = ~n13266 & n13270;
  assign n13272 = ~n13262 & ~n13271;
  assign n13273 = pi785 & ~n13272;
  assign n13274 = ~pi785 & ~n13249;
  assign n13275 = ~n13273 & ~n13274;
  assign n13276 = ~pi618 & ~n13275;
  assign n13277 = ~n62880 & n13254;
  assign n13278 = ~n13226 & ~n13277;
  assign n13279 = pi618 & ~n13278;
  assign n13280 = ~pi1154 & ~n13279;
  assign n13281 = ~n13276 & n13280;
  assign n13282 = ~n63011 & n13227;
  assign n13283 = n11386 & n13282;
  assign n13284 = pi1154 & ~n13226;
  assign n13285 = ~n13283 & n13284;
  assign n13286 = ~pi627 & ~n13285;
  assign n13287 = ~n13281 & n13286;
  assign n13288 = pi618 & ~n13275;
  assign n13289 = ~pi618 & ~n13278;
  assign n13290 = pi1154 & ~n13289;
  assign n13291 = ~n13288 & n13290;
  assign n13292 = n11388 & n13282;
  assign n13293 = ~pi1154 & ~n13226;
  assign n13294 = ~n13292 & n13293;
  assign n13295 = pi627 & ~n13294;
  assign n13296 = ~n13291 & n13295;
  assign n13297 = ~n13287 & ~n13296;
  assign n13298 = pi781 & ~n13297;
  assign n13299 = ~pi781 & ~n13275;
  assign n13300 = ~n11434 & ~n13299;
  assign n13301 = ~n13298 & n13300;
  assign n13302 = n10106 & n13254;
  assign n13303 = ~n11431 & ~n13302;
  assign n13304 = ~n8135 & n11305;
  assign n13305 = ~n63012 & n13304;
  assign n13306 = n13282 & n13305;
  assign n13307 = ~n63012 & n13282;
  assign n13308 = ~n62884 & ~n13307;
  assign n13309 = ~n62884 & ~n13304;
  assign n13310 = ~n13308 & ~n13309;
  assign n13311 = n11438 & n13307;
  assign n13312 = n8254 & ~n13311;
  assign n13313 = n11447 & n13307;
  assign n13314 = n8253 & ~n13313;
  assign n13315 = ~n13312 & ~n13314;
  assign n13316 = ~n62884 & ~n13306;
  assign n13317 = ~n13303 & n63117;
  assign n13318 = pi789 & ~n13226;
  assign n13319 = ~n13317 & n13318;
  assign n13320 = n62894 & ~n13319;
  assign n13321 = ~n13301 & n13320;
  assign n13322 = ~n8257 & n13302;
  assign n13323 = ~n13226 & ~n13322;
  assign n13324 = n8417 & ~n13323;
  assign n13325 = n63013 & n13282;
  assign n13326 = pi626 & n13325;
  assign n13327 = ~n13226 & ~n13326;
  assign n13328 = pi1158 & ~n13327;
  assign n13329 = ~pi641 & ~n13328;
  assign n13330 = ~n13324 & n13329;
  assign n13331 = n8416 & ~n13323;
  assign n13332 = ~pi626 & n13325;
  assign n13333 = ~n13226 & ~n13332;
  assign n13334 = ~pi1158 & ~n13333;
  assign n13335 = pi641 & ~n13334;
  assign n13336 = ~n13331 & n13335;
  assign n13337 = pi788 & ~n13336;
  assign n13338 = pi788 & ~n13330;
  assign n13339 = ~n13336 & n13338;
  assign n13340 = ~n13330 & n13337;
  assign n13341 = ~n63030 & ~n63118;
  assign n13342 = ~n13321 & n13341;
  assign n13343 = ~n8595 & ~n63011;
  assign n13344 = n63013 & n13343;
  assign n13345 = ~n8595 & n13325;
  assign n13346 = n13227 & n13344;
  assign n13347 = ~pi629 & n63119;
  assign n13348 = pi628 & ~n13347;
  assign n13349 = ~n8303 & n13322;
  assign n13350 = n10207 & n13254;
  assign n13351 = pi629 & ~n63120;
  assign n13352 = ~pi628 & n63120;
  assign n13353 = pi629 & ~n13352;
  assign n13354 = pi628 & ~n63119;
  assign n13355 = ~n13353 & ~n13354;
  assign n13356 = ~n13348 & ~n13351;
  assign n13357 = ~pi1156 & ~n63121;
  assign n13358 = pi628 & n63120;
  assign n13359 = ~pi628 & ~n63119;
  assign n13360 = pi629 & ~n13359;
  assign n13361 = pi1156 & ~n13360;
  assign n13362 = ~n13358 & n13361;
  assign n13363 = ~n13357 & ~n13362;
  assign n13364 = pi792 & ~n13226;
  assign n13365 = ~n13363 & n13364;
  assign n13366 = ~n13342 & ~n13365;
  assign n13367 = ~n8651 & ~n13366;
  assign n13368 = ~n62892 & n63120;
  assign n13369 = ~pi630 & ~n13368;
  assign n13370 = pi647 & ~n13369;
  assign n13371 = ~n8334 & n63119;
  assign n13372 = pi630 & n13371;
  assign n13373 = pi1157 & ~n13372;
  assign n13374 = ~n13370 & n13373;
  assign n13375 = pi630 & ~n13368;
  assign n13376 = ~pi647 & ~n13375;
  assign n13377 = ~pi630 & n13371;
  assign n13378 = ~pi1157 & ~n13377;
  assign n13379 = pi647 & ~n13377;
  assign n13380 = ~pi647 & n13368;
  assign n13381 = pi630 & ~n13380;
  assign n13382 = pi647 & ~n13371;
  assign n13383 = ~n13381 & ~n13382;
  assign n13384 = ~n13375 & ~n13379;
  assign n13385 = ~pi1157 & ~n63122;
  assign n13386 = ~n13376 & n13378;
  assign n13387 = ~n13374 & ~n63123;
  assign n13388 = pi787 & ~n13226;
  assign n13389 = ~n13387 & n13388;
  assign n13390 = ~n11547 & ~n13389;
  assign n13391 = ~n13367 & n13390;
  assign n13392 = n11556 & n13368;
  assign n13393 = n63013 & n11558;
  assign n13394 = n8685 & n63119;
  assign n13395 = n13282 & n13393;
  assign n13396 = ~pi1160 & n63124;
  assign n13397 = ~n13226 & ~n13396;
  assign n13398 = n11540 & ~n13397;
  assign n13399 = pi1160 & n63124;
  assign n13400 = ~n13226 & ~n13399;
  assign n13401 = n11542 & ~n13400;
  assign n13402 = ~n13398 & ~n13401;
  assign n13403 = ~n13392 & n13402;
  assign n13404 = pi790 & ~n13403;
  assign n13405 = pi832 & ~n13404;
  assign n13406 = ~n13367 & ~n13389;
  assign n13407 = pi644 & n13406;
  assign n13408 = ~n10298 & n13368;
  assign n13409 = ~n13226 & ~n13408;
  assign n13410 = ~pi644 & ~n13409;
  assign n13411 = pi715 & ~n13410;
  assign n13412 = ~n13407 & n13411;
  assign n13413 = pi644 & n11558;
  assign n13414 = pi644 & n63124;
  assign n13415 = n13325 & n13413;
  assign n13416 = ~pi715 & ~n13226;
  assign n13417 = ~n63125 & n13416;
  assign n13418 = pi1160 & ~n13417;
  assign n13419 = ~n13412 & n13418;
  assign n13420 = ~pi644 & n13406;
  assign n13421 = pi644 & ~n13409;
  assign n13422 = ~pi715 & ~n13421;
  assign n13423 = ~n13420 & n13422;
  assign n13424 = ~pi644 & n11558;
  assign n13425 = ~pi644 & n63124;
  assign n13426 = n13325 & n13424;
  assign n13427 = pi715 & ~n13226;
  assign n13428 = ~n63126 & n13427;
  assign n13429 = ~pi1160 & ~n13428;
  assign n13430 = ~n13423 & n13429;
  assign n13431 = ~n13419 & ~n13430;
  assign n13432 = pi790 & ~n13431;
  assign n13433 = ~pi790 & n13406;
  assign n13434 = pi832 & ~n13433;
  assign n13435 = ~n13432 & n13434;
  assign n13436 = ~n13391 & n13405;
  assign po331 = ~n13219 & ~n63127;
  assign n13438 = ~pi175 & ~n2923;
  assign n13439 = pi766 & n7316;
  assign n13440 = ~n13438 & ~n13439;
  assign n13441 = ~n8420 & ~n13440;
  assign n13442 = ~pi785 & ~n13441;
  assign n13443 = n8148 & n13439;
  assign n13444 = n13441 & ~n13443;
  assign n13445 = pi1155 & ~n13444;
  assign n13446 = ~pi1155 & ~n13438;
  assign n13447 = ~n13443 & n13446;
  assign n13448 = ~n13445 & ~n13447;
  assign n13449 = pi785 & ~n13448;
  assign n13450 = ~n13442 & ~n13449;
  assign n13451 = ~pi781 & ~n13450;
  assign n13452 = ~n8435 & n13450;
  assign n13453 = pi1154 & ~n13452;
  assign n13454 = ~n8438 & n13450;
  assign n13455 = ~pi1154 & ~n13454;
  assign n13456 = ~n13453 & ~n13455;
  assign n13457 = pi781 & ~n13456;
  assign n13458 = ~n13451 & ~n13457;
  assign n13459 = ~pi789 & ~n13458;
  assign n13460 = ~pi1159 & ~n12615;
  assign n13461 = n13458 & n13460;
  assign n13462 = pi1159 & ~n12612;
  assign n13463 = n13458 & n13462;
  assign n13464 = pi789 & ~n13463;
  assign n13465 = ~n12612 & n13458;
  assign n13466 = pi1159 & ~n13465;
  assign n13467 = ~n12615 & n13458;
  assign n13468 = ~pi1159 & ~n13467;
  assign n13469 = ~n13466 & ~n13468;
  assign n13470 = pi789 & ~n13469;
  assign n13471 = ~n13461 & n13464;
  assign n13472 = ~n13459 & ~n63128;
  assign n13473 = ~n8595 & n13472;
  assign n13474 = n8595 & n13438;
  assign n13475 = ~n8595 & ~n13472;
  assign n13476 = n8595 & ~n13438;
  assign n13477 = ~n13475 & ~n13476;
  assign n13478 = ~n13473 & ~n13474;
  assign n13479 = ~n8334 & n63129;
  assign n13480 = n8334 & n13438;
  assign n13481 = ~n8413 & ~n13480;
  assign n13482 = ~n13479 & ~n13480;
  assign n13483 = ~n8413 & n13482;
  assign n13484 = ~n13479 & n13481;
  assign n13485 = pi700 & n7564;
  assign n13486 = ~n13438 & ~n13485;
  assign n13487 = ~pi778 & ~n13486;
  assign n13488 = ~pi625 & n13485;
  assign n13489 = ~n13486 & ~n13488;
  assign n13490 = pi1153 & ~n13489;
  assign n13491 = ~pi1153 & ~n13438;
  assign n13492 = ~n13488 & n13491;
  assign n13493 = pi778 & ~n13492;
  assign n13494 = ~n13490 & n13493;
  assign n13495 = ~n13487 & ~n13494;
  assign n13496 = ~n8490 & ~n13495;
  assign n13497 = ~n8492 & n13496;
  assign n13498 = ~n8494 & n13497;
  assign n13499 = ~n8496 & n13498;
  assign n13500 = ~n8508 & n13499;
  assign n13501 = pi647 & ~n13500;
  assign n13502 = ~pi647 & ~n13438;
  assign n13503 = ~n13501 & ~n13502;
  assign n13504 = n8373 & ~n13503;
  assign n13505 = ~pi647 & n13500;
  assign n13506 = pi647 & n13438;
  assign n13507 = ~pi1157 & ~n13506;
  assign n13508 = ~n13505 & n13507;
  assign n13509 = pi630 & n13508;
  assign n13510 = ~n13504 & ~n13509;
  assign n13511 = ~n63130 & n13510;
  assign n13512 = pi787 & ~n13511;
  assign n13513 = ~pi626 & ~n13472;
  assign n13514 = pi626 & ~n13438;
  assign n13515 = n8301 & ~n13514;
  assign n13516 = ~n13513 & n13515;
  assign n13517 = n8525 & n13498;
  assign n13518 = pi626 & ~n13472;
  assign n13519 = ~pi626 & ~n13438;
  assign n13520 = n8300 & ~n13519;
  assign n13521 = ~n13518 & n13520;
  assign n13522 = ~n13517 & ~n13521;
  assign n13523 = ~n13516 & ~n13517;
  assign n13524 = ~n13521 & n13523;
  assign n13525 = ~n13516 & n13522;
  assign n13526 = pi788 & ~n63131;
  assign n13527 = n11303 & n13497;
  assign n13528 = pi648 & ~n13527;
  assign n13529 = ~n13461 & n13528;
  assign n13530 = n11304 & n13497;
  assign n13531 = ~pi648 & ~n13530;
  assign n13532 = ~n13463 & n13531;
  assign n13533 = pi789 & ~n13532;
  assign n13534 = ~n13529 & n13533;
  assign n13535 = ~n7187 & ~n13486;
  assign n13536 = pi625 & n13535;
  assign n13537 = n13440 & ~n13535;
  assign n13538 = ~n13536 & ~n13537;
  assign n13539 = n13491 & ~n13538;
  assign n13540 = ~pi608 & ~n13490;
  assign n13541 = ~n13539 & n13540;
  assign n13542 = pi1153 & n13440;
  assign n13543 = ~n13536 & n13542;
  assign n13544 = pi608 & ~n13492;
  assign n13545 = ~n13543 & n13544;
  assign n13546 = ~n13541 & ~n13545;
  assign n13547 = pi778 & ~n13546;
  assign n13548 = ~pi778 & ~n13537;
  assign n13549 = ~n13547 & ~n13548;
  assign n13550 = ~pi609 & ~n13549;
  assign n13551 = pi609 & ~n13495;
  assign n13552 = ~pi1155 & ~n13551;
  assign n13553 = ~n13550 & n13552;
  assign n13554 = ~pi660 & ~n13445;
  assign n13555 = ~n13553 & n13554;
  assign n13556 = pi609 & ~n13549;
  assign n13557 = ~pi609 & ~n13495;
  assign n13558 = pi1155 & ~n13557;
  assign n13559 = ~n13556 & n13558;
  assign n13560 = pi660 & ~n13447;
  assign n13561 = ~n13559 & n13560;
  assign n13562 = ~n13555 & ~n13561;
  assign n13563 = pi785 & ~n13562;
  assign n13564 = ~pi785 & ~n13549;
  assign n13565 = ~n13563 & ~n13564;
  assign n13566 = pi618 & ~n13565;
  assign n13567 = ~pi618 & n13496;
  assign n13568 = pi1154 & ~n13567;
  assign n13569 = ~n13566 & n13568;
  assign n13570 = pi627 & ~n13455;
  assign n13571 = ~n13569 & n13570;
  assign n13572 = ~pi618 & ~n13565;
  assign n13573 = pi618 & n13496;
  assign n13574 = ~pi1154 & ~n13573;
  assign n13575 = ~n13572 & n13574;
  assign n13576 = ~pi627 & ~n13453;
  assign n13577 = ~n13575 & n13576;
  assign n13578 = pi781 & ~n13577;
  assign n13579 = ~n13571 & n13578;
  assign n13580 = ~pi781 & n13565;
  assign n13581 = ~n11434 & ~n13580;
  assign n13582 = ~n13579 & n13581;
  assign n13583 = ~n13534 & ~n13582;
  assign n13584 = ~n13571 & ~n13577;
  assign n13585 = pi781 & ~n13584;
  assign n13586 = ~pi781 & ~n13565;
  assign n13587 = ~n13585 & ~n13586;
  assign n13588 = ~pi619 & ~n13587;
  assign n13589 = pi619 & n13497;
  assign n13590 = ~pi1159 & ~n13589;
  assign n13591 = ~n13588 & n13590;
  assign n13592 = ~pi648 & ~n13466;
  assign n13593 = ~n13591 & n13592;
  assign n13594 = pi619 & ~n13587;
  assign n13595 = ~pi619 & n13497;
  assign n13596 = pi1159 & ~n13595;
  assign n13597 = ~n13594 & n13596;
  assign n13598 = pi648 & ~n13468;
  assign n13599 = ~n13597 & n13598;
  assign n13600 = pi789 & ~n13599;
  assign n13601 = pi789 & ~n13593;
  assign n13602 = ~n13599 & n13601;
  assign n13603 = ~n13593 & n13600;
  assign n13604 = ~pi789 & n13587;
  assign n13605 = n62894 & ~n13604;
  assign n13606 = ~n63132 & n13605;
  assign n13607 = n62894 & ~n13583;
  assign n13608 = ~n13526 & ~n63133;
  assign n13609 = ~n63030 & ~n13608;
  assign n13610 = n8498 & n63129;
  assign n13611 = n8615 & n13499;
  assign n13612 = pi629 & ~n13611;
  assign n13613 = ~n13610 & n13612;
  assign n13614 = n8499 & n63129;
  assign n13615 = n8606 & n13499;
  assign n13616 = ~pi629 & ~n13615;
  assign n13617 = ~n13614 & n13616;
  assign n13618 = pi792 & ~n13617;
  assign n13619 = pi792 & ~n13613;
  assign n13620 = ~n13617 & n13619;
  assign n13621 = ~n13614 & ~n13615;
  assign n13622 = ~pi629 & ~n13621;
  assign n13623 = ~n13610 & ~n13611;
  assign n13624 = pi629 & ~n13623;
  assign n13625 = ~n13622 & ~n13624;
  assign n13626 = pi792 & ~n13625;
  assign n13627 = ~n13613 & n13618;
  assign n13628 = ~n8651 & ~n63134;
  assign n13629 = ~n13609 & n13628;
  assign n13630 = ~n13512 & ~n13629;
  assign n13631 = pi644 & n13630;
  assign n13632 = ~pi787 & ~n13500;
  assign n13633 = pi1157 & ~n13503;
  assign n13634 = ~n13508 & ~n13633;
  assign n13635 = pi787 & ~n13634;
  assign n13636 = ~n13632 & ~n13635;
  assign n13637 = ~pi644 & n13636;
  assign n13638 = pi715 & ~n13637;
  assign n13639 = ~n13631 & n13638;
  assign n13640 = ~n8685 & n13438;
  assign n13641 = ~n8376 & n13479;
  assign n13642 = ~n8376 & ~n13482;
  assign n13643 = n8376 & n13438;
  assign n13644 = ~n13642 & ~n13643;
  assign n13645 = ~n13640 & ~n13641;
  assign n13646 = pi644 & ~n63135;
  assign n13647 = ~pi644 & n13438;
  assign n13648 = ~pi715 & ~n13647;
  assign n13649 = ~n13646 & n13648;
  assign n13650 = pi1160 & ~n13649;
  assign n13651 = ~n13639 & n13650;
  assign n13652 = ~pi644 & n13630;
  assign n13653 = pi644 & n13636;
  assign n13654 = ~pi715 & ~n13653;
  assign n13655 = ~n13652 & n13654;
  assign n13656 = ~pi644 & ~n63135;
  assign n13657 = pi644 & n13438;
  assign n13658 = pi715 & ~n13657;
  assign n13659 = ~n13656 & n13658;
  assign n13660 = ~pi1160 & ~n13659;
  assign n13661 = ~n13655 & n13660;
  assign n13662 = ~n13651 & ~n13661;
  assign n13663 = pi790 & ~n13662;
  assign n13664 = ~pi790 & n13630;
  assign n13665 = pi832 & ~n13664;
  assign n13666 = ~n13663 & n13665;
  assign n13667 = ~pi175 & ~n8098;
  assign n13668 = ~n11558 & n13667;
  assign n13669 = pi175 & ~n62765;
  assign n13670 = ~pi766 & n7143;
  assign n13671 = pi175 & n7349;
  assign n13672 = ~n13670 & ~n13671;
  assign n13673 = pi39 & ~n13672;
  assign n13674 = ~pi175 & pi766;
  assign n13675 = n62802 & n13674;
  assign n13676 = ~pi766 & n6946;
  assign n13677 = pi766 & ~n7293;
  assign n13678 = pi175 & ~n13677;
  assign n13679 = ~n13676 & ~n13678;
  assign n13680 = ~n13675 & n13679;
  assign n13681 = ~n13673 & n13680;
  assign n13682 = ~pi38 & ~n13681;
  assign n13683 = pi766 & n7359;
  assign n13684 = ~pi175 & ~n7357;
  assign n13685 = pi38 & ~n13684;
  assign n13686 = ~n13683 & n13685;
  assign n13687 = ~n13682 & ~n13686;
  assign n13688 = n62765 & ~n13687;
  assign n13689 = ~n13669 & ~n13688;
  assign n13690 = ~n8135 & ~n13689;
  assign n13691 = n8135 & ~n13667;
  assign n13692 = ~n13690 & ~n13691;
  assign n13693 = ~pi785 & ~n13692;
  assign n13694 = ~n8136 & ~n13667;
  assign n13695 = pi609 & n13690;
  assign n13696 = ~n13694 & ~n13695;
  assign n13697 = pi1155 & ~n13696;
  assign n13698 = ~n8148 & ~n13667;
  assign n13699 = ~pi609 & n13690;
  assign n13700 = ~n13698 & ~n13699;
  assign n13701 = ~pi1155 & ~n13700;
  assign n13702 = ~n13697 & ~n13701;
  assign n13703 = pi785 & ~n13702;
  assign n13704 = ~n13693 & ~n13703;
  assign n13705 = ~pi781 & ~n13704;
  assign n13706 = pi618 & n13704;
  assign n13707 = ~pi618 & n13667;
  assign n13708 = pi1154 & ~n13707;
  assign n13709 = ~n13706 & n13708;
  assign n13710 = ~pi618 & n13704;
  assign n13711 = pi618 & n13667;
  assign n13712 = ~pi1154 & ~n13711;
  assign n13713 = ~n13710 & n13712;
  assign n13714 = ~n13709 & ~n13713;
  assign n13715 = pi781 & ~n13714;
  assign n13716 = ~n13705 & ~n13715;
  assign n13717 = ~pi619 & ~n13716;
  assign n13718 = pi619 & ~n13667;
  assign n13719 = ~pi1159 & ~n13718;
  assign n13720 = ~n13717 & n13719;
  assign n13721 = pi619 & ~n13716;
  assign n13722 = ~pi619 & ~n13667;
  assign n13723 = pi1159 & ~n13722;
  assign n13724 = ~n13721 & n13723;
  assign n13725 = pi619 & n13716;
  assign n13726 = ~pi619 & n13667;
  assign n13727 = pi1159 & ~n13726;
  assign n13728 = ~n13725 & n13727;
  assign n13729 = ~pi619 & n13716;
  assign n13730 = pi619 & n13667;
  assign n13731 = ~pi1159 & ~n13730;
  assign n13732 = ~n13729 & n13731;
  assign n13733 = ~n13728 & ~n13732;
  assign n13734 = ~n13720 & ~n13724;
  assign n13735 = pi789 & n63136;
  assign n13736 = ~pi789 & n13716;
  assign n13737 = ~pi789 & ~n13716;
  assign n13738 = pi789 & ~n63136;
  assign n13739 = ~n13737 & ~n13738;
  assign n13740 = ~n13735 & ~n13736;
  assign n13741 = ~n8595 & n63137;
  assign n13742 = n8685 & n13741;
  assign n13743 = n8376 & ~n13667;
  assign n13744 = n8595 & n13667;
  assign n13745 = ~n13741 & ~n13744;
  assign n13746 = ~n8334 & ~n13745;
  assign n13747 = n8334 & n13667;
  assign n13748 = ~n13746 & ~n13747;
  assign n13749 = ~n8376 & n13748;
  assign n13750 = ~n13743 & ~n13749;
  assign n13751 = ~n8376 & ~n13748;
  assign n13752 = n8376 & n13667;
  assign n13753 = ~n13751 & ~n13752;
  assign n13754 = ~n13668 & ~n13742;
  assign n13755 = pi644 & n63138;
  assign n13756 = ~pi644 & n13667;
  assign n13757 = ~pi715 & ~n13756;
  assign n13758 = ~n13755 & n13757;
  assign n13759 = n10298 & ~n13667;
  assign n13760 = n8257 & ~n13667;
  assign n13761 = ~pi175 & n8009;
  assign n13762 = pi175 & n62874;
  assign n13763 = ~pi38 & ~n13762;
  assign n13764 = ~n13761 & n13763;
  assign n13765 = n8085 & ~n13684;
  assign n13766 = pi700 & ~n13765;
  assign n13767 = ~n13764 & n13766;
  assign n13768 = ~pi175 & ~pi700;
  assign n13769 = ~n8091 & n13768;
  assign n13770 = n62765 & ~n13769;
  assign n13771 = ~n13767 & n13770;
  assign n13772 = ~n13669 & ~n13771;
  assign n13773 = ~pi778 & ~n13772;
  assign n13774 = pi625 & n13772;
  assign n13775 = ~pi625 & n13667;
  assign n13776 = pi1153 & ~n13775;
  assign n13777 = ~n13774 & n13776;
  assign n13778 = ~pi625 & n13772;
  assign n13779 = pi625 & n13667;
  assign n13780 = ~pi1153 & ~n13779;
  assign n13781 = ~n13778 & n13780;
  assign n13782 = ~n13777 & ~n13781;
  assign n13783 = pi778 & ~n13782;
  assign n13784 = ~n13773 & ~n13783;
  assign n13785 = ~n62880 & ~n13784;
  assign n13786 = n62880 & ~n13667;
  assign n13787 = ~n62880 & n13784;
  assign n13788 = n62880 & n13667;
  assign n13789 = ~n13787 & ~n13788;
  assign n13790 = ~n13785 & ~n13786;
  assign n13791 = ~n62882 & ~n63139;
  assign n13792 = n62882 & n13667;
  assign n13793 = n62882 & ~n13667;
  assign n13794 = ~n62882 & n63139;
  assign n13795 = ~n13793 & ~n13794;
  assign n13796 = ~n13791 & ~n13792;
  assign n13797 = ~n8257 & ~n63140;
  assign n13798 = ~n8257 & n63140;
  assign n13799 = n8257 & n13667;
  assign n13800 = ~n13798 & ~n13799;
  assign n13801 = ~n13760 & ~n13797;
  assign n13802 = ~n8303 & ~n63141;
  assign n13803 = n8303 & n13667;
  assign n13804 = ~n13802 & ~n13803;
  assign n13805 = ~n62892 & ~n13804;
  assign n13806 = n62892 & n13667;
  assign n13807 = n62892 & ~n13667;
  assign n13808 = ~n62892 & n13804;
  assign n13809 = ~n13807 & ~n13808;
  assign n13810 = ~pi628 & ~n13804;
  assign n13811 = pi628 & n13667;
  assign n13812 = ~n13810 & ~n13811;
  assign n13813 = ~pi1156 & ~n13812;
  assign n13814 = pi628 & ~n13804;
  assign n13815 = ~pi628 & n13667;
  assign n13816 = ~n13814 & ~n13815;
  assign n13817 = pi1156 & ~n13816;
  assign n13818 = ~n13813 & ~n13817;
  assign n13819 = pi792 & ~n13818;
  assign n13820 = ~pi792 & ~n13804;
  assign n13821 = ~n13819 & ~n13820;
  assign n13822 = ~n13805 & ~n13806;
  assign n13823 = ~n10298 & ~n63142;
  assign n13824 = ~n10298 & n63142;
  assign n13825 = n10298 & n13667;
  assign n13826 = ~n13824 & ~n13825;
  assign n13827 = ~pi647 & n63142;
  assign n13828 = pi647 & n13667;
  assign n13829 = ~n13827 & ~n13828;
  assign n13830 = ~pi1157 & ~n13829;
  assign n13831 = pi647 & n63142;
  assign n13832 = ~pi647 & n13667;
  assign n13833 = ~n13831 & ~n13832;
  assign n13834 = pi1157 & ~n13833;
  assign n13835 = ~n13830 & ~n13834;
  assign n13836 = pi787 & ~n13835;
  assign n13837 = ~pi787 & n63142;
  assign n13838 = ~n13836 & ~n13837;
  assign n13839 = ~n13759 & ~n13823;
  assign n13840 = ~pi644 & ~n63143;
  assign n13841 = pi715 & ~n13840;
  assign n13842 = pi1160 & ~n13841;
  assign n13843 = pi1160 & ~n13758;
  assign n13844 = ~n13841 & n13843;
  assign n13845 = ~n13758 & n13842;
  assign n13846 = pi644 & ~n63143;
  assign n13847 = ~pi715 & ~n13846;
  assign n13848 = ~pi644 & n63138;
  assign n13849 = pi644 & n13667;
  assign n13850 = pi715 & ~n13849;
  assign n13851 = ~n13848 & n13850;
  assign n13852 = ~pi1160 & ~n13851;
  assign n13853 = ~n13847 & n13852;
  assign n13854 = ~n63144 & ~n13853;
  assign n13855 = pi790 & ~n13854;
  assign n13856 = ~n63052 & n13745;
  assign n13857 = n8332 & ~n13811;
  assign n13858 = n8332 & n13812;
  assign n13859 = ~n13810 & n13857;
  assign n13860 = n8331 & ~n13815;
  assign n13861 = n8331 & n13816;
  assign n13862 = ~n13814 & n13860;
  assign n13863 = ~n63145 & ~n63146;
  assign n13864 = ~n13856 & n13863;
  assign n13865 = pi792 & ~n13864;
  assign n13866 = ~pi700 & n13687;
  assign n13867 = ~pi175 & ~n62821;
  assign n13868 = pi175 & n7632;
  assign n13869 = ~pi766 & ~n13868;
  assign n13870 = ~n13867 & n13869;
  assign n13871 = pi175 & n7709;
  assign n13872 = ~pi175 & n62851;
  assign n13873 = pi766 & ~n13872;
  assign n13874 = ~n13871 & n13873;
  assign n13875 = pi39 & ~n13874;
  assign n13876 = ~n13870 & n13875;
  assign n13877 = ~pi175 & n7832;
  assign n13878 = pi175 & n7855;
  assign n13879 = ~pi766 & ~n13878;
  assign n13880 = ~pi766 & ~n13877;
  assign n13881 = ~n13878 & n13880;
  assign n13882 = ~n13877 & n13879;
  assign n13883 = ~pi175 & ~n7861;
  assign n13884 = pi175 & ~n7868;
  assign n13885 = pi766 & ~n13884;
  assign n13886 = ~n13883 & n13885;
  assign n13887 = ~pi39 & ~n13886;
  assign n13888 = ~n63147 & n13887;
  assign n13889 = ~pi38 & ~n13888;
  assign n13890 = ~pi175 & n8759;
  assign n13891 = pi175 & n8763;
  assign n13892 = ~pi766 & ~n13891;
  assign n13893 = ~n13890 & n13892;
  assign n13894 = pi175 & n8775;
  assign n13895 = ~pi175 & ~n8779;
  assign n13896 = pi766 & ~n13895;
  assign n13897 = ~n13894 & n13896;
  assign n13898 = ~n13893 & ~n13897;
  assign n13899 = ~pi38 & ~n13898;
  assign n13900 = ~n13876 & n13889;
  assign n13901 = n6955 & ~n7367;
  assign n13902 = ~pi766 & n13901;
  assign n13903 = ~n7744 & ~n13902;
  assign n13904 = ~pi39 & ~n13903;
  assign n13905 = ~pi175 & ~n13904;
  assign n13906 = ~n7565 & ~n13439;
  assign n13907 = pi175 & ~n13906;
  assign n13908 = n7356 & n13907;
  assign n13909 = pi38 & ~n13908;
  assign n13910 = ~n13905 & n13909;
  assign n13911 = pi700 & ~n13910;
  assign n13912 = ~n63148 & n13911;
  assign n13913 = n62765 & ~n13912;
  assign n13914 = n62765 & ~n13866;
  assign n13915 = ~n13912 & n13914;
  assign n13916 = ~n13866 & n13913;
  assign n13917 = ~n13669 & ~n63149;
  assign n13918 = ~pi625 & n13917;
  assign n13919 = pi625 & n13689;
  assign n13920 = ~pi1153 & ~n13919;
  assign n13921 = ~n13918 & n13920;
  assign n13922 = ~pi608 & ~n13777;
  assign n13923 = ~n13921 & n13922;
  assign n13924 = pi625 & n13917;
  assign n13925 = ~pi625 & n13689;
  assign n13926 = pi1153 & ~n13925;
  assign n13927 = ~n13924 & n13926;
  assign n13928 = pi608 & ~n13781;
  assign n13929 = ~n13927 & n13928;
  assign n13930 = ~n13923 & ~n13929;
  assign n13931 = pi778 & ~n13930;
  assign n13932 = ~pi778 & n13917;
  assign n13933 = ~n13931 & ~n13932;
  assign n13934 = ~pi609 & ~n13933;
  assign n13935 = pi609 & n13784;
  assign n13936 = ~pi1155 & ~n13935;
  assign n13937 = ~n13934 & n13936;
  assign n13938 = ~pi660 & ~n13697;
  assign n13939 = ~n13937 & n13938;
  assign n13940 = pi609 & ~n13933;
  assign n13941 = ~pi609 & n13784;
  assign n13942 = pi1155 & ~n13941;
  assign n13943 = ~n13940 & n13942;
  assign n13944 = pi660 & ~n13701;
  assign n13945 = ~n13943 & n13944;
  assign n13946 = ~n13939 & ~n13945;
  assign n13947 = pi785 & ~n13946;
  assign n13948 = ~pi785 & ~n13933;
  assign n13949 = ~n13947 & ~n13948;
  assign n13950 = ~pi781 & n13949;
  assign n13951 = ~pi618 & ~n13949;
  assign n13952 = pi618 & ~n63139;
  assign n13953 = ~pi1154 & ~n13952;
  assign n13954 = ~n13951 & n13953;
  assign n13955 = ~pi627 & ~n13709;
  assign n13956 = ~n13954 & n13955;
  assign n13957 = pi618 & ~n13949;
  assign n13958 = ~pi618 & ~n63139;
  assign n13959 = pi1154 & ~n13958;
  assign n13960 = ~n13957 & n13959;
  assign n13961 = pi627 & ~n13713;
  assign n13962 = ~n13960 & n13961;
  assign n13963 = pi781 & ~n13962;
  assign n13964 = ~n13956 & n13963;
  assign n13965 = ~n13956 & ~n13962;
  assign n13966 = pi781 & ~n13965;
  assign n13967 = ~pi781 & ~n13949;
  assign n13968 = ~n13966 & ~n13967;
  assign n13969 = ~n13950 & ~n13964;
  assign n13970 = ~n11434 & n63150;
  assign n13971 = ~n11431 & ~n63140;
  assign n13972 = ~n62884 & ~n63136;
  assign n13973 = ~n13971 & ~n13972;
  assign n13974 = pi789 & ~n13973;
  assign n13975 = n62894 & ~n13974;
  assign n13976 = ~pi619 & ~n63150;
  assign n13977 = pi619 & n63140;
  assign n13978 = ~pi1159 & ~n13977;
  assign n13979 = ~n13976 & n13978;
  assign n13980 = ~pi648 & ~n13728;
  assign n13981 = ~n13979 & n13980;
  assign n13982 = pi619 & ~n63150;
  assign n13983 = ~pi619 & n63140;
  assign n13984 = pi1159 & ~n13983;
  assign n13985 = ~n13982 & n13984;
  assign n13986 = pi648 & ~n13732;
  assign n13987 = ~n13985 & n13986;
  assign n13988 = pi789 & ~n13987;
  assign n13989 = pi789 & ~n13981;
  assign n13990 = ~n13987 & n13989;
  assign n13991 = ~n13981 & n13988;
  assign n13992 = ~pi789 & n63150;
  assign n13993 = n62894 & ~n13992;
  assign n13994 = ~n63151 & n13993;
  assign n13995 = ~n13970 & n13975;
  assign n13996 = ~pi626 & ~n63137;
  assign n13997 = pi626 & ~n13667;
  assign n13998 = n8301 & ~n13997;
  assign n13999 = ~n13996 & n13998;
  assign n14000 = n8525 & ~n63141;
  assign n14001 = pi626 & ~n63137;
  assign n14002 = ~pi626 & ~n13667;
  assign n14003 = n8300 & ~n14002;
  assign n14004 = ~n14001 & n14003;
  assign n14005 = ~n14000 & ~n14004;
  assign n14006 = ~n13999 & ~n14000;
  assign n14007 = ~n14004 & n14006;
  assign n14008 = ~n13999 & n14005;
  assign n14009 = pi788 & ~n63153;
  assign n14010 = ~n63030 & ~n14009;
  assign n14011 = ~n63152 & n14010;
  assign n14012 = ~n13865 & ~n14011;
  assign n14013 = ~n8651 & ~n14012;
  assign n14014 = ~n8413 & ~n13747;
  assign n14015 = ~n8413 & n13748;
  assign n14016 = ~n13746 & n14014;
  assign n14017 = n8374 & ~n13828;
  assign n14018 = n8374 & n13829;
  assign n14019 = ~n13827 & n14017;
  assign n14020 = n8373 & ~n13832;
  assign n14021 = n8373 & n13833;
  assign n14022 = ~n13831 & n14020;
  assign n14023 = ~n63155 & ~n63156;
  assign n14024 = ~n63154 & ~n63155;
  assign n14025 = ~n63156 & n14024;
  assign n14026 = ~n63154 & n14023;
  assign n14027 = pi787 & ~n63157;
  assign n14028 = ~pi644 & n13852;
  assign n14029 = pi644 & pi1160;
  assign n14030 = pi644 & n13843;
  assign n14031 = ~n13758 & n14029;
  assign n14032 = pi790 & ~n63158;
  assign n14033 = pi790 & ~n14028;
  assign n14034 = ~n63158 & n14033;
  assign n14035 = ~n14028 & n14032;
  assign n14036 = ~n14027 & ~n63159;
  assign n14037 = ~n14013 & ~n14027;
  assign n14038 = ~n63159 & n14037;
  assign n14039 = ~n14013 & n14036;
  assign n14040 = ~n13855 & ~n63160;
  assign n14041 = n62455 & ~n14040;
  assign n14042 = ~pi175 & ~n62455;
  assign n14043 = ~pi832 & ~n14042;
  assign n14044 = ~n14041 & n14043;
  assign po332 = ~n13666 & ~n14044;
  assign n14046 = ~pi176 & ~n2923;
  assign n14047 = ~pi742 & n7316;
  assign n14048 = ~n14046 & ~n14047;
  assign n14049 = ~n8420 & ~n14048;
  assign n14050 = ~pi785 & ~n14049;
  assign n14051 = ~n8425 & ~n14048;
  assign n14052 = pi1155 & ~n14051;
  assign n14053 = ~n8428 & n14049;
  assign n14054 = ~pi1155 & ~n14053;
  assign n14055 = ~n14052 & ~n14054;
  assign n14056 = pi785 & ~n14055;
  assign n14057 = ~n14050 & ~n14056;
  assign n14058 = ~pi781 & ~n14057;
  assign n14059 = ~n8435 & n14057;
  assign n14060 = pi1154 & ~n14059;
  assign n14061 = ~n8438 & n14057;
  assign n14062 = ~pi1154 & ~n14061;
  assign n14063 = ~n14060 & ~n14062;
  assign n14064 = pi781 & ~n14063;
  assign n14065 = ~n14058 & ~n14064;
  assign n14066 = ~pi619 & ~n14065;
  assign n14067 = pi619 & ~n14046;
  assign n14068 = ~pi1159 & ~n14067;
  assign n14069 = ~n14066 & n14068;
  assign n14070 = pi619 & ~n14065;
  assign n14071 = ~pi619 & ~n14046;
  assign n14072 = pi1159 & ~n14071;
  assign n14073 = ~n14070 & n14072;
  assign n14074 = pi619 & n14065;
  assign n14075 = ~pi619 & n14046;
  assign n14076 = pi1159 & ~n14075;
  assign n14077 = ~n14074 & n14076;
  assign n14078 = ~pi619 & n14065;
  assign n14079 = pi619 & n14046;
  assign n14080 = ~pi1159 & ~n14079;
  assign n14081 = ~n14078 & n14080;
  assign n14082 = ~n14077 & ~n14081;
  assign n14083 = ~n14069 & ~n14073;
  assign n14084 = pi789 & n63161;
  assign n14085 = ~pi789 & n14065;
  assign n14086 = ~pi789 & ~n14065;
  assign n14087 = pi789 & ~n63161;
  assign n14088 = ~n14086 & ~n14087;
  assign n14089 = ~n14084 & ~n14085;
  assign n14090 = ~n8595 & n63162;
  assign n14091 = n8595 & n14046;
  assign n14092 = ~n8595 & ~n63162;
  assign n14093 = n8595 & ~n14046;
  assign n14094 = ~n14092 & ~n14093;
  assign n14095 = ~n14090 & ~n14091;
  assign n14096 = ~n8334 & n63163;
  assign n14097 = n8334 & n14046;
  assign n14098 = ~n8413 & ~n14097;
  assign n14099 = ~n14096 & ~n14097;
  assign n14100 = ~n8413 & n14099;
  assign n14101 = ~n14096 & n14098;
  assign n14102 = ~pi704 & n7564;
  assign n14103 = ~n14046 & ~n14102;
  assign n14104 = ~pi778 & n14103;
  assign n14105 = ~pi625 & n14102;
  assign n14106 = ~n14103 & ~n14105;
  assign n14107 = pi1153 & ~n14106;
  assign n14108 = ~pi1153 & ~n14046;
  assign n14109 = ~n14105 & n14108;
  assign n14110 = ~n14107 & ~n14109;
  assign n14111 = pi778 & ~n14110;
  assign n14112 = ~n14104 & ~n14111;
  assign n14113 = ~n8490 & n14112;
  assign n14114 = ~n8492 & n14113;
  assign n14115 = ~n8494 & n14114;
  assign n14116 = ~n8496 & n14115;
  assign n14117 = ~n8508 & n14116;
  assign n14118 = pi647 & ~n14117;
  assign n14119 = ~pi647 & ~n14046;
  assign n14120 = ~n14118 & ~n14119;
  assign n14121 = n8373 & ~n14120;
  assign n14122 = ~pi647 & n14117;
  assign n14123 = pi647 & n14046;
  assign n14124 = ~pi1157 & ~n14123;
  assign n14125 = ~n14122 & n14124;
  assign n14126 = pi630 & n14125;
  assign n14127 = ~n14121 & ~n14126;
  assign n14128 = ~n63164 & n14127;
  assign n14129 = pi787 & ~n14128;
  assign n14130 = ~pi626 & ~n63162;
  assign n14131 = pi626 & ~n14046;
  assign n14132 = n8301 & ~n14131;
  assign n14133 = ~n14130 & n14132;
  assign n14134 = n8525 & n14115;
  assign n14135 = pi626 & ~n63162;
  assign n14136 = ~pi626 & ~n14046;
  assign n14137 = n8300 & ~n14136;
  assign n14138 = ~n14135 & n14137;
  assign n14139 = ~n14134 & ~n14138;
  assign n14140 = ~n14133 & ~n14134;
  assign n14141 = ~n14138 & n14140;
  assign n14142 = ~n14133 & n14139;
  assign n14143 = pi788 & ~n63165;
  assign n14144 = ~n7187 & ~n14103;
  assign n14145 = pi625 & n14144;
  assign n14146 = n14048 & ~n14144;
  assign n14147 = ~n14145 & ~n14146;
  assign n14148 = n14108 & ~n14147;
  assign n14149 = ~pi608 & ~n14107;
  assign n14150 = ~n14148 & n14149;
  assign n14151 = pi1153 & n14048;
  assign n14152 = ~n14145 & n14151;
  assign n14153 = pi608 & ~n14109;
  assign n14154 = ~n14152 & n14153;
  assign n14155 = ~n14150 & ~n14154;
  assign n14156 = pi778 & ~n14155;
  assign n14157 = ~pi778 & ~n14146;
  assign n14158 = ~n14156 & ~n14157;
  assign n14159 = ~pi609 & ~n14158;
  assign n14160 = pi609 & n14112;
  assign n14161 = ~pi1155 & ~n14160;
  assign n14162 = ~n14159 & n14161;
  assign n14163 = ~pi660 & ~n14052;
  assign n14164 = ~n14162 & n14163;
  assign n14165 = pi609 & ~n14158;
  assign n14166 = ~pi609 & n14112;
  assign n14167 = pi1155 & ~n14166;
  assign n14168 = ~n14165 & n14167;
  assign n14169 = pi660 & ~n14054;
  assign n14170 = ~n14168 & n14169;
  assign n14171 = ~n14164 & ~n14170;
  assign n14172 = pi785 & ~n14171;
  assign n14173 = ~pi785 & ~n14158;
  assign n14174 = ~n14172 & ~n14173;
  assign n14175 = pi618 & ~n14174;
  assign n14176 = ~pi618 & n14113;
  assign n14177 = pi1154 & ~n14176;
  assign n14178 = ~n14175 & n14177;
  assign n14179 = pi627 & ~n14062;
  assign n14180 = ~n14178 & n14179;
  assign n14181 = ~pi618 & ~n14174;
  assign n14182 = pi618 & n14113;
  assign n14183 = ~pi1154 & ~n14182;
  assign n14184 = ~n14181 & n14183;
  assign n14185 = ~pi627 & ~n14060;
  assign n14186 = ~n14184 & n14185;
  assign n14187 = pi781 & ~n14186;
  assign n14188 = ~n14180 & n14187;
  assign n14189 = ~n11431 & ~n14114;
  assign n14190 = ~n62884 & ~n63161;
  assign n14191 = ~n14189 & ~n14190;
  assign n14192 = pi789 & ~n14191;
  assign n14193 = ~pi781 & n14174;
  assign n14194 = ~n14192 & ~n14193;
  assign n14195 = ~n14188 & n14194;
  assign n14196 = n11434 & n14191;
  assign n14197 = ~n14195 & ~n14196;
  assign n14198 = ~n14180 & ~n14186;
  assign n14199 = pi781 & ~n14198;
  assign n14200 = ~pi781 & ~n14174;
  assign n14201 = ~n14199 & ~n14200;
  assign n14202 = ~pi619 & ~n14201;
  assign n14203 = pi619 & n14114;
  assign n14204 = ~pi1159 & ~n14203;
  assign n14205 = ~n14202 & n14204;
  assign n14206 = ~pi648 & ~n14077;
  assign n14207 = ~n14205 & n14206;
  assign n14208 = pi619 & ~n14201;
  assign n14209 = ~pi619 & n14114;
  assign n14210 = pi1159 & ~n14209;
  assign n14211 = ~n14208 & n14210;
  assign n14212 = pi648 & ~n14081;
  assign n14213 = ~n14211 & n14212;
  assign n14214 = pi789 & ~n14213;
  assign n14215 = pi789 & ~n14207;
  assign n14216 = ~n14213 & n14215;
  assign n14217 = ~n14207 & n14214;
  assign n14218 = ~pi789 & n14201;
  assign n14219 = n62894 & ~n14218;
  assign n14220 = ~n63166 & n14219;
  assign n14221 = n62894 & ~n14197;
  assign n14222 = ~n14143 & ~n63167;
  assign n14223 = ~n63030 & ~n14222;
  assign n14224 = n8498 & n63163;
  assign n14225 = n8615 & n14116;
  assign n14226 = pi629 & ~n14225;
  assign n14227 = ~n14224 & n14226;
  assign n14228 = n8499 & n63163;
  assign n14229 = n8606 & n14116;
  assign n14230 = ~pi629 & ~n14229;
  assign n14231 = ~n14228 & n14230;
  assign n14232 = pi792 & ~n14231;
  assign n14233 = pi792 & ~n14227;
  assign n14234 = ~n14231 & n14233;
  assign n14235 = ~n14228 & ~n14229;
  assign n14236 = ~pi629 & ~n14235;
  assign n14237 = ~n14224 & ~n14225;
  assign n14238 = pi629 & ~n14237;
  assign n14239 = ~n14236 & ~n14238;
  assign n14240 = pi792 & ~n14239;
  assign n14241 = ~n14227 & n14232;
  assign n14242 = ~n8651 & ~n63168;
  assign n14243 = ~n14223 & n14242;
  assign n14244 = ~n14129 & ~n14243;
  assign n14245 = pi644 & n14244;
  assign n14246 = ~pi787 & ~n14117;
  assign n14247 = pi1157 & ~n14120;
  assign n14248 = ~n14125 & ~n14247;
  assign n14249 = pi787 & ~n14248;
  assign n14250 = ~n14246 & ~n14249;
  assign n14251 = ~pi644 & n14250;
  assign n14252 = pi715 & ~n14251;
  assign n14253 = ~n14245 & n14252;
  assign n14254 = ~n8685 & n14046;
  assign n14255 = ~n8376 & n14096;
  assign n14256 = ~n8376 & ~n14099;
  assign n14257 = n8376 & n14046;
  assign n14258 = ~n14256 & ~n14257;
  assign n14259 = ~n14254 & ~n14255;
  assign n14260 = pi644 & ~n63169;
  assign n14261 = ~pi644 & n14046;
  assign n14262 = ~pi715 & ~n14261;
  assign n14263 = ~n14260 & n14262;
  assign n14264 = pi1160 & ~n14263;
  assign n14265 = ~n14253 & n14264;
  assign n14266 = ~pi644 & n14244;
  assign n14267 = pi644 & n14250;
  assign n14268 = ~pi715 & ~n14267;
  assign n14269 = ~n14266 & n14268;
  assign n14270 = ~pi644 & ~n63169;
  assign n14271 = pi644 & n14046;
  assign n14272 = pi715 & ~n14271;
  assign n14273 = ~n14270 & n14272;
  assign n14274 = ~pi1160 & ~n14273;
  assign n14275 = ~n14269 & n14274;
  assign n14276 = ~n14265 & ~n14275;
  assign n14277 = pi790 & ~n14276;
  assign n14278 = ~pi790 & n14244;
  assign n14279 = pi832 & ~n14278;
  assign n14280 = ~n14277 & n14279;
  assign n14281 = ~pi176 & ~n8098;
  assign n14282 = ~n11558 & n14281;
  assign n14283 = pi176 & ~n62765;
  assign n14284 = ~pi176 & n10343;
  assign n14285 = ~n62977 & ~n10339;
  assign n14286 = pi176 & n14285;
  assign n14287 = ~n14284 & ~n14286;
  assign n14288 = ~pi742 & ~n14287;
  assign n14289 = ~pi176 & ~n8091;
  assign n14290 = pi742 & ~n14289;
  assign n14291 = ~n14288 & ~n14290;
  assign n14292 = n62765 & ~n14291;
  assign n14293 = ~n14283 & ~n14292;
  assign n14294 = ~n8135 & ~n14293;
  assign n14295 = n8135 & ~n14281;
  assign n14296 = ~n14294 & ~n14295;
  assign n14297 = ~pi785 & ~n14296;
  assign n14298 = ~n8136 & ~n14281;
  assign n14299 = pi609 & n14294;
  assign n14300 = ~n14298 & ~n14299;
  assign n14301 = pi1155 & ~n14300;
  assign n14302 = ~n8148 & ~n14281;
  assign n14303 = ~pi609 & n14294;
  assign n14304 = ~n14302 & ~n14303;
  assign n14305 = ~pi1155 & ~n14304;
  assign n14306 = ~n14301 & ~n14305;
  assign n14307 = pi785 & ~n14306;
  assign n14308 = ~n14297 & ~n14307;
  assign n14309 = ~pi781 & ~n14308;
  assign n14310 = pi618 & n14308;
  assign n14311 = ~pi618 & n14281;
  assign n14312 = pi1154 & ~n14311;
  assign n14313 = ~n14310 & n14312;
  assign n14314 = ~pi618 & n14308;
  assign n14315 = pi618 & n14281;
  assign n14316 = ~pi1154 & ~n14315;
  assign n14317 = ~n14314 & n14316;
  assign n14318 = ~n14313 & ~n14317;
  assign n14319 = pi781 & ~n14318;
  assign n14320 = ~n14309 & ~n14319;
  assign n14321 = ~pi619 & ~n14320;
  assign n14322 = pi619 & ~n14281;
  assign n14323 = ~pi1159 & ~n14322;
  assign n14324 = ~n14321 & n14323;
  assign n14325 = pi619 & ~n14320;
  assign n14326 = ~pi619 & ~n14281;
  assign n14327 = pi1159 & ~n14326;
  assign n14328 = ~n14325 & n14327;
  assign n14329 = pi619 & n14320;
  assign n14330 = ~pi619 & n14281;
  assign n14331 = pi1159 & ~n14330;
  assign n14332 = ~n14329 & n14331;
  assign n14333 = ~pi619 & n14320;
  assign n14334 = pi619 & n14281;
  assign n14335 = ~pi1159 & ~n14334;
  assign n14336 = ~n14333 & n14335;
  assign n14337 = ~n14332 & ~n14336;
  assign n14338 = ~n14324 & ~n14328;
  assign n14339 = pi789 & n63170;
  assign n14340 = ~pi789 & n14320;
  assign n14341 = ~pi789 & ~n14320;
  assign n14342 = pi789 & ~n63170;
  assign n14343 = ~n14341 & ~n14342;
  assign n14344 = ~n14339 & ~n14340;
  assign n14345 = ~n8595 & n63171;
  assign n14346 = n8685 & n14345;
  assign n14347 = n8376 & ~n14281;
  assign n14348 = n8595 & n14281;
  assign n14349 = ~n14345 & ~n14348;
  assign n14350 = ~n8334 & ~n14349;
  assign n14351 = n8334 & n14281;
  assign n14352 = ~n14350 & ~n14351;
  assign n14353 = ~n8376 & n14352;
  assign n14354 = ~n14347 & ~n14353;
  assign n14355 = ~n8376 & ~n14352;
  assign n14356 = n8376 & n14281;
  assign n14357 = ~n14355 & ~n14356;
  assign n14358 = ~n14282 & ~n14346;
  assign n14359 = pi644 & n63172;
  assign n14360 = ~pi644 & n14281;
  assign n14361 = ~pi715 & ~n14360;
  assign n14362 = ~n14359 & n14361;
  assign n14363 = n10298 & ~n14281;
  assign n14364 = n8257 & ~n14281;
  assign n14365 = ~pi38 & ~n62874;
  assign n14366 = n62765 & ~n8085;
  assign n14367 = ~n14365 & n14366;
  assign n14368 = pi176 & ~n14367;
  assign n14369 = ~pi38 & n8009;
  assign n14370 = ~n10997 & ~n14369;
  assign n14371 = ~pi176 & n14370;
  assign n14372 = ~pi704 & ~n14371;
  assign n14373 = pi704 & n14289;
  assign n14374 = n62765 & ~n14373;
  assign n14375 = ~n14372 & n14374;
  assign n14376 = ~n14368 & ~n14375;
  assign n14377 = ~pi778 & ~n14376;
  assign n14378 = pi625 & n14376;
  assign n14379 = ~pi625 & n14281;
  assign n14380 = pi1153 & ~n14379;
  assign n14381 = ~n14378 & n14380;
  assign n14382 = ~pi625 & n14376;
  assign n14383 = pi625 & n14281;
  assign n14384 = ~pi1153 & ~n14383;
  assign n14385 = ~n14382 & n14384;
  assign n14386 = ~n14381 & ~n14385;
  assign n14387 = pi778 & ~n14386;
  assign n14388 = ~n14377 & ~n14387;
  assign n14389 = ~n62880 & ~n14388;
  assign n14390 = n62880 & ~n14281;
  assign n14391 = ~n62880 & n14388;
  assign n14392 = n62880 & n14281;
  assign n14393 = ~n14391 & ~n14392;
  assign n14394 = ~n14389 & ~n14390;
  assign n14395 = ~n62882 & ~n63173;
  assign n14396 = n62882 & n14281;
  assign n14397 = n62882 & ~n14281;
  assign n14398 = ~n62882 & n63173;
  assign n14399 = ~n14397 & ~n14398;
  assign n14400 = ~n14395 & ~n14396;
  assign n14401 = ~n8257 & ~n63174;
  assign n14402 = ~n8257 & n63174;
  assign n14403 = n8257 & n14281;
  assign n14404 = ~n14402 & ~n14403;
  assign n14405 = ~n14364 & ~n14401;
  assign n14406 = ~n8303 & ~n63175;
  assign n14407 = n8303 & n14281;
  assign n14408 = ~n14406 & ~n14407;
  assign n14409 = ~n62892 & ~n14408;
  assign n14410 = n62892 & n14281;
  assign n14411 = n62892 & ~n14281;
  assign n14412 = ~n62892 & n14408;
  assign n14413 = ~n14411 & ~n14412;
  assign n14414 = ~pi628 & ~n14408;
  assign n14415 = pi628 & n14281;
  assign n14416 = ~n14414 & ~n14415;
  assign n14417 = ~pi1156 & ~n14416;
  assign n14418 = pi628 & ~n14408;
  assign n14419 = ~pi628 & n14281;
  assign n14420 = ~n14418 & ~n14419;
  assign n14421 = pi1156 & ~n14420;
  assign n14422 = ~n14417 & ~n14421;
  assign n14423 = pi792 & ~n14422;
  assign n14424 = ~pi792 & ~n14408;
  assign n14425 = ~n14423 & ~n14424;
  assign n14426 = ~n14409 & ~n14410;
  assign n14427 = ~n10298 & ~n63176;
  assign n14428 = ~n10298 & n63176;
  assign n14429 = n10298 & n14281;
  assign n14430 = ~n14428 & ~n14429;
  assign n14431 = ~pi647 & n63176;
  assign n14432 = pi647 & n14281;
  assign n14433 = ~n14431 & ~n14432;
  assign n14434 = ~pi1157 & ~n14433;
  assign n14435 = pi647 & n63176;
  assign n14436 = ~pi647 & n14281;
  assign n14437 = ~n14435 & ~n14436;
  assign n14438 = pi1157 & ~n14437;
  assign n14439 = ~n14434 & ~n14438;
  assign n14440 = pi787 & ~n14439;
  assign n14441 = ~pi787 & n63176;
  assign n14442 = ~n14440 & ~n14441;
  assign n14443 = ~n14363 & ~n14427;
  assign n14444 = ~pi644 & ~n63177;
  assign n14445 = pi715 & ~n14444;
  assign n14446 = pi1160 & ~n14445;
  assign n14447 = pi1160 & ~n14362;
  assign n14448 = ~n14445 & n14447;
  assign n14449 = ~n14362 & n14446;
  assign n14450 = pi644 & ~n63177;
  assign n14451 = ~pi715 & ~n14450;
  assign n14452 = ~pi644 & n63172;
  assign n14453 = pi644 & n14281;
  assign n14454 = pi715 & ~n14453;
  assign n14455 = ~n14452 & n14454;
  assign n14456 = ~pi1160 & ~n14455;
  assign n14457 = ~n14451 & n14456;
  assign n14458 = ~n63178 & ~n14457;
  assign n14459 = pi790 & ~n14458;
  assign n14460 = ~n63052 & n14349;
  assign n14461 = n8332 & ~n14415;
  assign n14462 = n8332 & n14416;
  assign n14463 = ~n14414 & n14461;
  assign n14464 = n8331 & ~n14419;
  assign n14465 = n8331 & n14420;
  assign n14466 = ~n14418 & n14464;
  assign n14467 = ~n63179 & ~n63180;
  assign n14468 = ~n14460 & n14467;
  assign n14469 = pi792 & ~n14468;
  assign n14470 = pi704 & n14291;
  assign n14471 = ~pi176 & n10353;
  assign n14472 = ~n10355 & ~n10357;
  assign n14473 = pi176 & ~n14472;
  assign n14474 = pi742 & ~n14473;
  assign n14475 = ~n14471 & n14474;
  assign n14476 = pi176 & n10363;
  assign n14477 = ~pi176 & ~n62980;
  assign n14478 = ~pi742 & ~n14477;
  assign n14479 = ~n14476 & n14478;
  assign n14480 = ~pi704 & ~n14479;
  assign n14481 = ~pi176 & ~n10353;
  assign n14482 = pi176 & n14472;
  assign n14483 = pi742 & ~n14482;
  assign n14484 = ~n14481 & n14483;
  assign n14485 = pi176 & ~n10363;
  assign n14486 = ~pi176 & n62980;
  assign n14487 = ~pi742 & ~n14486;
  assign n14488 = ~n14485 & n14487;
  assign n14489 = ~n14484 & ~n14488;
  assign n14490 = ~pi704 & ~n14489;
  assign n14491 = ~n14475 & n14480;
  assign n14492 = n62765 & ~n63181;
  assign n14493 = n62765 & ~n14470;
  assign n14494 = ~n63181 & n14493;
  assign n14495 = ~n14470 & n14492;
  assign n14496 = ~n14283 & ~n63182;
  assign n14497 = ~pi625 & n14496;
  assign n14498 = pi625 & n14293;
  assign n14499 = ~pi1153 & ~n14498;
  assign n14500 = ~n14497 & n14499;
  assign n14501 = ~pi608 & ~n14381;
  assign n14502 = ~n14500 & n14501;
  assign n14503 = pi625 & n14496;
  assign n14504 = ~pi625 & n14293;
  assign n14505 = pi1153 & ~n14504;
  assign n14506 = ~n14503 & n14505;
  assign n14507 = pi608 & ~n14385;
  assign n14508 = ~n14506 & n14507;
  assign n14509 = ~n14502 & ~n14508;
  assign n14510 = pi778 & ~n14509;
  assign n14511 = ~pi778 & n14496;
  assign n14512 = ~n14510 & ~n14511;
  assign n14513 = ~pi609 & ~n14512;
  assign n14514 = pi609 & n14388;
  assign n14515 = ~pi1155 & ~n14514;
  assign n14516 = ~n14513 & n14515;
  assign n14517 = ~pi660 & ~n14301;
  assign n14518 = ~n14516 & n14517;
  assign n14519 = pi609 & ~n14512;
  assign n14520 = ~pi609 & n14388;
  assign n14521 = pi1155 & ~n14520;
  assign n14522 = ~n14519 & n14521;
  assign n14523 = pi660 & ~n14305;
  assign n14524 = ~n14522 & n14523;
  assign n14525 = ~n14518 & ~n14524;
  assign n14526 = pi785 & ~n14525;
  assign n14527 = ~pi785 & ~n14512;
  assign n14528 = ~n14526 & ~n14527;
  assign n14529 = pi618 & ~n14528;
  assign n14530 = ~pi618 & ~n63173;
  assign n14531 = pi1154 & ~n14530;
  assign n14532 = ~n14529 & n14531;
  assign n14533 = pi627 & ~n14317;
  assign n14534 = ~n14532 & n14533;
  assign n14535 = ~pi618 & ~n14528;
  assign n14536 = pi618 & ~n63173;
  assign n14537 = ~pi1154 & ~n14536;
  assign n14538 = ~n14535 & n14537;
  assign n14539 = ~pi627 & ~n14313;
  assign n14540 = ~n14538 & n14539;
  assign n14541 = pi781 & ~n14540;
  assign n14542 = ~n14534 & n14541;
  assign n14543 = ~n11431 & ~n63174;
  assign n14544 = ~n62884 & ~n63170;
  assign n14545 = ~n14543 & ~n14544;
  assign n14546 = pi789 & ~n14545;
  assign n14547 = ~pi781 & n14528;
  assign n14548 = ~n14546 & ~n14547;
  assign n14549 = ~n14542 & n14548;
  assign n14550 = n11434 & n14545;
  assign n14551 = ~n14549 & ~n14550;
  assign n14552 = ~n14534 & ~n14540;
  assign n14553 = pi781 & ~n14552;
  assign n14554 = ~pi781 & ~n14528;
  assign n14555 = ~n14553 & ~n14554;
  assign n14556 = ~pi619 & ~n14555;
  assign n14557 = pi619 & n63174;
  assign n14558 = ~pi1159 & ~n14557;
  assign n14559 = ~n14556 & n14558;
  assign n14560 = ~pi648 & ~n14332;
  assign n14561 = ~n14559 & n14560;
  assign n14562 = pi619 & ~n14555;
  assign n14563 = ~pi619 & n63174;
  assign n14564 = pi1159 & ~n14563;
  assign n14565 = ~n14562 & n14564;
  assign n14566 = pi648 & ~n14336;
  assign n14567 = ~n14565 & n14566;
  assign n14568 = pi789 & ~n14567;
  assign n14569 = pi789 & ~n14561;
  assign n14570 = ~n14567 & n14569;
  assign n14571 = ~n14561 & n14568;
  assign n14572 = ~pi789 & n14555;
  assign n14573 = n62894 & ~n14572;
  assign n14574 = ~n63183 & n14573;
  assign n14575 = n62894 & ~n14551;
  assign n14576 = ~pi626 & ~n63171;
  assign n14577 = pi626 & ~n14281;
  assign n14578 = n8301 & ~n14577;
  assign n14579 = ~n14576 & n14578;
  assign n14580 = n8525 & ~n63175;
  assign n14581 = pi626 & ~n63171;
  assign n14582 = ~pi626 & ~n14281;
  assign n14583 = n8300 & ~n14582;
  assign n14584 = ~n14581 & n14583;
  assign n14585 = ~n14580 & ~n14584;
  assign n14586 = ~n14579 & ~n14580;
  assign n14587 = ~n14584 & n14586;
  assign n14588 = ~n14579 & n14585;
  assign n14589 = pi788 & ~n63185;
  assign n14590 = ~n63184 & ~n14589;
  assign n14591 = ~n14469 & ~n14590;
  assign n14592 = n63030 & n14468;
  assign n14593 = ~n8651 & ~n14592;
  assign n14594 = ~n63030 & ~n14589;
  assign n14595 = ~n63184 & n14594;
  assign n14596 = ~n14469 & ~n14595;
  assign n14597 = ~n8651 & ~n14596;
  assign n14598 = ~n14591 & n14593;
  assign n14599 = ~n8413 & ~n14351;
  assign n14600 = ~n8413 & n14352;
  assign n14601 = ~n14350 & n14599;
  assign n14602 = n8374 & ~n14432;
  assign n14603 = n8374 & n14433;
  assign n14604 = ~n14431 & n14602;
  assign n14605 = n8373 & ~n14436;
  assign n14606 = n8373 & n14437;
  assign n14607 = ~n14435 & n14605;
  assign n14608 = ~n63188 & ~n63189;
  assign n14609 = ~n63187 & ~n63188;
  assign n14610 = ~n63189 & n14609;
  assign n14611 = ~n63187 & n14608;
  assign n14612 = pi787 & ~n63190;
  assign n14613 = ~pi644 & n14456;
  assign n14614 = pi644 & n14447;
  assign n14615 = n14029 & ~n14362;
  assign n14616 = pi790 & ~n63191;
  assign n14617 = pi790 & ~n14613;
  assign n14618 = ~n63191 & n14617;
  assign n14619 = ~n14613 & n14616;
  assign n14620 = ~n14612 & ~n63192;
  assign n14621 = ~n63186 & ~n14612;
  assign n14622 = ~n63192 & n14621;
  assign n14623 = ~n63186 & n14620;
  assign n14624 = ~n14459 & ~n63193;
  assign n14625 = n62455 & ~n14624;
  assign n14626 = ~pi176 & ~n62455;
  assign n14627 = ~pi832 & ~n14626;
  assign n14628 = ~n14625 & n14627;
  assign po333 = ~n14280 & ~n14628;
  assign n14630 = ~pi177 & ~n2923;
  assign n14631 = ~pi757 & n7316;
  assign n14632 = ~n14630 & ~n14631;
  assign n14633 = ~n8420 & ~n14632;
  assign n14634 = ~pi785 & ~n14633;
  assign n14635 = ~n8425 & ~n14632;
  assign n14636 = pi1155 & ~n14635;
  assign n14637 = ~n8428 & n14633;
  assign n14638 = ~pi1155 & ~n14637;
  assign n14639 = ~n14636 & ~n14638;
  assign n14640 = pi785 & ~n14639;
  assign n14641 = ~n14634 & ~n14640;
  assign n14642 = ~pi781 & ~n14641;
  assign n14643 = ~n8435 & n14641;
  assign n14644 = pi1154 & ~n14643;
  assign n14645 = ~n8438 & n14641;
  assign n14646 = ~pi1154 & ~n14645;
  assign n14647 = ~n14644 & ~n14646;
  assign n14648 = pi781 & ~n14647;
  assign n14649 = ~n14642 & ~n14648;
  assign n14650 = ~pi619 & ~n14649;
  assign n14651 = pi619 & ~n14630;
  assign n14652 = ~pi1159 & ~n14651;
  assign n14653 = ~n14650 & n14652;
  assign n14654 = pi619 & ~n14649;
  assign n14655 = ~pi619 & ~n14630;
  assign n14656 = pi1159 & ~n14655;
  assign n14657 = ~n14654 & n14656;
  assign n14658 = pi619 & n14649;
  assign n14659 = ~pi619 & n14630;
  assign n14660 = pi1159 & ~n14659;
  assign n14661 = ~n14658 & n14660;
  assign n14662 = ~pi619 & n14649;
  assign n14663 = pi619 & n14630;
  assign n14664 = ~pi1159 & ~n14663;
  assign n14665 = ~n14662 & n14664;
  assign n14666 = ~n14661 & ~n14665;
  assign n14667 = ~n14653 & ~n14657;
  assign n14668 = pi789 & n63194;
  assign n14669 = ~pi789 & n14649;
  assign n14670 = ~pi789 & ~n14649;
  assign n14671 = pi789 & ~n63194;
  assign n14672 = ~n14670 & ~n14671;
  assign n14673 = ~n14668 & ~n14669;
  assign n14674 = ~n8595 & n63195;
  assign n14675 = n8595 & n14630;
  assign n14676 = ~n8595 & ~n63195;
  assign n14677 = n8595 & ~n14630;
  assign n14678 = ~n14676 & ~n14677;
  assign n14679 = ~n14674 & ~n14675;
  assign n14680 = ~n8334 & n63196;
  assign n14681 = n8334 & n14630;
  assign n14682 = ~n8413 & ~n14681;
  assign n14683 = ~n14680 & ~n14681;
  assign n14684 = ~n8413 & n14683;
  assign n14685 = ~n14680 & n14682;
  assign n14686 = ~pi686 & n7564;
  assign n14687 = ~n14630 & ~n14686;
  assign n14688 = ~pi778 & n14687;
  assign n14689 = ~pi625 & n14686;
  assign n14690 = ~n14687 & ~n14689;
  assign n14691 = pi1153 & ~n14690;
  assign n14692 = ~pi1153 & ~n14630;
  assign n14693 = ~n14689 & n14692;
  assign n14694 = ~n14691 & ~n14693;
  assign n14695 = pi778 & ~n14694;
  assign n14696 = ~n14688 & ~n14695;
  assign n14697 = ~n8490 & n14696;
  assign n14698 = ~n8492 & n14697;
  assign n14699 = ~n8494 & n14698;
  assign n14700 = ~n8496 & n14699;
  assign n14701 = ~n8508 & n14700;
  assign n14702 = pi647 & ~n14701;
  assign n14703 = ~pi647 & ~n14630;
  assign n14704 = ~n14702 & ~n14703;
  assign n14705 = n8373 & ~n14704;
  assign n14706 = ~pi647 & n14701;
  assign n14707 = pi647 & n14630;
  assign n14708 = ~pi1157 & ~n14707;
  assign n14709 = ~n14706 & n14708;
  assign n14710 = pi630 & n14709;
  assign n14711 = ~n14705 & ~n14710;
  assign n14712 = ~n63197 & n14711;
  assign n14713 = pi787 & ~n14712;
  assign n14714 = ~pi626 & ~n63195;
  assign n14715 = pi626 & ~n14630;
  assign n14716 = n8301 & ~n14715;
  assign n14717 = ~n14714 & n14716;
  assign n14718 = n8525 & n14699;
  assign n14719 = pi626 & ~n63195;
  assign n14720 = ~pi626 & ~n14630;
  assign n14721 = n8300 & ~n14720;
  assign n14722 = ~n14719 & n14721;
  assign n14723 = ~n14718 & ~n14722;
  assign n14724 = ~n14717 & ~n14718;
  assign n14725 = ~n14722 & n14724;
  assign n14726 = ~n14717 & n14723;
  assign n14727 = pi788 & ~n63198;
  assign n14728 = ~n7187 & ~n14687;
  assign n14729 = pi625 & n14728;
  assign n14730 = n14632 & ~n14728;
  assign n14731 = ~n14729 & ~n14730;
  assign n14732 = n14692 & ~n14731;
  assign n14733 = ~pi608 & ~n14691;
  assign n14734 = ~n14732 & n14733;
  assign n14735 = pi1153 & n14632;
  assign n14736 = ~n14729 & n14735;
  assign n14737 = pi608 & ~n14693;
  assign n14738 = ~n14736 & n14737;
  assign n14739 = ~n14734 & ~n14738;
  assign n14740 = pi778 & ~n14739;
  assign n14741 = ~pi778 & ~n14730;
  assign n14742 = ~n14740 & ~n14741;
  assign n14743 = ~pi609 & ~n14742;
  assign n14744 = pi609 & n14696;
  assign n14745 = ~pi1155 & ~n14744;
  assign n14746 = ~n14743 & n14745;
  assign n14747 = ~pi660 & ~n14636;
  assign n14748 = ~n14746 & n14747;
  assign n14749 = pi609 & ~n14742;
  assign n14750 = ~pi609 & n14696;
  assign n14751 = pi1155 & ~n14750;
  assign n14752 = ~n14749 & n14751;
  assign n14753 = pi660 & ~n14638;
  assign n14754 = ~n14752 & n14753;
  assign n14755 = ~n14748 & ~n14754;
  assign n14756 = pi785 & ~n14755;
  assign n14757 = ~pi785 & ~n14742;
  assign n14758 = ~n14756 & ~n14757;
  assign n14759 = pi618 & ~n14758;
  assign n14760 = ~pi618 & n14697;
  assign n14761 = pi1154 & ~n14760;
  assign n14762 = ~n14759 & n14761;
  assign n14763 = pi627 & ~n14646;
  assign n14764 = ~n14762 & n14763;
  assign n14765 = ~pi618 & ~n14758;
  assign n14766 = pi618 & n14697;
  assign n14767 = ~pi1154 & ~n14766;
  assign n14768 = ~n14765 & n14767;
  assign n14769 = ~pi627 & ~n14644;
  assign n14770 = ~n14768 & n14769;
  assign n14771 = pi781 & ~n14770;
  assign n14772 = ~n14764 & n14771;
  assign n14773 = ~n11431 & ~n14698;
  assign n14774 = ~n62884 & ~n63194;
  assign n14775 = ~n14773 & ~n14774;
  assign n14776 = pi789 & ~n14775;
  assign n14777 = ~pi781 & n14758;
  assign n14778 = ~n14776 & ~n14777;
  assign n14779 = ~n14772 & n14778;
  assign n14780 = n11434 & n14775;
  assign n14781 = ~n14779 & ~n14780;
  assign n14782 = ~n14764 & ~n14770;
  assign n14783 = pi781 & ~n14782;
  assign n14784 = ~pi781 & ~n14758;
  assign n14785 = ~n14783 & ~n14784;
  assign n14786 = ~pi619 & ~n14785;
  assign n14787 = pi619 & n14698;
  assign n14788 = ~pi1159 & ~n14787;
  assign n14789 = ~n14786 & n14788;
  assign n14790 = ~pi648 & ~n14661;
  assign n14791 = ~n14789 & n14790;
  assign n14792 = pi619 & ~n14785;
  assign n14793 = ~pi619 & n14698;
  assign n14794 = pi1159 & ~n14793;
  assign n14795 = ~n14792 & n14794;
  assign n14796 = pi648 & ~n14665;
  assign n14797 = ~n14795 & n14796;
  assign n14798 = pi789 & ~n14797;
  assign n14799 = pi789 & ~n14791;
  assign n14800 = ~n14797 & n14799;
  assign n14801 = ~n14791 & n14798;
  assign n14802 = ~pi789 & n14785;
  assign n14803 = n62894 & ~n14802;
  assign n14804 = ~n63199 & n14803;
  assign n14805 = n62894 & ~n14781;
  assign n14806 = ~n14727 & ~n63200;
  assign n14807 = ~n63030 & ~n14806;
  assign n14808 = n8498 & n63196;
  assign n14809 = n8615 & n14700;
  assign n14810 = pi629 & ~n14809;
  assign n14811 = ~n14808 & n14810;
  assign n14812 = n8499 & n63196;
  assign n14813 = n8606 & n14700;
  assign n14814 = ~pi629 & ~n14813;
  assign n14815 = ~n14812 & n14814;
  assign n14816 = pi792 & ~n14815;
  assign n14817 = pi792 & ~n14811;
  assign n14818 = ~n14815 & n14817;
  assign n14819 = ~n14812 & ~n14813;
  assign n14820 = ~pi629 & ~n14819;
  assign n14821 = ~n14808 & ~n14809;
  assign n14822 = pi629 & ~n14821;
  assign n14823 = ~n14820 & ~n14822;
  assign n14824 = pi792 & ~n14823;
  assign n14825 = ~n14811 & n14816;
  assign n14826 = ~n8651 & ~n63201;
  assign n14827 = ~n14807 & n14826;
  assign n14828 = ~n14713 & ~n14827;
  assign n14829 = pi644 & n14828;
  assign n14830 = ~pi787 & ~n14701;
  assign n14831 = pi1157 & ~n14704;
  assign n14832 = ~n14709 & ~n14831;
  assign n14833 = pi787 & ~n14832;
  assign n14834 = ~n14830 & ~n14833;
  assign n14835 = ~pi644 & n14834;
  assign n14836 = pi715 & ~n14835;
  assign n14837 = ~n14829 & n14836;
  assign n14838 = ~n8685 & n14630;
  assign n14839 = ~n8376 & n14680;
  assign n14840 = ~n8376 & ~n14683;
  assign n14841 = n8376 & n14630;
  assign n14842 = ~n14840 & ~n14841;
  assign n14843 = ~n14838 & ~n14839;
  assign n14844 = pi644 & ~n63202;
  assign n14845 = ~pi644 & n14630;
  assign n14846 = ~pi715 & ~n14845;
  assign n14847 = ~n14844 & n14846;
  assign n14848 = pi1160 & ~n14847;
  assign n14849 = ~n14837 & n14848;
  assign n14850 = ~pi644 & n14828;
  assign n14851 = pi644 & n14834;
  assign n14852 = ~pi715 & ~n14851;
  assign n14853 = ~n14850 & n14852;
  assign n14854 = ~pi644 & ~n63202;
  assign n14855 = pi644 & n14630;
  assign n14856 = pi715 & ~n14855;
  assign n14857 = ~n14854 & n14856;
  assign n14858 = ~pi1160 & ~n14857;
  assign n14859 = ~n14853 & n14858;
  assign n14860 = ~n14849 & ~n14859;
  assign n14861 = pi790 & ~n14860;
  assign n14862 = ~pi790 & n14828;
  assign n14863 = pi832 & ~n14862;
  assign n14864 = ~n14861 & n14863;
  assign n14865 = ~pi177 & ~n8098;
  assign n14866 = n8257 & ~n14865;
  assign n14867 = pi177 & ~n62765;
  assign n14868 = ~pi177 & n8009;
  assign n14869 = pi177 & n62874;
  assign n14870 = ~pi38 & ~n14869;
  assign n14871 = ~n14868 & n14870;
  assign n14872 = ~pi177 & ~n7357;
  assign n14873 = n8085 & ~n14872;
  assign n14874 = ~pi686 & ~n14873;
  assign n14875 = ~n14871 & n14874;
  assign n14876 = ~pi177 & pi686;
  assign n14877 = ~n8091 & n14876;
  assign n14878 = n62765 & ~n14877;
  assign n14879 = ~n14875 & n14878;
  assign n14880 = ~n14867 & ~n14879;
  assign n14881 = ~pi778 & ~n14880;
  assign n14882 = pi625 & n14880;
  assign n14883 = ~pi625 & n14865;
  assign n14884 = pi1153 & ~n14883;
  assign n14885 = ~n14882 & n14884;
  assign n14886 = ~pi625 & n14880;
  assign n14887 = pi625 & n14865;
  assign n14888 = ~pi1153 & ~n14887;
  assign n14889 = ~n14886 & n14888;
  assign n14890 = ~n14885 & ~n14889;
  assign n14891 = pi778 & ~n14890;
  assign n14892 = ~n14881 & ~n14891;
  assign n14893 = ~n62880 & ~n14892;
  assign n14894 = n62880 & ~n14865;
  assign n14895 = ~n62880 & n14892;
  assign n14896 = n62880 & n14865;
  assign n14897 = ~n14895 & ~n14896;
  assign n14898 = ~n14893 & ~n14894;
  assign n14899 = ~n62882 & ~n63203;
  assign n14900 = n62882 & n14865;
  assign n14901 = n62882 & ~n14865;
  assign n14902 = ~n62882 & n63203;
  assign n14903 = ~n14901 & ~n14902;
  assign n14904 = ~n14899 & ~n14900;
  assign n14905 = ~n8257 & ~n63204;
  assign n14906 = ~n14866 & ~n14905;
  assign n14907 = ~n8303 & n14906;
  assign n14908 = n8303 & n14865;
  assign n14909 = n8303 & ~n14865;
  assign n14910 = ~n8257 & n63204;
  assign n14911 = n8257 & n14865;
  assign n14912 = ~n14910 & ~n14911;
  assign n14913 = ~n8303 & n14912;
  assign n14914 = ~n14909 & ~n14913;
  assign n14915 = ~n14907 & ~n14908;
  assign n14916 = ~pi792 & ~n63205;
  assign n14917 = pi628 & n63205;
  assign n14918 = ~pi628 & n14865;
  assign n14919 = pi1156 & ~n14918;
  assign n14920 = ~pi628 & ~n14865;
  assign n14921 = pi628 & ~n63205;
  assign n14922 = ~n14920 & ~n14921;
  assign n14923 = pi1156 & ~n14922;
  assign n14924 = ~n14917 & n14919;
  assign n14925 = ~pi628 & n63205;
  assign n14926 = pi628 & n14865;
  assign n14927 = ~pi1156 & ~n14926;
  assign n14928 = ~n14925 & n14927;
  assign n14929 = ~n63206 & ~n14928;
  assign n14930 = pi792 & ~n14929;
  assign n14931 = ~n14916 & ~n14930;
  assign n14932 = ~pi787 & ~n14931;
  assign n14933 = ~pi647 & n14931;
  assign n14934 = pi647 & n14865;
  assign n14935 = ~pi1157 & ~n14934;
  assign n14936 = ~n14933 & n14935;
  assign n14937 = pi647 & n14931;
  assign n14938 = ~pi647 & n14865;
  assign n14939 = pi1157 & ~n14938;
  assign n14940 = ~pi647 & ~n14865;
  assign n14941 = pi647 & ~n14931;
  assign n14942 = ~n14940 & ~n14941;
  assign n14943 = ~n14937 & ~n14938;
  assign n14944 = pi1157 & ~n63207;
  assign n14945 = ~n14937 & n14939;
  assign n14946 = ~n14936 & ~n63208;
  assign n14947 = pi787 & ~n14946;
  assign n14948 = ~n14932 & ~n14947;
  assign n14949 = ~pi644 & pi715;
  assign n14950 = ~n14948 & n14949;
  assign n14951 = pi757 & n8091;
  assign n14952 = ~pi177 & ~pi757;
  assign n14953 = n10343 & n14952;
  assign n14954 = ~pi757 & ~n14285;
  assign n14955 = pi177 & ~n14954;
  assign n14956 = ~n14953 & ~n14955;
  assign n14957 = pi757 & ~n8091;
  assign n14958 = ~pi757 & ~n10343;
  assign n14959 = ~n14957 & ~n14958;
  assign n14960 = ~pi177 & ~n14959;
  assign n14961 = ~pi177 & ~n62977;
  assign n14962 = ~pi757 & ~n14961;
  assign n14963 = ~n14285 & n14962;
  assign n14964 = ~n14960 & ~n14963;
  assign n14965 = ~n14951 & n14956;
  assign n14966 = n62765 & n63209;
  assign n14967 = ~n14867 & ~n14966;
  assign n14968 = ~n8135 & ~n14967;
  assign n14969 = n8135 & ~n14865;
  assign n14970 = ~n14968 & ~n14969;
  assign n14971 = ~pi785 & ~n14970;
  assign n14972 = ~n8136 & ~n14865;
  assign n14973 = pi609 & n14968;
  assign n14974 = ~n14972 & ~n14973;
  assign n14975 = pi1155 & ~n14974;
  assign n14976 = ~n8148 & ~n14865;
  assign n14977 = ~pi609 & n14968;
  assign n14978 = ~n14976 & ~n14977;
  assign n14979 = ~pi1155 & ~n14978;
  assign n14980 = ~n14975 & ~n14979;
  assign n14981 = pi785 & ~n14980;
  assign n14982 = ~n14971 & ~n14981;
  assign n14983 = ~pi781 & ~n14982;
  assign n14984 = pi618 & n14982;
  assign n14985 = ~pi618 & n14865;
  assign n14986 = pi1154 & ~n14985;
  assign n14987 = ~n14984 & n14986;
  assign n14988 = ~pi618 & n14982;
  assign n14989 = pi618 & n14865;
  assign n14990 = ~pi1154 & ~n14989;
  assign n14991 = ~n14988 & n14990;
  assign n14992 = ~n14987 & ~n14991;
  assign n14993 = pi781 & ~n14992;
  assign n14994 = ~n14983 & ~n14993;
  assign n14995 = ~pi789 & ~n14994;
  assign n14996 = ~pi619 & n14994;
  assign n14997 = pi619 & n14865;
  assign n14998 = ~pi1159 & ~n14997;
  assign n14999 = ~n14996 & n14998;
  assign n15000 = pi619 & n14994;
  assign n15001 = ~pi619 & n14865;
  assign n15002 = pi1159 & ~n15001;
  assign n15003 = ~n15000 & n15002;
  assign n15004 = ~n14999 & ~n15003;
  assign n15005 = pi789 & ~n15004;
  assign n15006 = ~n14995 & ~n15005;
  assign n15007 = ~n8595 & n15006;
  assign n15008 = n8595 & n14865;
  assign n15009 = ~n15007 & ~n15008;
  assign n15010 = ~n8334 & ~n15009;
  assign n15011 = n8334 & n14865;
  assign n15012 = ~n15010 & ~n15011;
  assign n15013 = ~n8376 & ~n15012;
  assign n15014 = n8376 & n14865;
  assign n15015 = n8376 & ~n14865;
  assign n15016 = ~n8376 & n15012;
  assign n15017 = ~n15015 & ~n15016;
  assign n15018 = ~n15013 & ~n15014;
  assign n15019 = pi644 & n63210;
  assign n15020 = ~pi644 & n14865;
  assign n15021 = ~pi715 & ~n15020;
  assign n15022 = ~n15019 & n15021;
  assign n15023 = pi1160 & ~n15022;
  assign n15024 = ~n14950 & n15023;
  assign n15025 = pi644 & ~pi715;
  assign n15026 = ~n14948 & n15025;
  assign n15027 = ~pi644 & n63210;
  assign n15028 = pi644 & n14865;
  assign n15029 = pi715 & ~n15028;
  assign n15030 = ~n15027 & n15029;
  assign n15031 = ~pi1160 & ~n15030;
  assign n15032 = ~n15026 & n15031;
  assign n15033 = pi790 & ~n15032;
  assign n15034 = ~n15024 & n15033;
  assign n15035 = ~n63052 & n15009;
  assign n15036 = n8331 & ~n14922;
  assign n15037 = ~pi629 & n63206;
  assign n15038 = pi629 & n14928;
  assign n15039 = ~n63211 & ~n15038;
  assign n15040 = ~n15035 & n15039;
  assign n15041 = pi792 & ~n15040;
  assign n15042 = pi619 & n63204;
  assign n15043 = ~pi1159 & ~n15042;
  assign n15044 = ~pi648 & ~n15043;
  assign n15045 = ~pi648 & ~n15003;
  assign n15046 = ~n15043 & n15045;
  assign n15047 = ~n15003 & n15044;
  assign n15048 = ~pi619 & n63204;
  assign n15049 = pi1159 & ~n15048;
  assign n15050 = pi648 & ~n14999;
  assign n15051 = ~n15049 & n15050;
  assign n15052 = ~n63212 & ~n15051;
  assign n15053 = pi789 & ~n15052;
  assign n15054 = ~pi177 & n8759;
  assign n15055 = pi177 & n8763;
  assign n15056 = ~pi38 & ~n15055;
  assign n15057 = ~n15054 & n15056;
  assign n15058 = n8793 & ~n14872;
  assign n15059 = pi757 & ~n15058;
  assign n15060 = ~n15057 & n15059;
  assign n15061 = pi177 & n8775;
  assign n15062 = ~pi177 & ~n8779;
  assign n15063 = ~pi38 & ~n15062;
  assign n15064 = ~n15061 & n15063;
  assign n15065 = ~pi177 & ~n10366;
  assign n15066 = pi177 & n62856;
  assign n15067 = pi38 & ~n15066;
  assign n15068 = ~n15065 & n15067;
  assign n15069 = n10362 & ~n14872;
  assign n15070 = ~pi757 & ~n63213;
  assign n15071 = ~n15064 & n15070;
  assign n15072 = ~n15060 & ~n15071;
  assign n15073 = ~pi686 & ~n15072;
  assign n15074 = pi686 & ~n63209;
  assign n15075 = n62765 & ~n15074;
  assign n15076 = n62765 & ~n15073;
  assign n15077 = ~n15074 & n15076;
  assign n15078 = ~n15073 & n15075;
  assign n15079 = ~n14867 & ~n63214;
  assign n15080 = ~pi625 & n15079;
  assign n15081 = pi625 & n14967;
  assign n15082 = ~pi1153 & ~n15081;
  assign n15083 = ~n15080 & n15082;
  assign n15084 = ~pi608 & ~n14885;
  assign n15085 = ~n15083 & n15084;
  assign n15086 = pi625 & n15079;
  assign n15087 = ~pi625 & n14967;
  assign n15088 = pi1153 & ~n15087;
  assign n15089 = ~n15086 & n15088;
  assign n15090 = pi608 & ~n14889;
  assign n15091 = ~n15089 & n15090;
  assign n15092 = ~n15085 & ~n15091;
  assign n15093 = pi778 & ~n15092;
  assign n15094 = ~pi778 & n15079;
  assign n15095 = ~pi778 & ~n15079;
  assign n15096 = pi778 & ~n15091;
  assign n15097 = ~n15085 & n15096;
  assign n15098 = ~n15095 & ~n15097;
  assign n15099 = ~n15093 & ~n15094;
  assign n15100 = ~pi609 & n63215;
  assign n15101 = pi609 & n14892;
  assign n15102 = ~pi1155 & ~n15101;
  assign n15103 = ~n15100 & n15102;
  assign n15104 = ~pi660 & ~n14975;
  assign n15105 = ~n15103 & n15104;
  assign n15106 = pi609 & n63215;
  assign n15107 = ~pi609 & n14892;
  assign n15108 = pi1155 & ~n15107;
  assign n15109 = ~n15106 & n15108;
  assign n15110 = pi660 & ~n14979;
  assign n15111 = ~n15109 & n15110;
  assign n15112 = ~n15105 & ~n15111;
  assign n15113 = pi785 & ~n15112;
  assign n15114 = ~pi785 & n63215;
  assign n15115 = ~n15113 & ~n15114;
  assign n15116 = ~pi618 & ~n15115;
  assign n15117 = pi618 & ~n63203;
  assign n15118 = ~pi1154 & ~n15117;
  assign n15119 = ~n15116 & n15118;
  assign n15120 = ~pi627 & ~n14987;
  assign n15121 = ~n15119 & n15120;
  assign n15122 = pi618 & ~n15115;
  assign n15123 = ~pi618 & ~n63203;
  assign n15124 = pi1154 & ~n15123;
  assign n15125 = ~n15122 & n15124;
  assign n15126 = pi627 & ~n14991;
  assign n15127 = ~n15125 & n15126;
  assign n15128 = pi781 & ~n15127;
  assign n15129 = pi781 & ~n15121;
  assign n15130 = ~n15127 & n15129;
  assign n15131 = ~n15121 & n15128;
  assign n15132 = ~pi781 & n15115;
  assign n15133 = pi619 & n15050;
  assign n15134 = ~pi619 & n15045;
  assign n15135 = n11420 & ~n15003;
  assign n15136 = pi789 & ~n63217;
  assign n15137 = pi789 & ~n15133;
  assign n15138 = ~n63217 & n15137;
  assign n15139 = ~n15133 & n15136;
  assign n15140 = ~n15132 & ~n63218;
  assign n15141 = ~n63216 & n15140;
  assign n15142 = ~n15121 & ~n15127;
  assign n15143 = pi781 & ~n15142;
  assign n15144 = ~pi781 & ~n15115;
  assign n15145 = ~n15143 & ~n15144;
  assign n15146 = ~pi619 & ~n15145;
  assign n15147 = n15043 & ~n15146;
  assign n15148 = n15045 & ~n15147;
  assign n15149 = pi619 & ~n15145;
  assign n15150 = n15049 & ~n15149;
  assign n15151 = n15050 & ~n15150;
  assign n15152 = ~n15148 & ~n15151;
  assign n15153 = pi789 & ~n15152;
  assign n15154 = ~pi789 & ~n15145;
  assign n15155 = ~n15153 & ~n15154;
  assign n15156 = ~n15053 & ~n15141;
  assign n15157 = n62894 & ~n63219;
  assign n15158 = n12979 & n15006;
  assign n15159 = ~pi641 & n14912;
  assign n15160 = ~pi641 & ~n14906;
  assign n15161 = pi641 & ~n14865;
  assign n15162 = n8417 & ~n15161;
  assign n15163 = ~n63220 & n15162;
  assign n15164 = pi641 & n14912;
  assign n15165 = pi641 & ~n14906;
  assign n15166 = ~pi641 & ~n14865;
  assign n15167 = n8416 & ~n15166;
  assign n15168 = ~n63221 & n15167;
  assign n15169 = ~n15163 & ~n15168;
  assign n15170 = ~n15158 & n15169;
  assign n15171 = pi788 & ~n15170;
  assign n15172 = ~n63030 & ~n15171;
  assign n15173 = ~n15157 & n15172;
  assign n15174 = ~pi788 & n63219;
  assign n15175 = ~pi626 & n63219;
  assign n15176 = pi626 & ~n14906;
  assign n15177 = ~pi641 & ~n15176;
  assign n15178 = ~n15175 & n15177;
  assign n15179 = ~pi626 & ~n15006;
  assign n15180 = pi626 & ~n14865;
  assign n15181 = pi641 & ~n15180;
  assign n15182 = ~n15179 & n15181;
  assign n15183 = ~pi1158 & ~n15182;
  assign n15184 = ~n15178 & n15183;
  assign n15185 = pi626 & n63219;
  assign n15186 = ~pi626 & ~n14906;
  assign n15187 = pi641 & ~n15186;
  assign n15188 = ~n15185 & n15187;
  assign n15189 = pi626 & ~n15006;
  assign n15190 = ~pi626 & ~n14865;
  assign n15191 = ~pi641 & ~n15190;
  assign n15192 = ~n15189 & n15191;
  assign n15193 = pi1158 & ~n15192;
  assign n15194 = ~n15188 & n15193;
  assign n15195 = ~n15184 & ~n15194;
  assign n15196 = pi788 & ~n15195;
  assign n15197 = ~n15174 & ~n15196;
  assign n15198 = ~pi628 & n15197;
  assign n15199 = pi628 & ~n15009;
  assign n15200 = ~pi1156 & ~n15199;
  assign n15201 = ~n15198 & n15200;
  assign n15202 = ~pi629 & ~n63206;
  assign n15203 = ~n15201 & n15202;
  assign n15204 = pi628 & n15197;
  assign n15205 = ~pi628 & ~n15009;
  assign n15206 = pi1156 & ~n15205;
  assign n15207 = ~n15204 & n15206;
  assign n15208 = pi629 & ~n14928;
  assign n15209 = ~n15207 & n15208;
  assign n15210 = ~n15203 & ~n15209;
  assign n15211 = pi792 & ~n15210;
  assign n15212 = ~pi792 & n15197;
  assign n15213 = ~n15211 & ~n15212;
  assign n15214 = ~n15041 & ~n15173;
  assign n15215 = ~n8651 & n63222;
  assign n15216 = ~n8413 & n15012;
  assign n15217 = n8373 & ~n63207;
  assign n15218 = pi630 & n14936;
  assign n15219 = ~n15217 & ~n15218;
  assign n15220 = ~n15216 & n15219;
  assign n15221 = pi787 & ~n15220;
  assign n15222 = ~n62896 & n63222;
  assign n15223 = ~pi647 & ~n63222;
  assign n15224 = pi647 & ~n15012;
  assign n15225 = ~pi1157 & ~n15224;
  assign n15226 = ~n15223 & n15225;
  assign n15227 = ~pi630 & ~n63208;
  assign n15228 = ~n15226 & n15227;
  assign n15229 = pi647 & ~n63222;
  assign n15230 = ~pi647 & ~n15012;
  assign n15231 = pi1157 & ~n15230;
  assign n15232 = ~n15229 & n15231;
  assign n15233 = pi630 & ~n14936;
  assign n15234 = ~n15232 & n15233;
  assign n15235 = ~n15228 & ~n15234;
  assign n15236 = n15220 & ~n15222;
  assign n15237 = pi787 & n63223;
  assign n15238 = ~pi787 & n63222;
  assign n15239 = ~n15237 & ~n15238;
  assign n15240 = pi787 & ~n63223;
  assign n15241 = ~pi787 & ~n63222;
  assign n15242 = ~n15240 & ~n15241;
  assign n15243 = ~n15215 & ~n15221;
  assign n15244 = ~n11547 & ~n63224;
  assign n15245 = n62455 & ~n15244;
  assign n15246 = ~pi644 & n63224;
  assign n15247 = pi644 & n14948;
  assign n15248 = ~pi715 & ~n15247;
  assign n15249 = ~n15246 & n15248;
  assign n15250 = n15031 & ~n15249;
  assign n15251 = ~pi644 & n14948;
  assign n15252 = pi715 & ~n15251;
  assign n15253 = n15023 & ~n15252;
  assign n15254 = ~n15250 & ~n15253;
  assign n15255 = pi790 & ~n15254;
  assign n15256 = pi644 & n15023;
  assign n15257 = pi790 & ~n15256;
  assign n15258 = n63224 & ~n15257;
  assign n15259 = ~n15255 & ~n15258;
  assign n15260 = n62455 & ~n15259;
  assign n15261 = pi644 & n63224;
  assign n15262 = n15252 & ~n15261;
  assign n15263 = n15023 & ~n15262;
  assign n15264 = pi790 & ~n15250;
  assign n15265 = pi790 & ~n15263;
  assign n15266 = ~n15250 & n15265;
  assign n15267 = ~n15263 & n15264;
  assign n15268 = ~pi790 & ~n63224;
  assign n15269 = n62455 & ~n15268;
  assign n15270 = ~n63226 & n15269;
  assign n15271 = ~n15034 & n15245;
  assign n15272 = ~pi177 & ~n62455;
  assign n15273 = ~pi832 & ~n15272;
  assign n15274 = ~n63225 & n15273;
  assign po334 = ~n14864 & ~n15274;
  assign n15276 = ~pi178 & ~n2923;
  assign n15277 = ~pi760 & n7316;
  assign n15278 = ~n15276 & ~n15277;
  assign n15279 = ~n8420 & ~n15278;
  assign n15280 = ~pi785 & ~n15279;
  assign n15281 = n8148 & n15277;
  assign n15282 = n15279 & ~n15281;
  assign n15283 = pi1155 & ~n15282;
  assign n15284 = ~pi1155 & ~n15276;
  assign n15285 = ~n15281 & n15284;
  assign n15286 = ~n15283 & ~n15285;
  assign n15287 = pi785 & ~n15286;
  assign n15288 = ~n15280 & ~n15287;
  assign n15289 = ~pi781 & ~n15288;
  assign n15290 = ~n8435 & n15288;
  assign n15291 = pi1154 & ~n15290;
  assign n15292 = ~n8438 & n15288;
  assign n15293 = ~pi1154 & ~n15292;
  assign n15294 = ~n15291 & ~n15293;
  assign n15295 = pi781 & ~n15294;
  assign n15296 = ~n15289 & ~n15295;
  assign n15297 = pi789 & ~n13462;
  assign n15298 = ~n13460 & n15297;
  assign n15299 = ~pi789 & ~n15296;
  assign n15300 = ~n12612 & n15296;
  assign n15301 = pi1159 & ~n15300;
  assign n15302 = ~n12615 & n15296;
  assign n15303 = ~pi1159 & ~n15302;
  assign n15304 = ~n15301 & ~n15303;
  assign n15305 = pi789 & ~n15304;
  assign n15306 = ~n15299 & ~n15305;
  assign n15307 = n15296 & ~n15298;
  assign n15308 = ~n8595 & n63227;
  assign n15309 = n8595 & n15276;
  assign n15310 = ~n8595 & ~n63227;
  assign n15311 = n8595 & ~n15276;
  assign n15312 = ~n15310 & ~n15311;
  assign n15313 = ~n15308 & ~n15309;
  assign n15314 = ~n8334 & n63228;
  assign n15315 = n8334 & n15276;
  assign n15316 = ~n8413 & ~n15315;
  assign n15317 = ~n15314 & ~n15315;
  assign n15318 = ~n8413 & n15317;
  assign n15319 = ~n15314 & n15316;
  assign n15320 = ~pi688 & n7564;
  assign n15321 = ~n15276 & ~n15320;
  assign n15322 = ~pi778 & ~n15321;
  assign n15323 = ~pi625 & n15320;
  assign n15324 = ~n15321 & ~n15323;
  assign n15325 = pi1153 & ~n15324;
  assign n15326 = ~pi1153 & ~n15276;
  assign n15327 = ~n15323 & n15326;
  assign n15328 = pi778 & ~n15327;
  assign n15329 = ~n15325 & n15328;
  assign n15330 = ~n15322 & ~n15329;
  assign n15331 = ~n8490 & ~n15330;
  assign n15332 = ~n8492 & n15331;
  assign n15333 = ~n8494 & n15332;
  assign n15334 = ~n8496 & n15333;
  assign n15335 = ~n8508 & n15334;
  assign n15336 = pi647 & ~n15335;
  assign n15337 = ~pi647 & ~n15276;
  assign n15338 = ~n15336 & ~n15337;
  assign n15339 = n8373 & ~n15338;
  assign n15340 = ~pi647 & n15335;
  assign n15341 = pi647 & n15276;
  assign n15342 = ~pi1157 & ~n15341;
  assign n15343 = ~n15340 & n15342;
  assign n15344 = pi630 & n15343;
  assign n15345 = ~n15339 & ~n15344;
  assign n15346 = ~n63229 & n15345;
  assign n15347 = pi787 & ~n15346;
  assign n15348 = ~pi626 & ~n63227;
  assign n15349 = pi626 & ~n15276;
  assign n15350 = n8301 & ~n15349;
  assign n15351 = ~n15348 & n15350;
  assign n15352 = n8525 & n15333;
  assign n15353 = pi626 & ~n63227;
  assign n15354 = ~pi626 & ~n15276;
  assign n15355 = n8300 & ~n15354;
  assign n15356 = ~n15353 & n15355;
  assign n15357 = ~n15352 & ~n15356;
  assign n15358 = ~n15351 & ~n15352;
  assign n15359 = ~n15356 & n15358;
  assign n15360 = ~n15351 & n15357;
  assign n15361 = pi788 & ~n63230;
  assign n15362 = n13460 & n15296;
  assign n15363 = n11303 & n15332;
  assign n15364 = pi648 & ~n15363;
  assign n15365 = ~n15362 & n15364;
  assign n15366 = n13462 & n15296;
  assign n15367 = n11304 & n15332;
  assign n15368 = ~pi648 & ~n15367;
  assign n15369 = ~n15366 & n15368;
  assign n15370 = pi789 & ~n15369;
  assign n15371 = ~n15365 & n15370;
  assign n15372 = ~n7187 & ~n15321;
  assign n15373 = pi625 & n15372;
  assign n15374 = n15278 & ~n15372;
  assign n15375 = ~n15373 & ~n15374;
  assign n15376 = n15326 & ~n15375;
  assign n15377 = ~pi608 & ~n15325;
  assign n15378 = ~n15376 & n15377;
  assign n15379 = pi1153 & n15278;
  assign n15380 = ~n15373 & n15379;
  assign n15381 = pi608 & ~n15327;
  assign n15382 = ~n15380 & n15381;
  assign n15383 = ~n15378 & ~n15382;
  assign n15384 = pi778 & ~n15383;
  assign n15385 = ~pi778 & ~n15374;
  assign n15386 = ~n15384 & ~n15385;
  assign n15387 = ~pi609 & ~n15386;
  assign n15388 = pi609 & ~n15330;
  assign n15389 = ~pi1155 & ~n15388;
  assign n15390 = ~n15387 & n15389;
  assign n15391 = ~pi660 & ~n15283;
  assign n15392 = ~n15390 & n15391;
  assign n15393 = pi609 & ~n15386;
  assign n15394 = ~pi609 & ~n15330;
  assign n15395 = pi1155 & ~n15394;
  assign n15396 = ~n15393 & n15395;
  assign n15397 = pi660 & ~n15285;
  assign n15398 = ~n15396 & n15397;
  assign n15399 = ~n15392 & ~n15398;
  assign n15400 = pi785 & ~n15399;
  assign n15401 = ~pi785 & ~n15386;
  assign n15402 = ~n15400 & ~n15401;
  assign n15403 = pi618 & ~n15402;
  assign n15404 = ~pi618 & n15331;
  assign n15405 = pi1154 & ~n15404;
  assign n15406 = ~n15403 & n15405;
  assign n15407 = pi627 & ~n15293;
  assign n15408 = ~n15406 & n15407;
  assign n15409 = ~pi618 & ~n15402;
  assign n15410 = pi618 & n15331;
  assign n15411 = ~pi1154 & ~n15410;
  assign n15412 = ~n15409 & n15411;
  assign n15413 = ~pi627 & ~n15291;
  assign n15414 = ~n15412 & n15413;
  assign n15415 = pi781 & ~n15414;
  assign n15416 = ~n15408 & n15415;
  assign n15417 = ~pi781 & n15402;
  assign n15418 = ~n11434 & ~n15417;
  assign n15419 = ~n15416 & n15418;
  assign n15420 = ~n15371 & ~n15419;
  assign n15421 = ~n15408 & ~n15414;
  assign n15422 = pi781 & ~n15421;
  assign n15423 = ~pi781 & ~n15402;
  assign n15424 = ~n15422 & ~n15423;
  assign n15425 = ~pi619 & ~n15424;
  assign n15426 = pi619 & n15332;
  assign n15427 = ~pi1159 & ~n15426;
  assign n15428 = ~n15425 & n15427;
  assign n15429 = ~pi648 & ~n15301;
  assign n15430 = ~n15428 & n15429;
  assign n15431 = pi619 & ~n15424;
  assign n15432 = ~pi619 & n15332;
  assign n15433 = pi1159 & ~n15432;
  assign n15434 = ~n15431 & n15433;
  assign n15435 = pi648 & ~n15303;
  assign n15436 = ~n15434 & n15435;
  assign n15437 = pi789 & ~n15436;
  assign n15438 = pi789 & ~n15430;
  assign n15439 = ~n15436 & n15438;
  assign n15440 = ~n15430 & n15437;
  assign n15441 = ~pi789 & n15424;
  assign n15442 = n62894 & ~n15441;
  assign n15443 = ~n63231 & n15442;
  assign n15444 = n62894 & ~n15420;
  assign n15445 = ~n15361 & ~n63232;
  assign n15446 = ~n63030 & ~n15445;
  assign n15447 = n8498 & n63228;
  assign n15448 = n8615 & n15334;
  assign n15449 = pi629 & ~n15448;
  assign n15450 = ~n15447 & n15449;
  assign n15451 = n8499 & n63228;
  assign n15452 = n8606 & n15334;
  assign n15453 = ~pi629 & ~n15452;
  assign n15454 = ~n15451 & n15453;
  assign n15455 = pi792 & ~n15454;
  assign n15456 = pi792 & ~n15450;
  assign n15457 = ~n15454 & n15456;
  assign n15458 = ~n15451 & ~n15452;
  assign n15459 = ~pi629 & ~n15458;
  assign n15460 = ~n15447 & ~n15448;
  assign n15461 = pi629 & ~n15460;
  assign n15462 = ~n15459 & ~n15461;
  assign n15463 = pi792 & ~n15462;
  assign n15464 = ~n15450 & n15455;
  assign n15465 = ~n8651 & ~n63233;
  assign n15466 = ~n15446 & n15465;
  assign n15467 = ~n15347 & ~n15466;
  assign n15468 = pi644 & n15467;
  assign n15469 = ~pi787 & ~n15335;
  assign n15470 = pi1157 & ~n15338;
  assign n15471 = ~n15343 & ~n15470;
  assign n15472 = pi787 & ~n15471;
  assign n15473 = ~n15469 & ~n15472;
  assign n15474 = ~pi644 & n15473;
  assign n15475 = pi715 & ~n15474;
  assign n15476 = ~n15468 & n15475;
  assign n15477 = ~n8685 & n15276;
  assign n15478 = ~n8376 & n15314;
  assign n15479 = ~n8376 & ~n15317;
  assign n15480 = n8376 & n15276;
  assign n15481 = ~n15479 & ~n15480;
  assign n15482 = ~n15477 & ~n15478;
  assign n15483 = pi644 & ~n63234;
  assign n15484 = ~pi644 & n15276;
  assign n15485 = ~pi715 & ~n15484;
  assign n15486 = ~n15483 & n15485;
  assign n15487 = pi1160 & ~n15486;
  assign n15488 = ~n15476 & n15487;
  assign n15489 = ~pi644 & n15467;
  assign n15490 = pi644 & n15473;
  assign n15491 = ~pi715 & ~n15490;
  assign n15492 = ~n15489 & n15491;
  assign n15493 = ~pi644 & ~n63234;
  assign n15494 = pi644 & n15276;
  assign n15495 = pi715 & ~n15494;
  assign n15496 = ~n15493 & n15495;
  assign n15497 = ~pi1160 & ~n15496;
  assign n15498 = ~n15492 & n15497;
  assign n15499 = ~n15488 & ~n15498;
  assign n15500 = pi790 & ~n15499;
  assign n15501 = ~pi790 & n15467;
  assign n15502 = pi832 & ~n15501;
  assign n15503 = ~n15500 & n15502;
  assign n15504 = ~pi178 & ~n8098;
  assign n15505 = n8257 & ~n15504;
  assign n15506 = ~pi688 & n62765;
  assign n15507 = n15504 & ~n15506;
  assign n15508 = pi178 & n62874;
  assign n15509 = ~pi38 & ~n15508;
  assign n15510 = n62765 & ~n15509;
  assign n15511 = ~pi178 & n8009;
  assign n15512 = ~n15510 & ~n15511;
  assign n15513 = ~pi178 & ~n7357;
  assign n15514 = n8085 & ~n15513;
  assign n15515 = ~pi688 & ~n15514;
  assign n15516 = ~n15512 & n15515;
  assign n15517 = ~n15507 & ~n15516;
  assign n15518 = ~pi778 & n15517;
  assign n15519 = pi625 & ~n15517;
  assign n15520 = ~pi625 & n15504;
  assign n15521 = pi1153 & ~n15520;
  assign n15522 = ~n15519 & n15521;
  assign n15523 = ~pi625 & ~n15517;
  assign n15524 = pi625 & n15504;
  assign n15525 = ~pi1153 & ~n15524;
  assign n15526 = ~n15523 & n15525;
  assign n15527 = ~n15522 & ~n15526;
  assign n15528 = pi778 & ~n15527;
  assign n15529 = ~n15518 & ~n15528;
  assign n15530 = ~n62880 & ~n15529;
  assign n15531 = n62880 & ~n15504;
  assign n15532 = ~n62880 & n15529;
  assign n15533 = n62880 & n15504;
  assign n15534 = ~n15532 & ~n15533;
  assign n15535 = ~n15530 & ~n15531;
  assign n15536 = ~n62882 & ~n63235;
  assign n15537 = n62882 & n15504;
  assign n15538 = n62882 & ~n15504;
  assign n15539 = ~n62882 & n63235;
  assign n15540 = ~n15538 & ~n15539;
  assign n15541 = ~n15536 & ~n15537;
  assign n15542 = ~n8257 & ~n63236;
  assign n15543 = ~n8257 & n63236;
  assign n15544 = n8257 & n15504;
  assign n15545 = ~n15543 & ~n15544;
  assign n15546 = ~n15505 & ~n15542;
  assign n15547 = ~n8303 & ~n63237;
  assign n15548 = n8303 & n15504;
  assign n15549 = ~n15547 & ~n15548;
  assign n15550 = ~pi792 & n15549;
  assign n15551 = pi628 & ~n15549;
  assign n15552 = ~pi628 & n15504;
  assign n15553 = pi1156 & ~n15552;
  assign n15554 = ~n15551 & n15553;
  assign n15555 = ~pi628 & ~n15549;
  assign n15556 = pi628 & n15504;
  assign n15557 = ~pi1156 & ~n15556;
  assign n15558 = ~n15555 & n15557;
  assign n15559 = ~n15554 & ~n15558;
  assign n15560 = pi792 & ~n15559;
  assign n15561 = ~n15550 & ~n15560;
  assign n15562 = pi647 & n15561;
  assign n15563 = ~pi647 & n15504;
  assign n15564 = pi1157 & ~n15563;
  assign n15565 = pi647 & ~n15561;
  assign n15566 = ~pi647 & ~n15504;
  assign n15567 = ~n15562 & ~n15563;
  assign n15568 = ~n15565 & ~n15566;
  assign n15569 = pi1157 & n63238;
  assign n15570 = ~n15562 & n15564;
  assign n15571 = ~pi647 & n15561;
  assign n15572 = pi647 & n15504;
  assign n15573 = ~pi1157 & ~n15572;
  assign n15574 = ~n15571 & n15573;
  assign n15575 = ~pi647 & ~n15561;
  assign n15576 = pi647 & ~n15504;
  assign n15577 = ~n15575 & ~n15576;
  assign n15578 = ~pi1157 & n15577;
  assign n15579 = pi1157 & ~n63238;
  assign n15580 = ~n15578 & ~n15579;
  assign n15581 = ~n63239 & ~n15574;
  assign n15582 = pi787 & n63240;
  assign n15583 = ~pi787 & ~n15561;
  assign n15584 = pi787 & ~n63240;
  assign n15585 = ~pi787 & n15561;
  assign n15586 = ~n15584 & ~n15585;
  assign n15587 = ~n15582 & ~n15583;
  assign n15588 = ~pi644 & ~n63241;
  assign n15589 = pi715 & ~n15588;
  assign n15590 = ~n11558 & n15504;
  assign n15591 = pi178 & ~n62765;
  assign n15592 = ~pi760 & n7359;
  assign n15593 = ~n15513 & ~n15592;
  assign n15594 = pi38 & ~n15593;
  assign n15595 = ~pi178 & n62802;
  assign n15596 = pi178 & ~n7351;
  assign n15597 = ~pi760 & ~n15596;
  assign n15598 = ~n15595 & n15597;
  assign n15599 = ~pi178 & pi760;
  assign n15600 = ~n62792 & n15599;
  assign n15601 = pi760 & ~n62792;
  assign n15602 = ~pi760 & ~n15595;
  assign n15603 = ~n15601 & ~n15602;
  assign n15604 = ~pi178 & ~n15603;
  assign n15605 = n7351 & n15602;
  assign n15606 = ~n15604 & ~n15605;
  assign n15607 = ~n15598 & ~n15600;
  assign n15608 = ~pi38 & ~n63242;
  assign n15609 = ~n15594 & ~n15608;
  assign n15610 = n62765 & n15609;
  assign n15611 = ~n15591 & ~n15610;
  assign n15612 = ~n8135 & ~n15611;
  assign n15613 = n8135 & ~n15504;
  assign n15614 = ~n15612 & ~n15613;
  assign n15615 = ~pi785 & ~n15614;
  assign n15616 = ~n8136 & ~n15504;
  assign n15617 = pi609 & n15612;
  assign n15618 = ~n15616 & ~n15617;
  assign n15619 = pi1155 & ~n15618;
  assign n15620 = ~n8148 & ~n15504;
  assign n15621 = ~pi609 & n15612;
  assign n15622 = ~n15620 & ~n15621;
  assign n15623 = ~pi1155 & ~n15622;
  assign n15624 = ~n15619 & ~n15623;
  assign n15625 = pi785 & ~n15624;
  assign n15626 = ~n15615 & ~n15625;
  assign n15627 = ~pi781 & ~n15626;
  assign n15628 = pi618 & n15626;
  assign n15629 = ~pi618 & n15504;
  assign n15630 = pi1154 & ~n15629;
  assign n15631 = ~n15628 & n15630;
  assign n15632 = ~pi618 & n15626;
  assign n15633 = pi618 & n15504;
  assign n15634 = ~pi1154 & ~n15633;
  assign n15635 = ~n15632 & n15634;
  assign n15636 = ~n15631 & ~n15635;
  assign n15637 = pi781 & ~n15636;
  assign n15638 = ~n15627 & ~n15637;
  assign n15639 = ~pi619 & ~n15638;
  assign n15640 = pi619 & ~n15504;
  assign n15641 = ~pi1159 & ~n15640;
  assign n15642 = ~n15639 & n15641;
  assign n15643 = pi619 & ~n15638;
  assign n15644 = ~pi619 & ~n15504;
  assign n15645 = pi1159 & ~n15644;
  assign n15646 = ~n15643 & n15645;
  assign n15647 = pi619 & n15638;
  assign n15648 = ~pi619 & n15504;
  assign n15649 = pi1159 & ~n15648;
  assign n15650 = ~n15647 & n15649;
  assign n15651 = ~pi619 & n15638;
  assign n15652 = pi619 & n15504;
  assign n15653 = ~pi1159 & ~n15652;
  assign n15654 = ~n15651 & n15653;
  assign n15655 = ~n15650 & ~n15654;
  assign n15656 = ~n15642 & ~n15646;
  assign n15657 = pi789 & n63243;
  assign n15658 = ~pi789 & n15638;
  assign n15659 = ~pi789 & ~n15638;
  assign n15660 = pi789 & ~n63243;
  assign n15661 = ~n15659 & ~n15660;
  assign n15662 = ~n15657 & ~n15658;
  assign n15663 = ~n8595 & n63244;
  assign n15664 = n8685 & n15663;
  assign n15665 = n8376 & ~n15504;
  assign n15666 = n8595 & n15504;
  assign n15667 = ~n15663 & ~n15666;
  assign n15668 = ~n8334 & ~n15667;
  assign n15669 = n8334 & n15504;
  assign n15670 = ~n15668 & ~n15669;
  assign n15671 = ~n8376 & n15670;
  assign n15672 = ~n15665 & ~n15671;
  assign n15673 = ~n8376 & ~n15670;
  assign n15674 = n8376 & n15504;
  assign n15675 = ~n15673 & ~n15674;
  assign n15676 = ~n15590 & ~n15664;
  assign n15677 = pi644 & n63245;
  assign n15678 = ~pi644 & n15504;
  assign n15679 = ~pi715 & ~n15678;
  assign n15680 = ~n15677 & n15679;
  assign n15681 = pi1160 & ~n15680;
  assign n15682 = ~n15589 & n15681;
  assign n15683 = pi644 & ~n63241;
  assign n15684 = ~pi715 & ~n15683;
  assign n15685 = ~pi644 & n63245;
  assign n15686 = pi644 & n15504;
  assign n15687 = pi715 & ~n15686;
  assign n15688 = ~n15685 & n15687;
  assign n15689 = ~pi1160 & ~n15688;
  assign n15690 = ~n15684 & n15689;
  assign n15691 = ~n15682 & ~n15690;
  assign n15692 = pi790 & ~n15691;
  assign n15693 = ~n63052 & n15667;
  assign n15694 = ~pi629 & n15554;
  assign n15695 = pi629 & n15558;
  assign n15696 = ~n15694 & ~n15695;
  assign n15697 = ~n15693 & n15696;
  assign n15698 = pi792 & ~n15697;
  assign n15699 = pi688 & ~n15609;
  assign n15700 = ~pi178 & ~n62821;
  assign n15701 = pi178 & n7632;
  assign n15702 = pi760 & ~n15701;
  assign n15703 = ~n15700 & n15702;
  assign n15704 = pi178 & n7709;
  assign n15705 = ~pi178 & n62851;
  assign n15706 = ~pi760 & ~n15705;
  assign n15707 = ~n15704 & n15706;
  assign n15708 = pi39 & ~n15707;
  assign n15709 = ~n15703 & n15708;
  assign n15710 = pi178 & n7855;
  assign n15711 = ~pi178 & n7832;
  assign n15712 = pi760 & ~n15711;
  assign n15713 = ~n15710 & n15712;
  assign n15714 = ~pi178 & ~n7861;
  assign n15715 = pi178 & ~n7868;
  assign n15716 = ~pi760 & ~n15715;
  assign n15717 = ~n15714 & n15716;
  assign n15718 = ~pi39 & ~n15717;
  assign n15719 = pi178 & ~n7855;
  assign n15720 = ~pi178 & ~n7832;
  assign n15721 = pi760 & ~n15720;
  assign n15722 = pi760 & ~n15719;
  assign n15723 = ~n15720 & n15722;
  assign n15724 = ~n15719 & n15721;
  assign n15725 = ~pi178 & n7861;
  assign n15726 = pi178 & n7868;
  assign n15727 = ~pi760 & ~n15726;
  assign n15728 = ~n15725 & n15727;
  assign n15729 = ~n63246 & ~n15728;
  assign n15730 = ~pi39 & ~n15729;
  assign n15731 = ~n15713 & n15718;
  assign n15732 = ~pi38 & ~n63247;
  assign n15733 = ~n15709 & n15732;
  assign n15734 = ~pi760 & ~n7744;
  assign n15735 = n10350 & ~n15734;
  assign n15736 = ~pi178 & ~n15735;
  assign n15737 = ~n7565 & ~n15277;
  assign n15738 = pi178 & ~n15737;
  assign n15739 = n7356 & n15738;
  assign n15740 = pi38 & ~n15739;
  assign n15741 = ~n15736 & n15740;
  assign n15742 = ~pi688 & ~n15741;
  assign n15743 = ~n15733 & n15742;
  assign n15744 = n62765 & ~n15743;
  assign n15745 = ~n15699 & n15744;
  assign n15746 = ~n15591 & ~n15745;
  assign n15747 = ~pi625 & n15746;
  assign n15748 = pi625 & n15611;
  assign n15749 = ~pi1153 & ~n15748;
  assign n15750 = ~n15747 & n15749;
  assign n15751 = ~pi608 & ~n15522;
  assign n15752 = ~n15750 & n15751;
  assign n15753 = pi625 & n15746;
  assign n15754 = ~pi625 & n15611;
  assign n15755 = pi1153 & ~n15754;
  assign n15756 = ~n15753 & n15755;
  assign n15757 = pi608 & ~n15526;
  assign n15758 = ~n15756 & n15757;
  assign n15759 = ~n15752 & ~n15758;
  assign n15760 = pi778 & ~n15759;
  assign n15761 = ~pi778 & n15746;
  assign n15762 = ~n15760 & ~n15761;
  assign n15763 = ~pi609 & ~n15762;
  assign n15764 = pi609 & n15529;
  assign n15765 = ~pi1155 & ~n15764;
  assign n15766 = ~n15763 & n15765;
  assign n15767 = ~pi660 & ~n15619;
  assign n15768 = ~n15766 & n15767;
  assign n15769 = pi609 & ~n15762;
  assign n15770 = ~pi609 & n15529;
  assign n15771 = pi1155 & ~n15770;
  assign n15772 = ~n15769 & n15771;
  assign n15773 = pi660 & ~n15623;
  assign n15774 = ~n15772 & n15773;
  assign n15775 = ~n15768 & ~n15774;
  assign n15776 = pi785 & ~n15775;
  assign n15777 = ~pi785 & ~n15762;
  assign n15778 = ~n15776 & ~n15777;
  assign n15779 = pi618 & ~n15778;
  assign n15780 = ~pi618 & ~n63235;
  assign n15781 = pi1154 & ~n15780;
  assign n15782 = ~n15779 & n15781;
  assign n15783 = pi627 & ~n15635;
  assign n15784 = ~n15782 & n15783;
  assign n15785 = ~pi618 & ~n15778;
  assign n15786 = pi618 & ~n63235;
  assign n15787 = ~pi1154 & ~n15786;
  assign n15788 = ~n15785 & n15787;
  assign n15789 = ~pi627 & ~n15631;
  assign n15790 = ~n15788 & n15789;
  assign n15791 = pi781 & ~n15790;
  assign n15792 = ~n15784 & n15791;
  assign n15793 = ~n11431 & ~n63236;
  assign n15794 = ~n62884 & ~n63243;
  assign n15795 = ~n15793 & ~n15794;
  assign n15796 = pi789 & ~n15795;
  assign n15797 = ~pi781 & n15778;
  assign n15798 = ~n15796 & ~n15797;
  assign n15799 = ~n15792 & n15798;
  assign n15800 = n11434 & n15795;
  assign n15801 = ~n15799 & ~n15800;
  assign n15802 = ~n15784 & ~n15790;
  assign n15803 = pi781 & ~n15802;
  assign n15804 = ~pi781 & ~n15778;
  assign n15805 = ~n15803 & ~n15804;
  assign n15806 = ~pi619 & ~n15805;
  assign n15807 = pi619 & n63236;
  assign n15808 = ~pi1159 & ~n15807;
  assign n15809 = ~n15806 & n15808;
  assign n15810 = ~pi648 & ~n15650;
  assign n15811 = ~n15809 & n15810;
  assign n15812 = pi619 & ~n15805;
  assign n15813 = ~pi619 & n63236;
  assign n15814 = pi1159 & ~n15813;
  assign n15815 = ~n15812 & n15814;
  assign n15816 = pi648 & ~n15654;
  assign n15817 = ~n15815 & n15816;
  assign n15818 = pi789 & ~n15817;
  assign n15819 = pi789 & ~n15811;
  assign n15820 = ~n15817 & n15819;
  assign n15821 = ~n15811 & n15818;
  assign n15822 = ~pi789 & n15805;
  assign n15823 = n62894 & ~n15822;
  assign n15824 = ~n63248 & n15823;
  assign n15825 = n62894 & ~n15801;
  assign n15826 = ~pi626 & ~n63244;
  assign n15827 = pi626 & ~n15504;
  assign n15828 = n8301 & ~n15827;
  assign n15829 = ~n15826 & n15828;
  assign n15830 = n8525 & ~n63237;
  assign n15831 = pi626 & ~n63244;
  assign n15832 = ~pi626 & ~n15504;
  assign n15833 = n8300 & ~n15832;
  assign n15834 = ~n15831 & n15833;
  assign n15835 = ~n15830 & ~n15834;
  assign n15836 = ~n15829 & ~n15830;
  assign n15837 = ~n15834 & n15836;
  assign n15838 = ~n15829 & n15835;
  assign n15839 = pi788 & ~n63250;
  assign n15840 = ~n63030 & ~n15839;
  assign n15841 = ~n63249 & n15840;
  assign n15842 = ~n15698 & ~n15841;
  assign n15843 = ~n8651 & ~n15842;
  assign n15844 = ~n8413 & ~n15669;
  assign n15845 = ~n8413 & n15670;
  assign n15846 = ~n15668 & n15844;
  assign n15847 = n8373 & n63238;
  assign n15848 = ~pi630 & n63239;
  assign n15849 = n8374 & ~n15577;
  assign n15850 = pi630 & n15574;
  assign n15851 = ~n63252 & ~n63253;
  assign n15852 = ~n63251 & n15851;
  assign n15853 = pi787 & ~n15852;
  assign n15854 = ~pi644 & n15689;
  assign n15855 = pi644 & n15681;
  assign n15856 = n14029 & ~n15680;
  assign n15857 = pi790 & ~n63254;
  assign n15858 = pi790 & ~n15854;
  assign n15859 = ~n63254 & n15858;
  assign n15860 = ~n15854 & n15857;
  assign n15861 = ~n15853 & ~n63255;
  assign n15862 = ~n15843 & ~n15853;
  assign n15863 = ~n63255 & n15862;
  assign n15864 = ~n15843 & n15861;
  assign n15865 = ~n15692 & ~n63256;
  assign n15866 = n62455 & ~n15865;
  assign n15867 = ~pi178 & ~n62455;
  assign n15868 = ~pi832 & ~n15867;
  assign n15869 = ~n15866 & n15868;
  assign po335 = ~n15503 & ~n15869;
  assign n15871 = ~pi179 & ~n2923;
  assign n15872 = ~pi741 & n7316;
  assign n15873 = ~n15871 & ~n15872;
  assign n15874 = ~n8420 & ~n15873;
  assign n15875 = ~pi785 & ~n15874;
  assign n15876 = ~n8425 & ~n15873;
  assign n15877 = pi1155 & ~n15876;
  assign n15878 = ~n8428 & n15874;
  assign n15879 = ~pi1155 & ~n15878;
  assign n15880 = ~n15877 & ~n15879;
  assign n15881 = pi785 & ~n15880;
  assign n15882 = ~n15875 & ~n15881;
  assign n15883 = ~pi781 & ~n15882;
  assign n15884 = ~n8435 & n15882;
  assign n15885 = pi1154 & ~n15884;
  assign n15886 = ~n8438 & n15882;
  assign n15887 = ~pi1154 & ~n15886;
  assign n15888 = ~n15885 & ~n15887;
  assign n15889 = pi781 & ~n15888;
  assign n15890 = ~n15883 & ~n15889;
  assign n15891 = ~pi619 & ~n15890;
  assign n15892 = pi619 & ~n15871;
  assign n15893 = ~pi1159 & ~n15892;
  assign n15894 = ~n15891 & n15893;
  assign n15895 = pi619 & ~n15890;
  assign n15896 = ~pi619 & ~n15871;
  assign n15897 = pi1159 & ~n15896;
  assign n15898 = ~n15895 & n15897;
  assign n15899 = pi619 & n15890;
  assign n15900 = ~pi619 & n15871;
  assign n15901 = pi1159 & ~n15900;
  assign n15902 = ~n15899 & n15901;
  assign n15903 = ~pi619 & n15890;
  assign n15904 = pi619 & n15871;
  assign n15905 = ~pi1159 & ~n15904;
  assign n15906 = ~n15903 & n15905;
  assign n15907 = ~n15902 & ~n15906;
  assign n15908 = ~n15894 & ~n15898;
  assign n15909 = pi789 & n63257;
  assign n15910 = ~pi789 & n15890;
  assign n15911 = ~pi789 & ~n15890;
  assign n15912 = pi789 & ~n63257;
  assign n15913 = ~n15911 & ~n15912;
  assign n15914 = ~n15909 & ~n15910;
  assign n15915 = ~n8595 & n63258;
  assign n15916 = n8595 & n15871;
  assign n15917 = ~n8595 & ~n63258;
  assign n15918 = n8595 & ~n15871;
  assign n15919 = ~n15917 & ~n15918;
  assign n15920 = ~n15915 & ~n15916;
  assign n15921 = ~n8334 & n63259;
  assign n15922 = n8334 & n15871;
  assign n15923 = ~n8413 & ~n15922;
  assign n15924 = ~n15921 & ~n15922;
  assign n15925 = ~n8413 & n15924;
  assign n15926 = ~n15921 & n15923;
  assign n15927 = ~pi724 & n7564;
  assign n15928 = ~n15871 & ~n15927;
  assign n15929 = ~pi778 & n15928;
  assign n15930 = ~pi625 & n15927;
  assign n15931 = ~n15928 & ~n15930;
  assign n15932 = pi1153 & ~n15931;
  assign n15933 = ~pi1153 & ~n15871;
  assign n15934 = ~n15930 & n15933;
  assign n15935 = ~n15932 & ~n15934;
  assign n15936 = pi778 & ~n15935;
  assign n15937 = ~n15929 & ~n15936;
  assign n15938 = ~n8490 & n15937;
  assign n15939 = ~n8492 & n15938;
  assign n15940 = ~n8494 & n15939;
  assign n15941 = ~n8496 & n15940;
  assign n15942 = ~n8508 & n15941;
  assign n15943 = pi647 & ~n15942;
  assign n15944 = ~pi647 & ~n15871;
  assign n15945 = ~n15943 & ~n15944;
  assign n15946 = n8373 & ~n15945;
  assign n15947 = ~pi647 & n15942;
  assign n15948 = pi647 & n15871;
  assign n15949 = ~pi1157 & ~n15948;
  assign n15950 = ~n15947 & n15949;
  assign n15951 = pi630 & n15950;
  assign n15952 = ~n15946 & ~n15951;
  assign n15953 = ~n63260 & n15952;
  assign n15954 = pi787 & ~n15953;
  assign n15955 = ~pi626 & ~n63258;
  assign n15956 = pi626 & ~n15871;
  assign n15957 = n8301 & ~n15956;
  assign n15958 = ~n15955 & n15957;
  assign n15959 = n8525 & n15940;
  assign n15960 = pi626 & ~n63258;
  assign n15961 = ~pi626 & ~n15871;
  assign n15962 = n8300 & ~n15961;
  assign n15963 = ~n15960 & n15962;
  assign n15964 = ~n15959 & ~n15963;
  assign n15965 = ~n15958 & ~n15959;
  assign n15966 = ~n15963 & n15965;
  assign n15967 = ~n15958 & n15964;
  assign n15968 = pi788 & ~n63261;
  assign n15969 = ~n7187 & ~n15928;
  assign n15970 = pi625 & n15969;
  assign n15971 = n15873 & ~n15969;
  assign n15972 = ~n15970 & ~n15971;
  assign n15973 = n15933 & ~n15972;
  assign n15974 = ~pi608 & ~n15932;
  assign n15975 = ~n15973 & n15974;
  assign n15976 = pi1153 & n15873;
  assign n15977 = ~n15970 & n15976;
  assign n15978 = pi608 & ~n15934;
  assign n15979 = ~n15977 & n15978;
  assign n15980 = ~n15975 & ~n15979;
  assign n15981 = pi778 & ~n15980;
  assign n15982 = ~pi778 & ~n15971;
  assign n15983 = ~n15981 & ~n15982;
  assign n15984 = ~pi609 & ~n15983;
  assign n15985 = pi609 & n15937;
  assign n15986 = ~pi1155 & ~n15985;
  assign n15987 = ~n15984 & n15986;
  assign n15988 = ~pi660 & ~n15877;
  assign n15989 = ~n15987 & n15988;
  assign n15990 = pi609 & ~n15983;
  assign n15991 = ~pi609 & n15937;
  assign n15992 = pi1155 & ~n15991;
  assign n15993 = ~n15990 & n15992;
  assign n15994 = pi660 & ~n15879;
  assign n15995 = ~n15993 & n15994;
  assign n15996 = ~n15989 & ~n15995;
  assign n15997 = pi785 & ~n15996;
  assign n15998 = ~pi785 & ~n15983;
  assign n15999 = ~n15997 & ~n15998;
  assign n16000 = pi618 & ~n15999;
  assign n16001 = ~pi618 & n15938;
  assign n16002 = pi1154 & ~n16001;
  assign n16003 = ~n16000 & n16002;
  assign n16004 = pi627 & ~n15887;
  assign n16005 = ~n16003 & n16004;
  assign n16006 = ~pi618 & ~n15999;
  assign n16007 = pi618 & n15938;
  assign n16008 = ~pi1154 & ~n16007;
  assign n16009 = ~n16006 & n16008;
  assign n16010 = ~pi627 & ~n15885;
  assign n16011 = ~n16009 & n16010;
  assign n16012 = pi781 & ~n16011;
  assign n16013 = ~n16005 & n16012;
  assign n16014 = ~n11431 & ~n15939;
  assign n16015 = ~n62884 & ~n63257;
  assign n16016 = ~n16014 & ~n16015;
  assign n16017 = pi789 & ~n16016;
  assign n16018 = ~pi781 & n15999;
  assign n16019 = ~n16017 & ~n16018;
  assign n16020 = ~n16013 & n16019;
  assign n16021 = n11434 & n16016;
  assign n16022 = ~n16020 & ~n16021;
  assign n16023 = ~n16005 & ~n16011;
  assign n16024 = pi781 & ~n16023;
  assign n16025 = ~pi781 & ~n15999;
  assign n16026 = ~n16024 & ~n16025;
  assign n16027 = ~pi619 & ~n16026;
  assign n16028 = pi619 & n15939;
  assign n16029 = ~pi1159 & ~n16028;
  assign n16030 = ~n16027 & n16029;
  assign n16031 = ~pi648 & ~n15902;
  assign n16032 = ~n16030 & n16031;
  assign n16033 = pi619 & ~n16026;
  assign n16034 = ~pi619 & n15939;
  assign n16035 = pi1159 & ~n16034;
  assign n16036 = ~n16033 & n16035;
  assign n16037 = pi648 & ~n15906;
  assign n16038 = ~n16036 & n16037;
  assign n16039 = pi789 & ~n16038;
  assign n16040 = pi789 & ~n16032;
  assign n16041 = ~n16038 & n16040;
  assign n16042 = ~n16032 & n16039;
  assign n16043 = ~pi789 & n16026;
  assign n16044 = n62894 & ~n16043;
  assign n16045 = ~n63262 & n16044;
  assign n16046 = n62894 & ~n16022;
  assign n16047 = ~n15968 & ~n63263;
  assign n16048 = ~n63030 & ~n16047;
  assign n16049 = n8498 & n63259;
  assign n16050 = n8615 & n15941;
  assign n16051 = pi629 & ~n16050;
  assign n16052 = ~n16049 & n16051;
  assign n16053 = n8499 & n63259;
  assign n16054 = n8606 & n15941;
  assign n16055 = ~pi629 & ~n16054;
  assign n16056 = ~n16053 & n16055;
  assign n16057 = pi792 & ~n16056;
  assign n16058 = pi792 & ~n16052;
  assign n16059 = ~n16056 & n16058;
  assign n16060 = ~n16053 & ~n16054;
  assign n16061 = ~pi629 & ~n16060;
  assign n16062 = ~n16049 & ~n16050;
  assign n16063 = pi629 & ~n16062;
  assign n16064 = ~n16061 & ~n16063;
  assign n16065 = pi792 & ~n16064;
  assign n16066 = ~n16052 & n16057;
  assign n16067 = ~n8651 & ~n63264;
  assign n16068 = ~n16048 & n16067;
  assign n16069 = ~n15954 & ~n16068;
  assign n16070 = pi644 & n16069;
  assign n16071 = ~pi787 & ~n15942;
  assign n16072 = pi1157 & ~n15945;
  assign n16073 = ~n15950 & ~n16072;
  assign n16074 = pi787 & ~n16073;
  assign n16075 = ~n16071 & ~n16074;
  assign n16076 = ~pi644 & n16075;
  assign n16077 = pi715 & ~n16076;
  assign n16078 = ~n16070 & n16077;
  assign n16079 = ~n8685 & n15871;
  assign n16080 = ~n8376 & n15921;
  assign n16081 = ~n8376 & ~n15924;
  assign n16082 = n8376 & n15871;
  assign n16083 = ~n16081 & ~n16082;
  assign n16084 = ~n16079 & ~n16080;
  assign n16085 = pi644 & ~n63265;
  assign n16086 = ~pi644 & n15871;
  assign n16087 = ~pi715 & ~n16086;
  assign n16088 = ~n16085 & n16087;
  assign n16089 = pi1160 & ~n16088;
  assign n16090 = ~n16078 & n16089;
  assign n16091 = ~pi644 & n16069;
  assign n16092 = pi644 & n16075;
  assign n16093 = ~pi715 & ~n16092;
  assign n16094 = ~n16091 & n16093;
  assign n16095 = ~pi644 & ~n63265;
  assign n16096 = pi644 & n15871;
  assign n16097 = pi715 & ~n16096;
  assign n16098 = ~n16095 & n16097;
  assign n16099 = ~pi1160 & ~n16098;
  assign n16100 = ~n16094 & n16099;
  assign n16101 = ~n16090 & ~n16100;
  assign n16102 = pi790 & ~n16101;
  assign n16103 = ~pi790 & n16069;
  assign n16104 = pi832 & ~n16103;
  assign n16105 = ~n16102 & n16104;
  assign n16106 = pi179 & ~n62765;
  assign n16107 = pi741 & n8091;
  assign n16108 = ~pi741 & ~n14285;
  assign n16109 = pi179 & ~n16108;
  assign n16110 = ~pi179 & ~pi741;
  assign n16111 = ~n62977 & n16110;
  assign n16112 = n10343 & n16111;
  assign n16113 = n10343 & n16110;
  assign n16114 = ~n16109 & ~n63266;
  assign n16115 = ~n16107 & n16114;
  assign n16116 = n62765 & ~n16115;
  assign n16117 = ~n16106 & ~n16116;
  assign n16118 = ~n8135 & ~n16117;
  assign n16119 = ~pi179 & ~n8098;
  assign n16120 = n8135 & ~n16119;
  assign n16121 = ~n16118 & ~n16120;
  assign n16122 = ~pi785 & ~n16121;
  assign n16123 = ~n8136 & ~n16119;
  assign n16124 = pi609 & n16118;
  assign n16125 = ~n16123 & ~n16124;
  assign n16126 = pi1155 & ~n16125;
  assign n16127 = ~n8148 & ~n16119;
  assign n16128 = ~pi609 & n16118;
  assign n16129 = ~n16127 & ~n16128;
  assign n16130 = ~pi1155 & ~n16129;
  assign n16131 = ~n16126 & ~n16130;
  assign n16132 = pi785 & ~n16131;
  assign n16133 = ~n16122 & ~n16132;
  assign n16134 = ~pi781 & ~n16133;
  assign n16135 = pi618 & n16133;
  assign n16136 = ~pi618 & n16119;
  assign n16137 = pi1154 & ~n16136;
  assign n16138 = ~n16135 & n16137;
  assign n16139 = ~pi618 & n16133;
  assign n16140 = pi618 & n16119;
  assign n16141 = ~pi1154 & ~n16140;
  assign n16142 = ~n16139 & n16141;
  assign n16143 = ~n16138 & ~n16142;
  assign n16144 = pi781 & ~n16143;
  assign n16145 = ~n16134 & ~n16144;
  assign n16146 = ~pi789 & ~n16145;
  assign n16147 = ~pi619 & n16145;
  assign n16148 = pi619 & n16119;
  assign n16149 = ~pi1159 & ~n16148;
  assign n16150 = ~n16147 & n16149;
  assign n16151 = pi619 & n16145;
  assign n16152 = ~pi619 & n16119;
  assign n16153 = pi1159 & ~n16152;
  assign n16154 = ~n16151 & n16153;
  assign n16155 = ~n16150 & ~n16154;
  assign n16156 = pi789 & ~n16155;
  assign n16157 = ~n16146 & ~n16156;
  assign n16158 = ~n8595 & n16157;
  assign n16159 = n8595 & n16119;
  assign n16160 = ~n16158 & ~n16159;
  assign n16161 = ~n8334 & ~n16160;
  assign n16162 = n8334 & n16119;
  assign n16163 = ~n16161 & ~n16162;
  assign n16164 = ~n8376 & ~n16163;
  assign n16165 = n8376 & n16119;
  assign n16166 = n8376 & ~n16119;
  assign n16167 = ~n8376 & n16163;
  assign n16168 = ~n16166 & ~n16167;
  assign n16169 = ~n16164 & ~n16165;
  assign n16170 = ~pi644 & n63267;
  assign n16171 = pi644 & n16119;
  assign n16172 = pi715 & ~pi1160;
  assign n16173 = ~n16171 & n16172;
  assign n16174 = ~n16170 & n16173;
  assign n16175 = pi644 & n63267;
  assign n16176 = ~pi644 & n16119;
  assign n16177 = ~pi715 & pi1160;
  assign n16178 = ~n16176 & n16177;
  assign n16179 = ~n16175 & n16178;
  assign n16180 = n8257 & ~n16119;
  assign n16181 = ~pi724 & n62765;
  assign n16182 = n16119 & ~n16181;
  assign n16183 = ~pi179 & n8009;
  assign n16184 = pi179 & n62874;
  assign n16185 = ~pi38 & ~n16184;
  assign n16186 = n62765 & ~n16185;
  assign n16187 = ~n16183 & ~n16186;
  assign n16188 = ~pi179 & ~n7357;
  assign n16189 = n8085 & ~n16188;
  assign n16190 = ~pi724 & ~n16189;
  assign n16191 = ~n16187 & n16190;
  assign n16192 = ~n16182 & ~n16191;
  assign n16193 = ~pi778 & n16192;
  assign n16194 = ~pi625 & ~n16192;
  assign n16195 = pi625 & n16119;
  assign n16196 = ~pi1153 & ~n16195;
  assign n16197 = ~n16194 & n16196;
  assign n16198 = pi625 & ~n16192;
  assign n16199 = ~pi625 & n16119;
  assign n16200 = pi1153 & ~n16199;
  assign n16201 = ~n16198 & n16200;
  assign n16202 = ~n16197 & ~n16201;
  assign n16203 = pi778 & ~n16202;
  assign n16204 = ~n16193 & ~n16203;
  assign n16205 = ~n62880 & ~n16204;
  assign n16206 = n62880 & ~n16119;
  assign n16207 = ~n62880 & n16204;
  assign n16208 = n62880 & n16119;
  assign n16209 = ~n16207 & ~n16208;
  assign n16210 = ~n16205 & ~n16206;
  assign n16211 = ~n62882 & ~n63268;
  assign n16212 = n62882 & n16119;
  assign n16213 = n62882 & ~n16119;
  assign n16214 = ~n62882 & n63268;
  assign n16215 = ~n16213 & ~n16214;
  assign n16216 = ~n16211 & ~n16212;
  assign n16217 = ~n8257 & ~n63269;
  assign n16218 = ~n8257 & n63269;
  assign n16219 = n8257 & n16119;
  assign n16220 = ~n16218 & ~n16219;
  assign n16221 = ~n16180 & ~n16217;
  assign n16222 = ~n8303 & ~n63270;
  assign n16223 = n8303 & n16119;
  assign n16224 = n8303 & ~n16119;
  assign n16225 = ~n8303 & n63270;
  assign n16226 = ~n16224 & ~n16225;
  assign n16227 = ~n16222 & ~n16223;
  assign n16228 = ~n62892 & n63271;
  assign n16229 = n62892 & n16119;
  assign n16230 = pi628 & n63271;
  assign n16231 = ~pi628 & n16119;
  assign n16232 = pi1156 & ~n16231;
  assign n16233 = ~n16230 & n16232;
  assign n16234 = ~pi628 & n63271;
  assign n16235 = pi628 & n16119;
  assign n16236 = ~pi1156 & ~n16235;
  assign n16237 = ~n16234 & n16236;
  assign n16238 = pi628 & ~n16119;
  assign n16239 = ~pi628 & ~n63271;
  assign n16240 = ~n16238 & ~n16239;
  assign n16241 = ~pi1156 & n16240;
  assign n16242 = ~pi628 & ~n16119;
  assign n16243 = pi628 & ~n63271;
  assign n16244 = ~n16242 & ~n16243;
  assign n16245 = pi1156 & n16244;
  assign n16246 = ~n16241 & ~n16245;
  assign n16247 = ~n16233 & ~n16237;
  assign n16248 = pi792 & ~n63272;
  assign n16249 = ~pi792 & n63271;
  assign n16250 = ~n16248 & ~n16249;
  assign n16251 = ~pi792 & ~n63271;
  assign n16252 = pi792 & n63272;
  assign n16253 = ~n16251 & ~n16252;
  assign n16254 = ~n16228 & ~n16229;
  assign n16255 = ~pi647 & ~n63273;
  assign n16256 = pi647 & n16119;
  assign n16257 = ~pi1157 & ~n16256;
  assign n16258 = ~n16255 & n16257;
  assign n16259 = pi647 & ~n63273;
  assign n16260 = ~pi647 & n16119;
  assign n16261 = pi1157 & ~n16260;
  assign n16262 = ~n16259 & ~n16260;
  assign n16263 = pi1157 & n16262;
  assign n16264 = ~n16259 & n16261;
  assign n16265 = pi787 & ~n63274;
  assign n16266 = ~n16258 & n16265;
  assign n16267 = ~pi787 & ~n63273;
  assign n16268 = ~n63036 & ~n16267;
  assign n16269 = ~n16266 & n16268;
  assign n16270 = ~n16179 & ~n16269;
  assign n16271 = ~n16174 & n16270;
  assign n16272 = pi790 & ~n16271;
  assign n16273 = ~n8413 & n16163;
  assign n16274 = n8373 & n16262;
  assign n16275 = ~pi630 & n63274;
  assign n16276 = pi630 & n16258;
  assign n16277 = ~n63275 & ~n16276;
  assign n16278 = ~n16273 & ~n16276;
  assign n16279 = ~n63275 & n16278;
  assign n16280 = ~n16273 & n16277;
  assign n16281 = pi787 & ~n63276;
  assign n16282 = ~n63052 & n16160;
  assign n16283 = n8332 & ~n16235;
  assign n16284 = n8332 & ~n16240;
  assign n16285 = ~n16234 & n16283;
  assign n16286 = n8331 & ~n16231;
  assign n16287 = n8331 & ~n16244;
  assign n16288 = ~n16230 & n16286;
  assign n16289 = ~n63277 & ~n63278;
  assign n16290 = ~n16282 & n16289;
  assign n16291 = pi792 & ~n16290;
  assign n16292 = n12979 & n16157;
  assign n16293 = ~pi641 & n63270;
  assign n16294 = pi641 & ~n16119;
  assign n16295 = n8417 & ~n16294;
  assign n16296 = ~n16293 & n16295;
  assign n16297 = pi641 & n63270;
  assign n16298 = ~pi641 & ~n16119;
  assign n16299 = n8416 & ~n16298;
  assign n16300 = ~n16297 & n16299;
  assign n16301 = ~n16296 & ~n16300;
  assign n16302 = ~n16292 & n16301;
  assign n16303 = pi788 & ~n16302;
  assign n16304 = pi619 & n63269;
  assign n16305 = ~pi1159 & ~n16304;
  assign n16306 = ~pi648 & ~n16154;
  assign n16307 = ~n16305 & n16306;
  assign n16308 = ~pi619 & n63269;
  assign n16309 = pi1159 & ~n16308;
  assign n16310 = pi648 & ~n16309;
  assign n16311 = pi648 & ~n16150;
  assign n16312 = ~n16309 & n16311;
  assign n16313 = ~n16150 & n16310;
  assign n16314 = ~n16307 & ~n63279;
  assign n16315 = pi789 & ~n16314;
  assign n16316 = pi618 & ~n63268;
  assign n16317 = ~pi1154 & ~n16316;
  assign n16318 = ~pi627 & ~n16138;
  assign n16319 = ~n16317 & n16318;
  assign n16320 = ~pi618 & ~n63268;
  assign n16321 = pi1154 & ~n16320;
  assign n16322 = pi627 & ~n16142;
  assign n16323 = ~n16321 & n16322;
  assign n16324 = ~n16319 & ~n16323;
  assign n16325 = pi781 & ~n16324;
  assign n16326 = ~pi618 & n16318;
  assign n16327 = pi618 & n16322;
  assign n16328 = pi781 & ~n16327;
  assign n16329 = ~n16326 & n16328;
  assign n16330 = n8793 & ~n16188;
  assign n16331 = ~pi179 & n8759;
  assign n16332 = pi179 & n8763;
  assign n16333 = ~pi38 & ~n16332;
  assign n16334 = ~pi179 & ~n62821;
  assign n16335 = pi179 & n7632;
  assign n16336 = pi39 & ~n16335;
  assign n16337 = ~n16334 & n16336;
  assign n16338 = ~pi179 & n7832;
  assign n16339 = pi179 & n7855;
  assign n16340 = ~pi39 & ~n16339;
  assign n16341 = ~pi39 & ~n16338;
  assign n16342 = ~n16339 & n16341;
  assign n16343 = ~n16338 & n16340;
  assign n16344 = ~n16337 & ~n63280;
  assign n16345 = ~pi38 & ~n16344;
  assign n16346 = ~n16331 & n16333;
  assign n16347 = ~n16330 & ~n63281;
  assign n16348 = pi741 & ~n16347;
  assign n16349 = pi179 & n10363;
  assign n16350 = ~pi179 & ~n62980;
  assign n16351 = ~pi741 & ~n16350;
  assign n16352 = ~n16349 & n16351;
  assign n16353 = ~pi724 & ~n16352;
  assign n16354 = ~n16348 & n16353;
  assign n16355 = pi724 & n16115;
  assign n16356 = n62765 & ~n16355;
  assign n16357 = ~n16354 & n16356;
  assign n16358 = ~n16106 & ~n16357;
  assign n16359 = pi625 & n16358;
  assign n16360 = ~pi625 & n16117;
  assign n16361 = pi1153 & ~n16360;
  assign n16362 = ~n16359 & n16361;
  assign n16363 = pi608 & ~n16197;
  assign n16364 = ~n16362 & n16363;
  assign n16365 = ~pi625 & n16358;
  assign n16366 = pi625 & n16117;
  assign n16367 = ~pi1153 & ~n16366;
  assign n16368 = ~n16365 & n16367;
  assign n16369 = ~pi608 & ~n16201;
  assign n16370 = ~n16368 & n16369;
  assign n16371 = ~n16364 & ~n16370;
  assign n16372 = pi778 & ~n16371;
  assign n16373 = ~pi778 & n16358;
  assign n16374 = ~pi778 & ~n16358;
  assign n16375 = pi778 & ~n16370;
  assign n16376 = ~n16364 & n16375;
  assign n16377 = ~n16374 & ~n16376;
  assign n16378 = ~n16372 & ~n16373;
  assign n16379 = ~pi785 & ~n63282;
  assign n16380 = ~pi609 & n63282;
  assign n16381 = pi609 & n16204;
  assign n16382 = ~pi1155 & ~n16381;
  assign n16383 = ~n16380 & n16382;
  assign n16384 = ~pi660 & ~n16126;
  assign n16385 = ~n16383 & n16384;
  assign n16386 = pi609 & n63282;
  assign n16387 = ~pi609 & n16204;
  assign n16388 = pi1155 & ~n16387;
  assign n16389 = ~n16386 & n16388;
  assign n16390 = pi660 & ~n16130;
  assign n16391 = ~n16389 & n16390;
  assign n16392 = pi785 & ~n16391;
  assign n16393 = ~n16385 & n16392;
  assign n16394 = ~n16385 & ~n16391;
  assign n16395 = pi785 & ~n16394;
  assign n16396 = ~pi785 & n63282;
  assign n16397 = ~n16395 & ~n16396;
  assign n16398 = ~n16379 & ~n16393;
  assign n16399 = ~n16329 & ~n63283;
  assign n16400 = pi618 & ~n63283;
  assign n16401 = n16321 & ~n16400;
  assign n16402 = n16322 & ~n16401;
  assign n16403 = ~n16319 & ~n16402;
  assign n16404 = pi781 & ~n16403;
  assign n16405 = pi781 & ~n16326;
  assign n16406 = ~n63283 & ~n16405;
  assign n16407 = ~n16404 & ~n16406;
  assign n16408 = ~pi618 & ~n63283;
  assign n16409 = n16317 & ~n16408;
  assign n16410 = n16318 & ~n16409;
  assign n16411 = ~n16402 & ~n16410;
  assign n16412 = pi781 & ~n16411;
  assign n16413 = ~pi781 & ~n63283;
  assign n16414 = ~n16412 & ~n16413;
  assign n16415 = ~n16325 & ~n16399;
  assign n16416 = ~pi619 & n16306;
  assign n16417 = pi619 & n16311;
  assign n16418 = n11422 & ~n16150;
  assign n16419 = pi789 & ~n63285;
  assign n16420 = ~n16416 & n16419;
  assign n16421 = ~n63284 & ~n16420;
  assign n16422 = ~pi619 & ~n63284;
  assign n16423 = n16305 & ~n16422;
  assign n16424 = n16306 & ~n16423;
  assign n16425 = pi619 & ~n63284;
  assign n16426 = n16309 & ~n16425;
  assign n16427 = n16311 & ~n16426;
  assign n16428 = ~n16424 & ~n16427;
  assign n16429 = pi789 & ~n16428;
  assign n16430 = ~pi789 & ~n63284;
  assign n16431 = ~n16429 & ~n16430;
  assign n16432 = ~n16315 & ~n16421;
  assign n16433 = n62894 & ~n63286;
  assign n16434 = ~n63030 & ~n16433;
  assign n16435 = ~n16303 & n16434;
  assign n16436 = ~pi788 & n63286;
  assign n16437 = ~pi626 & n63286;
  assign n16438 = pi626 & n63270;
  assign n16439 = ~pi641 & ~n16438;
  assign n16440 = ~n16437 & n16439;
  assign n16441 = ~pi626 & ~n16157;
  assign n16442 = pi626 & ~n16119;
  assign n16443 = pi641 & ~n16442;
  assign n16444 = ~n16441 & n16443;
  assign n16445 = ~pi1158 & ~n16444;
  assign n16446 = ~n16440 & n16445;
  assign n16447 = pi626 & n63286;
  assign n16448 = ~pi626 & n63270;
  assign n16449 = pi641 & ~n16448;
  assign n16450 = ~n16447 & n16449;
  assign n16451 = pi626 & ~n16157;
  assign n16452 = ~pi626 & ~n16119;
  assign n16453 = ~pi641 & ~n16452;
  assign n16454 = ~n16451 & n16453;
  assign n16455 = pi1158 & ~n16454;
  assign n16456 = ~n16450 & n16455;
  assign n16457 = ~n16446 & ~n16456;
  assign n16458 = pi788 & ~n16457;
  assign n16459 = ~n16436 & ~n16458;
  assign n16460 = ~n16303 & ~n16433;
  assign n16461 = ~pi628 & n63287;
  assign n16462 = pi628 & ~n16160;
  assign n16463 = ~pi1156 & ~n16462;
  assign n16464 = ~n16461 & n16463;
  assign n16465 = ~pi629 & ~n16233;
  assign n16466 = ~n16464 & n16465;
  assign n16467 = pi628 & n63287;
  assign n16468 = ~pi628 & ~n16160;
  assign n16469 = pi1156 & ~n16468;
  assign n16470 = ~n16467 & n16469;
  assign n16471 = pi629 & ~n16237;
  assign n16472 = ~n16470 & n16471;
  assign n16473 = ~n16466 & ~n16472;
  assign n16474 = pi792 & ~n16473;
  assign n16475 = ~pi792 & n63287;
  assign n16476 = ~n16474 & ~n16475;
  assign n16477 = ~n16291 & ~n16435;
  assign n16478 = ~n16291 & n63287;
  assign n16479 = n63030 & n16290;
  assign n16480 = ~n8651 & ~n16479;
  assign n16481 = ~n16478 & n16480;
  assign n16482 = ~n8651 & n63288;
  assign n16483 = ~pi647 & ~n63288;
  assign n16484 = pi647 & ~n16163;
  assign n16485 = ~pi1157 & ~n16484;
  assign n16486 = ~n16483 & n16485;
  assign n16487 = ~pi630 & ~n63274;
  assign n16488 = ~n16486 & n16487;
  assign n16489 = pi647 & ~n63288;
  assign n16490 = ~pi647 & ~n16163;
  assign n16491 = pi1157 & ~n16490;
  assign n16492 = ~n16489 & n16491;
  assign n16493 = pi630 & ~n16258;
  assign n16494 = ~n16492 & n16493;
  assign n16495 = ~n16488 & ~n16494;
  assign n16496 = pi787 & ~n16495;
  assign n16497 = ~pi787 & ~n63288;
  assign n16498 = ~n16496 & ~n16497;
  assign n16499 = ~n16281 & ~n63289;
  assign n16500 = ~n11547 & n63290;
  assign n16501 = n62455 & ~n16500;
  assign n16502 = ~pi644 & ~n63290;
  assign n16503 = ~pi787 & n63273;
  assign n16504 = ~n16258 & ~n63274;
  assign n16505 = pi787 & ~n16504;
  assign n16506 = ~n16503 & ~n16505;
  assign n16507 = pi644 & n16506;
  assign n16508 = ~pi715 & ~n16507;
  assign n16509 = ~n16502 & n16508;
  assign n16510 = pi715 & ~n16171;
  assign n16511 = ~n16170 & n16510;
  assign n16512 = ~pi1160 & ~n16511;
  assign n16513 = ~n16509 & n16512;
  assign n16514 = ~pi644 & n16506;
  assign n16515 = pi715 & ~n16514;
  assign n16516 = ~pi715 & ~n16176;
  assign n16517 = ~n16175 & n16516;
  assign n16518 = pi1160 & ~n16517;
  assign n16519 = ~n16515 & n16518;
  assign n16520 = ~n16513 & ~n16519;
  assign n16521 = pi790 & ~n16520;
  assign n16522 = pi644 & n16518;
  assign n16523 = pi790 & ~n16522;
  assign n16524 = ~n63290 & ~n16523;
  assign n16525 = ~n16521 & ~n16524;
  assign n16526 = n62455 & ~n16525;
  assign n16527 = pi644 & ~n63290;
  assign n16528 = n16515 & ~n16527;
  assign n16529 = n16518 & ~n16528;
  assign n16530 = pi790 & ~n16513;
  assign n16531 = pi790 & ~n16529;
  assign n16532 = ~n16513 & n16531;
  assign n16533 = ~n16529 & n16530;
  assign n16534 = ~pi790 & n63290;
  assign n16535 = n62455 & ~n16534;
  assign n16536 = ~n63292 & n16535;
  assign n16537 = ~n16272 & n16501;
  assign n16538 = ~pi179 & ~n62455;
  assign n16539 = ~pi832 & ~n16538;
  assign n16540 = ~n63291 & n16539;
  assign po336 = ~n16105 & ~n16540;
  assign n16542 = ~pi180 & ~n2923;
  assign n16543 = ~pi753 & n7316;
  assign n16544 = ~n16542 & ~n16543;
  assign n16545 = ~n8420 & ~n16544;
  assign n16546 = ~pi785 & ~n16545;
  assign n16547 = n8148 & n16543;
  assign n16548 = n16545 & ~n16547;
  assign n16549 = pi1155 & ~n16548;
  assign n16550 = ~pi1155 & ~n16542;
  assign n16551 = ~n16547 & n16550;
  assign n16552 = ~n16549 & ~n16551;
  assign n16553 = pi785 & ~n16552;
  assign n16554 = ~n16546 & ~n16553;
  assign n16555 = ~pi781 & ~n16554;
  assign n16556 = ~n8435 & n16554;
  assign n16557 = pi1154 & ~n16556;
  assign n16558 = ~n8438 & n16554;
  assign n16559 = ~pi1154 & ~n16558;
  assign n16560 = ~n16557 & ~n16559;
  assign n16561 = pi781 & ~n16560;
  assign n16562 = ~n16555 & ~n16561;
  assign n16563 = ~pi789 & ~n16562;
  assign n16564 = ~n12612 & n16562;
  assign n16565 = pi1159 & ~n16564;
  assign n16566 = ~n12615 & n16562;
  assign n16567 = ~pi1159 & ~n16566;
  assign n16568 = ~n16565 & ~n16567;
  assign n16569 = pi789 & ~n16568;
  assign n16570 = ~n16563 & ~n16569;
  assign n16571 = ~n15298 & n16562;
  assign n16572 = ~n8595 & n63293;
  assign n16573 = n8595 & n16542;
  assign n16574 = ~n8595 & ~n63293;
  assign n16575 = n8595 & ~n16542;
  assign n16576 = ~n16574 & ~n16575;
  assign n16577 = ~n16572 & ~n16573;
  assign n16578 = ~n8334 & n63294;
  assign n16579 = n8334 & n16542;
  assign n16580 = ~n8413 & ~n16579;
  assign n16581 = ~n16578 & ~n16579;
  assign n16582 = ~n8413 & n16581;
  assign n16583 = ~n16578 & n16580;
  assign n16584 = ~pi702 & n7564;
  assign n16585 = ~n16542 & ~n16584;
  assign n16586 = ~pi778 & ~n16585;
  assign n16587 = ~pi625 & n16584;
  assign n16588 = ~n16585 & ~n16587;
  assign n16589 = pi1153 & ~n16588;
  assign n16590 = ~pi1153 & ~n16542;
  assign n16591 = ~n16587 & n16590;
  assign n16592 = pi778 & ~n16591;
  assign n16593 = ~n16589 & n16592;
  assign n16594 = ~n16586 & ~n16593;
  assign n16595 = ~n8490 & ~n16594;
  assign n16596 = ~n8492 & n16595;
  assign n16597 = ~n8494 & n16596;
  assign n16598 = ~n8496 & n16597;
  assign n16599 = ~n8508 & n16598;
  assign n16600 = pi647 & ~n16599;
  assign n16601 = ~pi647 & ~n16542;
  assign n16602 = ~n16600 & ~n16601;
  assign n16603 = n8373 & ~n16602;
  assign n16604 = ~pi647 & n16599;
  assign n16605 = pi647 & n16542;
  assign n16606 = ~pi1157 & ~n16605;
  assign n16607 = ~n16604 & n16606;
  assign n16608 = pi630 & n16607;
  assign n16609 = ~n16603 & ~n16608;
  assign n16610 = ~n63295 & n16609;
  assign n16611 = pi787 & ~n16610;
  assign n16612 = ~pi626 & ~n63293;
  assign n16613 = pi626 & ~n16542;
  assign n16614 = n8301 & ~n16613;
  assign n16615 = ~n16612 & n16614;
  assign n16616 = n8525 & n16597;
  assign n16617 = pi626 & ~n63293;
  assign n16618 = ~pi626 & ~n16542;
  assign n16619 = n8300 & ~n16618;
  assign n16620 = ~n16617 & n16619;
  assign n16621 = ~n16616 & ~n16620;
  assign n16622 = ~n16615 & ~n16616;
  assign n16623 = ~n16620 & n16622;
  assign n16624 = ~n16615 & n16621;
  assign n16625 = pi788 & ~n63296;
  assign n16626 = n13460 & n16562;
  assign n16627 = n11303 & n16596;
  assign n16628 = pi648 & ~n16627;
  assign n16629 = ~n16626 & n16628;
  assign n16630 = n13462 & n16562;
  assign n16631 = n11304 & n16596;
  assign n16632 = ~pi648 & ~n16631;
  assign n16633 = ~n16630 & n16632;
  assign n16634 = pi789 & ~n16633;
  assign n16635 = ~n16629 & n16634;
  assign n16636 = ~n7187 & ~n16585;
  assign n16637 = pi625 & n16636;
  assign n16638 = n16544 & ~n16636;
  assign n16639 = ~n16637 & ~n16638;
  assign n16640 = n16590 & ~n16639;
  assign n16641 = ~pi608 & ~n16589;
  assign n16642 = ~n16640 & n16641;
  assign n16643 = pi1153 & n16544;
  assign n16644 = ~n16637 & n16643;
  assign n16645 = pi608 & ~n16591;
  assign n16646 = ~n16644 & n16645;
  assign n16647 = ~n16642 & ~n16646;
  assign n16648 = pi778 & ~n16647;
  assign n16649 = ~pi778 & ~n16638;
  assign n16650 = ~n16648 & ~n16649;
  assign n16651 = ~pi609 & ~n16650;
  assign n16652 = pi609 & ~n16594;
  assign n16653 = ~pi1155 & ~n16652;
  assign n16654 = ~n16651 & n16653;
  assign n16655 = ~pi660 & ~n16549;
  assign n16656 = ~n16654 & n16655;
  assign n16657 = pi609 & ~n16650;
  assign n16658 = ~pi609 & ~n16594;
  assign n16659 = pi1155 & ~n16658;
  assign n16660 = ~n16657 & n16659;
  assign n16661 = pi660 & ~n16551;
  assign n16662 = ~n16660 & n16661;
  assign n16663 = ~n16656 & ~n16662;
  assign n16664 = pi785 & ~n16663;
  assign n16665 = ~pi785 & ~n16650;
  assign n16666 = ~n16664 & ~n16665;
  assign n16667 = pi618 & ~n16666;
  assign n16668 = ~pi618 & n16595;
  assign n16669 = pi1154 & ~n16668;
  assign n16670 = ~n16667 & n16669;
  assign n16671 = pi627 & ~n16559;
  assign n16672 = ~n16670 & n16671;
  assign n16673 = ~pi618 & ~n16666;
  assign n16674 = pi618 & n16595;
  assign n16675 = ~pi1154 & ~n16674;
  assign n16676 = ~n16673 & n16675;
  assign n16677 = ~pi627 & ~n16557;
  assign n16678 = ~n16676 & n16677;
  assign n16679 = pi781 & ~n16678;
  assign n16680 = ~n16672 & n16679;
  assign n16681 = ~pi781 & n16666;
  assign n16682 = ~n11434 & ~n16681;
  assign n16683 = ~n16680 & n16682;
  assign n16684 = ~n16635 & ~n16683;
  assign n16685 = ~n16672 & ~n16678;
  assign n16686 = pi781 & ~n16685;
  assign n16687 = ~pi781 & ~n16666;
  assign n16688 = ~n16686 & ~n16687;
  assign n16689 = ~pi619 & ~n16688;
  assign n16690 = pi619 & n16596;
  assign n16691 = ~pi1159 & ~n16690;
  assign n16692 = ~n16689 & n16691;
  assign n16693 = ~pi648 & ~n16565;
  assign n16694 = ~n16692 & n16693;
  assign n16695 = pi619 & ~n16688;
  assign n16696 = ~pi619 & n16596;
  assign n16697 = pi1159 & ~n16696;
  assign n16698 = ~n16695 & n16697;
  assign n16699 = pi648 & ~n16567;
  assign n16700 = ~n16698 & n16699;
  assign n16701 = pi789 & ~n16700;
  assign n16702 = pi789 & ~n16694;
  assign n16703 = ~n16700 & n16702;
  assign n16704 = ~n16694 & n16701;
  assign n16705 = ~pi789 & n16688;
  assign n16706 = n62894 & ~n16705;
  assign n16707 = ~n63297 & n16706;
  assign n16708 = n62894 & ~n16684;
  assign n16709 = ~n16625 & ~n63298;
  assign n16710 = ~n63030 & ~n16709;
  assign n16711 = n8498 & n63294;
  assign n16712 = n8615 & n16598;
  assign n16713 = pi629 & ~n16712;
  assign n16714 = ~n16711 & n16713;
  assign n16715 = n8499 & n63294;
  assign n16716 = n8606 & n16598;
  assign n16717 = ~pi629 & ~n16716;
  assign n16718 = ~n16715 & n16717;
  assign n16719 = pi792 & ~n16718;
  assign n16720 = pi792 & ~n16714;
  assign n16721 = ~n16718 & n16720;
  assign n16722 = ~n16715 & ~n16716;
  assign n16723 = ~pi629 & ~n16722;
  assign n16724 = ~n16711 & ~n16712;
  assign n16725 = pi629 & ~n16724;
  assign n16726 = ~n16723 & ~n16725;
  assign n16727 = pi792 & ~n16726;
  assign n16728 = ~n16714 & n16719;
  assign n16729 = ~n8651 & ~n63299;
  assign n16730 = ~n16710 & n16729;
  assign n16731 = ~n16611 & ~n16730;
  assign n16732 = pi644 & n16731;
  assign n16733 = ~pi787 & ~n16599;
  assign n16734 = pi1157 & ~n16602;
  assign n16735 = ~n16607 & ~n16734;
  assign n16736 = pi787 & ~n16735;
  assign n16737 = ~n16733 & ~n16736;
  assign n16738 = ~pi644 & n16737;
  assign n16739 = pi715 & ~n16738;
  assign n16740 = ~n16732 & n16739;
  assign n16741 = ~n8685 & n16542;
  assign n16742 = ~n8376 & n16578;
  assign n16743 = ~n8376 & ~n16581;
  assign n16744 = n8376 & n16542;
  assign n16745 = ~n16743 & ~n16744;
  assign n16746 = ~n16741 & ~n16742;
  assign n16747 = pi644 & ~n63300;
  assign n16748 = ~pi644 & n16542;
  assign n16749 = ~pi715 & ~n16748;
  assign n16750 = ~n16747 & n16749;
  assign n16751 = pi1160 & ~n16750;
  assign n16752 = ~n16740 & n16751;
  assign n16753 = ~pi644 & n16731;
  assign n16754 = pi644 & n16737;
  assign n16755 = ~pi715 & ~n16754;
  assign n16756 = ~n16753 & n16755;
  assign n16757 = ~pi644 & ~n63300;
  assign n16758 = pi644 & n16542;
  assign n16759 = pi715 & ~n16758;
  assign n16760 = ~n16757 & n16759;
  assign n16761 = ~pi1160 & ~n16760;
  assign n16762 = ~n16756 & n16761;
  assign n16763 = ~n16752 & ~n16762;
  assign n16764 = pi790 & ~n16763;
  assign n16765 = ~pi790 & n16731;
  assign n16766 = pi832 & ~n16765;
  assign n16767 = ~n16764 & n16766;
  assign n16768 = ~pi180 & ~n8098;
  assign n16769 = n8257 & ~n16768;
  assign n16770 = ~pi702 & n62765;
  assign n16771 = n16768 & ~n16770;
  assign n16772 = pi180 & n62874;
  assign n16773 = ~pi38 & ~n16772;
  assign n16774 = n62765 & ~n16773;
  assign n16775 = ~pi180 & n8009;
  assign n16776 = ~n16774 & ~n16775;
  assign n16777 = ~pi180 & ~n7357;
  assign n16778 = n8085 & ~n16777;
  assign n16779 = ~pi702 & ~n16778;
  assign n16780 = ~n16776 & n16779;
  assign n16781 = ~n16771 & ~n16780;
  assign n16782 = ~pi778 & n16781;
  assign n16783 = pi625 & ~n16781;
  assign n16784 = ~pi625 & n16768;
  assign n16785 = pi1153 & ~n16784;
  assign n16786 = ~n16783 & n16785;
  assign n16787 = ~pi625 & ~n16781;
  assign n16788 = pi625 & n16768;
  assign n16789 = ~pi1153 & ~n16788;
  assign n16790 = ~n16787 & n16789;
  assign n16791 = ~n16786 & ~n16790;
  assign n16792 = pi778 & ~n16791;
  assign n16793 = ~n16782 & ~n16792;
  assign n16794 = ~n62880 & ~n16793;
  assign n16795 = n62880 & ~n16768;
  assign n16796 = ~n62880 & n16793;
  assign n16797 = n62880 & n16768;
  assign n16798 = ~n16796 & ~n16797;
  assign n16799 = ~n16794 & ~n16795;
  assign n16800 = ~n62882 & ~n63301;
  assign n16801 = n62882 & n16768;
  assign n16802 = n62882 & ~n16768;
  assign n16803 = ~n62882 & n63301;
  assign n16804 = ~n16802 & ~n16803;
  assign n16805 = ~n16800 & ~n16801;
  assign n16806 = ~n8257 & ~n63302;
  assign n16807 = ~n8257 & n63302;
  assign n16808 = n8257 & n16768;
  assign n16809 = ~n16807 & ~n16808;
  assign n16810 = ~n16769 & ~n16806;
  assign n16811 = ~n8303 & ~n63303;
  assign n16812 = n8303 & n16768;
  assign n16813 = ~n16811 & ~n16812;
  assign n16814 = ~pi792 & n16813;
  assign n16815 = pi628 & ~n16813;
  assign n16816 = ~pi628 & n16768;
  assign n16817 = pi1156 & ~n16816;
  assign n16818 = ~n16815 & n16817;
  assign n16819 = ~pi628 & ~n16813;
  assign n16820 = pi628 & n16768;
  assign n16821 = ~pi1156 & ~n16820;
  assign n16822 = ~n16819 & n16821;
  assign n16823 = ~n16818 & ~n16822;
  assign n16824 = pi792 & ~n16823;
  assign n16825 = ~n16814 & ~n16824;
  assign n16826 = pi647 & n16825;
  assign n16827 = ~pi647 & n16768;
  assign n16828 = pi1157 & ~n16827;
  assign n16829 = pi647 & ~n16825;
  assign n16830 = ~pi647 & ~n16768;
  assign n16831 = ~n16826 & ~n16827;
  assign n16832 = ~n16829 & ~n16830;
  assign n16833 = pi1157 & n63304;
  assign n16834 = ~n16826 & n16828;
  assign n16835 = ~pi647 & n16825;
  assign n16836 = pi647 & n16768;
  assign n16837 = ~pi1157 & ~n16836;
  assign n16838 = ~n16835 & n16837;
  assign n16839 = ~pi647 & ~n16825;
  assign n16840 = pi647 & ~n16768;
  assign n16841 = ~n16839 & ~n16840;
  assign n16842 = ~pi1157 & n16841;
  assign n16843 = pi1157 & ~n63304;
  assign n16844 = ~n16842 & ~n16843;
  assign n16845 = ~n63305 & ~n16838;
  assign n16846 = pi787 & n63306;
  assign n16847 = ~pi787 & ~n16825;
  assign n16848 = pi787 & ~n63306;
  assign n16849 = ~pi787 & n16825;
  assign n16850 = ~n16848 & ~n16849;
  assign n16851 = ~n16846 & ~n16847;
  assign n16852 = ~pi644 & ~n63307;
  assign n16853 = pi715 & ~n16852;
  assign n16854 = ~n11558 & n16768;
  assign n16855 = pi180 & ~n62765;
  assign n16856 = pi753 & n7143;
  assign n16857 = pi180 & n7349;
  assign n16858 = ~n16856 & ~n16857;
  assign n16859 = pi39 & ~n16858;
  assign n16860 = ~pi180 & ~pi753;
  assign n16861 = n62802 & n16860;
  assign n16862 = pi180 & pi753;
  assign n16863 = pi753 & ~n62781;
  assign n16864 = pi180 & ~n7292;
  assign n16865 = ~n16863 & ~n16864;
  assign n16866 = ~pi39 & ~n16865;
  assign n16867 = ~n16862 & ~n16866;
  assign n16868 = ~n16861 & n16867;
  assign n16869 = ~n16859 & n16868;
  assign n16870 = ~pi38 & ~n16869;
  assign n16871 = ~pi753 & n7359;
  assign n16872 = pi38 & ~n16777;
  assign n16873 = ~n16871 & n16872;
  assign n16874 = ~n16870 & ~n16873;
  assign n16875 = n62765 & ~n16874;
  assign n16876 = ~n16855 & ~n16875;
  assign n16877 = ~n8135 & ~n16876;
  assign n16878 = n8135 & ~n16768;
  assign n16879 = ~n16877 & ~n16878;
  assign n16880 = ~pi785 & ~n16879;
  assign n16881 = ~n8136 & ~n16768;
  assign n16882 = pi609 & n16877;
  assign n16883 = ~n16881 & ~n16882;
  assign n16884 = pi1155 & ~n16883;
  assign n16885 = ~n8148 & ~n16768;
  assign n16886 = ~pi609 & n16877;
  assign n16887 = ~n16885 & ~n16886;
  assign n16888 = ~pi1155 & ~n16887;
  assign n16889 = ~n16884 & ~n16888;
  assign n16890 = pi785 & ~n16889;
  assign n16891 = ~n16880 & ~n16890;
  assign n16892 = ~pi781 & ~n16891;
  assign n16893 = pi618 & n16891;
  assign n16894 = ~pi618 & n16768;
  assign n16895 = pi1154 & ~n16894;
  assign n16896 = ~n16893 & n16895;
  assign n16897 = ~pi618 & n16891;
  assign n16898 = pi618 & n16768;
  assign n16899 = ~pi1154 & ~n16898;
  assign n16900 = ~n16897 & n16899;
  assign n16901 = ~n16896 & ~n16900;
  assign n16902 = pi781 & ~n16901;
  assign n16903 = ~n16892 & ~n16902;
  assign n16904 = ~pi619 & ~n16903;
  assign n16905 = pi619 & ~n16768;
  assign n16906 = ~pi1159 & ~n16905;
  assign n16907 = ~n16904 & n16906;
  assign n16908 = pi619 & ~n16903;
  assign n16909 = ~pi619 & ~n16768;
  assign n16910 = pi1159 & ~n16909;
  assign n16911 = ~n16908 & n16910;
  assign n16912 = pi619 & n16903;
  assign n16913 = ~pi619 & n16768;
  assign n16914 = pi1159 & ~n16913;
  assign n16915 = ~n16912 & n16914;
  assign n16916 = ~pi619 & n16903;
  assign n16917 = pi619 & n16768;
  assign n16918 = ~pi1159 & ~n16917;
  assign n16919 = ~n16916 & n16918;
  assign n16920 = ~n16915 & ~n16919;
  assign n16921 = ~n16907 & ~n16911;
  assign n16922 = pi789 & n63308;
  assign n16923 = ~pi789 & n16903;
  assign n16924 = ~pi789 & ~n16903;
  assign n16925 = pi789 & ~n63308;
  assign n16926 = ~n16924 & ~n16925;
  assign n16927 = ~n16922 & ~n16923;
  assign n16928 = ~n8595 & n63309;
  assign n16929 = n8685 & n16928;
  assign n16930 = n8376 & ~n16768;
  assign n16931 = n8595 & n16768;
  assign n16932 = ~n16928 & ~n16931;
  assign n16933 = ~n8334 & ~n16932;
  assign n16934 = n8334 & n16768;
  assign n16935 = ~n16933 & ~n16934;
  assign n16936 = ~n8376 & n16935;
  assign n16937 = ~n16930 & ~n16936;
  assign n16938 = ~n8376 & ~n16935;
  assign n16939 = n8376 & n16768;
  assign n16940 = ~n16938 & ~n16939;
  assign n16941 = ~n16854 & ~n16929;
  assign n16942 = pi644 & n63310;
  assign n16943 = ~pi644 & n16768;
  assign n16944 = ~pi715 & ~n16943;
  assign n16945 = ~n16942 & n16944;
  assign n16946 = pi1160 & ~n16945;
  assign n16947 = ~n16853 & n16946;
  assign n16948 = pi644 & ~n63307;
  assign n16949 = ~pi715 & ~n16948;
  assign n16950 = ~pi644 & n63310;
  assign n16951 = pi644 & n16768;
  assign n16952 = pi715 & ~n16951;
  assign n16953 = ~n16950 & n16952;
  assign n16954 = ~pi1160 & ~n16953;
  assign n16955 = ~n16949 & n16954;
  assign n16956 = ~n16947 & ~n16955;
  assign n16957 = pi790 & ~n16956;
  assign n16958 = ~n63052 & n16932;
  assign n16959 = ~pi629 & n16818;
  assign n16960 = pi629 & n16822;
  assign n16961 = ~n16959 & ~n16960;
  assign n16962 = ~n16958 & n16961;
  assign n16963 = pi792 & ~n16962;
  assign n16964 = ~pi626 & ~n63309;
  assign n16965 = pi626 & ~n16768;
  assign n16966 = n8301 & ~n16965;
  assign n16967 = ~n16964 & n16966;
  assign n16968 = n8525 & ~n63303;
  assign n16969 = pi626 & ~n63309;
  assign n16970 = ~pi626 & ~n16768;
  assign n16971 = n8300 & ~n16970;
  assign n16972 = ~n16969 & n16971;
  assign n16973 = ~n16968 & ~n16972;
  assign n16974 = ~n16967 & ~n16968;
  assign n16975 = ~n16972 & n16974;
  assign n16976 = ~n16967 & n16973;
  assign n16977 = pi788 & ~n63311;
  assign n16978 = pi702 & n16874;
  assign n16979 = ~pi180 & ~n62821;
  assign n16980 = pi180 & n7632;
  assign n16981 = pi753 & ~n16980;
  assign n16982 = ~n16979 & n16981;
  assign n16983 = pi180 & n7709;
  assign n16984 = ~pi180 & n62851;
  assign n16985 = ~pi753 & ~n16984;
  assign n16986 = ~n16983 & n16985;
  assign n16987 = pi39 & ~n16986;
  assign n16988 = ~n16982 & n16987;
  assign n16989 = pi180 & n7855;
  assign n16990 = ~pi180 & n7832;
  assign n16991 = pi753 & ~n16990;
  assign n16992 = ~n16989 & n16991;
  assign n16993 = ~pi180 & ~n7861;
  assign n16994 = pi180 & ~n7868;
  assign n16995 = ~pi753 & ~n16994;
  assign n16996 = ~n16993 & n16995;
  assign n16997 = ~pi39 & ~n16996;
  assign n16998 = pi180 & ~n7855;
  assign n16999 = ~pi180 & ~n7832;
  assign n17000 = pi753 & ~n16999;
  assign n17001 = pi753 & ~n16998;
  assign n17002 = ~n16999 & n17001;
  assign n17003 = ~n16998 & n17000;
  assign n17004 = ~pi180 & n7861;
  assign n17005 = pi180 & n7868;
  assign n17006 = ~pi753 & ~n17005;
  assign n17007 = ~n17004 & n17006;
  assign n17008 = ~n63312 & ~n17007;
  assign n17009 = ~pi39 & ~n17008;
  assign n17010 = ~n16992 & n16997;
  assign n17011 = ~pi38 & ~n63313;
  assign n17012 = ~n16988 & n17011;
  assign n17013 = ~pi753 & ~n7744;
  assign n17014 = n10350 & ~n17013;
  assign n17015 = ~pi180 & ~n17014;
  assign n17016 = ~n7565 & ~n16543;
  assign n17017 = pi180 & ~n17016;
  assign n17018 = n7356 & n17017;
  assign n17019 = pi38 & ~n17018;
  assign n17020 = ~n17015 & n17019;
  assign n17021 = ~pi702 & ~n17020;
  assign n17022 = ~n17012 & n17021;
  assign n17023 = n62765 & ~n17022;
  assign n17024 = ~n16978 & n17023;
  assign n17025 = ~n16855 & ~n17024;
  assign n17026 = ~pi625 & n17025;
  assign n17027 = pi625 & n16876;
  assign n17028 = ~pi1153 & ~n17027;
  assign n17029 = ~n17026 & n17028;
  assign n17030 = ~pi608 & ~n16786;
  assign n17031 = ~n17029 & n17030;
  assign n17032 = pi625 & n17025;
  assign n17033 = ~pi625 & n16876;
  assign n17034 = pi1153 & ~n17033;
  assign n17035 = ~n17032 & n17034;
  assign n17036 = pi608 & ~n16790;
  assign n17037 = ~n17035 & n17036;
  assign n17038 = ~n17031 & ~n17037;
  assign n17039 = pi778 & ~n17038;
  assign n17040 = ~pi778 & n17025;
  assign n17041 = ~n17039 & ~n17040;
  assign n17042 = ~pi609 & ~n17041;
  assign n17043 = pi609 & n16793;
  assign n17044 = ~pi1155 & ~n17043;
  assign n17045 = ~n17042 & n17044;
  assign n17046 = ~pi660 & ~n16884;
  assign n17047 = ~n17045 & n17046;
  assign n17048 = pi609 & ~n17041;
  assign n17049 = ~pi609 & n16793;
  assign n17050 = pi1155 & ~n17049;
  assign n17051 = ~n17048 & n17050;
  assign n17052 = pi660 & ~n16888;
  assign n17053 = ~n17051 & n17052;
  assign n17054 = ~n17047 & ~n17053;
  assign n17055 = pi785 & ~n17054;
  assign n17056 = ~pi785 & ~n17041;
  assign n17057 = ~n17055 & ~n17056;
  assign n17058 = ~pi781 & n17057;
  assign n17059 = ~pi618 & ~n17057;
  assign n17060 = pi618 & ~n63301;
  assign n17061 = ~pi1154 & ~n17060;
  assign n17062 = ~n17059 & n17061;
  assign n17063 = ~pi627 & ~n16896;
  assign n17064 = ~n17062 & n17063;
  assign n17065 = pi618 & ~n17057;
  assign n17066 = ~pi618 & ~n63301;
  assign n17067 = pi1154 & ~n17066;
  assign n17068 = ~n17065 & n17067;
  assign n17069 = pi627 & ~n16900;
  assign n17070 = ~n17068 & n17069;
  assign n17071 = pi781 & ~n17070;
  assign n17072 = ~n17064 & n17071;
  assign n17073 = ~n17064 & ~n17070;
  assign n17074 = pi781 & ~n17073;
  assign n17075 = ~pi781 & ~n17057;
  assign n17076 = ~n17074 & ~n17075;
  assign n17077 = ~n17058 & ~n17072;
  assign n17078 = ~n11434 & n63314;
  assign n17079 = ~n11431 & ~n63302;
  assign n17080 = ~n62884 & ~n63308;
  assign n17081 = ~n17079 & ~n17080;
  assign n17082 = pi789 & ~n17081;
  assign n17083 = n62894 & ~n17082;
  assign n17084 = ~pi619 & ~n63314;
  assign n17085 = pi619 & n63302;
  assign n17086 = ~pi1159 & ~n17085;
  assign n17087 = ~n17084 & n17086;
  assign n17088 = ~pi648 & ~n16915;
  assign n17089 = ~n17087 & n17088;
  assign n17090 = pi619 & ~n63314;
  assign n17091 = ~pi619 & n63302;
  assign n17092 = pi1159 & ~n17091;
  assign n17093 = ~n17090 & n17092;
  assign n17094 = pi648 & ~n16919;
  assign n17095 = ~n17093 & n17094;
  assign n17096 = pi789 & ~n17095;
  assign n17097 = pi789 & ~n17089;
  assign n17098 = ~n17095 & n17097;
  assign n17099 = ~n17089 & n17096;
  assign n17100 = ~pi789 & n63314;
  assign n17101 = n62894 & ~n17100;
  assign n17102 = ~n63315 & n17101;
  assign n17103 = ~n17078 & n17083;
  assign n17104 = ~n63030 & ~n63316;
  assign n17105 = ~n63030 & ~n16977;
  assign n17106 = ~n63316 & n17105;
  assign n17107 = ~n16977 & n17104;
  assign n17108 = ~n16963 & ~n63317;
  assign n17109 = ~n8651 & ~n17108;
  assign n17110 = ~n8413 & ~n16934;
  assign n17111 = ~n8413 & n16935;
  assign n17112 = ~n16933 & n17110;
  assign n17113 = n8373 & n63304;
  assign n17114 = ~pi630 & n63305;
  assign n17115 = n8374 & ~n16841;
  assign n17116 = pi630 & n16838;
  assign n17117 = ~n63319 & ~n63320;
  assign n17118 = ~n63318 & n17117;
  assign n17119 = pi787 & ~n17118;
  assign n17120 = ~pi644 & n16954;
  assign n17121 = pi644 & n16946;
  assign n17122 = n14029 & ~n16945;
  assign n17123 = pi790 & ~n63321;
  assign n17124 = pi790 & ~n17120;
  assign n17125 = ~n63321 & n17124;
  assign n17126 = ~n17120 & n17123;
  assign n17127 = ~n17119 & ~n63322;
  assign n17128 = ~n17109 & ~n17119;
  assign n17129 = ~n63322 & n17128;
  assign n17130 = ~n17109 & n17127;
  assign n17131 = ~n16957 & ~n63323;
  assign n17132 = n62455 & ~n17131;
  assign n17133 = ~pi180 & ~n62455;
  assign n17134 = ~pi832 & ~n17133;
  assign n17135 = ~n17132 & n17134;
  assign po337 = ~n16767 & ~n17135;
  assign n17137 = ~pi181 & ~n2923;
  assign n17138 = ~pi754 & n7316;
  assign n17139 = ~n17137 & ~n17138;
  assign n17140 = ~n8420 & ~n17139;
  assign n17141 = ~pi785 & ~n17140;
  assign n17142 = n8148 & n17138;
  assign n17143 = n17140 & ~n17142;
  assign n17144 = pi1155 & ~n17143;
  assign n17145 = ~pi1155 & ~n17137;
  assign n17146 = ~n17142 & n17145;
  assign n17147 = ~n17144 & ~n17146;
  assign n17148 = pi785 & ~n17147;
  assign n17149 = ~n17141 & ~n17148;
  assign n17150 = ~pi781 & ~n17149;
  assign n17151 = ~n8435 & n17149;
  assign n17152 = pi1154 & ~n17151;
  assign n17153 = ~n8438 & n17149;
  assign n17154 = ~pi1154 & ~n17153;
  assign n17155 = ~n17152 & ~n17154;
  assign n17156 = pi781 & ~n17155;
  assign n17157 = ~n17150 & ~n17156;
  assign n17158 = ~pi789 & ~n17157;
  assign n17159 = ~n12612 & n17157;
  assign n17160 = pi1159 & ~n17159;
  assign n17161 = ~n12615 & n17157;
  assign n17162 = ~pi1159 & ~n17161;
  assign n17163 = ~n17160 & ~n17162;
  assign n17164 = pi789 & ~n17163;
  assign n17165 = ~n17158 & ~n17164;
  assign n17166 = ~n15298 & n17157;
  assign n17167 = ~n8595 & n63324;
  assign n17168 = n8595 & n17137;
  assign n17169 = ~n8595 & ~n63324;
  assign n17170 = n8595 & ~n17137;
  assign n17171 = ~n17169 & ~n17170;
  assign n17172 = ~n17167 & ~n17168;
  assign n17173 = ~n8334 & n63325;
  assign n17174 = n8334 & n17137;
  assign n17175 = ~n8413 & ~n17174;
  assign n17176 = ~n17173 & ~n17174;
  assign n17177 = ~n8413 & n17176;
  assign n17178 = ~n17173 & n17175;
  assign n17179 = ~pi709 & n7564;
  assign n17180 = ~n17137 & ~n17179;
  assign n17181 = ~pi778 & ~n17180;
  assign n17182 = ~pi625 & n17179;
  assign n17183 = ~n17180 & ~n17182;
  assign n17184 = pi1153 & ~n17183;
  assign n17185 = ~pi1153 & ~n17137;
  assign n17186 = ~n17182 & n17185;
  assign n17187 = pi778 & ~n17186;
  assign n17188 = ~n17184 & n17187;
  assign n17189 = ~n17181 & ~n17188;
  assign n17190 = ~n8490 & ~n17189;
  assign n17191 = ~n8492 & n17190;
  assign n17192 = ~n8494 & n17191;
  assign n17193 = ~n8496 & n17192;
  assign n17194 = ~n8508 & n17193;
  assign n17195 = pi647 & ~n17194;
  assign n17196 = ~pi647 & ~n17137;
  assign n17197 = ~n17195 & ~n17196;
  assign n17198 = n8373 & ~n17197;
  assign n17199 = ~pi647 & n17194;
  assign n17200 = pi647 & n17137;
  assign n17201 = ~pi1157 & ~n17200;
  assign n17202 = ~n17199 & n17201;
  assign n17203 = pi630 & n17202;
  assign n17204 = ~n17198 & ~n17203;
  assign n17205 = ~n63326 & n17204;
  assign n17206 = pi787 & ~n17205;
  assign n17207 = ~pi626 & ~n63324;
  assign n17208 = pi626 & ~n17137;
  assign n17209 = n8301 & ~n17208;
  assign n17210 = ~n17207 & n17209;
  assign n17211 = n8525 & n17192;
  assign n17212 = pi626 & ~n63324;
  assign n17213 = ~pi626 & ~n17137;
  assign n17214 = n8300 & ~n17213;
  assign n17215 = ~n17212 & n17214;
  assign n17216 = ~n17211 & ~n17215;
  assign n17217 = ~n17210 & ~n17211;
  assign n17218 = ~n17215 & n17217;
  assign n17219 = ~n17210 & n17216;
  assign n17220 = pi788 & ~n63327;
  assign n17221 = n13460 & n17157;
  assign n17222 = n11303 & n17191;
  assign n17223 = pi648 & ~n17222;
  assign n17224 = ~n17221 & n17223;
  assign n17225 = n13462 & n17157;
  assign n17226 = n11304 & n17191;
  assign n17227 = ~pi648 & ~n17226;
  assign n17228 = ~n17225 & n17227;
  assign n17229 = pi789 & ~n17228;
  assign n17230 = ~n17224 & n17229;
  assign n17231 = ~n7187 & ~n17180;
  assign n17232 = pi625 & n17231;
  assign n17233 = n17139 & ~n17231;
  assign n17234 = ~n17232 & ~n17233;
  assign n17235 = n17185 & ~n17234;
  assign n17236 = ~pi608 & ~n17184;
  assign n17237 = ~n17235 & n17236;
  assign n17238 = pi1153 & n17139;
  assign n17239 = ~n17232 & n17238;
  assign n17240 = pi608 & ~n17186;
  assign n17241 = ~n17239 & n17240;
  assign n17242 = ~n17237 & ~n17241;
  assign n17243 = pi778 & ~n17242;
  assign n17244 = ~pi778 & ~n17233;
  assign n17245 = ~n17243 & ~n17244;
  assign n17246 = ~pi609 & ~n17245;
  assign n17247 = pi609 & ~n17189;
  assign n17248 = ~pi1155 & ~n17247;
  assign n17249 = ~n17246 & n17248;
  assign n17250 = ~pi660 & ~n17144;
  assign n17251 = ~n17249 & n17250;
  assign n17252 = pi609 & ~n17245;
  assign n17253 = ~pi609 & ~n17189;
  assign n17254 = pi1155 & ~n17253;
  assign n17255 = ~n17252 & n17254;
  assign n17256 = pi660 & ~n17146;
  assign n17257 = ~n17255 & n17256;
  assign n17258 = ~n17251 & ~n17257;
  assign n17259 = pi785 & ~n17258;
  assign n17260 = ~pi785 & ~n17245;
  assign n17261 = ~n17259 & ~n17260;
  assign n17262 = pi618 & ~n17261;
  assign n17263 = ~pi618 & n17190;
  assign n17264 = pi1154 & ~n17263;
  assign n17265 = ~n17262 & n17264;
  assign n17266 = pi627 & ~n17154;
  assign n17267 = ~n17265 & n17266;
  assign n17268 = ~pi618 & ~n17261;
  assign n17269 = pi618 & n17190;
  assign n17270 = ~pi1154 & ~n17269;
  assign n17271 = ~n17268 & n17270;
  assign n17272 = ~pi627 & ~n17152;
  assign n17273 = ~n17271 & n17272;
  assign n17274 = pi781 & ~n17273;
  assign n17275 = ~n17267 & n17274;
  assign n17276 = ~pi781 & n17261;
  assign n17277 = ~n11434 & ~n17276;
  assign n17278 = ~n17275 & n17277;
  assign n17279 = ~n17230 & ~n17278;
  assign n17280 = ~n17267 & ~n17273;
  assign n17281 = pi781 & ~n17280;
  assign n17282 = ~pi781 & ~n17261;
  assign n17283 = ~n17281 & ~n17282;
  assign n17284 = ~pi619 & ~n17283;
  assign n17285 = pi619 & n17191;
  assign n17286 = ~pi1159 & ~n17285;
  assign n17287 = ~n17284 & n17286;
  assign n17288 = ~pi648 & ~n17160;
  assign n17289 = ~n17287 & n17288;
  assign n17290 = pi619 & ~n17283;
  assign n17291 = ~pi619 & n17191;
  assign n17292 = pi1159 & ~n17291;
  assign n17293 = ~n17290 & n17292;
  assign n17294 = pi648 & ~n17162;
  assign n17295 = ~n17293 & n17294;
  assign n17296 = pi789 & ~n17295;
  assign n17297 = pi789 & ~n17289;
  assign n17298 = ~n17295 & n17297;
  assign n17299 = ~n17289 & n17296;
  assign n17300 = ~pi789 & n17283;
  assign n17301 = n62894 & ~n17300;
  assign n17302 = ~n63328 & n17301;
  assign n17303 = n62894 & ~n17279;
  assign n17304 = ~n17220 & ~n63329;
  assign n17305 = ~n63030 & ~n17304;
  assign n17306 = n8498 & n63325;
  assign n17307 = n8615 & n17193;
  assign n17308 = pi629 & ~n17307;
  assign n17309 = ~n17306 & n17308;
  assign n17310 = n8499 & n63325;
  assign n17311 = n8606 & n17193;
  assign n17312 = ~pi629 & ~n17311;
  assign n17313 = ~n17310 & n17312;
  assign n17314 = pi792 & ~n17313;
  assign n17315 = pi792 & ~n17309;
  assign n17316 = ~n17313 & n17315;
  assign n17317 = ~n17310 & ~n17311;
  assign n17318 = ~pi629 & ~n17317;
  assign n17319 = ~n17306 & ~n17307;
  assign n17320 = pi629 & ~n17319;
  assign n17321 = ~n17318 & ~n17320;
  assign n17322 = pi792 & ~n17321;
  assign n17323 = ~n17309 & n17314;
  assign n17324 = ~n8651 & ~n63330;
  assign n17325 = ~n17305 & n17324;
  assign n17326 = ~n17206 & ~n17325;
  assign n17327 = pi644 & n17326;
  assign n17328 = ~pi787 & ~n17194;
  assign n17329 = pi1157 & ~n17197;
  assign n17330 = ~n17202 & ~n17329;
  assign n17331 = pi787 & ~n17330;
  assign n17332 = ~n17328 & ~n17331;
  assign n17333 = ~pi644 & n17332;
  assign n17334 = pi715 & ~n17333;
  assign n17335 = ~n17327 & n17334;
  assign n17336 = ~n8685 & n17137;
  assign n17337 = ~n8376 & n17173;
  assign n17338 = ~n8376 & ~n17176;
  assign n17339 = n8376 & n17137;
  assign n17340 = ~n17338 & ~n17339;
  assign n17341 = ~n17336 & ~n17337;
  assign n17342 = pi644 & ~n63331;
  assign n17343 = ~pi644 & n17137;
  assign n17344 = ~pi715 & ~n17343;
  assign n17345 = ~n17342 & n17344;
  assign n17346 = pi1160 & ~n17345;
  assign n17347 = ~n17335 & n17346;
  assign n17348 = ~pi644 & n17326;
  assign n17349 = pi644 & n17332;
  assign n17350 = ~pi715 & ~n17349;
  assign n17351 = ~n17348 & n17350;
  assign n17352 = ~pi644 & ~n63331;
  assign n17353 = pi644 & n17137;
  assign n17354 = pi715 & ~n17353;
  assign n17355 = ~n17352 & n17354;
  assign n17356 = ~pi1160 & ~n17355;
  assign n17357 = ~n17351 & n17356;
  assign n17358 = ~n17347 & ~n17357;
  assign n17359 = pi790 & ~n17358;
  assign n17360 = ~pi790 & n17326;
  assign n17361 = pi832 & ~n17360;
  assign n17362 = ~n17359 & n17361;
  assign n17363 = ~pi181 & ~n8098;
  assign n17364 = n8257 & ~n17363;
  assign n17365 = ~pi709 & n62765;
  assign n17366 = n17363 & ~n17365;
  assign n17367 = pi181 & n62874;
  assign n17368 = ~pi38 & ~n17367;
  assign n17369 = n62765 & ~n17368;
  assign n17370 = ~pi181 & n8009;
  assign n17371 = ~n17369 & ~n17370;
  assign n17372 = ~pi181 & ~n7357;
  assign n17373 = n8085 & ~n17372;
  assign n17374 = ~pi709 & ~n17373;
  assign n17375 = ~n17371 & n17374;
  assign n17376 = ~n17366 & ~n17375;
  assign n17377 = ~pi778 & n17376;
  assign n17378 = pi625 & ~n17376;
  assign n17379 = ~pi625 & n17363;
  assign n17380 = pi1153 & ~n17379;
  assign n17381 = ~n17378 & n17380;
  assign n17382 = ~pi625 & ~n17376;
  assign n17383 = pi625 & n17363;
  assign n17384 = ~pi1153 & ~n17383;
  assign n17385 = ~n17382 & n17384;
  assign n17386 = ~n17381 & ~n17385;
  assign n17387 = pi778 & ~n17386;
  assign n17388 = ~n17377 & ~n17387;
  assign n17389 = ~n62880 & ~n17388;
  assign n17390 = n62880 & ~n17363;
  assign n17391 = ~n62880 & n17388;
  assign n17392 = n62880 & n17363;
  assign n17393 = ~n17391 & ~n17392;
  assign n17394 = ~n17389 & ~n17390;
  assign n17395 = ~n62882 & ~n63332;
  assign n17396 = n62882 & n17363;
  assign n17397 = n62882 & ~n17363;
  assign n17398 = ~n62882 & n63332;
  assign n17399 = ~n17397 & ~n17398;
  assign n17400 = ~n17395 & ~n17396;
  assign n17401 = ~n8257 & ~n63333;
  assign n17402 = ~n8257 & n63333;
  assign n17403 = n8257 & n17363;
  assign n17404 = ~n17402 & ~n17403;
  assign n17405 = ~n17364 & ~n17401;
  assign n17406 = ~n8303 & ~n63334;
  assign n17407 = n8303 & n17363;
  assign n17408 = ~n17406 & ~n17407;
  assign n17409 = ~pi792 & n17408;
  assign n17410 = pi628 & ~n17408;
  assign n17411 = ~pi628 & n17363;
  assign n17412 = pi1156 & ~n17411;
  assign n17413 = ~n17410 & n17412;
  assign n17414 = ~pi628 & ~n17408;
  assign n17415 = pi628 & n17363;
  assign n17416 = ~pi1156 & ~n17415;
  assign n17417 = ~n17414 & n17416;
  assign n17418 = ~n17413 & ~n17417;
  assign n17419 = pi792 & ~n17418;
  assign n17420 = ~n17409 & ~n17419;
  assign n17421 = pi647 & n17420;
  assign n17422 = ~pi647 & n17363;
  assign n17423 = pi1157 & ~n17422;
  assign n17424 = pi647 & ~n17420;
  assign n17425 = ~pi647 & ~n17363;
  assign n17426 = ~n17421 & ~n17422;
  assign n17427 = ~n17424 & ~n17425;
  assign n17428 = pi1157 & n63335;
  assign n17429 = ~n17421 & n17423;
  assign n17430 = ~pi647 & n17420;
  assign n17431 = pi647 & n17363;
  assign n17432 = ~pi1157 & ~n17431;
  assign n17433 = ~n17430 & n17432;
  assign n17434 = ~pi647 & ~n17420;
  assign n17435 = pi647 & ~n17363;
  assign n17436 = ~n17434 & ~n17435;
  assign n17437 = ~pi1157 & n17436;
  assign n17438 = pi1157 & ~n63335;
  assign n17439 = ~n17437 & ~n17438;
  assign n17440 = ~n63336 & ~n17433;
  assign n17441 = pi787 & n63337;
  assign n17442 = ~pi787 & ~n17420;
  assign n17443 = pi787 & ~n63337;
  assign n17444 = ~pi787 & n17420;
  assign n17445 = ~n17443 & ~n17444;
  assign n17446 = ~n17441 & ~n17442;
  assign n17447 = ~pi644 & ~n63338;
  assign n17448 = pi715 & ~n17447;
  assign n17449 = ~n11558 & n17363;
  assign n17450 = pi181 & ~n62765;
  assign n17451 = pi754 & n7143;
  assign n17452 = pi181 & n7349;
  assign n17453 = ~n17451 & ~n17452;
  assign n17454 = pi39 & ~n17453;
  assign n17455 = ~pi181 & ~pi754;
  assign n17456 = n62802 & n17455;
  assign n17457 = pi181 & pi754;
  assign n17458 = pi754 & ~n62781;
  assign n17459 = pi181 & ~n7292;
  assign n17460 = ~n17458 & ~n17459;
  assign n17461 = ~pi39 & ~n17460;
  assign n17462 = ~n17457 & ~n17461;
  assign n17463 = ~n17456 & n17462;
  assign n17464 = ~n17454 & n17463;
  assign n17465 = ~pi38 & ~n17464;
  assign n17466 = ~pi754 & n7359;
  assign n17467 = pi38 & ~n17372;
  assign n17468 = ~n17466 & n17467;
  assign n17469 = ~n17465 & ~n17468;
  assign n17470 = n62765 & ~n17469;
  assign n17471 = ~n17450 & ~n17470;
  assign n17472 = ~n8135 & ~n17471;
  assign n17473 = n8135 & ~n17363;
  assign n17474 = ~n17472 & ~n17473;
  assign n17475 = ~pi785 & ~n17474;
  assign n17476 = ~n8136 & ~n17363;
  assign n17477 = pi609 & n17472;
  assign n17478 = ~n17476 & ~n17477;
  assign n17479 = pi1155 & ~n17478;
  assign n17480 = ~n8148 & ~n17363;
  assign n17481 = ~pi609 & n17472;
  assign n17482 = ~n17480 & ~n17481;
  assign n17483 = ~pi1155 & ~n17482;
  assign n17484 = ~n17479 & ~n17483;
  assign n17485 = pi785 & ~n17484;
  assign n17486 = ~n17475 & ~n17485;
  assign n17487 = ~pi781 & ~n17486;
  assign n17488 = pi618 & n17486;
  assign n17489 = ~pi618 & n17363;
  assign n17490 = pi1154 & ~n17489;
  assign n17491 = ~n17488 & n17490;
  assign n17492 = ~pi618 & n17486;
  assign n17493 = pi618 & n17363;
  assign n17494 = ~pi1154 & ~n17493;
  assign n17495 = ~n17492 & n17494;
  assign n17496 = ~n17491 & ~n17495;
  assign n17497 = pi781 & ~n17496;
  assign n17498 = ~n17487 & ~n17497;
  assign n17499 = ~pi619 & ~n17498;
  assign n17500 = pi619 & ~n17363;
  assign n17501 = ~pi1159 & ~n17500;
  assign n17502 = ~n17499 & n17501;
  assign n17503 = pi619 & ~n17498;
  assign n17504 = ~pi619 & ~n17363;
  assign n17505 = pi1159 & ~n17504;
  assign n17506 = ~n17503 & n17505;
  assign n17507 = pi619 & n17498;
  assign n17508 = ~pi619 & n17363;
  assign n17509 = pi1159 & ~n17508;
  assign n17510 = ~n17507 & n17509;
  assign n17511 = ~pi619 & n17498;
  assign n17512 = pi619 & n17363;
  assign n17513 = ~pi1159 & ~n17512;
  assign n17514 = ~n17511 & n17513;
  assign n17515 = ~n17510 & ~n17514;
  assign n17516 = ~n17502 & ~n17506;
  assign n17517 = pi789 & n63339;
  assign n17518 = ~pi789 & n17498;
  assign n17519 = ~pi789 & ~n17498;
  assign n17520 = pi789 & ~n63339;
  assign n17521 = ~n17519 & ~n17520;
  assign n17522 = ~n17517 & ~n17518;
  assign n17523 = ~n8595 & n63340;
  assign n17524 = n8685 & n17523;
  assign n17525 = n8376 & ~n17363;
  assign n17526 = n8595 & n17363;
  assign n17527 = ~n17523 & ~n17526;
  assign n17528 = ~n8334 & ~n17527;
  assign n17529 = n8334 & n17363;
  assign n17530 = ~n17528 & ~n17529;
  assign n17531 = ~n8376 & n17530;
  assign n17532 = ~n17525 & ~n17531;
  assign n17533 = ~n8376 & ~n17530;
  assign n17534 = n8376 & n17363;
  assign n17535 = ~n17533 & ~n17534;
  assign n17536 = ~n17449 & ~n17524;
  assign n17537 = pi644 & n63341;
  assign n17538 = ~pi644 & n17363;
  assign n17539 = ~pi715 & ~n17538;
  assign n17540 = ~n17537 & n17539;
  assign n17541 = pi1160 & ~n17540;
  assign n17542 = ~n17448 & n17541;
  assign n17543 = pi644 & ~n63338;
  assign n17544 = ~pi715 & ~n17543;
  assign n17545 = ~pi644 & n63341;
  assign n17546 = pi644 & n17363;
  assign n17547 = pi715 & ~n17546;
  assign n17548 = ~n17545 & n17547;
  assign n17549 = ~pi1160 & ~n17548;
  assign n17550 = ~n17544 & n17549;
  assign n17551 = ~n17542 & ~n17550;
  assign n17552 = pi790 & ~n17551;
  assign n17553 = ~n63052 & n17527;
  assign n17554 = ~pi629 & n17413;
  assign n17555 = pi629 & n17417;
  assign n17556 = ~n17554 & ~n17555;
  assign n17557 = ~n17553 & n17556;
  assign n17558 = pi792 & ~n17557;
  assign n17559 = ~pi626 & ~n63340;
  assign n17560 = pi626 & ~n17363;
  assign n17561 = n8301 & ~n17560;
  assign n17562 = ~n17559 & n17561;
  assign n17563 = n8525 & ~n63334;
  assign n17564 = pi626 & ~n63340;
  assign n17565 = ~pi626 & ~n17363;
  assign n17566 = n8300 & ~n17565;
  assign n17567 = ~n17564 & n17566;
  assign n17568 = ~n17563 & ~n17567;
  assign n17569 = ~n17562 & ~n17563;
  assign n17570 = ~n17567 & n17569;
  assign n17571 = ~n17562 & n17568;
  assign n17572 = pi788 & ~n63342;
  assign n17573 = pi709 & n17469;
  assign n17574 = ~pi181 & ~n62821;
  assign n17575 = pi181 & n7632;
  assign n17576 = pi754 & ~n17575;
  assign n17577 = ~n17574 & n17576;
  assign n17578 = pi181 & n7709;
  assign n17579 = ~pi181 & n62851;
  assign n17580 = ~pi754 & ~n17579;
  assign n17581 = ~n17578 & n17580;
  assign n17582 = pi39 & ~n17581;
  assign n17583 = ~n17577 & n17582;
  assign n17584 = pi181 & n7855;
  assign n17585 = ~pi181 & n7832;
  assign n17586 = pi754 & ~n17585;
  assign n17587 = ~n17584 & n17586;
  assign n17588 = ~pi181 & ~n7861;
  assign n17589 = pi181 & ~n7868;
  assign n17590 = ~pi754 & ~n17589;
  assign n17591 = ~n17588 & n17590;
  assign n17592 = ~pi39 & ~n17591;
  assign n17593 = pi181 & ~n7855;
  assign n17594 = ~pi181 & ~n7832;
  assign n17595 = pi754 & ~n17594;
  assign n17596 = pi754 & ~n17593;
  assign n17597 = ~n17594 & n17596;
  assign n17598 = ~n17593 & n17595;
  assign n17599 = ~pi181 & n7861;
  assign n17600 = pi181 & n7868;
  assign n17601 = ~pi754 & ~n17600;
  assign n17602 = ~n17599 & n17601;
  assign n17603 = ~n63343 & ~n17602;
  assign n17604 = ~pi39 & ~n17603;
  assign n17605 = ~n17587 & n17592;
  assign n17606 = ~pi38 & ~n63344;
  assign n17607 = ~n17583 & n17606;
  assign n17608 = ~pi754 & ~n7744;
  assign n17609 = n10350 & ~n17608;
  assign n17610 = ~pi181 & ~n17609;
  assign n17611 = ~n7565 & ~n17138;
  assign n17612 = pi181 & ~n17611;
  assign n17613 = n7356 & n17612;
  assign n17614 = pi38 & ~n17613;
  assign n17615 = ~n17610 & n17614;
  assign n17616 = ~pi709 & ~n17615;
  assign n17617 = ~n17607 & n17616;
  assign n17618 = n62765 & ~n17617;
  assign n17619 = ~n17573 & n17618;
  assign n17620 = ~n17450 & ~n17619;
  assign n17621 = ~pi625 & n17620;
  assign n17622 = pi625 & n17471;
  assign n17623 = ~pi1153 & ~n17622;
  assign n17624 = ~n17621 & n17623;
  assign n17625 = ~pi608 & ~n17381;
  assign n17626 = ~n17624 & n17625;
  assign n17627 = pi625 & n17620;
  assign n17628 = ~pi625 & n17471;
  assign n17629 = pi1153 & ~n17628;
  assign n17630 = ~n17627 & n17629;
  assign n17631 = pi608 & ~n17385;
  assign n17632 = ~n17630 & n17631;
  assign n17633 = ~n17626 & ~n17632;
  assign n17634 = pi778 & ~n17633;
  assign n17635 = ~pi778 & n17620;
  assign n17636 = ~n17634 & ~n17635;
  assign n17637 = ~pi609 & ~n17636;
  assign n17638 = pi609 & n17388;
  assign n17639 = ~pi1155 & ~n17638;
  assign n17640 = ~n17637 & n17639;
  assign n17641 = ~pi660 & ~n17479;
  assign n17642 = ~n17640 & n17641;
  assign n17643 = pi609 & ~n17636;
  assign n17644 = ~pi609 & n17388;
  assign n17645 = pi1155 & ~n17644;
  assign n17646 = ~n17643 & n17645;
  assign n17647 = pi660 & ~n17483;
  assign n17648 = ~n17646 & n17647;
  assign n17649 = ~n17642 & ~n17648;
  assign n17650 = pi785 & ~n17649;
  assign n17651 = ~pi785 & ~n17636;
  assign n17652 = ~n17650 & ~n17651;
  assign n17653 = ~pi781 & n17652;
  assign n17654 = ~pi618 & ~n17652;
  assign n17655 = pi618 & ~n63332;
  assign n17656 = ~pi1154 & ~n17655;
  assign n17657 = ~n17654 & n17656;
  assign n17658 = ~pi627 & ~n17491;
  assign n17659 = ~n17657 & n17658;
  assign n17660 = pi618 & ~n17652;
  assign n17661 = ~pi618 & ~n63332;
  assign n17662 = pi1154 & ~n17661;
  assign n17663 = ~n17660 & n17662;
  assign n17664 = pi627 & ~n17495;
  assign n17665 = ~n17663 & n17664;
  assign n17666 = pi781 & ~n17665;
  assign n17667 = ~n17659 & n17666;
  assign n17668 = ~n17659 & ~n17665;
  assign n17669 = pi781 & ~n17668;
  assign n17670 = ~pi781 & ~n17652;
  assign n17671 = ~n17669 & ~n17670;
  assign n17672 = ~n17653 & ~n17667;
  assign n17673 = ~n11434 & n63345;
  assign n17674 = ~n11431 & ~n63333;
  assign n17675 = ~n62884 & ~n63339;
  assign n17676 = ~n17674 & ~n17675;
  assign n17677 = pi789 & ~n17676;
  assign n17678 = n62894 & ~n17677;
  assign n17679 = ~pi619 & ~n63345;
  assign n17680 = pi619 & n63333;
  assign n17681 = ~pi1159 & ~n17680;
  assign n17682 = ~n17679 & n17681;
  assign n17683 = ~pi648 & ~n17510;
  assign n17684 = ~n17682 & n17683;
  assign n17685 = pi619 & ~n63345;
  assign n17686 = ~pi619 & n63333;
  assign n17687 = pi1159 & ~n17686;
  assign n17688 = ~n17685 & n17687;
  assign n17689 = pi648 & ~n17514;
  assign n17690 = ~n17688 & n17689;
  assign n17691 = pi789 & ~n17690;
  assign n17692 = pi789 & ~n17684;
  assign n17693 = ~n17690 & n17692;
  assign n17694 = ~n17684 & n17691;
  assign n17695 = ~pi789 & n63345;
  assign n17696 = n62894 & ~n17695;
  assign n17697 = ~n63346 & n17696;
  assign n17698 = ~n17673 & n17678;
  assign n17699 = ~n63030 & ~n63347;
  assign n17700 = ~n63030 & ~n17572;
  assign n17701 = ~n63347 & n17700;
  assign n17702 = ~n17572 & n17699;
  assign n17703 = ~n17558 & ~n63348;
  assign n17704 = ~n8651 & ~n17703;
  assign n17705 = ~n8413 & ~n17529;
  assign n17706 = ~n8413 & n17530;
  assign n17707 = ~n17528 & n17705;
  assign n17708 = n8373 & n63335;
  assign n17709 = ~pi630 & n63336;
  assign n17710 = n8374 & ~n17436;
  assign n17711 = pi630 & n17433;
  assign n17712 = ~n63350 & ~n63351;
  assign n17713 = ~n63349 & n17712;
  assign n17714 = pi787 & ~n17713;
  assign n17715 = ~pi644 & n17549;
  assign n17716 = pi644 & n17541;
  assign n17717 = n14029 & ~n17540;
  assign n17718 = pi790 & ~n63352;
  assign n17719 = pi790 & ~n17715;
  assign n17720 = ~n63352 & n17719;
  assign n17721 = ~n17715 & n17718;
  assign n17722 = ~n17714 & ~n63353;
  assign n17723 = ~n17704 & ~n17714;
  assign n17724 = ~n63353 & n17723;
  assign n17725 = ~n17704 & n17722;
  assign n17726 = ~n17552 & ~n63354;
  assign n17727 = n62455 & ~n17726;
  assign n17728 = ~pi181 & ~n62455;
  assign n17729 = ~pi832 & ~n17728;
  assign n17730 = ~n17727 & n17729;
  assign po338 = ~n17362 & ~n17730;
  assign n17732 = ~pi182 & ~n2923;
  assign n17733 = ~pi756 & n7316;
  assign n17734 = ~n17732 & ~n17733;
  assign n17735 = ~n8420 & ~n17734;
  assign n17736 = ~pi785 & ~n17735;
  assign n17737 = n8148 & n17733;
  assign n17738 = n17735 & ~n17737;
  assign n17739 = pi1155 & ~n17738;
  assign n17740 = ~pi1155 & ~n17732;
  assign n17741 = ~n17737 & n17740;
  assign n17742 = ~n17739 & ~n17741;
  assign n17743 = pi785 & ~n17742;
  assign n17744 = ~n17736 & ~n17743;
  assign n17745 = ~pi781 & ~n17744;
  assign n17746 = ~n8435 & n17744;
  assign n17747 = pi1154 & ~n17746;
  assign n17748 = ~n8438 & n17744;
  assign n17749 = ~pi1154 & ~n17748;
  assign n17750 = ~n17747 & ~n17749;
  assign n17751 = pi781 & ~n17750;
  assign n17752 = ~n17745 & ~n17751;
  assign n17753 = ~pi789 & ~n17752;
  assign n17754 = ~n12612 & n17752;
  assign n17755 = pi1159 & ~n17754;
  assign n17756 = ~n12615 & n17752;
  assign n17757 = ~pi1159 & ~n17756;
  assign n17758 = ~n17755 & ~n17757;
  assign n17759 = pi789 & ~n17758;
  assign n17760 = ~n17753 & ~n17759;
  assign n17761 = ~n15298 & n17752;
  assign n17762 = ~n8595 & n63355;
  assign n17763 = n8595 & n17732;
  assign n17764 = ~n8595 & ~n63355;
  assign n17765 = n8595 & ~n17732;
  assign n17766 = ~n17764 & ~n17765;
  assign n17767 = ~n17762 & ~n17763;
  assign n17768 = ~n8334 & n63356;
  assign n17769 = n8334 & n17732;
  assign n17770 = ~n8413 & ~n17769;
  assign n17771 = ~n17768 & ~n17769;
  assign n17772 = ~n8413 & n17771;
  assign n17773 = ~n17768 & n17770;
  assign n17774 = ~pi734 & n7564;
  assign n17775 = ~n17732 & ~n17774;
  assign n17776 = ~pi778 & ~n17775;
  assign n17777 = ~pi625 & n17774;
  assign n17778 = ~n17775 & ~n17777;
  assign n17779 = pi1153 & ~n17778;
  assign n17780 = ~pi1153 & ~n17732;
  assign n17781 = ~n17777 & n17780;
  assign n17782 = pi778 & ~n17781;
  assign n17783 = ~n17779 & n17782;
  assign n17784 = ~n17776 & ~n17783;
  assign n17785 = ~n8490 & ~n17784;
  assign n17786 = ~n8492 & n17785;
  assign n17787 = ~n8494 & n17786;
  assign n17788 = ~n8496 & n17787;
  assign n17789 = ~n8508 & n17788;
  assign n17790 = pi647 & ~n17789;
  assign n17791 = ~pi647 & ~n17732;
  assign n17792 = ~n17790 & ~n17791;
  assign n17793 = n8373 & ~n17792;
  assign n17794 = ~pi647 & n17789;
  assign n17795 = pi647 & n17732;
  assign n17796 = ~pi1157 & ~n17795;
  assign n17797 = ~n17794 & n17796;
  assign n17798 = pi630 & n17797;
  assign n17799 = ~n17793 & ~n17798;
  assign n17800 = ~n63357 & n17799;
  assign n17801 = pi787 & ~n17800;
  assign n17802 = ~pi626 & ~n63355;
  assign n17803 = pi626 & ~n17732;
  assign n17804 = n8301 & ~n17803;
  assign n17805 = ~n17802 & n17804;
  assign n17806 = n8525 & n17787;
  assign n17807 = pi626 & ~n63355;
  assign n17808 = ~pi626 & ~n17732;
  assign n17809 = n8300 & ~n17808;
  assign n17810 = ~n17807 & n17809;
  assign n17811 = ~n17806 & ~n17810;
  assign n17812 = ~n17805 & ~n17806;
  assign n17813 = ~n17810 & n17812;
  assign n17814 = ~n17805 & n17811;
  assign n17815 = pi788 & ~n63358;
  assign n17816 = n13460 & n17752;
  assign n17817 = n11303 & n17786;
  assign n17818 = pi648 & ~n17817;
  assign n17819 = ~n17816 & n17818;
  assign n17820 = n13462 & n17752;
  assign n17821 = n11304 & n17786;
  assign n17822 = ~pi648 & ~n17821;
  assign n17823 = ~n17820 & n17822;
  assign n17824 = pi789 & ~n17823;
  assign n17825 = ~n17819 & n17824;
  assign n17826 = ~n7187 & ~n17775;
  assign n17827 = pi625 & n17826;
  assign n17828 = n17734 & ~n17826;
  assign n17829 = ~n17827 & ~n17828;
  assign n17830 = n17780 & ~n17829;
  assign n17831 = ~pi608 & ~n17779;
  assign n17832 = ~n17830 & n17831;
  assign n17833 = pi1153 & n17734;
  assign n17834 = ~n17827 & n17833;
  assign n17835 = pi608 & ~n17781;
  assign n17836 = ~n17834 & n17835;
  assign n17837 = ~n17832 & ~n17836;
  assign n17838 = pi778 & ~n17837;
  assign n17839 = ~pi778 & ~n17828;
  assign n17840 = ~n17838 & ~n17839;
  assign n17841 = ~pi609 & ~n17840;
  assign n17842 = pi609 & ~n17784;
  assign n17843 = ~pi1155 & ~n17842;
  assign n17844 = ~n17841 & n17843;
  assign n17845 = ~pi660 & ~n17739;
  assign n17846 = ~n17844 & n17845;
  assign n17847 = pi609 & ~n17840;
  assign n17848 = ~pi609 & ~n17784;
  assign n17849 = pi1155 & ~n17848;
  assign n17850 = ~n17847 & n17849;
  assign n17851 = pi660 & ~n17741;
  assign n17852 = ~n17850 & n17851;
  assign n17853 = ~n17846 & ~n17852;
  assign n17854 = pi785 & ~n17853;
  assign n17855 = ~pi785 & ~n17840;
  assign n17856 = ~n17854 & ~n17855;
  assign n17857 = pi618 & ~n17856;
  assign n17858 = ~pi618 & n17785;
  assign n17859 = pi1154 & ~n17858;
  assign n17860 = ~n17857 & n17859;
  assign n17861 = pi627 & ~n17749;
  assign n17862 = ~n17860 & n17861;
  assign n17863 = ~pi618 & ~n17856;
  assign n17864 = pi618 & n17785;
  assign n17865 = ~pi1154 & ~n17864;
  assign n17866 = ~n17863 & n17865;
  assign n17867 = ~pi627 & ~n17747;
  assign n17868 = ~n17866 & n17867;
  assign n17869 = pi781 & ~n17868;
  assign n17870 = ~n17862 & n17869;
  assign n17871 = ~pi781 & n17856;
  assign n17872 = ~n11434 & ~n17871;
  assign n17873 = ~n17870 & n17872;
  assign n17874 = ~n17825 & ~n17873;
  assign n17875 = ~n17862 & ~n17868;
  assign n17876 = pi781 & ~n17875;
  assign n17877 = ~pi781 & ~n17856;
  assign n17878 = ~n17876 & ~n17877;
  assign n17879 = ~pi619 & ~n17878;
  assign n17880 = pi619 & n17786;
  assign n17881 = ~pi1159 & ~n17880;
  assign n17882 = ~n17879 & n17881;
  assign n17883 = ~pi648 & ~n17755;
  assign n17884 = ~n17882 & n17883;
  assign n17885 = pi619 & ~n17878;
  assign n17886 = ~pi619 & n17786;
  assign n17887 = pi1159 & ~n17886;
  assign n17888 = ~n17885 & n17887;
  assign n17889 = pi648 & ~n17757;
  assign n17890 = ~n17888 & n17889;
  assign n17891 = pi789 & ~n17890;
  assign n17892 = pi789 & ~n17884;
  assign n17893 = ~n17890 & n17892;
  assign n17894 = ~n17884 & n17891;
  assign n17895 = ~pi789 & n17878;
  assign n17896 = n62894 & ~n17895;
  assign n17897 = ~n63359 & n17896;
  assign n17898 = n62894 & ~n17874;
  assign n17899 = ~n17815 & ~n63360;
  assign n17900 = ~n63030 & ~n17899;
  assign n17901 = n8498 & n63356;
  assign n17902 = n8615 & n17788;
  assign n17903 = pi629 & ~n17902;
  assign n17904 = ~n17901 & n17903;
  assign n17905 = n8499 & n63356;
  assign n17906 = n8606 & n17788;
  assign n17907 = ~pi629 & ~n17906;
  assign n17908 = ~n17905 & n17907;
  assign n17909 = pi792 & ~n17908;
  assign n17910 = pi792 & ~n17904;
  assign n17911 = ~n17908 & n17910;
  assign n17912 = ~n17905 & ~n17906;
  assign n17913 = ~pi629 & ~n17912;
  assign n17914 = ~n17901 & ~n17902;
  assign n17915 = pi629 & ~n17914;
  assign n17916 = ~n17913 & ~n17915;
  assign n17917 = pi792 & ~n17916;
  assign n17918 = ~n17904 & n17909;
  assign n17919 = ~n8651 & ~n63361;
  assign n17920 = ~n17900 & n17919;
  assign n17921 = ~n17801 & ~n17920;
  assign n17922 = pi644 & n17921;
  assign n17923 = ~pi787 & ~n17789;
  assign n17924 = pi1157 & ~n17792;
  assign n17925 = ~n17797 & ~n17924;
  assign n17926 = pi787 & ~n17925;
  assign n17927 = ~n17923 & ~n17926;
  assign n17928 = ~pi644 & n17927;
  assign n17929 = pi715 & ~n17928;
  assign n17930 = ~n17922 & n17929;
  assign n17931 = ~n8685 & n17732;
  assign n17932 = ~n8376 & n17768;
  assign n17933 = ~n8376 & ~n17771;
  assign n17934 = n8376 & n17732;
  assign n17935 = ~n17933 & ~n17934;
  assign n17936 = ~n17931 & ~n17932;
  assign n17937 = pi644 & ~n63362;
  assign n17938 = ~pi644 & n17732;
  assign n17939 = ~pi715 & ~n17938;
  assign n17940 = ~n17937 & n17939;
  assign n17941 = pi1160 & ~n17940;
  assign n17942 = ~n17930 & n17941;
  assign n17943 = ~pi644 & n17921;
  assign n17944 = pi644 & n17927;
  assign n17945 = ~pi715 & ~n17944;
  assign n17946 = ~n17943 & n17945;
  assign n17947 = ~pi644 & ~n63362;
  assign n17948 = pi644 & n17732;
  assign n17949 = pi715 & ~n17948;
  assign n17950 = ~n17947 & n17949;
  assign n17951 = ~pi1160 & ~n17950;
  assign n17952 = ~n17946 & n17951;
  assign n17953 = ~n17942 & ~n17952;
  assign n17954 = pi790 & ~n17953;
  assign n17955 = ~pi790 & n17921;
  assign n17956 = pi832 & ~n17955;
  assign n17957 = ~n17954 & n17956;
  assign n17958 = ~pi182 & ~n8098;
  assign n17959 = n8257 & ~n17958;
  assign n17960 = ~pi734 & n62765;
  assign n17961 = n17958 & ~n17960;
  assign n17962 = pi182 & n62874;
  assign n17963 = ~pi38 & ~n17962;
  assign n17964 = n62765 & ~n17963;
  assign n17965 = ~pi182 & n8009;
  assign n17966 = ~n17964 & ~n17965;
  assign n17967 = ~pi182 & ~n7357;
  assign n17968 = n8085 & ~n17967;
  assign n17969 = ~pi734 & ~n17968;
  assign n17970 = ~n17966 & n17969;
  assign n17971 = ~n17961 & ~n17970;
  assign n17972 = ~pi778 & n17971;
  assign n17973 = pi625 & ~n17971;
  assign n17974 = ~pi625 & n17958;
  assign n17975 = pi1153 & ~n17974;
  assign n17976 = ~n17973 & n17975;
  assign n17977 = ~pi625 & ~n17971;
  assign n17978 = pi625 & n17958;
  assign n17979 = ~pi1153 & ~n17978;
  assign n17980 = ~n17977 & n17979;
  assign n17981 = ~n17976 & ~n17980;
  assign n17982 = pi778 & ~n17981;
  assign n17983 = ~n17972 & ~n17982;
  assign n17984 = ~n62880 & ~n17983;
  assign n17985 = n62880 & ~n17958;
  assign n17986 = ~n62880 & n17983;
  assign n17987 = n62880 & n17958;
  assign n17988 = ~n17986 & ~n17987;
  assign n17989 = ~n17984 & ~n17985;
  assign n17990 = ~n62882 & ~n63363;
  assign n17991 = n62882 & n17958;
  assign n17992 = n62882 & ~n17958;
  assign n17993 = ~n62882 & n63363;
  assign n17994 = ~n17992 & ~n17993;
  assign n17995 = ~n17990 & ~n17991;
  assign n17996 = ~n8257 & ~n63364;
  assign n17997 = ~n8257 & n63364;
  assign n17998 = n8257 & n17958;
  assign n17999 = ~n17997 & ~n17998;
  assign n18000 = ~n17959 & ~n17996;
  assign n18001 = ~n8303 & ~n63365;
  assign n18002 = n8303 & n17958;
  assign n18003 = ~n18001 & ~n18002;
  assign n18004 = ~pi792 & n18003;
  assign n18005 = pi628 & ~n18003;
  assign n18006 = ~pi628 & n17958;
  assign n18007 = pi1156 & ~n18006;
  assign n18008 = ~n18005 & n18007;
  assign n18009 = ~pi628 & ~n18003;
  assign n18010 = pi628 & n17958;
  assign n18011 = ~pi1156 & ~n18010;
  assign n18012 = ~n18009 & n18011;
  assign n18013 = ~n18008 & ~n18012;
  assign n18014 = pi792 & ~n18013;
  assign n18015 = ~n18004 & ~n18014;
  assign n18016 = pi647 & n18015;
  assign n18017 = ~pi647 & n17958;
  assign n18018 = pi1157 & ~n18017;
  assign n18019 = pi647 & ~n18015;
  assign n18020 = ~pi647 & ~n17958;
  assign n18021 = ~n18016 & ~n18017;
  assign n18022 = ~n18019 & ~n18020;
  assign n18023 = pi1157 & n63366;
  assign n18024 = ~n18016 & n18018;
  assign n18025 = ~pi647 & n18015;
  assign n18026 = pi647 & n17958;
  assign n18027 = ~pi1157 & ~n18026;
  assign n18028 = ~n18025 & n18027;
  assign n18029 = ~pi647 & ~n18015;
  assign n18030 = pi647 & ~n17958;
  assign n18031 = ~n18029 & ~n18030;
  assign n18032 = ~pi1157 & n18031;
  assign n18033 = pi1157 & ~n63366;
  assign n18034 = ~n18032 & ~n18033;
  assign n18035 = ~n63367 & ~n18028;
  assign n18036 = pi787 & n63368;
  assign n18037 = ~pi787 & ~n18015;
  assign n18038 = pi787 & ~n63368;
  assign n18039 = ~pi787 & n18015;
  assign n18040 = ~n18038 & ~n18039;
  assign n18041 = ~n18036 & ~n18037;
  assign n18042 = ~pi644 & ~n63369;
  assign n18043 = pi715 & ~n18042;
  assign n18044 = ~n11558 & n17958;
  assign n18045 = pi182 & ~n62765;
  assign n18046 = ~pi756 & n7359;
  assign n18047 = ~n17967 & ~n18046;
  assign n18048 = pi38 & ~n18047;
  assign n18049 = ~pi182 & n62802;
  assign n18050 = pi182 & ~n7351;
  assign n18051 = ~pi756 & ~n18050;
  assign n18052 = ~n18049 & n18051;
  assign n18053 = ~pi182 & pi756;
  assign n18054 = ~n62792 & n18053;
  assign n18055 = pi756 & ~n62792;
  assign n18056 = ~pi756 & ~n18049;
  assign n18057 = ~n18055 & ~n18056;
  assign n18058 = ~pi182 & ~n18057;
  assign n18059 = n7351 & n18056;
  assign n18060 = ~n18058 & ~n18059;
  assign n18061 = ~n18052 & ~n18054;
  assign n18062 = ~pi38 & ~n63370;
  assign n18063 = ~n18048 & ~n18062;
  assign n18064 = n62765 & n18063;
  assign n18065 = ~n18045 & ~n18064;
  assign n18066 = ~n8135 & ~n18065;
  assign n18067 = n8135 & ~n17958;
  assign n18068 = ~n18066 & ~n18067;
  assign n18069 = ~pi785 & ~n18068;
  assign n18070 = ~n8136 & ~n17958;
  assign n18071 = pi609 & n18066;
  assign n18072 = ~n18070 & ~n18071;
  assign n18073 = pi1155 & ~n18072;
  assign n18074 = ~n8148 & ~n17958;
  assign n18075 = ~pi609 & n18066;
  assign n18076 = ~n18074 & ~n18075;
  assign n18077 = ~pi1155 & ~n18076;
  assign n18078 = ~n18073 & ~n18077;
  assign n18079 = pi785 & ~n18078;
  assign n18080 = ~n18069 & ~n18079;
  assign n18081 = ~pi781 & ~n18080;
  assign n18082 = pi618 & n18080;
  assign n18083 = ~pi618 & n17958;
  assign n18084 = pi1154 & ~n18083;
  assign n18085 = ~n18082 & n18084;
  assign n18086 = ~pi618 & n18080;
  assign n18087 = pi618 & n17958;
  assign n18088 = ~pi1154 & ~n18087;
  assign n18089 = ~n18086 & n18088;
  assign n18090 = ~n18085 & ~n18089;
  assign n18091 = pi781 & ~n18090;
  assign n18092 = ~n18081 & ~n18091;
  assign n18093 = ~pi619 & ~n18092;
  assign n18094 = pi619 & ~n17958;
  assign n18095 = ~pi1159 & ~n18094;
  assign n18096 = ~n18093 & n18095;
  assign n18097 = pi619 & ~n18092;
  assign n18098 = ~pi619 & ~n17958;
  assign n18099 = pi1159 & ~n18098;
  assign n18100 = ~n18097 & n18099;
  assign n18101 = pi619 & n18092;
  assign n18102 = ~pi619 & n17958;
  assign n18103 = pi1159 & ~n18102;
  assign n18104 = ~n18101 & n18103;
  assign n18105 = ~pi619 & n18092;
  assign n18106 = pi619 & n17958;
  assign n18107 = ~pi1159 & ~n18106;
  assign n18108 = ~n18105 & n18107;
  assign n18109 = ~n18104 & ~n18108;
  assign n18110 = ~n18096 & ~n18100;
  assign n18111 = pi789 & n63371;
  assign n18112 = ~pi789 & n18092;
  assign n18113 = ~pi789 & ~n18092;
  assign n18114 = pi789 & ~n63371;
  assign n18115 = ~n18113 & ~n18114;
  assign n18116 = ~n18111 & ~n18112;
  assign n18117 = ~n8595 & n63372;
  assign n18118 = n8685 & n18117;
  assign n18119 = n8376 & ~n17958;
  assign n18120 = n8595 & n17958;
  assign n18121 = ~n18117 & ~n18120;
  assign n18122 = ~n8334 & ~n18121;
  assign n18123 = n8334 & n17958;
  assign n18124 = ~n18122 & ~n18123;
  assign n18125 = ~n8376 & n18124;
  assign n18126 = ~n18119 & ~n18125;
  assign n18127 = ~n8376 & ~n18124;
  assign n18128 = n8376 & n17958;
  assign n18129 = ~n18127 & ~n18128;
  assign n18130 = ~n18044 & ~n18118;
  assign n18131 = pi644 & n63373;
  assign n18132 = ~pi644 & n17958;
  assign n18133 = ~pi715 & ~n18132;
  assign n18134 = ~n18131 & n18133;
  assign n18135 = pi1160 & ~n18134;
  assign n18136 = ~n18043 & n18135;
  assign n18137 = pi644 & ~n63369;
  assign n18138 = ~pi715 & ~n18137;
  assign n18139 = ~pi644 & n63373;
  assign n18140 = pi644 & n17958;
  assign n18141 = pi715 & ~n18140;
  assign n18142 = ~n18139 & n18141;
  assign n18143 = ~pi1160 & ~n18142;
  assign n18144 = ~n18138 & n18143;
  assign n18145 = ~n18136 & ~n18144;
  assign n18146 = pi790 & ~n18145;
  assign n18147 = ~n63052 & n18121;
  assign n18148 = ~pi629 & n18008;
  assign n18149 = pi629 & n18012;
  assign n18150 = ~n18148 & ~n18149;
  assign n18151 = ~n18147 & n18150;
  assign n18152 = pi792 & ~n18151;
  assign n18153 = pi734 & ~n18063;
  assign n18154 = ~pi182 & ~n62821;
  assign n18155 = pi182 & n7632;
  assign n18156 = pi756 & ~n18155;
  assign n18157 = ~n18154 & n18156;
  assign n18158 = pi182 & n7709;
  assign n18159 = ~pi182 & n62851;
  assign n18160 = ~pi756 & ~n18159;
  assign n18161 = ~n18158 & n18160;
  assign n18162 = pi39 & ~n18161;
  assign n18163 = ~n18157 & n18162;
  assign n18164 = pi182 & n7855;
  assign n18165 = ~pi182 & n7832;
  assign n18166 = pi756 & ~n18165;
  assign n18167 = ~n18164 & n18166;
  assign n18168 = ~pi182 & ~n7861;
  assign n18169 = pi182 & ~n7868;
  assign n18170 = ~pi756 & ~n18169;
  assign n18171 = ~n18168 & n18170;
  assign n18172 = ~pi39 & ~n18171;
  assign n18173 = pi182 & ~n7855;
  assign n18174 = ~pi182 & ~n7832;
  assign n18175 = pi756 & ~n18174;
  assign n18176 = pi756 & ~n18173;
  assign n18177 = ~n18174 & n18176;
  assign n18178 = ~n18173 & n18175;
  assign n18179 = ~pi182 & n7861;
  assign n18180 = pi182 & n7868;
  assign n18181 = ~pi756 & ~n18180;
  assign n18182 = ~n18179 & n18181;
  assign n18183 = ~n63374 & ~n18182;
  assign n18184 = ~pi39 & ~n18183;
  assign n18185 = ~n18167 & n18172;
  assign n18186 = ~pi38 & ~n63375;
  assign n18187 = ~n18163 & n18186;
  assign n18188 = ~pi756 & ~n7744;
  assign n18189 = n10350 & ~n18188;
  assign n18190 = ~pi182 & ~n18189;
  assign n18191 = ~n7565 & ~n17733;
  assign n18192 = pi182 & ~n18191;
  assign n18193 = n7356 & n18192;
  assign n18194 = pi38 & ~n18193;
  assign n18195 = ~n18190 & n18194;
  assign n18196 = ~pi734 & ~n18195;
  assign n18197 = ~n18187 & n18196;
  assign n18198 = n62765 & ~n18197;
  assign n18199 = ~n18153 & n18198;
  assign n18200 = ~n18045 & ~n18199;
  assign n18201 = ~pi625 & n18200;
  assign n18202 = pi625 & n18065;
  assign n18203 = ~pi1153 & ~n18202;
  assign n18204 = ~n18201 & n18203;
  assign n18205 = ~pi608 & ~n17976;
  assign n18206 = ~n18204 & n18205;
  assign n18207 = pi625 & n18200;
  assign n18208 = ~pi625 & n18065;
  assign n18209 = pi1153 & ~n18208;
  assign n18210 = ~n18207 & n18209;
  assign n18211 = pi608 & ~n17980;
  assign n18212 = ~n18210 & n18211;
  assign n18213 = ~n18206 & ~n18212;
  assign n18214 = pi778 & ~n18213;
  assign n18215 = ~pi778 & n18200;
  assign n18216 = ~n18214 & ~n18215;
  assign n18217 = ~pi609 & ~n18216;
  assign n18218 = pi609 & n17983;
  assign n18219 = ~pi1155 & ~n18218;
  assign n18220 = ~n18217 & n18219;
  assign n18221 = ~pi660 & ~n18073;
  assign n18222 = ~n18220 & n18221;
  assign n18223 = pi609 & ~n18216;
  assign n18224 = ~pi609 & n17983;
  assign n18225 = pi1155 & ~n18224;
  assign n18226 = ~n18223 & n18225;
  assign n18227 = pi660 & ~n18077;
  assign n18228 = ~n18226 & n18227;
  assign n18229 = ~n18222 & ~n18228;
  assign n18230 = pi785 & ~n18229;
  assign n18231 = ~pi785 & ~n18216;
  assign n18232 = ~n18230 & ~n18231;
  assign n18233 = pi618 & ~n18232;
  assign n18234 = ~pi618 & ~n63363;
  assign n18235 = pi1154 & ~n18234;
  assign n18236 = ~n18233 & n18235;
  assign n18237 = pi627 & ~n18089;
  assign n18238 = ~n18236 & n18237;
  assign n18239 = ~pi618 & ~n18232;
  assign n18240 = pi618 & ~n63363;
  assign n18241 = ~pi1154 & ~n18240;
  assign n18242 = ~n18239 & n18241;
  assign n18243 = ~pi627 & ~n18085;
  assign n18244 = ~n18242 & n18243;
  assign n18245 = pi781 & ~n18244;
  assign n18246 = ~n18238 & n18245;
  assign n18247 = ~n11431 & ~n63364;
  assign n18248 = ~n62884 & ~n63371;
  assign n18249 = ~n18247 & ~n18248;
  assign n18250 = pi789 & ~n18249;
  assign n18251 = ~pi781 & n18232;
  assign n18252 = ~n18250 & ~n18251;
  assign n18253 = ~n18246 & n18252;
  assign n18254 = n11434 & n18249;
  assign n18255 = ~n18253 & ~n18254;
  assign n18256 = ~n18238 & ~n18244;
  assign n18257 = pi781 & ~n18256;
  assign n18258 = ~pi781 & ~n18232;
  assign n18259 = ~n18257 & ~n18258;
  assign n18260 = ~pi619 & ~n18259;
  assign n18261 = pi619 & n63364;
  assign n18262 = ~pi1159 & ~n18261;
  assign n18263 = ~n18260 & n18262;
  assign n18264 = ~pi648 & ~n18104;
  assign n18265 = ~n18263 & n18264;
  assign n18266 = pi619 & ~n18259;
  assign n18267 = ~pi619 & n63364;
  assign n18268 = pi1159 & ~n18267;
  assign n18269 = ~n18266 & n18268;
  assign n18270 = pi648 & ~n18108;
  assign n18271 = ~n18269 & n18270;
  assign n18272 = pi789 & ~n18271;
  assign n18273 = pi789 & ~n18265;
  assign n18274 = ~n18271 & n18273;
  assign n18275 = ~n18265 & n18272;
  assign n18276 = ~pi789 & n18259;
  assign n18277 = n62894 & ~n18276;
  assign n18278 = ~n63376 & n18277;
  assign n18279 = n62894 & ~n18255;
  assign n18280 = ~pi626 & ~n63372;
  assign n18281 = pi626 & ~n17958;
  assign n18282 = n8301 & ~n18281;
  assign n18283 = ~n18280 & n18282;
  assign n18284 = n8525 & ~n63365;
  assign n18285 = pi626 & ~n63372;
  assign n18286 = ~pi626 & ~n17958;
  assign n18287 = n8300 & ~n18286;
  assign n18288 = ~n18285 & n18287;
  assign n18289 = ~n18284 & ~n18288;
  assign n18290 = ~n18283 & ~n18284;
  assign n18291 = ~n18288 & n18290;
  assign n18292 = ~n18283 & n18289;
  assign n18293 = pi788 & ~n63378;
  assign n18294 = ~n63030 & ~n18293;
  assign n18295 = ~n63377 & n18294;
  assign n18296 = ~n18152 & ~n18295;
  assign n18297 = ~n8651 & ~n18296;
  assign n18298 = ~n8413 & ~n18123;
  assign n18299 = ~n8413 & n18124;
  assign n18300 = ~n18122 & n18298;
  assign n18301 = n8373 & n63366;
  assign n18302 = ~pi630 & n63367;
  assign n18303 = n8374 & ~n18031;
  assign n18304 = pi630 & n18028;
  assign n18305 = ~n63380 & ~n63381;
  assign n18306 = ~n63379 & n18305;
  assign n18307 = pi787 & ~n18306;
  assign n18308 = ~pi644 & n18143;
  assign n18309 = pi644 & n18135;
  assign n18310 = n14029 & ~n18134;
  assign n18311 = pi790 & ~n63382;
  assign n18312 = pi790 & ~n18308;
  assign n18313 = ~n63382 & n18312;
  assign n18314 = ~n18308 & n18311;
  assign n18315 = ~n18307 & ~n63383;
  assign n18316 = ~n18297 & ~n18307;
  assign n18317 = ~n63383 & n18316;
  assign n18318 = ~n18297 & n18315;
  assign n18319 = ~n18146 & ~n63384;
  assign n18320 = n62455 & ~n18319;
  assign n18321 = ~pi182 & ~n62455;
  assign n18322 = ~pi832 & ~n18321;
  assign n18323 = ~n18320 & n18322;
  assign po339 = ~n17957 & ~n18323;
  assign n18325 = ~pi183 & ~n2923;
  assign n18326 = ~pi755 & n7316;
  assign n18327 = ~n18325 & ~n18326;
  assign n18328 = ~n8420 & ~n18327;
  assign n18329 = ~pi785 & ~n18328;
  assign n18330 = n8148 & n18326;
  assign n18331 = n18328 & ~n18330;
  assign n18332 = pi1155 & ~n18331;
  assign n18333 = ~pi1155 & ~n18325;
  assign n18334 = ~n18330 & n18333;
  assign n18335 = ~n18332 & ~n18334;
  assign n18336 = pi785 & ~n18335;
  assign n18337 = ~n18329 & ~n18336;
  assign n18338 = ~pi781 & ~n18337;
  assign n18339 = ~n8435 & n18337;
  assign n18340 = pi1154 & ~n18339;
  assign n18341 = ~n8438 & n18337;
  assign n18342 = ~pi1154 & ~n18341;
  assign n18343 = ~n18340 & ~n18342;
  assign n18344 = pi781 & ~n18343;
  assign n18345 = ~n18338 & ~n18344;
  assign n18346 = ~pi789 & ~n18345;
  assign n18347 = ~n12612 & n18345;
  assign n18348 = pi1159 & ~n18347;
  assign n18349 = ~n12615 & n18345;
  assign n18350 = ~pi1159 & ~n18349;
  assign n18351 = ~n18348 & ~n18350;
  assign n18352 = pi789 & ~n18351;
  assign n18353 = ~n18346 & ~n18352;
  assign n18354 = ~n15298 & n18345;
  assign n18355 = ~n8595 & n63385;
  assign n18356 = n8595 & n18325;
  assign n18357 = ~n8595 & ~n63385;
  assign n18358 = n8595 & ~n18325;
  assign n18359 = ~n18357 & ~n18358;
  assign n18360 = ~n18355 & ~n18356;
  assign n18361 = ~n8334 & n63386;
  assign n18362 = n8334 & n18325;
  assign n18363 = ~n8413 & ~n18362;
  assign n18364 = ~n18361 & ~n18362;
  assign n18365 = ~n8413 & n18364;
  assign n18366 = ~n18361 & n18363;
  assign n18367 = ~pi725 & n7564;
  assign n18368 = ~n18325 & ~n18367;
  assign n18369 = ~pi778 & ~n18368;
  assign n18370 = ~pi625 & n18367;
  assign n18371 = ~n18368 & ~n18370;
  assign n18372 = pi1153 & ~n18371;
  assign n18373 = ~pi1153 & ~n18325;
  assign n18374 = ~n18370 & n18373;
  assign n18375 = pi778 & ~n18374;
  assign n18376 = ~n18372 & n18375;
  assign n18377 = ~n18369 & ~n18376;
  assign n18378 = ~n8490 & ~n18377;
  assign n18379 = ~n8492 & n18378;
  assign n18380 = ~n8494 & n18379;
  assign n18381 = ~n8496 & n18380;
  assign n18382 = ~n8508 & n18381;
  assign n18383 = pi647 & ~n18382;
  assign n18384 = ~pi647 & ~n18325;
  assign n18385 = ~n18383 & ~n18384;
  assign n18386 = n8373 & ~n18385;
  assign n18387 = ~pi647 & n18382;
  assign n18388 = pi647 & n18325;
  assign n18389 = ~pi1157 & ~n18388;
  assign n18390 = ~n18387 & n18389;
  assign n18391 = pi630 & n18390;
  assign n18392 = ~n18386 & ~n18391;
  assign n18393 = ~n63387 & n18392;
  assign n18394 = pi787 & ~n18393;
  assign n18395 = ~pi626 & ~n63385;
  assign n18396 = pi626 & ~n18325;
  assign n18397 = n8301 & ~n18396;
  assign n18398 = ~n18395 & n18397;
  assign n18399 = n8525 & n18380;
  assign n18400 = pi626 & ~n63385;
  assign n18401 = ~pi626 & ~n18325;
  assign n18402 = n8300 & ~n18401;
  assign n18403 = ~n18400 & n18402;
  assign n18404 = ~n18399 & ~n18403;
  assign n18405 = ~n18398 & ~n18399;
  assign n18406 = ~n18403 & n18405;
  assign n18407 = ~n18398 & n18404;
  assign n18408 = pi788 & ~n63388;
  assign n18409 = n13460 & n18345;
  assign n18410 = n11303 & n18379;
  assign n18411 = pi648 & ~n18410;
  assign n18412 = ~n18409 & n18411;
  assign n18413 = n13462 & n18345;
  assign n18414 = n11304 & n18379;
  assign n18415 = ~pi648 & ~n18414;
  assign n18416 = ~n18413 & n18415;
  assign n18417 = pi789 & ~n18416;
  assign n18418 = ~n18412 & n18417;
  assign n18419 = ~n7187 & ~n18368;
  assign n18420 = pi625 & n18419;
  assign n18421 = n18327 & ~n18419;
  assign n18422 = ~n18420 & ~n18421;
  assign n18423 = n18373 & ~n18422;
  assign n18424 = ~pi608 & ~n18372;
  assign n18425 = ~n18423 & n18424;
  assign n18426 = pi1153 & n18327;
  assign n18427 = ~n18420 & n18426;
  assign n18428 = pi608 & ~n18374;
  assign n18429 = ~n18427 & n18428;
  assign n18430 = ~n18425 & ~n18429;
  assign n18431 = pi778 & ~n18430;
  assign n18432 = ~pi778 & ~n18421;
  assign n18433 = ~n18431 & ~n18432;
  assign n18434 = ~pi609 & ~n18433;
  assign n18435 = pi609 & ~n18377;
  assign n18436 = ~pi1155 & ~n18435;
  assign n18437 = ~n18434 & n18436;
  assign n18438 = ~pi660 & ~n18332;
  assign n18439 = ~n18437 & n18438;
  assign n18440 = pi609 & ~n18433;
  assign n18441 = ~pi609 & ~n18377;
  assign n18442 = pi1155 & ~n18441;
  assign n18443 = ~n18440 & n18442;
  assign n18444 = pi660 & ~n18334;
  assign n18445 = ~n18443 & n18444;
  assign n18446 = ~n18439 & ~n18445;
  assign n18447 = pi785 & ~n18446;
  assign n18448 = ~pi785 & ~n18433;
  assign n18449 = ~n18447 & ~n18448;
  assign n18450 = pi618 & ~n18449;
  assign n18451 = ~pi618 & n18378;
  assign n18452 = pi1154 & ~n18451;
  assign n18453 = ~n18450 & n18452;
  assign n18454 = pi627 & ~n18342;
  assign n18455 = ~n18453 & n18454;
  assign n18456 = ~pi618 & ~n18449;
  assign n18457 = pi618 & n18378;
  assign n18458 = ~pi1154 & ~n18457;
  assign n18459 = ~n18456 & n18458;
  assign n18460 = ~pi627 & ~n18340;
  assign n18461 = ~n18459 & n18460;
  assign n18462 = pi781 & ~n18461;
  assign n18463 = ~n18455 & n18462;
  assign n18464 = ~pi781 & n18449;
  assign n18465 = ~n11434 & ~n18464;
  assign n18466 = ~n18463 & n18465;
  assign n18467 = ~n18418 & ~n18466;
  assign n18468 = ~n18455 & ~n18461;
  assign n18469 = pi781 & ~n18468;
  assign n18470 = ~pi781 & ~n18449;
  assign n18471 = ~n18469 & ~n18470;
  assign n18472 = ~pi619 & ~n18471;
  assign n18473 = pi619 & n18379;
  assign n18474 = ~pi1159 & ~n18473;
  assign n18475 = ~n18472 & n18474;
  assign n18476 = ~pi648 & ~n18348;
  assign n18477 = ~n18475 & n18476;
  assign n18478 = pi619 & ~n18471;
  assign n18479 = ~pi619 & n18379;
  assign n18480 = pi1159 & ~n18479;
  assign n18481 = ~n18478 & n18480;
  assign n18482 = pi648 & ~n18350;
  assign n18483 = ~n18481 & n18482;
  assign n18484 = pi789 & ~n18483;
  assign n18485 = pi789 & ~n18477;
  assign n18486 = ~n18483 & n18485;
  assign n18487 = ~n18477 & n18484;
  assign n18488 = ~pi789 & n18471;
  assign n18489 = n62894 & ~n18488;
  assign n18490 = ~n63389 & n18489;
  assign n18491 = n62894 & ~n18467;
  assign n18492 = ~n18408 & ~n63390;
  assign n18493 = ~n63030 & ~n18492;
  assign n18494 = n8498 & n63386;
  assign n18495 = n8615 & n18381;
  assign n18496 = pi629 & ~n18495;
  assign n18497 = ~n18494 & n18496;
  assign n18498 = n8499 & n63386;
  assign n18499 = n8606 & n18381;
  assign n18500 = ~pi629 & ~n18499;
  assign n18501 = ~n18498 & n18500;
  assign n18502 = pi792 & ~n18501;
  assign n18503 = pi792 & ~n18497;
  assign n18504 = ~n18501 & n18503;
  assign n18505 = ~n18498 & ~n18499;
  assign n18506 = ~pi629 & ~n18505;
  assign n18507 = ~n18494 & ~n18495;
  assign n18508 = pi629 & ~n18507;
  assign n18509 = ~n18506 & ~n18508;
  assign n18510 = pi792 & ~n18509;
  assign n18511 = ~n18497 & n18502;
  assign n18512 = ~n8651 & ~n63391;
  assign n18513 = ~n18493 & n18512;
  assign n18514 = ~n18394 & ~n18513;
  assign n18515 = pi644 & n18514;
  assign n18516 = ~pi787 & ~n18382;
  assign n18517 = pi1157 & ~n18385;
  assign n18518 = ~n18390 & ~n18517;
  assign n18519 = pi787 & ~n18518;
  assign n18520 = ~n18516 & ~n18519;
  assign n18521 = ~pi644 & n18520;
  assign n18522 = pi715 & ~n18521;
  assign n18523 = ~n18515 & n18522;
  assign n18524 = ~n8685 & n18325;
  assign n18525 = ~n8376 & n18361;
  assign n18526 = ~n8376 & ~n18364;
  assign n18527 = n8376 & n18325;
  assign n18528 = ~n18526 & ~n18527;
  assign n18529 = ~n18524 & ~n18525;
  assign n18530 = pi644 & ~n63392;
  assign n18531 = ~pi644 & n18325;
  assign n18532 = ~pi715 & ~n18531;
  assign n18533 = ~n18530 & n18532;
  assign n18534 = pi1160 & ~n18533;
  assign n18535 = ~n18523 & n18534;
  assign n18536 = ~pi644 & n18514;
  assign n18537 = pi644 & n18520;
  assign n18538 = ~pi715 & ~n18537;
  assign n18539 = ~n18536 & n18538;
  assign n18540 = ~pi644 & ~n63392;
  assign n18541 = pi644 & n18325;
  assign n18542 = pi715 & ~n18541;
  assign n18543 = ~n18540 & n18542;
  assign n18544 = ~pi1160 & ~n18543;
  assign n18545 = ~n18539 & n18544;
  assign n18546 = ~n18535 & ~n18545;
  assign n18547 = pi790 & ~n18546;
  assign n18548 = ~pi790 & n18514;
  assign n18549 = pi832 & ~n18548;
  assign n18550 = ~n18547 & n18549;
  assign n18551 = ~pi183 & ~n8098;
  assign n18552 = n8257 & ~n18551;
  assign n18553 = ~pi725 & n62765;
  assign n18554 = n18551 & ~n18553;
  assign n18555 = pi183 & n62874;
  assign n18556 = ~pi38 & ~n18555;
  assign n18557 = n62765 & ~n18556;
  assign n18558 = ~pi183 & n8009;
  assign n18559 = ~n18557 & ~n18558;
  assign n18560 = ~pi183 & ~n7357;
  assign n18561 = n8085 & ~n18560;
  assign n18562 = ~pi725 & ~n18561;
  assign n18563 = ~n18559 & n18562;
  assign n18564 = ~n18554 & ~n18563;
  assign n18565 = ~pi778 & n18564;
  assign n18566 = pi625 & ~n18564;
  assign n18567 = ~pi625 & n18551;
  assign n18568 = pi1153 & ~n18567;
  assign n18569 = ~n18566 & n18568;
  assign n18570 = ~pi625 & ~n18564;
  assign n18571 = pi625 & n18551;
  assign n18572 = ~pi1153 & ~n18571;
  assign n18573 = ~n18570 & n18572;
  assign n18574 = ~n18569 & ~n18573;
  assign n18575 = pi778 & ~n18574;
  assign n18576 = ~n18565 & ~n18575;
  assign n18577 = ~n62880 & ~n18576;
  assign n18578 = n62880 & ~n18551;
  assign n18579 = ~n62880 & n18576;
  assign n18580 = n62880 & n18551;
  assign n18581 = ~n18579 & ~n18580;
  assign n18582 = ~n18577 & ~n18578;
  assign n18583 = ~n62882 & ~n63393;
  assign n18584 = n62882 & n18551;
  assign n18585 = n62882 & ~n18551;
  assign n18586 = ~n62882 & n63393;
  assign n18587 = ~n18585 & ~n18586;
  assign n18588 = ~n18583 & ~n18584;
  assign n18589 = ~n8257 & ~n63394;
  assign n18590 = ~n8257 & n63394;
  assign n18591 = n8257 & n18551;
  assign n18592 = ~n18590 & ~n18591;
  assign n18593 = ~n18552 & ~n18589;
  assign n18594 = ~n8303 & ~n63395;
  assign n18595 = n8303 & n18551;
  assign n18596 = ~n18594 & ~n18595;
  assign n18597 = ~pi792 & n18596;
  assign n18598 = pi628 & ~n18596;
  assign n18599 = ~pi628 & n18551;
  assign n18600 = pi1156 & ~n18599;
  assign n18601 = ~n18598 & n18600;
  assign n18602 = ~pi628 & ~n18596;
  assign n18603 = pi628 & n18551;
  assign n18604 = ~pi1156 & ~n18603;
  assign n18605 = ~n18602 & n18604;
  assign n18606 = ~n18601 & ~n18605;
  assign n18607 = pi792 & ~n18606;
  assign n18608 = ~n18597 & ~n18607;
  assign n18609 = pi647 & n18608;
  assign n18610 = ~pi647 & n18551;
  assign n18611 = pi1157 & ~n18610;
  assign n18612 = pi647 & ~n18608;
  assign n18613 = ~pi647 & ~n18551;
  assign n18614 = ~n18609 & ~n18610;
  assign n18615 = ~n18612 & ~n18613;
  assign n18616 = pi1157 & n63396;
  assign n18617 = ~n18609 & n18611;
  assign n18618 = ~pi647 & n18608;
  assign n18619 = pi647 & n18551;
  assign n18620 = ~pi1157 & ~n18619;
  assign n18621 = ~n18618 & n18620;
  assign n18622 = ~pi647 & ~n18608;
  assign n18623 = pi647 & ~n18551;
  assign n18624 = ~n18622 & ~n18623;
  assign n18625 = ~pi1157 & n18624;
  assign n18626 = pi1157 & ~n63396;
  assign n18627 = ~n18625 & ~n18626;
  assign n18628 = ~n63397 & ~n18621;
  assign n18629 = pi787 & n63398;
  assign n18630 = ~pi787 & ~n18608;
  assign n18631 = pi787 & ~n63398;
  assign n18632 = ~pi787 & n18608;
  assign n18633 = ~n18631 & ~n18632;
  assign n18634 = ~n18629 & ~n18630;
  assign n18635 = ~pi644 & ~n63399;
  assign n18636 = pi715 & ~n18635;
  assign n18637 = ~n11558 & n18551;
  assign n18638 = pi183 & ~n62765;
  assign n18639 = ~pi755 & n7359;
  assign n18640 = ~n18560 & ~n18639;
  assign n18641 = pi38 & ~n18640;
  assign n18642 = ~pi183 & n62802;
  assign n18643 = pi183 & ~n7351;
  assign n18644 = ~pi755 & ~n18643;
  assign n18645 = ~n18642 & n18644;
  assign n18646 = ~pi183 & pi755;
  assign n18647 = ~n62792 & n18646;
  assign n18648 = pi755 & ~n62792;
  assign n18649 = ~pi755 & ~n18642;
  assign n18650 = ~n18648 & ~n18649;
  assign n18651 = ~pi183 & ~n18650;
  assign n18652 = n7351 & n18649;
  assign n18653 = ~n18651 & ~n18652;
  assign n18654 = ~n18645 & ~n18647;
  assign n18655 = ~pi38 & ~n63400;
  assign n18656 = ~n18641 & ~n18655;
  assign n18657 = n62765 & n18656;
  assign n18658 = ~n18638 & ~n18657;
  assign n18659 = ~n8135 & ~n18658;
  assign n18660 = n8135 & ~n18551;
  assign n18661 = ~n18659 & ~n18660;
  assign n18662 = ~pi785 & ~n18661;
  assign n18663 = ~n8136 & ~n18551;
  assign n18664 = pi609 & n18659;
  assign n18665 = ~n18663 & ~n18664;
  assign n18666 = pi1155 & ~n18665;
  assign n18667 = ~n8148 & ~n18551;
  assign n18668 = ~pi609 & n18659;
  assign n18669 = ~n18667 & ~n18668;
  assign n18670 = ~pi1155 & ~n18669;
  assign n18671 = ~n18666 & ~n18670;
  assign n18672 = pi785 & ~n18671;
  assign n18673 = ~n18662 & ~n18672;
  assign n18674 = ~pi781 & ~n18673;
  assign n18675 = pi618 & n18673;
  assign n18676 = ~pi618 & n18551;
  assign n18677 = pi1154 & ~n18676;
  assign n18678 = ~n18675 & n18677;
  assign n18679 = ~pi618 & n18673;
  assign n18680 = pi618 & n18551;
  assign n18681 = ~pi1154 & ~n18680;
  assign n18682 = ~n18679 & n18681;
  assign n18683 = ~n18678 & ~n18682;
  assign n18684 = pi781 & ~n18683;
  assign n18685 = ~n18674 & ~n18684;
  assign n18686 = ~pi619 & ~n18685;
  assign n18687 = pi619 & ~n18551;
  assign n18688 = ~pi1159 & ~n18687;
  assign n18689 = ~n18686 & n18688;
  assign n18690 = pi619 & ~n18685;
  assign n18691 = ~pi619 & ~n18551;
  assign n18692 = pi1159 & ~n18691;
  assign n18693 = ~n18690 & n18692;
  assign n18694 = pi619 & n18685;
  assign n18695 = ~pi619 & n18551;
  assign n18696 = pi1159 & ~n18695;
  assign n18697 = ~n18694 & n18696;
  assign n18698 = ~pi619 & n18685;
  assign n18699 = pi619 & n18551;
  assign n18700 = ~pi1159 & ~n18699;
  assign n18701 = ~n18698 & n18700;
  assign n18702 = ~n18697 & ~n18701;
  assign n18703 = ~n18689 & ~n18693;
  assign n18704 = pi789 & n63401;
  assign n18705 = ~pi789 & n18685;
  assign n18706 = ~pi789 & ~n18685;
  assign n18707 = pi789 & ~n63401;
  assign n18708 = ~n18706 & ~n18707;
  assign n18709 = ~n18704 & ~n18705;
  assign n18710 = ~n8595 & n63402;
  assign n18711 = n8685 & n18710;
  assign n18712 = n8376 & ~n18551;
  assign n18713 = n8595 & n18551;
  assign n18714 = ~n18710 & ~n18713;
  assign n18715 = ~n8334 & ~n18714;
  assign n18716 = n8334 & n18551;
  assign n18717 = ~n18715 & ~n18716;
  assign n18718 = ~n8376 & n18717;
  assign n18719 = ~n18712 & ~n18718;
  assign n18720 = ~n8376 & ~n18717;
  assign n18721 = n8376 & n18551;
  assign n18722 = ~n18720 & ~n18721;
  assign n18723 = ~n18637 & ~n18711;
  assign n18724 = pi644 & n63403;
  assign n18725 = ~pi644 & n18551;
  assign n18726 = ~pi715 & ~n18725;
  assign n18727 = ~n18724 & n18726;
  assign n18728 = pi1160 & ~n18727;
  assign n18729 = ~n18636 & n18728;
  assign n18730 = pi644 & ~n63399;
  assign n18731 = ~pi715 & ~n18730;
  assign n18732 = ~pi644 & n63403;
  assign n18733 = pi644 & n18551;
  assign n18734 = pi715 & ~n18733;
  assign n18735 = ~n18732 & n18734;
  assign n18736 = ~pi1160 & ~n18735;
  assign n18737 = ~n18731 & n18736;
  assign n18738 = ~n18729 & ~n18737;
  assign n18739 = pi790 & ~n18738;
  assign n18740 = ~n63052 & n18714;
  assign n18741 = ~pi629 & n18601;
  assign n18742 = pi629 & n18605;
  assign n18743 = ~n18741 & ~n18742;
  assign n18744 = ~n18740 & n18743;
  assign n18745 = pi792 & ~n18744;
  assign n18746 = pi725 & ~n18656;
  assign n18747 = ~pi183 & ~n62821;
  assign n18748 = pi183 & n7632;
  assign n18749 = pi755 & ~n18748;
  assign n18750 = ~n18747 & n18749;
  assign n18751 = pi183 & n7709;
  assign n18752 = ~pi183 & n62851;
  assign n18753 = ~pi755 & ~n18752;
  assign n18754 = ~n18751 & n18753;
  assign n18755 = pi39 & ~n18754;
  assign n18756 = ~n18750 & n18755;
  assign n18757 = pi183 & n7855;
  assign n18758 = ~pi183 & n7832;
  assign n18759 = pi755 & ~n18758;
  assign n18760 = ~n18757 & n18759;
  assign n18761 = ~pi183 & ~n7861;
  assign n18762 = pi183 & ~n7868;
  assign n18763 = ~pi755 & ~n18762;
  assign n18764 = ~n18761 & n18763;
  assign n18765 = ~pi39 & ~n18764;
  assign n18766 = pi183 & ~n7855;
  assign n18767 = ~pi183 & ~n7832;
  assign n18768 = pi755 & ~n18767;
  assign n18769 = pi755 & ~n18766;
  assign n18770 = ~n18767 & n18769;
  assign n18771 = ~n18766 & n18768;
  assign n18772 = ~pi183 & n7861;
  assign n18773 = pi183 & n7868;
  assign n18774 = ~pi755 & ~n18773;
  assign n18775 = ~n18772 & n18774;
  assign n18776 = ~n63404 & ~n18775;
  assign n18777 = ~pi39 & ~n18776;
  assign n18778 = ~n18760 & n18765;
  assign n18779 = ~pi38 & ~n63405;
  assign n18780 = ~n18756 & n18779;
  assign n18781 = ~pi755 & ~n7744;
  assign n18782 = n10350 & ~n18781;
  assign n18783 = ~pi183 & ~n18782;
  assign n18784 = ~n7565 & ~n18326;
  assign n18785 = pi183 & ~n18784;
  assign n18786 = n7356 & n18785;
  assign n18787 = pi38 & ~n18786;
  assign n18788 = ~n18783 & n18787;
  assign n18789 = ~pi725 & ~n18788;
  assign n18790 = ~n18780 & n18789;
  assign n18791 = n62765 & ~n18790;
  assign n18792 = ~n18746 & n18791;
  assign n18793 = ~n18638 & ~n18792;
  assign n18794 = ~pi625 & n18793;
  assign n18795 = pi625 & n18658;
  assign n18796 = ~pi1153 & ~n18795;
  assign n18797 = ~n18794 & n18796;
  assign n18798 = ~pi608 & ~n18569;
  assign n18799 = ~n18797 & n18798;
  assign n18800 = pi625 & n18793;
  assign n18801 = ~pi625 & n18658;
  assign n18802 = pi1153 & ~n18801;
  assign n18803 = ~n18800 & n18802;
  assign n18804 = pi608 & ~n18573;
  assign n18805 = ~n18803 & n18804;
  assign n18806 = ~n18799 & ~n18805;
  assign n18807 = pi778 & ~n18806;
  assign n18808 = ~pi778 & n18793;
  assign n18809 = ~n18807 & ~n18808;
  assign n18810 = ~pi609 & ~n18809;
  assign n18811 = pi609 & n18576;
  assign n18812 = ~pi1155 & ~n18811;
  assign n18813 = ~n18810 & n18812;
  assign n18814 = ~pi660 & ~n18666;
  assign n18815 = ~n18813 & n18814;
  assign n18816 = pi609 & ~n18809;
  assign n18817 = ~pi609 & n18576;
  assign n18818 = pi1155 & ~n18817;
  assign n18819 = ~n18816 & n18818;
  assign n18820 = pi660 & ~n18670;
  assign n18821 = ~n18819 & n18820;
  assign n18822 = ~n18815 & ~n18821;
  assign n18823 = pi785 & ~n18822;
  assign n18824 = ~pi785 & ~n18809;
  assign n18825 = ~n18823 & ~n18824;
  assign n18826 = pi618 & ~n18825;
  assign n18827 = ~pi618 & ~n63393;
  assign n18828 = pi1154 & ~n18827;
  assign n18829 = ~n18826 & n18828;
  assign n18830 = pi627 & ~n18682;
  assign n18831 = ~n18829 & n18830;
  assign n18832 = ~pi618 & ~n18825;
  assign n18833 = pi618 & ~n63393;
  assign n18834 = ~pi1154 & ~n18833;
  assign n18835 = ~n18832 & n18834;
  assign n18836 = ~pi627 & ~n18678;
  assign n18837 = ~n18835 & n18836;
  assign n18838 = pi781 & ~n18837;
  assign n18839 = ~n18831 & n18838;
  assign n18840 = ~n11431 & ~n63394;
  assign n18841 = ~n62884 & ~n63401;
  assign n18842 = ~n18840 & ~n18841;
  assign n18843 = pi789 & ~n18842;
  assign n18844 = ~pi781 & n18825;
  assign n18845 = ~n18843 & ~n18844;
  assign n18846 = ~n18839 & n18845;
  assign n18847 = n11434 & n18842;
  assign n18848 = ~n18846 & ~n18847;
  assign n18849 = ~n18831 & ~n18837;
  assign n18850 = pi781 & ~n18849;
  assign n18851 = ~pi781 & ~n18825;
  assign n18852 = ~n18850 & ~n18851;
  assign n18853 = ~pi619 & ~n18852;
  assign n18854 = pi619 & n63394;
  assign n18855 = ~pi1159 & ~n18854;
  assign n18856 = ~n18853 & n18855;
  assign n18857 = ~pi648 & ~n18697;
  assign n18858 = ~n18856 & n18857;
  assign n18859 = pi619 & ~n18852;
  assign n18860 = ~pi619 & n63394;
  assign n18861 = pi1159 & ~n18860;
  assign n18862 = ~n18859 & n18861;
  assign n18863 = pi648 & ~n18701;
  assign n18864 = ~n18862 & n18863;
  assign n18865 = pi789 & ~n18864;
  assign n18866 = pi789 & ~n18858;
  assign n18867 = ~n18864 & n18866;
  assign n18868 = ~n18858 & n18865;
  assign n18869 = ~pi789 & n18852;
  assign n18870 = n62894 & ~n18869;
  assign n18871 = ~n63406 & n18870;
  assign n18872 = n62894 & ~n18848;
  assign n18873 = ~pi626 & ~n63402;
  assign n18874 = pi626 & ~n18551;
  assign n18875 = n8301 & ~n18874;
  assign n18876 = ~n18873 & n18875;
  assign n18877 = n8525 & ~n63395;
  assign n18878 = pi626 & ~n63402;
  assign n18879 = ~pi626 & ~n18551;
  assign n18880 = n8300 & ~n18879;
  assign n18881 = ~n18878 & n18880;
  assign n18882 = ~n18877 & ~n18881;
  assign n18883 = ~n18876 & ~n18877;
  assign n18884 = ~n18881 & n18883;
  assign n18885 = ~n18876 & n18882;
  assign n18886 = pi788 & ~n63408;
  assign n18887 = ~n63030 & ~n18886;
  assign n18888 = ~n63407 & n18887;
  assign n18889 = ~n18745 & ~n18888;
  assign n18890 = ~n8651 & ~n18889;
  assign n18891 = ~n8413 & ~n18716;
  assign n18892 = ~n8413 & n18717;
  assign n18893 = ~n18715 & n18891;
  assign n18894 = n8373 & n63396;
  assign n18895 = ~pi630 & n63397;
  assign n18896 = n8374 & ~n18624;
  assign n18897 = pi630 & n18621;
  assign n18898 = ~n63410 & ~n63411;
  assign n18899 = ~n63409 & n18898;
  assign n18900 = pi787 & ~n18899;
  assign n18901 = ~pi644 & n18736;
  assign n18902 = pi644 & n18728;
  assign n18903 = n14029 & ~n18727;
  assign n18904 = pi790 & ~n63412;
  assign n18905 = pi790 & ~n18901;
  assign n18906 = ~n63412 & n18905;
  assign n18907 = ~n18901 & n18904;
  assign n18908 = ~n18900 & ~n63413;
  assign n18909 = ~n18890 & ~n18900;
  assign n18910 = ~n63413 & n18909;
  assign n18911 = ~n18890 & n18908;
  assign n18912 = ~n18739 & ~n63414;
  assign n18913 = n62455 & ~n18912;
  assign n18914 = ~pi183 & ~n62455;
  assign n18915 = ~pi832 & ~n18914;
  assign n18916 = ~n18913 & n18915;
  assign po340 = ~n18550 & ~n18916;
  assign n18918 = ~pi184 & ~n2923;
  assign n18919 = ~pi777 & n7316;
  assign n18920 = ~n18918 & ~n18919;
  assign n18921 = ~n8420 & ~n18920;
  assign n18922 = ~pi785 & ~n18921;
  assign n18923 = n8148 & n18919;
  assign n18924 = n18921 & ~n18923;
  assign n18925 = pi1155 & ~n18924;
  assign n18926 = ~pi1155 & ~n18918;
  assign n18927 = ~n18923 & n18926;
  assign n18928 = ~n18925 & ~n18927;
  assign n18929 = pi785 & ~n18928;
  assign n18930 = ~n18922 & ~n18929;
  assign n18931 = ~pi781 & ~n18930;
  assign n18932 = ~n8435 & n18930;
  assign n18933 = pi1154 & ~n18932;
  assign n18934 = ~n8438 & n18930;
  assign n18935 = ~pi1154 & ~n18934;
  assign n18936 = ~n18933 & ~n18935;
  assign n18937 = pi781 & ~n18936;
  assign n18938 = ~n18931 & ~n18937;
  assign n18939 = ~pi789 & ~n18938;
  assign n18940 = ~n12612 & n18938;
  assign n18941 = pi1159 & ~n18940;
  assign n18942 = ~n12615 & n18938;
  assign n18943 = ~pi1159 & ~n18942;
  assign n18944 = ~n18941 & ~n18943;
  assign n18945 = pi789 & ~n18944;
  assign n18946 = ~n18939 & ~n18945;
  assign n18947 = ~n15298 & n18938;
  assign n18948 = ~n8595 & n63415;
  assign n18949 = n8595 & n18918;
  assign n18950 = ~n8595 & ~n63415;
  assign n18951 = n8595 & ~n18918;
  assign n18952 = ~n18950 & ~n18951;
  assign n18953 = ~n18948 & ~n18949;
  assign n18954 = ~n8334 & n63416;
  assign n18955 = n8334 & n18918;
  assign n18956 = ~n8413 & ~n18955;
  assign n18957 = ~n18954 & ~n18955;
  assign n18958 = ~n8413 & n18957;
  assign n18959 = ~n18954 & n18956;
  assign n18960 = ~pi737 & n7564;
  assign n18961 = ~n18918 & ~n18960;
  assign n18962 = ~pi778 & ~n18961;
  assign n18963 = ~pi625 & n18960;
  assign n18964 = ~n18961 & ~n18963;
  assign n18965 = pi1153 & ~n18964;
  assign n18966 = ~pi1153 & ~n18918;
  assign n18967 = ~n18963 & n18966;
  assign n18968 = pi778 & ~n18967;
  assign n18969 = ~n18965 & n18968;
  assign n18970 = ~n18962 & ~n18969;
  assign n18971 = ~n8490 & ~n18970;
  assign n18972 = ~n8492 & n18971;
  assign n18973 = ~n8494 & n18972;
  assign n18974 = ~n8496 & n18973;
  assign n18975 = ~n8508 & n18974;
  assign n18976 = pi647 & ~n18975;
  assign n18977 = ~pi647 & ~n18918;
  assign n18978 = ~n18976 & ~n18977;
  assign n18979 = n8373 & ~n18978;
  assign n18980 = ~pi647 & n18975;
  assign n18981 = pi647 & n18918;
  assign n18982 = ~pi1157 & ~n18981;
  assign n18983 = ~n18980 & n18982;
  assign n18984 = pi630 & n18983;
  assign n18985 = ~n18979 & ~n18984;
  assign n18986 = ~n63417 & n18985;
  assign n18987 = pi787 & ~n18986;
  assign n18988 = ~pi626 & ~n63415;
  assign n18989 = pi626 & ~n18918;
  assign n18990 = n8301 & ~n18989;
  assign n18991 = ~n18988 & n18990;
  assign n18992 = n8525 & n18973;
  assign n18993 = pi626 & ~n63415;
  assign n18994 = ~pi626 & ~n18918;
  assign n18995 = n8300 & ~n18994;
  assign n18996 = ~n18993 & n18995;
  assign n18997 = ~n18992 & ~n18996;
  assign n18998 = ~n18991 & ~n18992;
  assign n18999 = ~n18996 & n18998;
  assign n19000 = ~n18991 & n18997;
  assign n19001 = pi788 & ~n63418;
  assign n19002 = n13460 & n18938;
  assign n19003 = n11303 & n18972;
  assign n19004 = pi648 & ~n19003;
  assign n19005 = ~n19002 & n19004;
  assign n19006 = n13462 & n18938;
  assign n19007 = n11304 & n18972;
  assign n19008 = ~pi648 & ~n19007;
  assign n19009 = ~n19006 & n19008;
  assign n19010 = pi789 & ~n19009;
  assign n19011 = ~n19005 & n19010;
  assign n19012 = ~n7187 & ~n18961;
  assign n19013 = pi625 & n19012;
  assign n19014 = n18920 & ~n19012;
  assign n19015 = ~n19013 & ~n19014;
  assign n19016 = n18966 & ~n19015;
  assign n19017 = ~pi608 & ~n18965;
  assign n19018 = ~n19016 & n19017;
  assign n19019 = pi1153 & n18920;
  assign n19020 = ~n19013 & n19019;
  assign n19021 = pi608 & ~n18967;
  assign n19022 = ~n19020 & n19021;
  assign n19023 = ~n19018 & ~n19022;
  assign n19024 = pi778 & ~n19023;
  assign n19025 = ~pi778 & ~n19014;
  assign n19026 = ~n19024 & ~n19025;
  assign n19027 = ~pi609 & ~n19026;
  assign n19028 = pi609 & ~n18970;
  assign n19029 = ~pi1155 & ~n19028;
  assign n19030 = ~n19027 & n19029;
  assign n19031 = ~pi660 & ~n18925;
  assign n19032 = ~n19030 & n19031;
  assign n19033 = pi609 & ~n19026;
  assign n19034 = ~pi609 & ~n18970;
  assign n19035 = pi1155 & ~n19034;
  assign n19036 = ~n19033 & n19035;
  assign n19037 = pi660 & ~n18927;
  assign n19038 = ~n19036 & n19037;
  assign n19039 = ~n19032 & ~n19038;
  assign n19040 = pi785 & ~n19039;
  assign n19041 = ~pi785 & ~n19026;
  assign n19042 = ~n19040 & ~n19041;
  assign n19043 = pi618 & ~n19042;
  assign n19044 = ~pi618 & n18971;
  assign n19045 = pi1154 & ~n19044;
  assign n19046 = ~n19043 & n19045;
  assign n19047 = pi627 & ~n18935;
  assign n19048 = ~n19046 & n19047;
  assign n19049 = ~pi618 & ~n19042;
  assign n19050 = pi618 & n18971;
  assign n19051 = ~pi1154 & ~n19050;
  assign n19052 = ~n19049 & n19051;
  assign n19053 = ~pi627 & ~n18933;
  assign n19054 = ~n19052 & n19053;
  assign n19055 = pi781 & ~n19054;
  assign n19056 = ~n19048 & n19055;
  assign n19057 = ~pi781 & n19042;
  assign n19058 = ~n11434 & ~n19057;
  assign n19059 = ~n19056 & n19058;
  assign n19060 = ~n19011 & ~n19059;
  assign n19061 = ~n19048 & ~n19054;
  assign n19062 = pi781 & ~n19061;
  assign n19063 = ~pi781 & ~n19042;
  assign n19064 = ~n19062 & ~n19063;
  assign n19065 = ~pi619 & ~n19064;
  assign n19066 = pi619 & n18972;
  assign n19067 = ~pi1159 & ~n19066;
  assign n19068 = ~n19065 & n19067;
  assign n19069 = ~pi648 & ~n18941;
  assign n19070 = ~n19068 & n19069;
  assign n19071 = pi619 & ~n19064;
  assign n19072 = ~pi619 & n18972;
  assign n19073 = pi1159 & ~n19072;
  assign n19074 = ~n19071 & n19073;
  assign n19075 = pi648 & ~n18943;
  assign n19076 = ~n19074 & n19075;
  assign n19077 = pi789 & ~n19076;
  assign n19078 = pi789 & ~n19070;
  assign n19079 = ~n19076 & n19078;
  assign n19080 = ~n19070 & n19077;
  assign n19081 = ~pi789 & n19064;
  assign n19082 = n62894 & ~n19081;
  assign n19083 = ~n63419 & n19082;
  assign n19084 = n62894 & ~n19060;
  assign n19085 = ~n19001 & ~n63420;
  assign n19086 = ~n63030 & ~n19085;
  assign n19087 = n8498 & n63416;
  assign n19088 = n8615 & n18974;
  assign n19089 = pi629 & ~n19088;
  assign n19090 = ~n19087 & n19089;
  assign n19091 = n8499 & n63416;
  assign n19092 = n8606 & n18974;
  assign n19093 = ~pi629 & ~n19092;
  assign n19094 = ~n19091 & n19093;
  assign n19095 = pi792 & ~n19094;
  assign n19096 = pi792 & ~n19090;
  assign n19097 = ~n19094 & n19096;
  assign n19098 = ~n19091 & ~n19092;
  assign n19099 = ~pi629 & ~n19098;
  assign n19100 = ~n19087 & ~n19088;
  assign n19101 = pi629 & ~n19100;
  assign n19102 = ~n19099 & ~n19101;
  assign n19103 = pi792 & ~n19102;
  assign n19104 = ~n19090 & n19095;
  assign n19105 = ~n8651 & ~n63421;
  assign n19106 = ~n19086 & n19105;
  assign n19107 = ~n18987 & ~n19106;
  assign n19108 = pi644 & n19107;
  assign n19109 = ~pi787 & ~n18975;
  assign n19110 = pi1157 & ~n18978;
  assign n19111 = ~n18983 & ~n19110;
  assign n19112 = pi787 & ~n19111;
  assign n19113 = ~n19109 & ~n19112;
  assign n19114 = ~pi644 & n19113;
  assign n19115 = pi715 & ~n19114;
  assign n19116 = ~n19108 & n19115;
  assign n19117 = ~n8685 & n18918;
  assign n19118 = ~n8376 & n18954;
  assign n19119 = ~n8376 & ~n18957;
  assign n19120 = n8376 & n18918;
  assign n19121 = ~n19119 & ~n19120;
  assign n19122 = ~n19117 & ~n19118;
  assign n19123 = pi644 & ~n63422;
  assign n19124 = ~pi644 & n18918;
  assign n19125 = ~pi715 & ~n19124;
  assign n19126 = ~n19123 & n19125;
  assign n19127 = pi1160 & ~n19126;
  assign n19128 = ~n19116 & n19127;
  assign n19129 = ~pi644 & n19107;
  assign n19130 = pi644 & n19113;
  assign n19131 = ~pi715 & ~n19130;
  assign n19132 = ~n19129 & n19131;
  assign n19133 = ~pi644 & ~n63422;
  assign n19134 = pi644 & n18918;
  assign n19135 = pi715 & ~n19134;
  assign n19136 = ~n19133 & n19135;
  assign n19137 = ~pi1160 & ~n19136;
  assign n19138 = ~n19132 & n19137;
  assign n19139 = ~n19128 & ~n19138;
  assign n19140 = pi790 & ~n19139;
  assign n19141 = ~pi790 & n19107;
  assign n19142 = pi832 & ~n19141;
  assign n19143 = ~n19140 & n19142;
  assign n19144 = ~pi184 & ~n8098;
  assign n19145 = n8257 & ~n19144;
  assign n19146 = ~pi737 & n62765;
  assign n19147 = n19144 & ~n19146;
  assign n19148 = pi184 & n62874;
  assign n19149 = ~pi38 & ~n19148;
  assign n19150 = n62765 & ~n19149;
  assign n19151 = ~pi184 & n8009;
  assign n19152 = ~n19150 & ~n19151;
  assign n19153 = ~pi184 & ~n7357;
  assign n19154 = n8085 & ~n19153;
  assign n19155 = ~pi737 & ~n19154;
  assign n19156 = ~n19152 & n19155;
  assign n19157 = ~n19147 & ~n19156;
  assign n19158 = ~pi778 & n19157;
  assign n19159 = pi625 & ~n19157;
  assign n19160 = ~pi625 & n19144;
  assign n19161 = pi1153 & ~n19160;
  assign n19162 = ~n19159 & n19161;
  assign n19163 = ~pi625 & ~n19157;
  assign n19164 = pi625 & n19144;
  assign n19165 = ~pi1153 & ~n19164;
  assign n19166 = ~n19163 & n19165;
  assign n19167 = ~n19162 & ~n19166;
  assign n19168 = pi778 & ~n19167;
  assign n19169 = ~n19158 & ~n19168;
  assign n19170 = ~n62880 & ~n19169;
  assign n19171 = n62880 & ~n19144;
  assign n19172 = ~n62880 & n19169;
  assign n19173 = n62880 & n19144;
  assign n19174 = ~n19172 & ~n19173;
  assign n19175 = ~n19170 & ~n19171;
  assign n19176 = ~n62882 & ~n63423;
  assign n19177 = n62882 & n19144;
  assign n19178 = n62882 & ~n19144;
  assign n19179 = ~n62882 & n63423;
  assign n19180 = ~n19178 & ~n19179;
  assign n19181 = ~n19176 & ~n19177;
  assign n19182 = ~n8257 & ~n63424;
  assign n19183 = ~n8257 & n63424;
  assign n19184 = n8257 & n19144;
  assign n19185 = ~n19183 & ~n19184;
  assign n19186 = ~n19145 & ~n19182;
  assign n19187 = ~n8303 & ~n63425;
  assign n19188 = n8303 & n19144;
  assign n19189 = ~n19187 & ~n19188;
  assign n19190 = ~pi792 & n19189;
  assign n19191 = pi628 & ~n19189;
  assign n19192 = ~pi628 & n19144;
  assign n19193 = pi1156 & ~n19192;
  assign n19194 = ~n19191 & n19193;
  assign n19195 = ~pi628 & ~n19189;
  assign n19196 = pi628 & n19144;
  assign n19197 = ~pi1156 & ~n19196;
  assign n19198 = ~n19195 & n19197;
  assign n19199 = ~n19194 & ~n19198;
  assign n19200 = pi792 & ~n19199;
  assign n19201 = ~n19190 & ~n19200;
  assign n19202 = pi647 & n19201;
  assign n19203 = ~pi647 & n19144;
  assign n19204 = pi1157 & ~n19203;
  assign n19205 = pi647 & ~n19201;
  assign n19206 = ~pi647 & ~n19144;
  assign n19207 = ~n19202 & ~n19203;
  assign n19208 = ~n19205 & ~n19206;
  assign n19209 = pi1157 & n63426;
  assign n19210 = ~n19202 & n19204;
  assign n19211 = ~pi647 & n19201;
  assign n19212 = pi647 & n19144;
  assign n19213 = ~pi1157 & ~n19212;
  assign n19214 = ~n19211 & n19213;
  assign n19215 = ~pi647 & ~n19201;
  assign n19216 = pi647 & ~n19144;
  assign n19217 = ~n19215 & ~n19216;
  assign n19218 = ~pi1157 & n19217;
  assign n19219 = pi1157 & ~n63426;
  assign n19220 = ~n19218 & ~n19219;
  assign n19221 = ~n63427 & ~n19214;
  assign n19222 = pi787 & n63428;
  assign n19223 = ~pi787 & ~n19201;
  assign n19224 = pi787 & ~n63428;
  assign n19225 = ~pi787 & n19201;
  assign n19226 = ~n19224 & ~n19225;
  assign n19227 = ~n19222 & ~n19223;
  assign n19228 = ~pi644 & ~n63429;
  assign n19229 = pi715 & ~n19228;
  assign n19230 = ~n11558 & n19144;
  assign n19231 = pi184 & ~n62765;
  assign n19232 = ~pi777 & n7359;
  assign n19233 = ~n19153 & ~n19232;
  assign n19234 = pi38 & ~n19233;
  assign n19235 = ~pi184 & n62802;
  assign n19236 = pi184 & ~n7351;
  assign n19237 = ~pi777 & ~n19236;
  assign n19238 = ~n19235 & n19237;
  assign n19239 = ~pi184 & pi777;
  assign n19240 = ~n62792 & n19239;
  assign n19241 = pi777 & ~n62792;
  assign n19242 = ~pi777 & ~n19235;
  assign n19243 = ~n19241 & ~n19242;
  assign n19244 = ~pi184 & ~n19243;
  assign n19245 = n7351 & n19242;
  assign n19246 = ~n19244 & ~n19245;
  assign n19247 = ~n19238 & ~n19240;
  assign n19248 = ~pi38 & ~n63430;
  assign n19249 = ~n19234 & ~n19248;
  assign n19250 = n62765 & n19249;
  assign n19251 = ~n19231 & ~n19250;
  assign n19252 = ~n8135 & ~n19251;
  assign n19253 = n8135 & ~n19144;
  assign n19254 = ~n19252 & ~n19253;
  assign n19255 = ~pi785 & ~n19254;
  assign n19256 = ~n8136 & ~n19144;
  assign n19257 = pi609 & n19252;
  assign n19258 = ~n19256 & ~n19257;
  assign n19259 = pi1155 & ~n19258;
  assign n19260 = ~n8148 & ~n19144;
  assign n19261 = ~pi609 & n19252;
  assign n19262 = ~n19260 & ~n19261;
  assign n19263 = ~pi1155 & ~n19262;
  assign n19264 = ~n19259 & ~n19263;
  assign n19265 = pi785 & ~n19264;
  assign n19266 = ~n19255 & ~n19265;
  assign n19267 = ~pi781 & ~n19266;
  assign n19268 = pi618 & n19266;
  assign n19269 = ~pi618 & n19144;
  assign n19270 = pi1154 & ~n19269;
  assign n19271 = ~n19268 & n19270;
  assign n19272 = ~pi618 & n19266;
  assign n19273 = pi618 & n19144;
  assign n19274 = ~pi1154 & ~n19273;
  assign n19275 = ~n19272 & n19274;
  assign n19276 = ~n19271 & ~n19275;
  assign n19277 = pi781 & ~n19276;
  assign n19278 = ~n19267 & ~n19277;
  assign n19279 = ~pi619 & ~n19278;
  assign n19280 = pi619 & ~n19144;
  assign n19281 = ~pi1159 & ~n19280;
  assign n19282 = ~n19279 & n19281;
  assign n19283 = pi619 & ~n19278;
  assign n19284 = ~pi619 & ~n19144;
  assign n19285 = pi1159 & ~n19284;
  assign n19286 = ~n19283 & n19285;
  assign n19287 = pi619 & n19278;
  assign n19288 = ~pi619 & n19144;
  assign n19289 = pi1159 & ~n19288;
  assign n19290 = ~n19287 & n19289;
  assign n19291 = ~pi619 & n19278;
  assign n19292 = pi619 & n19144;
  assign n19293 = ~pi1159 & ~n19292;
  assign n19294 = ~n19291 & n19293;
  assign n19295 = ~n19290 & ~n19294;
  assign n19296 = ~n19282 & ~n19286;
  assign n19297 = pi789 & n63431;
  assign n19298 = ~pi789 & n19278;
  assign n19299 = ~pi789 & ~n19278;
  assign n19300 = pi789 & ~n63431;
  assign n19301 = ~n19299 & ~n19300;
  assign n19302 = ~n19297 & ~n19298;
  assign n19303 = ~n8595 & n63432;
  assign n19304 = n8685 & n19303;
  assign n19305 = n8376 & ~n19144;
  assign n19306 = n8595 & n19144;
  assign n19307 = ~n19303 & ~n19306;
  assign n19308 = ~n8334 & ~n19307;
  assign n19309 = n8334 & n19144;
  assign n19310 = ~n19308 & ~n19309;
  assign n19311 = ~n8376 & n19310;
  assign n19312 = ~n19305 & ~n19311;
  assign n19313 = ~n8376 & ~n19310;
  assign n19314 = n8376 & n19144;
  assign n19315 = ~n19313 & ~n19314;
  assign n19316 = ~n19230 & ~n19304;
  assign n19317 = pi644 & n63433;
  assign n19318 = ~pi644 & n19144;
  assign n19319 = ~pi715 & ~n19318;
  assign n19320 = ~n19317 & n19319;
  assign n19321 = pi1160 & ~n19320;
  assign n19322 = ~n19229 & n19321;
  assign n19323 = pi644 & ~n63429;
  assign n19324 = ~pi715 & ~n19323;
  assign n19325 = ~pi644 & n63433;
  assign n19326 = pi644 & n19144;
  assign n19327 = pi715 & ~n19326;
  assign n19328 = ~n19325 & n19327;
  assign n19329 = ~pi1160 & ~n19328;
  assign n19330 = ~n19324 & n19329;
  assign n19331 = ~n19322 & ~n19330;
  assign n19332 = pi790 & ~n19331;
  assign n19333 = ~n63052 & n19307;
  assign n19334 = ~pi629 & n19194;
  assign n19335 = pi629 & n19198;
  assign n19336 = ~n19334 & ~n19335;
  assign n19337 = ~n19333 & n19336;
  assign n19338 = pi792 & ~n19337;
  assign n19339 = pi737 & ~n19249;
  assign n19340 = ~pi184 & ~n62821;
  assign n19341 = pi184 & n7632;
  assign n19342 = pi777 & ~n19341;
  assign n19343 = ~n19340 & n19342;
  assign n19344 = pi184 & n7709;
  assign n19345 = ~pi184 & n62851;
  assign n19346 = ~pi777 & ~n19345;
  assign n19347 = ~n19344 & n19346;
  assign n19348 = pi39 & ~n19347;
  assign n19349 = ~n19343 & n19348;
  assign n19350 = pi184 & n7855;
  assign n19351 = ~pi184 & n7832;
  assign n19352 = pi777 & ~n19351;
  assign n19353 = ~n19350 & n19352;
  assign n19354 = ~pi184 & ~n7861;
  assign n19355 = pi184 & ~n7868;
  assign n19356 = ~pi777 & ~n19355;
  assign n19357 = ~n19354 & n19356;
  assign n19358 = ~pi39 & ~n19357;
  assign n19359 = pi184 & ~n7855;
  assign n19360 = ~pi184 & ~n7832;
  assign n19361 = pi777 & ~n19360;
  assign n19362 = pi777 & ~n19359;
  assign n19363 = ~n19360 & n19362;
  assign n19364 = ~n19359 & n19361;
  assign n19365 = ~pi184 & n7861;
  assign n19366 = pi184 & n7868;
  assign n19367 = ~pi777 & ~n19366;
  assign n19368 = ~n19365 & n19367;
  assign n19369 = ~n63434 & ~n19368;
  assign n19370 = ~pi39 & ~n19369;
  assign n19371 = ~n19353 & n19358;
  assign n19372 = ~pi38 & ~n63435;
  assign n19373 = ~n19349 & n19372;
  assign n19374 = ~pi777 & ~n7744;
  assign n19375 = n10350 & ~n19374;
  assign n19376 = ~pi184 & ~n19375;
  assign n19377 = ~n7565 & ~n18919;
  assign n19378 = pi184 & ~n19377;
  assign n19379 = n7356 & n19378;
  assign n19380 = pi38 & ~n19379;
  assign n19381 = ~n19376 & n19380;
  assign n19382 = ~pi737 & ~n19381;
  assign n19383 = ~n19373 & n19382;
  assign n19384 = n62765 & ~n19383;
  assign n19385 = ~n19339 & n19384;
  assign n19386 = ~n19231 & ~n19385;
  assign n19387 = ~pi625 & n19386;
  assign n19388 = pi625 & n19251;
  assign n19389 = ~pi1153 & ~n19388;
  assign n19390 = ~n19387 & n19389;
  assign n19391 = ~pi608 & ~n19162;
  assign n19392 = ~n19390 & n19391;
  assign n19393 = pi625 & n19386;
  assign n19394 = ~pi625 & n19251;
  assign n19395 = pi1153 & ~n19394;
  assign n19396 = ~n19393 & n19395;
  assign n19397 = pi608 & ~n19166;
  assign n19398 = ~n19396 & n19397;
  assign n19399 = ~n19392 & ~n19398;
  assign n19400 = pi778 & ~n19399;
  assign n19401 = ~pi778 & n19386;
  assign n19402 = ~n19400 & ~n19401;
  assign n19403 = ~pi609 & ~n19402;
  assign n19404 = pi609 & n19169;
  assign n19405 = ~pi1155 & ~n19404;
  assign n19406 = ~n19403 & n19405;
  assign n19407 = ~pi660 & ~n19259;
  assign n19408 = ~n19406 & n19407;
  assign n19409 = pi609 & ~n19402;
  assign n19410 = ~pi609 & n19169;
  assign n19411 = pi1155 & ~n19410;
  assign n19412 = ~n19409 & n19411;
  assign n19413 = pi660 & ~n19263;
  assign n19414 = ~n19412 & n19413;
  assign n19415 = ~n19408 & ~n19414;
  assign n19416 = pi785 & ~n19415;
  assign n19417 = ~pi785 & ~n19402;
  assign n19418 = ~n19416 & ~n19417;
  assign n19419 = pi618 & ~n19418;
  assign n19420 = ~pi618 & ~n63423;
  assign n19421 = pi1154 & ~n19420;
  assign n19422 = ~n19419 & n19421;
  assign n19423 = pi627 & ~n19275;
  assign n19424 = ~n19422 & n19423;
  assign n19425 = ~pi618 & ~n19418;
  assign n19426 = pi618 & ~n63423;
  assign n19427 = ~pi1154 & ~n19426;
  assign n19428 = ~n19425 & n19427;
  assign n19429 = ~pi627 & ~n19271;
  assign n19430 = ~n19428 & n19429;
  assign n19431 = pi781 & ~n19430;
  assign n19432 = ~n19424 & n19431;
  assign n19433 = ~n11431 & ~n63424;
  assign n19434 = ~n62884 & ~n63431;
  assign n19435 = ~n19433 & ~n19434;
  assign n19436 = pi789 & ~n19435;
  assign n19437 = ~pi781 & n19418;
  assign n19438 = ~n19436 & ~n19437;
  assign n19439 = ~n19432 & n19438;
  assign n19440 = n11434 & n19435;
  assign n19441 = ~n19439 & ~n19440;
  assign n19442 = ~n19424 & ~n19430;
  assign n19443 = pi781 & ~n19442;
  assign n19444 = ~pi781 & ~n19418;
  assign n19445 = ~n19443 & ~n19444;
  assign n19446 = ~pi619 & ~n19445;
  assign n19447 = pi619 & n63424;
  assign n19448 = ~pi1159 & ~n19447;
  assign n19449 = ~n19446 & n19448;
  assign n19450 = ~pi648 & ~n19290;
  assign n19451 = ~n19449 & n19450;
  assign n19452 = pi619 & ~n19445;
  assign n19453 = ~pi619 & n63424;
  assign n19454 = pi1159 & ~n19453;
  assign n19455 = ~n19452 & n19454;
  assign n19456 = pi648 & ~n19294;
  assign n19457 = ~n19455 & n19456;
  assign n19458 = pi789 & ~n19457;
  assign n19459 = pi789 & ~n19451;
  assign n19460 = ~n19457 & n19459;
  assign n19461 = ~n19451 & n19458;
  assign n19462 = ~pi789 & n19445;
  assign n19463 = n62894 & ~n19462;
  assign n19464 = ~n63436 & n19463;
  assign n19465 = n62894 & ~n19441;
  assign n19466 = ~pi626 & ~n63432;
  assign n19467 = pi626 & ~n19144;
  assign n19468 = n8301 & ~n19467;
  assign n19469 = ~n19466 & n19468;
  assign n19470 = n8525 & ~n63425;
  assign n19471 = pi626 & ~n63432;
  assign n19472 = ~pi626 & ~n19144;
  assign n19473 = n8300 & ~n19472;
  assign n19474 = ~n19471 & n19473;
  assign n19475 = ~n19470 & ~n19474;
  assign n19476 = ~n19469 & ~n19470;
  assign n19477 = ~n19474 & n19476;
  assign n19478 = ~n19469 & n19475;
  assign n19479 = pi788 & ~n63438;
  assign n19480 = ~n63030 & ~n19479;
  assign n19481 = ~n63437 & n19480;
  assign n19482 = ~n19338 & ~n19481;
  assign n19483 = ~n8651 & ~n19482;
  assign n19484 = ~n8413 & ~n19309;
  assign n19485 = ~n8413 & n19310;
  assign n19486 = ~n19308 & n19484;
  assign n19487 = n8373 & n63426;
  assign n19488 = ~pi630 & n63427;
  assign n19489 = n8374 & ~n19217;
  assign n19490 = pi630 & n19214;
  assign n19491 = ~n63440 & ~n63441;
  assign n19492 = ~n63439 & n19491;
  assign n19493 = pi787 & ~n19492;
  assign n19494 = ~pi644 & n19329;
  assign n19495 = pi644 & n19321;
  assign n19496 = n14029 & ~n19320;
  assign n19497 = pi790 & ~n63442;
  assign n19498 = pi790 & ~n19494;
  assign n19499 = ~n63442 & n19498;
  assign n19500 = ~n19494 & n19497;
  assign n19501 = ~n19493 & ~n63443;
  assign n19502 = ~n19483 & ~n19493;
  assign n19503 = ~n63443 & n19502;
  assign n19504 = ~n19483 & n19501;
  assign n19505 = ~n19332 & ~n63444;
  assign n19506 = n62455 & ~n19505;
  assign n19507 = ~pi184 & ~n62455;
  assign n19508 = ~pi832 & ~n19507;
  assign n19509 = ~n19506 & n19508;
  assign po341 = ~n19143 & ~n19509;
  assign n19511 = ~pi185 & ~n2923;
  assign n19512 = ~pi751 & n7316;
  assign n19513 = ~n19511 & ~n19512;
  assign n19514 = ~n8420 & ~n19513;
  assign n19515 = ~pi785 & ~n19514;
  assign n19516 = n8148 & n19512;
  assign n19517 = n19514 & ~n19516;
  assign n19518 = pi1155 & ~n19517;
  assign n19519 = ~pi1155 & ~n19511;
  assign n19520 = ~n19516 & n19519;
  assign n19521 = ~n19518 & ~n19520;
  assign n19522 = pi785 & ~n19521;
  assign n19523 = ~n19515 & ~n19522;
  assign n19524 = ~pi781 & ~n19523;
  assign n19525 = ~n8435 & n19523;
  assign n19526 = pi1154 & ~n19525;
  assign n19527 = ~n8438 & n19523;
  assign n19528 = ~pi1154 & ~n19527;
  assign n19529 = ~n19526 & ~n19528;
  assign n19530 = pi781 & ~n19529;
  assign n19531 = ~n19524 & ~n19530;
  assign n19532 = ~pi789 & ~n19531;
  assign n19533 = ~n12612 & n19531;
  assign n19534 = pi1159 & ~n19533;
  assign n19535 = ~n12615 & n19531;
  assign n19536 = ~pi1159 & ~n19535;
  assign n19537 = ~n19534 & ~n19536;
  assign n19538 = pi789 & ~n19537;
  assign n19539 = ~n19532 & ~n19538;
  assign n19540 = ~n15298 & n19531;
  assign n19541 = ~n8595 & n63445;
  assign n19542 = n8595 & n19511;
  assign n19543 = ~n8595 & ~n63445;
  assign n19544 = n8595 & ~n19511;
  assign n19545 = ~n19543 & ~n19544;
  assign n19546 = ~n19541 & ~n19542;
  assign n19547 = ~n8334 & n63446;
  assign n19548 = n8334 & n19511;
  assign n19549 = ~n8413 & ~n19548;
  assign n19550 = ~n19547 & ~n19548;
  assign n19551 = ~n8413 & n19550;
  assign n19552 = ~n19547 & n19549;
  assign n19553 = ~pi701 & n7564;
  assign n19554 = ~n19511 & ~n19553;
  assign n19555 = ~pi778 & ~n19554;
  assign n19556 = ~pi625 & n19553;
  assign n19557 = ~n19554 & ~n19556;
  assign n19558 = pi1153 & ~n19557;
  assign n19559 = ~pi1153 & ~n19511;
  assign n19560 = ~n19556 & n19559;
  assign n19561 = pi778 & ~n19560;
  assign n19562 = ~n19558 & n19561;
  assign n19563 = ~n19555 & ~n19562;
  assign n19564 = ~n8490 & ~n19563;
  assign n19565 = ~n8492 & n19564;
  assign n19566 = ~n8494 & n19565;
  assign n19567 = ~n8496 & n19566;
  assign n19568 = ~n8508 & n19567;
  assign n19569 = pi647 & ~n19568;
  assign n19570 = ~pi647 & ~n19511;
  assign n19571 = ~n19569 & ~n19570;
  assign n19572 = n8373 & ~n19571;
  assign n19573 = ~pi647 & n19568;
  assign n19574 = pi647 & n19511;
  assign n19575 = ~pi1157 & ~n19574;
  assign n19576 = ~n19573 & n19575;
  assign n19577 = pi630 & n19576;
  assign n19578 = ~n19572 & ~n19577;
  assign n19579 = ~n63447 & n19578;
  assign n19580 = pi787 & ~n19579;
  assign n19581 = ~pi626 & ~n63445;
  assign n19582 = pi626 & ~n19511;
  assign n19583 = n8301 & ~n19582;
  assign n19584 = ~n19581 & n19583;
  assign n19585 = n8525 & n19566;
  assign n19586 = pi626 & ~n63445;
  assign n19587 = ~pi626 & ~n19511;
  assign n19588 = n8300 & ~n19587;
  assign n19589 = ~n19586 & n19588;
  assign n19590 = ~n19585 & ~n19589;
  assign n19591 = ~n19584 & ~n19585;
  assign n19592 = ~n19589 & n19591;
  assign n19593 = ~n19584 & n19590;
  assign n19594 = pi788 & ~n63448;
  assign n19595 = n13460 & n19531;
  assign n19596 = n11303 & n19565;
  assign n19597 = pi648 & ~n19596;
  assign n19598 = ~n19595 & n19597;
  assign n19599 = n13462 & n19531;
  assign n19600 = n11304 & n19565;
  assign n19601 = ~pi648 & ~n19600;
  assign n19602 = ~n19599 & n19601;
  assign n19603 = pi789 & ~n19602;
  assign n19604 = ~n19598 & n19603;
  assign n19605 = ~n7187 & ~n19554;
  assign n19606 = pi625 & n19605;
  assign n19607 = n19513 & ~n19605;
  assign n19608 = ~n19606 & ~n19607;
  assign n19609 = n19559 & ~n19608;
  assign n19610 = ~pi608 & ~n19558;
  assign n19611 = ~n19609 & n19610;
  assign n19612 = pi1153 & n19513;
  assign n19613 = ~n19606 & n19612;
  assign n19614 = pi608 & ~n19560;
  assign n19615 = ~n19613 & n19614;
  assign n19616 = ~n19611 & ~n19615;
  assign n19617 = pi778 & ~n19616;
  assign n19618 = ~pi778 & ~n19607;
  assign n19619 = ~n19617 & ~n19618;
  assign n19620 = ~pi609 & ~n19619;
  assign n19621 = pi609 & ~n19563;
  assign n19622 = ~pi1155 & ~n19621;
  assign n19623 = ~n19620 & n19622;
  assign n19624 = ~pi660 & ~n19518;
  assign n19625 = ~n19623 & n19624;
  assign n19626 = pi609 & ~n19619;
  assign n19627 = ~pi609 & ~n19563;
  assign n19628 = pi1155 & ~n19627;
  assign n19629 = ~n19626 & n19628;
  assign n19630 = pi660 & ~n19520;
  assign n19631 = ~n19629 & n19630;
  assign n19632 = ~n19625 & ~n19631;
  assign n19633 = pi785 & ~n19632;
  assign n19634 = ~pi785 & ~n19619;
  assign n19635 = ~n19633 & ~n19634;
  assign n19636 = pi618 & ~n19635;
  assign n19637 = ~pi618 & n19564;
  assign n19638 = pi1154 & ~n19637;
  assign n19639 = ~n19636 & n19638;
  assign n19640 = pi627 & ~n19528;
  assign n19641 = ~n19639 & n19640;
  assign n19642 = ~pi618 & ~n19635;
  assign n19643 = pi618 & n19564;
  assign n19644 = ~pi1154 & ~n19643;
  assign n19645 = ~n19642 & n19644;
  assign n19646 = ~pi627 & ~n19526;
  assign n19647 = ~n19645 & n19646;
  assign n19648 = pi781 & ~n19647;
  assign n19649 = ~n19641 & n19648;
  assign n19650 = ~pi781 & n19635;
  assign n19651 = ~n11434 & ~n19650;
  assign n19652 = ~n19649 & n19651;
  assign n19653 = ~n19604 & ~n19652;
  assign n19654 = ~n19641 & ~n19647;
  assign n19655 = pi781 & ~n19654;
  assign n19656 = ~pi781 & ~n19635;
  assign n19657 = ~n19655 & ~n19656;
  assign n19658 = ~pi619 & ~n19657;
  assign n19659 = pi619 & n19565;
  assign n19660 = ~pi1159 & ~n19659;
  assign n19661 = ~n19658 & n19660;
  assign n19662 = ~pi648 & ~n19534;
  assign n19663 = ~n19661 & n19662;
  assign n19664 = pi619 & ~n19657;
  assign n19665 = ~pi619 & n19565;
  assign n19666 = pi1159 & ~n19665;
  assign n19667 = ~n19664 & n19666;
  assign n19668 = pi648 & ~n19536;
  assign n19669 = ~n19667 & n19668;
  assign n19670 = pi789 & ~n19669;
  assign n19671 = pi789 & ~n19663;
  assign n19672 = ~n19669 & n19671;
  assign n19673 = ~n19663 & n19670;
  assign n19674 = ~pi789 & n19657;
  assign n19675 = n62894 & ~n19674;
  assign n19676 = ~n63449 & n19675;
  assign n19677 = n62894 & ~n19653;
  assign n19678 = ~n19594 & ~n63450;
  assign n19679 = ~n63030 & ~n19678;
  assign n19680 = n8498 & n63446;
  assign n19681 = n8615 & n19567;
  assign n19682 = pi629 & ~n19681;
  assign n19683 = ~n19680 & n19682;
  assign n19684 = n8499 & n63446;
  assign n19685 = n8606 & n19567;
  assign n19686 = ~pi629 & ~n19685;
  assign n19687 = ~n19684 & n19686;
  assign n19688 = pi792 & ~n19687;
  assign n19689 = pi792 & ~n19683;
  assign n19690 = ~n19687 & n19689;
  assign n19691 = ~n19684 & ~n19685;
  assign n19692 = ~pi629 & ~n19691;
  assign n19693 = ~n19680 & ~n19681;
  assign n19694 = pi629 & ~n19693;
  assign n19695 = ~n19692 & ~n19694;
  assign n19696 = pi792 & ~n19695;
  assign n19697 = ~n19683 & n19688;
  assign n19698 = ~n8651 & ~n63451;
  assign n19699 = ~n19679 & n19698;
  assign n19700 = ~n19580 & ~n19699;
  assign n19701 = pi644 & n19700;
  assign n19702 = ~pi787 & ~n19568;
  assign n19703 = pi1157 & ~n19571;
  assign n19704 = ~n19576 & ~n19703;
  assign n19705 = pi787 & ~n19704;
  assign n19706 = ~n19702 & ~n19705;
  assign n19707 = ~pi644 & n19706;
  assign n19708 = pi715 & ~n19707;
  assign n19709 = ~n19701 & n19708;
  assign n19710 = ~n8685 & n19511;
  assign n19711 = ~n8376 & n19547;
  assign n19712 = ~n8376 & ~n19550;
  assign n19713 = n8376 & n19511;
  assign n19714 = ~n19712 & ~n19713;
  assign n19715 = ~n19710 & ~n19711;
  assign n19716 = pi644 & ~n63452;
  assign n19717 = ~pi644 & n19511;
  assign n19718 = ~pi715 & ~n19717;
  assign n19719 = ~n19716 & n19718;
  assign n19720 = pi1160 & ~n19719;
  assign n19721 = ~n19709 & n19720;
  assign n19722 = ~pi644 & n19700;
  assign n19723 = pi644 & n19706;
  assign n19724 = ~pi715 & ~n19723;
  assign n19725 = ~n19722 & n19724;
  assign n19726 = ~pi644 & ~n63452;
  assign n19727 = pi644 & n19511;
  assign n19728 = pi715 & ~n19727;
  assign n19729 = ~n19726 & n19728;
  assign n19730 = ~pi1160 & ~n19729;
  assign n19731 = ~n19725 & n19730;
  assign n19732 = ~n19721 & ~n19731;
  assign n19733 = pi790 & ~n19732;
  assign n19734 = ~pi790 & n19700;
  assign n19735 = pi832 & ~n19734;
  assign n19736 = ~n19733 & n19735;
  assign n19737 = ~pi185 & ~n8098;
  assign n19738 = n8257 & ~n19737;
  assign n19739 = ~pi701 & n62765;
  assign n19740 = n19737 & ~n19739;
  assign n19741 = pi185 & n62874;
  assign n19742 = ~pi38 & ~n19741;
  assign n19743 = n62765 & ~n19742;
  assign n19744 = ~pi185 & n8009;
  assign n19745 = ~n19743 & ~n19744;
  assign n19746 = ~pi185 & ~n7357;
  assign n19747 = n8085 & ~n19746;
  assign n19748 = ~pi701 & ~n19747;
  assign n19749 = ~n19745 & n19748;
  assign n19750 = ~n19740 & ~n19749;
  assign n19751 = ~pi778 & n19750;
  assign n19752 = pi625 & ~n19750;
  assign n19753 = ~pi625 & n19737;
  assign n19754 = pi1153 & ~n19753;
  assign n19755 = ~n19752 & n19754;
  assign n19756 = ~pi625 & ~n19750;
  assign n19757 = pi625 & n19737;
  assign n19758 = ~pi1153 & ~n19757;
  assign n19759 = ~n19756 & n19758;
  assign n19760 = ~n19755 & ~n19759;
  assign n19761 = pi778 & ~n19760;
  assign n19762 = ~n19751 & ~n19761;
  assign n19763 = ~n62880 & ~n19762;
  assign n19764 = n62880 & ~n19737;
  assign n19765 = ~n62880 & n19762;
  assign n19766 = n62880 & n19737;
  assign n19767 = ~n19765 & ~n19766;
  assign n19768 = ~n19763 & ~n19764;
  assign n19769 = ~n62882 & ~n63453;
  assign n19770 = n62882 & n19737;
  assign n19771 = n62882 & ~n19737;
  assign n19772 = ~n62882 & n63453;
  assign n19773 = ~n19771 & ~n19772;
  assign n19774 = ~n19769 & ~n19770;
  assign n19775 = ~n8257 & ~n63454;
  assign n19776 = ~n8257 & n63454;
  assign n19777 = n8257 & n19737;
  assign n19778 = ~n19776 & ~n19777;
  assign n19779 = ~n19738 & ~n19775;
  assign n19780 = ~n8303 & ~n63455;
  assign n19781 = n8303 & n19737;
  assign n19782 = ~n19780 & ~n19781;
  assign n19783 = ~pi792 & n19782;
  assign n19784 = pi628 & ~n19782;
  assign n19785 = ~pi628 & n19737;
  assign n19786 = pi1156 & ~n19785;
  assign n19787 = ~n19784 & n19786;
  assign n19788 = ~pi628 & ~n19782;
  assign n19789 = pi628 & n19737;
  assign n19790 = ~pi1156 & ~n19789;
  assign n19791 = ~n19788 & n19790;
  assign n19792 = ~n19787 & ~n19791;
  assign n19793 = pi792 & ~n19792;
  assign n19794 = ~n19783 & ~n19793;
  assign n19795 = pi647 & n19794;
  assign n19796 = ~pi647 & n19737;
  assign n19797 = pi1157 & ~n19796;
  assign n19798 = pi647 & ~n19794;
  assign n19799 = ~pi647 & ~n19737;
  assign n19800 = ~n19795 & ~n19796;
  assign n19801 = ~n19798 & ~n19799;
  assign n19802 = pi1157 & n63456;
  assign n19803 = ~n19795 & n19797;
  assign n19804 = ~pi647 & n19794;
  assign n19805 = pi647 & n19737;
  assign n19806 = ~pi1157 & ~n19805;
  assign n19807 = ~n19804 & n19806;
  assign n19808 = ~pi647 & ~n19794;
  assign n19809 = pi647 & ~n19737;
  assign n19810 = ~n19808 & ~n19809;
  assign n19811 = ~pi1157 & n19810;
  assign n19812 = pi1157 & ~n63456;
  assign n19813 = ~n19811 & ~n19812;
  assign n19814 = ~n63457 & ~n19807;
  assign n19815 = pi787 & n63458;
  assign n19816 = ~pi787 & ~n19794;
  assign n19817 = pi787 & ~n63458;
  assign n19818 = ~pi787 & n19794;
  assign n19819 = ~n19817 & ~n19818;
  assign n19820 = ~n19815 & ~n19816;
  assign n19821 = ~pi644 & ~n63459;
  assign n19822 = pi715 & ~n19821;
  assign n19823 = ~n11558 & n19737;
  assign n19824 = pi185 & ~n62765;
  assign n19825 = pi751 & n7143;
  assign n19826 = pi185 & n7349;
  assign n19827 = ~n19825 & ~n19826;
  assign n19828 = pi39 & ~n19827;
  assign n19829 = ~pi185 & ~pi751;
  assign n19830 = n62802 & n19829;
  assign n19831 = pi185 & pi751;
  assign n19832 = pi751 & ~n62781;
  assign n19833 = pi185 & ~n7292;
  assign n19834 = ~n19832 & ~n19833;
  assign n19835 = ~pi39 & ~n19834;
  assign n19836 = ~n19831 & ~n19835;
  assign n19837 = ~n19830 & n19836;
  assign n19838 = ~n19828 & n19837;
  assign n19839 = ~pi38 & ~n19838;
  assign n19840 = ~pi751 & n7359;
  assign n19841 = pi38 & ~n19746;
  assign n19842 = ~n19840 & n19841;
  assign n19843 = ~n19839 & ~n19842;
  assign n19844 = n62765 & ~n19843;
  assign n19845 = ~n19824 & ~n19844;
  assign n19846 = ~n8135 & ~n19845;
  assign n19847 = n8135 & ~n19737;
  assign n19848 = ~n19846 & ~n19847;
  assign n19849 = ~pi785 & ~n19848;
  assign n19850 = ~n8136 & ~n19737;
  assign n19851 = pi609 & n19846;
  assign n19852 = ~n19850 & ~n19851;
  assign n19853 = pi1155 & ~n19852;
  assign n19854 = ~n8148 & ~n19737;
  assign n19855 = ~pi609 & n19846;
  assign n19856 = ~n19854 & ~n19855;
  assign n19857 = ~pi1155 & ~n19856;
  assign n19858 = ~n19853 & ~n19857;
  assign n19859 = pi785 & ~n19858;
  assign n19860 = ~n19849 & ~n19859;
  assign n19861 = ~pi781 & ~n19860;
  assign n19862 = pi618 & n19860;
  assign n19863 = ~pi618 & n19737;
  assign n19864 = pi1154 & ~n19863;
  assign n19865 = ~n19862 & n19864;
  assign n19866 = ~pi618 & n19860;
  assign n19867 = pi618 & n19737;
  assign n19868 = ~pi1154 & ~n19867;
  assign n19869 = ~n19866 & n19868;
  assign n19870 = ~n19865 & ~n19869;
  assign n19871 = pi781 & ~n19870;
  assign n19872 = ~n19861 & ~n19871;
  assign n19873 = ~pi619 & ~n19872;
  assign n19874 = pi619 & ~n19737;
  assign n19875 = ~pi1159 & ~n19874;
  assign n19876 = ~n19873 & n19875;
  assign n19877 = pi619 & ~n19872;
  assign n19878 = ~pi619 & ~n19737;
  assign n19879 = pi1159 & ~n19878;
  assign n19880 = ~n19877 & n19879;
  assign n19881 = pi619 & n19872;
  assign n19882 = ~pi619 & n19737;
  assign n19883 = pi1159 & ~n19882;
  assign n19884 = ~n19881 & n19883;
  assign n19885 = ~pi619 & n19872;
  assign n19886 = pi619 & n19737;
  assign n19887 = ~pi1159 & ~n19886;
  assign n19888 = ~n19885 & n19887;
  assign n19889 = ~n19884 & ~n19888;
  assign n19890 = ~n19876 & ~n19880;
  assign n19891 = pi789 & n63460;
  assign n19892 = ~pi789 & n19872;
  assign n19893 = ~pi789 & ~n19872;
  assign n19894 = pi789 & ~n63460;
  assign n19895 = ~n19893 & ~n19894;
  assign n19896 = ~n19891 & ~n19892;
  assign n19897 = ~n8595 & n63461;
  assign n19898 = n8685 & n19897;
  assign n19899 = n8376 & ~n19737;
  assign n19900 = n8595 & n19737;
  assign n19901 = ~n19897 & ~n19900;
  assign n19902 = ~n8334 & ~n19901;
  assign n19903 = n8334 & n19737;
  assign n19904 = ~n19902 & ~n19903;
  assign n19905 = ~n8376 & n19904;
  assign n19906 = ~n19899 & ~n19905;
  assign n19907 = ~n8376 & ~n19904;
  assign n19908 = n8376 & n19737;
  assign n19909 = ~n19907 & ~n19908;
  assign n19910 = ~n19823 & ~n19898;
  assign n19911 = pi644 & n63462;
  assign n19912 = ~pi644 & n19737;
  assign n19913 = ~pi715 & ~n19912;
  assign n19914 = ~n19911 & n19913;
  assign n19915 = pi1160 & ~n19914;
  assign n19916 = ~n19822 & n19915;
  assign n19917 = pi644 & ~n63459;
  assign n19918 = ~pi715 & ~n19917;
  assign n19919 = ~pi644 & n63462;
  assign n19920 = pi644 & n19737;
  assign n19921 = pi715 & ~n19920;
  assign n19922 = ~n19919 & n19921;
  assign n19923 = ~pi1160 & ~n19922;
  assign n19924 = ~n19918 & n19923;
  assign n19925 = ~n19916 & ~n19924;
  assign n19926 = pi790 & ~n19925;
  assign n19927 = ~n63052 & n19901;
  assign n19928 = ~pi629 & n19787;
  assign n19929 = pi629 & n19791;
  assign n19930 = ~n19928 & ~n19929;
  assign n19931 = ~n19927 & n19930;
  assign n19932 = pi792 & ~n19931;
  assign n19933 = ~pi626 & ~n63461;
  assign n19934 = pi626 & ~n19737;
  assign n19935 = n8301 & ~n19934;
  assign n19936 = ~n19933 & n19935;
  assign n19937 = n8525 & ~n63455;
  assign n19938 = pi626 & ~n63461;
  assign n19939 = ~pi626 & ~n19737;
  assign n19940 = n8300 & ~n19939;
  assign n19941 = ~n19938 & n19940;
  assign n19942 = ~n19937 & ~n19941;
  assign n19943 = ~n19936 & ~n19937;
  assign n19944 = ~n19941 & n19943;
  assign n19945 = ~n19936 & n19942;
  assign n19946 = pi788 & ~n63463;
  assign n19947 = pi701 & n19843;
  assign n19948 = ~pi185 & ~n62821;
  assign n19949 = pi185 & n7632;
  assign n19950 = pi751 & ~n19949;
  assign n19951 = ~n19948 & n19950;
  assign n19952 = pi185 & n7709;
  assign n19953 = ~pi185 & n62851;
  assign n19954 = ~pi751 & ~n19953;
  assign n19955 = ~n19952 & n19954;
  assign n19956 = pi39 & ~n19955;
  assign n19957 = ~n19951 & n19956;
  assign n19958 = pi185 & n7855;
  assign n19959 = ~pi185 & n7832;
  assign n19960 = pi751 & ~n19959;
  assign n19961 = ~n19958 & n19960;
  assign n19962 = ~pi185 & ~n7861;
  assign n19963 = pi185 & ~n7868;
  assign n19964 = ~pi751 & ~n19963;
  assign n19965 = ~n19962 & n19964;
  assign n19966 = ~pi39 & ~n19965;
  assign n19967 = pi185 & ~n7855;
  assign n19968 = ~pi185 & ~n7832;
  assign n19969 = pi751 & ~n19968;
  assign n19970 = pi751 & ~n19967;
  assign n19971 = ~n19968 & n19970;
  assign n19972 = ~n19967 & n19969;
  assign n19973 = ~pi185 & n7861;
  assign n19974 = pi185 & n7868;
  assign n19975 = ~pi751 & ~n19974;
  assign n19976 = ~n19973 & n19975;
  assign n19977 = ~n63464 & ~n19976;
  assign n19978 = ~pi39 & ~n19977;
  assign n19979 = ~n19961 & n19966;
  assign n19980 = ~pi38 & ~n63465;
  assign n19981 = ~n19957 & n19980;
  assign n19982 = ~pi751 & ~n7744;
  assign n19983 = n10350 & ~n19982;
  assign n19984 = ~pi185 & ~n19983;
  assign n19985 = ~n7565 & ~n19512;
  assign n19986 = pi185 & ~n19985;
  assign n19987 = n7356 & n19986;
  assign n19988 = pi38 & ~n19987;
  assign n19989 = ~n19984 & n19988;
  assign n19990 = ~pi701 & ~n19989;
  assign n19991 = ~n19981 & n19990;
  assign n19992 = n62765 & ~n19991;
  assign n19993 = ~n19947 & n19992;
  assign n19994 = ~n19824 & ~n19993;
  assign n19995 = ~pi625 & n19994;
  assign n19996 = pi625 & n19845;
  assign n19997 = ~pi1153 & ~n19996;
  assign n19998 = ~n19995 & n19997;
  assign n19999 = ~pi608 & ~n19755;
  assign n20000 = ~n19998 & n19999;
  assign n20001 = pi625 & n19994;
  assign n20002 = ~pi625 & n19845;
  assign n20003 = pi1153 & ~n20002;
  assign n20004 = ~n20001 & n20003;
  assign n20005 = pi608 & ~n19759;
  assign n20006 = ~n20004 & n20005;
  assign n20007 = ~n20000 & ~n20006;
  assign n20008 = pi778 & ~n20007;
  assign n20009 = ~pi778 & n19994;
  assign n20010 = ~n20008 & ~n20009;
  assign n20011 = ~pi609 & ~n20010;
  assign n20012 = pi609 & n19762;
  assign n20013 = ~pi1155 & ~n20012;
  assign n20014 = ~n20011 & n20013;
  assign n20015 = ~pi660 & ~n19853;
  assign n20016 = ~n20014 & n20015;
  assign n20017 = pi609 & ~n20010;
  assign n20018 = ~pi609 & n19762;
  assign n20019 = pi1155 & ~n20018;
  assign n20020 = ~n20017 & n20019;
  assign n20021 = pi660 & ~n19857;
  assign n20022 = ~n20020 & n20021;
  assign n20023 = ~n20016 & ~n20022;
  assign n20024 = pi785 & ~n20023;
  assign n20025 = ~pi785 & ~n20010;
  assign n20026 = ~n20024 & ~n20025;
  assign n20027 = ~pi781 & n20026;
  assign n20028 = ~pi618 & ~n20026;
  assign n20029 = pi618 & ~n63453;
  assign n20030 = ~pi1154 & ~n20029;
  assign n20031 = ~n20028 & n20030;
  assign n20032 = ~pi627 & ~n19865;
  assign n20033 = ~n20031 & n20032;
  assign n20034 = pi618 & ~n20026;
  assign n20035 = ~pi618 & ~n63453;
  assign n20036 = pi1154 & ~n20035;
  assign n20037 = ~n20034 & n20036;
  assign n20038 = pi627 & ~n19869;
  assign n20039 = ~n20037 & n20038;
  assign n20040 = pi781 & ~n20039;
  assign n20041 = ~n20033 & n20040;
  assign n20042 = ~n20033 & ~n20039;
  assign n20043 = pi781 & ~n20042;
  assign n20044 = ~pi781 & ~n20026;
  assign n20045 = ~n20043 & ~n20044;
  assign n20046 = ~n20027 & ~n20041;
  assign n20047 = ~n11434 & n63466;
  assign n20048 = ~n11431 & ~n63454;
  assign n20049 = ~n62884 & ~n63460;
  assign n20050 = ~n20048 & ~n20049;
  assign n20051 = pi789 & ~n20050;
  assign n20052 = n62894 & ~n20051;
  assign n20053 = ~pi619 & ~n63466;
  assign n20054 = pi619 & n63454;
  assign n20055 = ~pi1159 & ~n20054;
  assign n20056 = ~n20053 & n20055;
  assign n20057 = ~pi648 & ~n19884;
  assign n20058 = ~n20056 & n20057;
  assign n20059 = pi619 & ~n63466;
  assign n20060 = ~pi619 & n63454;
  assign n20061 = pi1159 & ~n20060;
  assign n20062 = ~n20059 & n20061;
  assign n20063 = pi648 & ~n19888;
  assign n20064 = ~n20062 & n20063;
  assign n20065 = pi789 & ~n20064;
  assign n20066 = pi789 & ~n20058;
  assign n20067 = ~n20064 & n20066;
  assign n20068 = ~n20058 & n20065;
  assign n20069 = ~pi789 & n63466;
  assign n20070 = n62894 & ~n20069;
  assign n20071 = ~n63467 & n20070;
  assign n20072 = ~n20047 & n20052;
  assign n20073 = ~n63030 & ~n63468;
  assign n20074 = ~n63030 & ~n19946;
  assign n20075 = ~n63468 & n20074;
  assign n20076 = ~n19946 & n20073;
  assign n20077 = ~n19932 & ~n63469;
  assign n20078 = ~n8651 & ~n20077;
  assign n20079 = ~n8413 & ~n19903;
  assign n20080 = ~n8413 & n19904;
  assign n20081 = ~n19902 & n20079;
  assign n20082 = n8373 & n63456;
  assign n20083 = ~pi630 & n63457;
  assign n20084 = n8374 & ~n19810;
  assign n20085 = pi630 & n19807;
  assign n20086 = ~n63471 & ~n63472;
  assign n20087 = ~n63470 & n20086;
  assign n20088 = pi787 & ~n20087;
  assign n20089 = ~pi644 & n19923;
  assign n20090 = pi644 & n19915;
  assign n20091 = n14029 & ~n19914;
  assign n20092 = pi790 & ~n63473;
  assign n20093 = pi790 & ~n20089;
  assign n20094 = ~n63473 & n20093;
  assign n20095 = ~n20089 & n20092;
  assign n20096 = ~n20088 & ~n63474;
  assign n20097 = ~n20078 & ~n20088;
  assign n20098 = ~n63474 & n20097;
  assign n20099 = ~n20078 & n20096;
  assign n20100 = ~n19926 & ~n63475;
  assign n20101 = n62455 & ~n20100;
  assign n20102 = ~pi185 & ~n62455;
  assign n20103 = ~pi832 & ~n20102;
  assign n20104 = ~n20101 & n20103;
  assign po342 = ~n19736 & ~n20104;
  assign n20106 = ~pi186 & ~n2923;
  assign n20107 = ~pi752 & n7316;
  assign n20108 = ~n20106 & ~n20107;
  assign n20109 = ~n8420 & ~n20108;
  assign n20110 = ~pi785 & ~n20109;
  assign n20111 = ~n8425 & ~n20108;
  assign n20112 = pi1155 & ~n20111;
  assign n20113 = ~n8428 & n20109;
  assign n20114 = ~pi1155 & ~n20113;
  assign n20115 = ~n20112 & ~n20114;
  assign n20116 = pi785 & ~n20115;
  assign n20117 = ~n20110 & ~n20116;
  assign n20118 = ~pi781 & ~n20117;
  assign n20119 = ~n8435 & n20117;
  assign n20120 = pi1154 & ~n20119;
  assign n20121 = ~n8438 & n20117;
  assign n20122 = ~pi1154 & ~n20121;
  assign n20123 = ~n20120 & ~n20122;
  assign n20124 = pi781 & ~n20123;
  assign n20125 = ~n20118 & ~n20124;
  assign n20126 = ~pi619 & ~n20125;
  assign n20127 = pi619 & ~n20106;
  assign n20128 = ~pi1159 & ~n20127;
  assign n20129 = ~n20126 & n20128;
  assign n20130 = pi619 & ~n20125;
  assign n20131 = ~pi619 & ~n20106;
  assign n20132 = pi1159 & ~n20131;
  assign n20133 = ~n20130 & n20132;
  assign n20134 = pi619 & n20125;
  assign n20135 = ~pi619 & n20106;
  assign n20136 = pi1159 & ~n20135;
  assign n20137 = ~n20134 & n20136;
  assign n20138 = ~pi619 & n20125;
  assign n20139 = pi619 & n20106;
  assign n20140 = ~pi1159 & ~n20139;
  assign n20141 = ~n20138 & n20140;
  assign n20142 = ~n20137 & ~n20141;
  assign n20143 = ~n20129 & ~n20133;
  assign n20144 = pi789 & n63476;
  assign n20145 = ~pi789 & n20125;
  assign n20146 = ~pi789 & ~n20125;
  assign n20147 = pi789 & ~n63476;
  assign n20148 = ~n20146 & ~n20147;
  assign n20149 = ~n20144 & ~n20145;
  assign n20150 = ~n8595 & n63477;
  assign n20151 = n8595 & n20106;
  assign n20152 = ~n8595 & ~n63477;
  assign n20153 = n8595 & ~n20106;
  assign n20154 = ~n20152 & ~n20153;
  assign n20155 = ~n20150 & ~n20151;
  assign n20156 = ~n8334 & n63478;
  assign n20157 = n8334 & n20106;
  assign n20158 = ~n8413 & ~n20157;
  assign n20159 = ~n20156 & ~n20157;
  assign n20160 = ~n8413 & n20159;
  assign n20161 = ~n20156 & n20158;
  assign n20162 = pi703 & n7564;
  assign n20163 = ~n20106 & ~n20162;
  assign n20164 = ~pi778 & n20163;
  assign n20165 = ~pi625 & n20162;
  assign n20166 = ~n20163 & ~n20165;
  assign n20167 = pi1153 & ~n20166;
  assign n20168 = ~pi1153 & ~n20106;
  assign n20169 = ~n20165 & n20168;
  assign n20170 = ~n20167 & ~n20169;
  assign n20171 = pi778 & ~n20170;
  assign n20172 = ~n20164 & ~n20171;
  assign n20173 = ~n8490 & n20172;
  assign n20174 = ~n8492 & n20173;
  assign n20175 = ~n8494 & n20174;
  assign n20176 = ~n8496 & n20175;
  assign n20177 = ~n8508 & n20176;
  assign n20178 = pi647 & ~n20177;
  assign n20179 = ~pi647 & ~n20106;
  assign n20180 = ~n20178 & ~n20179;
  assign n20181 = n8373 & ~n20180;
  assign n20182 = ~pi647 & n20177;
  assign n20183 = pi647 & n20106;
  assign n20184 = ~pi1157 & ~n20183;
  assign n20185 = ~n20182 & n20184;
  assign n20186 = pi630 & n20185;
  assign n20187 = ~n20181 & ~n20186;
  assign n20188 = ~n63479 & n20187;
  assign n20189 = pi787 & ~n20188;
  assign n20190 = ~pi626 & ~n63477;
  assign n20191 = pi626 & ~n20106;
  assign n20192 = n8301 & ~n20191;
  assign n20193 = ~n20190 & n20192;
  assign n20194 = n8525 & n20175;
  assign n20195 = pi626 & ~n63477;
  assign n20196 = ~pi626 & ~n20106;
  assign n20197 = n8300 & ~n20196;
  assign n20198 = ~n20195 & n20197;
  assign n20199 = ~n20194 & ~n20198;
  assign n20200 = ~n20193 & ~n20194;
  assign n20201 = ~n20198 & n20200;
  assign n20202 = ~n20193 & n20199;
  assign n20203 = pi788 & ~n63480;
  assign n20204 = ~n7187 & ~n20163;
  assign n20205 = pi625 & n20204;
  assign n20206 = n20108 & ~n20204;
  assign n20207 = ~n20205 & ~n20206;
  assign n20208 = n20168 & ~n20207;
  assign n20209 = ~pi608 & ~n20167;
  assign n20210 = ~n20208 & n20209;
  assign n20211 = pi1153 & n20108;
  assign n20212 = ~n20205 & n20211;
  assign n20213 = pi608 & ~n20169;
  assign n20214 = ~n20212 & n20213;
  assign n20215 = ~n20210 & ~n20214;
  assign n20216 = pi778 & ~n20215;
  assign n20217 = ~pi778 & ~n20206;
  assign n20218 = ~n20216 & ~n20217;
  assign n20219 = ~pi609 & ~n20218;
  assign n20220 = pi609 & n20172;
  assign n20221 = ~pi1155 & ~n20220;
  assign n20222 = ~n20219 & n20221;
  assign n20223 = ~pi660 & ~n20112;
  assign n20224 = ~n20222 & n20223;
  assign n20225 = pi609 & ~n20218;
  assign n20226 = ~pi609 & n20172;
  assign n20227 = pi1155 & ~n20226;
  assign n20228 = ~n20225 & n20227;
  assign n20229 = pi660 & ~n20114;
  assign n20230 = ~n20228 & n20229;
  assign n20231 = ~n20224 & ~n20230;
  assign n20232 = pi785 & ~n20231;
  assign n20233 = ~pi785 & ~n20218;
  assign n20234 = ~n20232 & ~n20233;
  assign n20235 = pi618 & ~n20234;
  assign n20236 = ~pi618 & n20173;
  assign n20237 = pi1154 & ~n20236;
  assign n20238 = ~n20235 & n20237;
  assign n20239 = pi627 & ~n20122;
  assign n20240 = ~n20238 & n20239;
  assign n20241 = ~pi618 & ~n20234;
  assign n20242 = pi618 & n20173;
  assign n20243 = ~pi1154 & ~n20242;
  assign n20244 = ~n20241 & n20243;
  assign n20245 = ~pi627 & ~n20120;
  assign n20246 = ~n20244 & n20245;
  assign n20247 = pi781 & ~n20246;
  assign n20248 = ~n20240 & n20247;
  assign n20249 = ~n11431 & ~n20174;
  assign n20250 = ~n62884 & ~n63476;
  assign n20251 = ~n20249 & ~n20250;
  assign n20252 = pi789 & ~n20251;
  assign n20253 = ~pi781 & n20234;
  assign n20254 = ~n20252 & ~n20253;
  assign n20255 = ~n20248 & n20254;
  assign n20256 = n11434 & n20251;
  assign n20257 = ~n20255 & ~n20256;
  assign n20258 = ~n20240 & ~n20246;
  assign n20259 = pi781 & ~n20258;
  assign n20260 = ~pi781 & ~n20234;
  assign n20261 = ~n20259 & ~n20260;
  assign n20262 = ~pi619 & ~n20261;
  assign n20263 = pi619 & n20174;
  assign n20264 = ~pi1159 & ~n20263;
  assign n20265 = ~n20262 & n20264;
  assign n20266 = ~pi648 & ~n20137;
  assign n20267 = ~n20265 & n20266;
  assign n20268 = pi619 & ~n20261;
  assign n20269 = ~pi619 & n20174;
  assign n20270 = pi1159 & ~n20269;
  assign n20271 = ~n20268 & n20270;
  assign n20272 = pi648 & ~n20141;
  assign n20273 = ~n20271 & n20272;
  assign n20274 = pi789 & ~n20273;
  assign n20275 = pi789 & ~n20267;
  assign n20276 = ~n20273 & n20275;
  assign n20277 = ~n20267 & n20274;
  assign n20278 = ~pi789 & n20261;
  assign n20279 = n62894 & ~n20278;
  assign n20280 = ~n63481 & n20279;
  assign n20281 = n62894 & ~n20257;
  assign n20282 = ~n20203 & ~n63482;
  assign n20283 = ~n63030 & ~n20282;
  assign n20284 = n8498 & n63478;
  assign n20285 = n8615 & n20176;
  assign n20286 = pi629 & ~n20285;
  assign n20287 = ~n20284 & n20286;
  assign n20288 = n8499 & n63478;
  assign n20289 = n8606 & n20176;
  assign n20290 = ~pi629 & ~n20289;
  assign n20291 = ~n20288 & n20290;
  assign n20292 = pi792 & ~n20291;
  assign n20293 = pi792 & ~n20287;
  assign n20294 = ~n20291 & n20293;
  assign n20295 = ~n20288 & ~n20289;
  assign n20296 = ~pi629 & ~n20295;
  assign n20297 = ~n20284 & ~n20285;
  assign n20298 = pi629 & ~n20297;
  assign n20299 = ~n20296 & ~n20298;
  assign n20300 = pi792 & ~n20299;
  assign n20301 = ~n20287 & n20292;
  assign n20302 = ~n8651 & ~n63483;
  assign n20303 = ~n20283 & n20302;
  assign n20304 = ~n20189 & ~n20303;
  assign n20305 = pi644 & n20304;
  assign n20306 = ~pi787 & ~n20177;
  assign n20307 = pi1157 & ~n20180;
  assign n20308 = ~n20185 & ~n20307;
  assign n20309 = pi787 & ~n20308;
  assign n20310 = ~n20306 & ~n20309;
  assign n20311 = ~pi644 & n20310;
  assign n20312 = pi715 & ~n20311;
  assign n20313 = ~n20305 & n20312;
  assign n20314 = ~n8685 & n20106;
  assign n20315 = ~n8376 & n20156;
  assign n20316 = ~n8376 & ~n20159;
  assign n20317 = n8376 & n20106;
  assign n20318 = ~n20316 & ~n20317;
  assign n20319 = ~n20314 & ~n20315;
  assign n20320 = pi644 & ~n63484;
  assign n20321 = ~pi644 & n20106;
  assign n20322 = ~pi715 & ~n20321;
  assign n20323 = ~n20320 & n20322;
  assign n20324 = pi1160 & ~n20323;
  assign n20325 = ~n20313 & n20324;
  assign n20326 = ~pi644 & n20304;
  assign n20327 = pi644 & n20310;
  assign n20328 = ~pi715 & ~n20327;
  assign n20329 = ~n20326 & n20328;
  assign n20330 = ~pi644 & ~n63484;
  assign n20331 = pi644 & n20106;
  assign n20332 = pi715 & ~n20331;
  assign n20333 = ~n20330 & n20332;
  assign n20334 = ~pi1160 & ~n20333;
  assign n20335 = ~n20329 & n20334;
  assign n20336 = ~n20325 & ~n20335;
  assign n20337 = pi790 & ~n20336;
  assign n20338 = ~pi790 & n20304;
  assign n20339 = pi832 & ~n20338;
  assign n20340 = ~n20337 & n20339;
  assign n20341 = pi186 & ~n62765;
  assign n20342 = ~pi186 & ~n8091;
  assign n20343 = pi752 & ~n20342;
  assign n20344 = pi186 & ~n10339;
  assign n20345 = ~pi186 & ~pi752;
  assign n20346 = n10343 & n20345;
  assign n20347 = ~n20344 & ~n20346;
  assign n20348 = ~n62977 & ~n20347;
  assign n20349 = ~n20343 & ~n20348;
  assign n20350 = n62765 & ~n20349;
  assign n20351 = ~n20341 & ~n20350;
  assign n20352 = ~n8135 & ~n20351;
  assign n20353 = ~pi186 & ~n8098;
  assign n20354 = n8135 & ~n20353;
  assign n20355 = ~n20352 & ~n20354;
  assign n20356 = ~pi785 & ~n20355;
  assign n20357 = ~n8136 & ~n20353;
  assign n20358 = pi609 & n20352;
  assign n20359 = ~n20357 & ~n20358;
  assign n20360 = pi1155 & ~n20359;
  assign n20361 = ~n8148 & ~n20353;
  assign n20362 = ~pi609 & n20352;
  assign n20363 = ~n20361 & ~n20362;
  assign n20364 = ~pi1155 & ~n20363;
  assign n20365 = ~n20360 & ~n20364;
  assign n20366 = pi785 & ~n20365;
  assign n20367 = ~n20356 & ~n20366;
  assign n20368 = ~pi781 & ~n20367;
  assign n20369 = pi618 & n20367;
  assign n20370 = ~pi618 & n20353;
  assign n20371 = pi1154 & ~n20370;
  assign n20372 = ~n20369 & n20371;
  assign n20373 = ~pi618 & n20367;
  assign n20374 = pi618 & n20353;
  assign n20375 = ~pi1154 & ~n20374;
  assign n20376 = ~n20373 & n20375;
  assign n20377 = ~n20372 & ~n20376;
  assign n20378 = pi781 & ~n20377;
  assign n20379 = ~n20368 & ~n20378;
  assign n20380 = ~pi789 & ~n20379;
  assign n20381 = ~pi619 & n20379;
  assign n20382 = pi619 & n20353;
  assign n20383 = ~pi1159 & ~n20382;
  assign n20384 = ~n20381 & n20383;
  assign n20385 = pi619 & n20379;
  assign n20386 = ~pi619 & n20353;
  assign n20387 = pi1159 & ~n20386;
  assign n20388 = ~n20385 & n20387;
  assign n20389 = ~n20384 & ~n20388;
  assign n20390 = pi789 & ~n20389;
  assign n20391 = ~n20380 & ~n20390;
  assign n20392 = ~n8595 & n20391;
  assign n20393 = n8595 & n20353;
  assign n20394 = ~n20392 & ~n20393;
  assign n20395 = ~n8334 & ~n20394;
  assign n20396 = n8334 & n20353;
  assign n20397 = ~n20395 & ~n20396;
  assign n20398 = ~n8376 & ~n20397;
  assign n20399 = n8376 & n20353;
  assign n20400 = n8376 & ~n20353;
  assign n20401 = ~n8376 & n20397;
  assign n20402 = ~n20400 & ~n20401;
  assign n20403 = ~n20398 & ~n20399;
  assign n20404 = ~pi644 & n63485;
  assign n20405 = pi644 & n20353;
  assign n20406 = n16172 & ~n20405;
  assign n20407 = ~n20404 & n20406;
  assign n20408 = pi644 & n63485;
  assign n20409 = ~pi644 & n20353;
  assign n20410 = n16177 & ~n20409;
  assign n20411 = ~n20408 & n20410;
  assign n20412 = n8257 & ~n20353;
  assign n20413 = ~pi186 & n8009;
  assign n20414 = pi186 & n62874;
  assign n20415 = ~pi38 & ~n20414;
  assign n20416 = ~n20413 & n20415;
  assign n20417 = ~pi186 & ~n7357;
  assign n20418 = n8085 & ~n20417;
  assign n20419 = pi703 & ~n20418;
  assign n20420 = ~n20416 & n20419;
  assign n20421 = ~pi703 & n20342;
  assign n20422 = n62765 & ~n20421;
  assign n20423 = n62765 & ~n20420;
  assign n20424 = ~n20421 & n20423;
  assign n20425 = ~n20420 & n20422;
  assign n20426 = ~n20341 & ~n63486;
  assign n20427 = ~pi778 & ~n20426;
  assign n20428 = pi625 & n20426;
  assign n20429 = ~pi625 & n20353;
  assign n20430 = pi1153 & ~n20429;
  assign n20431 = ~n20428 & n20430;
  assign n20432 = ~pi625 & n20426;
  assign n20433 = pi625 & n20353;
  assign n20434 = ~pi1153 & ~n20433;
  assign n20435 = ~n20432 & n20434;
  assign n20436 = ~n20431 & ~n20435;
  assign n20437 = pi778 & ~n20436;
  assign n20438 = ~n20427 & ~n20437;
  assign n20439 = ~n62880 & ~n20438;
  assign n20440 = n62880 & ~n20353;
  assign n20441 = ~n62880 & n20438;
  assign n20442 = n62880 & n20353;
  assign n20443 = ~n20441 & ~n20442;
  assign n20444 = ~n20439 & ~n20440;
  assign n20445 = ~n62882 & ~n63487;
  assign n20446 = n62882 & n20353;
  assign n20447 = n62882 & ~n20353;
  assign n20448 = ~n62882 & n63487;
  assign n20449 = ~n20447 & ~n20448;
  assign n20450 = ~n20445 & ~n20446;
  assign n20451 = ~n8257 & ~n63488;
  assign n20452 = ~n8257 & n63488;
  assign n20453 = n8257 & n20353;
  assign n20454 = ~n20452 & ~n20453;
  assign n20455 = ~n20412 & ~n20451;
  assign n20456 = ~n8303 & ~n63489;
  assign n20457 = n8303 & n20353;
  assign n20458 = n8303 & ~n20353;
  assign n20459 = ~n8303 & n63489;
  assign n20460 = ~n20458 & ~n20459;
  assign n20461 = ~n20456 & ~n20457;
  assign n20462 = ~pi792 & ~n63490;
  assign n20463 = pi628 & n63490;
  assign n20464 = ~pi628 & n20353;
  assign n20465 = pi1156 & ~n20464;
  assign n20466 = ~pi628 & ~n20353;
  assign n20467 = pi628 & ~n63490;
  assign n20468 = ~n20466 & ~n20467;
  assign n20469 = pi1156 & ~n20468;
  assign n20470 = ~n20463 & n20465;
  assign n20471 = ~pi628 & n63490;
  assign n20472 = pi628 & n20353;
  assign n20473 = ~pi1156 & ~n20472;
  assign n20474 = ~n20471 & n20473;
  assign n20475 = ~n63491 & ~n20474;
  assign n20476 = pi792 & ~n20475;
  assign n20477 = ~n20462 & ~n20476;
  assign n20478 = pi647 & n20477;
  assign n20479 = ~pi647 & n20353;
  assign n20480 = pi1157 & ~n20479;
  assign n20481 = ~pi647 & ~n20353;
  assign n20482 = pi647 & ~n20477;
  assign n20483 = ~n20481 & ~n20482;
  assign n20484 = ~n20478 & ~n20479;
  assign n20485 = pi1157 & ~n63492;
  assign n20486 = ~n20478 & n20480;
  assign n20487 = ~pi647 & n20477;
  assign n20488 = pi647 & n20353;
  assign n20489 = ~pi1157 & ~n20488;
  assign n20490 = ~n20487 & n20489;
  assign n20491 = pi787 & ~n20490;
  assign n20492 = ~n63493 & n20491;
  assign n20493 = ~pi787 & n20477;
  assign n20494 = ~n63036 & ~n20493;
  assign n20495 = ~n20492 & n20494;
  assign n20496 = ~n20411 & ~n20495;
  assign n20497 = ~n20407 & n20496;
  assign n20498 = pi790 & ~n20497;
  assign n20499 = ~n63052 & n20394;
  assign n20500 = n8331 & ~n20468;
  assign n20501 = ~pi629 & n63491;
  assign n20502 = pi629 & n20474;
  assign n20503 = ~n63494 & ~n20502;
  assign n20504 = ~n20499 & n20503;
  assign n20505 = pi792 & ~n20504;
  assign n20506 = n12979 & n20391;
  assign n20507 = ~pi641 & n63489;
  assign n20508 = pi641 & ~n20353;
  assign n20509 = n8417 & ~n20508;
  assign n20510 = ~n20507 & n20509;
  assign n20511 = pi641 & n63489;
  assign n20512 = ~pi641 & ~n20353;
  assign n20513 = n8416 & ~n20512;
  assign n20514 = ~n20511 & n20513;
  assign n20515 = ~n20510 & ~n20514;
  assign n20516 = ~n20506 & n20515;
  assign n20517 = pi788 & ~n20516;
  assign n20518 = pi619 & n63488;
  assign n20519 = ~pi1159 & ~n20518;
  assign n20520 = ~pi648 & ~n20388;
  assign n20521 = ~n20519 & n20520;
  assign n20522 = ~pi619 & n63488;
  assign n20523 = pi1159 & ~n20522;
  assign n20524 = pi648 & ~n20523;
  assign n20525 = pi648 & ~n20384;
  assign n20526 = ~n20523 & n20525;
  assign n20527 = ~n20384 & n20524;
  assign n20528 = ~n20521 & ~n63495;
  assign n20529 = pi789 & ~n20528;
  assign n20530 = pi618 & ~n63487;
  assign n20531 = ~pi1154 & ~n20530;
  assign n20532 = ~pi627 & ~n20372;
  assign n20533 = ~n20531 & n20532;
  assign n20534 = ~pi618 & ~n63487;
  assign n20535 = pi1154 & ~n20534;
  assign n20536 = pi627 & ~n20376;
  assign n20537 = ~n20535 & n20536;
  assign n20538 = ~n20533 & ~n20537;
  assign n20539 = pi781 & ~n20538;
  assign n20540 = ~pi618 & n20532;
  assign n20541 = pi618 & n20536;
  assign n20542 = pi781 & ~n20541;
  assign n20543 = ~n20540 & n20542;
  assign n20544 = ~pi703 & n20349;
  assign n20545 = ~pi186 & n10353;
  assign n20546 = pi186 & n10355;
  assign n20547 = pi752 & ~n10357;
  assign n20548 = ~n20546 & n20547;
  assign n20549 = ~n20545 & n20548;
  assign n20550 = pi186 & n10363;
  assign n20551 = ~pi186 & ~n62980;
  assign n20552 = ~pi752 & ~n20551;
  assign n20553 = ~n20550 & n20552;
  assign n20554 = pi703 & ~n20553;
  assign n20555 = ~n20549 & n20554;
  assign n20556 = n62765 & ~n20555;
  assign n20557 = n62765 & ~n20544;
  assign n20558 = ~n20555 & n20557;
  assign n20559 = ~n20544 & n20556;
  assign n20560 = ~n20341 & ~n63496;
  assign n20561 = ~pi625 & n20560;
  assign n20562 = pi625 & n20351;
  assign n20563 = ~pi1153 & ~n20562;
  assign n20564 = ~n20561 & n20563;
  assign n20565 = ~pi608 & ~n20431;
  assign n20566 = ~n20564 & n20565;
  assign n20567 = pi625 & n20560;
  assign n20568 = ~pi625 & n20351;
  assign n20569 = pi1153 & ~n20568;
  assign n20570 = ~n20567 & n20569;
  assign n20571 = pi608 & ~n20435;
  assign n20572 = ~n20570 & n20571;
  assign n20573 = ~n20566 & ~n20572;
  assign n20574 = pi778 & ~n20573;
  assign n20575 = ~pi778 & n20560;
  assign n20576 = ~pi778 & ~n20560;
  assign n20577 = pi778 & ~n20572;
  assign n20578 = ~n20566 & n20577;
  assign n20579 = ~n20576 & ~n20578;
  assign n20580 = ~n20574 & ~n20575;
  assign n20581 = ~pi609 & n63497;
  assign n20582 = pi609 & n20438;
  assign n20583 = ~pi1155 & ~n20582;
  assign n20584 = ~n20581 & n20583;
  assign n20585 = ~pi660 & ~n20360;
  assign n20586 = ~n20584 & n20585;
  assign n20587 = pi609 & n63497;
  assign n20588 = ~pi609 & n20438;
  assign n20589 = pi1155 & ~n20588;
  assign n20590 = ~n20587 & n20589;
  assign n20591 = pi660 & ~n20364;
  assign n20592 = ~n20590 & n20591;
  assign n20593 = pi785 & ~n20592;
  assign n20594 = ~n20586 & n20593;
  assign n20595 = ~pi785 & ~n63497;
  assign n20596 = ~n20586 & ~n20592;
  assign n20597 = pi785 & ~n20596;
  assign n20598 = ~pi785 & n63497;
  assign n20599 = ~n20597 & ~n20598;
  assign n20600 = ~n20594 & ~n20595;
  assign n20601 = ~n20543 & ~n63498;
  assign n20602 = pi618 & ~n63498;
  assign n20603 = n20535 & ~n20602;
  assign n20604 = n20536 & ~n20603;
  assign n20605 = ~n20533 & ~n20604;
  assign n20606 = pi781 & ~n20605;
  assign n20607 = pi781 & ~n20540;
  assign n20608 = ~n63498 & ~n20607;
  assign n20609 = ~n20606 & ~n20608;
  assign n20610 = ~pi618 & ~n63498;
  assign n20611 = n20531 & ~n20610;
  assign n20612 = n20532 & ~n20611;
  assign n20613 = ~n20604 & ~n20612;
  assign n20614 = pi781 & ~n20613;
  assign n20615 = ~pi781 & ~n63498;
  assign n20616 = ~n20614 & ~n20615;
  assign n20617 = ~n20539 & ~n20601;
  assign n20618 = ~pi619 & n20520;
  assign n20619 = pi619 & n20525;
  assign n20620 = n11422 & ~n20384;
  assign n20621 = pi789 & ~n63500;
  assign n20622 = ~n20618 & n20621;
  assign n20623 = ~n63499 & ~n20622;
  assign n20624 = ~pi619 & ~n63499;
  assign n20625 = n20519 & ~n20624;
  assign n20626 = n20520 & ~n20625;
  assign n20627 = pi619 & ~n63499;
  assign n20628 = n20523 & ~n20627;
  assign n20629 = n20525 & ~n20628;
  assign n20630 = ~n20626 & ~n20629;
  assign n20631 = pi789 & ~n20630;
  assign n20632 = ~pi789 & ~n63499;
  assign n20633 = ~n20631 & ~n20632;
  assign n20634 = ~n20529 & ~n20623;
  assign n20635 = n62894 & ~n63501;
  assign n20636 = ~n63030 & ~n20635;
  assign n20637 = ~n63030 & ~n20517;
  assign n20638 = ~n20635 & n20637;
  assign n20639 = ~n20517 & n20636;
  assign n20640 = ~pi788 & n63501;
  assign n20641 = ~pi626 & n63501;
  assign n20642 = pi626 & n63489;
  assign n20643 = ~pi641 & ~n20642;
  assign n20644 = ~n20641 & n20643;
  assign n20645 = ~pi626 & ~n20391;
  assign n20646 = pi626 & ~n20353;
  assign n20647 = pi641 & ~n20646;
  assign n20648 = ~n20645 & n20647;
  assign n20649 = ~pi1158 & ~n20648;
  assign n20650 = ~n20644 & n20649;
  assign n20651 = pi626 & n63501;
  assign n20652 = ~pi626 & n63489;
  assign n20653 = pi641 & ~n20652;
  assign n20654 = ~n20651 & n20653;
  assign n20655 = pi626 & ~n20391;
  assign n20656 = ~pi626 & ~n20353;
  assign n20657 = ~pi641 & ~n20656;
  assign n20658 = ~n20655 & n20657;
  assign n20659 = pi1158 & ~n20658;
  assign n20660 = ~n20654 & n20659;
  assign n20661 = ~n20650 & ~n20660;
  assign n20662 = pi788 & ~n20661;
  assign n20663 = ~n20640 & ~n20662;
  assign n20664 = ~pi628 & n20663;
  assign n20665 = pi628 & ~n20394;
  assign n20666 = ~pi1156 & ~n20665;
  assign n20667 = ~n20664 & n20666;
  assign n20668 = ~pi629 & ~n63491;
  assign n20669 = ~n20667 & n20668;
  assign n20670 = pi628 & n20663;
  assign n20671 = ~pi628 & ~n20394;
  assign n20672 = pi1156 & ~n20671;
  assign n20673 = ~n20670 & n20672;
  assign n20674 = pi629 & ~n20474;
  assign n20675 = ~n20673 & n20674;
  assign n20676 = ~n20669 & ~n20675;
  assign n20677 = pi792 & ~n20676;
  assign n20678 = ~pi792 & n20663;
  assign n20679 = ~n20677 & ~n20678;
  assign n20680 = ~n20505 & ~n63502;
  assign n20681 = ~n8651 & n63503;
  assign n20682 = ~n8413 & n20397;
  assign n20683 = n8373 & ~n63492;
  assign n20684 = pi630 & n20490;
  assign n20685 = ~n20683 & ~n20684;
  assign n20686 = ~n20682 & ~n20684;
  assign n20687 = ~n20683 & n20686;
  assign n20688 = ~n20682 & n20685;
  assign n20689 = pi787 & ~n63504;
  assign n20690 = ~n62896 & n63503;
  assign n20691 = ~pi647 & ~n63503;
  assign n20692 = pi647 & ~n20397;
  assign n20693 = ~pi1157 & ~n20692;
  assign n20694 = ~n20691 & n20693;
  assign n20695 = ~pi630 & ~n63493;
  assign n20696 = ~n20694 & n20695;
  assign n20697 = pi647 & ~n63503;
  assign n20698 = ~pi647 & ~n20397;
  assign n20699 = pi1157 & ~n20698;
  assign n20700 = ~n20697 & n20699;
  assign n20701 = pi630 & ~n20490;
  assign n20702 = ~n20700 & n20701;
  assign n20703 = ~n20696 & ~n20702;
  assign n20704 = n63504 & ~n20690;
  assign n20705 = pi787 & n63505;
  assign n20706 = ~pi787 & n63503;
  assign n20707 = ~n20705 & ~n20706;
  assign n20708 = pi787 & ~n63505;
  assign n20709 = ~pi787 & ~n63503;
  assign n20710 = ~n20708 & ~n20709;
  assign n20711 = ~n20681 & ~n20689;
  assign n20712 = ~n11547 & ~n63506;
  assign n20713 = n62455 & ~n20712;
  assign n20714 = ~pi644 & n63506;
  assign n20715 = ~pi787 & ~n20477;
  assign n20716 = ~n63493 & ~n20490;
  assign n20717 = pi787 & ~n20716;
  assign n20718 = ~n20715 & ~n20717;
  assign n20719 = pi644 & n20718;
  assign n20720 = ~pi715 & ~n20719;
  assign n20721 = ~n20714 & n20720;
  assign n20722 = pi715 & ~n20405;
  assign n20723 = ~n20404 & n20722;
  assign n20724 = ~pi1160 & ~n20723;
  assign n20725 = ~n20721 & n20724;
  assign n20726 = ~pi644 & n20718;
  assign n20727 = pi715 & ~n20726;
  assign n20728 = ~pi715 & ~n20409;
  assign n20729 = ~n20408 & n20728;
  assign n20730 = pi1160 & ~n20729;
  assign n20731 = ~n20727 & n20730;
  assign n20732 = ~n20725 & ~n20731;
  assign n20733 = pi790 & ~n20732;
  assign n20734 = pi644 & n20730;
  assign n20735 = pi790 & ~n20734;
  assign n20736 = n63506 & ~n20735;
  assign n20737 = ~n20733 & ~n20736;
  assign n20738 = n62455 & ~n20737;
  assign n20739 = pi644 & n63506;
  assign n20740 = n20727 & ~n20739;
  assign n20741 = n20730 & ~n20740;
  assign n20742 = pi790 & ~n20725;
  assign n20743 = pi790 & ~n20741;
  assign n20744 = ~n20725 & n20743;
  assign n20745 = ~n20741 & n20742;
  assign n20746 = ~pi790 & ~n63506;
  assign n20747 = n62455 & ~n20746;
  assign n20748 = ~n63508 & n20747;
  assign n20749 = ~n20498 & n20713;
  assign n20750 = ~pi186 & ~n62455;
  assign n20751 = ~pi832 & ~n20750;
  assign n20752 = ~n63507 & n20751;
  assign po343 = ~n20340 & ~n20752;
  assign n20754 = ~pi187 & ~n2923;
  assign n20755 = ~pi770 & n7316;
  assign n20756 = ~n20754 & ~n20755;
  assign n20757 = ~n8420 & ~n20756;
  assign n20758 = ~pi785 & ~n20757;
  assign n20759 = ~n8425 & ~n20756;
  assign n20760 = pi1155 & ~n20759;
  assign n20761 = ~n8428 & n20757;
  assign n20762 = ~pi1155 & ~n20761;
  assign n20763 = ~n20760 & ~n20762;
  assign n20764 = pi785 & ~n20763;
  assign n20765 = ~n20758 & ~n20764;
  assign n20766 = ~pi781 & ~n20765;
  assign n20767 = ~n8435 & n20765;
  assign n20768 = pi1154 & ~n20767;
  assign n20769 = ~n8438 & n20765;
  assign n20770 = ~pi1154 & ~n20769;
  assign n20771 = ~n20768 & ~n20770;
  assign n20772 = pi781 & ~n20771;
  assign n20773 = ~n20766 & ~n20772;
  assign n20774 = ~pi619 & ~n20773;
  assign n20775 = pi619 & ~n20754;
  assign n20776 = ~pi1159 & ~n20775;
  assign n20777 = ~n20774 & n20776;
  assign n20778 = pi619 & ~n20773;
  assign n20779 = ~pi619 & ~n20754;
  assign n20780 = pi1159 & ~n20779;
  assign n20781 = ~n20778 & n20780;
  assign n20782 = pi619 & n20773;
  assign n20783 = ~pi619 & n20754;
  assign n20784 = pi1159 & ~n20783;
  assign n20785 = ~n20782 & n20784;
  assign n20786 = ~pi619 & n20773;
  assign n20787 = pi619 & n20754;
  assign n20788 = ~pi1159 & ~n20787;
  assign n20789 = ~n20786 & n20788;
  assign n20790 = ~n20785 & ~n20789;
  assign n20791 = ~n20777 & ~n20781;
  assign n20792 = pi789 & n63509;
  assign n20793 = ~pi789 & n20773;
  assign n20794 = ~pi789 & ~n20773;
  assign n20795 = pi789 & ~n63509;
  assign n20796 = ~n20794 & ~n20795;
  assign n20797 = ~n20792 & ~n20793;
  assign n20798 = ~n8595 & n63510;
  assign n20799 = n8595 & n20754;
  assign n20800 = ~n8595 & ~n63510;
  assign n20801 = n8595 & ~n20754;
  assign n20802 = ~n20800 & ~n20801;
  assign n20803 = ~n20798 & ~n20799;
  assign n20804 = ~n8334 & n63511;
  assign n20805 = n8334 & n20754;
  assign n20806 = ~n8413 & ~n20805;
  assign n20807 = ~n20804 & ~n20805;
  assign n20808 = ~n8413 & n20807;
  assign n20809 = ~n20804 & n20806;
  assign n20810 = pi726 & n7564;
  assign n20811 = ~n20754 & ~n20810;
  assign n20812 = ~pi778 & n20811;
  assign n20813 = ~pi625 & n20810;
  assign n20814 = ~n20811 & ~n20813;
  assign n20815 = pi1153 & ~n20814;
  assign n20816 = ~pi1153 & ~n20754;
  assign n20817 = ~n20813 & n20816;
  assign n20818 = ~n20815 & ~n20817;
  assign n20819 = pi778 & ~n20818;
  assign n20820 = ~n20812 & ~n20819;
  assign n20821 = ~n8490 & n20820;
  assign n20822 = ~n8492 & n20821;
  assign n20823 = ~n8494 & n20822;
  assign n20824 = ~n8496 & n20823;
  assign n20825 = ~n8508 & n20824;
  assign n20826 = pi647 & ~n20825;
  assign n20827 = ~pi647 & ~n20754;
  assign n20828 = ~n20826 & ~n20827;
  assign n20829 = n8373 & ~n20828;
  assign n20830 = ~pi647 & n20825;
  assign n20831 = pi647 & n20754;
  assign n20832 = ~pi1157 & ~n20831;
  assign n20833 = ~n20830 & n20832;
  assign n20834 = pi630 & n20833;
  assign n20835 = ~n20829 & ~n20834;
  assign n20836 = ~n63512 & n20835;
  assign n20837 = pi787 & ~n20836;
  assign n20838 = ~pi626 & ~n63510;
  assign n20839 = pi626 & ~n20754;
  assign n20840 = n8301 & ~n20839;
  assign n20841 = ~n20838 & n20840;
  assign n20842 = n8525 & n20823;
  assign n20843 = pi626 & ~n63510;
  assign n20844 = ~pi626 & ~n20754;
  assign n20845 = n8300 & ~n20844;
  assign n20846 = ~n20843 & n20845;
  assign n20847 = ~n20842 & ~n20846;
  assign n20848 = ~n20841 & ~n20842;
  assign n20849 = ~n20846 & n20848;
  assign n20850 = ~n20841 & n20847;
  assign n20851 = pi788 & ~n63513;
  assign n20852 = ~n7187 & ~n20811;
  assign n20853 = pi625 & n20852;
  assign n20854 = n20756 & ~n20852;
  assign n20855 = ~n20853 & ~n20854;
  assign n20856 = n20816 & ~n20855;
  assign n20857 = ~pi608 & ~n20815;
  assign n20858 = ~n20856 & n20857;
  assign n20859 = pi1153 & n20756;
  assign n20860 = ~n20853 & n20859;
  assign n20861 = pi608 & ~n20817;
  assign n20862 = ~n20860 & n20861;
  assign n20863 = ~n20858 & ~n20862;
  assign n20864 = pi778 & ~n20863;
  assign n20865 = ~pi778 & ~n20854;
  assign n20866 = ~n20864 & ~n20865;
  assign n20867 = ~pi609 & ~n20866;
  assign n20868 = pi609 & n20820;
  assign n20869 = ~pi1155 & ~n20868;
  assign n20870 = ~n20867 & n20869;
  assign n20871 = ~pi660 & ~n20760;
  assign n20872 = ~n20870 & n20871;
  assign n20873 = pi609 & ~n20866;
  assign n20874 = ~pi609 & n20820;
  assign n20875 = pi1155 & ~n20874;
  assign n20876 = ~n20873 & n20875;
  assign n20877 = pi660 & ~n20762;
  assign n20878 = ~n20876 & n20877;
  assign n20879 = ~n20872 & ~n20878;
  assign n20880 = pi785 & ~n20879;
  assign n20881 = ~pi785 & ~n20866;
  assign n20882 = ~n20880 & ~n20881;
  assign n20883 = pi618 & ~n20882;
  assign n20884 = ~pi618 & n20821;
  assign n20885 = pi1154 & ~n20884;
  assign n20886 = ~n20883 & n20885;
  assign n20887 = pi627 & ~n20770;
  assign n20888 = ~n20886 & n20887;
  assign n20889 = ~pi618 & ~n20882;
  assign n20890 = pi618 & n20821;
  assign n20891 = ~pi1154 & ~n20890;
  assign n20892 = ~n20889 & n20891;
  assign n20893 = ~pi627 & ~n20768;
  assign n20894 = ~n20892 & n20893;
  assign n20895 = pi781 & ~n20894;
  assign n20896 = ~n20888 & n20895;
  assign n20897 = ~n11431 & ~n20822;
  assign n20898 = ~n62884 & ~n63509;
  assign n20899 = ~n20897 & ~n20898;
  assign n20900 = pi789 & ~n20899;
  assign n20901 = ~pi781 & n20882;
  assign n20902 = ~n20900 & ~n20901;
  assign n20903 = ~n20896 & n20902;
  assign n20904 = n11434 & n20899;
  assign n20905 = ~n20903 & ~n20904;
  assign n20906 = ~n20888 & ~n20894;
  assign n20907 = pi781 & ~n20906;
  assign n20908 = ~pi781 & ~n20882;
  assign n20909 = ~n20907 & ~n20908;
  assign n20910 = ~pi619 & ~n20909;
  assign n20911 = pi619 & n20822;
  assign n20912 = ~pi1159 & ~n20911;
  assign n20913 = ~n20910 & n20912;
  assign n20914 = ~pi648 & ~n20785;
  assign n20915 = ~n20913 & n20914;
  assign n20916 = pi619 & ~n20909;
  assign n20917 = ~pi619 & n20822;
  assign n20918 = pi1159 & ~n20917;
  assign n20919 = ~n20916 & n20918;
  assign n20920 = pi648 & ~n20789;
  assign n20921 = ~n20919 & n20920;
  assign n20922 = pi789 & ~n20921;
  assign n20923 = pi789 & ~n20915;
  assign n20924 = ~n20921 & n20923;
  assign n20925 = ~n20915 & n20922;
  assign n20926 = ~pi789 & n20909;
  assign n20927 = n62894 & ~n20926;
  assign n20928 = ~n63514 & n20927;
  assign n20929 = n62894 & ~n20905;
  assign n20930 = ~n20851 & ~n63515;
  assign n20931 = ~n63030 & ~n20930;
  assign n20932 = n8498 & n63511;
  assign n20933 = n8615 & n20824;
  assign n20934 = pi629 & ~n20933;
  assign n20935 = ~n20932 & n20934;
  assign n20936 = n8499 & n63511;
  assign n20937 = n8606 & n20824;
  assign n20938 = ~pi629 & ~n20937;
  assign n20939 = ~n20936 & n20938;
  assign n20940 = pi792 & ~n20939;
  assign n20941 = pi792 & ~n20935;
  assign n20942 = ~n20939 & n20941;
  assign n20943 = ~n20936 & ~n20937;
  assign n20944 = ~pi629 & ~n20943;
  assign n20945 = ~n20932 & ~n20933;
  assign n20946 = pi629 & ~n20945;
  assign n20947 = ~n20944 & ~n20946;
  assign n20948 = pi792 & ~n20947;
  assign n20949 = ~n20935 & n20940;
  assign n20950 = ~n8651 & ~n63516;
  assign n20951 = ~n20931 & n20950;
  assign n20952 = ~n20837 & ~n20951;
  assign n20953 = pi644 & n20952;
  assign n20954 = ~pi787 & ~n20825;
  assign n20955 = pi1157 & ~n20828;
  assign n20956 = ~n20833 & ~n20955;
  assign n20957 = pi787 & ~n20956;
  assign n20958 = ~n20954 & ~n20957;
  assign n20959 = ~pi644 & n20958;
  assign n20960 = pi715 & ~n20959;
  assign n20961 = ~n20953 & n20960;
  assign n20962 = ~n8685 & n20754;
  assign n20963 = ~n8376 & n20804;
  assign n20964 = ~n8376 & ~n20807;
  assign n20965 = n8376 & n20754;
  assign n20966 = ~n20964 & ~n20965;
  assign n20967 = ~n20962 & ~n20963;
  assign n20968 = pi644 & ~n63517;
  assign n20969 = ~pi644 & n20754;
  assign n20970 = ~pi715 & ~n20969;
  assign n20971 = ~n20968 & n20970;
  assign n20972 = pi1160 & ~n20971;
  assign n20973 = ~n20961 & n20972;
  assign n20974 = ~pi644 & n20952;
  assign n20975 = pi644 & n20958;
  assign n20976 = ~pi715 & ~n20975;
  assign n20977 = ~n20974 & n20976;
  assign n20978 = ~pi644 & ~n63517;
  assign n20979 = pi644 & n20754;
  assign n20980 = pi715 & ~n20979;
  assign n20981 = ~n20978 & n20980;
  assign n20982 = ~pi1160 & ~n20981;
  assign n20983 = ~n20977 & n20982;
  assign n20984 = ~n20973 & ~n20983;
  assign n20985 = pi790 & ~n20984;
  assign n20986 = ~pi790 & n20952;
  assign n20987 = pi832 & ~n20986;
  assign n20988 = ~n20985 & n20987;
  assign n20989 = ~pi187 & ~n8098;
  assign n20990 = n8257 & ~n20989;
  assign n20991 = pi187 & ~n62765;
  assign n20992 = ~pi187 & n8009;
  assign n20993 = pi187 & n62874;
  assign n20994 = ~pi38 & ~n20993;
  assign n20995 = ~n20992 & n20994;
  assign n20996 = ~pi187 & ~n7357;
  assign n20997 = n8085 & ~n20996;
  assign n20998 = pi726 & ~n20997;
  assign n20999 = ~n20995 & n20998;
  assign n21000 = ~pi187 & ~pi726;
  assign n21001 = ~n8091 & n21000;
  assign n21002 = n62765 & ~n21001;
  assign n21003 = ~n20999 & n21002;
  assign n21004 = ~n20991 & ~n21003;
  assign n21005 = ~pi778 & ~n21004;
  assign n21006 = pi625 & n21004;
  assign n21007 = ~pi625 & n20989;
  assign n21008 = pi1153 & ~n21007;
  assign n21009 = ~n21006 & n21008;
  assign n21010 = ~pi625 & n21004;
  assign n21011 = pi625 & n20989;
  assign n21012 = ~pi1153 & ~n21011;
  assign n21013 = ~n21010 & n21012;
  assign n21014 = ~n21009 & ~n21013;
  assign n21015 = pi778 & ~n21014;
  assign n21016 = ~n21005 & ~n21015;
  assign n21017 = ~n62880 & ~n21016;
  assign n21018 = n62880 & ~n20989;
  assign n21019 = ~n62880 & n21016;
  assign n21020 = n62880 & n20989;
  assign n21021 = ~n21019 & ~n21020;
  assign n21022 = ~n21017 & ~n21018;
  assign n21023 = ~n62882 & ~n63518;
  assign n21024 = n62882 & n20989;
  assign n21025 = n62882 & ~n20989;
  assign n21026 = ~n62882 & n63518;
  assign n21027 = ~n21025 & ~n21026;
  assign n21028 = ~n21023 & ~n21024;
  assign n21029 = ~n8257 & ~n63519;
  assign n21030 = ~n8257 & n63519;
  assign n21031 = n8257 & n20989;
  assign n21032 = ~n21030 & ~n21031;
  assign n21033 = ~n20990 & ~n21029;
  assign n21034 = ~n8303 & ~n63520;
  assign n21035 = n8303 & n20989;
  assign n21036 = n8303 & ~n20989;
  assign n21037 = ~n8303 & n63520;
  assign n21038 = ~n21036 & ~n21037;
  assign n21039 = ~n21034 & ~n21035;
  assign n21040 = ~pi792 & ~n63521;
  assign n21041 = pi628 & n63521;
  assign n21042 = ~pi628 & n20989;
  assign n21043 = pi1156 & ~n21042;
  assign n21044 = ~pi628 & ~n20989;
  assign n21045 = pi628 & ~n63521;
  assign n21046 = ~n21044 & ~n21045;
  assign n21047 = pi1156 & ~n21046;
  assign n21048 = ~n21041 & n21043;
  assign n21049 = ~pi628 & n63521;
  assign n21050 = pi628 & n20989;
  assign n21051 = ~pi1156 & ~n21050;
  assign n21052 = ~n21049 & n21051;
  assign n21053 = ~n63522 & ~n21052;
  assign n21054 = pi792 & ~n21053;
  assign n21055 = ~n21040 & ~n21054;
  assign n21056 = ~pi787 & ~n21055;
  assign n21057 = pi647 & n21055;
  assign n21058 = ~pi647 & n20989;
  assign n21059 = pi1157 & ~n21058;
  assign n21060 = ~pi647 & ~n20989;
  assign n21061 = pi647 & ~n21055;
  assign n21062 = ~n21060 & ~n21061;
  assign n21063 = pi1157 & ~n21062;
  assign n21064 = ~n21057 & n21059;
  assign n21065 = ~pi647 & n21055;
  assign n21066 = pi647 & n20989;
  assign n21067 = ~pi1157 & ~n21066;
  assign n21068 = ~n21065 & n21067;
  assign n21069 = ~n63523 & ~n21068;
  assign n21070 = pi787 & ~n21069;
  assign n21071 = ~n21056 & ~n21070;
  assign n21072 = ~pi644 & n21071;
  assign n21073 = pi715 & ~n21072;
  assign n21074 = pi770 & n8091;
  assign n21075 = ~pi770 & ~n14285;
  assign n21076 = pi187 & ~n21075;
  assign n21077 = ~pi187 & ~pi770;
  assign n21078 = n10343 & n21077;
  assign n21079 = ~n21076 & ~n21078;
  assign n21080 = pi770 & ~n8091;
  assign n21081 = ~pi770 & ~n10343;
  assign n21082 = ~n21080 & ~n21081;
  assign n21083 = ~pi187 & ~n21082;
  assign n21084 = ~pi187 & ~n62977;
  assign n21085 = ~pi770 & ~n21084;
  assign n21086 = ~n14285 & n21085;
  assign n21087 = ~n21083 & ~n21086;
  assign n21088 = ~n21074 & n21079;
  assign n21089 = n62765 & n63524;
  assign n21090 = ~n20991 & ~n21089;
  assign n21091 = ~n8135 & ~n21090;
  assign n21092 = n8135 & ~n20989;
  assign n21093 = ~n21091 & ~n21092;
  assign n21094 = ~pi785 & ~n21093;
  assign n21095 = ~n8136 & ~n20989;
  assign n21096 = pi609 & n21091;
  assign n21097 = ~n21095 & ~n21096;
  assign n21098 = pi1155 & ~n21097;
  assign n21099 = ~n8148 & ~n20989;
  assign n21100 = ~pi609 & n21091;
  assign n21101 = ~n21099 & ~n21100;
  assign n21102 = ~pi1155 & ~n21101;
  assign n21103 = ~n21098 & ~n21102;
  assign n21104 = pi785 & ~n21103;
  assign n21105 = ~n21094 & ~n21104;
  assign n21106 = ~pi781 & ~n21105;
  assign n21107 = pi618 & n21105;
  assign n21108 = ~pi618 & n20989;
  assign n21109 = pi1154 & ~n21108;
  assign n21110 = ~n21107 & n21109;
  assign n21111 = ~pi618 & n21105;
  assign n21112 = pi618 & n20989;
  assign n21113 = ~pi1154 & ~n21112;
  assign n21114 = ~n21111 & n21113;
  assign n21115 = ~n21110 & ~n21114;
  assign n21116 = pi781 & ~n21115;
  assign n21117 = ~n21106 & ~n21116;
  assign n21118 = ~pi789 & ~n21117;
  assign n21119 = ~pi619 & n21117;
  assign n21120 = pi619 & n20989;
  assign n21121 = ~pi1159 & ~n21120;
  assign n21122 = ~n21119 & n21121;
  assign n21123 = pi619 & n21117;
  assign n21124 = ~pi619 & n20989;
  assign n21125 = pi1159 & ~n21124;
  assign n21126 = ~n21123 & n21125;
  assign n21127 = ~n21122 & ~n21126;
  assign n21128 = pi789 & ~n21127;
  assign n21129 = ~n21118 & ~n21128;
  assign n21130 = ~n8595 & n21129;
  assign n21131 = n8595 & n20989;
  assign n21132 = ~n21130 & ~n21131;
  assign n21133 = ~n8334 & ~n21132;
  assign n21134 = n8334 & n20989;
  assign n21135 = ~n21133 & ~n21134;
  assign n21136 = ~n8376 & ~n21135;
  assign n21137 = n8376 & n20989;
  assign n21138 = n8376 & ~n20989;
  assign n21139 = ~n8376 & n21135;
  assign n21140 = ~n21138 & ~n21139;
  assign n21141 = ~n21136 & ~n21137;
  assign n21142 = pi644 & n63525;
  assign n21143 = ~pi644 & n20989;
  assign n21144 = ~pi715 & ~n21143;
  assign n21145 = ~n21142 & n21144;
  assign n21146 = pi1160 & ~n21145;
  assign n21147 = ~n21073 & n21146;
  assign n21148 = pi644 & n21071;
  assign n21149 = ~pi715 & ~n21148;
  assign n21150 = ~pi644 & n63525;
  assign n21151 = pi644 & n20989;
  assign n21152 = pi715 & ~n21151;
  assign n21153 = ~n21150 & n21152;
  assign n21154 = ~pi1160 & ~n21153;
  assign n21155 = ~n21149 & n21154;
  assign n21156 = ~n21147 & ~n21155;
  assign n21157 = pi790 & ~n21156;
  assign n21158 = ~pi644 & n21154;
  assign n21159 = pi644 & n21146;
  assign n21160 = n14029 & ~n21145;
  assign n21161 = pi790 & ~n63526;
  assign n21162 = ~n21158 & n21161;
  assign n21163 = ~n63052 & n21132;
  assign n21164 = n8331 & ~n21046;
  assign n21165 = ~pi629 & n63522;
  assign n21166 = pi629 & n21052;
  assign n21167 = ~n63527 & ~n21166;
  assign n21168 = ~n21163 & n21167;
  assign n21169 = pi792 & ~n21168;
  assign n21170 = n12979 & n21129;
  assign n21171 = ~pi641 & n63520;
  assign n21172 = pi641 & ~n20989;
  assign n21173 = n8417 & ~n21172;
  assign n21174 = ~n21171 & n21173;
  assign n21175 = pi641 & n63520;
  assign n21176 = ~pi641 & ~n20989;
  assign n21177 = n8416 & ~n21176;
  assign n21178 = ~n21175 & n21177;
  assign n21179 = ~n21174 & ~n21178;
  assign n21180 = ~n21170 & n21179;
  assign n21181 = pi788 & ~n21180;
  assign n21182 = pi619 & n63519;
  assign n21183 = ~pi1159 & ~n21182;
  assign n21184 = ~pi648 & ~n21126;
  assign n21185 = ~n21183 & n21184;
  assign n21186 = ~pi619 & n63519;
  assign n21187 = pi1159 & ~n21186;
  assign n21188 = pi648 & ~n21187;
  assign n21189 = pi648 & ~n21122;
  assign n21190 = ~n21187 & n21189;
  assign n21191 = ~n21122 & n21188;
  assign n21192 = ~n21185 & ~n63528;
  assign n21193 = pi789 & ~n21192;
  assign n21194 = pi618 & ~n63518;
  assign n21195 = ~pi1154 & ~n21194;
  assign n21196 = ~pi627 & ~n21110;
  assign n21197 = ~n21195 & n21196;
  assign n21198 = ~pi618 & ~n63518;
  assign n21199 = pi1154 & ~n21198;
  assign n21200 = pi627 & ~n21114;
  assign n21201 = ~n21199 & n21200;
  assign n21202 = ~n21197 & ~n21201;
  assign n21203 = pi781 & ~n21202;
  assign n21204 = ~pi618 & n21196;
  assign n21205 = pi618 & n21200;
  assign n21206 = pi781 & ~n21205;
  assign n21207 = ~n21204 & n21206;
  assign n21208 = ~pi187 & n10353;
  assign n21209 = pi187 & n10355;
  assign n21210 = pi770 & ~n10357;
  assign n21211 = ~n21209 & n21210;
  assign n21212 = ~n21208 & n21211;
  assign n21213 = pi187 & n10363;
  assign n21214 = ~pi187 & ~n62980;
  assign n21215 = ~pi770 & ~n21214;
  assign n21216 = ~n21213 & n21215;
  assign n21217 = pi726 & ~n21216;
  assign n21218 = ~n21212 & n21217;
  assign n21219 = ~pi726 & ~n63524;
  assign n21220 = n62765 & ~n21219;
  assign n21221 = n62765 & ~n21218;
  assign n21222 = ~n21219 & n21221;
  assign n21223 = ~n21218 & n21220;
  assign n21224 = ~n20991 & ~n63529;
  assign n21225 = ~pi625 & n21224;
  assign n21226 = pi625 & n21090;
  assign n21227 = ~pi1153 & ~n21226;
  assign n21228 = ~n21225 & n21227;
  assign n21229 = ~pi608 & ~n21009;
  assign n21230 = ~n21228 & n21229;
  assign n21231 = pi625 & n21224;
  assign n21232 = ~pi625 & n21090;
  assign n21233 = pi1153 & ~n21232;
  assign n21234 = ~n21231 & n21233;
  assign n21235 = pi608 & ~n21013;
  assign n21236 = ~n21234 & n21235;
  assign n21237 = ~n21230 & ~n21236;
  assign n21238 = pi778 & ~n21237;
  assign n21239 = ~pi778 & n21224;
  assign n21240 = ~pi778 & ~n21224;
  assign n21241 = pi778 & ~n21236;
  assign n21242 = ~n21230 & n21241;
  assign n21243 = ~n21240 & ~n21242;
  assign n21244 = ~n21238 & ~n21239;
  assign n21245 = ~pi785 & ~n63530;
  assign n21246 = ~pi609 & n63530;
  assign n21247 = pi609 & n21016;
  assign n21248 = ~pi1155 & ~n21247;
  assign n21249 = ~n21246 & n21248;
  assign n21250 = ~pi660 & ~n21098;
  assign n21251 = ~n21249 & n21250;
  assign n21252 = pi609 & n63530;
  assign n21253 = ~pi609 & n21016;
  assign n21254 = pi1155 & ~n21253;
  assign n21255 = ~n21252 & n21254;
  assign n21256 = pi660 & ~n21102;
  assign n21257 = ~n21255 & n21256;
  assign n21258 = pi785 & ~n21257;
  assign n21259 = ~n21251 & n21258;
  assign n21260 = ~n21251 & ~n21257;
  assign n21261 = pi785 & ~n21260;
  assign n21262 = ~pi785 & n63530;
  assign n21263 = ~n21261 & ~n21262;
  assign n21264 = ~n21245 & ~n21259;
  assign n21265 = ~n21207 & ~n63531;
  assign n21266 = pi618 & ~n63531;
  assign n21267 = n21199 & ~n21266;
  assign n21268 = n21200 & ~n21267;
  assign n21269 = ~n21197 & ~n21268;
  assign n21270 = pi781 & ~n21269;
  assign n21271 = pi781 & ~n21204;
  assign n21272 = ~n63531 & ~n21271;
  assign n21273 = ~n21270 & ~n21272;
  assign n21274 = ~pi618 & ~n63531;
  assign n21275 = n21195 & ~n21274;
  assign n21276 = n21196 & ~n21275;
  assign n21277 = ~n21268 & ~n21276;
  assign n21278 = pi781 & ~n21277;
  assign n21279 = ~pi781 & ~n63531;
  assign n21280 = ~n21278 & ~n21279;
  assign n21281 = ~n21203 & ~n21265;
  assign n21282 = ~pi619 & n21184;
  assign n21283 = pi619 & n21189;
  assign n21284 = n11422 & ~n21122;
  assign n21285 = pi789 & ~n63533;
  assign n21286 = ~n21282 & n21285;
  assign n21287 = ~n63532 & ~n21286;
  assign n21288 = ~pi619 & ~n63532;
  assign n21289 = n21183 & ~n21288;
  assign n21290 = n21184 & ~n21289;
  assign n21291 = pi619 & ~n63532;
  assign n21292 = n21187 & ~n21291;
  assign n21293 = n21189 & ~n21292;
  assign n21294 = ~n21290 & ~n21293;
  assign n21295 = pi789 & ~n21294;
  assign n21296 = ~pi789 & ~n63532;
  assign n21297 = ~n21295 & ~n21296;
  assign n21298 = ~n21193 & ~n21287;
  assign n21299 = n62894 & ~n63534;
  assign n21300 = ~n63030 & ~n21299;
  assign n21301 = ~n63030 & ~n21181;
  assign n21302 = ~n21299 & n21301;
  assign n21303 = ~n21181 & n21300;
  assign n21304 = ~pi788 & n63534;
  assign n21305 = ~pi626 & n63534;
  assign n21306 = pi626 & n63520;
  assign n21307 = ~pi641 & ~n21306;
  assign n21308 = ~n21305 & n21307;
  assign n21309 = ~pi626 & ~n21129;
  assign n21310 = pi626 & ~n20989;
  assign n21311 = pi641 & ~n21310;
  assign n21312 = ~n21309 & n21311;
  assign n21313 = ~pi1158 & ~n21312;
  assign n21314 = ~n21308 & n21313;
  assign n21315 = pi626 & n63534;
  assign n21316 = ~pi626 & n63520;
  assign n21317 = pi641 & ~n21316;
  assign n21318 = ~n21315 & n21317;
  assign n21319 = pi626 & ~n21129;
  assign n21320 = ~pi626 & ~n20989;
  assign n21321 = ~pi641 & ~n21320;
  assign n21322 = ~n21319 & n21321;
  assign n21323 = pi1158 & ~n21322;
  assign n21324 = ~n21318 & n21323;
  assign n21325 = ~n21314 & ~n21324;
  assign n21326 = pi788 & ~n21325;
  assign n21327 = ~n21304 & ~n21326;
  assign n21328 = ~pi628 & n21327;
  assign n21329 = pi628 & ~n21132;
  assign n21330 = ~pi1156 & ~n21329;
  assign n21331 = ~n21328 & n21330;
  assign n21332 = ~pi629 & ~n63522;
  assign n21333 = ~n21331 & n21332;
  assign n21334 = pi628 & n21327;
  assign n21335 = ~pi628 & ~n21132;
  assign n21336 = pi1156 & ~n21335;
  assign n21337 = ~n21334 & n21336;
  assign n21338 = pi629 & ~n21052;
  assign n21339 = ~n21337 & n21338;
  assign n21340 = ~n21333 & ~n21339;
  assign n21341 = pi792 & ~n21340;
  assign n21342 = ~pi792 & n21327;
  assign n21343 = ~n21341 & ~n21342;
  assign n21344 = ~n21169 & ~n63535;
  assign n21345 = ~n8651 & n63536;
  assign n21346 = ~n8413 & n21135;
  assign n21347 = n8373 & ~n21062;
  assign n21348 = ~pi630 & n63523;
  assign n21349 = pi630 & n21068;
  assign n21350 = ~n63537 & ~n21349;
  assign n21351 = ~n21346 & ~n21349;
  assign n21352 = ~n63537 & n21351;
  assign n21353 = ~n21346 & n21350;
  assign n21354 = pi787 & ~n63538;
  assign n21355 = ~n62896 & n63536;
  assign n21356 = ~pi647 & ~n63536;
  assign n21357 = pi647 & ~n21135;
  assign n21358 = ~pi1157 & ~n21357;
  assign n21359 = ~n21356 & n21358;
  assign n21360 = ~pi630 & ~n63523;
  assign n21361 = ~n21359 & n21360;
  assign n21362 = pi647 & ~n63536;
  assign n21363 = ~pi647 & ~n21135;
  assign n21364 = pi1157 & ~n21363;
  assign n21365 = ~n21362 & n21364;
  assign n21366 = pi630 & ~n21068;
  assign n21367 = ~n21365 & n21366;
  assign n21368 = ~n21361 & ~n21367;
  assign n21369 = n63538 & ~n21355;
  assign n21370 = pi787 & n63539;
  assign n21371 = ~pi787 & n63536;
  assign n21372 = ~n21370 & ~n21371;
  assign n21373 = pi787 & ~n63539;
  assign n21374 = ~pi787 & ~n63536;
  assign n21375 = ~n21373 & ~n21374;
  assign n21376 = ~n21345 & ~n21354;
  assign n21377 = ~n21162 & n63540;
  assign n21378 = ~pi644 & n63540;
  assign n21379 = n21149 & ~n21378;
  assign n21380 = n21154 & ~n21379;
  assign n21381 = ~n21147 & ~n21380;
  assign n21382 = pi790 & ~n21381;
  assign n21383 = ~n21161 & n63540;
  assign n21384 = ~n21382 & ~n21383;
  assign n21385 = ~n21157 & ~n21377;
  assign n21386 = pi644 & n63540;
  assign n21387 = n21073 & ~n21386;
  assign n21388 = n21146 & ~n21387;
  assign n21389 = pi790 & ~n21380;
  assign n21390 = pi790 & ~n21388;
  assign n21391 = ~n21380 & n21390;
  assign n21392 = ~n21388 & n21389;
  assign n21393 = ~pi790 & ~n63540;
  assign n21394 = n62455 & ~n21393;
  assign n21395 = ~n63542 & n21394;
  assign n21396 = n62455 & ~n63541;
  assign n21397 = ~pi187 & ~n62455;
  assign n21398 = ~pi832 & ~n21397;
  assign n21399 = ~n63543 & n21398;
  assign po344 = ~n20988 & ~n21399;
  assign n21401 = ~pi188 & ~n2923;
  assign n21402 = ~pi768 & n7316;
  assign n21403 = ~n21401 & ~n21402;
  assign n21404 = ~n8420 & ~n21403;
  assign n21405 = ~pi785 & ~n21404;
  assign n21406 = ~n8425 & ~n21403;
  assign n21407 = pi1155 & ~n21406;
  assign n21408 = ~n8428 & n21404;
  assign n21409 = ~pi1155 & ~n21408;
  assign n21410 = ~n21407 & ~n21409;
  assign n21411 = pi785 & ~n21410;
  assign n21412 = ~n21405 & ~n21411;
  assign n21413 = ~pi781 & ~n21412;
  assign n21414 = ~n8435 & n21412;
  assign n21415 = pi1154 & ~n21414;
  assign n21416 = ~n8438 & n21412;
  assign n21417 = ~pi1154 & ~n21416;
  assign n21418 = ~n21415 & ~n21417;
  assign n21419 = pi781 & ~n21418;
  assign n21420 = ~n21413 & ~n21419;
  assign n21421 = ~pi619 & ~n21420;
  assign n21422 = pi619 & ~n21401;
  assign n21423 = ~pi1159 & ~n21422;
  assign n21424 = ~n21421 & n21423;
  assign n21425 = pi619 & ~n21420;
  assign n21426 = ~pi619 & ~n21401;
  assign n21427 = pi1159 & ~n21426;
  assign n21428 = ~n21425 & n21427;
  assign n21429 = pi619 & n21420;
  assign n21430 = ~pi619 & n21401;
  assign n21431 = pi1159 & ~n21430;
  assign n21432 = ~n21429 & n21431;
  assign n21433 = ~pi619 & n21420;
  assign n21434 = pi619 & n21401;
  assign n21435 = ~pi1159 & ~n21434;
  assign n21436 = ~n21433 & n21435;
  assign n21437 = ~n21432 & ~n21436;
  assign n21438 = ~n21424 & ~n21428;
  assign n21439 = pi789 & n63544;
  assign n21440 = ~pi789 & n21420;
  assign n21441 = ~pi789 & ~n21420;
  assign n21442 = pi789 & ~n63544;
  assign n21443 = ~n21441 & ~n21442;
  assign n21444 = ~n21439 & ~n21440;
  assign n21445 = ~n8595 & n63545;
  assign n21446 = n8595 & n21401;
  assign n21447 = ~n8595 & ~n63545;
  assign n21448 = n8595 & ~n21401;
  assign n21449 = ~n21447 & ~n21448;
  assign n21450 = ~n21445 & ~n21446;
  assign n21451 = ~n8334 & n63546;
  assign n21452 = n8334 & n21401;
  assign n21453 = ~n8413 & ~n21452;
  assign n21454 = ~n21451 & ~n21452;
  assign n21455 = ~n8413 & n21454;
  assign n21456 = ~n21451 & n21453;
  assign n21457 = pi705 & n7564;
  assign n21458 = ~n21401 & ~n21457;
  assign n21459 = ~pi778 & n21458;
  assign n21460 = ~pi625 & n21457;
  assign n21461 = ~n21458 & ~n21460;
  assign n21462 = pi1153 & ~n21461;
  assign n21463 = ~pi1153 & ~n21401;
  assign n21464 = ~n21460 & n21463;
  assign n21465 = ~n21462 & ~n21464;
  assign n21466 = pi778 & ~n21465;
  assign n21467 = ~n21459 & ~n21466;
  assign n21468 = ~n8490 & n21467;
  assign n21469 = ~n8492 & n21468;
  assign n21470 = ~n8494 & n21469;
  assign n21471 = ~n8496 & n21470;
  assign n21472 = ~n8508 & n21471;
  assign n21473 = pi647 & ~n21472;
  assign n21474 = ~pi647 & ~n21401;
  assign n21475 = ~n21473 & ~n21474;
  assign n21476 = n8373 & ~n21475;
  assign n21477 = ~pi647 & n21472;
  assign n21478 = pi647 & n21401;
  assign n21479 = ~pi1157 & ~n21478;
  assign n21480 = ~n21477 & n21479;
  assign n21481 = pi630 & n21480;
  assign n21482 = ~n21476 & ~n21481;
  assign n21483 = ~n63547 & n21482;
  assign n21484 = pi787 & ~n21483;
  assign n21485 = ~pi626 & ~n63545;
  assign n21486 = pi626 & ~n21401;
  assign n21487 = n8301 & ~n21486;
  assign n21488 = ~n21485 & n21487;
  assign n21489 = n8525 & n21470;
  assign n21490 = pi626 & ~n63545;
  assign n21491 = ~pi626 & ~n21401;
  assign n21492 = n8300 & ~n21491;
  assign n21493 = ~n21490 & n21492;
  assign n21494 = ~n21489 & ~n21493;
  assign n21495 = ~n21488 & ~n21489;
  assign n21496 = ~n21493 & n21495;
  assign n21497 = ~n21488 & n21494;
  assign n21498 = pi788 & ~n63548;
  assign n21499 = ~n7187 & ~n21458;
  assign n21500 = pi625 & n21499;
  assign n21501 = n21403 & ~n21499;
  assign n21502 = ~n21500 & ~n21501;
  assign n21503 = n21463 & ~n21502;
  assign n21504 = ~pi608 & ~n21462;
  assign n21505 = ~n21503 & n21504;
  assign n21506 = pi1153 & n21403;
  assign n21507 = ~n21500 & n21506;
  assign n21508 = pi608 & ~n21464;
  assign n21509 = ~n21507 & n21508;
  assign n21510 = ~n21505 & ~n21509;
  assign n21511 = pi778 & ~n21510;
  assign n21512 = ~pi778 & ~n21501;
  assign n21513 = ~n21511 & ~n21512;
  assign n21514 = ~pi609 & ~n21513;
  assign n21515 = pi609 & n21467;
  assign n21516 = ~pi1155 & ~n21515;
  assign n21517 = ~n21514 & n21516;
  assign n21518 = ~pi660 & ~n21407;
  assign n21519 = ~n21517 & n21518;
  assign n21520 = pi609 & ~n21513;
  assign n21521 = ~pi609 & n21467;
  assign n21522 = pi1155 & ~n21521;
  assign n21523 = ~n21520 & n21522;
  assign n21524 = pi660 & ~n21409;
  assign n21525 = ~n21523 & n21524;
  assign n21526 = ~n21519 & ~n21525;
  assign n21527 = pi785 & ~n21526;
  assign n21528 = ~pi785 & ~n21513;
  assign n21529 = ~n21527 & ~n21528;
  assign n21530 = pi618 & ~n21529;
  assign n21531 = ~pi618 & n21468;
  assign n21532 = pi1154 & ~n21531;
  assign n21533 = ~n21530 & n21532;
  assign n21534 = pi627 & ~n21417;
  assign n21535 = ~n21533 & n21534;
  assign n21536 = ~pi618 & ~n21529;
  assign n21537 = pi618 & n21468;
  assign n21538 = ~pi1154 & ~n21537;
  assign n21539 = ~n21536 & n21538;
  assign n21540 = ~pi627 & ~n21415;
  assign n21541 = ~n21539 & n21540;
  assign n21542 = pi781 & ~n21541;
  assign n21543 = ~n21535 & n21542;
  assign n21544 = ~n11431 & ~n21469;
  assign n21545 = ~n62884 & ~n63544;
  assign n21546 = ~n21544 & ~n21545;
  assign n21547 = pi789 & ~n21546;
  assign n21548 = ~pi781 & n21529;
  assign n21549 = ~n21547 & ~n21548;
  assign n21550 = ~n21543 & n21549;
  assign n21551 = n11434 & n21546;
  assign n21552 = ~n21550 & ~n21551;
  assign n21553 = ~n21535 & ~n21541;
  assign n21554 = pi781 & ~n21553;
  assign n21555 = ~pi781 & ~n21529;
  assign n21556 = ~n21554 & ~n21555;
  assign n21557 = ~pi619 & ~n21556;
  assign n21558 = pi619 & n21469;
  assign n21559 = ~pi1159 & ~n21558;
  assign n21560 = ~n21557 & n21559;
  assign n21561 = ~pi648 & ~n21432;
  assign n21562 = ~n21560 & n21561;
  assign n21563 = pi619 & ~n21556;
  assign n21564 = ~pi619 & n21469;
  assign n21565 = pi1159 & ~n21564;
  assign n21566 = ~n21563 & n21565;
  assign n21567 = pi648 & ~n21436;
  assign n21568 = ~n21566 & n21567;
  assign n21569 = pi789 & ~n21568;
  assign n21570 = pi789 & ~n21562;
  assign n21571 = ~n21568 & n21570;
  assign n21572 = ~n21562 & n21569;
  assign n21573 = ~pi789 & n21556;
  assign n21574 = n62894 & ~n21573;
  assign n21575 = ~n63549 & n21574;
  assign n21576 = n62894 & ~n21552;
  assign n21577 = ~n21498 & ~n63550;
  assign n21578 = ~n63030 & ~n21577;
  assign n21579 = n8498 & n63546;
  assign n21580 = n8615 & n21471;
  assign n21581 = pi629 & ~n21580;
  assign n21582 = ~n21579 & n21581;
  assign n21583 = n8499 & n63546;
  assign n21584 = n8606 & n21471;
  assign n21585 = ~pi629 & ~n21584;
  assign n21586 = ~n21583 & n21585;
  assign n21587 = pi792 & ~n21586;
  assign n21588 = pi792 & ~n21582;
  assign n21589 = ~n21586 & n21588;
  assign n21590 = ~n21583 & ~n21584;
  assign n21591 = ~pi629 & ~n21590;
  assign n21592 = ~n21579 & ~n21580;
  assign n21593 = pi629 & ~n21592;
  assign n21594 = ~n21591 & ~n21593;
  assign n21595 = pi792 & ~n21594;
  assign n21596 = ~n21582 & n21587;
  assign n21597 = ~n8651 & ~n63551;
  assign n21598 = ~n21578 & n21597;
  assign n21599 = ~n21484 & ~n21598;
  assign n21600 = pi644 & n21599;
  assign n21601 = ~pi787 & ~n21472;
  assign n21602 = pi1157 & ~n21475;
  assign n21603 = ~n21480 & ~n21602;
  assign n21604 = pi787 & ~n21603;
  assign n21605 = ~n21601 & ~n21604;
  assign n21606 = ~pi644 & n21605;
  assign n21607 = pi715 & ~n21606;
  assign n21608 = ~n21600 & n21607;
  assign n21609 = ~n8685 & n21401;
  assign n21610 = ~n8376 & n21451;
  assign n21611 = ~n8376 & ~n21454;
  assign n21612 = n8376 & n21401;
  assign n21613 = ~n21611 & ~n21612;
  assign n21614 = ~n21609 & ~n21610;
  assign n21615 = pi644 & ~n63552;
  assign n21616 = ~pi644 & n21401;
  assign n21617 = ~pi715 & ~n21616;
  assign n21618 = ~n21615 & n21617;
  assign n21619 = pi1160 & ~n21618;
  assign n21620 = ~n21608 & n21619;
  assign n21621 = ~pi644 & n21599;
  assign n21622 = pi644 & n21605;
  assign n21623 = ~pi715 & ~n21622;
  assign n21624 = ~n21621 & n21623;
  assign n21625 = ~pi644 & ~n63552;
  assign n21626 = pi644 & n21401;
  assign n21627 = pi715 & ~n21626;
  assign n21628 = ~n21625 & n21627;
  assign n21629 = ~pi1160 & ~n21628;
  assign n21630 = ~n21624 & n21629;
  assign n21631 = ~n21620 & ~n21630;
  assign n21632 = pi790 & ~n21631;
  assign n21633 = ~pi790 & n21599;
  assign n21634 = pi832 & ~n21633;
  assign n21635 = ~n21632 & n21634;
  assign n21636 = ~pi188 & ~n8098;
  assign n21637 = n8257 & ~n21636;
  assign n21638 = pi188 & ~n62765;
  assign n21639 = ~pi188 & n8009;
  assign n21640 = pi188 & n62874;
  assign n21641 = ~pi38 & ~n21640;
  assign n21642 = ~n21639 & n21641;
  assign n21643 = ~pi188 & ~n7357;
  assign n21644 = n8085 & ~n21643;
  assign n21645 = pi705 & ~n21644;
  assign n21646 = ~n21642 & n21645;
  assign n21647 = ~pi188 & ~pi705;
  assign n21648 = ~n8091 & n21647;
  assign n21649 = n62765 & ~n21648;
  assign n21650 = ~n21646 & n21649;
  assign n21651 = ~n21638 & ~n21650;
  assign n21652 = ~pi778 & ~n21651;
  assign n21653 = pi625 & n21651;
  assign n21654 = ~pi625 & n21636;
  assign n21655 = pi1153 & ~n21654;
  assign n21656 = ~n21653 & n21655;
  assign n21657 = ~pi625 & n21651;
  assign n21658 = pi625 & n21636;
  assign n21659 = ~pi1153 & ~n21658;
  assign n21660 = ~n21657 & n21659;
  assign n21661 = ~n21656 & ~n21660;
  assign n21662 = pi778 & ~n21661;
  assign n21663 = ~n21652 & ~n21662;
  assign n21664 = ~n62880 & ~n21663;
  assign n21665 = n62880 & ~n21636;
  assign n21666 = ~n62880 & n21663;
  assign n21667 = n62880 & n21636;
  assign n21668 = ~n21666 & ~n21667;
  assign n21669 = ~n21664 & ~n21665;
  assign n21670 = ~n62882 & ~n63553;
  assign n21671 = n62882 & n21636;
  assign n21672 = n62882 & ~n21636;
  assign n21673 = ~n62882 & n63553;
  assign n21674 = ~n21672 & ~n21673;
  assign n21675 = ~n21670 & ~n21671;
  assign n21676 = ~n8257 & ~n63554;
  assign n21677 = ~n8257 & n63554;
  assign n21678 = n8257 & n21636;
  assign n21679 = ~n21677 & ~n21678;
  assign n21680 = ~n21637 & ~n21676;
  assign n21681 = ~n8303 & ~n63555;
  assign n21682 = n8303 & n21636;
  assign n21683 = n8303 & ~n21636;
  assign n21684 = ~n8303 & n63555;
  assign n21685 = ~n21683 & ~n21684;
  assign n21686 = ~n21681 & ~n21682;
  assign n21687 = ~pi792 & ~n63556;
  assign n21688 = pi628 & n63556;
  assign n21689 = ~pi628 & n21636;
  assign n21690 = pi1156 & ~n21689;
  assign n21691 = ~pi628 & ~n21636;
  assign n21692 = pi628 & ~n63556;
  assign n21693 = ~n21691 & ~n21692;
  assign n21694 = pi1156 & ~n21693;
  assign n21695 = ~n21688 & n21690;
  assign n21696 = ~pi628 & n63556;
  assign n21697 = pi628 & n21636;
  assign n21698 = ~pi1156 & ~n21697;
  assign n21699 = ~n21696 & n21698;
  assign n21700 = ~n63557 & ~n21699;
  assign n21701 = pi792 & ~n21700;
  assign n21702 = ~n21687 & ~n21701;
  assign n21703 = ~pi787 & ~n21702;
  assign n21704 = pi647 & n21702;
  assign n21705 = ~pi647 & n21636;
  assign n21706 = pi1157 & ~n21705;
  assign n21707 = ~pi647 & ~n21636;
  assign n21708 = pi647 & ~n21702;
  assign n21709 = ~n21707 & ~n21708;
  assign n21710 = pi1157 & ~n21709;
  assign n21711 = ~n21704 & n21706;
  assign n21712 = ~pi647 & n21702;
  assign n21713 = pi647 & n21636;
  assign n21714 = ~pi1157 & ~n21713;
  assign n21715 = ~n21712 & n21714;
  assign n21716 = ~n63558 & ~n21715;
  assign n21717 = pi787 & ~n21716;
  assign n21718 = ~n21703 & ~n21717;
  assign n21719 = ~pi644 & n21718;
  assign n21720 = pi715 & ~n21719;
  assign n21721 = pi768 & n8091;
  assign n21722 = ~pi768 & ~n14285;
  assign n21723 = pi188 & ~n21722;
  assign n21724 = ~pi188 & ~pi768;
  assign n21725 = n10343 & n21724;
  assign n21726 = ~n21723 & ~n21725;
  assign n21727 = pi768 & ~n8091;
  assign n21728 = ~pi768 & ~n10343;
  assign n21729 = ~n21727 & ~n21728;
  assign n21730 = ~pi188 & ~n21729;
  assign n21731 = ~pi188 & ~n62977;
  assign n21732 = ~pi768 & ~n21731;
  assign n21733 = ~n14285 & n21732;
  assign n21734 = ~n21730 & ~n21733;
  assign n21735 = ~n21721 & n21726;
  assign n21736 = n62765 & n63559;
  assign n21737 = ~n21638 & ~n21736;
  assign n21738 = ~n8135 & ~n21737;
  assign n21739 = n8135 & ~n21636;
  assign n21740 = ~n21738 & ~n21739;
  assign n21741 = ~pi785 & ~n21740;
  assign n21742 = ~n8136 & ~n21636;
  assign n21743 = pi609 & n21738;
  assign n21744 = ~n21742 & ~n21743;
  assign n21745 = pi1155 & ~n21744;
  assign n21746 = ~n8148 & ~n21636;
  assign n21747 = ~pi609 & n21738;
  assign n21748 = ~n21746 & ~n21747;
  assign n21749 = ~pi1155 & ~n21748;
  assign n21750 = ~n21745 & ~n21749;
  assign n21751 = pi785 & ~n21750;
  assign n21752 = ~n21741 & ~n21751;
  assign n21753 = ~pi781 & ~n21752;
  assign n21754 = pi618 & n21752;
  assign n21755 = ~pi618 & n21636;
  assign n21756 = pi1154 & ~n21755;
  assign n21757 = ~n21754 & n21756;
  assign n21758 = ~pi618 & n21752;
  assign n21759 = pi618 & n21636;
  assign n21760 = ~pi1154 & ~n21759;
  assign n21761 = ~n21758 & n21760;
  assign n21762 = ~n21757 & ~n21761;
  assign n21763 = pi781 & ~n21762;
  assign n21764 = ~n21753 & ~n21763;
  assign n21765 = ~pi789 & ~n21764;
  assign n21766 = ~pi619 & n21764;
  assign n21767 = pi619 & n21636;
  assign n21768 = ~pi1159 & ~n21767;
  assign n21769 = ~n21766 & n21768;
  assign n21770 = pi619 & n21764;
  assign n21771 = ~pi619 & n21636;
  assign n21772 = pi1159 & ~n21771;
  assign n21773 = ~n21770 & n21772;
  assign n21774 = ~n21769 & ~n21773;
  assign n21775 = pi789 & ~n21774;
  assign n21776 = ~n21765 & ~n21775;
  assign n21777 = ~n8595 & n21776;
  assign n21778 = n8595 & n21636;
  assign n21779 = ~n21777 & ~n21778;
  assign n21780 = ~n8334 & ~n21779;
  assign n21781 = n8334 & n21636;
  assign n21782 = ~n21780 & ~n21781;
  assign n21783 = ~n8376 & ~n21782;
  assign n21784 = n8376 & n21636;
  assign n21785 = n8376 & ~n21636;
  assign n21786 = ~n8376 & n21782;
  assign n21787 = ~n21785 & ~n21786;
  assign n21788 = ~n21783 & ~n21784;
  assign n21789 = pi644 & n63560;
  assign n21790 = ~pi644 & n21636;
  assign n21791 = ~pi715 & ~n21790;
  assign n21792 = ~n21789 & n21791;
  assign n21793 = pi1160 & ~n21792;
  assign n21794 = ~n21720 & n21793;
  assign n21795 = pi644 & n21718;
  assign n21796 = ~pi715 & ~n21795;
  assign n21797 = ~pi644 & n63560;
  assign n21798 = pi644 & n21636;
  assign n21799 = pi715 & ~n21798;
  assign n21800 = ~n21797 & n21799;
  assign n21801 = ~pi1160 & ~n21800;
  assign n21802 = ~n21796 & n21801;
  assign n21803 = ~n21794 & ~n21802;
  assign n21804 = pi790 & ~n21803;
  assign n21805 = ~pi644 & n21801;
  assign n21806 = pi644 & n21793;
  assign n21807 = n14029 & ~n21792;
  assign n21808 = pi790 & ~n63561;
  assign n21809 = ~n21805 & n21808;
  assign n21810 = ~n63052 & n21779;
  assign n21811 = n8331 & ~n21693;
  assign n21812 = ~pi629 & n63557;
  assign n21813 = pi629 & n21699;
  assign n21814 = ~n63562 & ~n21813;
  assign n21815 = ~n21810 & n21814;
  assign n21816 = pi792 & ~n21815;
  assign n21817 = n12979 & n21776;
  assign n21818 = ~pi641 & n63555;
  assign n21819 = pi641 & ~n21636;
  assign n21820 = n8417 & ~n21819;
  assign n21821 = ~n21818 & n21820;
  assign n21822 = pi641 & n63555;
  assign n21823 = ~pi641 & ~n21636;
  assign n21824 = n8416 & ~n21823;
  assign n21825 = ~n21822 & n21824;
  assign n21826 = ~n21821 & ~n21825;
  assign n21827 = ~n21817 & n21826;
  assign n21828 = pi788 & ~n21827;
  assign n21829 = pi619 & n63554;
  assign n21830 = ~pi1159 & ~n21829;
  assign n21831 = ~pi648 & ~n21773;
  assign n21832 = ~n21830 & n21831;
  assign n21833 = ~pi619 & n63554;
  assign n21834 = pi1159 & ~n21833;
  assign n21835 = pi648 & ~n21834;
  assign n21836 = pi648 & ~n21769;
  assign n21837 = ~n21834 & n21836;
  assign n21838 = ~n21769 & n21835;
  assign n21839 = ~n21832 & ~n63563;
  assign n21840 = pi789 & ~n21839;
  assign n21841 = pi618 & ~n63553;
  assign n21842 = ~pi1154 & ~n21841;
  assign n21843 = ~pi627 & ~n21757;
  assign n21844 = ~n21842 & n21843;
  assign n21845 = ~pi618 & ~n63553;
  assign n21846 = pi1154 & ~n21845;
  assign n21847 = pi627 & ~n21761;
  assign n21848 = ~n21846 & n21847;
  assign n21849 = ~n21844 & ~n21848;
  assign n21850 = pi781 & ~n21849;
  assign n21851 = ~pi618 & n21843;
  assign n21852 = pi618 & n21847;
  assign n21853 = pi781 & ~n21852;
  assign n21854 = ~n21851 & n21853;
  assign n21855 = ~pi188 & n10353;
  assign n21856 = pi188 & n10355;
  assign n21857 = pi768 & ~n10357;
  assign n21858 = ~n21856 & n21857;
  assign n21859 = ~n21855 & n21858;
  assign n21860 = pi188 & n10363;
  assign n21861 = ~pi188 & ~n62980;
  assign n21862 = ~pi768 & ~n21861;
  assign n21863 = ~n21860 & n21862;
  assign n21864 = pi705 & ~n21863;
  assign n21865 = ~n21859 & n21864;
  assign n21866 = ~pi705 & ~n63559;
  assign n21867 = n62765 & ~n21866;
  assign n21868 = n62765 & ~n21865;
  assign n21869 = ~n21866 & n21868;
  assign n21870 = ~n21865 & n21867;
  assign n21871 = ~n21638 & ~n63564;
  assign n21872 = ~pi625 & n21871;
  assign n21873 = pi625 & n21737;
  assign n21874 = ~pi1153 & ~n21873;
  assign n21875 = ~n21872 & n21874;
  assign n21876 = ~pi608 & ~n21656;
  assign n21877 = ~n21875 & n21876;
  assign n21878 = pi625 & n21871;
  assign n21879 = ~pi625 & n21737;
  assign n21880 = pi1153 & ~n21879;
  assign n21881 = ~n21878 & n21880;
  assign n21882 = pi608 & ~n21660;
  assign n21883 = ~n21881 & n21882;
  assign n21884 = ~n21877 & ~n21883;
  assign n21885 = pi778 & ~n21884;
  assign n21886 = ~pi778 & n21871;
  assign n21887 = ~pi778 & ~n21871;
  assign n21888 = pi778 & ~n21883;
  assign n21889 = ~n21877 & n21888;
  assign n21890 = ~n21887 & ~n21889;
  assign n21891 = ~n21885 & ~n21886;
  assign n21892 = ~pi785 & ~n63565;
  assign n21893 = ~pi609 & n63565;
  assign n21894 = pi609 & n21663;
  assign n21895 = ~pi1155 & ~n21894;
  assign n21896 = ~n21893 & n21895;
  assign n21897 = ~pi660 & ~n21745;
  assign n21898 = ~n21896 & n21897;
  assign n21899 = pi609 & n63565;
  assign n21900 = ~pi609 & n21663;
  assign n21901 = pi1155 & ~n21900;
  assign n21902 = ~n21899 & n21901;
  assign n21903 = pi660 & ~n21749;
  assign n21904 = ~n21902 & n21903;
  assign n21905 = pi785 & ~n21904;
  assign n21906 = ~n21898 & n21905;
  assign n21907 = ~n21898 & ~n21904;
  assign n21908 = pi785 & ~n21907;
  assign n21909 = ~pi785 & n63565;
  assign n21910 = ~n21908 & ~n21909;
  assign n21911 = ~n21892 & ~n21906;
  assign n21912 = ~n21854 & ~n63566;
  assign n21913 = pi618 & ~n63566;
  assign n21914 = n21846 & ~n21913;
  assign n21915 = n21847 & ~n21914;
  assign n21916 = ~n21844 & ~n21915;
  assign n21917 = pi781 & ~n21916;
  assign n21918 = pi781 & ~n21851;
  assign n21919 = ~n63566 & ~n21918;
  assign n21920 = ~n21917 & ~n21919;
  assign n21921 = ~pi618 & ~n63566;
  assign n21922 = n21842 & ~n21921;
  assign n21923 = n21843 & ~n21922;
  assign n21924 = ~n21915 & ~n21923;
  assign n21925 = pi781 & ~n21924;
  assign n21926 = ~pi781 & ~n63566;
  assign n21927 = ~n21925 & ~n21926;
  assign n21928 = ~n21850 & ~n21912;
  assign n21929 = ~pi619 & n21831;
  assign n21930 = pi619 & n21836;
  assign n21931 = n11422 & ~n21769;
  assign n21932 = pi789 & ~n63568;
  assign n21933 = ~n21929 & n21932;
  assign n21934 = ~n63567 & ~n21933;
  assign n21935 = ~pi619 & ~n63567;
  assign n21936 = n21830 & ~n21935;
  assign n21937 = n21831 & ~n21936;
  assign n21938 = pi619 & ~n63567;
  assign n21939 = n21834 & ~n21938;
  assign n21940 = n21836 & ~n21939;
  assign n21941 = ~n21937 & ~n21940;
  assign n21942 = pi789 & ~n21941;
  assign n21943 = ~pi789 & ~n63567;
  assign n21944 = ~n21942 & ~n21943;
  assign n21945 = ~n21840 & ~n21934;
  assign n21946 = n62894 & ~n63569;
  assign n21947 = ~n63030 & ~n21946;
  assign n21948 = ~n63030 & ~n21828;
  assign n21949 = ~n21946 & n21948;
  assign n21950 = ~n21828 & n21947;
  assign n21951 = ~pi788 & n63569;
  assign n21952 = ~pi626 & n63569;
  assign n21953 = pi626 & n63555;
  assign n21954 = ~pi641 & ~n21953;
  assign n21955 = ~n21952 & n21954;
  assign n21956 = ~pi626 & ~n21776;
  assign n21957 = pi626 & ~n21636;
  assign n21958 = pi641 & ~n21957;
  assign n21959 = ~n21956 & n21958;
  assign n21960 = ~pi1158 & ~n21959;
  assign n21961 = ~n21955 & n21960;
  assign n21962 = pi626 & n63569;
  assign n21963 = ~pi626 & n63555;
  assign n21964 = pi641 & ~n21963;
  assign n21965 = ~n21962 & n21964;
  assign n21966 = pi626 & ~n21776;
  assign n21967 = ~pi626 & ~n21636;
  assign n21968 = ~pi641 & ~n21967;
  assign n21969 = ~n21966 & n21968;
  assign n21970 = pi1158 & ~n21969;
  assign n21971 = ~n21965 & n21970;
  assign n21972 = ~n21961 & ~n21971;
  assign n21973 = pi788 & ~n21972;
  assign n21974 = ~n21951 & ~n21973;
  assign n21975 = ~pi628 & n21974;
  assign n21976 = pi628 & ~n21779;
  assign n21977 = ~pi1156 & ~n21976;
  assign n21978 = ~n21975 & n21977;
  assign n21979 = ~pi629 & ~n63557;
  assign n21980 = ~n21978 & n21979;
  assign n21981 = pi628 & n21974;
  assign n21982 = ~pi628 & ~n21779;
  assign n21983 = pi1156 & ~n21982;
  assign n21984 = ~n21981 & n21983;
  assign n21985 = pi629 & ~n21699;
  assign n21986 = ~n21984 & n21985;
  assign n21987 = ~n21980 & ~n21986;
  assign n21988 = pi792 & ~n21987;
  assign n21989 = ~pi792 & n21974;
  assign n21990 = ~n21988 & ~n21989;
  assign n21991 = ~n21816 & ~n63570;
  assign n21992 = ~n8651 & n63571;
  assign n21993 = ~n8413 & n21782;
  assign n21994 = n8373 & ~n21709;
  assign n21995 = ~pi630 & n63558;
  assign n21996 = pi630 & n21715;
  assign n21997 = ~n63572 & ~n21996;
  assign n21998 = ~n21993 & ~n21996;
  assign n21999 = ~n63572 & n21998;
  assign n22000 = ~n21993 & n21997;
  assign n22001 = pi787 & ~n63573;
  assign n22002 = ~n62896 & n63571;
  assign n22003 = ~pi647 & ~n63571;
  assign n22004 = pi647 & ~n21782;
  assign n22005 = ~pi1157 & ~n22004;
  assign n22006 = ~n22003 & n22005;
  assign n22007 = ~pi630 & ~n63558;
  assign n22008 = ~n22006 & n22007;
  assign n22009 = pi647 & ~n63571;
  assign n22010 = ~pi647 & ~n21782;
  assign n22011 = pi1157 & ~n22010;
  assign n22012 = ~n22009 & n22011;
  assign n22013 = pi630 & ~n21715;
  assign n22014 = ~n22012 & n22013;
  assign n22015 = ~n22008 & ~n22014;
  assign n22016 = n63573 & ~n22002;
  assign n22017 = pi787 & n63574;
  assign n22018 = ~pi787 & n63571;
  assign n22019 = ~n22017 & ~n22018;
  assign n22020 = pi787 & ~n63574;
  assign n22021 = ~pi787 & ~n63571;
  assign n22022 = ~n22020 & ~n22021;
  assign n22023 = ~n21992 & ~n22001;
  assign n22024 = ~n21809 & n63575;
  assign n22025 = ~pi644 & n63575;
  assign n22026 = n21796 & ~n22025;
  assign n22027 = n21801 & ~n22026;
  assign n22028 = ~n21794 & ~n22027;
  assign n22029 = pi790 & ~n22028;
  assign n22030 = ~n21808 & n63575;
  assign n22031 = ~n22029 & ~n22030;
  assign n22032 = ~n21804 & ~n22024;
  assign n22033 = pi644 & n63575;
  assign n22034 = n21720 & ~n22033;
  assign n22035 = n21793 & ~n22034;
  assign n22036 = pi790 & ~n22027;
  assign n22037 = pi790 & ~n22035;
  assign n22038 = ~n22027 & n22037;
  assign n22039 = ~n22035 & n22036;
  assign n22040 = ~pi790 & ~n63575;
  assign n22041 = n62455 & ~n22040;
  assign n22042 = ~n63577 & n22041;
  assign n22043 = n62455 & ~n63576;
  assign n22044 = ~pi188 & ~n62455;
  assign n22045 = ~pi832 & ~n22044;
  assign n22046 = ~n63578 & n22045;
  assign po345 = ~n21635 & ~n22046;
  assign n22048 = pi189 & ~n62765;
  assign n22049 = ~pi772 & ~n7143;
  assign n22050 = pi772 & ~n62801;
  assign n22051 = ~n22049 & ~n22050;
  assign n22052 = pi39 & ~n22051;
  assign n22053 = pi772 & n62793;
  assign n22054 = ~pi772 & ~n62781;
  assign n22055 = ~pi39 & ~n22054;
  assign n22056 = ~n22053 & n22055;
  assign n22057 = ~n22052 & ~n22056;
  assign n22058 = pi189 & ~n22057;
  assign n22059 = ~pi189 & pi772;
  assign n22060 = n7351 & n22059;
  assign n22061 = ~n22058 & ~n22060;
  assign n22062 = ~pi38 & ~n22061;
  assign n22063 = pi772 & n7187;
  assign n22064 = n7357 & ~n22063;
  assign n22065 = ~pi189 & ~n7357;
  assign n22066 = pi38 & ~n22065;
  assign n22067 = pi38 & ~n22064;
  assign n22068 = ~n22065 & n22067;
  assign n22069 = ~n22064 & n22066;
  assign n22070 = ~n22062 & ~n63579;
  assign n22071 = n62765 & ~n22070;
  assign n22072 = ~n22048 & ~n22071;
  assign n22073 = ~n8135 & ~n22072;
  assign n22074 = pi189 & ~n8098;
  assign n22075 = n8135 & n22074;
  assign n22076 = n8135 & ~n22074;
  assign n22077 = ~n8135 & n22072;
  assign n22078 = ~n22076 & ~n22077;
  assign n22079 = ~n22073 & ~n22075;
  assign n22080 = ~pi785 & n63580;
  assign n22081 = pi609 & ~n63580;
  assign n22082 = ~pi609 & ~n22074;
  assign n22083 = pi1155 & ~n22082;
  assign n22084 = ~n22081 & n22083;
  assign n22085 = ~pi609 & ~n63580;
  assign n22086 = pi609 & ~n22074;
  assign n22087 = ~pi1155 & ~n22086;
  assign n22088 = ~n22085 & n22087;
  assign n22089 = ~n22084 & ~n22088;
  assign n22090 = pi785 & ~n22089;
  assign n22091 = ~n22080 & ~n22090;
  assign n22092 = ~pi781 & ~n22091;
  assign n22093 = pi618 & n22091;
  assign n22094 = ~pi618 & ~n22074;
  assign n22095 = pi1154 & ~n22094;
  assign n22096 = ~n22093 & n22095;
  assign n22097 = ~pi618 & n22091;
  assign n22098 = pi618 & ~n22074;
  assign n22099 = ~pi1154 & ~n22098;
  assign n22100 = ~n22097 & n22099;
  assign n22101 = ~n22096 & ~n22100;
  assign n22102 = pi781 & ~n22101;
  assign n22103 = ~n22092 & ~n22102;
  assign n22104 = ~pi789 & ~n22103;
  assign n22105 = ~pi619 & n22103;
  assign n22106 = pi619 & ~n22074;
  assign n22107 = ~pi1159 & ~n22106;
  assign n22108 = ~n22105 & n22107;
  assign n22109 = pi619 & n22103;
  assign n22110 = ~pi619 & ~n22074;
  assign n22111 = pi1159 & ~n22110;
  assign n22112 = ~n22109 & n22111;
  assign n22113 = ~n22108 & ~n22112;
  assign n22114 = pi789 & ~n22113;
  assign n22115 = ~n22104 & ~n22114;
  assign n22116 = ~n8595 & ~n22115;
  assign n22117 = n8595 & n22074;
  assign n22118 = ~n22116 & ~n22117;
  assign n22119 = ~n8334 & ~n22118;
  assign n22120 = n8334 & n22074;
  assign n22121 = ~n22119 & ~n22120;
  assign n22122 = ~n8376 & ~n22121;
  assign n22123 = n8376 & n22074;
  assign n22124 = n8376 & ~n22074;
  assign n22125 = ~n8376 & n22121;
  assign n22126 = ~n22124 & ~n22125;
  assign n22127 = ~n22122 & ~n22123;
  assign n22128 = ~pi644 & ~n63581;
  assign n22129 = pi644 & ~n22074;
  assign n22130 = pi715 & ~n22129;
  assign n22131 = ~n22128 & n22130;
  assign n22132 = n8257 & ~n22074;
  assign n22133 = n62880 & ~n22074;
  assign n22134 = pi727 & n62765;
  assign n22135 = n10997 & ~n22065;
  assign n22136 = pi189 & ~n8009;
  assign n22137 = ~pi189 & ~n62874;
  assign n22138 = ~pi38 & ~n22137;
  assign n22139 = ~n22136 & n22138;
  assign n22140 = ~n22135 & ~n22139;
  assign n22141 = n22134 & ~n22140;
  assign n22142 = n22074 & ~n22134;
  assign n22143 = ~n22074 & ~n22134;
  assign n22144 = n22134 & ~n22135;
  assign n22145 = ~n22139 & n22144;
  assign n22146 = ~n22143 & ~n22145;
  assign n22147 = ~n22141 & ~n22142;
  assign n22148 = ~pi778 & n63582;
  assign n22149 = pi625 & ~n63582;
  assign n22150 = ~pi625 & ~n22074;
  assign n22151 = pi1153 & ~n22150;
  assign n22152 = ~n22149 & n22151;
  assign n22153 = ~pi625 & ~n63582;
  assign n22154 = pi625 & ~n22074;
  assign n22155 = ~pi1153 & ~n22154;
  assign n22156 = ~n22153 & n22155;
  assign n22157 = ~n22152 & ~n22156;
  assign n22158 = pi778 & ~n22157;
  assign n22159 = ~n22148 & ~n22158;
  assign n22160 = ~n62880 & n22159;
  assign n22161 = ~n62880 & ~n22159;
  assign n22162 = n62880 & n22074;
  assign n22163 = ~n22161 & ~n22162;
  assign n22164 = ~n22133 & ~n22160;
  assign n22165 = ~n62882 & ~n63583;
  assign n22166 = n62882 & n22074;
  assign n22167 = n62882 & ~n22074;
  assign n22168 = ~n62882 & n63583;
  assign n22169 = ~n22167 & ~n22168;
  assign n22170 = ~n22165 & ~n22166;
  assign n22171 = ~n8257 & ~n63584;
  assign n22172 = ~n8257 & n63584;
  assign n22173 = n8257 & n22074;
  assign n22174 = ~n22172 & ~n22173;
  assign n22175 = ~n22132 & ~n22171;
  assign n22176 = ~n8303 & ~n63585;
  assign n22177 = n8303 & n22074;
  assign n22178 = n8303 & ~n22074;
  assign n22179 = ~n8303 & n63585;
  assign n22180 = ~n22178 & ~n22179;
  assign n22181 = ~n22176 & ~n22177;
  assign n22182 = pi628 & ~n63586;
  assign n22183 = ~pi628 & ~n22074;
  assign n22184 = pi1156 & ~n22183;
  assign n22185 = pi628 & n63586;
  assign n22186 = ~pi628 & n22074;
  assign n22187 = ~n22185 & ~n22186;
  assign n22188 = pi1156 & ~n22187;
  assign n22189 = ~n22182 & n22184;
  assign n22190 = ~pi628 & ~n63586;
  assign n22191 = pi628 & ~n22074;
  assign n22192 = ~pi1156 & ~n22191;
  assign n22193 = ~n22190 & n22192;
  assign n22194 = ~n22190 & ~n22191;
  assign n22195 = ~pi1156 & ~n22194;
  assign n22196 = pi1156 & n22187;
  assign n22197 = ~n22195 & ~n22196;
  assign n22198 = ~n63587 & ~n22193;
  assign n22199 = pi792 & n63588;
  assign n22200 = ~pi792 & n63586;
  assign n22201 = pi792 & ~n63588;
  assign n22202 = ~pi792 & ~n63586;
  assign n22203 = ~n22201 & ~n22202;
  assign n22204 = ~n22199 & ~n22200;
  assign n22205 = ~pi787 & n63589;
  assign n22206 = pi647 & ~n63589;
  assign n22207 = ~pi647 & ~n22074;
  assign n22208 = pi1157 & ~n22207;
  assign n22209 = pi647 & n63589;
  assign n22210 = ~pi647 & n22074;
  assign n22211 = ~n22209 & ~n22210;
  assign n22212 = pi1157 & ~n22211;
  assign n22213 = ~n22206 & n22208;
  assign n22214 = ~pi647 & ~n63589;
  assign n22215 = pi647 & ~n22074;
  assign n22216 = ~pi1157 & ~n22215;
  assign n22217 = ~n22214 & n22216;
  assign n22218 = ~n63590 & ~n22217;
  assign n22219 = pi787 & ~n22218;
  assign n22220 = ~n22205 & ~n22219;
  assign n22221 = n15025 & ~n22220;
  assign n22222 = ~pi1160 & ~n22221;
  assign n22223 = ~n22131 & n22222;
  assign n22224 = pi644 & ~n63581;
  assign n22225 = ~pi644 & ~n22074;
  assign n22226 = ~pi715 & ~n22225;
  assign n22227 = ~n22224 & n22226;
  assign n22228 = n14949 & ~n22220;
  assign n22229 = pi1160 & ~n22228;
  assign n22230 = ~n22227 & n22229;
  assign n22231 = pi790 & ~n22230;
  assign n22232 = ~n22223 & n22231;
  assign n22233 = ~n8413 & ~n22121;
  assign n22234 = n8373 & ~n22211;
  assign n22235 = pi630 & n22217;
  assign n22236 = ~n22234 & ~n22235;
  assign n22237 = ~n22233 & n22236;
  assign n22238 = pi787 & ~n22237;
  assign n22239 = ~n63052 & ~n22118;
  assign n22240 = n8331 & ~n22187;
  assign n22241 = n8332 & n22194;
  assign n22242 = pi629 & n22193;
  assign n22243 = ~n22240 & ~n63591;
  assign n22244 = ~n22239 & n22243;
  assign n22245 = pi792 & ~n22244;
  assign n22246 = pi619 & ~n63584;
  assign n22247 = ~pi1159 & ~n22246;
  assign n22248 = ~pi648 & ~n22112;
  assign n22249 = ~n22247 & n22248;
  assign n22250 = ~pi619 & ~n63584;
  assign n22251 = pi1159 & ~n22250;
  assign n22252 = pi648 & ~n22251;
  assign n22253 = pi648 & ~n22108;
  assign n22254 = ~n22251 & n22253;
  assign n22255 = ~n22108 & n22252;
  assign n22256 = ~n22249 & ~n63592;
  assign n22257 = pi789 & ~n22256;
  assign n22258 = ~pi727 & n22062;
  assign n22259 = pi189 & ~n62821;
  assign n22260 = ~pi189 & n7632;
  assign n22261 = ~pi772 & ~n22260;
  assign n22262 = ~n22259 & n22261;
  assign n22263 = ~pi189 & n7709;
  assign n22264 = pi189 & n62851;
  assign n22265 = pi772 & ~n22264;
  assign n22266 = ~n22263 & n22265;
  assign n22267 = pi39 & ~n22266;
  assign n22268 = ~n22262 & n22267;
  assign n22269 = pi189 & ~n7832;
  assign n22270 = ~pi189 & ~n7855;
  assign n22271 = ~pi772 & ~n22270;
  assign n22272 = ~pi772 & ~n22269;
  assign n22273 = ~n22270 & n22272;
  assign n22274 = ~n22269 & n22271;
  assign n22275 = pi189 & n7861;
  assign n22276 = ~pi189 & n7868;
  assign n22277 = pi772 & ~n22276;
  assign n22278 = ~n22275 & n22277;
  assign n22279 = ~n63593 & ~n22278;
  assign n22280 = ~pi39 & ~n22279;
  assign n22281 = ~pi38 & ~n22280;
  assign n22282 = ~n22268 & n22281;
  assign n22283 = pi727 & ~n8793;
  assign n22284 = pi189 & n62821;
  assign n22285 = ~pi189 & ~n7632;
  assign n22286 = ~pi772 & ~n22285;
  assign n22287 = ~n22284 & n22286;
  assign n22288 = ~pi189 & ~n7709;
  assign n22289 = pi189 & ~n62851;
  assign n22290 = pi772 & ~n22289;
  assign n22291 = ~n22288 & n22290;
  assign n22292 = pi39 & ~n22291;
  assign n22293 = ~n22287 & n22292;
  assign n22294 = ~pi39 & ~n22278;
  assign n22295 = ~n63593 & n22294;
  assign n22296 = ~pi38 & ~n22295;
  assign n22297 = ~n22293 & n22296;
  assign n22298 = ~n10357 & ~n22297;
  assign n22299 = pi727 & ~n22298;
  assign n22300 = ~n22282 & n22283;
  assign n22301 = ~n63579 & ~n63594;
  assign n22302 = ~n22258 & n22301;
  assign n22303 = ~pi727 & n22070;
  assign n22304 = pi727 & ~n10357;
  assign n22305 = ~n63579 & n22304;
  assign n22306 = ~n22297 & n22305;
  assign n22307 = n62765 & ~n22306;
  assign n22308 = ~n22303 & n22307;
  assign n22309 = n62765 & ~n22302;
  assign n22310 = ~n22048 & ~n63595;
  assign n22311 = ~pi625 & n22310;
  assign n22312 = pi625 & n22072;
  assign n22313 = ~pi1153 & ~n22312;
  assign n22314 = ~n22311 & n22313;
  assign n22315 = ~pi608 & ~n22152;
  assign n22316 = ~n22314 & n22315;
  assign n22317 = pi625 & n22310;
  assign n22318 = ~pi625 & n22072;
  assign n22319 = pi1153 & ~n22318;
  assign n22320 = ~n22317 & n22319;
  assign n22321 = pi608 & ~n22156;
  assign n22322 = ~n22320 & n22321;
  assign n22323 = ~n22316 & ~n22322;
  assign n22324 = pi778 & ~n22323;
  assign n22325 = ~pi778 & n22310;
  assign n22326 = ~n22324 & ~n22325;
  assign n22327 = ~pi609 & ~n22326;
  assign n22328 = pi609 & n22159;
  assign n22329 = ~pi1155 & ~n22328;
  assign n22330 = ~n22327 & n22329;
  assign n22331 = ~pi660 & ~n22084;
  assign n22332 = ~n22330 & n22331;
  assign n22333 = pi609 & ~n22326;
  assign n22334 = ~pi609 & n22159;
  assign n22335 = pi1155 & ~n22334;
  assign n22336 = ~n22333 & n22335;
  assign n22337 = pi660 & ~n22088;
  assign n22338 = ~n22336 & n22337;
  assign n22339 = ~n22332 & ~n22338;
  assign n22340 = pi785 & ~n22339;
  assign n22341 = ~pi785 & ~n22326;
  assign n22342 = ~n22340 & ~n22341;
  assign n22343 = pi618 & ~n22342;
  assign n22344 = ~pi618 & n63583;
  assign n22345 = pi1154 & ~n22344;
  assign n22346 = ~n22343 & n22345;
  assign n22347 = pi627 & ~n22100;
  assign n22348 = ~n22346 & n22347;
  assign n22349 = ~pi618 & ~n22342;
  assign n22350 = pi618 & n63583;
  assign n22351 = ~pi1154 & ~n22350;
  assign n22352 = ~n22349 & n22351;
  assign n22353 = ~pi627 & ~n22096;
  assign n22354 = ~n22352 & n22353;
  assign n22355 = pi781 & ~n22354;
  assign n22356 = ~n22348 & n22355;
  assign n22357 = ~pi619 & n22248;
  assign n22358 = pi619 & n22253;
  assign n22359 = n11422 & ~n22108;
  assign n22360 = pi789 & ~n63596;
  assign n22361 = ~n22357 & n22360;
  assign n22362 = ~pi781 & n22342;
  assign n22363 = ~n22361 & ~n22362;
  assign n22364 = ~n22356 & n22363;
  assign n22365 = ~n22348 & ~n22354;
  assign n22366 = pi781 & ~n22365;
  assign n22367 = ~pi781 & ~n22342;
  assign n22368 = ~n22366 & ~n22367;
  assign n22369 = ~pi619 & ~n22368;
  assign n22370 = n22247 & ~n22369;
  assign n22371 = n22248 & ~n22370;
  assign n22372 = pi619 & ~n22368;
  assign n22373 = n22251 & ~n22372;
  assign n22374 = n22253 & ~n22373;
  assign n22375 = ~n22371 & ~n22374;
  assign n22376 = pi789 & ~n22375;
  assign n22377 = ~pi789 & ~n22368;
  assign n22378 = ~n22376 & ~n22377;
  assign n22379 = ~n22257 & ~n22364;
  assign n22380 = n62894 & ~n63597;
  assign n22381 = n12979 & n22115;
  assign n22382 = ~pi641 & ~n63585;
  assign n22383 = pi641 & n22074;
  assign n22384 = n8417 & ~n22383;
  assign n22385 = ~n22382 & n22384;
  assign n22386 = pi641 & ~n63585;
  assign n22387 = ~pi641 & n22074;
  assign n22388 = n8416 & ~n22387;
  assign n22389 = ~n22386 & n22388;
  assign n22390 = ~n22385 & ~n22389;
  assign n22391 = ~n22381 & n22390;
  assign n22392 = pi788 & ~n22391;
  assign n22393 = ~n63030 & ~n22392;
  assign n22394 = ~n22380 & n22393;
  assign n22395 = ~pi788 & n63597;
  assign n22396 = ~pi626 & n63597;
  assign n22397 = pi626 & ~n63585;
  assign n22398 = ~pi641 & ~n22397;
  assign n22399 = ~n22396 & n22398;
  assign n22400 = ~pi626 & ~n22115;
  assign n22401 = pi626 & n22074;
  assign n22402 = pi641 & ~n22401;
  assign n22403 = ~n22400 & n22402;
  assign n22404 = ~pi1158 & ~n22403;
  assign n22405 = ~n22399 & n22404;
  assign n22406 = pi626 & n63597;
  assign n22407 = ~pi626 & ~n63585;
  assign n22408 = pi641 & ~n22407;
  assign n22409 = ~n22406 & n22408;
  assign n22410 = pi626 & ~n22115;
  assign n22411 = ~pi626 & n22074;
  assign n22412 = ~pi641 & ~n22411;
  assign n22413 = ~n22410 & n22412;
  assign n22414 = pi1158 & ~n22413;
  assign n22415 = ~n22409 & n22414;
  assign n22416 = ~n22405 & ~n22415;
  assign n22417 = pi788 & ~n22416;
  assign n22418 = ~n22395 & ~n22417;
  assign n22419 = ~pi628 & n22418;
  assign n22420 = pi628 & n22118;
  assign n22421 = ~pi1156 & ~n22420;
  assign n22422 = ~n22419 & n22421;
  assign n22423 = ~pi629 & ~n63587;
  assign n22424 = ~n22422 & n22423;
  assign n22425 = pi628 & n22418;
  assign n22426 = ~pi628 & n22118;
  assign n22427 = pi1156 & ~n22426;
  assign n22428 = ~n22425 & n22427;
  assign n22429 = pi629 & ~n22193;
  assign n22430 = ~n22428 & n22429;
  assign n22431 = ~n22424 & ~n22430;
  assign n22432 = pi792 & ~n22431;
  assign n22433 = ~pi792 & n22418;
  assign n22434 = ~n22432 & ~n22433;
  assign n22435 = ~n22245 & ~n22394;
  assign n22436 = ~n8651 & n63598;
  assign n22437 = n8651 & n22237;
  assign n22438 = ~n22238 & ~n63598;
  assign n22439 = ~n22437 & ~n22438;
  assign n22440 = ~pi647 & ~n63598;
  assign n22441 = pi647 & n22121;
  assign n22442 = ~pi1157 & ~n22441;
  assign n22443 = ~n22440 & n22442;
  assign n22444 = ~pi630 & ~n63590;
  assign n22445 = ~n22443 & n22444;
  assign n22446 = pi647 & ~n63598;
  assign n22447 = ~pi647 & n22121;
  assign n22448 = pi1157 & ~n22447;
  assign n22449 = ~n22446 & n22448;
  assign n22450 = pi630 & ~n22217;
  assign n22451 = ~n22449 & n22450;
  assign n22452 = ~n22445 & ~n22451;
  assign n22453 = pi787 & ~n22452;
  assign n22454 = ~pi787 & ~n63598;
  assign n22455 = ~n22453 & ~n22454;
  assign n22456 = ~n22238 & ~n22436;
  assign n22457 = ~n11547 & n63599;
  assign n22458 = n3475 & ~n22457;
  assign n22459 = ~pi644 & ~n63599;
  assign n22460 = pi644 & n22220;
  assign n22461 = ~pi715 & ~n22460;
  assign n22462 = ~n22459 & n22461;
  assign n22463 = ~pi1160 & ~n22131;
  assign n22464 = ~n22462 & n22463;
  assign n22465 = ~pi644 & n22220;
  assign n22466 = pi715 & ~n22465;
  assign n22467 = pi1160 & ~n22227;
  assign n22468 = ~n22466 & n22467;
  assign n22469 = ~n22464 & ~n22468;
  assign n22470 = pi790 & ~n22469;
  assign n22471 = pi644 & n22467;
  assign n22472 = pi790 & ~n22471;
  assign n22473 = ~n63599 & ~n22472;
  assign n22474 = ~n22470 & ~n22473;
  assign n22475 = n3475 & ~n22474;
  assign n22476 = pi644 & ~n63599;
  assign n22477 = n22466 & ~n22476;
  assign n22478 = n22467 & ~n22477;
  assign n22479 = pi790 & ~n22464;
  assign n22480 = pi790 & ~n22478;
  assign n22481 = ~n22464 & n22480;
  assign n22482 = ~n22478 & n22479;
  assign n22483 = ~pi790 & n63599;
  assign n22484 = n3475 & ~n22483;
  assign n22485 = ~n63601 & n22484;
  assign n22486 = ~n22232 & n22458;
  assign n22487 = ~pi189 & ~n3475;
  assign n22488 = ~pi57 & ~n22487;
  assign n22489 = ~n63600 & n22488;
  assign n22490 = pi57 & pi189;
  assign n22491 = ~pi832 & ~n22490;
  assign n22492 = ~n22489 & n22491;
  assign n22493 = pi727 & n7564;
  assign n22494 = pi727 & n7565;
  assign n22495 = ~n7187 & n22493;
  assign n22496 = pi625 & n22493;
  assign n22497 = ~n7187 & n22496;
  assign n22498 = pi625 & n63602;
  assign n22499 = pi189 & ~n2923;
  assign n22500 = pi772 & n7316;
  assign n22501 = ~n22499 & ~n22500;
  assign n22502 = ~n63602 & n22501;
  assign n22503 = ~n63603 & ~n22502;
  assign n22504 = ~pi1153 & ~n22503;
  assign n22505 = pi1153 & ~n22499;
  assign n22506 = ~n22496 & n22505;
  assign n22507 = ~pi608 & ~n22506;
  assign n22508 = ~n22504 & n22507;
  assign n22509 = pi1153 & n22501;
  assign n22510 = ~n22500 & n22505;
  assign n22511 = ~n63603 & n63604;
  assign n22512 = ~n22493 & ~n22499;
  assign n22513 = ~n22496 & ~n22512;
  assign n22514 = ~pi1153 & ~n22513;
  assign n22515 = pi608 & ~n22514;
  assign n22516 = pi608 & ~n22511;
  assign n22517 = ~n22514 & n22516;
  assign n22518 = ~n22511 & n22515;
  assign n22519 = ~n22508 & ~n63605;
  assign n22520 = pi778 & ~n22519;
  assign n22521 = ~pi778 & ~n22502;
  assign n22522 = ~n22520 & ~n22521;
  assign n22523 = ~pi609 & ~n22522;
  assign n22524 = ~pi778 & n22512;
  assign n22525 = ~n22506 & ~n22514;
  assign n22526 = pi778 & ~n22525;
  assign n22527 = ~n22524 & ~n22526;
  assign n22528 = pi609 & n22527;
  assign n22529 = ~pi1155 & ~n22528;
  assign n22530 = ~n22523 & n22529;
  assign n22531 = n8136 & n22500;
  assign n22532 = pi1155 & ~n22499;
  assign n22533 = ~n22531 & n22532;
  assign n22534 = ~pi660 & ~n22533;
  assign n22535 = ~n22530 & n22534;
  assign n22536 = pi609 & ~n22522;
  assign n22537 = ~pi609 & n22527;
  assign n22538 = pi1155 & ~n22537;
  assign n22539 = ~n22536 & n22538;
  assign n22540 = n8148 & n22500;
  assign n22541 = ~pi1155 & ~n22499;
  assign n22542 = ~n22540 & n22541;
  assign n22543 = pi660 & ~n22542;
  assign n22544 = ~n22539 & n22543;
  assign n22545 = ~n22535 & ~n22544;
  assign n22546 = pi785 & ~n22545;
  assign n22547 = ~pi785 & ~n22522;
  assign n22548 = ~n22546 & ~n22547;
  assign n22549 = pi618 & ~n22548;
  assign n22550 = ~n62880 & n22527;
  assign n22551 = ~n22499 & ~n22550;
  assign n22552 = ~pi618 & ~n22551;
  assign n22553 = pi1154 & ~n22552;
  assign n22554 = ~n22549 & n22553;
  assign n22555 = ~n63011 & n22500;
  assign n22556 = n11388 & n22555;
  assign n22557 = ~pi1154 & ~n22499;
  assign n22558 = ~n22556 & n22557;
  assign n22559 = pi627 & ~n22558;
  assign n22560 = ~n22554 & n22559;
  assign n22561 = ~pi618 & ~n22548;
  assign n22562 = pi618 & ~n22551;
  assign n22563 = ~pi1154 & ~n22562;
  assign n22564 = ~n22561 & n22563;
  assign n22565 = n11386 & n22555;
  assign n22566 = pi1154 & ~n22499;
  assign n22567 = ~n22565 & n22566;
  assign n22568 = ~pi627 & ~n22567;
  assign n22569 = ~n22564 & n22568;
  assign n22570 = ~n22560 & ~n22569;
  assign n22571 = pi781 & ~n22570;
  assign n22572 = ~pi781 & ~n22548;
  assign n22573 = ~n11434 & ~n22572;
  assign n22574 = ~n22571 & n22573;
  assign n22575 = n10106 & n22527;
  assign n22576 = ~n11431 & ~n22575;
  assign n22577 = n13305 & n22555;
  assign n22578 = ~n63012 & n22555;
  assign n22579 = ~n62884 & ~n22578;
  assign n22580 = ~n13309 & ~n22579;
  assign n22581 = n11438 & n22578;
  assign n22582 = n8254 & ~n22581;
  assign n22583 = n11447 & n22578;
  assign n22584 = n8253 & ~n22583;
  assign n22585 = ~n22582 & ~n22584;
  assign n22586 = ~n62884 & ~n22577;
  assign n22587 = ~n22576 & n63606;
  assign n22588 = pi789 & ~n22499;
  assign n22589 = ~n22587 & n22588;
  assign n22590 = n62894 & ~n22589;
  assign n22591 = ~n22574 & n22590;
  assign n22592 = ~n8257 & n22575;
  assign n22593 = ~n22499 & ~n22592;
  assign n22594 = n8417 & ~n22593;
  assign n22595 = n63013 & n22555;
  assign n22596 = pi626 & n22595;
  assign n22597 = ~n22499 & ~n22596;
  assign n22598 = pi1158 & ~n22597;
  assign n22599 = ~pi641 & ~n22598;
  assign n22600 = ~n22594 & n22599;
  assign n22601 = n8416 & ~n22593;
  assign n22602 = ~pi626 & n22595;
  assign n22603 = ~n22499 & ~n22602;
  assign n22604 = ~pi1158 & ~n22603;
  assign n22605 = pi641 & ~n22604;
  assign n22606 = ~n22601 & n22605;
  assign n22607 = pi788 & ~n22606;
  assign n22608 = pi788 & ~n22600;
  assign n22609 = ~n22606 & n22608;
  assign n22610 = ~n22600 & n22607;
  assign n22611 = ~n63030 & ~n63607;
  assign n22612 = ~n22591 & n22611;
  assign n22613 = ~n8595 & n22595;
  assign n22614 = n13344 & n22500;
  assign n22615 = ~pi629 & n63608;
  assign n22616 = pi628 & ~n22615;
  assign n22617 = ~n8303 & n22592;
  assign n22618 = n10207 & n22527;
  assign n22619 = pi629 & ~n63609;
  assign n22620 = ~pi628 & n63609;
  assign n22621 = pi629 & ~n22620;
  assign n22622 = pi628 & ~n63608;
  assign n22623 = ~n22621 & ~n22622;
  assign n22624 = ~n22616 & ~n22619;
  assign n22625 = ~pi1156 & ~n63610;
  assign n22626 = pi628 & n63609;
  assign n22627 = ~pi628 & ~n63608;
  assign n22628 = pi629 & ~n22627;
  assign n22629 = pi1156 & ~n22628;
  assign n22630 = ~n22626 & n22629;
  assign n22631 = ~n22625 & ~n22630;
  assign n22632 = pi792 & ~n22499;
  assign n22633 = ~n22631 & n22632;
  assign n22634 = ~n22612 & ~n22633;
  assign n22635 = ~n8651 & ~n22634;
  assign n22636 = ~n62892 & n63609;
  assign n22637 = ~pi630 & ~n22636;
  assign n22638 = pi647 & ~n22637;
  assign n22639 = ~n8334 & n63608;
  assign n22640 = pi630 & n22639;
  assign n22641 = pi1157 & ~n22640;
  assign n22642 = ~n22638 & n22641;
  assign n22643 = pi630 & ~n22636;
  assign n22644 = ~pi647 & ~n22643;
  assign n22645 = ~pi630 & n22639;
  assign n22646 = ~pi1157 & ~n22645;
  assign n22647 = pi647 & ~n22645;
  assign n22648 = ~n22643 & ~n22647;
  assign n22649 = ~pi1157 & ~n22648;
  assign n22650 = ~n22644 & n22646;
  assign n22651 = ~n22642 & ~n63611;
  assign n22652 = pi787 & ~n22499;
  assign n22653 = ~n22651 & n22652;
  assign n22654 = ~n11547 & ~n22653;
  assign n22655 = ~n22635 & n22654;
  assign n22656 = n11556 & n22636;
  assign n22657 = n11558 & n22595;
  assign n22658 = n13393 & n22555;
  assign n22659 = ~pi1160 & n63612;
  assign n22660 = ~n22499 & ~n22659;
  assign n22661 = n11540 & ~n22660;
  assign n22662 = pi1160 & n63612;
  assign n22663 = ~n22499 & ~n22662;
  assign n22664 = n11542 & ~n22663;
  assign n22665 = ~n22661 & ~n22664;
  assign n22666 = ~n22656 & n22665;
  assign n22667 = pi790 & ~n22666;
  assign n22668 = pi832 & ~n22667;
  assign n22669 = ~n22635 & ~n22653;
  assign n22670 = pi644 & n22669;
  assign n22671 = ~n10298 & n22636;
  assign n22672 = ~n22499 & ~n22671;
  assign n22673 = ~pi644 & ~n22672;
  assign n22674 = pi715 & ~n22673;
  assign n22675 = ~n22670 & n22674;
  assign n22676 = pi644 & n63612;
  assign n22677 = ~pi715 & ~n22499;
  assign n22678 = ~n22676 & n22677;
  assign n22679 = pi1160 & ~n22678;
  assign n22680 = ~n22675 & n22679;
  assign n22681 = ~pi644 & n22669;
  assign n22682 = pi644 & ~n22672;
  assign n22683 = ~pi715 & ~n22682;
  assign n22684 = ~n22681 & n22683;
  assign n22685 = ~pi644 & n63612;
  assign n22686 = pi715 & ~n22499;
  assign n22687 = ~n22685 & n22686;
  assign n22688 = ~pi1160 & ~n22687;
  assign n22689 = ~n22684 & n22688;
  assign n22690 = ~n22680 & ~n22689;
  assign n22691 = pi790 & ~n22690;
  assign n22692 = ~pi790 & n22669;
  assign n22693 = pi832 & ~n22692;
  assign n22694 = ~n22691 & n22693;
  assign n22695 = ~n22655 & n22668;
  assign po346 = ~n22492 & ~n63613;
  assign n22697 = ~pi190 & ~n2923;
  assign n22698 = pi763 & n7316;
  assign n22699 = ~n22697 & ~n22698;
  assign n22700 = ~n8420 & ~n22699;
  assign n22701 = ~pi785 & ~n22700;
  assign n22702 = n8148 & n22698;
  assign n22703 = n22700 & ~n22702;
  assign n22704 = pi1155 & ~n22703;
  assign n22705 = ~pi1155 & ~n22697;
  assign n22706 = ~n22702 & n22705;
  assign n22707 = ~n22704 & ~n22706;
  assign n22708 = pi785 & ~n22707;
  assign n22709 = ~n22701 & ~n22708;
  assign n22710 = ~pi781 & ~n22709;
  assign n22711 = ~n8435 & n22709;
  assign n22712 = pi1154 & ~n22711;
  assign n22713 = ~n8438 & n22709;
  assign n22714 = ~pi1154 & ~n22713;
  assign n22715 = ~n22712 & ~n22714;
  assign n22716 = pi781 & ~n22715;
  assign n22717 = ~n22710 & ~n22716;
  assign n22718 = ~pi789 & ~n22717;
  assign n22719 = ~n12612 & n22717;
  assign n22720 = pi1159 & ~n22719;
  assign n22721 = ~n12615 & n22717;
  assign n22722 = ~pi1159 & ~n22721;
  assign n22723 = ~n22720 & ~n22722;
  assign n22724 = pi789 & ~n22723;
  assign n22725 = ~n22718 & ~n22724;
  assign n22726 = ~n15298 & n22717;
  assign n22727 = ~n8595 & n63614;
  assign n22728 = n8595 & n22697;
  assign n22729 = ~n8595 & ~n63614;
  assign n22730 = n8595 & ~n22697;
  assign n22731 = ~n22729 & ~n22730;
  assign n22732 = ~n22727 & ~n22728;
  assign n22733 = ~n8334 & n63615;
  assign n22734 = n8334 & n22697;
  assign n22735 = ~n8413 & ~n22734;
  assign n22736 = ~n22733 & ~n22734;
  assign n22737 = ~n8413 & n22736;
  assign n22738 = ~n22733 & n22735;
  assign n22739 = pi699 & n7564;
  assign n22740 = ~n22697 & ~n22739;
  assign n22741 = ~pi778 & ~n22740;
  assign n22742 = ~pi625 & n22739;
  assign n22743 = ~n22740 & ~n22742;
  assign n22744 = pi1153 & ~n22743;
  assign n22745 = ~pi1153 & ~n22697;
  assign n22746 = ~n22742 & n22745;
  assign n22747 = pi778 & ~n22746;
  assign n22748 = ~n22744 & n22747;
  assign n22749 = ~n22741 & ~n22748;
  assign n22750 = ~n8490 & ~n22749;
  assign n22751 = ~n8492 & n22750;
  assign n22752 = ~n8494 & n22751;
  assign n22753 = ~n8496 & n22752;
  assign n22754 = ~n8508 & n22753;
  assign n22755 = pi647 & ~n22754;
  assign n22756 = ~pi647 & ~n22697;
  assign n22757 = ~n22755 & ~n22756;
  assign n22758 = n8373 & ~n22757;
  assign n22759 = ~pi647 & n22754;
  assign n22760 = pi647 & n22697;
  assign n22761 = ~pi1157 & ~n22760;
  assign n22762 = ~n22759 & n22761;
  assign n22763 = pi630 & n22762;
  assign n22764 = ~n22758 & ~n22763;
  assign n22765 = ~n63616 & n22764;
  assign n22766 = pi787 & ~n22765;
  assign n22767 = ~pi626 & ~n63614;
  assign n22768 = pi626 & ~n22697;
  assign n22769 = n8301 & ~n22768;
  assign n22770 = ~n22767 & n22769;
  assign n22771 = n8525 & n22752;
  assign n22772 = pi626 & ~n63614;
  assign n22773 = ~pi626 & ~n22697;
  assign n22774 = n8300 & ~n22773;
  assign n22775 = ~n22772 & n22774;
  assign n22776 = ~n22771 & ~n22775;
  assign n22777 = ~n22770 & ~n22771;
  assign n22778 = ~n22775 & n22777;
  assign n22779 = ~n22770 & n22776;
  assign n22780 = pi788 & ~n63617;
  assign n22781 = n13460 & n22717;
  assign n22782 = n11303 & n22751;
  assign n22783 = pi648 & ~n22782;
  assign n22784 = ~n22781 & n22783;
  assign n22785 = n13462 & n22717;
  assign n22786 = n11304 & n22751;
  assign n22787 = ~pi648 & ~n22786;
  assign n22788 = ~n22785 & n22787;
  assign n22789 = pi789 & ~n22788;
  assign n22790 = ~n22784 & n22789;
  assign n22791 = ~n7187 & ~n22740;
  assign n22792 = pi625 & n22791;
  assign n22793 = n22699 & ~n22791;
  assign n22794 = ~n22792 & ~n22793;
  assign n22795 = n22745 & ~n22794;
  assign n22796 = ~pi608 & ~n22744;
  assign n22797 = ~n22795 & n22796;
  assign n22798 = pi1153 & n22699;
  assign n22799 = ~n22792 & n22798;
  assign n22800 = pi608 & ~n22746;
  assign n22801 = ~n22799 & n22800;
  assign n22802 = ~n22797 & ~n22801;
  assign n22803 = pi778 & ~n22802;
  assign n22804 = ~pi778 & ~n22793;
  assign n22805 = ~n22803 & ~n22804;
  assign n22806 = ~pi609 & ~n22805;
  assign n22807 = pi609 & ~n22749;
  assign n22808 = ~pi1155 & ~n22807;
  assign n22809 = ~n22806 & n22808;
  assign n22810 = ~pi660 & ~n22704;
  assign n22811 = ~n22809 & n22810;
  assign n22812 = pi609 & ~n22805;
  assign n22813 = ~pi609 & ~n22749;
  assign n22814 = pi1155 & ~n22813;
  assign n22815 = ~n22812 & n22814;
  assign n22816 = pi660 & ~n22706;
  assign n22817 = ~n22815 & n22816;
  assign n22818 = ~n22811 & ~n22817;
  assign n22819 = pi785 & ~n22818;
  assign n22820 = ~pi785 & ~n22805;
  assign n22821 = ~n22819 & ~n22820;
  assign n22822 = pi618 & ~n22821;
  assign n22823 = ~pi618 & n22750;
  assign n22824 = pi1154 & ~n22823;
  assign n22825 = ~n22822 & n22824;
  assign n22826 = pi627 & ~n22714;
  assign n22827 = ~n22825 & n22826;
  assign n22828 = ~pi618 & ~n22821;
  assign n22829 = pi618 & n22750;
  assign n22830 = ~pi1154 & ~n22829;
  assign n22831 = ~n22828 & n22830;
  assign n22832 = ~pi627 & ~n22712;
  assign n22833 = ~n22831 & n22832;
  assign n22834 = pi781 & ~n22833;
  assign n22835 = ~n22827 & n22834;
  assign n22836 = ~pi781 & n22821;
  assign n22837 = ~n11434 & ~n22836;
  assign n22838 = ~n22835 & n22837;
  assign n22839 = ~n22790 & ~n22838;
  assign n22840 = ~n22827 & ~n22833;
  assign n22841 = pi781 & ~n22840;
  assign n22842 = ~pi781 & ~n22821;
  assign n22843 = ~n22841 & ~n22842;
  assign n22844 = ~pi619 & ~n22843;
  assign n22845 = pi619 & n22751;
  assign n22846 = ~pi1159 & ~n22845;
  assign n22847 = ~n22844 & n22846;
  assign n22848 = ~pi648 & ~n22720;
  assign n22849 = ~n22847 & n22848;
  assign n22850 = pi619 & ~n22843;
  assign n22851 = ~pi619 & n22751;
  assign n22852 = pi1159 & ~n22851;
  assign n22853 = ~n22850 & n22852;
  assign n22854 = pi648 & ~n22722;
  assign n22855 = ~n22853 & n22854;
  assign n22856 = pi789 & ~n22855;
  assign n22857 = pi789 & ~n22849;
  assign n22858 = ~n22855 & n22857;
  assign n22859 = ~n22849 & n22856;
  assign n22860 = ~pi789 & n22843;
  assign n22861 = n62894 & ~n22860;
  assign n22862 = ~n63618 & n22861;
  assign n22863 = n62894 & ~n22839;
  assign n22864 = ~n22780 & ~n63619;
  assign n22865 = ~n63030 & ~n22864;
  assign n22866 = n8498 & n63615;
  assign n22867 = n8615 & n22753;
  assign n22868 = pi629 & ~n22867;
  assign n22869 = ~n22866 & n22868;
  assign n22870 = n8499 & n63615;
  assign n22871 = n8606 & n22753;
  assign n22872 = ~pi629 & ~n22871;
  assign n22873 = ~n22870 & n22872;
  assign n22874 = pi792 & ~n22873;
  assign n22875 = pi792 & ~n22869;
  assign n22876 = ~n22873 & n22875;
  assign n22877 = ~n22870 & ~n22871;
  assign n22878 = ~pi629 & ~n22877;
  assign n22879 = ~n22866 & ~n22867;
  assign n22880 = pi629 & ~n22879;
  assign n22881 = ~n22878 & ~n22880;
  assign n22882 = pi792 & ~n22881;
  assign n22883 = ~n22869 & n22874;
  assign n22884 = ~n8651 & ~n63620;
  assign n22885 = ~n22865 & n22884;
  assign n22886 = ~n22766 & ~n22885;
  assign n22887 = pi644 & n22886;
  assign n22888 = ~pi787 & ~n22754;
  assign n22889 = pi1157 & ~n22757;
  assign n22890 = ~n22762 & ~n22889;
  assign n22891 = pi787 & ~n22890;
  assign n22892 = ~n22888 & ~n22891;
  assign n22893 = ~pi644 & n22892;
  assign n22894 = pi715 & ~n22893;
  assign n22895 = ~n22887 & n22894;
  assign n22896 = ~n8685 & n22697;
  assign n22897 = ~n8376 & n22733;
  assign n22898 = ~n8376 & ~n22736;
  assign n22899 = n8376 & n22697;
  assign n22900 = ~n22898 & ~n22899;
  assign n22901 = ~n22896 & ~n22897;
  assign n22902 = pi644 & ~n63621;
  assign n22903 = ~pi644 & n22697;
  assign n22904 = ~pi715 & ~n22903;
  assign n22905 = ~n22902 & n22904;
  assign n22906 = pi1160 & ~n22905;
  assign n22907 = ~n22895 & n22906;
  assign n22908 = ~pi644 & n22886;
  assign n22909 = pi644 & n22892;
  assign n22910 = ~pi715 & ~n22909;
  assign n22911 = ~n22908 & n22910;
  assign n22912 = ~pi644 & ~n63621;
  assign n22913 = pi644 & n22697;
  assign n22914 = pi715 & ~n22913;
  assign n22915 = ~n22912 & n22914;
  assign n22916 = ~pi1160 & ~n22915;
  assign n22917 = ~n22911 & n22916;
  assign n22918 = ~n22907 & ~n22917;
  assign n22919 = pi790 & ~n22918;
  assign n22920 = ~pi790 & n22886;
  assign n22921 = pi832 & ~n22920;
  assign n22922 = ~n22919 & n22921;
  assign n22923 = ~pi190 & ~n8098;
  assign n22924 = ~n11558 & n22923;
  assign n22925 = pi190 & ~n62765;
  assign n22926 = ~pi763 & n7143;
  assign n22927 = pi190 & n7349;
  assign n22928 = ~n22926 & ~n22927;
  assign n22929 = pi39 & ~n22928;
  assign n22930 = ~pi190 & pi763;
  assign n22931 = n62802 & n22930;
  assign n22932 = ~pi763 & n6946;
  assign n22933 = pi763 & ~n7293;
  assign n22934 = pi190 & ~n22933;
  assign n22935 = ~n22932 & ~n22934;
  assign n22936 = ~n22931 & n22935;
  assign n22937 = ~n22929 & n22936;
  assign n22938 = ~pi38 & ~n22937;
  assign n22939 = pi763 & n7359;
  assign n22940 = ~pi190 & ~n7357;
  assign n22941 = pi38 & ~n22940;
  assign n22942 = ~n22939 & n22941;
  assign n22943 = ~n22938 & ~n22942;
  assign n22944 = n62765 & ~n22943;
  assign n22945 = ~n22925 & ~n22944;
  assign n22946 = ~n8135 & ~n22945;
  assign n22947 = n8135 & ~n22923;
  assign n22948 = ~n22946 & ~n22947;
  assign n22949 = ~pi785 & ~n22948;
  assign n22950 = ~n8136 & ~n22923;
  assign n22951 = pi609 & n22946;
  assign n22952 = ~n22950 & ~n22951;
  assign n22953 = pi1155 & ~n22952;
  assign n22954 = ~n8148 & ~n22923;
  assign n22955 = ~pi609 & n22946;
  assign n22956 = ~n22954 & ~n22955;
  assign n22957 = ~pi1155 & ~n22956;
  assign n22958 = ~n22953 & ~n22957;
  assign n22959 = pi785 & ~n22958;
  assign n22960 = ~n22949 & ~n22959;
  assign n22961 = ~pi781 & ~n22960;
  assign n22962 = pi618 & n22960;
  assign n22963 = ~pi618 & n22923;
  assign n22964 = pi1154 & ~n22963;
  assign n22965 = ~n22962 & n22964;
  assign n22966 = ~pi618 & n22960;
  assign n22967 = pi618 & n22923;
  assign n22968 = ~pi1154 & ~n22967;
  assign n22969 = ~n22966 & n22968;
  assign n22970 = ~n22965 & ~n22969;
  assign n22971 = pi781 & ~n22970;
  assign n22972 = ~n22961 & ~n22971;
  assign n22973 = ~pi619 & ~n22972;
  assign n22974 = pi619 & ~n22923;
  assign n22975 = ~pi1159 & ~n22974;
  assign n22976 = ~n22973 & n22975;
  assign n22977 = pi619 & ~n22972;
  assign n22978 = ~pi619 & ~n22923;
  assign n22979 = pi1159 & ~n22978;
  assign n22980 = ~n22977 & n22979;
  assign n22981 = pi619 & n22972;
  assign n22982 = ~pi619 & n22923;
  assign n22983 = pi1159 & ~n22982;
  assign n22984 = ~n22981 & n22983;
  assign n22985 = ~pi619 & n22972;
  assign n22986 = pi619 & n22923;
  assign n22987 = ~pi1159 & ~n22986;
  assign n22988 = ~n22985 & n22987;
  assign n22989 = ~n22984 & ~n22988;
  assign n22990 = ~n22976 & ~n22980;
  assign n22991 = pi789 & n63622;
  assign n22992 = ~pi789 & n22972;
  assign n22993 = ~pi789 & ~n22972;
  assign n22994 = pi789 & ~n63622;
  assign n22995 = ~n22993 & ~n22994;
  assign n22996 = ~n22991 & ~n22992;
  assign n22997 = ~n8595 & n63623;
  assign n22998 = n8685 & n22997;
  assign n22999 = n8376 & ~n22923;
  assign n23000 = n8595 & n22923;
  assign n23001 = ~n22997 & ~n23000;
  assign n23002 = ~n8334 & ~n23001;
  assign n23003 = n8334 & n22923;
  assign n23004 = ~n23002 & ~n23003;
  assign n23005 = ~n8376 & n23004;
  assign n23006 = ~n22999 & ~n23005;
  assign n23007 = ~n8376 & ~n23004;
  assign n23008 = n8376 & n22923;
  assign n23009 = ~n23007 & ~n23008;
  assign n23010 = ~n22924 & ~n22998;
  assign n23011 = pi644 & n63624;
  assign n23012 = ~pi644 & n22923;
  assign n23013 = ~pi715 & ~n23012;
  assign n23014 = ~n23011 & n23013;
  assign n23015 = n10298 & ~n22923;
  assign n23016 = n8257 & ~n22923;
  assign n23017 = ~pi190 & n8009;
  assign n23018 = pi190 & n62874;
  assign n23019 = ~pi38 & ~n23018;
  assign n23020 = ~n23017 & n23019;
  assign n23021 = n8085 & ~n22940;
  assign n23022 = pi699 & ~n23021;
  assign n23023 = ~n23020 & n23022;
  assign n23024 = ~pi190 & ~pi699;
  assign n23025 = ~n8091 & n23024;
  assign n23026 = n62765 & ~n23025;
  assign n23027 = ~n23023 & n23026;
  assign n23028 = ~n22925 & ~n23027;
  assign n23029 = ~pi778 & ~n23028;
  assign n23030 = pi625 & n23028;
  assign n23031 = ~pi625 & n22923;
  assign n23032 = pi1153 & ~n23031;
  assign n23033 = ~n23030 & n23032;
  assign n23034 = ~pi625 & n23028;
  assign n23035 = pi625 & n22923;
  assign n23036 = ~pi1153 & ~n23035;
  assign n23037 = ~n23034 & n23036;
  assign n23038 = ~n23033 & ~n23037;
  assign n23039 = pi778 & ~n23038;
  assign n23040 = ~n23029 & ~n23039;
  assign n23041 = ~n62880 & ~n23040;
  assign n23042 = n62880 & ~n22923;
  assign n23043 = ~n62880 & n23040;
  assign n23044 = n62880 & n22923;
  assign n23045 = ~n23043 & ~n23044;
  assign n23046 = ~n23041 & ~n23042;
  assign n23047 = ~n62882 & ~n63625;
  assign n23048 = n62882 & n22923;
  assign n23049 = n62882 & ~n22923;
  assign n23050 = ~n62882 & n63625;
  assign n23051 = ~n23049 & ~n23050;
  assign n23052 = ~n23047 & ~n23048;
  assign n23053 = ~n8257 & ~n63626;
  assign n23054 = ~n8257 & n63626;
  assign n23055 = n8257 & n22923;
  assign n23056 = ~n23054 & ~n23055;
  assign n23057 = ~n23016 & ~n23053;
  assign n23058 = ~n8303 & ~n63627;
  assign n23059 = n8303 & n22923;
  assign n23060 = ~n23058 & ~n23059;
  assign n23061 = ~n62892 & ~n23060;
  assign n23062 = n62892 & n22923;
  assign n23063 = n62892 & ~n22923;
  assign n23064 = ~n62892 & n23060;
  assign n23065 = ~n23063 & ~n23064;
  assign n23066 = ~pi628 & ~n23060;
  assign n23067 = pi628 & n22923;
  assign n23068 = ~n23066 & ~n23067;
  assign n23069 = ~pi1156 & ~n23068;
  assign n23070 = pi628 & ~n23060;
  assign n23071 = ~pi628 & n22923;
  assign n23072 = ~n23070 & ~n23071;
  assign n23073 = pi1156 & ~n23072;
  assign n23074 = ~n23069 & ~n23073;
  assign n23075 = pi792 & ~n23074;
  assign n23076 = ~pi792 & ~n23060;
  assign n23077 = ~n23075 & ~n23076;
  assign n23078 = ~n23061 & ~n23062;
  assign n23079 = ~n10298 & ~n63628;
  assign n23080 = ~n10298 & n63628;
  assign n23081 = n10298 & n22923;
  assign n23082 = ~n23080 & ~n23081;
  assign n23083 = ~pi647 & n63628;
  assign n23084 = pi647 & n22923;
  assign n23085 = ~n23083 & ~n23084;
  assign n23086 = ~pi1157 & ~n23085;
  assign n23087 = pi647 & n63628;
  assign n23088 = ~pi647 & n22923;
  assign n23089 = ~n23087 & ~n23088;
  assign n23090 = pi1157 & ~n23089;
  assign n23091 = ~n23086 & ~n23090;
  assign n23092 = pi787 & ~n23091;
  assign n23093 = ~pi787 & n63628;
  assign n23094 = ~n23092 & ~n23093;
  assign n23095 = ~n23015 & ~n23079;
  assign n23096 = ~pi644 & ~n63629;
  assign n23097 = pi715 & ~n23096;
  assign n23098 = pi1160 & ~n23097;
  assign n23099 = pi1160 & ~n23014;
  assign n23100 = ~n23097 & n23099;
  assign n23101 = ~n23014 & n23098;
  assign n23102 = pi644 & ~n63629;
  assign n23103 = ~pi715 & ~n23102;
  assign n23104 = ~pi644 & n63624;
  assign n23105 = pi644 & n22923;
  assign n23106 = pi715 & ~n23105;
  assign n23107 = ~n23104 & n23106;
  assign n23108 = ~pi1160 & ~n23107;
  assign n23109 = ~n23103 & n23108;
  assign n23110 = ~n63630 & ~n23109;
  assign n23111 = pi790 & ~n23110;
  assign n23112 = ~n63052 & n23001;
  assign n23113 = n8332 & ~n23067;
  assign n23114 = n8332 & n23068;
  assign n23115 = ~n23066 & n23113;
  assign n23116 = n8331 & ~n23071;
  assign n23117 = n8331 & n23072;
  assign n23118 = ~n23070 & n23116;
  assign n23119 = ~n63631 & ~n63632;
  assign n23120 = ~n23112 & n23119;
  assign n23121 = pi792 & ~n23120;
  assign n23122 = ~pi699 & n22943;
  assign n23123 = ~pi190 & ~n62821;
  assign n23124 = pi190 & n7632;
  assign n23125 = ~pi763 & ~n23124;
  assign n23126 = ~n23123 & n23125;
  assign n23127 = pi190 & n7709;
  assign n23128 = ~pi190 & n62851;
  assign n23129 = pi763 & ~n23128;
  assign n23130 = ~n23127 & n23129;
  assign n23131 = pi39 & ~n23130;
  assign n23132 = ~n23126 & n23131;
  assign n23133 = ~pi190 & n7832;
  assign n23134 = pi190 & n7855;
  assign n23135 = ~pi763 & ~n23134;
  assign n23136 = ~pi763 & ~n23133;
  assign n23137 = ~n23134 & n23136;
  assign n23138 = ~n23133 & n23135;
  assign n23139 = ~pi190 & ~n7861;
  assign n23140 = pi190 & ~n7868;
  assign n23141 = pi763 & ~n23140;
  assign n23142 = ~n23139 & n23141;
  assign n23143 = ~pi39 & ~n23142;
  assign n23144 = ~n63633 & n23143;
  assign n23145 = ~pi38 & ~n23144;
  assign n23146 = ~pi190 & n8759;
  assign n23147 = pi190 & n8763;
  assign n23148 = ~pi763 & ~n23147;
  assign n23149 = ~n23146 & n23148;
  assign n23150 = pi190 & n8775;
  assign n23151 = ~pi190 & ~n8779;
  assign n23152 = pi763 & ~n23151;
  assign n23153 = ~n23150 & n23152;
  assign n23154 = ~n23149 & ~n23153;
  assign n23155 = ~pi38 & ~n23154;
  assign n23156 = ~n23132 & n23145;
  assign n23157 = ~pi763 & n13901;
  assign n23158 = ~n7744 & ~n23157;
  assign n23159 = ~pi39 & ~n23158;
  assign n23160 = ~pi190 & ~n23159;
  assign n23161 = ~n7565 & ~n22698;
  assign n23162 = pi190 & ~n23161;
  assign n23163 = n7356 & n23162;
  assign n23164 = pi38 & ~n23163;
  assign n23165 = ~n23160 & n23164;
  assign n23166 = pi699 & ~n23165;
  assign n23167 = ~n63634 & n23166;
  assign n23168 = n62765 & ~n23167;
  assign n23169 = n62765 & ~n23122;
  assign n23170 = ~n23167 & n23169;
  assign n23171 = ~n23122 & n23168;
  assign n23172 = ~n22925 & ~n63635;
  assign n23173 = ~pi625 & n23172;
  assign n23174 = pi625 & n22945;
  assign n23175 = ~pi1153 & ~n23174;
  assign n23176 = ~n23173 & n23175;
  assign n23177 = ~pi608 & ~n23033;
  assign n23178 = ~n23176 & n23177;
  assign n23179 = pi625 & n23172;
  assign n23180 = ~pi625 & n22945;
  assign n23181 = pi1153 & ~n23180;
  assign n23182 = ~n23179 & n23181;
  assign n23183 = pi608 & ~n23037;
  assign n23184 = ~n23182 & n23183;
  assign n23185 = ~n23178 & ~n23184;
  assign n23186 = pi778 & ~n23185;
  assign n23187 = ~pi778 & n23172;
  assign n23188 = ~n23186 & ~n23187;
  assign n23189 = ~pi609 & ~n23188;
  assign n23190 = pi609 & n23040;
  assign n23191 = ~pi1155 & ~n23190;
  assign n23192 = ~n23189 & n23191;
  assign n23193 = ~pi660 & ~n22953;
  assign n23194 = ~n23192 & n23193;
  assign n23195 = pi609 & ~n23188;
  assign n23196 = ~pi609 & n23040;
  assign n23197 = pi1155 & ~n23196;
  assign n23198 = ~n23195 & n23197;
  assign n23199 = pi660 & ~n22957;
  assign n23200 = ~n23198 & n23199;
  assign n23201 = ~n23194 & ~n23200;
  assign n23202 = pi785 & ~n23201;
  assign n23203 = ~pi785 & ~n23188;
  assign n23204 = ~n23202 & ~n23203;
  assign n23205 = ~pi781 & n23204;
  assign n23206 = ~pi618 & ~n23204;
  assign n23207 = pi618 & ~n63625;
  assign n23208 = ~pi1154 & ~n23207;
  assign n23209 = ~n23206 & n23208;
  assign n23210 = ~pi627 & ~n22965;
  assign n23211 = ~n23209 & n23210;
  assign n23212 = pi618 & ~n23204;
  assign n23213 = ~pi618 & ~n63625;
  assign n23214 = pi1154 & ~n23213;
  assign n23215 = ~n23212 & n23214;
  assign n23216 = pi627 & ~n22969;
  assign n23217 = ~n23215 & n23216;
  assign n23218 = pi781 & ~n23217;
  assign n23219 = ~n23211 & n23218;
  assign n23220 = ~n23211 & ~n23217;
  assign n23221 = pi781 & ~n23220;
  assign n23222 = ~pi781 & ~n23204;
  assign n23223 = ~n23221 & ~n23222;
  assign n23224 = ~n23205 & ~n23219;
  assign n23225 = ~n11434 & n63636;
  assign n23226 = ~n11431 & ~n63626;
  assign n23227 = ~n62884 & ~n63622;
  assign n23228 = ~n23226 & ~n23227;
  assign n23229 = pi789 & ~n23228;
  assign n23230 = n62894 & ~n23229;
  assign n23231 = ~pi619 & ~n63636;
  assign n23232 = pi619 & n63626;
  assign n23233 = ~pi1159 & ~n23232;
  assign n23234 = ~n23231 & n23233;
  assign n23235 = ~pi648 & ~n22984;
  assign n23236 = ~n23234 & n23235;
  assign n23237 = pi619 & ~n63636;
  assign n23238 = ~pi619 & n63626;
  assign n23239 = pi1159 & ~n23238;
  assign n23240 = ~n23237 & n23239;
  assign n23241 = pi648 & ~n22988;
  assign n23242 = ~n23240 & n23241;
  assign n23243 = pi789 & ~n23242;
  assign n23244 = pi789 & ~n23236;
  assign n23245 = ~n23242 & n23244;
  assign n23246 = ~n23236 & n23243;
  assign n23247 = ~pi789 & n63636;
  assign n23248 = n62894 & ~n23247;
  assign n23249 = ~n63637 & n23248;
  assign n23250 = ~n23225 & n23230;
  assign n23251 = ~pi626 & ~n63623;
  assign n23252 = pi626 & ~n22923;
  assign n23253 = n8301 & ~n23252;
  assign n23254 = ~n23251 & n23253;
  assign n23255 = n8525 & ~n63627;
  assign n23256 = pi626 & ~n63623;
  assign n23257 = ~pi626 & ~n22923;
  assign n23258 = n8300 & ~n23257;
  assign n23259 = ~n23256 & n23258;
  assign n23260 = ~n23255 & ~n23259;
  assign n23261 = ~n23254 & ~n23255;
  assign n23262 = ~n23259 & n23261;
  assign n23263 = ~n23254 & n23260;
  assign n23264 = pi788 & ~n63639;
  assign n23265 = ~n63030 & ~n23264;
  assign n23266 = ~n63638 & n23265;
  assign n23267 = ~n23121 & ~n23266;
  assign n23268 = ~n8651 & ~n23267;
  assign n23269 = ~n8413 & ~n23003;
  assign n23270 = ~n8413 & n23004;
  assign n23271 = ~n23002 & n23269;
  assign n23272 = n8374 & ~n23084;
  assign n23273 = n8374 & n23085;
  assign n23274 = ~n23083 & n23272;
  assign n23275 = n8373 & ~n23088;
  assign n23276 = n8373 & n23089;
  assign n23277 = ~n23087 & n23275;
  assign n23278 = ~n63641 & ~n63642;
  assign n23279 = ~n63640 & ~n63641;
  assign n23280 = ~n63642 & n23279;
  assign n23281 = ~n63640 & n23278;
  assign n23282 = pi787 & ~n63643;
  assign n23283 = ~pi644 & n23108;
  assign n23284 = pi644 & n23099;
  assign n23285 = n14029 & ~n23014;
  assign n23286 = pi790 & ~n63644;
  assign n23287 = pi790 & ~n23283;
  assign n23288 = ~n63644 & n23287;
  assign n23289 = ~n23283 & n23286;
  assign n23290 = ~n23282 & ~n63645;
  assign n23291 = ~n23268 & ~n23282;
  assign n23292 = ~n63645 & n23291;
  assign n23293 = ~n23268 & n23290;
  assign n23294 = ~n23111 & ~n63646;
  assign n23295 = n62455 & ~n23294;
  assign n23296 = ~pi190 & ~n62455;
  assign n23297 = ~pi832 & ~n23296;
  assign n23298 = ~n23295 & n23297;
  assign po347 = ~n22922 & ~n23298;
  assign n23300 = ~pi191 & ~n2923;
  assign n23301 = pi746 & n7316;
  assign n23302 = ~n23300 & ~n23301;
  assign n23303 = ~n8420 & ~n23302;
  assign n23304 = ~pi785 & ~n23303;
  assign n23305 = n8148 & n23301;
  assign n23306 = n23303 & ~n23305;
  assign n23307 = pi1155 & ~n23306;
  assign n23308 = ~pi1155 & ~n23300;
  assign n23309 = ~n23305 & n23308;
  assign n23310 = ~n23307 & ~n23309;
  assign n23311 = pi785 & ~n23310;
  assign n23312 = ~n23304 & ~n23311;
  assign n23313 = ~pi781 & ~n23312;
  assign n23314 = ~n8435 & n23312;
  assign n23315 = pi1154 & ~n23314;
  assign n23316 = ~n8438 & n23312;
  assign n23317 = ~pi1154 & ~n23316;
  assign n23318 = ~n23315 & ~n23317;
  assign n23319 = pi781 & ~n23318;
  assign n23320 = ~n23313 & ~n23319;
  assign n23321 = ~pi789 & ~n23320;
  assign n23322 = ~n12612 & n23320;
  assign n23323 = pi1159 & ~n23322;
  assign n23324 = ~n12615 & n23320;
  assign n23325 = ~pi1159 & ~n23324;
  assign n23326 = ~n23323 & ~n23325;
  assign n23327 = pi789 & ~n23326;
  assign n23328 = ~n23321 & ~n23327;
  assign n23329 = ~n15298 & n23320;
  assign n23330 = ~n8595 & n63647;
  assign n23331 = n8595 & n23300;
  assign n23332 = ~n8595 & ~n63647;
  assign n23333 = n8595 & ~n23300;
  assign n23334 = ~n23332 & ~n23333;
  assign n23335 = ~n23330 & ~n23331;
  assign n23336 = ~n8334 & n63648;
  assign n23337 = n8334 & n23300;
  assign n23338 = ~n8413 & ~n23337;
  assign n23339 = ~n23336 & ~n23337;
  assign n23340 = ~n8413 & n23339;
  assign n23341 = ~n23336 & n23338;
  assign n23342 = pi729 & n7564;
  assign n23343 = ~n23300 & ~n23342;
  assign n23344 = ~pi778 & ~n23343;
  assign n23345 = ~pi625 & n23342;
  assign n23346 = ~n23343 & ~n23345;
  assign n23347 = pi1153 & ~n23346;
  assign n23348 = ~pi1153 & ~n23300;
  assign n23349 = ~n23345 & n23348;
  assign n23350 = pi778 & ~n23349;
  assign n23351 = ~n23347 & n23350;
  assign n23352 = ~n23344 & ~n23351;
  assign n23353 = ~n8490 & ~n23352;
  assign n23354 = ~n8492 & n23353;
  assign n23355 = ~n8494 & n23354;
  assign n23356 = ~n8496 & n23355;
  assign n23357 = ~n8508 & n23356;
  assign n23358 = pi647 & ~n23357;
  assign n23359 = ~pi647 & ~n23300;
  assign n23360 = ~n23358 & ~n23359;
  assign n23361 = n8373 & ~n23360;
  assign n23362 = ~pi647 & n23357;
  assign n23363 = pi647 & n23300;
  assign n23364 = ~pi1157 & ~n23363;
  assign n23365 = ~n23362 & n23364;
  assign n23366 = pi630 & n23365;
  assign n23367 = ~n23361 & ~n23366;
  assign n23368 = ~n63649 & n23367;
  assign n23369 = pi787 & ~n23368;
  assign n23370 = ~pi626 & ~n63647;
  assign n23371 = pi626 & ~n23300;
  assign n23372 = n8301 & ~n23371;
  assign n23373 = ~n23370 & n23372;
  assign n23374 = n8525 & n23355;
  assign n23375 = pi626 & ~n63647;
  assign n23376 = ~pi626 & ~n23300;
  assign n23377 = n8300 & ~n23376;
  assign n23378 = ~n23375 & n23377;
  assign n23379 = ~n23374 & ~n23378;
  assign n23380 = ~n23373 & ~n23374;
  assign n23381 = ~n23378 & n23380;
  assign n23382 = ~n23373 & n23379;
  assign n23383 = pi788 & ~n63650;
  assign n23384 = n13460 & n23320;
  assign n23385 = n11303 & n23354;
  assign n23386 = pi648 & ~n23385;
  assign n23387 = ~n23384 & n23386;
  assign n23388 = n13462 & n23320;
  assign n23389 = n11304 & n23354;
  assign n23390 = ~pi648 & ~n23389;
  assign n23391 = ~n23388 & n23390;
  assign n23392 = pi789 & ~n23391;
  assign n23393 = ~n23387 & n23392;
  assign n23394 = ~n7187 & ~n23343;
  assign n23395 = pi625 & n23394;
  assign n23396 = n23302 & ~n23394;
  assign n23397 = ~n23395 & ~n23396;
  assign n23398 = n23348 & ~n23397;
  assign n23399 = ~pi608 & ~n23347;
  assign n23400 = ~n23398 & n23399;
  assign n23401 = pi1153 & n23302;
  assign n23402 = ~n23395 & n23401;
  assign n23403 = pi608 & ~n23349;
  assign n23404 = ~n23402 & n23403;
  assign n23405 = ~n23400 & ~n23404;
  assign n23406 = pi778 & ~n23405;
  assign n23407 = ~pi778 & ~n23396;
  assign n23408 = ~n23406 & ~n23407;
  assign n23409 = ~pi609 & ~n23408;
  assign n23410 = pi609 & ~n23352;
  assign n23411 = ~pi1155 & ~n23410;
  assign n23412 = ~n23409 & n23411;
  assign n23413 = ~pi660 & ~n23307;
  assign n23414 = ~n23412 & n23413;
  assign n23415 = pi609 & ~n23408;
  assign n23416 = ~pi609 & ~n23352;
  assign n23417 = pi1155 & ~n23416;
  assign n23418 = ~n23415 & n23417;
  assign n23419 = pi660 & ~n23309;
  assign n23420 = ~n23418 & n23419;
  assign n23421 = ~n23414 & ~n23420;
  assign n23422 = pi785 & ~n23421;
  assign n23423 = ~pi785 & ~n23408;
  assign n23424 = ~n23422 & ~n23423;
  assign n23425 = pi618 & ~n23424;
  assign n23426 = ~pi618 & n23353;
  assign n23427 = pi1154 & ~n23426;
  assign n23428 = ~n23425 & n23427;
  assign n23429 = pi627 & ~n23317;
  assign n23430 = ~n23428 & n23429;
  assign n23431 = ~pi618 & ~n23424;
  assign n23432 = pi618 & n23353;
  assign n23433 = ~pi1154 & ~n23432;
  assign n23434 = ~n23431 & n23433;
  assign n23435 = ~pi627 & ~n23315;
  assign n23436 = ~n23434 & n23435;
  assign n23437 = pi781 & ~n23436;
  assign n23438 = ~n23430 & n23437;
  assign n23439 = ~pi781 & n23424;
  assign n23440 = ~n11434 & ~n23439;
  assign n23441 = ~n23438 & n23440;
  assign n23442 = ~n23393 & ~n23441;
  assign n23443 = ~n23430 & ~n23436;
  assign n23444 = pi781 & ~n23443;
  assign n23445 = ~pi781 & ~n23424;
  assign n23446 = ~n23444 & ~n23445;
  assign n23447 = ~pi619 & ~n23446;
  assign n23448 = pi619 & n23354;
  assign n23449 = ~pi1159 & ~n23448;
  assign n23450 = ~n23447 & n23449;
  assign n23451 = ~pi648 & ~n23323;
  assign n23452 = ~n23450 & n23451;
  assign n23453 = pi619 & ~n23446;
  assign n23454 = ~pi619 & n23354;
  assign n23455 = pi1159 & ~n23454;
  assign n23456 = ~n23453 & n23455;
  assign n23457 = pi648 & ~n23325;
  assign n23458 = ~n23456 & n23457;
  assign n23459 = pi789 & ~n23458;
  assign n23460 = pi789 & ~n23452;
  assign n23461 = ~n23458 & n23460;
  assign n23462 = ~n23452 & n23459;
  assign n23463 = ~pi789 & n23446;
  assign n23464 = n62894 & ~n23463;
  assign n23465 = ~n63651 & n23464;
  assign n23466 = n62894 & ~n23442;
  assign n23467 = ~n23383 & ~n63652;
  assign n23468 = ~n63030 & ~n23467;
  assign n23469 = n8498 & n63648;
  assign n23470 = n8615 & n23356;
  assign n23471 = pi629 & ~n23470;
  assign n23472 = ~n23469 & n23471;
  assign n23473 = n8499 & n63648;
  assign n23474 = n8606 & n23356;
  assign n23475 = ~pi629 & ~n23474;
  assign n23476 = ~n23473 & n23475;
  assign n23477 = pi792 & ~n23476;
  assign n23478 = pi792 & ~n23472;
  assign n23479 = ~n23476 & n23478;
  assign n23480 = ~n23473 & ~n23474;
  assign n23481 = ~pi629 & ~n23480;
  assign n23482 = ~n23469 & ~n23470;
  assign n23483 = pi629 & ~n23482;
  assign n23484 = ~n23481 & ~n23483;
  assign n23485 = pi792 & ~n23484;
  assign n23486 = ~n23472 & n23477;
  assign n23487 = ~n8651 & ~n63653;
  assign n23488 = ~n23468 & n23487;
  assign n23489 = ~n23369 & ~n23488;
  assign n23490 = pi644 & n23489;
  assign n23491 = ~pi787 & ~n23357;
  assign n23492 = pi1157 & ~n23360;
  assign n23493 = ~n23365 & ~n23492;
  assign n23494 = pi787 & ~n23493;
  assign n23495 = ~n23491 & ~n23494;
  assign n23496 = ~pi644 & n23495;
  assign n23497 = pi715 & ~n23496;
  assign n23498 = ~n23490 & n23497;
  assign n23499 = ~n8685 & n23300;
  assign n23500 = ~n8376 & n23336;
  assign n23501 = ~n8376 & ~n23339;
  assign n23502 = n8376 & n23300;
  assign n23503 = ~n23501 & ~n23502;
  assign n23504 = ~n23499 & ~n23500;
  assign n23505 = pi644 & ~n63654;
  assign n23506 = ~pi644 & n23300;
  assign n23507 = ~pi715 & ~n23506;
  assign n23508 = ~n23505 & n23507;
  assign n23509 = pi1160 & ~n23508;
  assign n23510 = ~n23498 & n23509;
  assign n23511 = ~pi644 & n23489;
  assign n23512 = pi644 & n23495;
  assign n23513 = ~pi715 & ~n23512;
  assign n23514 = ~n23511 & n23513;
  assign n23515 = ~pi644 & ~n63654;
  assign n23516 = pi644 & n23300;
  assign n23517 = pi715 & ~n23516;
  assign n23518 = ~n23515 & n23517;
  assign n23519 = ~pi1160 & ~n23518;
  assign n23520 = ~n23514 & n23519;
  assign n23521 = ~n23510 & ~n23520;
  assign n23522 = pi790 & ~n23521;
  assign n23523 = ~pi790 & n23489;
  assign n23524 = pi832 & ~n23523;
  assign n23525 = ~n23522 & n23524;
  assign n23526 = ~pi191 & ~n8098;
  assign n23527 = ~n11558 & n23526;
  assign n23528 = pi191 & ~n62765;
  assign n23529 = ~pi746 & n7143;
  assign n23530 = pi191 & n7349;
  assign n23531 = ~n23529 & ~n23530;
  assign n23532 = pi39 & ~n23531;
  assign n23533 = ~pi191 & pi746;
  assign n23534 = n62802 & n23533;
  assign n23535 = ~pi746 & n6946;
  assign n23536 = pi746 & ~n7293;
  assign n23537 = pi191 & ~n23536;
  assign n23538 = ~n23535 & ~n23537;
  assign n23539 = ~n23534 & n23538;
  assign n23540 = ~n23532 & n23539;
  assign n23541 = ~pi38 & ~n23540;
  assign n23542 = pi746 & n7359;
  assign n23543 = ~pi191 & ~n7357;
  assign n23544 = pi38 & ~n23543;
  assign n23545 = ~n23542 & n23544;
  assign n23546 = ~n23541 & ~n23545;
  assign n23547 = n62765 & ~n23546;
  assign n23548 = ~n23528 & ~n23547;
  assign n23549 = ~n8135 & ~n23548;
  assign n23550 = n8135 & ~n23526;
  assign n23551 = ~n23549 & ~n23550;
  assign n23552 = ~pi785 & ~n23551;
  assign n23553 = ~n8136 & ~n23526;
  assign n23554 = pi609 & n23549;
  assign n23555 = ~n23553 & ~n23554;
  assign n23556 = pi1155 & ~n23555;
  assign n23557 = ~n8148 & ~n23526;
  assign n23558 = ~pi609 & n23549;
  assign n23559 = ~n23557 & ~n23558;
  assign n23560 = ~pi1155 & ~n23559;
  assign n23561 = ~n23556 & ~n23560;
  assign n23562 = pi785 & ~n23561;
  assign n23563 = ~n23552 & ~n23562;
  assign n23564 = ~pi781 & ~n23563;
  assign n23565 = pi618 & n23563;
  assign n23566 = ~pi618 & n23526;
  assign n23567 = pi1154 & ~n23566;
  assign n23568 = ~n23565 & n23567;
  assign n23569 = ~pi618 & n23563;
  assign n23570 = pi618 & n23526;
  assign n23571 = ~pi1154 & ~n23570;
  assign n23572 = ~n23569 & n23571;
  assign n23573 = ~n23568 & ~n23572;
  assign n23574 = pi781 & ~n23573;
  assign n23575 = ~n23564 & ~n23574;
  assign n23576 = ~pi619 & ~n23575;
  assign n23577 = pi619 & ~n23526;
  assign n23578 = ~pi1159 & ~n23577;
  assign n23579 = ~n23576 & n23578;
  assign n23580 = pi619 & ~n23575;
  assign n23581 = ~pi619 & ~n23526;
  assign n23582 = pi1159 & ~n23581;
  assign n23583 = ~n23580 & n23582;
  assign n23584 = pi619 & n23575;
  assign n23585 = ~pi619 & n23526;
  assign n23586 = pi1159 & ~n23585;
  assign n23587 = ~n23584 & n23586;
  assign n23588 = ~pi619 & n23575;
  assign n23589 = pi619 & n23526;
  assign n23590 = ~pi1159 & ~n23589;
  assign n23591 = ~n23588 & n23590;
  assign n23592 = ~n23587 & ~n23591;
  assign n23593 = ~n23579 & ~n23583;
  assign n23594 = pi789 & n63655;
  assign n23595 = ~pi789 & n23575;
  assign n23596 = ~pi789 & ~n23575;
  assign n23597 = pi789 & ~n63655;
  assign n23598 = ~n23596 & ~n23597;
  assign n23599 = ~n23594 & ~n23595;
  assign n23600 = ~n8595 & n63656;
  assign n23601 = n8685 & n23600;
  assign n23602 = n8376 & ~n23526;
  assign n23603 = n8595 & n23526;
  assign n23604 = ~n23600 & ~n23603;
  assign n23605 = ~n8334 & ~n23604;
  assign n23606 = n8334 & n23526;
  assign n23607 = ~n23605 & ~n23606;
  assign n23608 = ~n8376 & n23607;
  assign n23609 = ~n23602 & ~n23608;
  assign n23610 = ~n8376 & ~n23607;
  assign n23611 = n8376 & n23526;
  assign n23612 = ~n23610 & ~n23611;
  assign n23613 = ~n23527 & ~n23601;
  assign n23614 = pi644 & n63657;
  assign n23615 = ~pi644 & n23526;
  assign n23616 = ~pi715 & ~n23615;
  assign n23617 = ~n23614 & n23616;
  assign n23618 = n10298 & ~n23526;
  assign n23619 = n8257 & ~n23526;
  assign n23620 = ~pi191 & n8009;
  assign n23621 = pi191 & n62874;
  assign n23622 = ~pi38 & ~n23621;
  assign n23623 = ~n23620 & n23622;
  assign n23624 = n8085 & ~n23543;
  assign n23625 = pi729 & ~n23624;
  assign n23626 = ~n23623 & n23625;
  assign n23627 = ~pi191 & ~pi729;
  assign n23628 = ~n8091 & n23627;
  assign n23629 = n62765 & ~n23628;
  assign n23630 = ~n23626 & n23629;
  assign n23631 = ~n23528 & ~n23630;
  assign n23632 = ~pi778 & ~n23631;
  assign n23633 = pi625 & n23631;
  assign n23634 = ~pi625 & n23526;
  assign n23635 = pi1153 & ~n23634;
  assign n23636 = ~n23633 & n23635;
  assign n23637 = ~pi625 & n23631;
  assign n23638 = pi625 & n23526;
  assign n23639 = ~pi1153 & ~n23638;
  assign n23640 = ~n23637 & n23639;
  assign n23641 = ~n23636 & ~n23640;
  assign n23642 = pi778 & ~n23641;
  assign n23643 = ~n23632 & ~n23642;
  assign n23644 = ~n62880 & ~n23643;
  assign n23645 = n62880 & ~n23526;
  assign n23646 = ~n62880 & n23643;
  assign n23647 = n62880 & n23526;
  assign n23648 = ~n23646 & ~n23647;
  assign n23649 = ~n23644 & ~n23645;
  assign n23650 = ~n62882 & ~n63658;
  assign n23651 = n62882 & n23526;
  assign n23652 = n62882 & ~n23526;
  assign n23653 = ~n62882 & n63658;
  assign n23654 = ~n23652 & ~n23653;
  assign n23655 = ~n23650 & ~n23651;
  assign n23656 = ~n8257 & ~n63659;
  assign n23657 = ~n8257 & n63659;
  assign n23658 = n8257 & n23526;
  assign n23659 = ~n23657 & ~n23658;
  assign n23660 = ~n23619 & ~n23656;
  assign n23661 = ~n8303 & ~n63660;
  assign n23662 = n8303 & n23526;
  assign n23663 = ~n23661 & ~n23662;
  assign n23664 = ~n62892 & ~n23663;
  assign n23665 = n62892 & n23526;
  assign n23666 = n62892 & ~n23526;
  assign n23667 = ~n62892 & n23663;
  assign n23668 = ~n23666 & ~n23667;
  assign n23669 = ~pi628 & ~n23663;
  assign n23670 = pi628 & n23526;
  assign n23671 = ~n23669 & ~n23670;
  assign n23672 = ~pi1156 & ~n23671;
  assign n23673 = pi628 & ~n23663;
  assign n23674 = ~pi628 & n23526;
  assign n23675 = ~n23673 & ~n23674;
  assign n23676 = pi1156 & ~n23675;
  assign n23677 = ~n23672 & ~n23676;
  assign n23678 = pi792 & ~n23677;
  assign n23679 = ~pi792 & ~n23663;
  assign n23680 = ~n23678 & ~n23679;
  assign n23681 = ~n23664 & ~n23665;
  assign n23682 = ~n10298 & ~n63661;
  assign n23683 = ~n10298 & n63661;
  assign n23684 = n10298 & n23526;
  assign n23685 = ~n23683 & ~n23684;
  assign n23686 = ~pi647 & n63661;
  assign n23687 = pi647 & n23526;
  assign n23688 = ~n23686 & ~n23687;
  assign n23689 = ~pi1157 & ~n23688;
  assign n23690 = pi647 & n63661;
  assign n23691 = ~pi647 & n23526;
  assign n23692 = ~n23690 & ~n23691;
  assign n23693 = pi1157 & ~n23692;
  assign n23694 = ~n23689 & ~n23693;
  assign n23695 = pi787 & ~n23694;
  assign n23696 = ~pi787 & n63661;
  assign n23697 = ~n23695 & ~n23696;
  assign n23698 = ~n23618 & ~n23682;
  assign n23699 = ~pi644 & ~n63662;
  assign n23700 = pi715 & ~n23699;
  assign n23701 = pi1160 & ~n23700;
  assign n23702 = pi1160 & ~n23617;
  assign n23703 = ~n23700 & n23702;
  assign n23704 = ~n23617 & n23701;
  assign n23705 = pi644 & ~n63662;
  assign n23706 = ~pi715 & ~n23705;
  assign n23707 = ~pi644 & n63657;
  assign n23708 = pi644 & n23526;
  assign n23709 = pi715 & ~n23708;
  assign n23710 = ~n23707 & n23709;
  assign n23711 = ~pi1160 & ~n23710;
  assign n23712 = ~n23706 & n23711;
  assign n23713 = ~n63663 & ~n23712;
  assign n23714 = pi790 & ~n23713;
  assign n23715 = ~n63052 & n23604;
  assign n23716 = n8332 & ~n23670;
  assign n23717 = n8332 & n23671;
  assign n23718 = ~n23669 & n23716;
  assign n23719 = n8331 & ~n23674;
  assign n23720 = n8331 & n23675;
  assign n23721 = ~n23673 & n23719;
  assign n23722 = ~n63664 & ~n63665;
  assign n23723 = ~n23715 & n23722;
  assign n23724 = pi792 & ~n23723;
  assign n23725 = ~pi729 & n23546;
  assign n23726 = ~pi191 & ~n62821;
  assign n23727 = pi191 & n7632;
  assign n23728 = ~pi746 & ~n23727;
  assign n23729 = ~n23726 & n23728;
  assign n23730 = pi191 & n7709;
  assign n23731 = ~pi191 & n62851;
  assign n23732 = pi746 & ~n23731;
  assign n23733 = ~n23730 & n23732;
  assign n23734 = pi39 & ~n23733;
  assign n23735 = ~n23729 & n23734;
  assign n23736 = ~pi191 & n7832;
  assign n23737 = pi191 & n7855;
  assign n23738 = ~pi746 & ~n23737;
  assign n23739 = ~pi746 & ~n23736;
  assign n23740 = ~n23737 & n23739;
  assign n23741 = ~n23736 & n23738;
  assign n23742 = ~pi191 & ~n7861;
  assign n23743 = pi191 & ~n7868;
  assign n23744 = pi746 & ~n23743;
  assign n23745 = ~n23742 & n23744;
  assign n23746 = ~pi39 & ~n23745;
  assign n23747 = ~n63666 & n23746;
  assign n23748 = ~pi38 & ~n23747;
  assign n23749 = ~pi191 & n8759;
  assign n23750 = pi191 & n8763;
  assign n23751 = ~pi746 & ~n23750;
  assign n23752 = ~n23749 & n23751;
  assign n23753 = pi191 & n8775;
  assign n23754 = ~pi191 & ~n8779;
  assign n23755 = pi746 & ~n23754;
  assign n23756 = ~n23753 & n23755;
  assign n23757 = ~n23752 & ~n23756;
  assign n23758 = ~pi38 & ~n23757;
  assign n23759 = ~n23735 & n23748;
  assign n23760 = ~pi746 & n13901;
  assign n23761 = ~n7744 & ~n23760;
  assign n23762 = ~pi39 & ~n23761;
  assign n23763 = ~pi191 & ~n23762;
  assign n23764 = ~n7565 & ~n23301;
  assign n23765 = pi191 & ~n23764;
  assign n23766 = n7356 & n23765;
  assign n23767 = pi38 & ~n23766;
  assign n23768 = ~n23763 & n23767;
  assign n23769 = pi729 & ~n23768;
  assign n23770 = ~n63667 & n23769;
  assign n23771 = n62765 & ~n23770;
  assign n23772 = n62765 & ~n23725;
  assign n23773 = ~n23770 & n23772;
  assign n23774 = ~n23725 & n23771;
  assign n23775 = ~n23528 & ~n63668;
  assign n23776 = ~pi625 & n23775;
  assign n23777 = pi625 & n23548;
  assign n23778 = ~pi1153 & ~n23777;
  assign n23779 = ~n23776 & n23778;
  assign n23780 = ~pi608 & ~n23636;
  assign n23781 = ~n23779 & n23780;
  assign n23782 = pi625 & n23775;
  assign n23783 = ~pi625 & n23548;
  assign n23784 = pi1153 & ~n23783;
  assign n23785 = ~n23782 & n23784;
  assign n23786 = pi608 & ~n23640;
  assign n23787 = ~n23785 & n23786;
  assign n23788 = ~n23781 & ~n23787;
  assign n23789 = pi778 & ~n23788;
  assign n23790 = ~pi778 & n23775;
  assign n23791 = ~n23789 & ~n23790;
  assign n23792 = ~pi609 & ~n23791;
  assign n23793 = pi609 & n23643;
  assign n23794 = ~pi1155 & ~n23793;
  assign n23795 = ~n23792 & n23794;
  assign n23796 = ~pi660 & ~n23556;
  assign n23797 = ~n23795 & n23796;
  assign n23798 = pi609 & ~n23791;
  assign n23799 = ~pi609 & n23643;
  assign n23800 = pi1155 & ~n23799;
  assign n23801 = ~n23798 & n23800;
  assign n23802 = pi660 & ~n23560;
  assign n23803 = ~n23801 & n23802;
  assign n23804 = ~n23797 & ~n23803;
  assign n23805 = pi785 & ~n23804;
  assign n23806 = ~pi785 & ~n23791;
  assign n23807 = ~n23805 & ~n23806;
  assign n23808 = ~pi781 & n23807;
  assign n23809 = ~pi618 & ~n23807;
  assign n23810 = pi618 & ~n63658;
  assign n23811 = ~pi1154 & ~n23810;
  assign n23812 = ~n23809 & n23811;
  assign n23813 = ~pi627 & ~n23568;
  assign n23814 = ~n23812 & n23813;
  assign n23815 = pi618 & ~n23807;
  assign n23816 = ~pi618 & ~n63658;
  assign n23817 = pi1154 & ~n23816;
  assign n23818 = ~n23815 & n23817;
  assign n23819 = pi627 & ~n23572;
  assign n23820 = ~n23818 & n23819;
  assign n23821 = pi781 & ~n23820;
  assign n23822 = ~n23814 & n23821;
  assign n23823 = ~n23814 & ~n23820;
  assign n23824 = pi781 & ~n23823;
  assign n23825 = ~pi781 & ~n23807;
  assign n23826 = ~n23824 & ~n23825;
  assign n23827 = ~n23808 & ~n23822;
  assign n23828 = ~n11434 & n63669;
  assign n23829 = ~n11431 & ~n63659;
  assign n23830 = ~n62884 & ~n63655;
  assign n23831 = ~n23829 & ~n23830;
  assign n23832 = pi789 & ~n23831;
  assign n23833 = n62894 & ~n23832;
  assign n23834 = ~pi619 & ~n63669;
  assign n23835 = pi619 & n63659;
  assign n23836 = ~pi1159 & ~n23835;
  assign n23837 = ~n23834 & n23836;
  assign n23838 = ~pi648 & ~n23587;
  assign n23839 = ~n23837 & n23838;
  assign n23840 = pi619 & ~n63669;
  assign n23841 = ~pi619 & n63659;
  assign n23842 = pi1159 & ~n23841;
  assign n23843 = ~n23840 & n23842;
  assign n23844 = pi648 & ~n23591;
  assign n23845 = ~n23843 & n23844;
  assign n23846 = pi789 & ~n23845;
  assign n23847 = pi789 & ~n23839;
  assign n23848 = ~n23845 & n23847;
  assign n23849 = ~n23839 & n23846;
  assign n23850 = ~pi789 & n63669;
  assign n23851 = n62894 & ~n23850;
  assign n23852 = ~n63670 & n23851;
  assign n23853 = ~n23828 & n23833;
  assign n23854 = ~pi626 & ~n63656;
  assign n23855 = pi626 & ~n23526;
  assign n23856 = n8301 & ~n23855;
  assign n23857 = ~n23854 & n23856;
  assign n23858 = n8525 & ~n63660;
  assign n23859 = pi626 & ~n63656;
  assign n23860 = ~pi626 & ~n23526;
  assign n23861 = n8300 & ~n23860;
  assign n23862 = ~n23859 & n23861;
  assign n23863 = ~n23858 & ~n23862;
  assign n23864 = ~n23857 & ~n23858;
  assign n23865 = ~n23862 & n23864;
  assign n23866 = ~n23857 & n23863;
  assign n23867 = pi788 & ~n63672;
  assign n23868 = ~n63030 & ~n23867;
  assign n23869 = ~n63671 & n23868;
  assign n23870 = ~n23724 & ~n23869;
  assign n23871 = ~n8651 & ~n23870;
  assign n23872 = ~n8413 & ~n23606;
  assign n23873 = ~n8413 & n23607;
  assign n23874 = ~n23605 & n23872;
  assign n23875 = n8374 & ~n23687;
  assign n23876 = n8374 & n23688;
  assign n23877 = ~n23686 & n23875;
  assign n23878 = n8373 & ~n23691;
  assign n23879 = n8373 & n23692;
  assign n23880 = ~n23690 & n23878;
  assign n23881 = ~n63674 & ~n63675;
  assign n23882 = ~n63673 & ~n63674;
  assign n23883 = ~n63675 & n23882;
  assign n23884 = ~n63673 & n23881;
  assign n23885 = pi787 & ~n63676;
  assign n23886 = ~pi644 & n23711;
  assign n23887 = pi644 & n23702;
  assign n23888 = n14029 & ~n23617;
  assign n23889 = pi790 & ~n63677;
  assign n23890 = pi790 & ~n23886;
  assign n23891 = ~n63677 & n23890;
  assign n23892 = ~n23886 & n23889;
  assign n23893 = ~n23885 & ~n63678;
  assign n23894 = ~n23871 & ~n23885;
  assign n23895 = ~n63678 & n23894;
  assign n23896 = ~n23871 & n23893;
  assign n23897 = ~n23714 & ~n63679;
  assign n23898 = n62455 & ~n23897;
  assign n23899 = ~pi191 & ~n62455;
  assign n23900 = ~pi832 & ~n23899;
  assign n23901 = ~n23898 & n23900;
  assign po348 = ~n23525 & ~n23901;
  assign n23903 = ~pi192 & ~n2923;
  assign n23904 = pi764 & n7316;
  assign n23905 = ~n23903 & ~n23904;
  assign n23906 = ~n8420 & ~n23905;
  assign n23907 = ~pi785 & ~n23906;
  assign n23908 = n8148 & n23904;
  assign n23909 = n23906 & ~n23908;
  assign n23910 = pi1155 & ~n23909;
  assign n23911 = ~pi1155 & ~n23903;
  assign n23912 = ~n23908 & n23911;
  assign n23913 = ~n23910 & ~n23912;
  assign n23914 = pi785 & ~n23913;
  assign n23915 = ~n23907 & ~n23914;
  assign n23916 = ~pi781 & ~n23915;
  assign n23917 = ~n8435 & n23915;
  assign n23918 = pi1154 & ~n23917;
  assign n23919 = ~n8438 & n23915;
  assign n23920 = ~pi1154 & ~n23919;
  assign n23921 = ~n23918 & ~n23920;
  assign n23922 = pi781 & ~n23921;
  assign n23923 = ~n23916 & ~n23922;
  assign n23924 = ~pi789 & ~n23923;
  assign n23925 = ~n12612 & n23923;
  assign n23926 = pi1159 & ~n23925;
  assign n23927 = ~n12615 & n23923;
  assign n23928 = ~pi1159 & ~n23927;
  assign n23929 = ~n23926 & ~n23928;
  assign n23930 = pi789 & ~n23929;
  assign n23931 = ~n23924 & ~n23930;
  assign n23932 = ~n15298 & n23923;
  assign n23933 = ~n8595 & n63680;
  assign n23934 = n8595 & n23903;
  assign n23935 = ~n8595 & ~n63680;
  assign n23936 = n8595 & ~n23903;
  assign n23937 = ~n23935 & ~n23936;
  assign n23938 = ~n23933 & ~n23934;
  assign n23939 = ~n8334 & n63681;
  assign n23940 = n8334 & n23903;
  assign n23941 = ~n8413 & ~n23940;
  assign n23942 = ~n23939 & ~n23940;
  assign n23943 = ~n8413 & n23942;
  assign n23944 = ~n23939 & n23941;
  assign n23945 = pi691 & n7564;
  assign n23946 = ~n23903 & ~n23945;
  assign n23947 = ~pi778 & ~n23946;
  assign n23948 = ~pi625 & n23945;
  assign n23949 = ~n23946 & ~n23948;
  assign n23950 = pi1153 & ~n23949;
  assign n23951 = ~pi1153 & ~n23903;
  assign n23952 = ~n23948 & n23951;
  assign n23953 = pi778 & ~n23952;
  assign n23954 = ~n23950 & n23953;
  assign n23955 = ~n23947 & ~n23954;
  assign n23956 = ~n8490 & ~n23955;
  assign n23957 = ~n8492 & n23956;
  assign n23958 = ~n8494 & n23957;
  assign n23959 = ~n8496 & n23958;
  assign n23960 = ~n8508 & n23959;
  assign n23961 = pi647 & ~n23960;
  assign n23962 = ~pi647 & ~n23903;
  assign n23963 = ~n23961 & ~n23962;
  assign n23964 = n8373 & ~n23963;
  assign n23965 = ~pi647 & n23960;
  assign n23966 = pi647 & n23903;
  assign n23967 = ~pi1157 & ~n23966;
  assign n23968 = ~n23965 & n23967;
  assign n23969 = pi630 & n23968;
  assign n23970 = ~n23964 & ~n23969;
  assign n23971 = ~n63682 & n23970;
  assign n23972 = pi787 & ~n23971;
  assign n23973 = ~pi626 & ~n63680;
  assign n23974 = pi626 & ~n23903;
  assign n23975 = n8301 & ~n23974;
  assign n23976 = ~n23973 & n23975;
  assign n23977 = n8525 & n23958;
  assign n23978 = pi626 & ~n63680;
  assign n23979 = ~pi626 & ~n23903;
  assign n23980 = n8300 & ~n23979;
  assign n23981 = ~n23978 & n23980;
  assign n23982 = ~n23977 & ~n23981;
  assign n23983 = ~n23976 & ~n23977;
  assign n23984 = ~n23981 & n23983;
  assign n23985 = ~n23976 & n23982;
  assign n23986 = pi788 & ~n63683;
  assign n23987 = n13460 & n23923;
  assign n23988 = n11303 & n23957;
  assign n23989 = pi648 & ~n23988;
  assign n23990 = ~n23987 & n23989;
  assign n23991 = n13462 & n23923;
  assign n23992 = n11304 & n23957;
  assign n23993 = ~pi648 & ~n23992;
  assign n23994 = ~n23991 & n23993;
  assign n23995 = pi789 & ~n23994;
  assign n23996 = ~n23990 & n23995;
  assign n23997 = ~n7187 & ~n23946;
  assign n23998 = pi625 & n23997;
  assign n23999 = n23905 & ~n23997;
  assign n24000 = ~n23998 & ~n23999;
  assign n24001 = n23951 & ~n24000;
  assign n24002 = ~pi608 & ~n23950;
  assign n24003 = ~n24001 & n24002;
  assign n24004 = pi1153 & n23905;
  assign n24005 = ~n23998 & n24004;
  assign n24006 = pi608 & ~n23952;
  assign n24007 = ~n24005 & n24006;
  assign n24008 = ~n24003 & ~n24007;
  assign n24009 = pi778 & ~n24008;
  assign n24010 = ~pi778 & ~n23999;
  assign n24011 = ~n24009 & ~n24010;
  assign n24012 = ~pi609 & ~n24011;
  assign n24013 = pi609 & ~n23955;
  assign n24014 = ~pi1155 & ~n24013;
  assign n24015 = ~n24012 & n24014;
  assign n24016 = ~pi660 & ~n23910;
  assign n24017 = ~n24015 & n24016;
  assign n24018 = pi609 & ~n24011;
  assign n24019 = ~pi609 & ~n23955;
  assign n24020 = pi1155 & ~n24019;
  assign n24021 = ~n24018 & n24020;
  assign n24022 = pi660 & ~n23912;
  assign n24023 = ~n24021 & n24022;
  assign n24024 = ~n24017 & ~n24023;
  assign n24025 = pi785 & ~n24024;
  assign n24026 = ~pi785 & ~n24011;
  assign n24027 = ~n24025 & ~n24026;
  assign n24028 = pi618 & ~n24027;
  assign n24029 = ~pi618 & n23956;
  assign n24030 = pi1154 & ~n24029;
  assign n24031 = ~n24028 & n24030;
  assign n24032 = pi627 & ~n23920;
  assign n24033 = ~n24031 & n24032;
  assign n24034 = ~pi618 & ~n24027;
  assign n24035 = pi618 & n23956;
  assign n24036 = ~pi1154 & ~n24035;
  assign n24037 = ~n24034 & n24036;
  assign n24038 = ~pi627 & ~n23918;
  assign n24039 = ~n24037 & n24038;
  assign n24040 = pi781 & ~n24039;
  assign n24041 = ~n24033 & n24040;
  assign n24042 = ~pi781 & n24027;
  assign n24043 = ~n11434 & ~n24042;
  assign n24044 = ~n24041 & n24043;
  assign n24045 = ~n23996 & ~n24044;
  assign n24046 = ~n24033 & ~n24039;
  assign n24047 = pi781 & ~n24046;
  assign n24048 = ~pi781 & ~n24027;
  assign n24049 = ~n24047 & ~n24048;
  assign n24050 = ~pi619 & ~n24049;
  assign n24051 = pi619 & n23957;
  assign n24052 = ~pi1159 & ~n24051;
  assign n24053 = ~n24050 & n24052;
  assign n24054 = ~pi648 & ~n23926;
  assign n24055 = ~n24053 & n24054;
  assign n24056 = pi619 & ~n24049;
  assign n24057 = ~pi619 & n23957;
  assign n24058 = pi1159 & ~n24057;
  assign n24059 = ~n24056 & n24058;
  assign n24060 = pi648 & ~n23928;
  assign n24061 = ~n24059 & n24060;
  assign n24062 = pi789 & ~n24061;
  assign n24063 = pi789 & ~n24055;
  assign n24064 = ~n24061 & n24063;
  assign n24065 = ~n24055 & n24062;
  assign n24066 = ~pi789 & n24049;
  assign n24067 = n62894 & ~n24066;
  assign n24068 = ~n63684 & n24067;
  assign n24069 = n62894 & ~n24045;
  assign n24070 = ~n23986 & ~n63685;
  assign n24071 = ~n63030 & ~n24070;
  assign n24072 = n8498 & n63681;
  assign n24073 = n8615 & n23959;
  assign n24074 = pi629 & ~n24073;
  assign n24075 = ~n24072 & n24074;
  assign n24076 = n8499 & n63681;
  assign n24077 = n8606 & n23959;
  assign n24078 = ~pi629 & ~n24077;
  assign n24079 = ~n24076 & n24078;
  assign n24080 = pi792 & ~n24079;
  assign n24081 = pi792 & ~n24075;
  assign n24082 = ~n24079 & n24081;
  assign n24083 = ~n24076 & ~n24077;
  assign n24084 = ~pi629 & ~n24083;
  assign n24085 = ~n24072 & ~n24073;
  assign n24086 = pi629 & ~n24085;
  assign n24087 = ~n24084 & ~n24086;
  assign n24088 = pi792 & ~n24087;
  assign n24089 = ~n24075 & n24080;
  assign n24090 = ~n8651 & ~n63686;
  assign n24091 = ~n24071 & n24090;
  assign n24092 = ~n23972 & ~n24091;
  assign n24093 = pi644 & n24092;
  assign n24094 = ~pi787 & ~n23960;
  assign n24095 = pi1157 & ~n23963;
  assign n24096 = ~n23968 & ~n24095;
  assign n24097 = pi787 & ~n24096;
  assign n24098 = ~n24094 & ~n24097;
  assign n24099 = ~pi644 & n24098;
  assign n24100 = pi715 & ~n24099;
  assign n24101 = ~n24093 & n24100;
  assign n24102 = ~n8685 & n23903;
  assign n24103 = ~n8376 & n23939;
  assign n24104 = ~n8376 & ~n23942;
  assign n24105 = n8376 & n23903;
  assign n24106 = ~n24104 & ~n24105;
  assign n24107 = ~n24102 & ~n24103;
  assign n24108 = pi644 & ~n63687;
  assign n24109 = ~pi644 & n23903;
  assign n24110 = ~pi715 & ~n24109;
  assign n24111 = ~n24108 & n24110;
  assign n24112 = pi1160 & ~n24111;
  assign n24113 = ~n24101 & n24112;
  assign n24114 = ~pi644 & n24092;
  assign n24115 = pi644 & n24098;
  assign n24116 = ~pi715 & ~n24115;
  assign n24117 = ~n24114 & n24116;
  assign n24118 = ~pi644 & ~n63687;
  assign n24119 = pi644 & n23903;
  assign n24120 = pi715 & ~n24119;
  assign n24121 = ~n24118 & n24120;
  assign n24122 = ~pi1160 & ~n24121;
  assign n24123 = ~n24117 & n24122;
  assign n24124 = ~n24113 & ~n24123;
  assign n24125 = pi790 & ~n24124;
  assign n24126 = ~pi790 & n24092;
  assign n24127 = pi832 & ~n24126;
  assign n24128 = ~n24125 & n24127;
  assign n24129 = ~pi192 & ~n8098;
  assign n24130 = ~n11558 & n24129;
  assign n24131 = pi192 & ~n62765;
  assign n24132 = ~pi764 & n7143;
  assign n24133 = pi192 & n7349;
  assign n24134 = ~n24132 & ~n24133;
  assign n24135 = pi39 & ~n24134;
  assign n24136 = ~pi192 & pi764;
  assign n24137 = n62802 & n24136;
  assign n24138 = ~pi764 & n6946;
  assign n24139 = pi764 & ~n7293;
  assign n24140 = pi192 & ~n24139;
  assign n24141 = ~n24138 & ~n24140;
  assign n24142 = ~n24137 & n24141;
  assign n24143 = ~n24135 & n24142;
  assign n24144 = ~pi38 & ~n24143;
  assign n24145 = pi764 & n7359;
  assign n24146 = ~pi192 & ~n7357;
  assign n24147 = pi38 & ~n24146;
  assign n24148 = ~n24145 & n24147;
  assign n24149 = ~n24144 & ~n24148;
  assign n24150 = n62765 & ~n24149;
  assign n24151 = ~n24131 & ~n24150;
  assign n24152 = ~n8135 & ~n24151;
  assign n24153 = n8135 & ~n24129;
  assign n24154 = ~n24152 & ~n24153;
  assign n24155 = ~pi785 & ~n24154;
  assign n24156 = ~n8136 & ~n24129;
  assign n24157 = pi609 & n24152;
  assign n24158 = ~n24156 & ~n24157;
  assign n24159 = pi1155 & ~n24158;
  assign n24160 = ~n8148 & ~n24129;
  assign n24161 = ~pi609 & n24152;
  assign n24162 = ~n24160 & ~n24161;
  assign n24163 = ~pi1155 & ~n24162;
  assign n24164 = ~n24159 & ~n24163;
  assign n24165 = pi785 & ~n24164;
  assign n24166 = ~n24155 & ~n24165;
  assign n24167 = ~pi781 & ~n24166;
  assign n24168 = pi618 & n24166;
  assign n24169 = ~pi618 & n24129;
  assign n24170 = pi1154 & ~n24169;
  assign n24171 = ~n24168 & n24170;
  assign n24172 = ~pi618 & n24166;
  assign n24173 = pi618 & n24129;
  assign n24174 = ~pi1154 & ~n24173;
  assign n24175 = ~n24172 & n24174;
  assign n24176 = ~n24171 & ~n24175;
  assign n24177 = pi781 & ~n24176;
  assign n24178 = ~n24167 & ~n24177;
  assign n24179 = ~pi619 & ~n24178;
  assign n24180 = pi619 & ~n24129;
  assign n24181 = ~pi1159 & ~n24180;
  assign n24182 = ~n24179 & n24181;
  assign n24183 = pi619 & ~n24178;
  assign n24184 = ~pi619 & ~n24129;
  assign n24185 = pi1159 & ~n24184;
  assign n24186 = ~n24183 & n24185;
  assign n24187 = pi619 & n24178;
  assign n24188 = ~pi619 & n24129;
  assign n24189 = pi1159 & ~n24188;
  assign n24190 = ~n24187 & n24189;
  assign n24191 = ~pi619 & n24178;
  assign n24192 = pi619 & n24129;
  assign n24193 = ~pi1159 & ~n24192;
  assign n24194 = ~n24191 & n24193;
  assign n24195 = ~n24190 & ~n24194;
  assign n24196 = ~n24182 & ~n24186;
  assign n24197 = pi789 & n63688;
  assign n24198 = ~pi789 & n24178;
  assign n24199 = ~pi789 & ~n24178;
  assign n24200 = pi789 & ~n63688;
  assign n24201 = ~n24199 & ~n24200;
  assign n24202 = ~n24197 & ~n24198;
  assign n24203 = ~n8595 & n63689;
  assign n24204 = n8685 & n24203;
  assign n24205 = n8376 & ~n24129;
  assign n24206 = n8595 & n24129;
  assign n24207 = ~n24203 & ~n24206;
  assign n24208 = ~n8334 & ~n24207;
  assign n24209 = n8334 & n24129;
  assign n24210 = ~n24208 & ~n24209;
  assign n24211 = ~n8376 & n24210;
  assign n24212 = ~n24205 & ~n24211;
  assign n24213 = ~n8376 & ~n24210;
  assign n24214 = n8376 & n24129;
  assign n24215 = ~n24213 & ~n24214;
  assign n24216 = ~n24130 & ~n24204;
  assign n24217 = pi644 & n63690;
  assign n24218 = ~pi644 & n24129;
  assign n24219 = ~pi715 & ~n24218;
  assign n24220 = ~n24217 & n24219;
  assign n24221 = n10298 & ~n24129;
  assign n24222 = n8257 & ~n24129;
  assign n24223 = ~pi192 & n8009;
  assign n24224 = pi192 & n62874;
  assign n24225 = ~pi38 & ~n24224;
  assign n24226 = ~n24223 & n24225;
  assign n24227 = n8085 & ~n24146;
  assign n24228 = pi691 & ~n24227;
  assign n24229 = ~n24226 & n24228;
  assign n24230 = ~pi192 & ~pi691;
  assign n24231 = ~n8091 & n24230;
  assign n24232 = n62765 & ~n24231;
  assign n24233 = ~n24229 & n24232;
  assign n24234 = ~n24131 & ~n24233;
  assign n24235 = ~pi778 & ~n24234;
  assign n24236 = pi625 & n24234;
  assign n24237 = ~pi625 & n24129;
  assign n24238 = pi1153 & ~n24237;
  assign n24239 = ~n24236 & n24238;
  assign n24240 = ~pi625 & n24234;
  assign n24241 = pi625 & n24129;
  assign n24242 = ~pi1153 & ~n24241;
  assign n24243 = ~n24240 & n24242;
  assign n24244 = ~n24239 & ~n24243;
  assign n24245 = pi778 & ~n24244;
  assign n24246 = ~n24235 & ~n24245;
  assign n24247 = ~n62880 & ~n24246;
  assign n24248 = n62880 & ~n24129;
  assign n24249 = ~n62880 & n24246;
  assign n24250 = n62880 & n24129;
  assign n24251 = ~n24249 & ~n24250;
  assign n24252 = ~n24247 & ~n24248;
  assign n24253 = ~n62882 & ~n63691;
  assign n24254 = n62882 & n24129;
  assign n24255 = n62882 & ~n24129;
  assign n24256 = ~n62882 & n63691;
  assign n24257 = ~n24255 & ~n24256;
  assign n24258 = ~n24253 & ~n24254;
  assign n24259 = ~n8257 & ~n63692;
  assign n24260 = ~n8257 & n63692;
  assign n24261 = n8257 & n24129;
  assign n24262 = ~n24260 & ~n24261;
  assign n24263 = ~n24222 & ~n24259;
  assign n24264 = ~n8303 & ~n63693;
  assign n24265 = n8303 & n24129;
  assign n24266 = ~n24264 & ~n24265;
  assign n24267 = ~n62892 & ~n24266;
  assign n24268 = n62892 & n24129;
  assign n24269 = n62892 & ~n24129;
  assign n24270 = ~n62892 & n24266;
  assign n24271 = ~n24269 & ~n24270;
  assign n24272 = ~pi628 & ~n24266;
  assign n24273 = pi628 & n24129;
  assign n24274 = ~n24272 & ~n24273;
  assign n24275 = ~pi1156 & ~n24274;
  assign n24276 = pi628 & ~n24266;
  assign n24277 = ~pi628 & n24129;
  assign n24278 = ~n24276 & ~n24277;
  assign n24279 = pi1156 & ~n24278;
  assign n24280 = ~n24275 & ~n24279;
  assign n24281 = pi792 & ~n24280;
  assign n24282 = ~pi792 & ~n24266;
  assign n24283 = ~n24281 & ~n24282;
  assign n24284 = ~n24267 & ~n24268;
  assign n24285 = ~n10298 & ~n63694;
  assign n24286 = ~n10298 & n63694;
  assign n24287 = n10298 & n24129;
  assign n24288 = ~n24286 & ~n24287;
  assign n24289 = ~pi647 & n63694;
  assign n24290 = pi647 & n24129;
  assign n24291 = ~n24289 & ~n24290;
  assign n24292 = ~pi1157 & ~n24291;
  assign n24293 = pi647 & n63694;
  assign n24294 = ~pi647 & n24129;
  assign n24295 = ~n24293 & ~n24294;
  assign n24296 = pi1157 & ~n24295;
  assign n24297 = ~n24292 & ~n24296;
  assign n24298 = pi787 & ~n24297;
  assign n24299 = ~pi787 & n63694;
  assign n24300 = ~n24298 & ~n24299;
  assign n24301 = ~n24221 & ~n24285;
  assign n24302 = ~pi644 & ~n63695;
  assign n24303 = pi715 & ~n24302;
  assign n24304 = pi1160 & ~n24303;
  assign n24305 = pi1160 & ~n24220;
  assign n24306 = ~n24303 & n24305;
  assign n24307 = ~n24220 & n24304;
  assign n24308 = pi644 & ~n63695;
  assign n24309 = ~pi715 & ~n24308;
  assign n24310 = ~pi644 & n63690;
  assign n24311 = pi644 & n24129;
  assign n24312 = pi715 & ~n24311;
  assign n24313 = ~n24310 & n24312;
  assign n24314 = ~pi1160 & ~n24313;
  assign n24315 = ~n24309 & n24314;
  assign n24316 = ~n63696 & ~n24315;
  assign n24317 = pi790 & ~n24316;
  assign n24318 = ~n63052 & n24207;
  assign n24319 = n8332 & ~n24273;
  assign n24320 = n8332 & n24274;
  assign n24321 = ~n24272 & n24319;
  assign n24322 = n8331 & ~n24277;
  assign n24323 = n8331 & n24278;
  assign n24324 = ~n24276 & n24322;
  assign n24325 = ~n63697 & ~n63698;
  assign n24326 = ~n24318 & n24325;
  assign n24327 = pi792 & ~n24326;
  assign n24328 = ~pi691 & n24149;
  assign n24329 = ~pi192 & ~n62821;
  assign n24330 = pi192 & n7632;
  assign n24331 = ~pi764 & ~n24330;
  assign n24332 = ~n24329 & n24331;
  assign n24333 = pi192 & n7709;
  assign n24334 = ~pi192 & n62851;
  assign n24335 = pi764 & ~n24334;
  assign n24336 = ~n24333 & n24335;
  assign n24337 = pi39 & ~n24336;
  assign n24338 = ~n24332 & n24337;
  assign n24339 = ~pi192 & n7832;
  assign n24340 = pi192 & n7855;
  assign n24341 = ~pi764 & ~n24340;
  assign n24342 = ~pi764 & ~n24339;
  assign n24343 = ~n24340 & n24342;
  assign n24344 = ~n24339 & n24341;
  assign n24345 = ~pi192 & ~n7861;
  assign n24346 = pi192 & ~n7868;
  assign n24347 = pi764 & ~n24346;
  assign n24348 = ~n24345 & n24347;
  assign n24349 = ~pi39 & ~n24348;
  assign n24350 = ~n63699 & n24349;
  assign n24351 = ~pi38 & ~n24350;
  assign n24352 = ~pi192 & n8759;
  assign n24353 = pi192 & n8763;
  assign n24354 = ~pi764 & ~n24353;
  assign n24355 = ~n24352 & n24354;
  assign n24356 = pi192 & n8775;
  assign n24357 = ~pi192 & ~n8779;
  assign n24358 = pi764 & ~n24357;
  assign n24359 = ~n24356 & n24358;
  assign n24360 = ~n24355 & ~n24359;
  assign n24361 = ~pi38 & ~n24360;
  assign n24362 = ~n24338 & n24351;
  assign n24363 = ~pi764 & n13901;
  assign n24364 = ~n7744 & ~n24363;
  assign n24365 = ~pi39 & ~n24364;
  assign n24366 = ~pi192 & ~n24365;
  assign n24367 = ~n7565 & ~n23904;
  assign n24368 = pi192 & ~n24367;
  assign n24369 = n7356 & n24368;
  assign n24370 = pi38 & ~n24369;
  assign n24371 = ~n24366 & n24370;
  assign n24372 = pi691 & ~n24371;
  assign n24373 = ~n63700 & n24372;
  assign n24374 = n62765 & ~n24373;
  assign n24375 = n62765 & ~n24328;
  assign n24376 = ~n24373 & n24375;
  assign n24377 = ~n24328 & n24374;
  assign n24378 = ~n24131 & ~n63701;
  assign n24379 = ~pi625 & n24378;
  assign n24380 = pi625 & n24151;
  assign n24381 = ~pi1153 & ~n24380;
  assign n24382 = ~n24379 & n24381;
  assign n24383 = ~pi608 & ~n24239;
  assign n24384 = ~n24382 & n24383;
  assign n24385 = pi625 & n24378;
  assign n24386 = ~pi625 & n24151;
  assign n24387 = pi1153 & ~n24386;
  assign n24388 = ~n24385 & n24387;
  assign n24389 = pi608 & ~n24243;
  assign n24390 = ~n24388 & n24389;
  assign n24391 = ~n24384 & ~n24390;
  assign n24392 = pi778 & ~n24391;
  assign n24393 = ~pi778 & n24378;
  assign n24394 = ~n24392 & ~n24393;
  assign n24395 = ~pi609 & ~n24394;
  assign n24396 = pi609 & n24246;
  assign n24397 = ~pi1155 & ~n24396;
  assign n24398 = ~n24395 & n24397;
  assign n24399 = ~pi660 & ~n24159;
  assign n24400 = ~n24398 & n24399;
  assign n24401 = pi609 & ~n24394;
  assign n24402 = ~pi609 & n24246;
  assign n24403 = pi1155 & ~n24402;
  assign n24404 = ~n24401 & n24403;
  assign n24405 = pi660 & ~n24163;
  assign n24406 = ~n24404 & n24405;
  assign n24407 = ~n24400 & ~n24406;
  assign n24408 = pi785 & ~n24407;
  assign n24409 = ~pi785 & ~n24394;
  assign n24410 = ~n24408 & ~n24409;
  assign n24411 = ~pi781 & n24410;
  assign n24412 = ~pi618 & ~n24410;
  assign n24413 = pi618 & ~n63691;
  assign n24414 = ~pi1154 & ~n24413;
  assign n24415 = ~n24412 & n24414;
  assign n24416 = ~pi627 & ~n24171;
  assign n24417 = ~n24415 & n24416;
  assign n24418 = pi618 & ~n24410;
  assign n24419 = ~pi618 & ~n63691;
  assign n24420 = pi1154 & ~n24419;
  assign n24421 = ~n24418 & n24420;
  assign n24422 = pi627 & ~n24175;
  assign n24423 = ~n24421 & n24422;
  assign n24424 = pi781 & ~n24423;
  assign n24425 = ~n24417 & n24424;
  assign n24426 = ~n24417 & ~n24423;
  assign n24427 = pi781 & ~n24426;
  assign n24428 = ~pi781 & ~n24410;
  assign n24429 = ~n24427 & ~n24428;
  assign n24430 = ~n24411 & ~n24425;
  assign n24431 = ~n11434 & n63702;
  assign n24432 = ~n11431 & ~n63692;
  assign n24433 = ~n62884 & ~n63688;
  assign n24434 = ~n24432 & ~n24433;
  assign n24435 = pi789 & ~n24434;
  assign n24436 = n62894 & ~n24435;
  assign n24437 = ~pi619 & ~n63702;
  assign n24438 = pi619 & n63692;
  assign n24439 = ~pi1159 & ~n24438;
  assign n24440 = ~n24437 & n24439;
  assign n24441 = ~pi648 & ~n24190;
  assign n24442 = ~n24440 & n24441;
  assign n24443 = pi619 & ~n63702;
  assign n24444 = ~pi619 & n63692;
  assign n24445 = pi1159 & ~n24444;
  assign n24446 = ~n24443 & n24445;
  assign n24447 = pi648 & ~n24194;
  assign n24448 = ~n24446 & n24447;
  assign n24449 = pi789 & ~n24448;
  assign n24450 = pi789 & ~n24442;
  assign n24451 = ~n24448 & n24450;
  assign n24452 = ~n24442 & n24449;
  assign n24453 = ~pi789 & n63702;
  assign n24454 = n62894 & ~n24453;
  assign n24455 = ~n63703 & n24454;
  assign n24456 = ~n24431 & n24436;
  assign n24457 = ~pi626 & ~n63689;
  assign n24458 = pi626 & ~n24129;
  assign n24459 = n8301 & ~n24458;
  assign n24460 = ~n24457 & n24459;
  assign n24461 = n8525 & ~n63693;
  assign n24462 = pi626 & ~n63689;
  assign n24463 = ~pi626 & ~n24129;
  assign n24464 = n8300 & ~n24463;
  assign n24465 = ~n24462 & n24464;
  assign n24466 = ~n24461 & ~n24465;
  assign n24467 = ~n24460 & ~n24461;
  assign n24468 = ~n24465 & n24467;
  assign n24469 = ~n24460 & n24466;
  assign n24470 = pi788 & ~n63705;
  assign n24471 = ~n63030 & ~n24470;
  assign n24472 = ~n63704 & n24471;
  assign n24473 = ~n24327 & ~n24472;
  assign n24474 = ~n8651 & ~n24473;
  assign n24475 = ~n8413 & ~n24209;
  assign n24476 = ~n8413 & n24210;
  assign n24477 = ~n24208 & n24475;
  assign n24478 = n8374 & ~n24290;
  assign n24479 = n8374 & n24291;
  assign n24480 = ~n24289 & n24478;
  assign n24481 = n8373 & ~n24294;
  assign n24482 = n8373 & n24295;
  assign n24483 = ~n24293 & n24481;
  assign n24484 = ~n63707 & ~n63708;
  assign n24485 = ~n63706 & ~n63707;
  assign n24486 = ~n63708 & n24485;
  assign n24487 = ~n63706 & n24484;
  assign n24488 = pi787 & ~n63709;
  assign n24489 = ~pi644 & n24314;
  assign n24490 = pi644 & n24305;
  assign n24491 = n14029 & ~n24220;
  assign n24492 = pi790 & ~n63710;
  assign n24493 = pi790 & ~n24489;
  assign n24494 = ~n63710 & n24493;
  assign n24495 = ~n24489 & n24492;
  assign n24496 = ~n24488 & ~n63711;
  assign n24497 = ~n24474 & ~n24488;
  assign n24498 = ~n63711 & n24497;
  assign n24499 = ~n24474 & n24496;
  assign n24500 = ~n24317 & ~n63712;
  assign n24501 = n62455 & ~n24500;
  assign n24502 = ~pi192 & ~n62455;
  assign n24503 = ~pi832 & ~n24502;
  assign n24504 = ~n24501 & n24503;
  assign po349 = ~n24128 & ~n24504;
  assign n24506 = ~pi193 & ~n2923;
  assign n24507 = pi739 & n7316;
  assign n24508 = ~n24506 & ~n24507;
  assign n24509 = ~n8420 & ~n24508;
  assign n24510 = ~pi785 & ~n24509;
  assign n24511 = n8148 & n24507;
  assign n24512 = n24509 & ~n24511;
  assign n24513 = pi1155 & ~n24512;
  assign n24514 = ~pi1155 & ~n24506;
  assign n24515 = ~n24511 & n24514;
  assign n24516 = ~n24513 & ~n24515;
  assign n24517 = pi785 & ~n24516;
  assign n24518 = ~n24510 & ~n24517;
  assign n24519 = ~pi781 & ~n24518;
  assign n24520 = ~n8435 & n24518;
  assign n24521 = pi1154 & ~n24520;
  assign n24522 = ~n8438 & n24518;
  assign n24523 = ~pi1154 & ~n24522;
  assign n24524 = ~n24521 & ~n24523;
  assign n24525 = pi781 & ~n24524;
  assign n24526 = ~n24519 & ~n24525;
  assign n24527 = ~pi789 & ~n24526;
  assign n24528 = ~n12612 & n24526;
  assign n24529 = pi1159 & ~n24528;
  assign n24530 = ~n12615 & n24526;
  assign n24531 = ~pi1159 & ~n24530;
  assign n24532 = ~n24529 & ~n24531;
  assign n24533 = pi789 & ~n24532;
  assign n24534 = ~n24527 & ~n24533;
  assign n24535 = ~n15298 & n24526;
  assign n24536 = ~n8595 & n63713;
  assign n24537 = n8595 & n24506;
  assign n24538 = ~n8595 & ~n63713;
  assign n24539 = n8595 & ~n24506;
  assign n24540 = ~n24538 & ~n24539;
  assign n24541 = ~n24536 & ~n24537;
  assign n24542 = ~n8334 & n63714;
  assign n24543 = n8334 & n24506;
  assign n24544 = ~n8413 & ~n24543;
  assign n24545 = ~n24542 & ~n24543;
  assign n24546 = ~n8413 & n24545;
  assign n24547 = ~n24542 & n24544;
  assign n24548 = pi690 & n7564;
  assign n24549 = ~n24506 & ~n24548;
  assign n24550 = ~pi778 & ~n24549;
  assign n24551 = ~pi625 & n24548;
  assign n24552 = ~n24549 & ~n24551;
  assign n24553 = pi1153 & ~n24552;
  assign n24554 = ~pi1153 & ~n24506;
  assign n24555 = ~n24551 & n24554;
  assign n24556 = pi778 & ~n24555;
  assign n24557 = ~n24553 & n24556;
  assign n24558 = ~n24550 & ~n24557;
  assign n24559 = ~n8490 & ~n24558;
  assign n24560 = ~n8492 & n24559;
  assign n24561 = ~n8494 & n24560;
  assign n24562 = ~n8496 & n24561;
  assign n24563 = ~n8508 & n24562;
  assign n24564 = pi647 & ~n24563;
  assign n24565 = ~pi647 & ~n24506;
  assign n24566 = ~n24564 & ~n24565;
  assign n24567 = n8373 & ~n24566;
  assign n24568 = ~pi647 & n24563;
  assign n24569 = pi647 & n24506;
  assign n24570 = ~pi1157 & ~n24569;
  assign n24571 = ~n24568 & n24570;
  assign n24572 = pi630 & n24571;
  assign n24573 = ~n24567 & ~n24572;
  assign n24574 = ~n63715 & n24573;
  assign n24575 = pi787 & ~n24574;
  assign n24576 = ~pi626 & ~n63713;
  assign n24577 = pi626 & ~n24506;
  assign n24578 = n8301 & ~n24577;
  assign n24579 = ~n24576 & n24578;
  assign n24580 = n8525 & n24561;
  assign n24581 = pi626 & ~n63713;
  assign n24582 = ~pi626 & ~n24506;
  assign n24583 = n8300 & ~n24582;
  assign n24584 = ~n24581 & n24583;
  assign n24585 = ~n24580 & ~n24584;
  assign n24586 = ~n24579 & ~n24580;
  assign n24587 = ~n24584 & n24586;
  assign n24588 = ~n24579 & n24585;
  assign n24589 = pi788 & ~n63716;
  assign n24590 = n13460 & n24526;
  assign n24591 = n11303 & n24560;
  assign n24592 = pi648 & ~n24591;
  assign n24593 = ~n24590 & n24592;
  assign n24594 = n13462 & n24526;
  assign n24595 = n11304 & n24560;
  assign n24596 = ~pi648 & ~n24595;
  assign n24597 = ~n24594 & n24596;
  assign n24598 = pi789 & ~n24597;
  assign n24599 = ~n24593 & n24598;
  assign n24600 = ~n7187 & ~n24549;
  assign n24601 = pi625 & n24600;
  assign n24602 = n24508 & ~n24600;
  assign n24603 = ~n24601 & ~n24602;
  assign n24604 = n24554 & ~n24603;
  assign n24605 = ~pi608 & ~n24553;
  assign n24606 = ~n24604 & n24605;
  assign n24607 = pi1153 & n24508;
  assign n24608 = ~n24601 & n24607;
  assign n24609 = pi608 & ~n24555;
  assign n24610 = ~n24608 & n24609;
  assign n24611 = ~n24606 & ~n24610;
  assign n24612 = pi778 & ~n24611;
  assign n24613 = ~pi778 & ~n24602;
  assign n24614 = ~n24612 & ~n24613;
  assign n24615 = ~pi609 & ~n24614;
  assign n24616 = pi609 & ~n24558;
  assign n24617 = ~pi1155 & ~n24616;
  assign n24618 = ~n24615 & n24617;
  assign n24619 = ~pi660 & ~n24513;
  assign n24620 = ~n24618 & n24619;
  assign n24621 = pi609 & ~n24614;
  assign n24622 = ~pi609 & ~n24558;
  assign n24623 = pi1155 & ~n24622;
  assign n24624 = ~n24621 & n24623;
  assign n24625 = pi660 & ~n24515;
  assign n24626 = ~n24624 & n24625;
  assign n24627 = ~n24620 & ~n24626;
  assign n24628 = pi785 & ~n24627;
  assign n24629 = ~pi785 & ~n24614;
  assign n24630 = ~n24628 & ~n24629;
  assign n24631 = pi618 & ~n24630;
  assign n24632 = ~pi618 & n24559;
  assign n24633 = pi1154 & ~n24632;
  assign n24634 = ~n24631 & n24633;
  assign n24635 = pi627 & ~n24523;
  assign n24636 = ~n24634 & n24635;
  assign n24637 = ~pi618 & ~n24630;
  assign n24638 = pi618 & n24559;
  assign n24639 = ~pi1154 & ~n24638;
  assign n24640 = ~n24637 & n24639;
  assign n24641 = ~pi627 & ~n24521;
  assign n24642 = ~n24640 & n24641;
  assign n24643 = pi781 & ~n24642;
  assign n24644 = ~n24636 & n24643;
  assign n24645 = ~pi781 & n24630;
  assign n24646 = ~n11434 & ~n24645;
  assign n24647 = ~n24644 & n24646;
  assign n24648 = ~n24599 & ~n24647;
  assign n24649 = ~n24636 & ~n24642;
  assign n24650 = pi781 & ~n24649;
  assign n24651 = ~pi781 & ~n24630;
  assign n24652 = ~n24650 & ~n24651;
  assign n24653 = ~pi619 & ~n24652;
  assign n24654 = pi619 & n24560;
  assign n24655 = ~pi1159 & ~n24654;
  assign n24656 = ~n24653 & n24655;
  assign n24657 = ~pi648 & ~n24529;
  assign n24658 = ~n24656 & n24657;
  assign n24659 = pi619 & ~n24652;
  assign n24660 = ~pi619 & n24560;
  assign n24661 = pi1159 & ~n24660;
  assign n24662 = ~n24659 & n24661;
  assign n24663 = pi648 & ~n24531;
  assign n24664 = ~n24662 & n24663;
  assign n24665 = pi789 & ~n24664;
  assign n24666 = pi789 & ~n24658;
  assign n24667 = ~n24664 & n24666;
  assign n24668 = ~n24658 & n24665;
  assign n24669 = ~pi789 & n24652;
  assign n24670 = n62894 & ~n24669;
  assign n24671 = ~n63717 & n24670;
  assign n24672 = n62894 & ~n24648;
  assign n24673 = ~n24589 & ~n63718;
  assign n24674 = ~n63030 & ~n24673;
  assign n24675 = n8498 & n63714;
  assign n24676 = n8615 & n24562;
  assign n24677 = pi629 & ~n24676;
  assign n24678 = ~n24675 & n24677;
  assign n24679 = n8499 & n63714;
  assign n24680 = n8606 & n24562;
  assign n24681 = ~pi629 & ~n24680;
  assign n24682 = ~n24679 & n24681;
  assign n24683 = pi792 & ~n24682;
  assign n24684 = pi792 & ~n24678;
  assign n24685 = ~n24682 & n24684;
  assign n24686 = ~n24679 & ~n24680;
  assign n24687 = ~pi629 & ~n24686;
  assign n24688 = ~n24675 & ~n24676;
  assign n24689 = pi629 & ~n24688;
  assign n24690 = ~n24687 & ~n24689;
  assign n24691 = pi792 & ~n24690;
  assign n24692 = ~n24678 & n24683;
  assign n24693 = ~n8651 & ~n63719;
  assign n24694 = ~n24674 & n24693;
  assign n24695 = ~n24575 & ~n24694;
  assign n24696 = pi644 & n24695;
  assign n24697 = ~pi787 & ~n24563;
  assign n24698 = pi1157 & ~n24566;
  assign n24699 = ~n24571 & ~n24698;
  assign n24700 = pi787 & ~n24699;
  assign n24701 = ~n24697 & ~n24700;
  assign n24702 = ~pi644 & n24701;
  assign n24703 = pi715 & ~n24702;
  assign n24704 = ~n24696 & n24703;
  assign n24705 = ~n8685 & n24506;
  assign n24706 = ~n8376 & n24542;
  assign n24707 = ~n8376 & ~n24545;
  assign n24708 = n8376 & n24506;
  assign n24709 = ~n24707 & ~n24708;
  assign n24710 = ~n24705 & ~n24706;
  assign n24711 = pi644 & ~n63720;
  assign n24712 = ~pi644 & n24506;
  assign n24713 = ~pi715 & ~n24712;
  assign n24714 = ~n24711 & n24713;
  assign n24715 = pi1160 & ~n24714;
  assign n24716 = ~n24704 & n24715;
  assign n24717 = ~pi644 & n24695;
  assign n24718 = pi644 & n24701;
  assign n24719 = ~pi715 & ~n24718;
  assign n24720 = ~n24717 & n24719;
  assign n24721 = ~pi644 & ~n63720;
  assign n24722 = pi644 & n24506;
  assign n24723 = pi715 & ~n24722;
  assign n24724 = ~n24721 & n24723;
  assign n24725 = ~pi1160 & ~n24724;
  assign n24726 = ~n24720 & n24725;
  assign n24727 = ~n24716 & ~n24726;
  assign n24728 = pi790 & ~n24727;
  assign n24729 = ~pi790 & n24695;
  assign n24730 = pi832 & ~n24729;
  assign n24731 = ~n24728 & n24730;
  assign n24732 = ~pi193 & ~n8098;
  assign n24733 = n8257 & ~n24732;
  assign n24734 = pi690 & n62765;
  assign n24735 = n24732 & ~n24734;
  assign n24736 = pi193 & n62874;
  assign n24737 = ~pi38 & ~n24736;
  assign n24738 = n62765 & ~n24737;
  assign n24739 = ~pi193 & n8009;
  assign n24740 = ~n24738 & ~n24739;
  assign n24741 = ~pi193 & ~n7357;
  assign n24742 = n8085 & ~n24741;
  assign n24743 = pi690 & ~n24742;
  assign n24744 = ~n24740 & n24743;
  assign n24745 = ~n24735 & ~n24744;
  assign n24746 = ~pi778 & n24745;
  assign n24747 = pi625 & ~n24745;
  assign n24748 = ~pi625 & n24732;
  assign n24749 = pi1153 & ~n24748;
  assign n24750 = ~n24747 & n24749;
  assign n24751 = ~pi625 & ~n24745;
  assign n24752 = pi625 & n24732;
  assign n24753 = ~pi1153 & ~n24752;
  assign n24754 = ~n24751 & n24753;
  assign n24755 = ~n24750 & ~n24754;
  assign n24756 = pi778 & ~n24755;
  assign n24757 = ~n24746 & ~n24756;
  assign n24758 = ~n62880 & ~n24757;
  assign n24759 = n62880 & ~n24732;
  assign n24760 = ~n62880 & n24757;
  assign n24761 = n62880 & n24732;
  assign n24762 = ~n24760 & ~n24761;
  assign n24763 = ~n24758 & ~n24759;
  assign n24764 = ~n62882 & ~n63721;
  assign n24765 = n62882 & n24732;
  assign n24766 = n62882 & ~n24732;
  assign n24767 = ~n62882 & n63721;
  assign n24768 = ~n24766 & ~n24767;
  assign n24769 = ~n24764 & ~n24765;
  assign n24770 = ~n8257 & ~n63722;
  assign n24771 = ~n8257 & n63722;
  assign n24772 = n8257 & n24732;
  assign n24773 = ~n24771 & ~n24772;
  assign n24774 = ~n24733 & ~n24770;
  assign n24775 = ~n8303 & ~n63723;
  assign n24776 = n8303 & n24732;
  assign n24777 = ~n24775 & ~n24776;
  assign n24778 = ~pi792 & n24777;
  assign n24779 = pi628 & ~n24777;
  assign n24780 = ~pi628 & n24732;
  assign n24781 = pi1156 & ~n24780;
  assign n24782 = ~n24779 & n24781;
  assign n24783 = ~pi628 & ~n24777;
  assign n24784 = pi628 & n24732;
  assign n24785 = ~pi1156 & ~n24784;
  assign n24786 = ~n24783 & n24785;
  assign n24787 = ~n24782 & ~n24786;
  assign n24788 = pi792 & ~n24787;
  assign n24789 = ~n24778 & ~n24788;
  assign n24790 = pi647 & n24789;
  assign n24791 = ~pi647 & n24732;
  assign n24792 = pi1157 & ~n24791;
  assign n24793 = pi647 & ~n24789;
  assign n24794 = ~pi647 & ~n24732;
  assign n24795 = ~n24790 & ~n24791;
  assign n24796 = ~n24793 & ~n24794;
  assign n24797 = pi1157 & n63724;
  assign n24798 = ~n24790 & n24792;
  assign n24799 = ~pi647 & n24789;
  assign n24800 = pi647 & n24732;
  assign n24801 = ~pi1157 & ~n24800;
  assign n24802 = ~n24799 & n24801;
  assign n24803 = ~pi647 & ~n24789;
  assign n24804 = pi647 & ~n24732;
  assign n24805 = ~n24803 & ~n24804;
  assign n24806 = ~pi1157 & n24805;
  assign n24807 = pi1157 & ~n63724;
  assign n24808 = ~n24806 & ~n24807;
  assign n24809 = ~n63725 & ~n24802;
  assign n24810 = pi787 & n63726;
  assign n24811 = ~pi787 & ~n24789;
  assign n24812 = pi787 & ~n63726;
  assign n24813 = ~pi787 & n24789;
  assign n24814 = ~n24812 & ~n24813;
  assign n24815 = ~n24810 & ~n24811;
  assign n24816 = ~pi644 & ~n63727;
  assign n24817 = pi715 & ~n24816;
  assign n24818 = ~n11558 & n24732;
  assign n24819 = pi193 & ~n62765;
  assign n24820 = pi739 & n7359;
  assign n24821 = ~n24741 & ~n24820;
  assign n24822 = pi38 & ~n24821;
  assign n24823 = ~pi193 & n62802;
  assign n24824 = pi193 & ~n7351;
  assign n24825 = pi739 & ~n24824;
  assign n24826 = ~n24823 & n24825;
  assign n24827 = ~pi193 & ~pi739;
  assign n24828 = ~n62792 & n24827;
  assign n24829 = ~n24826 & ~n24828;
  assign n24830 = ~pi38 & ~n24829;
  assign n24831 = ~n24822 & ~n24830;
  assign n24832 = n62765 & n24831;
  assign n24833 = ~n24819 & ~n24832;
  assign n24834 = ~n8135 & ~n24833;
  assign n24835 = n8135 & ~n24732;
  assign n24836 = ~n24834 & ~n24835;
  assign n24837 = ~pi785 & ~n24836;
  assign n24838 = ~n8136 & ~n24732;
  assign n24839 = pi609 & n24834;
  assign n24840 = ~n24838 & ~n24839;
  assign n24841 = pi1155 & ~n24840;
  assign n24842 = ~n8148 & ~n24732;
  assign n24843 = ~pi609 & n24834;
  assign n24844 = ~n24842 & ~n24843;
  assign n24845 = ~pi1155 & ~n24844;
  assign n24846 = ~n24841 & ~n24845;
  assign n24847 = pi785 & ~n24846;
  assign n24848 = ~n24837 & ~n24847;
  assign n24849 = ~pi781 & ~n24848;
  assign n24850 = pi618 & n24848;
  assign n24851 = ~pi618 & n24732;
  assign n24852 = pi1154 & ~n24851;
  assign n24853 = ~n24850 & n24852;
  assign n24854 = ~pi618 & n24848;
  assign n24855 = pi618 & n24732;
  assign n24856 = ~pi1154 & ~n24855;
  assign n24857 = ~n24854 & n24856;
  assign n24858 = ~n24853 & ~n24857;
  assign n24859 = pi781 & ~n24858;
  assign n24860 = ~n24849 & ~n24859;
  assign n24861 = ~pi619 & ~n24860;
  assign n24862 = pi619 & ~n24732;
  assign n24863 = ~pi1159 & ~n24862;
  assign n24864 = ~n24861 & n24863;
  assign n24865 = pi619 & ~n24860;
  assign n24866 = ~pi619 & ~n24732;
  assign n24867 = pi1159 & ~n24866;
  assign n24868 = ~n24865 & n24867;
  assign n24869 = pi619 & n24860;
  assign n24870 = ~pi619 & n24732;
  assign n24871 = pi1159 & ~n24870;
  assign n24872 = ~n24869 & n24871;
  assign n24873 = ~pi619 & n24860;
  assign n24874 = pi619 & n24732;
  assign n24875 = ~pi1159 & ~n24874;
  assign n24876 = ~n24873 & n24875;
  assign n24877 = ~n24872 & ~n24876;
  assign n24878 = ~n24864 & ~n24868;
  assign n24879 = pi789 & n63728;
  assign n24880 = ~pi789 & n24860;
  assign n24881 = ~pi789 & ~n24860;
  assign n24882 = pi789 & ~n63728;
  assign n24883 = ~n24881 & ~n24882;
  assign n24884 = ~n24879 & ~n24880;
  assign n24885 = ~n8595 & n63729;
  assign n24886 = n8685 & n24885;
  assign n24887 = n8376 & ~n24732;
  assign n24888 = n8595 & n24732;
  assign n24889 = ~n24885 & ~n24888;
  assign n24890 = ~n8334 & ~n24889;
  assign n24891 = n8334 & n24732;
  assign n24892 = ~n24890 & ~n24891;
  assign n24893 = ~n8376 & n24892;
  assign n24894 = ~n24887 & ~n24893;
  assign n24895 = ~n8376 & ~n24892;
  assign n24896 = n8376 & n24732;
  assign n24897 = ~n24895 & ~n24896;
  assign n24898 = ~n24818 & ~n24886;
  assign n24899 = pi644 & n63730;
  assign n24900 = ~pi644 & n24732;
  assign n24901 = ~pi715 & ~n24900;
  assign n24902 = ~n24899 & n24901;
  assign n24903 = pi1160 & ~n24902;
  assign n24904 = ~n24817 & n24903;
  assign n24905 = pi644 & ~n63727;
  assign n24906 = ~pi715 & ~n24905;
  assign n24907 = ~pi644 & n63730;
  assign n24908 = pi644 & n24732;
  assign n24909 = pi715 & ~n24908;
  assign n24910 = ~n24907 & n24909;
  assign n24911 = ~pi1160 & ~n24910;
  assign n24912 = ~n24906 & n24911;
  assign n24913 = ~n24904 & ~n24912;
  assign n24914 = pi790 & ~n24913;
  assign n24915 = ~n63052 & n24889;
  assign n24916 = ~pi629 & n24782;
  assign n24917 = pi629 & n24786;
  assign n24918 = ~n24916 & ~n24917;
  assign n24919 = ~n24915 & n24918;
  assign n24920 = pi792 & ~n24919;
  assign n24921 = ~pi690 & ~n24831;
  assign n24922 = ~pi193 & ~n62821;
  assign n24923 = pi193 & n7632;
  assign n24924 = ~pi739 & ~n24923;
  assign n24925 = ~n24922 & n24924;
  assign n24926 = pi193 & n7709;
  assign n24927 = ~pi193 & n62851;
  assign n24928 = pi739 & ~n24927;
  assign n24929 = ~n24926 & n24928;
  assign n24930 = pi39 & ~n24929;
  assign n24931 = ~n24925 & n24930;
  assign n24932 = pi193 & n7855;
  assign n24933 = ~pi193 & n7832;
  assign n24934 = ~pi739 & ~n24933;
  assign n24935 = ~n24932 & n24934;
  assign n24936 = ~pi193 & ~n7861;
  assign n24937 = pi193 & ~n7868;
  assign n24938 = pi739 & ~n24937;
  assign n24939 = ~n24936 & n24938;
  assign n24940 = ~pi39 & ~n24939;
  assign n24941 = ~pi193 & n7861;
  assign n24942 = pi193 & n7868;
  assign n24943 = pi739 & ~n24942;
  assign n24944 = ~n24941 & n24943;
  assign n24945 = pi193 & ~n7855;
  assign n24946 = ~pi193 & ~n7832;
  assign n24947 = ~pi739 & ~n24946;
  assign n24948 = ~pi739 & ~n24945;
  assign n24949 = ~n24946 & n24948;
  assign n24950 = ~n24945 & n24947;
  assign n24951 = ~n24944 & ~n63731;
  assign n24952 = ~pi39 & ~n24951;
  assign n24953 = ~n24935 & n24940;
  assign n24954 = ~pi38 & ~n63732;
  assign n24955 = ~n24931 & n24954;
  assign n24956 = ~pi739 & n13901;
  assign n24957 = ~n7744 & ~n24956;
  assign n24958 = ~pi39 & ~n24957;
  assign n24959 = ~pi193 & ~n24958;
  assign n24960 = ~n7565 & ~n24507;
  assign n24961 = pi193 & ~n24960;
  assign n24962 = n7356 & n24961;
  assign n24963 = pi38 & ~n24962;
  assign n24964 = ~n24959 & n24963;
  assign n24965 = pi690 & ~n24964;
  assign n24966 = ~n24955 & n24965;
  assign n24967 = n62765 & ~n24966;
  assign n24968 = ~n24921 & n24967;
  assign n24969 = ~n24819 & ~n24968;
  assign n24970 = ~pi625 & n24969;
  assign n24971 = pi625 & n24833;
  assign n24972 = ~pi1153 & ~n24971;
  assign n24973 = ~n24970 & n24972;
  assign n24974 = ~pi608 & ~n24750;
  assign n24975 = ~n24973 & n24974;
  assign n24976 = pi625 & n24969;
  assign n24977 = ~pi625 & n24833;
  assign n24978 = pi1153 & ~n24977;
  assign n24979 = ~n24976 & n24978;
  assign n24980 = pi608 & ~n24754;
  assign n24981 = ~n24979 & n24980;
  assign n24982 = ~n24975 & ~n24981;
  assign n24983 = pi778 & ~n24982;
  assign n24984 = ~pi778 & n24969;
  assign n24985 = ~n24983 & ~n24984;
  assign n24986 = ~pi609 & ~n24985;
  assign n24987 = pi609 & n24757;
  assign n24988 = ~pi1155 & ~n24987;
  assign n24989 = ~n24986 & n24988;
  assign n24990 = ~pi660 & ~n24841;
  assign n24991 = ~n24989 & n24990;
  assign n24992 = pi609 & ~n24985;
  assign n24993 = ~pi609 & n24757;
  assign n24994 = pi1155 & ~n24993;
  assign n24995 = ~n24992 & n24994;
  assign n24996 = pi660 & ~n24845;
  assign n24997 = ~n24995 & n24996;
  assign n24998 = ~n24991 & ~n24997;
  assign n24999 = pi785 & ~n24998;
  assign n25000 = ~pi785 & ~n24985;
  assign n25001 = ~n24999 & ~n25000;
  assign n25002 = pi618 & ~n25001;
  assign n25003 = ~pi618 & ~n63721;
  assign n25004 = pi1154 & ~n25003;
  assign n25005 = ~n25002 & n25004;
  assign n25006 = pi627 & ~n24857;
  assign n25007 = ~n25005 & n25006;
  assign n25008 = ~pi618 & ~n25001;
  assign n25009 = pi618 & ~n63721;
  assign n25010 = ~pi1154 & ~n25009;
  assign n25011 = ~n25008 & n25010;
  assign n25012 = ~pi627 & ~n24853;
  assign n25013 = ~n25011 & n25012;
  assign n25014 = pi781 & ~n25013;
  assign n25015 = ~n25007 & n25014;
  assign n25016 = ~n11431 & ~n63722;
  assign n25017 = ~n62884 & ~n63728;
  assign n25018 = ~n25016 & ~n25017;
  assign n25019 = pi789 & ~n25018;
  assign n25020 = ~pi781 & n25001;
  assign n25021 = ~n25019 & ~n25020;
  assign n25022 = ~n25015 & n25021;
  assign n25023 = n11434 & n25018;
  assign n25024 = ~n25022 & ~n25023;
  assign n25025 = ~n25007 & ~n25013;
  assign n25026 = pi781 & ~n25025;
  assign n25027 = ~pi781 & ~n25001;
  assign n25028 = ~n25026 & ~n25027;
  assign n25029 = ~pi619 & ~n25028;
  assign n25030 = pi619 & n63722;
  assign n25031 = ~pi1159 & ~n25030;
  assign n25032 = ~n25029 & n25031;
  assign n25033 = ~pi648 & ~n24872;
  assign n25034 = ~n25032 & n25033;
  assign n25035 = pi619 & ~n25028;
  assign n25036 = ~pi619 & n63722;
  assign n25037 = pi1159 & ~n25036;
  assign n25038 = ~n25035 & n25037;
  assign n25039 = pi648 & ~n24876;
  assign n25040 = ~n25038 & n25039;
  assign n25041 = pi789 & ~n25040;
  assign n25042 = pi789 & ~n25034;
  assign n25043 = ~n25040 & n25042;
  assign n25044 = ~n25034 & n25041;
  assign n25045 = ~pi789 & n25028;
  assign n25046 = n62894 & ~n25045;
  assign n25047 = ~n63733 & n25046;
  assign n25048 = n62894 & ~n25024;
  assign n25049 = ~pi626 & ~n63729;
  assign n25050 = pi626 & ~n24732;
  assign n25051 = n8301 & ~n25050;
  assign n25052 = ~n25049 & n25051;
  assign n25053 = n8525 & ~n63723;
  assign n25054 = pi626 & ~n63729;
  assign n25055 = ~pi626 & ~n24732;
  assign n25056 = n8300 & ~n25055;
  assign n25057 = ~n25054 & n25056;
  assign n25058 = ~n25053 & ~n25057;
  assign n25059 = ~n25052 & ~n25053;
  assign n25060 = ~n25057 & n25059;
  assign n25061 = ~n25052 & n25058;
  assign n25062 = pi788 & ~n63735;
  assign n25063 = ~n63030 & ~n25062;
  assign n25064 = ~n63734 & n25063;
  assign n25065 = ~n24920 & ~n25064;
  assign n25066 = ~n8651 & ~n25065;
  assign n25067 = ~n8413 & ~n24891;
  assign n25068 = ~n8413 & n24892;
  assign n25069 = ~n24890 & n25067;
  assign n25070 = n8373 & n63724;
  assign n25071 = ~pi630 & n63725;
  assign n25072 = n8374 & ~n24805;
  assign n25073 = pi630 & n24802;
  assign n25074 = ~n63737 & ~n63738;
  assign n25075 = ~n63736 & n25074;
  assign n25076 = pi787 & ~n25075;
  assign n25077 = ~pi644 & n24911;
  assign n25078 = pi644 & n24903;
  assign n25079 = n14029 & ~n24902;
  assign n25080 = pi790 & ~n63739;
  assign n25081 = pi790 & ~n25077;
  assign n25082 = ~n63739 & n25081;
  assign n25083 = ~n25077 & n25080;
  assign n25084 = ~n25076 & ~n63740;
  assign n25085 = ~n25066 & ~n25076;
  assign n25086 = ~n63740 & n25085;
  assign n25087 = ~n25066 & n25084;
  assign n25088 = ~n24914 & ~n63741;
  assign n25089 = n62455 & ~n25088;
  assign n25090 = ~pi193 & ~n62455;
  assign n25091 = ~pi832 & ~n25090;
  assign n25092 = ~n25089 & n25091;
  assign po350 = ~n24731 & ~n25092;
  assign n25094 = pi194 & ~n62765;
  assign n25095 = ~pi194 & n10343;
  assign n25096 = pi194 & n14285;
  assign n25097 = ~n25095 & ~n25096;
  assign n25098 = pi748 & ~n25097;
  assign n25099 = ~pi194 & ~n8091;
  assign n25100 = ~pi748 & ~n25099;
  assign n25101 = ~n25098 & ~n25100;
  assign n25102 = n62765 & ~n25101;
  assign n25103 = ~n25094 & ~n25102;
  assign n25104 = ~n8135 & ~n25103;
  assign n25105 = ~pi194 & ~n8098;
  assign n25106 = n8135 & ~n25105;
  assign n25107 = ~n25104 & ~n25106;
  assign n25108 = ~pi785 & ~n25107;
  assign n25109 = ~n8136 & ~n25105;
  assign n25110 = pi609 & n25104;
  assign n25111 = ~n25109 & ~n25110;
  assign n25112 = pi1155 & ~n25111;
  assign n25113 = ~n8148 & ~n25105;
  assign n25114 = ~pi609 & n25104;
  assign n25115 = ~n25113 & ~n25114;
  assign n25116 = ~pi1155 & ~n25115;
  assign n25117 = ~n25112 & ~n25116;
  assign n25118 = pi785 & ~n25117;
  assign n25119 = ~n25108 & ~n25118;
  assign n25120 = ~pi781 & ~n25119;
  assign n25121 = pi618 & n25119;
  assign n25122 = ~pi618 & n25105;
  assign n25123 = pi1154 & ~n25122;
  assign n25124 = ~n25121 & n25123;
  assign n25125 = ~pi618 & n25119;
  assign n25126 = pi618 & n25105;
  assign n25127 = ~pi1154 & ~n25126;
  assign n25128 = ~n25125 & n25127;
  assign n25129 = ~n25124 & ~n25128;
  assign n25130 = pi781 & ~n25129;
  assign n25131 = ~n25120 & ~n25130;
  assign n25132 = ~pi789 & ~n25131;
  assign n25133 = ~pi619 & n25131;
  assign n25134 = pi619 & n25105;
  assign n25135 = ~pi1159 & ~n25134;
  assign n25136 = ~n25133 & n25135;
  assign n25137 = pi619 & n25131;
  assign n25138 = ~pi619 & n25105;
  assign n25139 = pi1159 & ~n25138;
  assign n25140 = ~n25137 & n25139;
  assign n25141 = ~n25136 & ~n25140;
  assign n25142 = pi789 & ~n25141;
  assign n25143 = ~n25132 & ~n25142;
  assign n25144 = ~n8595 & n25143;
  assign n25145 = n8595 & n25105;
  assign n25146 = ~n25144 & ~n25145;
  assign n25147 = ~n8334 & ~n25146;
  assign n25148 = n8334 & n25105;
  assign n25149 = ~n25147 & ~n25148;
  assign n25150 = ~n8376 & ~n25149;
  assign n25151 = n8376 & n25105;
  assign n25152 = n8376 & ~n25105;
  assign n25153 = ~n8376 & n25149;
  assign n25154 = ~n25152 & ~n25153;
  assign n25155 = ~n25150 & ~n25151;
  assign n25156 = pi644 & n63742;
  assign n25157 = ~pi644 & n25105;
  assign n25158 = n16177 & ~n25157;
  assign n25159 = ~n25156 & n25158;
  assign n25160 = ~pi644 & n63742;
  assign n25161 = pi644 & n25105;
  assign n25162 = n16172 & ~n25161;
  assign n25163 = ~n25160 & n25162;
  assign n25164 = n8257 & ~n25105;
  assign n25165 = pi194 & ~n14367;
  assign n25166 = ~pi194 & n14370;
  assign n25167 = pi730 & ~n25166;
  assign n25168 = ~pi730 & n25099;
  assign n25169 = n62765 & ~n25168;
  assign n25170 = ~n25167 & n25169;
  assign n25171 = ~n25165 & ~n25170;
  assign n25172 = ~pi778 & ~n25171;
  assign n25173 = ~pi625 & n25171;
  assign n25174 = pi625 & n25105;
  assign n25175 = ~pi1153 & ~n25174;
  assign n25176 = ~n25173 & n25175;
  assign n25177 = pi625 & n25171;
  assign n25178 = ~pi625 & n25105;
  assign n25179 = pi1153 & ~n25178;
  assign n25180 = ~n25177 & n25179;
  assign n25181 = ~n25176 & ~n25180;
  assign n25182 = pi778 & ~n25181;
  assign n25183 = ~n25172 & ~n25182;
  assign n25184 = ~n62880 & ~n25183;
  assign n25185 = n62880 & ~n25105;
  assign n25186 = ~n62880 & n25183;
  assign n25187 = n62880 & n25105;
  assign n25188 = ~n25186 & ~n25187;
  assign n25189 = ~n25184 & ~n25185;
  assign n25190 = ~n62882 & ~n63743;
  assign n25191 = n62882 & n25105;
  assign n25192 = n62882 & ~n25105;
  assign n25193 = ~n62882 & n63743;
  assign n25194 = ~n25192 & ~n25193;
  assign n25195 = ~n25190 & ~n25191;
  assign n25196 = ~n8257 & ~n63744;
  assign n25197 = ~n8257 & n63744;
  assign n25198 = n8257 & n25105;
  assign n25199 = ~n25197 & ~n25198;
  assign n25200 = ~n25164 & ~n25196;
  assign n25201 = ~n8303 & ~n63745;
  assign n25202 = n8303 & n25105;
  assign n25203 = n8303 & ~n25105;
  assign n25204 = ~n8303 & n63745;
  assign n25205 = ~n25203 & ~n25204;
  assign n25206 = ~n25201 & ~n25202;
  assign n25207 = ~n62892 & n63746;
  assign n25208 = n62892 & n25105;
  assign n25209 = pi628 & n63746;
  assign n25210 = ~pi628 & n25105;
  assign n25211 = pi1156 & ~n25210;
  assign n25212 = ~n25209 & n25211;
  assign n25213 = ~pi628 & n63746;
  assign n25214 = pi628 & n25105;
  assign n25215 = ~pi1156 & ~n25214;
  assign n25216 = ~n25213 & n25215;
  assign n25217 = pi628 & ~n25105;
  assign n25218 = ~pi628 & ~n63746;
  assign n25219 = ~n25217 & ~n25218;
  assign n25220 = ~pi1156 & n25219;
  assign n25221 = ~pi628 & ~n25105;
  assign n25222 = pi628 & ~n63746;
  assign n25223 = ~n25221 & ~n25222;
  assign n25224 = pi1156 & n25223;
  assign n25225 = ~n25220 & ~n25224;
  assign n25226 = ~n25212 & ~n25216;
  assign n25227 = pi792 & ~n63747;
  assign n25228 = ~pi792 & n63746;
  assign n25229 = ~n25227 & ~n25228;
  assign n25230 = ~pi792 & ~n63746;
  assign n25231 = pi792 & n63747;
  assign n25232 = ~n25230 & ~n25231;
  assign n25233 = ~n25207 & ~n25208;
  assign n25234 = ~pi647 & ~n63748;
  assign n25235 = pi647 & n25105;
  assign n25236 = ~pi1157 & ~n25235;
  assign n25237 = pi647 & ~n25105;
  assign n25238 = ~pi647 & n63748;
  assign n25239 = ~n25234 & ~n25235;
  assign n25240 = ~n25237 & ~n25238;
  assign n25241 = ~pi1157 & n63749;
  assign n25242 = ~n25234 & n25236;
  assign n25243 = pi647 & ~n63748;
  assign n25244 = ~pi647 & n25105;
  assign n25245 = pi1157 & ~n25244;
  assign n25246 = ~n25243 & n25245;
  assign n25247 = pi787 & ~n25246;
  assign n25248 = ~pi1157 & ~n63749;
  assign n25249 = ~n25243 & ~n25244;
  assign n25250 = pi1157 & ~n25249;
  assign n25251 = ~n25248 & ~n25250;
  assign n25252 = ~n63750 & ~n25246;
  assign n25253 = pi787 & ~n63751;
  assign n25254 = ~n63750 & n25247;
  assign n25255 = ~pi787 & ~n63748;
  assign n25256 = ~n63036 & ~n25255;
  assign n25257 = ~n63752 & n25256;
  assign n25258 = ~n25163 & ~n25257;
  assign n25259 = ~n25159 & ~n25163;
  assign n25260 = ~n25257 & n25259;
  assign n25261 = ~n25159 & n25258;
  assign n25262 = pi790 & ~n63753;
  assign n25263 = ~n8413 & n25149;
  assign n25264 = n8374 & n63749;
  assign n25265 = n8373 & n25249;
  assign n25266 = ~pi630 & n25246;
  assign n25267 = ~n25264 & ~n63754;
  assign n25268 = ~n25263 & ~n25264;
  assign n25269 = ~n63754 & n25268;
  assign n25270 = ~n25263 & n25267;
  assign n25271 = pi787 & ~n63755;
  assign n25272 = ~n63052 & n25146;
  assign n25273 = n8332 & ~n25214;
  assign n25274 = n8332 & ~n25219;
  assign n25275 = ~n25213 & n25273;
  assign n25276 = n8331 & ~n25210;
  assign n25277 = n8331 & ~n25223;
  assign n25278 = ~n25209 & n25276;
  assign n25279 = ~n63756 & ~n63757;
  assign n25280 = ~n25272 & n25279;
  assign n25281 = pi792 & ~n25280;
  assign n25282 = n12979 & n25143;
  assign n25283 = ~pi641 & n63745;
  assign n25284 = pi641 & ~n25105;
  assign n25285 = n8417 & ~n25284;
  assign n25286 = ~n25283 & n25285;
  assign n25287 = pi641 & n63745;
  assign n25288 = ~pi641 & ~n25105;
  assign n25289 = n8416 & ~n25288;
  assign n25290 = ~n25287 & n25289;
  assign n25291 = ~n25286 & ~n25290;
  assign n25292 = ~n25282 & n25291;
  assign n25293 = pi788 & ~n25292;
  assign n25294 = pi619 & n63744;
  assign n25295 = ~pi1159 & ~n25294;
  assign n25296 = ~pi648 & ~n25140;
  assign n25297 = ~n25295 & n25296;
  assign n25298 = ~pi619 & n63744;
  assign n25299 = pi1159 & ~n25298;
  assign n25300 = pi648 & ~n25299;
  assign n25301 = pi648 & ~n25136;
  assign n25302 = ~n25299 & n25301;
  assign n25303 = ~n25136 & n25300;
  assign n25304 = ~n25297 & ~n63758;
  assign n25305 = pi789 & ~n25304;
  assign n25306 = pi618 & ~n63743;
  assign n25307 = ~pi1154 & ~n25306;
  assign n25308 = ~pi627 & ~n25124;
  assign n25309 = ~n25307 & n25308;
  assign n25310 = ~pi618 & ~n63743;
  assign n25311 = pi1154 & ~n25310;
  assign n25312 = pi627 & ~n25128;
  assign n25313 = ~n25311 & n25312;
  assign n25314 = ~n25309 & ~n25313;
  assign n25315 = pi781 & ~n25314;
  assign n25316 = ~pi618 & n25308;
  assign n25317 = pi618 & n25312;
  assign n25318 = pi781 & ~n25317;
  assign n25319 = ~n25316 & n25318;
  assign n25320 = ~pi730 & n25101;
  assign n25321 = ~pi194 & n10353;
  assign n25322 = pi194 & ~n14472;
  assign n25323 = ~pi748 & ~n25322;
  assign n25324 = ~n25321 & n25323;
  assign n25325 = pi194 & n10363;
  assign n25326 = ~pi194 & ~n62980;
  assign n25327 = pi748 & ~n25326;
  assign n25328 = ~n25325 & n25327;
  assign n25329 = pi730 & ~n25328;
  assign n25330 = pi194 & ~n10363;
  assign n25331 = ~pi194 & n62980;
  assign n25332 = pi748 & ~n25331;
  assign n25333 = ~n25330 & n25332;
  assign n25334 = ~pi194 & ~n10353;
  assign n25335 = pi194 & n14472;
  assign n25336 = ~pi748 & ~n25335;
  assign n25337 = ~n25334 & n25336;
  assign n25338 = ~n25333 & ~n25337;
  assign n25339 = pi730 & ~n25338;
  assign n25340 = ~n25324 & n25329;
  assign n25341 = n62765 & ~n63759;
  assign n25342 = n62765 & ~n25320;
  assign n25343 = ~n63759 & n25342;
  assign n25344 = ~n25320 & n25341;
  assign n25345 = ~n25094 & ~n63760;
  assign n25346 = pi625 & n25345;
  assign n25347 = ~pi625 & n25103;
  assign n25348 = pi1153 & ~n25347;
  assign n25349 = ~n25346 & n25348;
  assign n25350 = pi608 & ~n25176;
  assign n25351 = ~n25349 & n25350;
  assign n25352 = ~pi625 & n25345;
  assign n25353 = pi625 & n25103;
  assign n25354 = ~pi1153 & ~n25353;
  assign n25355 = ~n25352 & n25354;
  assign n25356 = ~pi608 & ~n25180;
  assign n25357 = ~n25355 & n25356;
  assign n25358 = ~n25351 & ~n25357;
  assign n25359 = pi778 & ~n25358;
  assign n25360 = ~pi778 & n25345;
  assign n25361 = ~pi778 & ~n25345;
  assign n25362 = pi778 & ~n25357;
  assign n25363 = ~n25351 & n25362;
  assign n25364 = ~n25361 & ~n25363;
  assign n25365 = ~n25359 & ~n25360;
  assign n25366 = ~pi609 & n63761;
  assign n25367 = pi609 & n25183;
  assign n25368 = ~pi1155 & ~n25367;
  assign n25369 = ~n25366 & n25368;
  assign n25370 = ~pi660 & ~n25112;
  assign n25371 = ~n25369 & n25370;
  assign n25372 = pi609 & n63761;
  assign n25373 = ~pi609 & n25183;
  assign n25374 = pi1155 & ~n25373;
  assign n25375 = ~n25372 & n25374;
  assign n25376 = pi660 & ~n25116;
  assign n25377 = ~n25375 & n25376;
  assign n25378 = pi785 & ~n25377;
  assign n25379 = ~n25371 & n25378;
  assign n25380 = ~pi785 & ~n63761;
  assign n25381 = ~n25371 & ~n25377;
  assign n25382 = pi785 & ~n25381;
  assign n25383 = ~pi785 & n63761;
  assign n25384 = ~n25382 & ~n25383;
  assign n25385 = ~n25379 & ~n25380;
  assign n25386 = ~n25319 & ~n63762;
  assign n25387 = pi618 & ~n63762;
  assign n25388 = n25311 & ~n25387;
  assign n25389 = n25312 & ~n25388;
  assign n25390 = ~n25309 & ~n25389;
  assign n25391 = pi781 & ~n25390;
  assign n25392 = pi781 & ~n25316;
  assign n25393 = ~n63762 & ~n25392;
  assign n25394 = ~n25391 & ~n25393;
  assign n25395 = ~pi618 & ~n63762;
  assign n25396 = n25307 & ~n25395;
  assign n25397 = n25308 & ~n25396;
  assign n25398 = ~n25389 & ~n25397;
  assign n25399 = pi781 & ~n25398;
  assign n25400 = ~pi781 & ~n63762;
  assign n25401 = ~n25399 & ~n25400;
  assign n25402 = ~n25315 & ~n25386;
  assign n25403 = ~pi619 & n25296;
  assign n25404 = pi619 & n25301;
  assign n25405 = n11422 & ~n25136;
  assign n25406 = pi789 & ~n63764;
  assign n25407 = ~n25403 & n25406;
  assign n25408 = ~n63763 & ~n25407;
  assign n25409 = ~pi619 & ~n63763;
  assign n25410 = n25295 & ~n25409;
  assign n25411 = n25296 & ~n25410;
  assign n25412 = pi619 & ~n63763;
  assign n25413 = n25299 & ~n25412;
  assign n25414 = n25301 & ~n25413;
  assign n25415 = ~n25411 & ~n25414;
  assign n25416 = pi789 & ~n25415;
  assign n25417 = ~pi789 & ~n63763;
  assign n25418 = ~n25416 & ~n25417;
  assign n25419 = ~n25305 & ~n25408;
  assign n25420 = n62894 & ~n63765;
  assign n25421 = ~n63030 & ~n25420;
  assign n25422 = ~n25293 & n25421;
  assign n25423 = ~pi788 & n63765;
  assign n25424 = ~pi626 & n63765;
  assign n25425 = pi626 & n63745;
  assign n25426 = ~pi641 & ~n25425;
  assign n25427 = ~n25424 & n25426;
  assign n25428 = ~pi626 & ~n25143;
  assign n25429 = pi626 & ~n25105;
  assign n25430 = pi641 & ~n25429;
  assign n25431 = ~n25428 & n25430;
  assign n25432 = ~pi1158 & ~n25431;
  assign n25433 = ~n25427 & n25432;
  assign n25434 = pi626 & n63765;
  assign n25435 = ~pi626 & n63745;
  assign n25436 = pi641 & ~n25435;
  assign n25437 = ~n25434 & n25436;
  assign n25438 = pi626 & ~n25143;
  assign n25439 = ~pi626 & ~n25105;
  assign n25440 = ~pi641 & ~n25439;
  assign n25441 = ~n25438 & n25440;
  assign n25442 = pi1158 & ~n25441;
  assign n25443 = ~n25437 & n25442;
  assign n25444 = ~n25433 & ~n25443;
  assign n25445 = pi788 & ~n25444;
  assign n25446 = ~n25423 & ~n25445;
  assign n25447 = ~n25293 & ~n25420;
  assign n25448 = ~pi628 & n63766;
  assign n25449 = pi628 & ~n25146;
  assign n25450 = ~pi1156 & ~n25449;
  assign n25451 = ~n25448 & n25450;
  assign n25452 = ~pi629 & ~n25212;
  assign n25453 = ~n25451 & n25452;
  assign n25454 = pi628 & n63766;
  assign n25455 = ~pi628 & ~n25146;
  assign n25456 = pi1156 & ~n25455;
  assign n25457 = ~n25454 & n25456;
  assign n25458 = pi629 & ~n25216;
  assign n25459 = ~n25457 & n25458;
  assign n25460 = ~n25453 & ~n25459;
  assign n25461 = pi792 & ~n25460;
  assign n25462 = ~pi792 & n63766;
  assign n25463 = ~n25461 & ~n25462;
  assign n25464 = ~n25281 & ~n25422;
  assign n25465 = ~n25281 & n63766;
  assign n25466 = n63030 & n25280;
  assign n25467 = ~n8651 & ~n25466;
  assign n25468 = ~n25465 & n25467;
  assign n25469 = ~n8651 & n63767;
  assign n25470 = ~pi647 & ~n63767;
  assign n25471 = pi647 & ~n25149;
  assign n25472 = ~pi1157 & ~n25471;
  assign n25473 = ~n25470 & n25472;
  assign n25474 = ~pi630 & ~n25246;
  assign n25475 = ~n25473 & n25474;
  assign n25476 = pi647 & ~n63767;
  assign n25477 = ~pi647 & ~n25149;
  assign n25478 = pi1157 & ~n25477;
  assign n25479 = ~n25476 & n25478;
  assign n25480 = pi630 & ~n63750;
  assign n25481 = ~n25479 & n25480;
  assign n25482 = ~n25475 & ~n25481;
  assign n25483 = pi787 & ~n25482;
  assign n25484 = ~pi787 & ~n63767;
  assign n25485 = ~n25483 & ~n25484;
  assign n25486 = ~n25271 & ~n63768;
  assign n25487 = ~n11547 & n63769;
  assign n25488 = n62455 & ~n25487;
  assign n25489 = n62455 & ~n25262;
  assign n25490 = ~n25487 & n25489;
  assign n25491 = pi644 & ~n63769;
  assign n25492 = ~pi787 & n63748;
  assign n25493 = pi787 & n63751;
  assign n25494 = ~n25492 & ~n25493;
  assign n25495 = ~pi644 & n25494;
  assign n25496 = pi715 & ~n25495;
  assign n25497 = ~n25491 & n25496;
  assign n25498 = ~pi715 & ~n25157;
  assign n25499 = ~n25156 & n25498;
  assign n25500 = pi1160 & ~n25499;
  assign n25501 = ~n25497 & n25500;
  assign n25502 = ~pi644 & ~n63769;
  assign n25503 = pi644 & n25494;
  assign n25504 = ~pi715 & ~n25503;
  assign n25505 = ~n25502 & n25504;
  assign n25506 = pi715 & ~n25161;
  assign n25507 = ~n25160 & n25506;
  assign n25508 = ~pi1160 & ~n25507;
  assign n25509 = ~n25505 & n25508;
  assign n25510 = pi790 & ~n25509;
  assign n25511 = pi790 & ~n25501;
  assign n25512 = ~n25509 & n25511;
  assign n25513 = ~n25501 & n25510;
  assign n25514 = ~pi790 & n63769;
  assign n25515 = n62455 & ~n25514;
  assign n25516 = ~n63771 & n25515;
  assign n25517 = ~n25262 & n25488;
  assign n25518 = ~pi194 & ~n62455;
  assign n25519 = ~pi832 & ~n25518;
  assign n25520 = ~n63770 & n25519;
  assign n25521 = ~pi194 & ~n2923;
  assign n25522 = pi748 & n7316;
  assign n25523 = ~n25521 & ~n25522;
  assign n25524 = ~n8420 & ~n25523;
  assign n25525 = ~pi785 & ~n25524;
  assign n25526 = ~n8425 & ~n25523;
  assign n25527 = pi1155 & ~n25526;
  assign n25528 = ~n8428 & n25524;
  assign n25529 = ~pi1155 & ~n25528;
  assign n25530 = ~n25527 & ~n25529;
  assign n25531 = pi785 & ~n25530;
  assign n25532 = ~n25525 & ~n25531;
  assign n25533 = ~pi781 & ~n25532;
  assign n25534 = ~n8435 & n25532;
  assign n25535 = pi1154 & ~n25534;
  assign n25536 = ~n8438 & n25532;
  assign n25537 = ~pi1154 & ~n25536;
  assign n25538 = ~n25535 & ~n25537;
  assign n25539 = pi781 & ~n25538;
  assign n25540 = ~n25533 & ~n25539;
  assign n25541 = ~pi619 & ~n25540;
  assign n25542 = pi619 & ~n25521;
  assign n25543 = ~pi1159 & ~n25542;
  assign n25544 = ~n25541 & n25543;
  assign n25545 = pi619 & ~n25540;
  assign n25546 = ~pi619 & ~n25521;
  assign n25547 = pi1159 & ~n25546;
  assign n25548 = ~n25545 & n25547;
  assign n25549 = pi619 & n25540;
  assign n25550 = ~pi619 & n25521;
  assign n25551 = pi1159 & ~n25550;
  assign n25552 = ~n25549 & n25551;
  assign n25553 = ~pi619 & n25540;
  assign n25554 = pi619 & n25521;
  assign n25555 = ~pi1159 & ~n25554;
  assign n25556 = ~n25553 & n25555;
  assign n25557 = ~n25552 & ~n25556;
  assign n25558 = ~n25544 & ~n25548;
  assign n25559 = pi789 & n63772;
  assign n25560 = ~pi789 & n25540;
  assign n25561 = ~pi789 & ~n25540;
  assign n25562 = pi789 & ~n63772;
  assign n25563 = ~n25561 & ~n25562;
  assign n25564 = ~n25559 & ~n25560;
  assign n25565 = ~n8595 & n63773;
  assign n25566 = n8595 & n25521;
  assign n25567 = ~n8595 & ~n63773;
  assign n25568 = n8595 & ~n25521;
  assign n25569 = ~n25567 & ~n25568;
  assign n25570 = ~n25565 & ~n25566;
  assign n25571 = ~n8334 & n63774;
  assign n25572 = n8334 & n25521;
  assign n25573 = ~n8413 & ~n25572;
  assign n25574 = ~n25571 & ~n25572;
  assign n25575 = ~n8413 & n25574;
  assign n25576 = ~n25571 & n25573;
  assign n25577 = pi730 & n7564;
  assign n25578 = ~n25521 & ~n25577;
  assign n25579 = ~pi778 & n25578;
  assign n25580 = ~pi625 & n25577;
  assign n25581 = ~n25578 & ~n25580;
  assign n25582 = pi1153 & ~n25581;
  assign n25583 = ~pi1153 & ~n25521;
  assign n25584 = ~n25580 & n25583;
  assign n25585 = ~n25582 & ~n25584;
  assign n25586 = pi778 & ~n25585;
  assign n25587 = ~n25579 & ~n25586;
  assign n25588 = ~n8490 & n25587;
  assign n25589 = ~n8492 & n25588;
  assign n25590 = ~n8494 & n25589;
  assign n25591 = ~n8496 & n25590;
  assign n25592 = ~n8508 & n25591;
  assign n25593 = pi647 & ~n25592;
  assign n25594 = ~pi647 & ~n25521;
  assign n25595 = ~n25593 & ~n25594;
  assign n25596 = n8373 & ~n25595;
  assign n25597 = ~pi647 & n25592;
  assign n25598 = pi647 & n25521;
  assign n25599 = ~pi1157 & ~n25598;
  assign n25600 = ~n25597 & n25599;
  assign n25601 = pi630 & n25600;
  assign n25602 = ~n25596 & ~n25601;
  assign n25603 = ~n63775 & n25602;
  assign n25604 = pi787 & ~n25603;
  assign n25605 = ~pi626 & ~n63773;
  assign n25606 = pi626 & ~n25521;
  assign n25607 = n8301 & ~n25606;
  assign n25608 = ~n25605 & n25607;
  assign n25609 = n8525 & n25590;
  assign n25610 = pi626 & ~n63773;
  assign n25611 = ~pi626 & ~n25521;
  assign n25612 = n8300 & ~n25611;
  assign n25613 = ~n25610 & n25612;
  assign n25614 = ~n25609 & ~n25613;
  assign n25615 = ~n25608 & ~n25609;
  assign n25616 = ~n25613 & n25615;
  assign n25617 = ~n25608 & n25614;
  assign n25618 = pi788 & ~n63776;
  assign n25619 = ~n7187 & ~n25578;
  assign n25620 = pi625 & n25619;
  assign n25621 = n25523 & ~n25619;
  assign n25622 = ~n25620 & ~n25621;
  assign n25623 = n25583 & ~n25622;
  assign n25624 = ~pi608 & ~n25582;
  assign n25625 = ~n25623 & n25624;
  assign n25626 = pi1153 & n25523;
  assign n25627 = ~n25620 & n25626;
  assign n25628 = pi608 & ~n25584;
  assign n25629 = ~n25627 & n25628;
  assign n25630 = ~n25625 & ~n25629;
  assign n25631 = pi778 & ~n25630;
  assign n25632 = ~pi778 & ~n25621;
  assign n25633 = ~n25631 & ~n25632;
  assign n25634 = ~pi609 & ~n25633;
  assign n25635 = pi609 & n25587;
  assign n25636 = ~pi1155 & ~n25635;
  assign n25637 = ~n25634 & n25636;
  assign n25638 = ~pi660 & ~n25527;
  assign n25639 = ~n25637 & n25638;
  assign n25640 = pi609 & ~n25633;
  assign n25641 = ~pi609 & n25587;
  assign n25642 = pi1155 & ~n25641;
  assign n25643 = ~n25640 & n25642;
  assign n25644 = pi660 & ~n25529;
  assign n25645 = ~n25643 & n25644;
  assign n25646 = ~n25639 & ~n25645;
  assign n25647 = pi785 & ~n25646;
  assign n25648 = ~pi785 & ~n25633;
  assign n25649 = ~n25647 & ~n25648;
  assign n25650 = pi618 & ~n25649;
  assign n25651 = ~pi618 & n25588;
  assign n25652 = pi1154 & ~n25651;
  assign n25653 = ~n25650 & n25652;
  assign n25654 = pi627 & ~n25537;
  assign n25655 = ~n25653 & n25654;
  assign n25656 = ~pi618 & ~n25649;
  assign n25657 = pi618 & n25588;
  assign n25658 = ~pi1154 & ~n25657;
  assign n25659 = ~n25656 & n25658;
  assign n25660 = ~pi627 & ~n25535;
  assign n25661 = ~n25659 & n25660;
  assign n25662 = pi781 & ~n25661;
  assign n25663 = ~n25655 & n25662;
  assign n25664 = ~n11431 & ~n25589;
  assign n25665 = ~n62884 & ~n63772;
  assign n25666 = ~n25664 & ~n25665;
  assign n25667 = pi789 & ~n25666;
  assign n25668 = ~pi781 & n25649;
  assign n25669 = ~n25667 & ~n25668;
  assign n25670 = ~n25663 & n25669;
  assign n25671 = n11434 & n25666;
  assign n25672 = ~n25670 & ~n25671;
  assign n25673 = ~n25655 & ~n25661;
  assign n25674 = pi781 & ~n25673;
  assign n25675 = ~pi781 & ~n25649;
  assign n25676 = ~n25674 & ~n25675;
  assign n25677 = ~pi619 & ~n25676;
  assign n25678 = pi619 & n25589;
  assign n25679 = ~pi1159 & ~n25678;
  assign n25680 = ~n25677 & n25679;
  assign n25681 = ~pi648 & ~n25552;
  assign n25682 = ~n25680 & n25681;
  assign n25683 = pi619 & ~n25676;
  assign n25684 = ~pi619 & n25589;
  assign n25685 = pi1159 & ~n25684;
  assign n25686 = ~n25683 & n25685;
  assign n25687 = pi648 & ~n25556;
  assign n25688 = ~n25686 & n25687;
  assign n25689 = pi789 & ~n25688;
  assign n25690 = pi789 & ~n25682;
  assign n25691 = ~n25688 & n25690;
  assign n25692 = ~n25682 & n25689;
  assign n25693 = ~pi789 & n25676;
  assign n25694 = n62894 & ~n25693;
  assign n25695 = ~n63777 & n25694;
  assign n25696 = n62894 & ~n25672;
  assign n25697 = ~n25618 & ~n63778;
  assign n25698 = ~n63030 & ~n25697;
  assign n25699 = n8498 & n63774;
  assign n25700 = n8615 & n25591;
  assign n25701 = pi629 & ~n25700;
  assign n25702 = ~n25699 & n25701;
  assign n25703 = n8499 & n63774;
  assign n25704 = n8606 & n25591;
  assign n25705 = ~pi629 & ~n25704;
  assign n25706 = ~n25703 & n25705;
  assign n25707 = pi792 & ~n25706;
  assign n25708 = pi792 & ~n25702;
  assign n25709 = ~n25706 & n25708;
  assign n25710 = ~n25703 & ~n25704;
  assign n25711 = ~pi629 & ~n25710;
  assign n25712 = ~n25699 & ~n25700;
  assign n25713 = pi629 & ~n25712;
  assign n25714 = ~n25711 & ~n25713;
  assign n25715 = pi792 & ~n25714;
  assign n25716 = ~n25702 & n25707;
  assign n25717 = ~n8651 & ~n63779;
  assign n25718 = ~n25698 & n25717;
  assign n25719 = ~n25604 & ~n25718;
  assign n25720 = pi644 & n25719;
  assign n25721 = ~pi787 & ~n25592;
  assign n25722 = pi1157 & ~n25595;
  assign n25723 = ~n25600 & ~n25722;
  assign n25724 = pi787 & ~n25723;
  assign n25725 = ~n25721 & ~n25724;
  assign n25726 = ~pi644 & n25725;
  assign n25727 = pi715 & ~n25726;
  assign n25728 = ~n25720 & n25727;
  assign n25729 = ~n8685 & n25521;
  assign n25730 = ~n8376 & n25571;
  assign n25731 = ~n8376 & ~n25574;
  assign n25732 = n8376 & n25521;
  assign n25733 = ~n25731 & ~n25732;
  assign n25734 = ~n25729 & ~n25730;
  assign n25735 = pi644 & ~n63780;
  assign n25736 = ~pi644 & n25521;
  assign n25737 = ~pi715 & ~n25736;
  assign n25738 = ~n25735 & n25737;
  assign n25739 = pi1160 & ~n25738;
  assign n25740 = ~n25728 & n25739;
  assign n25741 = ~pi644 & n25719;
  assign n25742 = pi644 & n25725;
  assign n25743 = ~pi715 & ~n25742;
  assign n25744 = ~n25741 & n25743;
  assign n25745 = ~pi644 & ~n63780;
  assign n25746 = pi644 & n25521;
  assign n25747 = pi715 & ~n25746;
  assign n25748 = ~n25745 & n25747;
  assign n25749 = ~pi1160 & ~n25748;
  assign n25750 = ~n25744 & n25749;
  assign n25751 = ~n25740 & ~n25750;
  assign n25752 = pi790 & ~n25751;
  assign n25753 = ~pi790 & n25719;
  assign n25754 = pi832 & ~n25753;
  assign n25755 = ~n25752 & n25754;
  assign po351 = ~n25520 & ~n25755;
  assign n25757 = pi199 & ~n62455;
  assign n25758 = pi199 & ~n8098;
  assign n25759 = n8257 & ~n25758;
  assign n25760 = n62880 & ~n25758;
  assign n25761 = ~pi637 & ~n25758;
  assign n25762 = ~pi199 & ~n7357;
  assign n25763 = n10997 & ~n25762;
  assign n25764 = pi199 & ~n62869;
  assign n25765 = ~pi199 & ~n8058;
  assign n25766 = pi39 & ~n25765;
  assign n25767 = ~n25764 & n25766;
  assign n25768 = ~pi199 & n7867;
  assign n25769 = pi199 & ~n7830;
  assign n25770 = ~pi39 & ~n25769;
  assign n25771 = ~pi39 & ~n25768;
  assign n25772 = ~n25769 & n25771;
  assign n25773 = ~n25768 & n25770;
  assign n25774 = ~pi38 & ~n63781;
  assign n25775 = ~n25767 & n25774;
  assign n25776 = ~n25763 & ~n25775;
  assign n25777 = n62765 & ~n25776;
  assign n25778 = pi199 & ~n62765;
  assign n25779 = pi637 & ~n25778;
  assign n25780 = ~n25777 & n25779;
  assign n25781 = ~n25761 & ~n25780;
  assign n25782 = ~pi778 & n25781;
  assign n25783 = pi625 & ~n25781;
  assign n25784 = ~pi625 & ~n25758;
  assign n25785 = pi1153 & ~n25784;
  assign n25786 = ~n25783 & n25785;
  assign n25787 = ~pi625 & ~n25781;
  assign n25788 = pi625 & ~n25758;
  assign n25789 = ~pi1153 & ~n25788;
  assign n25790 = ~n25787 & n25789;
  assign n25791 = ~n25786 & ~n25790;
  assign n25792 = pi778 & ~n25791;
  assign n25793 = ~n25782 & ~n25792;
  assign n25794 = ~n62880 & n25793;
  assign n25795 = ~n62880 & ~n25793;
  assign n25796 = n62880 & n25758;
  assign n25797 = ~n25795 & ~n25796;
  assign n25798 = ~n25760 & ~n25794;
  assign n25799 = ~n62882 & ~n63782;
  assign n25800 = n62882 & n25758;
  assign n25801 = n62882 & ~n25758;
  assign n25802 = ~n62882 & n63782;
  assign n25803 = ~n25801 & ~n25802;
  assign n25804 = ~n25799 & ~n25800;
  assign n25805 = ~n8257 & ~n63783;
  assign n25806 = ~n8257 & n63783;
  assign n25807 = n8257 & n25758;
  assign n25808 = ~n25806 & ~n25807;
  assign n25809 = ~n25759 & ~n25805;
  assign n25810 = ~n8303 & ~n63784;
  assign n25811 = n8303 & n25758;
  assign n25812 = n8303 & ~n25758;
  assign n25813 = ~n8303 & n63784;
  assign n25814 = ~n25812 & ~n25813;
  assign n25815 = ~n25810 & ~n25811;
  assign n25816 = pi628 & ~n63785;
  assign n25817 = ~pi628 & ~n25758;
  assign n25818 = pi1156 & ~n25817;
  assign n25819 = pi628 & n63785;
  assign n25820 = ~pi628 & n25758;
  assign n25821 = ~n25819 & ~n25820;
  assign n25822 = pi1156 & ~n25821;
  assign n25823 = ~n25816 & n25818;
  assign n25824 = ~pi628 & ~n63785;
  assign n25825 = pi628 & ~n25758;
  assign n25826 = ~pi1156 & ~n25825;
  assign n25827 = ~n25824 & n25826;
  assign n25828 = ~n25824 & ~n25825;
  assign n25829 = ~pi1156 & ~n25828;
  assign n25830 = pi1156 & n25821;
  assign n25831 = ~n25829 & ~n25830;
  assign n25832 = ~n63786 & ~n25827;
  assign n25833 = pi792 & n63787;
  assign n25834 = ~pi792 & n63785;
  assign n25835 = pi792 & ~n63787;
  assign n25836 = ~pi792 & ~n63785;
  assign n25837 = ~n25835 & ~n25836;
  assign n25838 = ~n25833 & ~n25834;
  assign n25839 = pi647 & ~n63788;
  assign n25840 = ~pi647 & ~n25758;
  assign n25841 = pi1157 & ~n25840;
  assign n25842 = pi647 & n63788;
  assign n25843 = ~pi647 & n25758;
  assign n25844 = ~n25842 & ~n25843;
  assign n25845 = pi1157 & ~n25844;
  assign n25846 = ~n25839 & n25841;
  assign n25847 = ~pi647 & ~n63788;
  assign n25848 = pi647 & ~n25758;
  assign n25849 = ~pi1157 & ~n25848;
  assign n25850 = ~n25847 & n25849;
  assign n25851 = ~n63789 & ~n25850;
  assign n25852 = pi787 & ~n25851;
  assign n25853 = ~pi787 & n63788;
  assign n25854 = ~n63036 & ~n25853;
  assign n25855 = ~n25852 & n25854;
  assign n25856 = ~pi617 & ~n25758;
  assign n25857 = n62765 & n10343;
  assign n25858 = pi199 & ~n25857;
  assign n25859 = n62765 & ~n14285;
  assign n25860 = pi199 & ~n62977;
  assign n25861 = n25859 & ~n25860;
  assign n25862 = pi617 & ~n25861;
  assign n25863 = ~pi199 & ~n7359;
  assign n25864 = n10342 & ~n25863;
  assign n25865 = pi199 & n62802;
  assign n25866 = ~pi199 & ~n7351;
  assign n25867 = ~pi38 & ~n25866;
  assign n25868 = ~n25865 & n25867;
  assign n25869 = ~n25864 & ~n25868;
  assign n25870 = n62765 & ~n25869;
  assign n25871 = pi617 & ~n25778;
  assign n25872 = ~n25870 & n25871;
  assign n25873 = ~n25858 & n25862;
  assign n25874 = ~n25856 & ~n63790;
  assign n25875 = ~n8135 & n25874;
  assign n25876 = n8135 & n25758;
  assign n25877 = ~n8135 & ~n25874;
  assign n25878 = n8135 & ~n25758;
  assign n25879 = ~n25877 & ~n25878;
  assign n25880 = ~n25875 & ~n25876;
  assign n25881 = ~pi785 & n63791;
  assign n25882 = pi609 & ~n63791;
  assign n25883 = ~pi609 & ~n25758;
  assign n25884 = pi1155 & ~n25883;
  assign n25885 = ~n25882 & n25884;
  assign n25886 = ~pi609 & ~n63791;
  assign n25887 = pi609 & ~n25758;
  assign n25888 = ~pi1155 & ~n25887;
  assign n25889 = ~n25886 & n25888;
  assign n25890 = ~n25885 & ~n25889;
  assign n25891 = pi785 & ~n25890;
  assign n25892 = ~n25881 & ~n25891;
  assign n25893 = ~pi781 & ~n25892;
  assign n25894 = pi618 & n25892;
  assign n25895 = ~pi618 & ~n25758;
  assign n25896 = pi1154 & ~n25895;
  assign n25897 = ~n25894 & n25896;
  assign n25898 = ~pi618 & n25892;
  assign n25899 = pi618 & ~n25758;
  assign n25900 = ~pi1154 & ~n25899;
  assign n25901 = ~n25898 & n25900;
  assign n25902 = ~n25897 & ~n25901;
  assign n25903 = pi781 & ~n25902;
  assign n25904 = ~n25893 & ~n25903;
  assign n25905 = ~pi789 & ~n25904;
  assign n25906 = pi619 & n25904;
  assign n25907 = ~pi619 & ~n25758;
  assign n25908 = pi1159 & ~n25907;
  assign n25909 = ~n25906 & n25908;
  assign n25910 = ~pi619 & n25904;
  assign n25911 = pi619 & ~n25758;
  assign n25912 = ~pi1159 & ~n25911;
  assign n25913 = ~n25910 & n25912;
  assign n25914 = ~n25909 & ~n25913;
  assign n25915 = pi789 & ~n25914;
  assign n25916 = ~n25905 & ~n25915;
  assign n25917 = ~n8595 & ~n25916;
  assign n25918 = n8595 & n25758;
  assign n25919 = ~n25917 & ~n25918;
  assign n25920 = ~n8334 & ~n25919;
  assign n25921 = n8334 & n25758;
  assign n25922 = ~n25920 & ~n25921;
  assign n25923 = ~n8376 & ~n25922;
  assign n25924 = n8376 & n25758;
  assign n25925 = pi644 & ~n16177;
  assign n25926 = ~pi644 & ~n16172;
  assign n25927 = ~pi644 & ~pi1160;
  assign n25928 = ~pi644 & pi1160;
  assign n25929 = pi644 & ~pi1160;
  assign n25930 = ~n25928 & ~n25929;
  assign n25931 = ~n14029 & ~n25927;
  assign n25932 = ~n16172 & ~n16177;
  assign n25933 = n63792 & ~n25932;
  assign n25934 = ~n25925 & ~n25926;
  assign n25935 = ~n25924 & n63793;
  assign n25936 = ~n25923 & n25935;
  assign n25937 = ~n63792 & ~n25932;
  assign n25938 = ~n25758 & n25937;
  assign n25939 = ~n25936 & ~n25938;
  assign n25940 = ~n25855 & n25939;
  assign n25941 = pi790 & ~n25940;
  assign n25942 = n8373 & ~n25844;
  assign n25943 = pi630 & n25850;
  assign n25944 = ~n8413 & ~n25922;
  assign n25945 = ~n25943 & ~n25944;
  assign n25946 = ~n25942 & n25945;
  assign n25947 = pi787 & ~n25946;
  assign n25948 = ~n63052 & ~n25919;
  assign n25949 = n8331 & ~n25821;
  assign n25950 = n8332 & n25828;
  assign n25951 = pi629 & n25827;
  assign n25952 = ~n25949 & ~n63794;
  assign n25953 = ~n25948 & n25952;
  assign n25954 = pi792 & ~n25953;
  assign n25955 = pi619 & ~n63783;
  assign n25956 = ~pi1159 & ~n25955;
  assign n25957 = ~pi648 & ~n25956;
  assign n25958 = ~pi648 & ~n25909;
  assign n25959 = ~n25956 & n25958;
  assign n25960 = ~n25909 & n25957;
  assign n25961 = ~pi619 & ~n63783;
  assign n25962 = pi1159 & ~n25961;
  assign n25963 = pi648 & ~n25913;
  assign n25964 = ~n25962 & n25963;
  assign n25965 = ~n63795 & ~n25964;
  assign n25966 = pi789 & ~n25965;
  assign n25967 = ~pi637 & n25874;
  assign n25968 = pi199 & n10352;
  assign n25969 = n62765 & ~n14472;
  assign n25970 = ~pi199 & ~n25969;
  assign n25971 = ~pi617 & ~n10351;
  assign n25972 = ~n25970 & n25971;
  assign n25973 = ~n25968 & n25971;
  assign n25974 = ~n25970 & n25973;
  assign n25975 = ~n25968 & n25972;
  assign n25976 = n62765 & ~n10362;
  assign n25977 = n2764 & n7868;
  assign n25978 = n25976 & ~n25977;
  assign n25979 = ~n10361 & n25976;
  assign n25980 = n62765 & n10363;
  assign n25981 = ~n8772 & n25978;
  assign n25982 = ~pi199 & ~n63797;
  assign n25983 = pi199 & n62980;
  assign n25984 = pi617 & ~n25983;
  assign n25985 = ~n25982 & n25984;
  assign n25986 = ~n25778 & ~n25985;
  assign n25987 = ~n63796 & n25986;
  assign n25988 = pi637 & ~n25987;
  assign n25989 = ~n25967 & ~n25988;
  assign n25990 = ~pi625 & n25989;
  assign n25991 = pi625 & ~n25874;
  assign n25992 = ~pi1153 & ~n25991;
  assign n25993 = ~n25990 & n25992;
  assign n25994 = ~pi608 & ~n25786;
  assign n25995 = ~n25993 & n25994;
  assign n25996 = pi625 & n25989;
  assign n25997 = ~pi625 & ~n25874;
  assign n25998 = pi1153 & ~n25997;
  assign n25999 = ~n25996 & n25998;
  assign n26000 = pi608 & ~n25790;
  assign n26001 = ~n25999 & n26000;
  assign n26002 = ~n25995 & ~n26001;
  assign n26003 = pi778 & ~n26002;
  assign n26004 = ~pi778 & n25989;
  assign n26005 = ~n26003 & ~n26004;
  assign n26006 = ~pi609 & ~n26005;
  assign n26007 = pi609 & n25793;
  assign n26008 = ~pi1155 & ~n26007;
  assign n26009 = ~n26006 & n26008;
  assign n26010 = ~pi660 & ~n25885;
  assign n26011 = ~n26009 & n26010;
  assign n26012 = pi609 & ~n26005;
  assign n26013 = ~pi609 & n25793;
  assign n26014 = pi1155 & ~n26013;
  assign n26015 = ~n26012 & n26014;
  assign n26016 = pi660 & ~n25889;
  assign n26017 = ~n26015 & n26016;
  assign n26018 = ~n26011 & ~n26017;
  assign n26019 = pi785 & ~n26018;
  assign n26020 = ~pi785 & ~n26005;
  assign n26021 = ~n26019 & ~n26020;
  assign n26022 = ~pi618 & ~n26021;
  assign n26023 = pi618 & n63782;
  assign n26024 = ~pi1154 & ~n26023;
  assign n26025 = ~n26022 & n26024;
  assign n26026 = ~pi627 & ~n25897;
  assign n26027 = ~n26025 & n26026;
  assign n26028 = pi618 & ~n26021;
  assign n26029 = ~pi618 & n63782;
  assign n26030 = pi1154 & ~n26029;
  assign n26031 = ~n26028 & n26030;
  assign n26032 = pi627 & ~n25901;
  assign n26033 = ~n26031 & n26032;
  assign n26034 = pi781 & ~n26033;
  assign n26035 = pi781 & ~n26027;
  assign n26036 = ~n26033 & n26035;
  assign n26037 = ~n26027 & n26034;
  assign n26038 = ~pi781 & n26021;
  assign n26039 = pi619 & n25963;
  assign n26040 = ~pi619 & n25958;
  assign n26041 = n11420 & ~n25909;
  assign n26042 = pi789 & ~n63799;
  assign n26043 = pi789 & ~n26039;
  assign n26044 = ~n63799 & n26043;
  assign n26045 = ~n26039 & n26042;
  assign n26046 = ~n26038 & ~n63800;
  assign n26047 = ~n63798 & n26046;
  assign n26048 = ~n26027 & ~n26033;
  assign n26049 = pi781 & ~n26048;
  assign n26050 = ~pi781 & ~n26021;
  assign n26051 = ~n26049 & ~n26050;
  assign n26052 = ~pi619 & ~n26051;
  assign n26053 = n25956 & ~n26052;
  assign n26054 = n25958 & ~n26053;
  assign n26055 = pi619 & ~n26051;
  assign n26056 = n25962 & ~n26055;
  assign n26057 = n25963 & ~n26056;
  assign n26058 = ~n26054 & ~n26057;
  assign n26059 = pi789 & ~n26058;
  assign n26060 = ~pi789 & ~n26051;
  assign n26061 = ~n26059 & ~n26060;
  assign n26062 = ~n25966 & ~n26047;
  assign n26063 = n62894 & ~n63801;
  assign n26064 = n12979 & n25916;
  assign n26065 = ~pi641 & ~n63784;
  assign n26066 = pi641 & n25758;
  assign n26067 = n8417 & ~n26066;
  assign n26068 = ~n26065 & n26067;
  assign n26069 = pi641 & ~n63784;
  assign n26070 = ~pi641 & n25758;
  assign n26071 = n8416 & ~n26070;
  assign n26072 = ~n26069 & n26071;
  assign n26073 = ~n26068 & ~n26072;
  assign n26074 = ~n26064 & n26073;
  assign n26075 = pi788 & ~n26074;
  assign n26076 = ~n63030 & ~n26075;
  assign n26077 = ~n26063 & n26076;
  assign n26078 = ~pi788 & n63801;
  assign n26079 = ~pi626 & n63801;
  assign n26080 = pi626 & ~n63784;
  assign n26081 = ~pi641 & ~n26080;
  assign n26082 = ~n26079 & n26081;
  assign n26083 = ~pi626 & ~n25916;
  assign n26084 = pi626 & n25758;
  assign n26085 = pi641 & ~n26084;
  assign n26086 = ~n26083 & n26085;
  assign n26087 = ~pi1158 & ~n26086;
  assign n26088 = ~n26082 & n26087;
  assign n26089 = pi626 & n63801;
  assign n26090 = ~pi626 & ~n63784;
  assign n26091 = pi641 & ~n26090;
  assign n26092 = ~n26089 & n26091;
  assign n26093 = pi626 & ~n25916;
  assign n26094 = ~pi626 & n25758;
  assign n26095 = ~pi641 & ~n26094;
  assign n26096 = ~n26093 & n26095;
  assign n26097 = pi1158 & ~n26096;
  assign n26098 = ~n26092 & n26097;
  assign n26099 = ~n26088 & ~n26098;
  assign n26100 = pi788 & ~n26099;
  assign n26101 = ~n26078 & ~n26100;
  assign n26102 = ~n26063 & ~n26075;
  assign n26103 = ~pi628 & n63802;
  assign n26104 = pi628 & n25919;
  assign n26105 = ~pi1156 & ~n26104;
  assign n26106 = ~n26103 & n26105;
  assign n26107 = ~pi629 & ~n63786;
  assign n26108 = ~n26106 & n26107;
  assign n26109 = pi628 & n63802;
  assign n26110 = ~pi628 & n25919;
  assign n26111 = pi1156 & ~n26110;
  assign n26112 = ~n26109 & n26111;
  assign n26113 = pi629 & ~n25827;
  assign n26114 = ~n26112 & n26113;
  assign n26115 = ~n26108 & ~n26114;
  assign n26116 = pi792 & ~n26115;
  assign n26117 = ~pi792 & n63802;
  assign n26118 = ~n26116 & ~n26117;
  assign n26119 = ~n25954 & ~n26077;
  assign n26120 = ~n25954 & n63802;
  assign n26121 = n63030 & n25953;
  assign n26122 = ~n8651 & ~n26121;
  assign n26123 = ~n26120 & n26122;
  assign n26124 = ~n8651 & n63803;
  assign n26125 = ~n11547 & ~n63804;
  assign n26126 = ~n25947 & n26125;
  assign n26127 = n62455 & ~n26126;
  assign n26128 = ~pi647 & ~n63803;
  assign n26129 = pi647 & n25922;
  assign n26130 = ~pi1157 & ~n26129;
  assign n26131 = ~n26128 & n26130;
  assign n26132 = ~pi630 & ~n63789;
  assign n26133 = ~n26131 & n26132;
  assign n26134 = pi647 & ~n63803;
  assign n26135 = ~pi647 & n25922;
  assign n26136 = pi1157 & ~n26135;
  assign n26137 = ~n26134 & n26136;
  assign n26138 = pi630 & ~n25850;
  assign n26139 = ~n26137 & n26138;
  assign n26140 = ~n26133 & ~n26139;
  assign n26141 = pi787 & ~n26140;
  assign n26142 = ~pi787 & ~n63803;
  assign n26143 = ~n26141 & ~n26142;
  assign n26144 = ~n25947 & ~n63804;
  assign n26145 = ~pi790 & n63805;
  assign n26146 = pi644 & ~n63805;
  assign n26147 = ~n25852 & ~n25853;
  assign n26148 = ~pi644 & n26147;
  assign n26149 = pi715 & ~n26148;
  assign n26150 = ~n26146 & n26149;
  assign n26151 = n8376 & ~n25758;
  assign n26152 = ~n8376 & n25922;
  assign n26153 = ~n25923 & ~n25924;
  assign n26154 = ~n26151 & ~n26152;
  assign n26155 = pi644 & n63806;
  assign n26156 = ~pi644 & ~n25758;
  assign n26157 = ~pi715 & ~n26156;
  assign n26158 = ~n26155 & n26157;
  assign n26159 = pi1160 & ~n26158;
  assign n26160 = ~n26150 & n26159;
  assign n26161 = ~pi644 & ~n63805;
  assign n26162 = pi644 & n26147;
  assign n26163 = ~pi715 & ~n26162;
  assign n26164 = ~n26161 & n26163;
  assign n26165 = ~pi644 & n63806;
  assign n26166 = pi644 & ~n25758;
  assign n26167 = pi715 & ~n26166;
  assign n26168 = ~n26165 & n26167;
  assign n26169 = ~pi1160 & ~n26168;
  assign n26170 = ~n26164 & n26169;
  assign n26171 = pi790 & ~n26170;
  assign n26172 = pi790 & ~n26160;
  assign n26173 = ~n26170 & n26172;
  assign n26174 = ~n26160 & n26171;
  assign n26175 = ~n26160 & ~n26170;
  assign n26176 = pi790 & ~n26175;
  assign n26177 = ~pi790 & ~n63805;
  assign n26178 = ~n26176 & ~n26177;
  assign n26179 = ~n26145 & ~n63807;
  assign n26180 = n62455 & n63808;
  assign n26181 = ~n25941 & n26127;
  assign n26182 = n62455 & ~n63808;
  assign n26183 = ~pi199 & ~n62455;
  assign n26184 = ~n26182 & ~n26183;
  assign n26185 = ~n25757 & ~n63809;
  assign n26186 = pi200 & ~n62455;
  assign n26187 = pi200 & ~n8098;
  assign n26188 = n8257 & ~n26187;
  assign n26189 = n62880 & ~n26187;
  assign n26190 = ~pi643 & ~n26187;
  assign n26191 = ~pi200 & ~n7357;
  assign n26192 = n10997 & ~n26191;
  assign n26193 = pi200 & ~n62868;
  assign n26194 = ~pi200 & n8034;
  assign n26195 = ~pi299 & ~n26194;
  assign n26196 = ~n26193 & n26195;
  assign n26197 = pi200 & ~n62865;
  assign n26198 = ~pi200 & n8056;
  assign n26199 = pi299 & ~n26198;
  assign n26200 = ~n26197 & n26199;
  assign n26201 = ~n26196 & ~n26200;
  assign n26202 = pi39 & ~n26201;
  assign n26203 = ~pi200 & ~n7867;
  assign n26204 = pi200 & n7830;
  assign n26205 = ~pi39 & ~n26204;
  assign n26206 = ~pi39 & ~n26203;
  assign n26207 = ~n26204 & n26206;
  assign n26208 = ~n26203 & n26205;
  assign n26209 = ~n26202 & ~n63811;
  assign n26210 = ~pi38 & ~n26209;
  assign n26211 = ~n26192 & ~n26210;
  assign n26212 = n62765 & ~n26211;
  assign n26213 = pi200 & ~n62765;
  assign n26214 = pi643 & ~n26213;
  assign n26215 = ~n26212 & n26214;
  assign n26216 = ~n26212 & ~n26213;
  assign n26217 = pi643 & ~n26216;
  assign n26218 = ~pi643 & n26187;
  assign n26219 = ~n26217 & ~n26218;
  assign n26220 = ~n26190 & ~n26215;
  assign n26221 = ~pi778 & ~n63812;
  assign n26222 = pi625 & n63812;
  assign n26223 = ~pi625 & ~n26187;
  assign n26224 = pi1153 & ~n26223;
  assign n26225 = ~n26222 & n26224;
  assign n26226 = ~pi625 & n63812;
  assign n26227 = pi625 & ~n26187;
  assign n26228 = ~pi1153 & ~n26227;
  assign n26229 = ~n26226 & n26228;
  assign n26230 = ~n26225 & ~n26229;
  assign n26231 = pi778 & ~n26230;
  assign n26232 = ~n26221 & ~n26231;
  assign n26233 = ~n62880 & n26232;
  assign n26234 = ~n62880 & ~n26232;
  assign n26235 = n62880 & n26187;
  assign n26236 = ~n26234 & ~n26235;
  assign n26237 = ~n26189 & ~n26233;
  assign n26238 = ~n62882 & ~n63813;
  assign n26239 = n62882 & n26187;
  assign n26240 = n62882 & ~n26187;
  assign n26241 = ~n62882 & n63813;
  assign n26242 = ~n26240 & ~n26241;
  assign n26243 = ~n26238 & ~n26239;
  assign n26244 = ~n8257 & ~n63814;
  assign n26245 = ~n8257 & n63814;
  assign n26246 = n8257 & n26187;
  assign n26247 = ~n26245 & ~n26246;
  assign n26248 = ~n26188 & ~n26244;
  assign n26249 = ~n8303 & ~n63815;
  assign n26250 = n8303 & n26187;
  assign n26251 = ~n26249 & ~n26250;
  assign n26252 = ~pi792 & ~n26251;
  assign n26253 = pi628 & n26251;
  assign n26254 = ~pi628 & ~n26187;
  assign n26255 = pi1156 & ~n26254;
  assign n26256 = ~n26253 & n26255;
  assign n26257 = ~pi628 & n26251;
  assign n26258 = pi628 & ~n26187;
  assign n26259 = ~pi1156 & ~n26258;
  assign n26260 = ~n26257 & n26259;
  assign n26261 = ~n26256 & ~n26260;
  assign n26262 = pi792 & ~n26261;
  assign n26263 = ~n26252 & ~n26262;
  assign n26264 = pi647 & ~n26263;
  assign n26265 = ~pi647 & n26187;
  assign n26266 = ~n26264 & ~n26265;
  assign n26267 = pi1157 & ~n26266;
  assign n26268 = ~pi647 & n26263;
  assign n26269 = pi647 & ~n26187;
  assign n26270 = ~pi1157 & ~n26269;
  assign n26271 = ~n26268 & n26270;
  assign n26272 = pi787 & ~n26271;
  assign n26273 = ~n26267 & n26272;
  assign n26274 = ~pi787 & n26263;
  assign n26275 = ~n63036 & ~n26274;
  assign n26276 = ~n26273 & n26275;
  assign n26277 = ~n11558 & n26187;
  assign n26278 = ~pi606 & ~n26187;
  assign n26279 = pi200 & ~n25857;
  assign n26280 = pi200 & ~n62977;
  assign n26281 = n25859 & ~n26280;
  assign n26282 = pi606 & ~n26281;
  assign n26283 = ~pi200 & ~n7359;
  assign n26284 = n10342 & ~n26283;
  assign n26285 = pi200 & n62802;
  assign n26286 = ~pi200 & ~n7351;
  assign n26287 = ~pi38 & ~n26286;
  assign n26288 = ~n26285 & n26287;
  assign n26289 = ~n26284 & ~n26288;
  assign n26290 = n62765 & ~n26289;
  assign n26291 = pi606 & ~n26213;
  assign n26292 = ~n26290 & n26291;
  assign n26293 = ~n26279 & n26282;
  assign n26294 = ~n26278 & ~n63816;
  assign n26295 = ~n8135 & n26294;
  assign n26296 = n8135 & n26187;
  assign n26297 = ~n8135 & ~n26294;
  assign n26298 = n8135 & ~n26187;
  assign n26299 = ~n26297 & ~n26298;
  assign n26300 = ~n26295 & ~n26296;
  assign n26301 = ~pi785 & n63817;
  assign n26302 = pi609 & ~n63817;
  assign n26303 = ~pi609 & ~n26187;
  assign n26304 = pi1155 & ~n26303;
  assign n26305 = ~n26302 & n26304;
  assign n26306 = ~pi609 & ~n63817;
  assign n26307 = pi609 & ~n26187;
  assign n26308 = ~pi1155 & ~n26307;
  assign n26309 = ~n26306 & n26308;
  assign n26310 = ~n26305 & ~n26309;
  assign n26311 = pi785 & ~n26310;
  assign n26312 = ~n26301 & ~n26311;
  assign n26313 = ~pi781 & ~n26312;
  assign n26314 = pi618 & n26312;
  assign n26315 = ~pi618 & ~n26187;
  assign n26316 = pi1154 & ~n26315;
  assign n26317 = ~n26314 & n26316;
  assign n26318 = ~pi618 & n26312;
  assign n26319 = pi618 & ~n26187;
  assign n26320 = ~pi1154 & ~n26319;
  assign n26321 = ~n26318 & n26320;
  assign n26322 = ~n26317 & ~n26321;
  assign n26323 = pi781 & ~n26322;
  assign n26324 = ~n26313 & ~n26323;
  assign n26325 = ~n11306 & n26324;
  assign n26326 = n11306 & ~n26187;
  assign n26327 = ~pi789 & ~n26324;
  assign n26328 = pi619 & n26324;
  assign n26329 = ~pi619 & ~n26187;
  assign n26330 = pi1159 & ~n26329;
  assign n26331 = ~n26328 & n26330;
  assign n26332 = ~pi619 & n26324;
  assign n26333 = pi619 & ~n26187;
  assign n26334 = ~pi1159 & ~n26333;
  assign n26335 = ~n26332 & n26334;
  assign n26336 = ~n26331 & ~n26335;
  assign n26337 = pi789 & ~n26336;
  assign n26338 = ~n26327 & ~n26337;
  assign n26339 = ~n26325 & ~n26326;
  assign n26340 = ~n8595 & ~n63818;
  assign n26341 = n8685 & n26340;
  assign n26342 = n8376 & ~n26187;
  assign n26343 = n8595 & n26187;
  assign n26344 = ~n26340 & ~n26343;
  assign n26345 = ~n8334 & ~n26344;
  assign n26346 = n8334 & n26187;
  assign n26347 = ~n26345 & ~n26346;
  assign n26348 = ~n8376 & n26347;
  assign n26349 = ~n26342 & ~n26348;
  assign n26350 = ~n8376 & ~n26347;
  assign n26351 = n8376 & n26187;
  assign n26352 = ~n26350 & ~n26351;
  assign n26353 = ~n26277 & ~n26341;
  assign n26354 = ~pi644 & ~n63819;
  assign n26355 = pi644 & ~n26187;
  assign n26356 = n16172 & ~n26355;
  assign n26357 = ~n26354 & n26356;
  assign n26358 = pi644 & ~n63819;
  assign n26359 = ~pi644 & ~n26187;
  assign n26360 = n16177 & ~n26359;
  assign n26361 = ~n26358 & n26360;
  assign n26362 = ~n26357 & ~n26361;
  assign n26363 = ~n26276 & n26362;
  assign n26364 = pi790 & ~n26363;
  assign n26365 = n8373 & ~n26266;
  assign n26366 = pi630 & n26271;
  assign n26367 = ~n8334 & n26344;
  assign n26368 = n8334 & ~n26187;
  assign n26369 = ~n8413 & ~n26368;
  assign n26370 = ~n8413 & ~n26347;
  assign n26371 = ~n26367 & n26369;
  assign n26372 = ~n26366 & ~n63820;
  assign n26373 = ~n26365 & ~n26366;
  assign n26374 = ~n63820 & n26373;
  assign n26375 = ~n26365 & n26372;
  assign n26376 = pi787 & ~n63821;
  assign n26377 = pi629 & n26260;
  assign n26378 = ~n63052 & ~n26344;
  assign n26379 = ~pi629 & n26256;
  assign n26380 = ~n26378 & ~n26379;
  assign n26381 = ~n26377 & ~n26379;
  assign n26382 = ~n26378 & n26381;
  assign n26383 = ~n26377 & n26380;
  assign n26384 = pi792 & ~n63822;
  assign n26385 = ~pi643 & n26294;
  assign n26386 = ~n7408 & ~n8085;
  assign n26387 = n26192 & ~n26386;
  assign n26388 = pi200 & ~n8759;
  assign n26389 = ~pi200 & ~n8763;
  assign n26390 = ~pi38 & ~n26389;
  assign n26391 = ~n26388 & n26390;
  assign n26392 = ~n26387 & ~n26391;
  assign n26393 = ~pi606 & n62765;
  assign n26394 = ~n26392 & n26393;
  assign n26395 = pi200 & ~n8779;
  assign n26396 = ~pi200 & ~n62901;
  assign n26397 = ~pi38 & ~n26396;
  assign n26398 = ~n26395 & n26397;
  assign n26399 = ~n8772 & ~n10362;
  assign n26400 = ~pi200 & ~n26399;
  assign n26401 = pi200 & n10335;
  assign n26402 = pi38 & pi200;
  assign n26403 = n10366 & n26402;
  assign n26404 = n7744 & n26401;
  assign n26405 = pi606 & n62765;
  assign n26406 = ~n63823 & n26405;
  assign n26407 = ~n26400 & n26406;
  assign n26408 = ~n26398 & n26406;
  assign n26409 = ~n26400 & n26408;
  assign n26410 = ~n26398 & n26407;
  assign n26411 = pi200 & n62980;
  assign n26412 = pi606 & ~n26411;
  assign n26413 = n62765 & ~n26412;
  assign n26414 = ~pi200 & ~n63797;
  assign n26415 = ~n26413 & ~n26414;
  assign n26416 = ~n26213 & ~n63824;
  assign n26417 = ~n26394 & ~n63825;
  assign n26418 = pi643 & ~n26417;
  assign n26419 = ~n26385 & ~n26418;
  assign n26420 = ~pi625 & n26419;
  assign n26421 = pi625 & ~n26294;
  assign n26422 = ~pi1153 & ~n26421;
  assign n26423 = ~n26420 & n26422;
  assign n26424 = ~pi608 & ~n26225;
  assign n26425 = ~pi608 & ~n26423;
  assign n26426 = ~n26225 & n26425;
  assign n26427 = ~n26423 & n26424;
  assign n26428 = pi625 & n26419;
  assign n26429 = ~pi625 & ~n26294;
  assign n26430 = pi1153 & ~n26429;
  assign n26431 = ~n26428 & n26430;
  assign n26432 = pi608 & ~n26229;
  assign n26433 = pi608 & ~n26431;
  assign n26434 = ~n26229 & n26433;
  assign n26435 = ~n26431 & n26432;
  assign n26436 = ~n63826 & ~n63827;
  assign n26437 = pi778 & ~n26436;
  assign n26438 = ~pi778 & n26419;
  assign n26439 = ~n26437 & ~n26438;
  assign n26440 = ~pi609 & ~n26439;
  assign n26441 = pi609 & n26232;
  assign n26442 = ~pi1155 & ~n26441;
  assign n26443 = ~n26440 & n26442;
  assign n26444 = ~pi660 & ~n26305;
  assign n26445 = ~n26443 & n26444;
  assign n26446 = pi609 & ~n26439;
  assign n26447 = ~pi609 & n26232;
  assign n26448 = pi1155 & ~n26447;
  assign n26449 = ~n26446 & n26448;
  assign n26450 = pi660 & ~n26309;
  assign n26451 = ~n26449 & n26450;
  assign n26452 = ~n26445 & ~n26451;
  assign n26453 = pi785 & ~n26452;
  assign n26454 = ~pi785 & ~n26439;
  assign n26455 = ~n26453 & ~n26454;
  assign n26456 = pi618 & ~n26455;
  assign n26457 = ~pi618 & n63813;
  assign n26458 = pi1154 & ~n26457;
  assign n26459 = ~n26456 & n26458;
  assign n26460 = pi627 & ~n26321;
  assign n26461 = ~n26459 & n26460;
  assign n26462 = ~pi618 & ~n26455;
  assign n26463 = pi618 & n63813;
  assign n26464 = ~pi1154 & ~n26463;
  assign n26465 = ~n26462 & n26464;
  assign n26466 = ~pi627 & ~n26317;
  assign n26467 = ~n26465 & n26466;
  assign n26468 = pi781 & ~n26467;
  assign n26469 = ~n26461 & n26468;
  assign n26470 = n8253 & ~n26329;
  assign n26471 = ~n26328 & n26470;
  assign n26472 = n8254 & ~n26333;
  assign n26473 = ~n26332 & n26472;
  assign n26474 = ~n11431 & n63814;
  assign n26475 = ~n26473 & ~n26474;
  assign n26476 = ~n26471 & n26475;
  assign n26477 = pi789 & ~n26476;
  assign n26478 = ~pi781 & n26455;
  assign n26479 = ~n26477 & ~n26478;
  assign n26480 = ~n26469 & n26479;
  assign n26481 = n11434 & n26476;
  assign n26482 = ~n26480 & ~n26481;
  assign n26483 = ~n26461 & ~n26467;
  assign n26484 = pi781 & ~n26483;
  assign n26485 = ~pi781 & ~n26455;
  assign n26486 = ~n26484 & ~n26485;
  assign n26487 = ~pi619 & ~n26486;
  assign n26488 = pi619 & ~n63814;
  assign n26489 = ~pi1159 & ~n26488;
  assign n26490 = ~n26487 & n26489;
  assign n26491 = ~pi648 & ~n26331;
  assign n26492 = ~n26490 & n26491;
  assign n26493 = pi619 & ~n26486;
  assign n26494 = ~pi619 & ~n63814;
  assign n26495 = pi1159 & ~n26494;
  assign n26496 = ~n26493 & n26495;
  assign n26497 = pi648 & ~n26335;
  assign n26498 = ~n26496 & n26497;
  assign n26499 = pi789 & ~n26498;
  assign n26500 = pi789 & ~n26492;
  assign n26501 = ~n26498 & n26500;
  assign n26502 = ~n26492 & n26499;
  assign n26503 = ~pi789 & n26486;
  assign n26504 = n62894 & ~n26503;
  assign n26505 = ~n63828 & n26504;
  assign n26506 = n62894 & ~n26482;
  assign n26507 = ~pi626 & ~n63818;
  assign n26508 = pi626 & n26187;
  assign n26509 = n8301 & ~n26508;
  assign n26510 = ~n26507 & n26509;
  assign n26511 = n8525 & n63815;
  assign n26512 = pi626 & ~n63818;
  assign n26513 = ~pi626 & n26187;
  assign n26514 = n8300 & ~n26513;
  assign n26515 = ~n26512 & n26514;
  assign n26516 = ~n26511 & ~n26515;
  assign n26517 = ~n26510 & ~n26511;
  assign n26518 = ~n26515 & n26517;
  assign n26519 = ~n26510 & n26516;
  assign n26520 = pi788 & ~n63830;
  assign n26521 = ~n63030 & ~n26520;
  assign n26522 = ~n63829 & n26521;
  assign n26523 = ~n26384 & ~n26522;
  assign n26524 = ~n8651 & ~n26523;
  assign n26525 = ~n26376 & ~n26524;
  assign n26526 = ~n11547 & ~n26525;
  assign n26527 = ~pi644 & n26525;
  assign n26528 = ~pi787 & ~n26263;
  assign n26529 = ~n26267 & ~n26271;
  assign n26530 = pi787 & ~n26529;
  assign n26531 = ~n26528 & ~n26530;
  assign n26532 = pi644 & n26531;
  assign n26533 = ~pi715 & ~n26532;
  assign n26534 = ~n26527 & n26533;
  assign n26535 = pi715 & ~n26355;
  assign n26536 = ~n26354 & n26535;
  assign n26537 = ~pi1160 & ~n26536;
  assign n26538 = ~n26534 & n26537;
  assign n26539 = pi644 & n26525;
  assign n26540 = ~pi644 & n26531;
  assign n26541 = pi715 & ~n26540;
  assign n26542 = ~n26539 & n26541;
  assign n26543 = ~pi715 & ~n26359;
  assign n26544 = ~n26358 & n26543;
  assign n26545 = pi1160 & ~n26544;
  assign n26546 = ~n26542 & n26545;
  assign n26547 = ~n26538 & ~n26546;
  assign n26548 = pi790 & ~n26547;
  assign n26549 = ~pi790 & n26525;
  assign n26550 = ~n26548 & ~n26549;
  assign n26551 = ~n26364 & ~n26526;
  assign n26552 = n62455 & n63831;
  assign n26553 = n62455 & ~n63831;
  assign n26554 = ~pi200 & ~n62455;
  assign n26555 = ~n26553 & ~n26554;
  assign n26556 = ~n26186 & ~n26552;
  assign n26557 = ~n8098 & n8257;
  assign n26558 = n62765 & n14370;
  assign n26559 = ~pi778 & ~n26558;
  assign n26560 = ~pi625 & ~n8098;
  assign n26561 = pi625 & ~n26558;
  assign n26562 = ~n26560 & ~n26561;
  assign n26563 = pi1153 & ~n26562;
  assign n26564 = ~pi625 & ~n26558;
  assign n26565 = ~n8099 & ~n26564;
  assign n26566 = ~pi1153 & ~n26565;
  assign n26567 = ~n26563 & ~n26566;
  assign n26568 = pi778 & ~n26567;
  assign n26569 = ~n26559 & ~n26568;
  assign n26570 = ~n62880 & ~n26569;
  assign n26571 = ~n8098 & n62880;
  assign n26572 = ~n62880 & n26569;
  assign n26573 = n8098 & n62880;
  assign n26574 = ~n26572 & ~n26573;
  assign n26575 = ~n26570 & ~n26571;
  assign n26576 = ~n62882 & ~n63833;
  assign n26577 = n8098 & n62882;
  assign n26578 = ~n8098 & n62882;
  assign n26579 = ~n62882 & n63833;
  assign n26580 = ~n26578 & ~n26579;
  assign n26581 = ~n26576 & ~n26577;
  assign n26582 = ~n8257 & ~n63834;
  assign n26583 = ~n8257 & n63834;
  assign n26584 = n8098 & n8257;
  assign n26585 = ~n26583 & ~n26584;
  assign n26586 = ~n26557 & ~n26582;
  assign n26587 = ~n8303 & ~n63835;
  assign n26588 = n8098 & n8303;
  assign n26589 = ~n8098 & n8303;
  assign n26590 = ~n8303 & n63835;
  assign n26591 = ~n26589 & ~n26590;
  assign n26592 = ~n26587 & ~n26588;
  assign n26593 = ~n62892 & n63836;
  assign n26594 = n8098 & n62892;
  assign n26595 = ~n62892 & ~n63836;
  assign n26596 = ~n8098 & n62892;
  assign n26597 = ~n26595 & ~n26596;
  assign n26598 = ~n26593 & ~n26594;
  assign n26599 = ~pi207 & n63837;
  assign n26600 = ~n62964 & n14367;
  assign n26601 = n10106 & n26600;
  assign n26602 = ~n8257 & n26601;
  assign n26603 = ~n8303 & n26602;
  assign n26604 = n10207 & n26600;
  assign n26605 = ~n62892 & n63838;
  assign n26606 = pi207 & ~n26605;
  assign n26607 = ~n26599 & ~n26606;
  assign n26608 = pi710 & ~n26607;
  assign n26609 = ~pi207 & ~n8098;
  assign n26610 = ~pi710 & ~n26609;
  assign n26611 = ~n26608 & ~n26610;
  assign n26612 = ~pi647 & n26611;
  assign n26613 = pi647 & n26609;
  assign n26614 = ~pi1157 & ~n26613;
  assign n26615 = ~n26612 & n26614;
  assign n26616 = pi630 & n26615;
  assign n26617 = pi647 & n26611;
  assign n26618 = ~pi647 & n26609;
  assign n26619 = pi1157 & ~n26618;
  assign n26620 = ~n26617 & n26619;
  assign n26621 = ~pi630 & n26620;
  assign n26622 = ~n8098 & n8135;
  assign n26623 = ~n8135 & ~n25857;
  assign n26624 = ~n26622 & ~n26623;
  assign n26625 = ~pi785 & ~n26624;
  assign n26626 = ~n8098 & ~n8148;
  assign n26627 = ~pi609 & n26623;
  assign n26628 = ~n26626 & ~n26627;
  assign n26629 = ~pi1155 & ~n26628;
  assign n26630 = ~n8098 & ~n8136;
  assign n26631 = pi609 & n26623;
  assign n26632 = ~n26630 & ~n26631;
  assign n26633 = pi1155 & ~n26632;
  assign n26634 = ~n26629 & ~n26633;
  assign n26635 = pi785 & ~n26634;
  assign n26636 = ~n26625 & ~n26635;
  assign n26637 = ~pi781 & ~n26636;
  assign n26638 = ~pi618 & n26636;
  assign n26639 = pi618 & n8098;
  assign n26640 = ~pi1154 & ~n26639;
  assign n26641 = ~n26638 & n26640;
  assign n26642 = pi618 & n26636;
  assign n26643 = ~pi618 & n8098;
  assign n26644 = pi1154 & ~n26643;
  assign n26645 = ~n26642 & n26644;
  assign n26646 = ~n26641 & ~n26645;
  assign n26647 = pi781 & ~n26646;
  assign n26648 = ~n26637 & ~n26647;
  assign n26649 = ~n11306 & n26648;
  assign n26650 = n8098 & n11306;
  assign n26651 = ~pi789 & ~n26648;
  assign n26652 = ~pi619 & n26648;
  assign n26653 = pi619 & n8098;
  assign n26654 = ~pi1159 & ~n26653;
  assign n26655 = ~n26652 & n26654;
  assign n26656 = pi619 & n26648;
  assign n26657 = ~pi619 & n8098;
  assign n26658 = pi1159 & ~n26657;
  assign n26659 = ~n26656 & n26658;
  assign n26660 = ~n26655 & ~n26659;
  assign n26661 = pi789 & ~n26660;
  assign n26662 = ~n26651 & ~n26661;
  assign n26663 = ~n26649 & ~n26650;
  assign n26664 = ~n8595 & n63839;
  assign n26665 = n8098 & n8595;
  assign n26666 = ~n26664 & ~n26665;
  assign n26667 = ~n8334 & ~n26666;
  assign n26668 = n8098 & n8334;
  assign n26669 = ~n26667 & ~n26668;
  assign n26670 = ~pi207 & ~n26669;
  assign n26671 = ~n8135 & n25859;
  assign n26672 = ~n63011 & n26671;
  assign n26673 = ~n63012 & n26672;
  assign n26674 = ~n11306 & n26673;
  assign n26675 = ~n8595 & n26674;
  assign n26676 = ~n8334 & n26675;
  assign n26677 = pi207 & ~n26676;
  assign n26678 = pi623 & ~n26677;
  assign n26679 = ~pi207 & n26669;
  assign n26680 = pi207 & n26676;
  assign n26681 = ~n26679 & ~n26680;
  assign n26682 = pi623 & ~n26681;
  assign n26683 = ~n26670 & n26678;
  assign n26684 = ~pi623 & n26609;
  assign n26685 = ~n63840 & ~n26684;
  assign n26686 = ~n8413 & n26685;
  assign n26687 = ~n26621 & ~n26686;
  assign n26688 = ~n26616 & ~n26621;
  assign n26689 = ~n26686 & n26688;
  assign n26690 = ~n26616 & n26687;
  assign n26691 = pi787 & ~n63841;
  assign n26692 = pi641 & ~n8098;
  assign n26693 = ~pi1158 & ~n26692;
  assign n26694 = pi618 & n63833;
  assign n26695 = pi609 & ~n26569;
  assign n26696 = n62765 & ~n10353;
  assign n26697 = ~pi778 & ~n26696;
  assign n26698 = ~pi608 & ~n26563;
  assign n26699 = ~pi625 & ~n26696;
  assign n26700 = ~n8099 & ~n26699;
  assign n26701 = ~pi1153 & ~n26700;
  assign n26702 = n26698 & ~n26701;
  assign n26703 = pi608 & ~n26566;
  assign n26704 = pi625 & ~n26696;
  assign n26705 = ~n26560 & ~n26704;
  assign n26706 = pi1153 & ~n26705;
  assign n26707 = n26703 & ~n26706;
  assign n26708 = pi778 & ~n26707;
  assign n26709 = pi778 & ~n26702;
  assign n26710 = ~n26707 & n26709;
  assign n26711 = ~n26702 & n26708;
  assign n26712 = ~n26697 & ~n63842;
  assign n26713 = ~pi609 & ~n26712;
  assign n26714 = ~n26695 & ~n26713;
  assign n26715 = ~pi1155 & ~n26714;
  assign n26716 = pi1155 & ~n8098;
  assign n26717 = ~pi660 & ~n26716;
  assign n26718 = ~n26715 & n26717;
  assign n26719 = ~pi609 & ~n26569;
  assign n26720 = pi609 & ~n26712;
  assign n26721 = ~n26719 & ~n26720;
  assign n26722 = pi1155 & ~n26721;
  assign n26723 = ~pi1155 & ~n8098;
  assign n26724 = pi660 & ~n26723;
  assign n26725 = ~n26722 & n26724;
  assign n26726 = ~n26718 & ~n26725;
  assign n26727 = pi785 & ~n26726;
  assign n26728 = ~pi785 & n26712;
  assign n26729 = ~n26727 & ~n26728;
  assign n26730 = ~pi618 & n26729;
  assign n26731 = ~n26694 & ~n26730;
  assign n26732 = ~pi1154 & ~n26731;
  assign n26733 = pi1154 & ~n8098;
  assign n26734 = ~pi627 & ~n26733;
  assign n26735 = ~n26732 & n26734;
  assign n26736 = ~pi618 & n63833;
  assign n26737 = pi618 & n26729;
  assign n26738 = ~n26736 & ~n26737;
  assign n26739 = pi1154 & ~n26738;
  assign n26740 = ~pi1154 & ~n8098;
  assign n26741 = pi627 & ~n26740;
  assign n26742 = ~n26739 & n26741;
  assign n26743 = ~n26735 & ~n26742;
  assign n26744 = pi781 & ~n26743;
  assign n26745 = ~pi781 & ~n26729;
  assign n26746 = ~n26744 & ~n26745;
  assign n26747 = ~pi619 & ~n26746;
  assign n26748 = pi619 & n63834;
  assign n26749 = ~pi1159 & ~n26748;
  assign n26750 = pi619 & ~n63834;
  assign n26751 = ~pi619 & n26746;
  assign n26752 = ~n26750 & ~n26751;
  assign n26753 = ~pi1159 & ~n26752;
  assign n26754 = ~n26747 & n26749;
  assign n26755 = pi1159 & ~n8098;
  assign n26756 = ~pi648 & ~n26755;
  assign n26757 = ~n63843 & n26756;
  assign n26758 = pi619 & ~n26746;
  assign n26759 = ~pi619 & n63834;
  assign n26760 = pi1159 & ~n26759;
  assign n26761 = ~pi619 & ~n63834;
  assign n26762 = pi619 & n26746;
  assign n26763 = ~n26761 & ~n26762;
  assign n26764 = pi1159 & ~n26763;
  assign n26765 = ~n26758 & n26760;
  assign n26766 = ~pi1159 & ~n8098;
  assign n26767 = pi648 & ~n26766;
  assign n26768 = ~n63844 & n26767;
  assign n26769 = ~n26757 & ~n26768;
  assign n26770 = pi789 & ~n26769;
  assign n26771 = ~pi789 & ~n26746;
  assign n26772 = ~n26770 & ~n26771;
  assign n26773 = ~pi626 & ~n26772;
  assign n26774 = pi626 & ~n63835;
  assign n26775 = ~pi641 & ~n26774;
  assign n26776 = ~n26773 & n26775;
  assign n26777 = n26693 & ~n26776;
  assign n26778 = ~pi641 & ~n8098;
  assign n26779 = pi1158 & ~n26778;
  assign n26780 = pi626 & ~n26772;
  assign n26781 = ~pi626 & ~n63835;
  assign n26782 = pi641 & ~n26781;
  assign n26783 = ~n26780 & n26782;
  assign n26784 = n26779 & ~n26783;
  assign n26785 = ~n26777 & ~n26784;
  assign n26786 = pi788 & ~n26785;
  assign n26787 = ~pi788 & ~n26772;
  assign n26788 = ~n63030 & ~n26787;
  assign n26789 = ~n26786 & n26788;
  assign n26790 = ~pi628 & ~n8098;
  assign n26791 = pi628 & ~n63836;
  assign n26792 = ~n26790 & ~n26791;
  assign n26793 = ~pi629 & ~n26792;
  assign n26794 = ~n26790 & ~n26793;
  assign n26795 = pi1156 & ~n26794;
  assign n26796 = ~pi628 & n63836;
  assign n26797 = pi628 & n8098;
  assign n26798 = n8332 & ~n26797;
  assign n26799 = pi628 & ~n8098;
  assign n26800 = ~pi628 & ~n63836;
  assign n26801 = ~n26799 & ~n26800;
  assign n26802 = n8332 & ~n26801;
  assign n26803 = ~n26796 & n26798;
  assign n26804 = ~pi1156 & n26799;
  assign n26805 = n8499 & ~n26797;
  assign n26806 = ~n63845 & ~n63846;
  assign n26807 = ~n26795 & n26806;
  assign n26808 = pi792 & ~n26807;
  assign n26809 = ~n26789 & ~n26808;
  assign n26810 = ~pi207 & ~n26809;
  assign n26811 = ~pi609 & ~n26600;
  assign n26812 = pi1155 & ~n26811;
  assign n26813 = pi660 & n26812;
  assign n26814 = n8164 & ~n26811;
  assign n26815 = ~pi609 & ~n63847;
  assign n26816 = pi609 & ~n26600;
  assign n26817 = ~pi1155 & ~n26816;
  assign n26818 = ~pi660 & n26817;
  assign n26819 = n8163 & ~n26816;
  assign n26820 = pi609 & ~n63848;
  assign n26821 = pi785 & ~n26820;
  assign n26822 = ~n26815 & n26821;
  assign n26823 = pi625 & n14367;
  assign n26824 = pi1153 & ~n26823;
  assign n26825 = ~pi608 & ~n26824;
  assign n26826 = ~pi625 & n25969;
  assign n26827 = ~pi1153 & ~n26826;
  assign n26828 = n26825 & ~n26827;
  assign n26829 = ~pi625 & n14367;
  assign n26830 = ~pi1153 & ~n26829;
  assign n26831 = pi608 & ~n26830;
  assign n26832 = pi625 & n25969;
  assign n26833 = pi1153 & ~n26832;
  assign n26834 = n26831 & ~n26833;
  assign n26835 = pi778 & ~n26834;
  assign n26836 = pi778 & ~n26828;
  assign n26837 = ~n26834 & n26836;
  assign n26838 = ~n26828 & n26835;
  assign n26839 = ~pi778 & ~n25969;
  assign n26840 = pi785 & ~n63848;
  assign n26841 = ~n63847 & n26840;
  assign n26842 = ~n26839 & ~n26841;
  assign n26843 = ~n63849 & n26842;
  assign n26844 = ~n63849 & ~n26839;
  assign n26845 = ~pi609 & ~n26844;
  assign n26846 = n63848 & ~n26845;
  assign n26847 = pi609 & ~n26844;
  assign n26848 = n63847 & ~n26847;
  assign n26849 = ~n26846 & ~n26848;
  assign n26850 = pi785 & ~n26849;
  assign n26851 = ~pi785 & n26844;
  assign n26852 = ~n26850 & ~n26851;
  assign n26853 = ~n26822 & ~n26843;
  assign n26854 = ~n11376 & ~n63850;
  assign n26855 = ~n62880 & n26600;
  assign n26856 = pi781 & ~n11383;
  assign n26857 = n26855 & n26856;
  assign n26858 = ~n26854 & ~n26857;
  assign n26859 = ~pi618 & n63850;
  assign n26860 = pi618 & ~n26855;
  assign n26861 = n8209 & ~n26860;
  assign n26862 = ~n26859 & n26861;
  assign n26863 = pi618 & n63850;
  assign n26864 = ~pi618 & ~n26855;
  assign n26865 = n8210 & ~n26864;
  assign n26866 = ~n26863 & n26865;
  assign n26867 = pi781 & ~n26866;
  assign n26868 = pi781 & ~n26862;
  assign n26869 = ~n26866 & n26868;
  assign n26870 = ~n26862 & n26867;
  assign n26871 = ~pi781 & n63850;
  assign n26872 = ~n11434 & ~n26871;
  assign n26873 = ~n63851 & n26872;
  assign n26874 = ~n11434 & ~n26858;
  assign n26875 = n62884 & n11306;
  assign n26876 = n26601 & n26875;
  assign n26877 = ~n63852 & ~n26876;
  assign n26878 = n62894 & ~n26877;
  assign n26879 = ~n8524 & n8595;
  assign n26880 = n26602 & n26879;
  assign n26881 = ~n26878 & ~n26880;
  assign n26882 = ~pi626 & n26877;
  assign n26883 = pi626 & ~n26602;
  assign n26884 = ~pi641 & ~n26883;
  assign n26885 = ~pi1158 & n26884;
  assign n26886 = ~n26882 & n26885;
  assign n26887 = pi626 & n26877;
  assign n26888 = ~pi626 & ~n26602;
  assign n26889 = pi641 & ~n26888;
  assign n26890 = pi1158 & n26889;
  assign n26891 = ~n26887 & n26890;
  assign n26892 = pi788 & ~n26891;
  assign n26893 = pi788 & ~n26886;
  assign n26894 = ~n26891 & n26893;
  assign n26895 = ~n26886 & n26892;
  assign n26896 = ~pi788 & n26877;
  assign n26897 = ~n63030 & ~n26896;
  assign n26898 = ~n63853 & n26897;
  assign n26899 = ~n63030 & ~n26881;
  assign n26900 = n8334 & n8500;
  assign n26901 = n63838 & n26900;
  assign n26902 = ~n63854 & ~n26901;
  assign n26903 = pi207 & ~n26902;
  assign n26904 = ~pi623 & ~n26903;
  assign n26905 = ~n26810 & n26904;
  assign n26906 = pi1156 & n26793;
  assign n26907 = ~n63052 & n26666;
  assign n26908 = ~n63845 & ~n26907;
  assign n26909 = ~n63845 & ~n26906;
  assign n26910 = ~n26907 & n26909;
  assign n26911 = ~n26906 & n26908;
  assign n26912 = pi792 & ~n63855;
  assign n26913 = n8253 & ~n26657;
  assign n26914 = ~n26656 & n26913;
  assign n26915 = n8254 & ~n26653;
  assign n26916 = ~n26652 & n26915;
  assign n26917 = ~n11431 & ~n63834;
  assign n26918 = ~n26916 & ~n26917;
  assign n26919 = ~n26914 & n26918;
  assign n26920 = n11434 & n26919;
  assign n26921 = n62765 & n62980;
  assign n26922 = ~pi778 & ~n26921;
  assign n26923 = pi625 & n26921;
  assign n26924 = ~pi625 & n25857;
  assign n26925 = pi1153 & ~n26924;
  assign n26926 = pi1153 & ~n26923;
  assign n26927 = ~n26924 & n26926;
  assign n26928 = ~n26923 & n26925;
  assign n26929 = n26703 & ~n63856;
  assign n26930 = ~pi625 & n26921;
  assign n26931 = pi625 & n25857;
  assign n26932 = ~pi1153 & ~n26931;
  assign n26933 = ~pi1153 & ~n26930;
  assign n26934 = ~n26931 & n26933;
  assign n26935 = ~n26930 & n26932;
  assign n26936 = n26698 & ~n63857;
  assign n26937 = pi778 & ~n26936;
  assign n26938 = pi778 & ~n26929;
  assign n26939 = ~n26936 & n26938;
  assign n26940 = ~n26929 & n26937;
  assign n26941 = ~n26922 & ~n63858;
  assign n26942 = ~pi609 & ~n26941;
  assign n26943 = ~n26695 & ~n26942;
  assign n26944 = ~pi1155 & ~n26943;
  assign n26945 = ~pi660 & ~n26633;
  assign n26946 = ~n26944 & n26945;
  assign n26947 = pi609 & ~n26941;
  assign n26948 = ~n26719 & ~n26947;
  assign n26949 = pi1155 & ~n26948;
  assign n26950 = pi660 & ~n26629;
  assign n26951 = ~n26949 & n26950;
  assign n26952 = ~n26946 & ~n26951;
  assign n26953 = pi785 & ~n26952;
  assign n26954 = ~pi785 & n26941;
  assign n26955 = ~n26953 & ~n26954;
  assign n26956 = ~pi618 & n26955;
  assign n26957 = ~n26694 & ~n26956;
  assign n26958 = ~pi1154 & ~n26957;
  assign n26959 = ~pi627 & ~n26645;
  assign n26960 = ~n26958 & n26959;
  assign n26961 = pi618 & n26955;
  assign n26962 = ~n26736 & ~n26961;
  assign n26963 = pi1154 & ~n26962;
  assign n26964 = pi627 & ~n26641;
  assign n26965 = ~n26963 & n26964;
  assign n26966 = pi781 & ~n26965;
  assign n26967 = ~n26960 & n26966;
  assign n26968 = ~pi781 & n26955;
  assign n26969 = pi789 & ~n26919;
  assign n26970 = ~n26968 & ~n26969;
  assign n26971 = ~n26960 & ~n26965;
  assign n26972 = pi781 & ~n26971;
  assign n26973 = ~pi781 & ~n26955;
  assign n26974 = ~n26972 & ~n26973;
  assign n26975 = ~n26967 & n26970;
  assign n26976 = ~n26920 & n63859;
  assign n26977 = ~pi619 & n63859;
  assign n26978 = ~n26750 & ~n26977;
  assign n26979 = ~pi1159 & ~n26978;
  assign n26980 = ~pi648 & ~n26659;
  assign n26981 = ~n26979 & n26980;
  assign n26982 = pi619 & n63859;
  assign n26983 = ~n26761 & ~n26982;
  assign n26984 = pi1159 & ~n26983;
  assign n26985 = pi648 & ~n26655;
  assign n26986 = ~n26984 & n26985;
  assign n26987 = pi789 & ~n26986;
  assign n26988 = pi789 & ~n26981;
  assign n26989 = ~n26986 & n26988;
  assign n26990 = ~n26981 & n26987;
  assign n26991 = ~pi789 & n63859;
  assign n26992 = n62894 & ~n26991;
  assign n26993 = ~n63860 & n26992;
  assign n26994 = n62894 & ~n26976;
  assign n26995 = ~pi641 & n63835;
  assign n26996 = pi626 & n26693;
  assign n26997 = n8417 & ~n26692;
  assign n26998 = ~n26995 & n63862;
  assign n26999 = n12979 & n63839;
  assign n27000 = pi641 & n63835;
  assign n27001 = ~pi626 & n26779;
  assign n27002 = n8416 & ~n26778;
  assign n27003 = ~n27000 & n63863;
  assign n27004 = ~n26999 & ~n27003;
  assign n27005 = ~n26998 & ~n27003;
  assign n27006 = ~n26999 & n27005;
  assign n27007 = ~n26998 & n27004;
  assign n27008 = pi788 & ~n63864;
  assign n27009 = ~n63030 & ~n27008;
  assign n27010 = ~n63861 & n27009;
  assign n27011 = ~n26912 & ~n27010;
  assign n27012 = ~pi207 & ~n27011;
  assign n27013 = ~pi778 & ~n63797;
  assign n27014 = ~pi625 & n63797;
  assign n27015 = pi625 & n25859;
  assign n27016 = ~pi1153 & ~n27015;
  assign n27017 = ~n27014 & n27016;
  assign n27018 = n26825 & ~n27017;
  assign n27019 = pi625 & n63797;
  assign n27020 = ~pi625 & n25859;
  assign n27021 = pi1153 & ~n27020;
  assign n27022 = ~n27019 & n27021;
  assign n27023 = n26831 & ~n27022;
  assign n27024 = pi778 & ~n27023;
  assign n27025 = pi778 & ~n27018;
  assign n27026 = ~n27023 & n27025;
  assign n27027 = ~n27018 & n27024;
  assign n27028 = ~n27013 & ~n63865;
  assign n27029 = ~pi785 & ~n27028;
  assign n27030 = ~pi609 & ~n27028;
  assign n27031 = n26817 & ~n27030;
  assign n27032 = n11295 & n26671;
  assign n27033 = ~pi660 & ~n27032;
  assign n27034 = ~n27031 & n27033;
  assign n27035 = pi609 & ~n27028;
  assign n27036 = n26812 & ~n27035;
  assign n27037 = n11296 & n26671;
  assign n27038 = pi660 & ~n27037;
  assign n27039 = ~n27036 & n27038;
  assign n27040 = ~n27034 & ~n27039;
  assign n27041 = pi785 & ~n27040;
  assign n27042 = ~n27029 & ~n27041;
  assign n27043 = pi618 & ~n27042;
  assign n27044 = pi1154 & ~n26864;
  assign n27045 = ~n27043 & n27044;
  assign n27046 = n11308 & n26672;
  assign n27047 = pi627 & ~n27046;
  assign n27048 = ~n27045 & n27047;
  assign n27049 = ~pi1154 & ~n26860;
  assign n27050 = n11307 & n26672;
  assign n27051 = ~pi627 & ~n27050;
  assign n27052 = ~n27049 & n27051;
  assign n27053 = ~n27048 & ~n27052;
  assign n27054 = pi781 & ~n27053;
  assign n27055 = ~pi618 & ~pi627;
  assign n27056 = pi781 & ~n27055;
  assign n27057 = ~n27042 & ~n27056;
  assign n27058 = ~pi1159 & ~n26673;
  assign n27059 = pi1159 & ~n26601;
  assign n27060 = n11428 & ~n27059;
  assign n27061 = n11428 & ~n27058;
  assign n27062 = ~n27059 & n27061;
  assign n27063 = ~n27058 & n27060;
  assign n27064 = pi1159 & ~n26673;
  assign n27065 = ~pi1159 & ~n26601;
  assign n27066 = n11425 & ~n27065;
  assign n27067 = n11425 & ~n27064;
  assign n27068 = ~n27065 & n27067;
  assign n27069 = ~n27064 & n27066;
  assign n27070 = pi789 & ~n63867;
  assign n27071 = pi789 & ~n63866;
  assign n27072 = ~n63867 & n27071;
  assign n27073 = ~n63866 & n27070;
  assign n27074 = ~n63021 & n63868;
  assign n27075 = ~n27057 & ~n27074;
  assign n27076 = n11425 & n26673;
  assign n27077 = n11428 & n26601;
  assign n27078 = pi1159 & ~n27077;
  assign n27079 = ~n27076 & n27078;
  assign n27080 = n11428 & n26673;
  assign n27081 = n11425 & n26601;
  assign n27082 = ~pi1159 & ~n27081;
  assign n27083 = ~n27080 & n27082;
  assign n27084 = pi789 & ~n27083;
  assign n27085 = ~n63866 & ~n63867;
  assign n27086 = pi789 & ~n27085;
  assign n27087 = pi789 & ~n63868;
  assign n27088 = ~n27079 & n27084;
  assign n27089 = ~n11434 & ~n27057;
  assign n27090 = ~n27054 & n27089;
  assign n27091 = ~n63869 & ~n27090;
  assign n27092 = ~n27054 & n27075;
  assign n27093 = n62894 & ~n63870;
  assign n27094 = n8523 & n26674;
  assign n27095 = n8522 & n26602;
  assign n27096 = pi1158 & ~n27095;
  assign n27097 = pi1158 & ~n27094;
  assign n27098 = ~n27095 & n27097;
  assign n27099 = ~n27094 & n27096;
  assign n27100 = n8522 & n26674;
  assign n27101 = n8523 & n26602;
  assign n27102 = ~pi1158 & ~n27101;
  assign n27103 = ~n27100 & n27102;
  assign n27104 = pi788 & ~n27103;
  assign n27105 = ~n63871 & n27104;
  assign n27106 = ~n27093 & ~n27105;
  assign n27107 = ~pi626 & n63870;
  assign n27108 = n26884 & ~n27107;
  assign n27109 = ~pi1158 & ~n27100;
  assign n27110 = ~n27108 & n27109;
  assign n27111 = pi626 & n63870;
  assign n27112 = n26889 & ~n27111;
  assign n27113 = n27097 & ~n27112;
  assign n27114 = ~n27110 & ~n27113;
  assign n27115 = pi788 & ~n27114;
  assign n27116 = ~pi788 & n63870;
  assign n27117 = ~n63030 & ~n27116;
  assign n27118 = ~n27115 & n27117;
  assign n27119 = ~n63030 & ~n27106;
  assign n27120 = n11801 & n26675;
  assign n27121 = n11799 & n63838;
  assign n27122 = pi1156 & ~n27121;
  assign n27123 = ~n27120 & n27122;
  assign n27124 = n11799 & n26675;
  assign n27125 = n11801 & n63838;
  assign n27126 = ~pi1156 & ~n27125;
  assign n27127 = ~pi1156 & ~n27124;
  assign n27128 = ~n27125 & n27127;
  assign n27129 = ~n27124 & n27126;
  assign n27130 = pi792 & ~n63873;
  assign n27131 = pi1156 & ~n26675;
  assign n27132 = ~pi1156 & ~n63838;
  assign n27133 = n11801 & ~n27132;
  assign n27134 = ~n27131 & n27133;
  assign n27135 = ~pi1156 & ~n26675;
  assign n27136 = pi1156 & ~n63838;
  assign n27137 = n11799 & ~n27136;
  assign n27138 = ~n27135 & n27137;
  assign n27139 = ~n27134 & ~n27138;
  assign n27140 = pi792 & ~n27139;
  assign n27141 = ~n27123 & n27130;
  assign n27142 = ~n63872 & ~n63874;
  assign n27143 = pi207 & ~n27142;
  assign n27144 = pi623 & ~n27143;
  assign n27145 = ~n27012 & n27144;
  assign n27146 = pi710 & ~n27145;
  assign n27147 = ~n26905 & n27146;
  assign n27148 = ~pi710 & ~n26685;
  assign n27149 = ~n8651 & ~n27148;
  assign n27150 = ~n27147 & n27149;
  assign n27151 = ~n26691 & ~n27150;
  assign n27152 = pi644 & n27151;
  assign n27153 = ~pi787 & ~n26611;
  assign n27154 = ~n26615 & ~n26620;
  assign n27155 = pi787 & ~n27154;
  assign n27156 = ~n27153 & ~n27155;
  assign n27157 = ~pi644 & n27156;
  assign n27158 = pi715 & ~n27157;
  assign n27159 = ~n27152 & n27158;
  assign n27160 = n8376 & ~n26609;
  assign n27161 = ~n8376 & n26685;
  assign n27162 = ~n8376 & ~n26685;
  assign n27163 = n8376 & n26609;
  assign n27164 = ~n27162 & ~n27163;
  assign n27165 = ~n27160 & ~n27161;
  assign n27166 = pi644 & ~n63875;
  assign n27167 = ~pi644 & n26609;
  assign n27168 = ~pi715 & ~n27167;
  assign n27169 = ~n27166 & n27168;
  assign n27170 = pi1160 & ~n27169;
  assign n27171 = ~n27159 & n27170;
  assign n27172 = ~pi644 & n27151;
  assign n27173 = pi644 & n27156;
  assign n27174 = ~pi715 & ~n27173;
  assign n27175 = ~n27172 & n27174;
  assign n27176 = ~pi644 & ~n63875;
  assign n27177 = pi644 & n26609;
  assign n27178 = pi715 & ~n27177;
  assign n27179 = ~n27176 & n27178;
  assign n27180 = ~pi1160 & ~n27179;
  assign n27181 = ~n27175 & n27180;
  assign n27182 = ~n27171 & ~n27181;
  assign n27183 = pi790 & ~n27182;
  assign n27184 = ~pi790 & n27151;
  assign n27185 = ~pi790 & ~n27151;
  assign n27186 = pi790 & ~n27181;
  assign n27187 = pi790 & ~n27171;
  assign n27188 = ~n27181 & n27187;
  assign n27189 = ~n27171 & n27186;
  assign n27190 = ~n27185 & ~n63876;
  assign n27191 = ~n27183 & ~n27184;
  assign n27192 = n62455 & n63877;
  assign n27193 = ~pi207 & ~n62455;
  assign n27194 = n62455 & ~n63877;
  assign n27195 = pi207 & ~n62455;
  assign n27196 = ~n27194 & ~n27195;
  assign n27197 = ~n27192 & ~n27193;
  assign n27198 = ~pi208 & n63837;
  assign n27199 = pi208 & ~n26605;
  assign n27200 = ~n27198 & ~n27199;
  assign n27201 = pi638 & ~n27200;
  assign n27202 = ~pi208 & ~n8098;
  assign n27203 = ~pi638 & ~n27202;
  assign n27204 = ~n27201 & ~n27203;
  assign n27205 = ~pi647 & n27204;
  assign n27206 = pi647 & n27202;
  assign n27207 = ~pi1157 & ~n27206;
  assign n27208 = ~n27205 & n27207;
  assign n27209 = pi630 & n27208;
  assign n27210 = pi647 & n27204;
  assign n27211 = ~pi647 & n27202;
  assign n27212 = pi1157 & ~n27211;
  assign n27213 = ~n27210 & n27212;
  assign n27214 = ~pi630 & n27213;
  assign n27215 = ~pi208 & ~n26669;
  assign n27216 = pi208 & ~n26676;
  assign n27217 = pi607 & ~n27216;
  assign n27218 = ~pi208 & n26669;
  assign n27219 = pi208 & n26676;
  assign n27220 = ~n27218 & ~n27219;
  assign n27221 = pi607 & ~n27220;
  assign n27222 = ~n27215 & n27217;
  assign n27223 = ~pi607 & n27202;
  assign n27224 = ~n63879 & ~n27223;
  assign n27225 = ~n8413 & n27224;
  assign n27226 = ~n27214 & ~n27225;
  assign n27227 = ~n27209 & ~n27214;
  assign n27228 = ~n27225 & n27227;
  assign n27229 = ~n27209 & n27226;
  assign n27230 = pi787 & ~n63880;
  assign n27231 = ~pi208 & ~n26809;
  assign n27232 = pi208 & ~n26902;
  assign n27233 = ~pi607 & ~n27232;
  assign n27234 = ~n27231 & n27233;
  assign n27235 = ~pi208 & ~n27011;
  assign n27236 = pi208 & ~n27142;
  assign n27237 = pi607 & ~n27236;
  assign n27238 = ~n27235 & n27237;
  assign n27239 = pi638 & ~n27238;
  assign n27240 = ~n27234 & n27239;
  assign n27241 = ~pi638 & ~n27224;
  assign n27242 = ~n8651 & ~n27241;
  assign n27243 = ~n27240 & n27242;
  assign n27244 = ~n27230 & ~n27243;
  assign n27245 = pi644 & n27244;
  assign n27246 = ~pi787 & ~n27204;
  assign n27247 = ~n27208 & ~n27213;
  assign n27248 = pi787 & ~n27247;
  assign n27249 = ~n27246 & ~n27248;
  assign n27250 = ~pi644 & n27249;
  assign n27251 = pi715 & ~n27250;
  assign n27252 = ~n27245 & n27251;
  assign n27253 = n8376 & ~n27202;
  assign n27254 = ~n8376 & n27224;
  assign n27255 = ~n8376 & ~n27224;
  assign n27256 = n8376 & n27202;
  assign n27257 = ~n27255 & ~n27256;
  assign n27258 = ~n27253 & ~n27254;
  assign n27259 = pi644 & ~n63881;
  assign n27260 = ~pi644 & n27202;
  assign n27261 = ~pi715 & ~n27260;
  assign n27262 = ~n27259 & n27261;
  assign n27263 = pi1160 & ~n27262;
  assign n27264 = ~n27252 & n27263;
  assign n27265 = ~pi644 & n27244;
  assign n27266 = pi644 & n27249;
  assign n27267 = ~pi715 & ~n27266;
  assign n27268 = ~n27265 & n27267;
  assign n27269 = ~pi644 & ~n63881;
  assign n27270 = pi644 & n27202;
  assign n27271 = pi715 & ~n27270;
  assign n27272 = ~n27269 & n27271;
  assign n27273 = ~pi1160 & ~n27272;
  assign n27274 = ~n27268 & n27273;
  assign n27275 = ~n27264 & ~n27274;
  assign n27276 = pi790 & ~n27275;
  assign n27277 = ~pi790 & n27244;
  assign n27278 = ~pi790 & ~n27244;
  assign n27279 = pi790 & ~n27274;
  assign n27280 = pi790 & ~n27264;
  assign n27281 = ~n27274 & n27280;
  assign n27282 = ~n27264 & n27279;
  assign n27283 = ~n27278 & ~n63882;
  assign n27284 = ~n27276 & ~n27277;
  assign n27285 = n62455 & n63883;
  assign n27286 = ~pi208 & ~n62455;
  assign n27287 = n62455 & ~n63883;
  assign n27288 = pi208 & ~n62455;
  assign n27289 = ~n27287 & ~n27288;
  assign n27290 = ~n27285 & ~n27286;
  assign n27291 = ~n8651 & ~n26809;
  assign n27292 = ~pi647 & ~n8098;
  assign n27293 = pi647 & ~n63837;
  assign n27294 = ~n27292 & ~n27293;
  assign n27295 = ~pi630 & ~n27294;
  assign n27296 = ~n27292 & ~n27295;
  assign n27297 = pi1157 & ~n27296;
  assign n27298 = pi647 & n8098;
  assign n27299 = pi647 & ~n8098;
  assign n27300 = ~pi1157 & n27299;
  assign n27301 = n8643 & ~n27298;
  assign n27302 = ~pi647 & n63837;
  assign n27303 = n8374 & ~n27298;
  assign n27304 = ~pi647 & ~n63837;
  assign n27305 = ~n27299 & ~n27304;
  assign n27306 = n8374 & ~n27305;
  assign n27307 = ~n27302 & n27303;
  assign n27308 = ~n63885 & ~n63886;
  assign n27309 = ~n27297 & n27308;
  assign n27310 = pi787 & ~n27309;
  assign n27311 = ~n27291 & ~n27310;
  assign n27312 = ~pi644 & ~n27311;
  assign n27313 = ~n8098 & n10298;
  assign n27314 = ~n10298 & ~n63837;
  assign n27315 = ~n10298 & n63837;
  assign n27316 = n8098 & n10298;
  assign n27317 = ~n27315 & ~n27316;
  assign n27318 = ~n27313 & ~n27314;
  assign n27319 = pi644 & n63887;
  assign n27320 = ~pi715 & ~n27319;
  assign n27321 = ~n27312 & n27320;
  assign n27322 = pi715 & n8098;
  assign n27323 = ~pi1160 & ~n27322;
  assign n27324 = ~n27321 & n27323;
  assign n27325 = pi644 & ~n27311;
  assign n27326 = ~pi644 & n63887;
  assign n27327 = pi715 & ~n27326;
  assign n27328 = ~n27325 & n27327;
  assign n27329 = ~pi715 & n8098;
  assign n27330 = pi1160 & ~n27329;
  assign n27331 = ~n27328 & n27330;
  assign n27332 = ~n27324 & ~n27331;
  assign n27333 = pi790 & ~n27332;
  assign n27334 = ~pi790 & ~n27311;
  assign n27335 = n62455 & ~n27334;
  assign n27336 = ~n27333 & n27335;
  assign n27337 = pi639 & n27336;
  assign n27338 = n3475 & n62765;
  assign n27339 = ~pi57 & n27338;
  assign n27340 = n62455 & n62765;
  assign n27341 = n62455 & n8098;
  assign n27342 = n8091 & n63888;
  assign n27343 = ~pi639 & n63889;
  assign n27344 = ~pi622 & ~n27343;
  assign n27345 = ~n27337 & n27344;
  assign n27346 = ~n8651 & ~n27011;
  assign n27347 = pi1157 & n27295;
  assign n27348 = ~n8413 & n26669;
  assign n27349 = ~n63886 & ~n27348;
  assign n27350 = ~n63886 & ~n27347;
  assign n27351 = ~n27348 & n27350;
  assign n27352 = ~n27347 & n27349;
  assign n27353 = pi787 & ~n63890;
  assign n27354 = ~n27346 & ~n27353;
  assign n27355 = ~pi644 & ~n27354;
  assign n27356 = n27320 & ~n27355;
  assign n27357 = ~n8098 & n8376;
  assign n27358 = ~n8376 & n26669;
  assign n27359 = ~n8376 & ~n26669;
  assign n27360 = n8098 & n8376;
  assign n27361 = ~n27359 & ~n27360;
  assign n27362 = ~n27357 & ~n27358;
  assign n27363 = ~pi644 & n63891;
  assign n27364 = pi644 & ~n8098;
  assign n27365 = ~pi644 & ~n63891;
  assign n27366 = pi644 & n8098;
  assign n27367 = ~n27365 & ~n27366;
  assign n27368 = ~n27363 & ~n27364;
  assign n27369 = pi715 & ~n63892;
  assign n27370 = ~pi1160 & ~n27369;
  assign n27371 = ~n27356 & n27370;
  assign n27372 = pi644 & ~n27354;
  assign n27373 = n27327 & ~n27372;
  assign n27374 = pi644 & n63891;
  assign n27375 = ~pi644 & ~n8098;
  assign n27376 = pi644 & ~n63891;
  assign n27377 = ~pi644 & n8098;
  assign n27378 = ~n27376 & ~n27377;
  assign n27379 = ~n27374 & ~n27375;
  assign n27380 = ~pi715 & ~n63893;
  assign n27381 = pi1160 & ~n27380;
  assign n27382 = ~n27373 & n27381;
  assign n27383 = ~n27371 & ~n27382;
  assign n27384 = pi790 & ~n27383;
  assign n27385 = ~pi790 & ~n27354;
  assign n27386 = n62455 & ~n27385;
  assign n27387 = ~n27384 & n27386;
  assign n27388 = pi639 & n27387;
  assign n27389 = ~pi1160 & ~n63892;
  assign n27390 = pi1160 & ~n63893;
  assign n27391 = pi790 & ~n27390;
  assign n27392 = pi790 & ~n27389;
  assign n27393 = ~n27390 & n27392;
  assign n27394 = ~n27389 & n27391;
  assign n27395 = ~pi790 & n63891;
  assign n27396 = n62455 & ~n27395;
  assign n27397 = ~n63894 & n27396;
  assign n27398 = ~pi639 & n27397;
  assign n27399 = pi622 & ~n27398;
  assign n27400 = ~n27388 & n27399;
  assign n27401 = ~n27345 & ~n27400;
  assign n27402 = ~pi209 & ~n27401;
  assign n27403 = n8685 & n26675;
  assign n27404 = n11558 & n26674;
  assign n27405 = pi1160 & ~n63895;
  assign n27406 = ~n10298 & n26605;
  assign n27407 = ~pi1160 & ~n27406;
  assign n27408 = n15025 & ~n27407;
  assign n27409 = ~n27405 & n27408;
  assign n27410 = ~pi1160 & ~n63895;
  assign n27411 = pi1160 & ~n27406;
  assign n27412 = n14949 & ~n27411;
  assign n27413 = ~n27410 & n27412;
  assign n27414 = ~n27409 & ~n27413;
  assign n27415 = pi790 & ~n27414;
  assign n27416 = ~n8651 & ~n27142;
  assign n27417 = n8409 & n26676;
  assign n27418 = n8411 & n26605;
  assign n27419 = pi1157 & ~n27418;
  assign n27420 = ~n27417 & n27419;
  assign n27421 = n8411 & n26676;
  assign n27422 = n8409 & n26605;
  assign n27423 = ~pi1157 & ~n27422;
  assign n27424 = ~n27421 & n27423;
  assign n27425 = pi787 & ~n27424;
  assign n27426 = ~pi1157 & ~n26605;
  assign n27427 = pi1157 & ~n26676;
  assign n27428 = n8409 & ~n27427;
  assign n27429 = ~n27426 & n27428;
  assign n27430 = pi1157 & ~n26605;
  assign n27431 = ~pi1157 & ~n26676;
  assign n27432 = n8411 & ~n27431;
  assign n27433 = ~n27430 & n27432;
  assign n27434 = ~n27429 & ~n27433;
  assign n27435 = pi787 & ~n27434;
  assign n27436 = ~n27420 & n27425;
  assign n27437 = ~pi647 & ~n27142;
  assign n27438 = pi647 & n26676;
  assign n27439 = ~pi1157 & ~n27438;
  assign n27440 = ~n27437 & n27439;
  assign n27441 = pi647 & n26605;
  assign n27442 = pi1157 & ~n27441;
  assign n27443 = ~pi630 & ~n27442;
  assign n27444 = ~n27440 & n27443;
  assign n27445 = pi647 & ~n27142;
  assign n27446 = ~pi647 & n26676;
  assign n27447 = pi1157 & ~n27446;
  assign n27448 = ~n27445 & n27447;
  assign n27449 = ~pi647 & n26605;
  assign n27450 = ~pi1157 & ~n27449;
  assign n27451 = pi630 & ~n27450;
  assign n27452 = ~n27448 & n27451;
  assign n27453 = ~n27444 & ~n27452;
  assign n27454 = pi787 & ~n27453;
  assign n27455 = ~pi787 & ~n27142;
  assign n27456 = ~n27454 & ~n27455;
  assign n27457 = ~n27416 & ~n63896;
  assign n27458 = ~n11547 & ~n63897;
  assign n27459 = ~n27415 & ~n27458;
  assign n27460 = pi644 & ~n27406;
  assign n27461 = ~pi715 & ~n27460;
  assign n27462 = ~pi644 & n63897;
  assign n27463 = n27461 & ~n27462;
  assign n27464 = pi715 & n13424;
  assign n27465 = n14949 & n63895;
  assign n27466 = n26674 & n27464;
  assign n27467 = ~pi1160 & ~n63898;
  assign n27468 = ~n27463 & n27467;
  assign n27469 = ~pi644 & ~n27406;
  assign n27470 = pi715 & ~n27469;
  assign n27471 = pi644 & n63897;
  assign n27472 = n27470 & ~n27471;
  assign n27473 = ~pi715 & n13413;
  assign n27474 = n15025 & n63895;
  assign n27475 = n26674 & n27473;
  assign n27476 = pi1160 & ~n63899;
  assign n27477 = ~n27472 & n27476;
  assign n27478 = ~n27468 & ~n27477;
  assign n27479 = pi790 & ~n27478;
  assign n27480 = ~pi790 & n63897;
  assign n27481 = n62455 & ~n27480;
  assign n27482 = ~n27479 & n27481;
  assign n27483 = n62455 & ~n27459;
  assign n27484 = pi622 & pi639;
  assign n27485 = ~n63900 & n27484;
  assign n27486 = ~n8651 & ~n26902;
  assign n27487 = n8376 & n8644;
  assign n27488 = n26605 & n27487;
  assign n27489 = ~n27486 & ~n27488;
  assign n27490 = ~n11547 & ~n27489;
  assign n27491 = pi790 & ~n63036;
  assign n27492 = n27406 & n27491;
  assign n27493 = ~n27490 & ~n27492;
  assign n27494 = pi644 & n27489;
  assign n27495 = pi1160 & n27470;
  assign n27496 = ~n27494 & n27495;
  assign n27497 = ~pi644 & n27489;
  assign n27498 = ~pi1160 & n27461;
  assign n27499 = ~n27497 & n27498;
  assign n27500 = pi790 & ~n27499;
  assign n27501 = pi790 & ~n27496;
  assign n27502 = ~n27499 & n27501;
  assign n27503 = ~n27496 & n27500;
  assign n27504 = ~pi790 & n27489;
  assign n27505 = n62455 & ~n27504;
  assign n27506 = ~n63901 & n27505;
  assign n27507 = n62455 & ~n27493;
  assign n27508 = ~pi622 & ~n63902;
  assign n27509 = pi790 & ~n63792;
  assign n27510 = n62455 & ~n27509;
  assign n27511 = n11558 & n27510;
  assign n27512 = n63895 & n27510;
  assign n27513 = n26674 & n27511;
  assign n27514 = pi622 & n63903;
  assign n27515 = ~pi639 & ~n27514;
  assign n27516 = pi209 & ~n27515;
  assign n27517 = pi639 & ~n27508;
  assign n27518 = ~n27514 & ~n27517;
  assign n27519 = pi209 & ~n27518;
  assign n27520 = ~n27508 & n27516;
  assign n27521 = ~n27485 & n63904;
  assign n27522 = ~n27402 & ~n27521;
  assign n27523 = ~pi695 & ~n27336;
  assign n27524 = pi695 & ~n63889;
  assign n27525 = ~pi217 & ~n27524;
  assign n27526 = ~n27523 & n27525;
  assign n27527 = ~pi695 & n63902;
  assign n27528 = pi217 & ~n27527;
  assign n27529 = ~pi612 & ~n27528;
  assign n27530 = ~n27526 & n27529;
  assign n27531 = ~pi695 & ~n27387;
  assign n27532 = pi695 & ~n27397;
  assign n27533 = ~pi217 & ~n27532;
  assign n27534 = ~n27531 & n27533;
  assign n27535 = ~pi695 & n63900;
  assign n27536 = pi695 & n63903;
  assign n27537 = pi217 & ~n27536;
  assign n27538 = ~n27535 & n27537;
  assign n27539 = pi612 & ~n27538;
  assign n27540 = ~n27534 & n27539;
  assign n27541 = ~n27530 & ~n27540;
  assign n27542 = pi198 & ~n62455;
  assign n27543 = n2764 & n62781;
  assign n27544 = n9733 & ~n27543;
  assign n27545 = pi198 & ~n27544;
  assign n27546 = pi198 & ~n62787;
  assign n27547 = ~n2971 & n27546;
  assign n27548 = pi198 & ~n6951;
  assign n27549 = n2908 & ~n27548;
  assign n27550 = pi198 & ~n7076;
  assign n27551 = ~n2908 & ~n27550;
  assign n27552 = ~n27549 & ~n27551;
  assign n27553 = n2971 & n27552;
  assign n27554 = ~n7034 & ~n27553;
  assign n27555 = ~n27547 & n27554;
  assign n27556 = n7034 & ~n27548;
  assign n27557 = ~pi223 & ~n27556;
  assign n27558 = ~n27555 & n27557;
  assign n27559 = pi198 & ~n6979;
  assign n27560 = ~n27549 & n27559;
  assign n27561 = ~n2904 & ~n6973;
  assign n27562 = n2904 & ~n6971;
  assign n27563 = pi198 & ~n27562;
  assign n27564 = pi198 & ~n62783;
  assign n27565 = ~n27561 & n27563;
  assign n27566 = ~n2971 & n63905;
  assign n27567 = ~n27560 & ~n27566;
  assign n27568 = pi223 & ~n27567;
  assign n27569 = ~pi299 & ~n27568;
  assign n27570 = ~n27558 & n27569;
  assign n27571 = ~n62393 & n27546;
  assign n27572 = n62393 & n27552;
  assign n27573 = ~n7118 & ~n27572;
  assign n27574 = ~n27571 & n27573;
  assign n27575 = n7118 & ~n27548;
  assign n27576 = ~pi215 & ~n27575;
  assign n27577 = ~n27574 & n27576;
  assign n27578 = ~n62393 & n63905;
  assign n27579 = ~n27560 & ~n27578;
  assign n27580 = pi215 & ~n27579;
  assign n27581 = pi299 & ~n27580;
  assign n27582 = ~n27577 & n27581;
  assign n27583 = ~pi38 & pi39;
  assign n27584 = pi39 & n62952;
  assign n27585 = n62765 & n27583;
  assign n27586 = ~n27582 & n63906;
  assign n27587 = ~n27570 & n63906;
  assign n27588 = ~n27582 & n27587;
  assign n27589 = ~n27570 & n27586;
  assign n27590 = ~n27545 & ~n63907;
  assign n27591 = n8595 & ~n27590;
  assign n27592 = pi198 & ~n62765;
  assign n27593 = pi633 & n6951;
  assign n27594 = ~n7176 & n27593;
  assign n27595 = ~n27548 & ~n27594;
  assign n27596 = pi603 & ~n27595;
  assign n27597 = ~pi603 & n27548;
  assign n27598 = ~n27596 & ~n27597;
  assign n27599 = ~n7186 & n27598;
  assign n27600 = n2814 & ~n27595;
  assign n27601 = ~n6971 & n27594;
  assign n27602 = ~n27559 & ~n27601;
  assign n27603 = ~n27600 & n27602;
  assign n27604 = pi603 & ~n27603;
  assign n27605 = n7186 & ~n27597;
  assign n27606 = ~n27604 & n27605;
  assign n27607 = ~n27599 & ~n27606;
  assign n27608 = ~n2907 & n27607;
  assign n27609 = ~n27559 & ~n27604;
  assign n27610 = n2907 & ~n27609;
  assign n27611 = ~n27608 & ~n27610;
  assign n27612 = n62393 & n27611;
  assign n27613 = pi633 & n7325;
  assign n27614 = ~n63905 & ~n27613;
  assign n27615 = ~n2907 & ~n27614;
  assign n27616 = pi198 & n6971;
  assign n27617 = ~n27601 & ~n27616;
  assign n27618 = n62796 & ~n27617;
  assign n27619 = ~n27615 & ~n27618;
  assign n27620 = ~n62393 & n27619;
  assign n27621 = pi215 & ~n27620;
  assign n27622 = ~n27612 & n27621;
  assign n27623 = pi198 & n7055;
  assign n27624 = pi633 & n7197;
  assign n27625 = ~n27623 & ~n27624;
  assign n27626 = ~n2814 & ~n27625;
  assign n27627 = ~n27600 & ~n27626;
  assign n27628 = pi603 & ~n27627;
  assign n27629 = ~pi642 & ~n27628;
  assign n27630 = pi642 & ~n27596;
  assign n27631 = n2903 & ~n27630;
  assign n27632 = ~n27629 & n27631;
  assign n27633 = ~n2903 & n27596;
  assign n27634 = ~n27597 & ~n27633;
  assign n27635 = ~n27632 & n27634;
  assign n27636 = ~n2907 & n27635;
  assign n27637 = ~pi603 & n27550;
  assign n27638 = n2907 & ~n27637;
  assign n27639 = ~n27628 & n27638;
  assign n27640 = ~n27636 & ~n27639;
  assign n27641 = n62393 & n27640;
  assign n27642 = n2814 & n27625;
  assign n27643 = ~n2814 & n27595;
  assign n27644 = pi603 & ~n7186;
  assign n27645 = ~n27643 & n27644;
  assign n27646 = ~n27642 & n27645;
  assign n27647 = pi603 & ~n27625;
  assign n27648 = n7186 & n27647;
  assign n27649 = pi198 & n7514;
  assign n27650 = ~n27648 & ~n27649;
  assign n27651 = ~n27646 & ~n27649;
  assign n27652 = ~n27648 & n27651;
  assign n27653 = ~n27646 & n27650;
  assign n27654 = ~n2907 & n63908;
  assign n27655 = n2907 & ~n27623;
  assign n27656 = ~n27647 & n27655;
  assign n27657 = ~n27654 & ~n27656;
  assign n27658 = ~n62393 & n27657;
  assign n27659 = ~n7118 & ~n27658;
  assign n27660 = ~n27641 & n27659;
  assign n27661 = n7118 & n27598;
  assign n27662 = ~pi215 & ~n27661;
  assign n27663 = ~n27660 & n27662;
  assign n27664 = ~n27622 & ~n27663;
  assign n27665 = pi299 & ~n27664;
  assign n27666 = n2971 & n27611;
  assign n27667 = ~n2971 & n27619;
  assign n27668 = pi223 & ~n27667;
  assign n27669 = ~n27666 & n27668;
  assign n27670 = n2971 & n27640;
  assign n27671 = ~n2971 & n27657;
  assign n27672 = ~n7034 & ~n27671;
  assign n27673 = ~n27670 & n27672;
  assign n27674 = n7034 & n27598;
  assign n27675 = ~pi223 & ~n27674;
  assign n27676 = ~n27673 & n27675;
  assign n27677 = ~n27669 & ~n27676;
  assign n27678 = ~pi299 & ~n27677;
  assign n27679 = pi39 & ~n27678;
  assign n27680 = pi39 & ~n27665;
  assign n27681 = ~n27678 & n27680;
  assign n27682 = ~n27665 & n27679;
  assign n27683 = pi198 & ~n6936;
  assign n27684 = pi603 & pi633;
  assign n27685 = ~n27683 & ~n27684;
  assign n27686 = pi198 & ~n7167;
  assign n27687 = ~pi198 & n7289;
  assign n27688 = ~pi198 & ~n7289;
  assign n27689 = pi198 & n7167;
  assign n27690 = ~n27688 & ~n27689;
  assign n27691 = ~n27686 & ~n27687;
  assign n27692 = n27684 & ~n63910;
  assign n27693 = ~n27685 & ~n27692;
  assign n27694 = pi299 & n27693;
  assign n27695 = ~n7153 & ~n7157;
  assign n27696 = pi633 & ~n27695;
  assign n27697 = ~n6939 & ~n27696;
  assign n27698 = ~n7162 & ~n27697;
  assign n27699 = ~pi299 & n27698;
  assign n27700 = ~pi39 & ~n27699;
  assign n27701 = ~n27694 & n27700;
  assign n27702 = ~n63909 & ~n27701;
  assign n27703 = ~pi38 & ~n27702;
  assign n27704 = pi39 & pi198;
  assign n27705 = pi38 & ~n27704;
  assign n27706 = pi198 & ~n6955;
  assign n27707 = pi633 & n7187;
  assign n27708 = n6955 & n27707;
  assign n27709 = ~n27706 & ~n27708;
  assign n27710 = ~pi39 & ~n27709;
  assign n27711 = n27705 & ~n27710;
  assign n27712 = n62765 & ~n27711;
  assign n27713 = ~n27703 & n27712;
  assign n27714 = ~n27592 & ~n27713;
  assign n27715 = ~n8135 & ~n27714;
  assign n27716 = n8135 & ~n27590;
  assign n27717 = ~n27715 & ~n27716;
  assign n27718 = ~pi785 & ~n27717;
  assign n27719 = ~n8136 & ~n27590;
  assign n27720 = pi609 & n27715;
  assign n27721 = ~n27719 & ~n27720;
  assign n27722 = pi1155 & ~n27721;
  assign n27723 = ~n8148 & ~n27590;
  assign n27724 = ~pi609 & n27715;
  assign n27725 = ~n27723 & ~n27724;
  assign n27726 = ~pi1155 & ~n27725;
  assign n27727 = ~n27722 & ~n27726;
  assign n27728 = pi785 & ~n27727;
  assign n27729 = ~n27718 & ~n27728;
  assign n27730 = ~pi781 & ~n27729;
  assign n27731 = pi618 & n27729;
  assign n27732 = ~pi618 & n27590;
  assign n27733 = pi1154 & ~n27732;
  assign n27734 = ~n27731 & n27733;
  assign n27735 = ~pi618 & n27729;
  assign n27736 = pi618 & n27590;
  assign n27737 = ~pi1154 & ~n27736;
  assign n27738 = ~n27735 & n27737;
  assign n27739 = ~n27734 & ~n27738;
  assign n27740 = pi781 & ~n27739;
  assign n27741 = ~n27730 & ~n27740;
  assign n27742 = ~n11306 & n27741;
  assign n27743 = n11306 & n27590;
  assign n27744 = ~pi789 & ~n27741;
  assign n27745 = pi619 & n27741;
  assign n27746 = ~pi619 & n27590;
  assign n27747 = pi1159 & ~n27746;
  assign n27748 = ~n27745 & n27747;
  assign n27749 = ~pi619 & n27741;
  assign n27750 = pi619 & n27590;
  assign n27751 = ~pi1159 & ~n27750;
  assign n27752 = ~n27749 & n27751;
  assign n27753 = ~n27748 & ~n27752;
  assign n27754 = pi789 & ~n27753;
  assign n27755 = ~n27744 & ~n27754;
  assign n27756 = ~n27742 & ~n27743;
  assign n27757 = ~n8595 & ~n63911;
  assign n27758 = ~n8595 & n63911;
  assign n27759 = n8595 & n27590;
  assign n27760 = ~n27758 & ~n27759;
  assign n27761 = ~n27591 & ~n27757;
  assign n27762 = ~n63052 & n63912;
  assign n27763 = ~n10206 & n27590;
  assign n27764 = n62882 & ~n27590;
  assign n27765 = ~n7544 & ~n27548;
  assign n27766 = pi634 & ~n27765;
  assign n27767 = ~n27548 & ~n27766;
  assign n27768 = ~n2904 & n27767;
  assign n27769 = n7365 & ~n27768;
  assign n27770 = n2814 & ~n27767;
  assign n27771 = pi634 & n62822;
  assign n27772 = ~n27623 & ~n27771;
  assign n27773 = ~n2814 & ~n27772;
  assign n27774 = ~n27770 & ~n27773;
  assign n27775 = n2904 & n27774;
  assign n27776 = n27769 & ~n27775;
  assign n27777 = n2907 & ~n27774;
  assign n27778 = n2904 & ~n27550;
  assign n27779 = ~n2904 & ~n27548;
  assign n27780 = ~pi680 & ~n27779;
  assign n27781 = ~n27778 & n27780;
  assign n27782 = ~n27777 & ~n27781;
  assign n27783 = ~n27776 & n27782;
  assign n27784 = n2971 & ~n27783;
  assign n27785 = ~n2814 & n27767;
  assign n27786 = n2814 & n27772;
  assign n27787 = ~n27785 & ~n27786;
  assign n27788 = ~n2904 & ~n27787;
  assign n27789 = n2904 & n27772;
  assign n27790 = n7365 & ~n27789;
  assign n27791 = ~n27788 & n27790;
  assign n27792 = pi198 & n7397;
  assign n27793 = n2907 & ~n27772;
  assign n27794 = ~n27792 & ~n27793;
  assign n27795 = ~n27791 & n27794;
  assign n27796 = ~n2971 & ~n27795;
  assign n27797 = ~n7034 & ~n27796;
  assign n27798 = ~n7034 & ~n27784;
  assign n27799 = ~n27796 & n27798;
  assign n27800 = ~n27784 & n27797;
  assign n27801 = pi634 & n6951;
  assign n27802 = n7563 & n27801;
  assign n27803 = pi634 & pi680;
  assign n27804 = pi680 & n27766;
  assign n27805 = ~n27765 & n27803;
  assign n27806 = ~n27548 & ~n63914;
  assign n27807 = n7034 & n27806;
  assign n27808 = n27556 & ~n27802;
  assign n27809 = ~pi223 & ~n63915;
  assign n27810 = ~n63913 & n27809;
  assign n27811 = pi634 & ~n6971;
  assign n27812 = n7544 & n27811;
  assign n27813 = ~n27616 & ~n27812;
  assign n27814 = ~n2814 & ~n27813;
  assign n27815 = ~n27770 & ~n27814;
  assign n27816 = n2904 & n27815;
  assign n27817 = n27769 & ~n27816;
  assign n27818 = ~pi680 & n63905;
  assign n27819 = n27559 & n27818;
  assign n27820 = ~n6979 & n27818;
  assign n27821 = n2907 & ~n27815;
  assign n27822 = ~n63916 & ~n27821;
  assign n27823 = ~n27817 & n27822;
  assign n27824 = n2971 & n27823;
  assign n27825 = n2814 & n27813;
  assign n27826 = ~n27785 & ~n27825;
  assign n27827 = ~n2904 & ~n27826;
  assign n27828 = n2904 & n27813;
  assign n27829 = n7365 & ~n27828;
  assign n27830 = ~n27827 & n27829;
  assign n27831 = n2907 & ~n27813;
  assign n27832 = ~n27818 & ~n27831;
  assign n27833 = ~n27830 & n27832;
  assign n27834 = ~n2971 & n27833;
  assign n27835 = pi223 & ~n27834;
  assign n27836 = pi223 & ~n27824;
  assign n27837 = ~n27834 & n27836;
  assign n27838 = ~n27824 & n27835;
  assign n27839 = ~pi299 & ~n63917;
  assign n27840 = ~n27810 & n27839;
  assign n27841 = ~n62393 & ~n27795;
  assign n27842 = n62393 & ~n27783;
  assign n27843 = ~n7118 & ~n27842;
  assign n27844 = ~n7118 & ~n27841;
  assign n27845 = ~n27842 & n27844;
  assign n27846 = ~n27841 & n27843;
  assign n27847 = n7118 & n27806;
  assign n27848 = n27575 & ~n27802;
  assign n27849 = ~pi215 & ~n63919;
  assign n27850 = ~n63918 & n27849;
  assign n27851 = n62393 & n27823;
  assign n27852 = ~n62393 & n27833;
  assign n27853 = pi215 & ~n27852;
  assign n27854 = pi215 & ~n27851;
  assign n27855 = ~n27852 & n27854;
  assign n27856 = ~n27851 & n27853;
  assign n27857 = pi299 & ~n63920;
  assign n27858 = ~n27850 & n27857;
  assign n27859 = ~n27840 & ~n27858;
  assign n27860 = ~n27850 & ~n63920;
  assign n27861 = pi299 & ~n27860;
  assign n27862 = ~n27810 & ~n63917;
  assign n27863 = ~pi299 & ~n27862;
  assign n27864 = pi39 & ~n27863;
  assign n27865 = ~n27861 & n27864;
  assign n27866 = pi39 & ~n27859;
  assign n27867 = ~pi198 & n7849;
  assign n27868 = pi198 & ~n7826;
  assign n27869 = ~n27867 & ~n27868;
  assign n27870 = n27803 & n27869;
  assign n27871 = ~n27683 & ~n27803;
  assign n27872 = pi299 & ~n27871;
  assign n27873 = n27803 & ~n27869;
  assign n27874 = n27683 & ~n27803;
  assign n27875 = ~n27873 & ~n27874;
  assign n27876 = pi299 & ~n27875;
  assign n27877 = ~n27870 & n27872;
  assign n27878 = pi198 & n7816;
  assign n27879 = ~n7836 & n27803;
  assign n27880 = ~n27878 & n27879;
  assign n27881 = ~n6939 & ~n27880;
  assign n27882 = ~pi299 & ~n27881;
  assign n27883 = ~pi39 & ~n27882;
  assign n27884 = ~n63922 & n27883;
  assign n27885 = ~n63921 & ~n27884;
  assign n27886 = ~pi38 & ~n27885;
  assign n27887 = pi634 & n7563;
  assign n27888 = n6955 & n27887;
  assign n27889 = ~n27706 & ~n27888;
  assign n27890 = ~pi39 & ~n27889;
  assign n27891 = n27705 & ~n27890;
  assign n27892 = n62765 & ~n27891;
  assign n27893 = ~n27886 & n27892;
  assign n27894 = ~n27592 & ~n27893;
  assign n27895 = ~pi778 & ~n27894;
  assign n27896 = pi625 & n27894;
  assign n27897 = ~pi625 & n27590;
  assign n27898 = pi1153 & ~n27897;
  assign n27899 = ~n27896 & n27898;
  assign n27900 = ~pi625 & n27894;
  assign n27901 = pi625 & n27590;
  assign n27902 = ~pi1153 & ~n27901;
  assign n27903 = ~n27900 & n27902;
  assign n27904 = ~n27899 & ~n27903;
  assign n27905 = pi778 & ~n27904;
  assign n27906 = ~n27895 & ~n27905;
  assign n27907 = ~n62880 & n27906;
  assign n27908 = n62880 & n27590;
  assign n27909 = ~n62880 & ~n27906;
  assign n27910 = n62880 & ~n27590;
  assign n27911 = ~n27909 & ~n27910;
  assign n27912 = ~n27907 & ~n27908;
  assign n27913 = ~n62882 & ~n63923;
  assign n27914 = ~n62882 & n63923;
  assign n27915 = n62882 & n27590;
  assign n27916 = ~n27914 & ~n27915;
  assign n27917 = ~n27764 & ~n27913;
  assign n27918 = ~n8257 & ~n63924;
  assign n27919 = ~n8303 & n27918;
  assign n27920 = ~n27763 & ~n27919;
  assign n27921 = pi628 & ~n27920;
  assign n27922 = ~pi628 & n27590;
  assign n27923 = pi1156 & ~n27922;
  assign n27924 = ~n27921 & ~n27922;
  assign n27925 = pi1156 & n27924;
  assign n27926 = ~n27921 & n27923;
  assign n27927 = n8331 & n27924;
  assign n27928 = ~pi629 & n63925;
  assign n27929 = ~pi628 & ~n27920;
  assign n27930 = pi628 & n27590;
  assign n27931 = ~pi1156 & ~n27930;
  assign n27932 = ~n27929 & n27931;
  assign n27933 = pi629 & n27932;
  assign n27934 = ~n63926 & ~n27933;
  assign n27935 = ~n27762 & n27934;
  assign n27936 = pi792 & ~n27935;
  assign n27937 = pi626 & ~n63911;
  assign n27938 = ~pi626 & ~n27590;
  assign n27939 = n8300 & ~n27938;
  assign n27940 = ~n27937 & n27939;
  assign n27941 = n8257 & n27590;
  assign n27942 = ~n27918 & ~n27941;
  assign n27943 = n8525 & ~n27942;
  assign n27944 = ~pi626 & ~n63911;
  assign n27945 = pi626 & ~n27590;
  assign n27946 = n8301 & ~n27945;
  assign n27947 = ~n27944 & n27946;
  assign n27948 = ~n27943 & ~n27947;
  assign n27949 = ~n27940 & ~n27943;
  assign n27950 = ~n27947 & n27949;
  assign n27951 = ~n27940 & n27948;
  assign n27952 = pi788 & ~n63927;
  assign n27953 = ~n7159 & n7817;
  assign n27954 = pi634 & ~n27953;
  assign n27955 = ~pi634 & ~n6939;
  assign n27956 = ~pi633 & ~n27955;
  assign n27957 = ~pi634 & n6939;
  assign n27958 = pi634 & n7817;
  assign n27959 = ~n7159 & n27958;
  assign n27960 = ~n27957 & ~n27959;
  assign n27961 = ~pi633 & ~n27960;
  assign n27962 = ~n27954 & n27956;
  assign n27963 = pi634 & ~pi665;
  assign n27964 = pi198 & ~pi633;
  assign n27965 = n27963 & ~n27964;
  assign n27966 = ~n7151 & n27965;
  assign n27967 = pi603 & ~n27966;
  assign n27968 = ~n27696 & n27967;
  assign n27969 = ~n63928 & n27968;
  assign n27970 = ~pi603 & n27881;
  assign n27971 = pi680 & ~n27970;
  assign n27972 = ~n27969 & n27971;
  assign n27973 = ~pi680 & n27698;
  assign n27974 = ~pi299 & ~n27973;
  assign n27975 = ~n27972 & n27974;
  assign n27976 = ~pi603 & ~n27869;
  assign n27977 = pi198 & ~pi665;
  assign n27978 = pi633 & ~n27977;
  assign n27979 = ~n27867 & n27978;
  assign n27980 = ~n63910 & n27979;
  assign n27981 = ~n7289 & n27868;
  assign n27982 = ~pi198 & ~pi665;
  assign n27983 = n7167 & n27982;
  assign n27984 = ~pi633 & ~n27983;
  assign n27985 = ~n27981 & n27984;
  assign n27986 = pi603 & ~n27985;
  assign n27987 = ~n27980 & n27986;
  assign n27988 = ~n27976 & ~n27987;
  assign n27989 = ~n27980 & ~n27985;
  assign n27990 = pi603 & ~n27989;
  assign n27991 = ~pi603 & n27869;
  assign n27992 = n27803 & ~n27991;
  assign n27993 = ~n27990 & n27992;
  assign n27994 = n27803 & ~n27988;
  assign n27995 = n27693 & ~n27803;
  assign n27996 = pi299 & ~n27995;
  assign n27997 = ~n63929 & n27996;
  assign n27998 = ~n27975 & ~n27997;
  assign n27999 = ~pi39 & ~n27998;
  assign n28000 = ~pi680 & n27635;
  assign n28001 = n7177 & n27963;
  assign n28002 = n27595 & ~n28001;
  assign n28003 = n2814 & ~n28002;
  assign n28004 = pi634 & n62824;
  assign n28005 = n27625 & ~n28004;
  assign n28006 = ~n2814 & ~n28005;
  assign n28007 = ~n28003 & ~n28006;
  assign n28008 = pi603 & ~n28007;
  assign n28009 = ~pi642 & n28008;
  assign n28010 = ~pi603 & ~n27767;
  assign n28011 = pi603 & ~n28002;
  assign n28012 = pi642 & n28011;
  assign n28013 = ~n28010 & ~n28012;
  assign n28014 = ~n28009 & n28013;
  assign n28015 = n2903 & ~n28014;
  assign n28016 = ~n28010 & ~n28011;
  assign n28017 = ~n2903 & ~n28016;
  assign n28018 = ~n7008 & ~n28017;
  assign n28019 = ~n28015 & n28018;
  assign n28020 = ~pi603 & ~n27774;
  assign n28021 = n7008 & ~n28020;
  assign n28022 = ~n28008 & n28021;
  assign n28023 = ~n28019 & ~n28022;
  assign n28024 = pi680 & ~n28023;
  assign n28025 = ~n28000 & ~n28024;
  assign n28026 = n62393 & n28025;
  assign n28027 = ~pi603 & n27787;
  assign n28028 = ~n7186 & n28011;
  assign n28029 = ~n27645 & ~n28028;
  assign n28030 = ~n2904 & n28029;
  assign n28031 = ~n2814 & ~n28029;
  assign n28032 = n28005 & ~n28031;
  assign n28033 = ~n28030 & ~n28032;
  assign n28034 = ~n28027 & ~n28033;
  assign n28035 = n7365 & ~n28034;
  assign n28036 = ~pi680 & ~n63908;
  assign n28037 = ~n7187 & ~n27772;
  assign n28038 = ~n27647 & ~n28037;
  assign n28039 = n2907 & ~n28038;
  assign n28040 = ~n28036 & ~n28039;
  assign n28041 = ~n28035 & ~n28039;
  assign n28042 = ~n28036 & n28041;
  assign n28043 = ~n28035 & n28040;
  assign n28044 = ~n62393 & ~n63930;
  assign n28045 = ~n7118 & ~n28044;
  assign n28046 = ~n28026 & n28045;
  assign n28047 = n7408 & n27766;
  assign n28048 = n27598 & ~n28047;
  assign n28049 = n7118 & n28048;
  assign n28050 = ~pi215 & ~n28049;
  assign n28051 = ~n28046 & n28050;
  assign n28052 = n7214 & n27982;
  assign n28053 = n7176 & n27977;
  assign n28054 = ~n27616 & ~n28053;
  assign n28055 = ~n28052 & n28054;
  assign n28056 = pi634 & ~n28055;
  assign n28057 = ~pi634 & n27616;
  assign n28058 = ~n27601 & ~n28057;
  assign n28059 = ~n28056 & n28058;
  assign n28060 = ~n2814 & ~n28059;
  assign n28061 = ~n28003 & ~n28060;
  assign n28062 = pi603 & ~n28061;
  assign n28063 = n7186 & ~n28010;
  assign n28064 = ~n28062 & n28063;
  assign n28065 = ~n7186 & n28016;
  assign n28066 = n7365 & ~n28065;
  assign n28067 = ~n28064 & n28066;
  assign n28068 = ~pi680 & n27607;
  assign n28069 = ~pi603 & ~n27815;
  assign n28070 = ~n28062 & ~n28069;
  assign n28071 = n2907 & ~n28070;
  assign n28072 = ~n28068 & ~n28071;
  assign n28073 = ~n28067 & ~n28068;
  assign n28074 = ~n28071 & n28073;
  assign n28075 = ~n28067 & n28072;
  assign n28076 = n62393 & n63931;
  assign n28077 = pi603 & ~n28059;
  assign n28078 = n7186 & n28077;
  assign n28079 = ~n28029 & ~n28059;
  assign n28080 = ~n28078 & ~n28079;
  assign n28081 = ~n28030 & ~n28059;
  assign n28082 = ~pi603 & n27826;
  assign n28083 = ~n28031 & ~n28082;
  assign n28084 = n63932 & n28083;
  assign n28085 = n7365 & ~n28084;
  assign n28086 = ~pi680 & ~n27614;
  assign n28087 = pi603 & n28059;
  assign n28088 = ~pi603 & n27813;
  assign n28089 = n2907 & ~n28088;
  assign n28090 = ~pi603 & ~n27813;
  assign n28091 = ~n28077 & ~n28090;
  assign n28092 = n2907 & ~n28091;
  assign n28093 = ~n28087 & n28089;
  assign n28094 = ~n28086 & ~n63933;
  assign n28095 = ~n28085 & n28094;
  assign n28096 = ~n62393 & n28095;
  assign n28097 = pi215 & ~n28096;
  assign n28098 = ~n28076 & n28097;
  assign n28099 = ~n28051 & ~n28098;
  assign n28100 = pi299 & ~n28099;
  assign n28101 = n2971 & n28025;
  assign n28102 = ~n2971 & ~n63930;
  assign n28103 = ~n7034 & ~n28102;
  assign n28104 = ~n28101 & n28103;
  assign n28105 = n7034 & n28048;
  assign n28106 = ~pi223 & ~n28105;
  assign n28107 = ~n28104 & n28106;
  assign n28108 = n2971 & n63931;
  assign n28109 = ~n2971 & n28095;
  assign n28110 = pi223 & ~n28109;
  assign n28111 = ~n28108 & n28110;
  assign n28112 = ~n28107 & ~n28111;
  assign n28113 = ~pi299 & ~n28112;
  assign n28114 = pi39 & ~n28113;
  assign n28115 = pi39 & ~n28100;
  assign n28116 = ~n28113 & n28115;
  assign n28117 = ~n28100 & n28114;
  assign n28118 = ~n27999 & ~n63934;
  assign n28119 = ~pi38 & ~n28118;
  assign n28120 = pi634 & n62857;
  assign n28121 = n27709 & ~n28120;
  assign n28122 = ~pi39 & ~n28121;
  assign n28123 = n27705 & ~n28122;
  assign n28124 = n62765 & ~n28123;
  assign n28125 = ~n28119 & n28124;
  assign n28126 = ~n27592 & ~n28125;
  assign n28127 = ~pi625 & n28126;
  assign n28128 = pi625 & n27714;
  assign n28129 = ~pi1153 & ~n28128;
  assign n28130 = ~n28127 & n28129;
  assign n28131 = ~pi608 & ~n27899;
  assign n28132 = ~n28130 & n28131;
  assign n28133 = pi625 & n28126;
  assign n28134 = ~pi625 & n27714;
  assign n28135 = pi1153 & ~n28134;
  assign n28136 = ~n28133 & n28135;
  assign n28137 = pi608 & ~n27903;
  assign n28138 = ~n28136 & n28137;
  assign n28139 = ~n28132 & ~n28138;
  assign n28140 = pi778 & ~n28139;
  assign n28141 = ~pi778 & n28126;
  assign n28142 = ~n28140 & ~n28141;
  assign n28143 = ~pi609 & ~n28142;
  assign n28144 = pi609 & n27906;
  assign n28145 = ~pi1155 & ~n28144;
  assign n28146 = ~n28143 & n28145;
  assign n28147 = ~pi660 & ~n27722;
  assign n28148 = ~n28146 & n28147;
  assign n28149 = pi609 & ~n28142;
  assign n28150 = ~pi609 & n27906;
  assign n28151 = pi1155 & ~n28150;
  assign n28152 = ~n28149 & n28151;
  assign n28153 = pi660 & ~n27726;
  assign n28154 = ~n28152 & n28153;
  assign n28155 = ~n28148 & ~n28154;
  assign n28156 = pi785 & ~n28155;
  assign n28157 = ~pi785 & ~n28142;
  assign n28158 = ~n28156 & ~n28157;
  assign n28159 = pi618 & ~n28158;
  assign n28160 = ~pi618 & n63923;
  assign n28161 = pi1154 & ~n28160;
  assign n28162 = ~n28159 & n28161;
  assign n28163 = pi627 & ~n27738;
  assign n28164 = ~n28162 & n28163;
  assign n28165 = ~pi618 & ~n28158;
  assign n28166 = pi618 & n63923;
  assign n28167 = ~pi1154 & ~n28166;
  assign n28168 = ~n28165 & n28167;
  assign n28169 = ~pi627 & ~n27734;
  assign n28170 = ~n28168 & n28169;
  assign n28171 = pi781 & ~n28170;
  assign n28172 = ~n28164 & n28171;
  assign n28173 = n8253 & ~n27746;
  assign n28174 = ~n27745 & n28173;
  assign n28175 = n8254 & ~n27750;
  assign n28176 = ~n27749 & n28175;
  assign n28177 = ~n11431 & n63924;
  assign n28178 = ~n28176 & ~n28177;
  assign n28179 = ~n28174 & n28178;
  assign n28180 = pi789 & ~n28179;
  assign n28181 = ~pi781 & n28158;
  assign n28182 = ~n28180 & ~n28181;
  assign n28183 = ~n28172 & n28182;
  assign n28184 = n11434 & n28179;
  assign n28185 = ~n28183 & ~n28184;
  assign n28186 = ~n28164 & ~n28170;
  assign n28187 = pi781 & ~n28186;
  assign n28188 = ~pi781 & ~n28158;
  assign n28189 = ~n28187 & ~n28188;
  assign n28190 = ~pi619 & ~n28189;
  assign n28191 = pi619 & ~n63924;
  assign n28192 = ~pi1159 & ~n28191;
  assign n28193 = ~n28190 & n28192;
  assign n28194 = ~pi648 & ~n27748;
  assign n28195 = ~n28193 & n28194;
  assign n28196 = pi619 & ~n28189;
  assign n28197 = ~pi619 & ~n63924;
  assign n28198 = pi1159 & ~n28197;
  assign n28199 = ~n28196 & n28198;
  assign n28200 = pi648 & ~n27752;
  assign n28201 = ~n28199 & n28200;
  assign n28202 = pi789 & ~n28201;
  assign n28203 = pi789 & ~n28195;
  assign n28204 = ~n28201 & n28203;
  assign n28205 = ~n28195 & n28202;
  assign n28206 = ~pi789 & n28189;
  assign n28207 = n62894 & ~n28206;
  assign n28208 = ~n63935 & n28207;
  assign n28209 = n62894 & ~n28185;
  assign n28210 = ~n27952 & ~n63936;
  assign n28211 = ~n27936 & ~n28210;
  assign n28212 = n63030 & n27935;
  assign n28213 = ~n8651 & ~n28212;
  assign n28214 = ~n28211 & n28213;
  assign n28215 = ~pi792 & n27920;
  assign n28216 = ~n63925 & ~n27932;
  assign n28217 = pi792 & ~n28216;
  assign n28218 = ~n28215 & ~n28217;
  assign n28219 = ~pi647 & n28218;
  assign n28220 = pi647 & n27590;
  assign n28221 = ~pi1157 & ~n28220;
  assign n28222 = ~n28219 & n28221;
  assign n28223 = pi630 & n28222;
  assign n28224 = pi647 & ~n28218;
  assign n28225 = ~pi647 & ~n27590;
  assign n28226 = ~n28224 & ~n28225;
  assign n28227 = n8373 & ~n28226;
  assign n28228 = ~n8334 & ~n63912;
  assign n28229 = n8334 & n27590;
  assign n28230 = ~n8413 & ~n28229;
  assign n28231 = n8334 & ~n27590;
  assign n28232 = ~n8334 & n63912;
  assign n28233 = ~n28231 & ~n28232;
  assign n28234 = ~n8413 & ~n28233;
  assign n28235 = ~n28228 & n28230;
  assign n28236 = ~n28227 & ~n63937;
  assign n28237 = ~n28223 & ~n28227;
  assign n28238 = ~n63937 & n28237;
  assign n28239 = ~n28223 & n28236;
  assign n28240 = pi787 & ~n63938;
  assign n28241 = ~n11547 & ~n28240;
  assign n28242 = ~n28214 & ~n28240;
  assign n28243 = ~n11547 & n28242;
  assign n28244 = ~n28214 & n28241;
  assign n28245 = pi1157 & ~n28226;
  assign n28246 = ~n28222 & ~n28245;
  assign n28247 = pi787 & ~n28246;
  assign n28248 = ~pi787 & ~n28218;
  assign n28249 = ~n63036 & ~n28248;
  assign n28250 = ~n28247 & n28249;
  assign n28251 = n11558 & n63792;
  assign n28252 = ~n63911 & n28251;
  assign n28253 = ~n27590 & ~n28251;
  assign n28254 = ~n25932 & ~n28253;
  assign n28255 = ~n25932 & ~n28251;
  assign n28256 = n27590 & n28255;
  assign n28257 = n11558 & n63793;
  assign n28258 = n63911 & n28257;
  assign n28259 = ~n28256 & ~n28258;
  assign n28260 = ~n28252 & n28254;
  assign n28261 = ~n28250 & n63940;
  assign n28262 = pi790 & ~n28261;
  assign n28263 = n62455 & ~n28262;
  assign n28264 = ~pi790 & ~n28242;
  assign n28265 = ~n63939 & n28261;
  assign n28266 = pi644 & n28242;
  assign n28267 = ~n28247 & ~n28248;
  assign n28268 = ~pi644 & n28267;
  assign n28269 = pi715 & ~n28268;
  assign n28270 = ~n28266 & n28269;
  assign n28271 = ~n8376 & n28233;
  assign n28272 = n8376 & n27590;
  assign n28273 = ~n28271 & ~n28272;
  assign n28274 = pi644 & ~n28273;
  assign n28275 = ~pi644 & n27590;
  assign n28276 = ~pi715 & ~n28275;
  assign n28277 = ~n28274 & n28276;
  assign n28278 = pi1160 & ~n28277;
  assign n28279 = ~n28270 & n28278;
  assign n28280 = ~pi644 & n28242;
  assign n28281 = pi644 & n28267;
  assign n28282 = ~pi715 & ~n28281;
  assign n28283 = ~n28280 & n28282;
  assign n28284 = ~pi644 & ~n28273;
  assign n28285 = pi644 & n27590;
  assign n28286 = pi715 & ~n28285;
  assign n28287 = ~n28284 & n28286;
  assign n28288 = ~pi1160 & ~n28287;
  assign n28289 = ~n28283 & n28288;
  assign n28290 = pi790 & ~n28289;
  assign n28291 = pi790 & ~n28279;
  assign n28292 = ~n28289 & n28291;
  assign n28293 = ~n28279 & n28290;
  assign n28294 = ~n28264 & ~n63941;
  assign n28295 = ~n28264 & ~n28265;
  assign n28296 = n62455 & ~n63942;
  assign n28297 = ~n63939 & n28263;
  assign n28298 = ~n27542 & ~n63943;
  assign n28299 = pi222 & ~n62455;
  assign n28300 = pi222 & ~n62765;
  assign n28301 = pi616 & ~n7523;
  assign n28302 = ~n2814 & n7082;
  assign n28303 = ~n7056 & ~n28302;
  assign n28304 = ~pi616 & n28303;
  assign n28305 = ~n28301 & ~n28304;
  assign n28306 = ~n7007 & ~n28305;
  assign n28307 = ~n2905 & n28305;
  assign n28308 = pi616 & n7187;
  assign n28309 = n7197 & ~n28308;
  assign n28310 = ~n7179 & ~n28309;
  assign n28311 = n2905 & ~n28310;
  assign n28312 = n7007 & ~n28311;
  assign n28313 = ~n28307 & n28312;
  assign n28314 = ~n28306 & ~n28313;
  assign n28315 = ~n2971 & n28314;
  assign n28316 = pi616 & ~n7188;
  assign n28317 = ~n7083 & ~n28316;
  assign n28318 = ~n7007 & ~n28317;
  assign n28319 = ~n2905 & n28317;
  assign n28320 = n2905 & ~n28308;
  assign n28321 = n7076 & n28320;
  assign n28322 = n7007 & ~n28321;
  assign n28323 = ~n28319 & n28322;
  assign n28324 = ~n28318 & ~n28323;
  assign n28325 = n2971 & n28324;
  assign n28326 = pi222 & ~n28325;
  assign n28327 = ~n28315 & n28326;
  assign n28328 = ~n7057 & n28308;
  assign n28329 = ~n7007 & ~n28328;
  assign n28330 = ~n2905 & n28328;
  assign n28331 = pi616 & n2905;
  assign n28332 = n7398 & n28331;
  assign n28333 = n7007 & ~n28332;
  assign n28334 = ~n28330 & n28333;
  assign n28335 = ~n28329 & ~n28334;
  assign n28336 = ~n2971 & n28335;
  assign n28337 = ~n2907 & ~n7298;
  assign n28338 = ~n2907 & n7298;
  assign n28339 = ~n7306 & ~n28338;
  assign n28340 = ~n7297 & ~n28337;
  assign n28341 = pi616 & ~n63944;
  assign n28342 = n2971 & n28341;
  assign n28343 = pi224 & ~n28342;
  assign n28344 = pi224 & ~n28336;
  assign n28345 = ~n28342 & n28344;
  assign n28346 = ~n28336 & n28343;
  assign n28347 = n7021 & n7187;
  assign n28348 = ~pi224 & ~n28347;
  assign n28349 = ~pi222 & ~n28348;
  assign n28350 = ~n63945 & n28349;
  assign n28351 = ~pi223 & ~n28350;
  assign n28352 = ~n28327 & n28351;
  assign n28353 = ~n6991 & ~n28316;
  assign n28354 = ~n7007 & ~n28353;
  assign n28355 = ~n2905 & n28353;
  assign n28356 = n6979 & n28320;
  assign n28357 = n7007 & ~n28356;
  assign n28358 = ~n28355 & n28357;
  assign n28359 = ~n28354 & ~n28358;
  assign n28360 = n2971 & n28359;
  assign n28361 = pi616 & ~n7224;
  assign n28362 = n62783 & ~n28361;
  assign n28363 = ~n7007 & ~n28362;
  assign n28364 = ~n2905 & ~n62783;
  assign n28365 = ~n6994 & ~n28361;
  assign n28366 = ~n28364 & n28365;
  assign n28367 = n7007 & ~n28366;
  assign n28368 = ~n28363 & ~n28367;
  assign n28369 = ~n2971 & n28368;
  assign n28370 = pi222 & ~n28369;
  assign n28371 = pi222 & ~n28360;
  assign n28372 = ~n28369 & n28371;
  assign n28373 = ~n28360 & n28370;
  assign n28374 = n6994 & n7007;
  assign n28375 = ~n2814 & n28374;
  assign n28376 = n2907 & n6978;
  assign n28377 = ~n7322 & ~n28338;
  assign n28378 = pi616 & ~n28377;
  assign n28379 = n28347 & ~n63947;
  assign n28380 = ~pi222 & n63948;
  assign n28381 = ~n7344 & n28380;
  assign n28382 = pi223 & ~n28381;
  assign n28383 = ~n63946 & n28382;
  assign n28384 = ~n28352 & ~n28383;
  assign n28385 = ~pi299 & ~n28384;
  assign n28386 = ~n62393 & n28314;
  assign n28387 = n62393 & n28324;
  assign n28388 = pi222 & ~n28387;
  assign n28389 = ~n28386 & n28388;
  assign n28390 = n62393 & ~n28341;
  assign n28391 = ~n62393 & ~n28335;
  assign n28392 = ~pi222 & ~n28391;
  assign n28393 = ~pi222 & ~n28390;
  assign n28394 = ~n28391 & n28393;
  assign n28395 = ~n28390 & n28392;
  assign n28396 = ~n7118 & ~n63949;
  assign n28397 = ~n28389 & n28396;
  assign n28398 = pi222 & ~n6951;
  assign n28399 = n7118 & ~n28398;
  assign n28400 = ~n28347 & n28399;
  assign n28401 = ~pi215 & ~n28400;
  assign n28402 = ~n28397 & n28401;
  assign n28403 = ~n7328 & n28380;
  assign n28404 = n62393 & n28359;
  assign n28405 = ~n62393 & n28368;
  assign n28406 = pi222 & ~n28405;
  assign n28407 = pi222 & ~n28404;
  assign n28408 = ~n28405 & n28407;
  assign n28409 = ~n28404 & n28406;
  assign n28410 = ~n28403 & ~n63950;
  assign n28411 = pi215 & ~n28410;
  assign n28412 = pi299 & ~n28411;
  assign n28413 = ~n28402 & n28412;
  assign n28414 = pi39 & ~n28413;
  assign n28415 = pi39 & ~n28385;
  assign n28416 = ~n28413 & n28415;
  assign n28417 = ~n28385 & n28414;
  assign n28418 = pi222 & n62793;
  assign n28419 = ~pi616 & n7292;
  assign n28420 = ~pi222 & ~n7292;
  assign n28421 = ~pi39 & ~n28420;
  assign n28422 = ~pi39 & ~n28419;
  assign n28423 = ~n28420 & n28422;
  assign n28424 = ~n28419 & n28421;
  assign n28425 = ~n28418 & n63952;
  assign n28426 = ~pi38 & ~n28425;
  assign n28427 = ~n63951 & n28426;
  assign n28428 = pi222 & ~n7357;
  assign n28429 = pi38 & ~n28428;
  assign n28430 = pi616 & n7359;
  assign n28431 = n7357 & n28308;
  assign n28432 = n28429 & ~n63953;
  assign n28433 = n62765 & ~n28432;
  assign n28434 = ~n28427 & n28433;
  assign n28435 = ~n28300 & ~n28434;
  assign n28436 = ~n8135 & ~n28435;
  assign n28437 = ~pi223 & ~n62789;
  assign n28438 = ~n7033 & ~n28437;
  assign n28439 = ~pi299 & ~n28438;
  assign n28440 = pi39 & ~n28439;
  assign n28441 = ~n7142 & n28440;
  assign n28442 = ~pi38 & ~n6946;
  assign n28443 = ~n28441 & n28442;
  assign n28444 = n9733 & ~n28443;
  assign n28445 = pi222 & ~n28444;
  assign n28446 = n8135 & n28445;
  assign n28447 = n8135 & ~n28445;
  assign n28448 = ~n8135 & n28435;
  assign n28449 = ~n28447 & ~n28448;
  assign n28450 = ~n28436 & ~n28446;
  assign n28451 = ~pi785 & n63954;
  assign n28452 = pi609 & ~n63954;
  assign n28453 = ~pi609 & ~n28445;
  assign n28454 = pi1155 & ~n28453;
  assign n28455 = ~n28452 & n28454;
  assign n28456 = ~pi609 & ~n63954;
  assign n28457 = pi609 & ~n28445;
  assign n28458 = ~pi1155 & ~n28457;
  assign n28459 = ~n28456 & n28458;
  assign n28460 = ~n28455 & ~n28459;
  assign n28461 = pi785 & ~n28460;
  assign n28462 = ~n28451 & ~n28461;
  assign n28463 = ~pi781 & ~n28462;
  assign n28464 = pi618 & n28462;
  assign n28465 = ~pi618 & ~n28445;
  assign n28466 = pi1154 & ~n28465;
  assign n28467 = ~n28464 & n28466;
  assign n28468 = ~pi618 & n28462;
  assign n28469 = pi618 & ~n28445;
  assign n28470 = ~pi1154 & ~n28469;
  assign n28471 = ~n28468 & n28470;
  assign n28472 = ~n28467 & ~n28471;
  assign n28473 = pi781 & ~n28472;
  assign n28474 = ~n28463 & ~n28473;
  assign n28475 = pi619 & n28474;
  assign n28476 = ~pi619 & ~n28445;
  assign n28477 = pi1159 & ~n28476;
  assign n28478 = ~n28475 & n28477;
  assign n28479 = ~pi619 & n28474;
  assign n28480 = pi619 & ~n28445;
  assign n28481 = ~pi1159 & ~n28480;
  assign n28482 = ~n28479 & n28481;
  assign n28483 = ~n28479 & ~n28480;
  assign n28484 = ~pi1159 & ~n28483;
  assign n28485 = ~n28475 & ~n28476;
  assign n28486 = pi1159 & ~n28485;
  assign n28487 = ~n28484 & ~n28486;
  assign n28488 = ~n28478 & ~n28482;
  assign n28489 = pi789 & ~n63955;
  assign n28490 = ~pi789 & n28474;
  assign n28491 = ~pi789 & ~n28474;
  assign n28492 = pi789 & n63955;
  assign n28493 = ~n28491 & ~n28492;
  assign n28494 = ~n28489 & ~n28490;
  assign n28495 = ~n8595 & n63956;
  assign n28496 = n8595 & ~n28445;
  assign n28497 = ~n28495 & ~n28496;
  assign n28498 = ~n63052 & n28497;
  assign n28499 = ~n10206 & ~n28445;
  assign n28500 = ~pi222 & ~n7849;
  assign n28501 = pi661 & pi680;
  assign n28502 = n7849 & ~n28501;
  assign n28503 = pi222 & n7826;
  assign n28504 = pi299 & ~n28503;
  assign n28505 = ~n28502 & n28504;
  assign n28506 = ~n28500 & n28504;
  assign n28507 = ~n28502 & n28506;
  assign n28508 = ~n28500 & n28505;
  assign n28509 = ~pi222 & ~n7840;
  assign n28510 = n7840 & ~n28501;
  assign n28511 = pi222 & n7820;
  assign n28512 = ~pi299 & ~n28511;
  assign n28513 = ~n28510 & n28512;
  assign n28514 = ~n28509 & n28512;
  assign n28515 = ~n28510 & n28514;
  assign n28516 = ~n28509 & n28513;
  assign n28517 = ~pi39 & ~n63958;
  assign n28518 = ~pi39 & ~n63957;
  assign n28519 = ~n63958 & n28518;
  assign n28520 = ~n63957 & n28517;
  assign n28521 = ~n2905 & ~n7084;
  assign n28522 = ~pi662 & n7095;
  assign n28523 = ~n28521 & ~n28522;
  assign n28524 = n7007 & ~n28523;
  assign n28525 = ~pi661 & n7085;
  assign n28526 = pi661 & ~n7937;
  assign n28527 = ~n28525 & ~n28526;
  assign n28528 = ~n28524 & ~n28525;
  assign n28529 = ~n28526 & n28528;
  assign n28530 = ~n28524 & n28527;
  assign n28531 = n2971 & n63960;
  assign n28532 = ~pi661 & ~n62787;
  assign n28533 = pi680 & n7731;
  assign n28534 = ~n7397 & ~n28533;
  assign n28535 = pi661 & ~n28534;
  assign n28536 = ~n28532 & ~n28535;
  assign n28537 = ~n2971 & n28536;
  assign n28538 = pi222 & ~n28537;
  assign n28539 = ~n28531 & n28538;
  assign n28540 = pi661 & n8013;
  assign n28541 = ~n2971 & n28540;
  assign n28542 = ~n8018 & n28501;
  assign n28543 = n2971 & n28542;
  assign n28544 = pi224 & ~n28543;
  assign n28545 = pi224 & ~n28541;
  assign n28546 = ~n28543 & n28545;
  assign n28547 = ~n28541 & n28544;
  assign n28548 = pi661 & n62828;
  assign n28549 = n7544 & n28501;
  assign n28550 = ~pi224 & ~n63962;
  assign n28551 = ~pi222 & ~n28550;
  assign n28552 = ~n63961 & n28551;
  assign n28553 = ~pi223 & ~n28552;
  assign n28554 = ~n28539 & n28553;
  assign n28555 = ~pi661 & ~n62784;
  assign n28556 = pi661 & ~n7959;
  assign n28557 = ~n28555 & ~n28556;
  assign n28558 = n2971 & n28557;
  assign n28559 = n6997 & n7007;
  assign n28560 = ~pi661 & n6987;
  assign n28561 = pi661 & ~n7964;
  assign n28562 = ~n28560 & ~n28561;
  assign n28563 = ~n28559 & n28562;
  assign n28564 = ~n2971 & n28563;
  assign n28565 = pi222 & ~n28564;
  assign n28566 = ~n28558 & n28565;
  assign n28567 = ~pi222 & pi661;
  assign n28568 = n8031 & n28567;
  assign n28569 = pi223 & ~n28568;
  assign n28570 = ~n28566 & n28569;
  assign n28571 = ~n28554 & ~n28570;
  assign n28572 = ~pi299 & ~n28571;
  assign n28573 = n62393 & n63960;
  assign n28574 = ~n62393 & n28536;
  assign n28575 = pi222 & ~n28574;
  assign n28576 = ~n28573 & n28575;
  assign n28577 = n62393 & ~n28542;
  assign n28578 = ~n62393 & ~n28540;
  assign n28579 = ~pi222 & ~n28578;
  assign n28580 = ~pi222 & ~n28577;
  assign n28581 = ~n28578 & n28580;
  assign n28582 = ~n28577 & n28579;
  assign n28583 = ~n7118 & ~n63963;
  assign n28584 = ~n28576 & n28583;
  assign n28585 = n28399 & ~n63962;
  assign n28586 = ~pi215 & ~n28585;
  assign n28587 = ~n28584 & n28586;
  assign n28588 = n8052 & n28567;
  assign n28589 = n62393 & n28557;
  assign n28590 = ~n62393 & n28563;
  assign n28591 = pi222 & ~n28590;
  assign n28592 = ~n28589 & n28591;
  assign n28593 = ~n28588 & ~n28592;
  assign n28594 = pi215 & ~n28593;
  assign n28595 = pi299 & ~n28594;
  assign n28596 = ~n28587 & n28595;
  assign n28597 = ~n28572 & ~n28596;
  assign n28598 = pi39 & ~n28597;
  assign n28599 = ~n63959 & ~n28598;
  assign n28600 = ~pi38 & ~n28599;
  assign n28601 = pi661 & n8084;
  assign n28602 = n28429 & ~n28601;
  assign n28603 = n62765 & ~n28602;
  assign n28604 = ~n28600 & n28603;
  assign n28605 = ~n28300 & ~n28604;
  assign n28606 = ~pi778 & ~n28605;
  assign n28607 = pi625 & n28605;
  assign n28608 = ~pi625 & ~n28445;
  assign n28609 = pi1153 & ~n28608;
  assign n28610 = ~n28607 & n28609;
  assign n28611 = ~pi625 & n28605;
  assign n28612 = pi625 & ~n28445;
  assign n28613 = ~pi1153 & ~n28612;
  assign n28614 = ~n28611 & n28613;
  assign n28615 = ~n28610 & ~n28614;
  assign n28616 = pi778 & ~n28615;
  assign n28617 = ~n28606 & ~n28616;
  assign n28618 = ~n62880 & ~n28617;
  assign n28619 = n62880 & n28445;
  assign n28620 = n62880 & ~n28445;
  assign n28621 = ~n62880 & n28617;
  assign n28622 = ~n28620 & ~n28621;
  assign n28623 = ~n28618 & ~n28619;
  assign n28624 = ~n62882 & n63964;
  assign n28625 = n62882 & n28445;
  assign n28626 = ~n62882 & ~n63964;
  assign n28627 = n62882 & ~n28445;
  assign n28628 = ~n28626 & ~n28627;
  assign n28629 = ~n28624 & ~n28625;
  assign n28630 = ~n8257 & ~n63965;
  assign n28631 = ~n8303 & n28630;
  assign n28632 = ~n28499 & ~n28631;
  assign n28633 = ~pi628 & ~n28632;
  assign n28634 = pi628 & ~n28445;
  assign n28635 = n8332 & ~n28634;
  assign n28636 = ~n28633 & n28635;
  assign n28637 = pi628 & ~n28632;
  assign n28638 = ~pi628 & ~n28445;
  assign n28639 = n8331 & ~n28638;
  assign n28640 = ~n28637 & n28639;
  assign n28641 = ~n28636 & ~n28640;
  assign n28642 = ~n28498 & n28641;
  assign n28643 = pi792 & ~n28642;
  assign n28644 = n8253 & n28485;
  assign n28645 = ~n11431 & n63965;
  assign n28646 = n8254 & n28483;
  assign n28647 = ~n28645 & ~n28646;
  assign n28648 = ~n28644 & n28647;
  assign n28649 = pi789 & ~n28648;
  assign n28650 = pi616 & ~n7712;
  assign n28651 = pi680 & ~n28650;
  assign n28652 = ~n7377 & n28651;
  assign n28653 = ~pi680 & n28317;
  assign n28654 = pi661 & ~n28653;
  assign n28655 = pi661 & ~n28652;
  assign n28656 = ~n28653 & n28655;
  assign n28657 = ~n28652 & n28654;
  assign n28658 = ~pi661 & pi681;
  assign n28659 = ~n28317 & n28658;
  assign n28660 = ~n28323 & ~n28659;
  assign n28661 = ~n63966 & n28660;
  assign n28662 = pi222 & ~n28661;
  assign n28663 = pi616 & ~n7653;
  assign n28664 = pi680 & ~n7556;
  assign n28665 = ~n28663 & n28664;
  assign n28666 = ~pi680 & n28347;
  assign n28667 = pi661 & ~n28666;
  assign n28668 = ~n28665 & n28667;
  assign n28669 = ~pi661 & ~n28347;
  assign n28670 = ~n2907 & ~n28669;
  assign n28671 = ~pi681 & n28331;
  assign n28672 = n7296 & n28671;
  assign n28673 = n7296 & n28331;
  assign n28674 = ~n2905 & n28347;
  assign n28675 = n7007 & ~n28674;
  assign n28676 = ~n28673 & n28675;
  assign n28677 = ~n28347 & n28658;
  assign n28678 = ~n28676 & ~n28677;
  assign n28679 = ~n28670 & ~n28672;
  assign n28680 = ~n28668 & n63967;
  assign n28681 = ~pi222 & n28680;
  assign n28682 = n62393 & ~n28681;
  assign n28683 = ~n28662 & n28682;
  assign n28684 = ~pi680 & n28305;
  assign n28685 = n2814 & n7383;
  assign n28686 = ~n7427 & ~n28685;
  assign n28687 = n7366 & ~n7519;
  assign n28688 = ~n7638 & n63968;
  assign n28689 = pi642 & ~n28688;
  assign n28690 = ~pi603 & n63968;
  assign n28691 = pi603 & n7055;
  assign n28692 = ~n7388 & ~n28691;
  assign n28693 = ~n28690 & n28692;
  assign n28694 = ~pi642 & n28693;
  assign n28695 = n2903 & ~n28694;
  assign n28696 = n2903 & ~n28689;
  assign n28697 = ~n28694 & n28696;
  assign n28698 = ~n28689 & n28695;
  assign n28699 = n7591 & n28688;
  assign n28700 = n7652 & ~n63968;
  assign n28701 = ~n7519 & n7652;
  assign n28702 = pi616 & ~n63970;
  assign n28703 = pi680 & ~n28702;
  assign n28704 = ~n28699 & n28703;
  assign n28705 = ~n63969 & n28704;
  assign n28706 = pi661 & ~n28705;
  assign n28707 = ~n28684 & n28706;
  assign n28708 = ~n28305 & n28658;
  assign n28709 = ~n28313 & ~n28708;
  assign n28710 = ~n28707 & n28709;
  assign n28711 = pi222 & ~n28710;
  assign n28712 = pi616 & n7639;
  assign n28713 = pi680 & ~n28712;
  assign n28714 = ~n62825 & n28713;
  assign n28715 = ~pi680 & n28328;
  assign n28716 = pi661 & ~n28715;
  assign n28717 = ~n28714 & n28716;
  assign n28718 = ~n28328 & n28658;
  assign n28719 = ~n28334 & ~n28718;
  assign n28720 = ~n28717 & n28719;
  assign n28721 = ~pi222 & n28720;
  assign n28722 = ~n62393 & ~n28721;
  assign n28723 = ~n28711 & n28722;
  assign n28724 = ~n62393 & ~n28710;
  assign n28725 = n62393 & ~n28661;
  assign n28726 = pi222 & ~n28725;
  assign n28727 = ~n28724 & n28726;
  assign n28728 = ~n62393 & n28720;
  assign n28729 = n62393 & n28680;
  assign n28730 = ~pi222 & ~n28729;
  assign n28731 = ~n28728 & n28730;
  assign n28732 = ~n28727 & ~n28731;
  assign n28733 = ~n28683 & ~n28723;
  assign n28734 = ~n7118 & ~n63971;
  assign n28735 = ~n28308 & ~n28501;
  assign n28736 = ~pi616 & ~n62826;
  assign n28737 = ~n28663 & ~n28736;
  assign n28738 = ~n28347 & ~n28501;
  assign n28739 = n28501 & ~n28737;
  assign n28740 = ~n28738 & ~n28739;
  assign n28741 = ~n28735 & n28737;
  assign n28742 = n28399 & ~n63972;
  assign n28743 = ~pi215 & ~n28742;
  assign n28744 = ~n28734 & n28743;
  assign n28745 = ~n7440 & n28651;
  assign n28746 = ~pi680 & n28353;
  assign n28747 = pi661 & ~n28746;
  assign n28748 = ~n28745 & n28747;
  assign n28749 = ~n28353 & n28658;
  assign n28750 = ~n28358 & ~n28749;
  assign n28751 = ~n28748 & n28750;
  assign n28752 = n62393 & ~n28751;
  assign n28753 = ~pi680 & n28362;
  assign n28754 = ~n7449 & n7652;
  assign n28755 = pi616 & ~n28754;
  assign n28756 = pi680 & ~n28755;
  assign n28757 = n7453 & n28756;
  assign n28758 = pi661 & ~n28757;
  assign n28759 = ~n28753 & n28758;
  assign n28760 = ~n28362 & n28658;
  assign n28761 = ~n28367 & ~n28760;
  assign n28762 = ~n28759 & n28761;
  assign n28763 = ~n62393 & ~n28762;
  assign n28764 = pi222 & ~n28763;
  assign n28765 = pi222 & ~n28752;
  assign n28766 = ~n28763 & n28765;
  assign n28767 = ~n28752 & n28764;
  assign n28768 = ~n7323 & ~n7690;
  assign n28769 = pi616 & n28768;
  assign n28770 = ~n6971 & n28347;
  assign n28771 = pi616 & n7425;
  assign n28772 = n2907 & ~n63974;
  assign n28773 = n6973 & ~n28501;
  assign n28774 = ~n28738 & ~n28773;
  assign n28775 = ~n28772 & n28774;
  assign n28776 = ~n28769 & n28775;
  assign n28777 = pi680 & ~n28769;
  assign n28778 = n62832 & n28777;
  assign n28779 = pi616 & n7323;
  assign n28780 = ~n6973 & n28347;
  assign n28781 = ~pi680 & n63975;
  assign n28782 = pi661 & ~n28781;
  assign n28783 = ~n28778 & n28782;
  assign n28784 = ~pi661 & ~n63975;
  assign n28785 = ~n28772 & ~n28784;
  assign n28786 = ~n28783 & n28785;
  assign n28787 = n62832 & n28776;
  assign n28788 = ~n62393 & n63976;
  assign n28789 = n7576 & n28501;
  assign n28790 = ~n63948 & ~n28789;
  assign n28791 = n62393 & ~n28790;
  assign n28792 = ~pi222 & ~n28791;
  assign n28793 = ~n28788 & n28792;
  assign n28794 = pi215 & ~n28793;
  assign n28795 = ~n63973 & n28794;
  assign n28796 = pi299 & ~n28795;
  assign n28797 = ~n28744 & n28796;
  assign n28798 = ~n2971 & n28710;
  assign n28799 = n2971 & n28661;
  assign n28800 = pi222 & ~n28799;
  assign n28801 = ~n28798 & n28800;
  assign n28802 = ~n2971 & n28720;
  assign n28803 = n2971 & n28680;
  assign n28804 = pi224 & ~n28803;
  assign n28805 = ~n28802 & n28804;
  assign n28806 = n28501 & n28737;
  assign n28807 = n28347 & ~n28501;
  assign n28808 = ~pi224 & ~n28807;
  assign n28809 = ~n28806 & n28808;
  assign n28810 = ~pi224 & ~n63972;
  assign n28811 = ~pi222 & pi224;
  assign n28812 = ~pi222 & ~n28738;
  assign n28813 = ~n28739 & n28812;
  assign n28814 = ~n28811 & ~n28813;
  assign n28815 = ~pi222 & ~n63977;
  assign n28816 = ~n28805 & ~n63978;
  assign n28817 = ~n28801 & ~n28816;
  assign n28818 = ~pi223 & ~n28817;
  assign n28819 = n2971 & ~n28751;
  assign n28820 = ~n2971 & ~n28762;
  assign n28821 = pi222 & ~n28820;
  assign n28822 = pi222 & ~n28819;
  assign n28823 = ~n28820 & n28822;
  assign n28824 = ~n28819 & n28821;
  assign n28825 = ~n2971 & n63976;
  assign n28826 = n2971 & ~n28790;
  assign n28827 = ~pi222 & ~n28826;
  assign n28828 = ~n28825 & n28827;
  assign n28829 = pi223 & ~n28828;
  assign n28830 = ~n63979 & n28829;
  assign n28831 = ~pi299 & ~n28830;
  assign n28832 = ~n28818 & n28831;
  assign n28833 = pi39 & ~n28832;
  assign n28834 = ~n28797 & n28833;
  assign n28835 = n7852 & ~n28501;
  assign n28836 = ~pi603 & ~n7826;
  assign n28837 = ~n7168 & ~n7387;
  assign n28838 = ~n28836 & n28837;
  assign n28839 = ~pi616 & n7290;
  assign n28840 = pi299 & ~n28839;
  assign n28841 = ~n28838 & n28840;
  assign n28842 = ~n28835 & n28841;
  assign n28843 = n7844 & ~n28501;
  assign n28844 = ~pi603 & ~n7820;
  assign n28845 = ~n7387 & ~n7842;
  assign n28846 = ~n28844 & n28845;
  assign n28847 = ~pi616 & n7285;
  assign n28848 = ~pi299 & ~n28847;
  assign n28849 = ~n28846 & n28848;
  assign n28850 = ~n28843 & n28849;
  assign n28851 = pi222 & ~n28850;
  assign n28852 = ~n28842 & n28851;
  assign n28853 = pi661 & n7845;
  assign n28854 = pi616 & n7285;
  assign n28855 = ~pi299 & ~n28854;
  assign n28856 = ~n28853 & n28855;
  assign n28857 = pi661 & n7853;
  assign n28858 = pi616 & n7290;
  assign n28859 = pi299 & ~n28858;
  assign n28860 = ~n28857 & n28859;
  assign n28861 = ~n28856 & ~n28860;
  assign n28862 = ~pi222 & ~n28861;
  assign n28863 = ~pi39 & ~n28862;
  assign n28864 = ~n28838 & ~n28839;
  assign n28865 = ~n28835 & n28864;
  assign n28866 = pi222 & ~n28865;
  assign n28867 = ~pi222 & ~n28858;
  assign n28868 = ~n28857 & n28867;
  assign n28869 = ~n28866 & ~n28868;
  assign n28870 = pi299 & ~n28869;
  assign n28871 = ~pi222 & ~n28854;
  assign n28872 = ~n28853 & n28871;
  assign n28873 = ~n28846 & ~n28847;
  assign n28874 = ~n28843 & n28873;
  assign n28875 = pi222 & ~n28874;
  assign n28876 = ~n28872 & ~n28875;
  assign n28877 = ~pi299 & ~n28876;
  assign n28878 = ~pi39 & ~n28877;
  assign n28879 = ~n28870 & n28878;
  assign n28880 = pi299 & ~n28866;
  assign n28881 = ~n28868 & n28880;
  assign n28882 = ~pi299 & ~n28875;
  assign n28883 = ~n28872 & n28882;
  assign n28884 = ~n28881 & ~n28883;
  assign n28885 = ~pi39 & ~n28884;
  assign n28886 = ~pi39 & ~n28870;
  assign n28887 = ~n28877 & n28886;
  assign n28888 = ~n28852 & n28863;
  assign n28889 = ~pi38 & ~n63980;
  assign n28890 = ~n28834 & n28889;
  assign n28891 = n6955 & n7652;
  assign n28892 = ~pi222 & ~pi616;
  assign n28893 = ~pi39 & pi616;
  assign n28894 = n28501 & n28893;
  assign n28895 = ~n28892 & ~n28894;
  assign n28896 = n28891 & ~n28895;
  assign n28897 = ~pi616 & ~n7408;
  assign n28898 = ~n28735 & ~n28897;
  assign n28899 = n7357 & n28898;
  assign n28900 = ~n28428 & ~n28899;
  assign n28901 = ~n28896 & ~n28900;
  assign n28902 = pi38 & ~n28901;
  assign n28903 = n62765 & ~n28902;
  assign n28904 = ~n28890 & n28903;
  assign n28905 = ~n28300 & ~n28904;
  assign n28906 = ~pi625 & n28905;
  assign n28907 = pi625 & n28435;
  assign n28908 = ~pi1153 & ~n28907;
  assign n28909 = ~n28906 & n28908;
  assign n28910 = ~pi608 & ~n28610;
  assign n28911 = ~n28909 & n28910;
  assign n28912 = pi625 & n28905;
  assign n28913 = ~pi625 & n28435;
  assign n28914 = pi1153 & ~n28913;
  assign n28915 = ~n28912 & n28914;
  assign n28916 = pi608 & ~n28614;
  assign n28917 = ~n28915 & n28916;
  assign n28918 = ~n28911 & ~n28917;
  assign n28919 = pi778 & ~n28918;
  assign n28920 = ~pi778 & n28905;
  assign n28921 = ~n28919 & ~n28920;
  assign n28922 = ~pi609 & ~n28921;
  assign n28923 = pi609 & n28617;
  assign n28924 = ~pi1155 & ~n28923;
  assign n28925 = ~n28922 & n28924;
  assign n28926 = ~pi660 & ~n28455;
  assign n28927 = ~n28925 & n28926;
  assign n28928 = pi609 & ~n28921;
  assign n28929 = ~pi609 & n28617;
  assign n28930 = pi1155 & ~n28929;
  assign n28931 = ~n28928 & n28930;
  assign n28932 = pi660 & ~n28459;
  assign n28933 = ~n28931 & n28932;
  assign n28934 = ~n28927 & ~n28933;
  assign n28935 = pi785 & ~n28934;
  assign n28936 = ~pi785 & ~n28921;
  assign n28937 = ~n28935 & ~n28936;
  assign n28938 = ~pi618 & ~n28937;
  assign n28939 = pi618 & ~n63964;
  assign n28940 = ~pi1154 & ~n28939;
  assign n28941 = ~n28938 & n28940;
  assign n28942 = ~pi627 & ~n28467;
  assign n28943 = ~n28941 & n28942;
  assign n28944 = pi618 & ~n28937;
  assign n28945 = ~pi618 & ~n63964;
  assign n28946 = pi1154 & ~n28945;
  assign n28947 = ~n28944 & n28946;
  assign n28948 = pi627 & ~n28471;
  assign n28949 = ~n28947 & n28948;
  assign n28950 = ~n28943 & ~n28949;
  assign n28951 = pi781 & ~n28950;
  assign n28952 = ~pi781 & ~n28937;
  assign n28953 = ~n11434 & ~n28952;
  assign n28954 = ~n28951 & n28953;
  assign n28955 = ~n28649 & ~n28954;
  assign n28956 = ~n28951 & ~n28952;
  assign n28957 = ~pi619 & ~n28956;
  assign n28958 = pi619 & ~n63965;
  assign n28959 = ~pi1159 & ~n28958;
  assign n28960 = ~n28957 & n28959;
  assign n28961 = ~pi648 & ~n28478;
  assign n28962 = ~n28960 & n28961;
  assign n28963 = pi619 & ~n28956;
  assign n28964 = ~pi619 & ~n63965;
  assign n28965 = pi1159 & ~n28964;
  assign n28966 = ~n28963 & n28965;
  assign n28967 = pi648 & ~n28482;
  assign n28968 = ~n28966 & n28967;
  assign n28969 = ~n28962 & ~n28968;
  assign n28970 = pi789 & ~n28969;
  assign n28971 = ~pi789 & ~n28956;
  assign n28972 = n62894 & ~n28971;
  assign n28973 = ~n28970 & n28972;
  assign n28974 = n62894 & ~n28955;
  assign n28975 = pi626 & n63956;
  assign n28976 = ~pi626 & ~n28445;
  assign n28977 = n8300 & ~n28976;
  assign n28978 = ~n28975 & n28977;
  assign n28979 = ~pi626 & n63956;
  assign n28980 = pi626 & ~n28445;
  assign n28981 = n8301 & ~n28980;
  assign n28982 = ~n28979 & n28981;
  assign n28983 = n8257 & ~n28445;
  assign n28984 = n8525 & ~n28983;
  assign n28985 = ~n28630 & n28984;
  assign n28986 = ~n28982 & ~n28985;
  assign n28987 = ~n28978 & ~n28985;
  assign n28988 = ~n28982 & n28987;
  assign n28989 = ~n28978 & n28986;
  assign n28990 = pi788 & ~n63982;
  assign n28991 = ~n63981 & ~n28990;
  assign n28992 = pi789 & ~n28968;
  assign n28993 = pi789 & ~n28962;
  assign n28994 = ~n28968 & n28993;
  assign n28995 = ~n28962 & n28992;
  assign n28996 = ~pi789 & n28956;
  assign n28997 = ~n28990 & ~n28996;
  assign n28998 = ~n63983 & n28997;
  assign n28999 = ~n62894 & n63982;
  assign n29000 = ~n63030 & ~n28999;
  assign n29001 = ~n28998 & n29000;
  assign n29002 = ~n63030 & ~n28991;
  assign n29003 = ~n28643 & ~n63984;
  assign n29004 = ~n8651 & ~n29003;
  assign n29005 = ~n8334 & ~n28497;
  assign n29006 = n8334 & ~n28445;
  assign n29007 = ~n8413 & ~n29006;
  assign n29008 = ~n8334 & n28497;
  assign n29009 = n8334 & n28445;
  assign n29010 = ~n29008 & ~n29009;
  assign n29011 = ~n8413 & ~n29010;
  assign n29012 = ~n29005 & n29007;
  assign n29013 = ~n62892 & ~n28632;
  assign n29014 = n62892 & ~n28445;
  assign n29015 = ~n29013 & ~n29014;
  assign n29016 = ~n62892 & n28632;
  assign n29017 = n62892 & n28445;
  assign n29018 = ~n29016 & ~n29017;
  assign n29019 = pi647 & n29018;
  assign n29020 = pi647 & ~n29015;
  assign n29021 = ~pi647 & ~n28445;
  assign n29022 = pi1157 & ~n29021;
  assign n29023 = ~n63986 & n29022;
  assign n29024 = ~pi630 & n29023;
  assign n29025 = ~pi647 & n29018;
  assign n29026 = ~pi647 & ~n29015;
  assign n29027 = pi647 & ~n28445;
  assign n29028 = ~pi1157 & ~n29027;
  assign n29029 = ~n63987 & n29028;
  assign n29030 = pi630 & n29029;
  assign n29031 = ~n29024 & ~n29030;
  assign n29032 = ~n63985 & n29031;
  assign n29033 = pi787 & ~n29032;
  assign n29034 = ~n11547 & ~n29033;
  assign n29035 = ~n29004 & n29034;
  assign n29036 = n8685 & n63793;
  assign n29037 = n28495 & n29036;
  assign n29038 = ~n29023 & ~n29029;
  assign n29039 = pi787 & ~n29038;
  assign n29040 = ~pi787 & ~n29018;
  assign n29041 = ~pi787 & n29015;
  assign n29042 = ~n63036 & ~n63988;
  assign n29043 = ~n29039 & n29042;
  assign n29044 = n28255 & ~n28445;
  assign n29045 = ~n29043 & ~n29044;
  assign n29046 = ~n29037 & n29045;
  assign n29047 = pi790 & ~n29046;
  assign n29048 = n62455 & ~n29047;
  assign n29049 = ~n29035 & n29048;
  assign n29050 = ~n29004 & ~n29033;
  assign n29051 = pi644 & n29050;
  assign n29052 = ~n29039 & ~n63988;
  assign n29053 = ~pi644 & n29052;
  assign n29054 = pi715 & ~n29053;
  assign n29055 = ~n29051 & n29054;
  assign n29056 = ~n11558 & ~n28445;
  assign n29057 = n8685 & n28495;
  assign n29058 = n8376 & ~n28445;
  assign n29059 = ~n8376 & n29010;
  assign n29060 = ~n29058 & ~n29059;
  assign n29061 = ~n29056 & ~n29057;
  assign n29062 = pi644 & ~n63989;
  assign n29063 = ~pi644 & ~n28445;
  assign n29064 = ~pi715 & ~n29063;
  assign n29065 = ~n29062 & n29064;
  assign n29066 = pi1160 & ~n29065;
  assign n29067 = ~n29055 & n29066;
  assign n29068 = ~pi644 & n29050;
  assign n29069 = pi644 & n29052;
  assign n29070 = ~pi715 & ~n29069;
  assign n29071 = ~n29068 & n29070;
  assign n29072 = ~pi644 & ~n63989;
  assign n29073 = pi644 & ~n28445;
  assign n29074 = pi715 & ~n29073;
  assign n29075 = ~n29072 & n29074;
  assign n29076 = ~pi1160 & ~n29075;
  assign n29077 = ~n29071 & n29076;
  assign n29078 = ~n29067 & ~n29077;
  assign n29079 = pi790 & ~n29078;
  assign n29080 = ~pi790 & n29050;
  assign n29081 = ~n29079 & ~n29080;
  assign n29082 = n62455 & ~n29081;
  assign n29083 = ~pi222 & ~n62455;
  assign n29084 = ~n29082 & ~n29083;
  assign n29085 = ~n28299 & ~n29049;
  assign n29086 = ~pi299 & n62785;
  assign n29087 = pi39 & ~n29086;
  assign n29088 = ~n7142 & n29087;
  assign n29089 = ~n6946 & n62952;
  assign n29090 = ~n29088 & n29089;
  assign n29091 = n9733 & ~n29090;
  assign n29092 = pi223 & ~n29091;
  assign n29093 = n16172 & ~n29092;
  assign n29094 = n8135 & ~n29092;
  assign n29095 = pi223 & ~n62765;
  assign n29096 = ~pi223 & pi642;
  assign n29097 = n7285 & n29096;
  assign n29098 = ~pi299 & ~n29097;
  assign n29099 = ~pi642 & n7285;
  assign n29100 = pi223 & ~n29099;
  assign n29101 = n7163 & n29100;
  assign n29102 = n29098 & ~n29101;
  assign n29103 = n7290 & n29096;
  assign n29104 = pi299 & ~n29103;
  assign n29105 = n2902 & n7289;
  assign n29106 = pi223 & ~n29105;
  assign n29107 = pi223 & ~n7169;
  assign n29108 = ~n29105 & n29107;
  assign n29109 = ~n7169 & n29106;
  assign n29110 = n29104 & ~n63991;
  assign n29111 = ~pi39 & ~n29110;
  assign n29112 = ~n29102 & n29111;
  assign n29113 = pi642 & n7187;
  assign n29114 = ~n2903 & n6951;
  assign n29115 = ~n29113 & n29114;
  assign n29116 = pi642 & ~n7188;
  assign n29117 = n2903 & ~n29116;
  assign n29118 = ~n7079 & n29117;
  assign n29119 = ~n29115 & ~n29118;
  assign n29120 = pi681 & n29119;
  assign n29121 = ~n2906 & ~n29119;
  assign n29122 = ~pi642 & n7076;
  assign n29123 = ~n7183 & ~n29122;
  assign n29124 = n2906 & ~n29123;
  assign n29125 = ~pi681 & ~n29124;
  assign n29126 = ~n29121 & n29125;
  assign n29127 = n62393 & ~n29126;
  assign n29128 = ~n29120 & n29127;
  assign n29129 = pi642 & ~n7523;
  assign n29130 = ~pi642 & n62786;
  assign n29131 = ~n29129 & ~n29130;
  assign n29132 = pi681 & ~n29131;
  assign n29133 = ~n2906 & n29131;
  assign n29134 = n7067 & ~n29113;
  assign n29135 = ~pi681 & ~n29134;
  assign n29136 = ~n29133 & n29135;
  assign n29137 = ~n62393 & ~n29136;
  assign n29138 = ~n29132 & n29137;
  assign n29139 = pi223 & ~n29138;
  assign n29140 = ~n29128 & n29139;
  assign n29141 = ~n7057 & n29113;
  assign n29142 = pi681 & ~n29141;
  assign n29143 = ~n2906 & n29141;
  assign n29144 = pi642 & n2906;
  assign n29145 = n7398 & n29144;
  assign n29146 = ~pi681 & ~n29145;
  assign n29147 = ~n29143 & n29146;
  assign n29148 = ~n29142 & ~n29147;
  assign n29149 = ~n2916 & n29148;
  assign n29150 = pi642 & n7298;
  assign n29151 = ~n2906 & n29150;
  assign n29152 = ~pi681 & ~n29151;
  assign n29153 = n7296 & n29144;
  assign n29154 = n29152 & ~n29153;
  assign n29155 = pi681 & ~n29150;
  assign n29156 = ~n29154 & ~n29155;
  assign n29157 = n2916 & n29156;
  assign n29158 = ~pi947 & ~n29157;
  assign n29159 = ~pi947 & ~n29149;
  assign n29160 = ~n29157 & n29159;
  assign n29161 = ~n29149 & n29158;
  assign n29162 = pi947 & ~n29148;
  assign n29163 = ~pi223 & ~n29162;
  assign n29164 = ~n63992 & n29163;
  assign n29165 = ~n7118 & ~n29164;
  assign n29166 = ~n29140 & n29165;
  assign n29167 = pi223 & ~n6951;
  assign n29168 = n7118 & ~n29167;
  assign n29169 = ~n29150 & n29168;
  assign n29170 = ~pi215 & ~n29169;
  assign n29171 = ~n29166 & n29170;
  assign n29172 = n7322 & n29144;
  assign n29173 = n29152 & ~n29172;
  assign n29174 = pi642 & ~n7224;
  assign n29175 = n2906 & ~n29174;
  assign n29176 = ~n6971 & n29175;
  assign n29177 = ~pi681 & ~n29176;
  assign n29178 = n6973 & n29177;
  assign n29179 = ~n29173 & ~n29178;
  assign n29180 = pi642 & n7323;
  assign n29181 = pi681 & ~n29180;
  assign n29182 = n29179 & ~n29181;
  assign n29183 = ~n2916 & n29182;
  assign n29184 = n62393 & ~n29173;
  assign n29185 = n29150 & n29184;
  assign n29186 = ~pi947 & ~n29185;
  assign n29187 = ~n29183 & n29186;
  assign n29188 = pi947 & ~n29182;
  assign n29189 = ~pi223 & ~n29188;
  assign n29190 = ~n29187 & n29189;
  assign n29191 = n28353 & ~n29116;
  assign n29192 = ~n29115 & ~n29191;
  assign n29193 = pi681 & n29192;
  assign n29194 = ~n2906 & ~n29192;
  assign n29195 = n6955 & ~n29113;
  assign n29196 = n2906 & n29195;
  assign n29197 = n6979 & n29196;
  assign n29198 = ~pi681 & ~n29197;
  assign n29199 = ~n29194 & n29198;
  assign n29200 = ~n29193 & ~n29199;
  assign n29201 = n62393 & n29200;
  assign n29202 = ~n6981 & n7186;
  assign n29203 = ~n6973 & ~n29174;
  assign n29204 = ~pi642 & ~n62783;
  assign n29205 = pi642 & ~n7225;
  assign n29206 = ~n29204 & ~n29205;
  assign n29207 = ~n29202 & n29203;
  assign n29208 = ~n2906 & n63993;
  assign n29209 = n29177 & ~n29208;
  assign n29210 = pi681 & ~n63993;
  assign n29211 = ~n29209 & ~n29210;
  assign n29212 = ~n62393 & n29211;
  assign n29213 = pi223 & ~n29212;
  assign n29214 = ~n29201 & n29213;
  assign n29215 = ~n29190 & ~n29214;
  assign n29216 = pi215 & ~n29215;
  assign n29217 = pi299 & ~n29216;
  assign n29218 = ~n29171 & n29217;
  assign n29219 = ~n2971 & n29148;
  assign n29220 = n2971 & n29156;
  assign n29221 = ~n7034 & ~n29220;
  assign n29222 = ~n7034 & ~n29219;
  assign n29223 = ~n29220 & n29222;
  assign n29224 = ~n29219 & n29221;
  assign n29225 = n7034 & ~n29150;
  assign n29226 = ~pi223 & ~n29225;
  assign n29227 = ~n63994 & n29226;
  assign n29228 = n2971 & n29200;
  assign n29229 = ~n2971 & n29211;
  assign n29230 = pi223 & ~n29229;
  assign n29231 = ~n29228 & n29230;
  assign n29232 = ~pi299 & ~n29231;
  assign n29233 = ~n29227 & n29232;
  assign n29234 = pi39 & ~n29233;
  assign n29235 = ~n29218 & n29234;
  assign n29236 = ~pi38 & ~n29235;
  assign n29237 = ~pi38 & ~n29112;
  assign n29238 = ~n29235 & n29237;
  assign n29239 = ~n29112 & n29236;
  assign n29240 = pi39 & pi223;
  assign n29241 = pi38 & ~n29240;
  assign n29242 = ~pi223 & ~n6955;
  assign n29243 = ~pi39 & ~n29242;
  assign n29244 = ~n29195 & n29243;
  assign n29245 = n29241 & ~n29244;
  assign n29246 = n62765 & ~n29245;
  assign n29247 = ~n63995 & n29246;
  assign n29248 = ~n29095 & ~n29247;
  assign n29249 = ~n8135 & n29248;
  assign n29250 = ~n8135 & ~n29248;
  assign n29251 = n8135 & n29092;
  assign n29252 = ~n29250 & ~n29251;
  assign n29253 = ~n29094 & ~n29249;
  assign n29254 = ~pi785 & ~n63996;
  assign n29255 = pi609 & n63996;
  assign n29256 = ~pi609 & ~n29092;
  assign n29257 = pi1155 & ~n29256;
  assign n29258 = ~n29255 & n29257;
  assign n29259 = ~pi609 & n63996;
  assign n29260 = pi609 & ~n29092;
  assign n29261 = ~pi1155 & ~n29260;
  assign n29262 = ~n29259 & n29261;
  assign n29263 = ~n29258 & ~n29262;
  assign n29264 = pi785 & ~n29263;
  assign n29265 = ~n29254 & ~n29264;
  assign n29266 = ~pi781 & ~n29265;
  assign n29267 = pi618 & n29265;
  assign n29268 = ~pi618 & ~n29092;
  assign n29269 = pi1154 & ~n29268;
  assign n29270 = ~n29267 & n29269;
  assign n29271 = ~pi618 & n29265;
  assign n29272 = pi618 & ~n29092;
  assign n29273 = ~pi1154 & ~n29272;
  assign n29274 = ~n29271 & n29273;
  assign n29275 = ~n29270 & ~n29274;
  assign n29276 = pi781 & ~n29275;
  assign n29277 = ~n29266 & ~n29276;
  assign n29278 = pi619 & n29277;
  assign n29279 = ~pi619 & ~n29092;
  assign n29280 = pi1159 & ~n29279;
  assign n29281 = ~n29278 & n29280;
  assign n29282 = ~pi619 & n29277;
  assign n29283 = pi619 & ~n29092;
  assign n29284 = ~pi1159 & ~n29283;
  assign n29285 = ~n29282 & n29284;
  assign n29286 = ~n29282 & ~n29283;
  assign n29287 = ~pi1159 & ~n29286;
  assign n29288 = ~n29278 & ~n29279;
  assign n29289 = pi1159 & ~n29288;
  assign n29290 = ~n29287 & ~n29289;
  assign n29291 = ~n29281 & ~n29285;
  assign n29292 = pi789 & ~n63997;
  assign n29293 = ~pi789 & n29277;
  assign n29294 = ~pi789 & ~n29277;
  assign n29295 = pi789 & n63997;
  assign n29296 = ~n29294 & ~n29295;
  assign n29297 = ~n29292 & ~n29293;
  assign n29298 = ~n8595 & n63998;
  assign n29299 = n8685 & n16177;
  assign n29300 = n11558 & n63998;
  assign n29301 = n16177 & n29300;
  assign n29302 = n29298 & n29299;
  assign n29303 = ~n29093 & ~n63999;
  assign n29304 = pi644 & ~n29303;
  assign n29305 = ~n11558 & ~n25932;
  assign n29306 = ~n29092 & n29305;
  assign n29307 = pi790 & ~n29306;
  assign n29308 = ~n29304 & n29307;
  assign n29309 = n16177 & ~n29092;
  assign n29310 = n8685 & n16172;
  assign n29311 = n16172 & n29300;
  assign n29312 = n29298 & n29310;
  assign n29313 = ~n29309 & ~n64000;
  assign n29314 = ~pi644 & ~n29313;
  assign n29315 = ~n10206 & ~n29092;
  assign n29316 = n62880 & ~n29092;
  assign n29317 = ~pi223 & ~n7849;
  assign n29318 = pi680 & pi681;
  assign n29319 = n7849 & ~n29318;
  assign n29320 = pi223 & n7826;
  assign n29321 = pi299 & ~n29320;
  assign n29322 = ~n29319 & n29321;
  assign n29323 = ~n29317 & n29321;
  assign n29324 = ~n29319 & n29323;
  assign n29325 = ~n29317 & n29322;
  assign n29326 = ~pi223 & ~n7840;
  assign n29327 = n7840 & ~n29318;
  assign n29328 = pi223 & n7820;
  assign n29329 = ~pi299 & ~n29328;
  assign n29330 = ~n29327 & n29329;
  assign n29331 = ~n29326 & n29329;
  assign n29332 = ~n29327 & n29331;
  assign n29333 = ~n29326 & n29330;
  assign n29334 = ~pi39 & ~n64002;
  assign n29335 = ~pi39 & ~n64001;
  assign n29336 = ~n64002 & n29335;
  assign n29337 = ~n64001 & n29334;
  assign n29338 = pi681 & n62828;
  assign n29339 = n7544 & n29318;
  assign n29340 = n29168 & ~n64004;
  assign n29341 = pi681 & ~n7937;
  assign n29342 = n62393 & ~n7103;
  assign n29343 = ~n29341 & n29342;
  assign n29344 = pi681 & ~n28534;
  assign n29345 = ~n62393 & ~n7069;
  assign n29346 = ~n29344 & n29345;
  assign n29347 = pi223 & ~n29346;
  assign n29348 = ~n29343 & n29347;
  assign n29349 = pi681 & n8013;
  assign n29350 = ~n62393 & ~n29349;
  assign n29351 = ~n8018 & n29318;
  assign n29352 = n62393 & ~n29351;
  assign n29353 = ~pi223 & ~n29352;
  assign n29354 = ~pi223 & ~n29350;
  assign n29355 = ~n29352 & n29354;
  assign n29356 = ~n29350 & n29353;
  assign n29357 = ~n7118 & ~n64005;
  assign n29358 = ~n29348 & n29357;
  assign n29359 = ~n29340 & ~n29358;
  assign n29360 = ~pi215 & ~n29359;
  assign n29361 = pi681 & ~n7964;
  assign n29362 = ~n7001 & ~n29361;
  assign n29363 = ~n62393 & n29362;
  assign n29364 = pi681 & ~n7959;
  assign n29365 = ~n7025 & ~n29364;
  assign n29366 = n62393 & n29365;
  assign n29367 = pi223 & ~n29366;
  assign n29368 = ~n29363 & n29367;
  assign n29369 = ~pi223 & pi681;
  assign n29370 = n8052 & n29369;
  assign n29371 = pi215 & ~n29370;
  assign n29372 = ~n29368 & n29371;
  assign n29373 = pi299 & ~n29372;
  assign n29374 = ~n29360 & n29373;
  assign n29375 = n2971 & ~n29351;
  assign n29376 = ~n2971 & ~n29349;
  assign n29377 = ~n7034 & ~n29376;
  assign n29378 = n2971 & n29351;
  assign n29379 = ~n2971 & n29349;
  assign n29380 = ~n29378 & ~n29379;
  assign n29381 = ~n7034 & ~n29380;
  assign n29382 = ~n29375 & n29377;
  assign n29383 = n7034 & n64004;
  assign n29384 = ~pi223 & ~n29383;
  assign n29385 = n7034 & ~n64004;
  assign n29386 = ~n7034 & ~n29379;
  assign n29387 = ~n7034 & ~n29378;
  assign n29388 = ~n29379 & n29387;
  assign n29389 = ~n29378 & n29386;
  assign n29390 = ~n29385 & ~n64007;
  assign n29391 = ~pi223 & ~n29390;
  assign n29392 = ~n64006 & n29384;
  assign n29393 = ~n2971 & ~n29362;
  assign n29394 = n2971 & ~n29365;
  assign n29395 = pi223 & ~n29394;
  assign n29396 = ~n29393 & n29395;
  assign n29397 = ~pi299 & ~n29396;
  assign n29398 = ~n64008 & n29397;
  assign n29399 = pi39 & ~n29398;
  assign n29400 = ~n29374 & n29399;
  assign n29401 = ~n64003 & ~n29400;
  assign n29402 = ~pi38 & ~n29401;
  assign n29403 = pi223 & ~n7357;
  assign n29404 = pi681 & n8084;
  assign n29405 = pi38 & ~n29404;
  assign n29406 = pi38 & ~n29403;
  assign n29407 = ~n29404 & n29406;
  assign n29408 = ~n29403 & n29405;
  assign n29409 = n62765 & ~n64009;
  assign n29410 = ~n29402 & n29409;
  assign n29411 = ~n29095 & ~n29410;
  assign n29412 = ~pi778 & ~n29411;
  assign n29413 = pi625 & n29411;
  assign n29414 = ~pi625 & ~n29092;
  assign n29415 = pi1153 & ~n29414;
  assign n29416 = ~n29413 & n29415;
  assign n29417 = ~pi625 & n29411;
  assign n29418 = pi625 & ~n29092;
  assign n29419 = ~pi1153 & ~n29418;
  assign n29420 = ~n29417 & n29419;
  assign n29421 = ~n29416 & ~n29420;
  assign n29422 = pi778 & ~n29421;
  assign n29423 = ~n29412 & ~n29422;
  assign n29424 = ~n62880 & n29423;
  assign n29425 = ~n62880 & ~n29423;
  assign n29426 = n62880 & n29092;
  assign n29427 = ~n29425 & ~n29426;
  assign n29428 = ~n29316 & ~n29424;
  assign n29429 = ~n62882 & ~n64010;
  assign n29430 = n62882 & n29092;
  assign n29431 = n62882 & ~n29092;
  assign n29432 = ~n62882 & n64010;
  assign n29433 = ~n29431 & ~n29432;
  assign n29434 = ~n29429 & ~n29430;
  assign n29435 = ~n8257 & ~n64011;
  assign n29436 = ~n8303 & n29435;
  assign n29437 = ~n29315 & ~n29436;
  assign n29438 = ~n62892 & ~n29437;
  assign n29439 = n62892 & ~n29092;
  assign n29440 = ~n62892 & n29437;
  assign n29441 = n62892 & n29092;
  assign n29442 = ~n29440 & ~n29441;
  assign n29443 = ~n29438 & ~n29439;
  assign n29444 = pi647 & n64012;
  assign n29445 = ~pi647 & ~n29092;
  assign n29446 = pi1157 & ~n29445;
  assign n29447 = ~n29444 & n29446;
  assign n29448 = ~pi647 & n64012;
  assign n29449 = pi647 & ~n29092;
  assign n29450 = ~pi1157 & ~n29449;
  assign n29451 = ~n29448 & n29450;
  assign n29452 = ~n29447 & ~n29451;
  assign n29453 = pi787 & ~n29452;
  assign n29454 = ~pi787 & ~n64012;
  assign n29455 = ~n63036 & ~n29454;
  assign n29456 = ~n29453 & n29455;
  assign n29457 = ~n29314 & ~n29456;
  assign n29458 = n29307 & ~n29456;
  assign n29459 = ~n29304 & n29458;
  assign n29460 = ~n29314 & n29459;
  assign n29461 = n29308 & n29457;
  assign n29462 = pi790 & ~n64013;
  assign n29463 = n8595 & ~n29092;
  assign n29464 = ~n8595 & ~n63998;
  assign n29465 = n8595 & n29092;
  assign n29466 = ~n29464 & ~n29465;
  assign n29467 = ~n29298 & ~n29463;
  assign n29468 = ~n63052 & ~n64014;
  assign n29469 = ~pi628 & ~n29437;
  assign n29470 = pi628 & ~n29092;
  assign n29471 = n8332 & ~n29470;
  assign n29472 = ~n29469 & n29471;
  assign n29473 = pi628 & ~n29437;
  assign n29474 = ~pi628 & ~n29092;
  assign n29475 = n8331 & ~n29474;
  assign n29476 = ~n29473 & n29475;
  assign n29477 = ~n29472 & ~n29476;
  assign n29478 = ~n29468 & n29477;
  assign n29479 = pi792 & ~n29478;
  assign n29480 = ~pi626 & ~n63998;
  assign n29481 = pi626 & n29092;
  assign n29482 = n8301 & ~n29481;
  assign n29483 = ~n29480 & n29482;
  assign n29484 = n8257 & ~n29092;
  assign n29485 = ~n29435 & ~n29484;
  assign n29486 = n8525 & ~n29485;
  assign n29487 = pi626 & ~n63998;
  assign n29488 = ~pi626 & n29092;
  assign n29489 = n8300 & ~n29488;
  assign n29490 = ~n29487 & n29489;
  assign n29491 = ~n29486 & ~n29490;
  assign n29492 = ~n29483 & ~n29486;
  assign n29493 = ~n29490 & n29492;
  assign n29494 = ~n29483 & n29491;
  assign n29495 = pi788 & ~n64015;
  assign n29496 = n7844 & ~n29318;
  assign n29497 = ~n28846 & n29100;
  assign n29498 = ~n29496 & n29497;
  assign n29499 = n7845 & n29369;
  assign n29500 = n29098 & ~n29499;
  assign n29501 = ~n29498 & n29500;
  assign n29502 = n7853 & n29369;
  assign n29503 = n7852 & ~n29318;
  assign n29504 = ~n28838 & n29106;
  assign n29505 = ~n29503 & n29504;
  assign n29506 = n29104 & ~n29505;
  assign n29507 = n29104 & ~n29502;
  assign n29508 = ~n29505 & n29507;
  assign n29509 = ~n29502 & n29506;
  assign n29510 = ~pi39 & ~n64016;
  assign n29511 = ~pi39 & ~n29501;
  assign n29512 = ~n64016 & n29511;
  assign n29513 = ~n29501 & n29510;
  assign n29514 = ~pi680 & ~n29150;
  assign n29515 = pi642 & ~n7712;
  assign n29516 = ~n7367 & ~n29515;
  assign n29517 = n29114 & ~n29516;
  assign n29518 = pi680 & ~n29517;
  assign n29519 = pi642 & ~n7653;
  assign n29520 = n2903 & ~n29519;
  assign n29521 = ~pi642 & ~n7552;
  assign n29522 = n29520 & ~n29521;
  assign n29523 = n29518 & ~n29522;
  assign n29524 = ~n29514 & ~n29523;
  assign n29525 = pi681 & ~n29524;
  assign n29526 = ~n29154 & ~n29525;
  assign n29527 = n62393 & ~n29526;
  assign n29528 = ~n29142 & ~n29318;
  assign n29529 = ~pi642 & ~n2903;
  assign n29530 = ~n7524 & n29529;
  assign n29531 = pi642 & n7639;
  assign n29532 = pi680 & ~n29531;
  assign n29533 = ~n7643 & n29532;
  assign n29534 = ~n29530 & n29533;
  assign n29535 = ~n29528 & ~n29534;
  assign n29536 = ~n29147 & ~n29535;
  assign n29537 = ~n62393 & ~n29536;
  assign n29538 = ~pi223 & ~n29537;
  assign n29539 = ~pi223 & ~n29527;
  assign n29540 = ~n29537 & n29539;
  assign n29541 = ~n29527 & n29538;
  assign n29542 = ~n29120 & ~n29318;
  assign n29543 = ~pi642 & ~n7367;
  assign n29544 = pi642 & n7652;
  assign n29545 = ~n29543 & ~n29544;
  assign n29546 = pi642 & ~n7652;
  assign n29547 = n13901 & ~n29546;
  assign n29548 = n6955 & ~n29545;
  assign n29549 = ~n6948 & n64019;
  assign n29550 = ~n2903 & ~n29549;
  assign n29551 = pi680 & ~n29550;
  assign n29552 = ~n7373 & ~n29515;
  assign n29553 = n2903 & ~n29552;
  assign n29554 = n29551 & ~n29553;
  assign n29555 = ~n29542 & ~n29554;
  assign n29556 = n29127 & ~n29555;
  assign n29557 = ~n29132 & ~n29318;
  assign n29558 = n28688 & n29529;
  assign n29559 = n7186 & ~n28693;
  assign n29560 = pi642 & ~n63970;
  assign n29561 = pi680 & ~n29560;
  assign n29562 = ~n29559 & n29561;
  assign n29563 = ~n29558 & n29561;
  assign n29564 = ~n29559 & n29563;
  assign n29565 = ~n29558 & n29562;
  assign n29566 = ~n29557 & ~n64020;
  assign n29567 = n29137 & ~n29566;
  assign n29568 = pi223 & ~n29567;
  assign n29569 = ~n29556 & n29568;
  assign n29570 = ~n7118 & ~n29569;
  assign n29571 = ~n29556 & ~n29567;
  assign n29572 = pi223 & ~n29571;
  assign n29573 = n62393 & n29526;
  assign n29574 = ~n62393 & n29536;
  assign n29575 = ~pi223 & ~n29574;
  assign n29576 = ~n29573 & n29575;
  assign n29577 = ~n29572 & ~n29576;
  assign n29578 = ~n7118 & ~n29577;
  assign n29579 = ~n64018 & n29570;
  assign n29580 = n29318 & n64019;
  assign n29581 = n29195 & ~n29318;
  assign n29582 = pi223 & ~n29581;
  assign n29583 = pi223 & ~n29580;
  assign n29584 = ~n29581 & n29583;
  assign n29585 = ~n29580 & n29582;
  assign n29586 = n29113 & ~n29318;
  assign n29587 = n29318 & ~n29543;
  assign n29588 = ~n28891 & n29587;
  assign n29589 = ~n29586 & ~n29588;
  assign n29590 = ~pi223 & ~n29589;
  assign n29591 = n6951 & ~n29589;
  assign n29592 = ~pi223 & n29591;
  assign n29593 = n6951 & n29590;
  assign n29594 = ~n64022 & ~n64023;
  assign n29595 = n29168 & ~n64022;
  assign n29596 = ~n64023 & n29595;
  assign n29597 = n29168 & n29594;
  assign n29598 = ~pi215 & ~n64024;
  assign n29599 = ~n64021 & n29598;
  assign n29600 = ~n29193 & ~n29318;
  assign n29601 = ~pi614 & n7436;
  assign n29602 = ~n29515 & ~n29601;
  assign n29603 = ~pi616 & ~n29602;
  assign n29604 = n29551 & ~n29603;
  assign n29605 = ~n29600 & ~n29604;
  assign n29606 = ~n29199 & ~n29605;
  assign n29607 = n62393 & ~n29606;
  assign n29608 = ~n2903 & n7450;
  assign n29609 = pi642 & ~n28754;
  assign n29610 = pi680 & ~n7452;
  assign n29611 = ~n29609 & n29610;
  assign n29612 = ~n29608 & n29611;
  assign n29613 = ~pi680 & n63993;
  assign n29614 = pi681 & ~n29613;
  assign n29615 = pi681 & ~n29612;
  assign n29616 = ~n29613 & n29615;
  assign n29617 = ~n29612 & n29614;
  assign n29618 = ~n29209 & ~n64025;
  assign n29619 = ~n62393 & ~n29618;
  assign n29620 = pi223 & ~n29619;
  assign n29621 = ~n29607 & n29620;
  assign n29622 = ~n7586 & n29520;
  assign n29623 = n29518 & ~n29622;
  assign n29624 = ~n29514 & ~n29623;
  assign n29625 = pi681 & ~n29624;
  assign n29626 = n29184 & ~n29625;
  assign n29627 = ~n29181 & ~n29318;
  assign n29628 = n7579 & n7690;
  assign n29629 = n7186 & ~n29628;
  assign n29630 = pi642 & n28768;
  assign n29631 = ~n7584 & n29529;
  assign n29632 = pi680 & ~n29631;
  assign n29633 = pi680 & ~n29630;
  assign n29634 = ~n29631 & n29633;
  assign n29635 = ~n29630 & n29632;
  assign n29636 = ~n29629 & n64026;
  assign n29637 = ~n29627 & ~n29636;
  assign n29638 = ~n62393 & n29179;
  assign n29639 = ~n29637 & n29638;
  assign n29640 = ~pi223 & ~n29639;
  assign n29641 = ~pi223 & ~n29626;
  assign n29642 = ~n29639 & n29641;
  assign n29643 = ~n29626 & n29640;
  assign n29644 = pi215 & ~n64027;
  assign n29645 = ~n29621 & n29644;
  assign n29646 = pi299 & ~n29645;
  assign n29647 = ~n29599 & n29646;
  assign n29648 = ~n2971 & n29536;
  assign n29649 = n2971 & n29526;
  assign n29650 = ~n7034 & ~n29649;
  assign n29651 = ~n7034 & ~n29648;
  assign n29652 = ~n29649 & n29651;
  assign n29653 = ~n29648 & n29650;
  assign n29654 = n7034 & ~n29591;
  assign n29655 = ~pi223 & ~n29654;
  assign n29656 = ~n64028 & n29655;
  assign n29657 = n2971 & n29606;
  assign n29658 = ~n2971 & n29618;
  assign n29659 = pi223 & ~n29658;
  assign n29660 = ~n29657 & n29659;
  assign n29661 = ~pi299 & ~n29660;
  assign n29662 = n2971 & ~n29606;
  assign n29663 = ~n2971 & ~n29618;
  assign n29664 = pi223 & ~n29663;
  assign n29665 = ~n29662 & n29664;
  assign n29666 = n2971 & ~n29526;
  assign n29667 = ~n2971 & ~n29536;
  assign n29668 = ~n7034 & ~n29667;
  assign n29669 = ~n29648 & ~n29649;
  assign n29670 = ~n7034 & ~n29669;
  assign n29671 = ~n29666 & n29668;
  assign n29672 = n7034 & n29591;
  assign n29673 = n62790 & ~n29589;
  assign n29674 = ~pi223 & ~n64030;
  assign n29675 = ~n64029 & n29674;
  assign n29676 = ~n29665 & ~n29675;
  assign n29677 = ~pi299 & ~n29676;
  assign n29678 = ~n29656 & n29661;
  assign n29679 = pi39 & ~n64031;
  assign n29680 = ~n29647 & n29679;
  assign n29681 = ~pi38 & ~n29680;
  assign n29682 = ~pi38 & ~n64017;
  assign n29683 = ~n29680 & n29682;
  assign n29684 = ~n64017 & n29681;
  assign n29685 = ~n64022 & n29589;
  assign n29686 = n29243 & ~n29685;
  assign n29687 = n29241 & ~n29686;
  assign n29688 = n62765 & ~n29687;
  assign n29689 = ~n64032 & n29688;
  assign n29690 = ~n29095 & ~n29689;
  assign n29691 = ~pi625 & n29690;
  assign n29692 = pi625 & n29248;
  assign n29693 = ~pi1153 & ~n29692;
  assign n29694 = ~n29691 & n29693;
  assign n29695 = ~pi608 & ~n29694;
  assign n29696 = ~n29416 & n29695;
  assign n29697 = pi625 & n29690;
  assign n29698 = ~pi625 & n29248;
  assign n29699 = pi1153 & ~n29698;
  assign n29700 = ~n29697 & n29699;
  assign n29701 = pi608 & ~n29700;
  assign n29702 = ~n29420 & n29701;
  assign n29703 = ~n29696 & ~n29702;
  assign n29704 = pi778 & ~n29703;
  assign n29705 = ~pi778 & n29690;
  assign n29706 = ~n29704 & ~n29705;
  assign n29707 = ~pi609 & ~n29706;
  assign n29708 = pi609 & n29423;
  assign n29709 = ~pi1155 & ~n29708;
  assign n29710 = ~n29707 & n29709;
  assign n29711 = ~pi660 & ~n29258;
  assign n29712 = ~n29710 & n29711;
  assign n29713 = pi609 & ~n29706;
  assign n29714 = ~pi609 & n29423;
  assign n29715 = pi1155 & ~n29714;
  assign n29716 = ~n29713 & n29715;
  assign n29717 = pi660 & ~n29262;
  assign n29718 = ~n29716 & n29717;
  assign n29719 = ~n29712 & ~n29718;
  assign n29720 = pi785 & ~n29719;
  assign n29721 = ~pi785 & ~n29706;
  assign n29722 = ~n29720 & ~n29721;
  assign n29723 = pi618 & ~n29722;
  assign n29724 = ~pi618 & n64010;
  assign n29725 = pi1154 & ~n29724;
  assign n29726 = ~n29723 & n29725;
  assign n29727 = pi627 & ~n29274;
  assign n29728 = ~n29726 & n29727;
  assign n29729 = ~pi618 & ~n29722;
  assign n29730 = pi618 & n64010;
  assign n29731 = ~pi1154 & ~n29730;
  assign n29732 = ~n29729 & n29731;
  assign n29733 = ~pi627 & ~n29270;
  assign n29734 = ~n29732 & n29733;
  assign n29735 = pi781 & ~n29734;
  assign n29736 = ~n29728 & n29735;
  assign n29737 = ~n11431 & n64011;
  assign n29738 = ~n62884 & n63997;
  assign n29739 = ~n29737 & ~n29738;
  assign n29740 = pi789 & ~n29739;
  assign n29741 = ~pi781 & n29722;
  assign n29742 = ~n29740 & ~n29741;
  assign n29743 = ~n29736 & n29742;
  assign n29744 = n11434 & n29739;
  assign n29745 = ~n29743 & ~n29744;
  assign n29746 = ~n29728 & ~n29734;
  assign n29747 = pi781 & ~n29746;
  assign n29748 = ~pi781 & ~n29722;
  assign n29749 = ~n29747 & ~n29748;
  assign n29750 = ~pi619 & ~n29749;
  assign n29751 = pi619 & ~n64011;
  assign n29752 = ~pi1159 & ~n29751;
  assign n29753 = ~n29750 & n29752;
  assign n29754 = ~pi648 & ~n29281;
  assign n29755 = ~n29753 & n29754;
  assign n29756 = pi619 & ~n29749;
  assign n29757 = ~pi619 & ~n64011;
  assign n29758 = pi1159 & ~n29757;
  assign n29759 = ~n29756 & n29758;
  assign n29760 = pi648 & ~n29285;
  assign n29761 = ~n29759 & n29760;
  assign n29762 = pi789 & ~n29761;
  assign n29763 = pi789 & ~n29755;
  assign n29764 = ~n29761 & n29763;
  assign n29765 = ~n29755 & n29762;
  assign n29766 = ~pi789 & n29749;
  assign n29767 = n62894 & ~n29766;
  assign n29768 = ~n64033 & n29767;
  assign n29769 = n62894 & ~n29745;
  assign n29770 = ~n29495 & ~n64034;
  assign n29771 = ~n29479 & ~n29770;
  assign n29772 = n63030 & n29478;
  assign n29773 = ~n8651 & ~n29772;
  assign n29774 = ~n29771 & n29773;
  assign n29775 = n63035 & n64013;
  assign n29776 = ~n8334 & n64014;
  assign n29777 = n8334 & ~n29092;
  assign n29778 = ~n8413 & ~n29777;
  assign n29779 = ~n8334 & ~n64014;
  assign n29780 = n8334 & n29092;
  assign n29781 = ~n29779 & ~n29780;
  assign n29782 = ~n8413 & ~n29781;
  assign n29783 = ~n29776 & n29778;
  assign n29784 = ~pi630 & n29447;
  assign n29785 = pi630 & n29451;
  assign n29786 = ~n29784 & ~n29785;
  assign n29787 = ~n64035 & n29786;
  assign n29788 = pi787 & ~n29787;
  assign n29789 = ~n29775 & ~n29788;
  assign n29790 = ~n29774 & n29789;
  assign n29791 = ~n29774 & ~n29788;
  assign n29792 = ~n63035 & n29791;
  assign n29793 = n64013 & ~n29792;
  assign n29794 = ~pi790 & ~n29791;
  assign n29795 = ~n29793 & ~n29794;
  assign n29796 = pi644 & n29791;
  assign n29797 = ~n29453 & ~n29454;
  assign n29798 = ~pi644 & n29797;
  assign n29799 = pi715 & ~n29798;
  assign n29800 = ~n29796 & n29799;
  assign n29801 = n8376 & ~n29092;
  assign n29802 = ~n8376 & n29781;
  assign n29803 = ~n29801 & ~n29802;
  assign n29804 = pi644 & ~n29803;
  assign n29805 = ~pi644 & ~n29092;
  assign n29806 = ~pi715 & ~n29805;
  assign n29807 = ~n29804 & n29806;
  assign n29808 = pi1160 & ~n29807;
  assign n29809 = ~n29800 & n29808;
  assign n29810 = ~pi644 & n29791;
  assign n29811 = pi644 & n29797;
  assign n29812 = ~pi715 & ~n29811;
  assign n29813 = ~n29810 & n29812;
  assign n29814 = ~pi644 & ~n29803;
  assign n29815 = pi644 & ~n29092;
  assign n29816 = pi715 & ~n29815;
  assign n29817 = ~n29814 & n29816;
  assign n29818 = ~pi1160 & ~n29817;
  assign n29819 = ~n29813 & n29818;
  assign n29820 = ~n29809 & ~n29819;
  assign n29821 = pi790 & ~n29820;
  assign n29822 = ~pi790 & n29791;
  assign n29823 = ~n29821 & ~n29822;
  assign n29824 = ~n29462 & ~n29790;
  assign n29825 = n62455 & n64036;
  assign n29826 = ~pi223 & ~n62455;
  assign n29827 = n62455 & ~n64036;
  assign n29828 = pi223 & ~n62455;
  assign n29829 = ~n29827 & ~n29828;
  assign n29830 = ~n29825 & ~n29826;
  assign n29831 = pi224 & ~n28444;
  assign n29832 = n16177 & ~n29831;
  assign n29833 = pi224 & ~n62765;
  assign n29834 = pi614 & n7187;
  assign n29835 = n6951 & ~n29834;
  assign n29836 = ~n2904 & ~n29835;
  assign n29837 = ~n7083 & ~n29836;
  assign n29838 = ~n7008 & ~n29837;
  assign n29839 = ~pi680 & ~n29837;
  assign n29840 = pi680 & n29834;
  assign n29841 = ~n7095 & ~n29840;
  assign n29842 = ~n29839 & n29841;
  assign n29843 = n7008 & ~n29842;
  assign n29844 = ~n29838 & ~n29843;
  assign n29845 = n62393 & n29844;
  assign n29846 = ~n2814 & n7080;
  assign n29847 = n2903 & ~n7056;
  assign n29848 = ~n29846 & n29847;
  assign n29849 = pi614 & ~n7523;
  assign n29850 = ~pi614 & pi616;
  assign n29851 = n7057 & n29850;
  assign n29852 = ~n29849 & ~n29851;
  assign n29853 = ~n2814 & n7089;
  assign n29854 = ~pi614 & ~n7056;
  assign n29855 = ~n29853 & n29854;
  assign n29856 = ~n29849 & ~n29855;
  assign n29857 = ~n29848 & n29852;
  assign n29858 = ~n7008 & ~n64038;
  assign n29859 = ~pi680 & ~n64038;
  assign n29860 = pi614 & n7398;
  assign n29861 = pi680 & ~n29860;
  assign n29862 = n7055 & n29861;
  assign n29863 = ~n29840 & ~n29862;
  assign n29864 = ~n29859 & n29863;
  assign n29865 = n7008 & ~n29864;
  assign n29866 = ~n29858 & ~n29865;
  assign n29867 = ~n62393 & n29866;
  assign n29868 = pi224 & ~n29867;
  assign n29869 = pi224 & ~n29845;
  assign n29870 = ~n29867 & n29869;
  assign n29871 = ~n29845 & n29868;
  assign n29872 = ~n7057 & n29834;
  assign n29873 = ~pi680 & ~n29872;
  assign n29874 = ~n29861 & ~n29873;
  assign n29875 = n7008 & ~n29874;
  assign n29876 = ~n7008 & ~n29872;
  assign n29877 = ~n29875 & ~n29876;
  assign n29878 = ~n62393 & ~n29877;
  assign n29879 = pi614 & ~n63944;
  assign n29880 = n62393 & ~n29879;
  assign n29881 = ~pi224 & ~n29880;
  assign n29882 = ~n29878 & n29881;
  assign n29883 = ~n7118 & ~n29882;
  assign n29884 = ~n64039 & n29883;
  assign n29885 = n7099 & n7187;
  assign n29886 = pi224 & ~n6951;
  assign n29887 = n7118 & ~n29886;
  assign n29888 = ~n29885 & n29887;
  assign n29889 = ~pi215 & ~n29888;
  assign n29890 = ~n29884 & n29889;
  assign n29891 = pi614 & ~n28377;
  assign n29892 = ~n63947 & n29885;
  assign n29893 = ~pi224 & n64040;
  assign n29894 = ~n7328 & n29893;
  assign n29895 = ~n6991 & ~n29836;
  assign n29896 = ~n7008 & ~n29895;
  assign n29897 = ~pi680 & ~n29895;
  assign n29898 = ~n7012 & ~n29840;
  assign n29899 = ~n29897 & n29898;
  assign n29900 = n7008 & ~n29899;
  assign n29901 = ~n29896 & ~n29900;
  assign n29902 = n62393 & n29901;
  assign n29903 = pi614 & ~n7225;
  assign n29904 = ~n7591 & ~n27562;
  assign n29905 = ~n62783 & ~n7591;
  assign n29906 = ~n27561 & n29904;
  assign n29907 = ~n29903 & ~n64041;
  assign n29908 = ~pi680 & ~n29907;
  assign n29909 = ~pi614 & ~n6971;
  assign n29910 = n7230 & ~n29909;
  assign n29911 = ~n29908 & ~n29910;
  assign n29912 = n7008 & ~n29911;
  assign n29913 = ~n7008 & ~n29907;
  assign n29914 = ~n29912 & ~n29913;
  assign n29915 = ~n62393 & n29914;
  assign n29916 = pi224 & ~n29915;
  assign n29917 = ~n29902 & n29916;
  assign n29918 = ~n29894 & ~n29917;
  assign n29919 = pi215 & ~n29918;
  assign n29920 = pi299 & ~n29919;
  assign n29921 = ~n29890 & n29920;
  assign n29922 = n2971 & n29901;
  assign n29923 = ~n2971 & n29914;
  assign n29924 = pi224 & ~n29923;
  assign n29925 = ~n29922 & n29924;
  assign n29926 = ~n7344 & n29893;
  assign n29927 = pi223 & ~n29926;
  assign n29928 = ~n29925 & n29927;
  assign n29929 = n2971 & n29844;
  assign n29930 = ~n2971 & n29866;
  assign n29931 = pi224 & ~n29930;
  assign n29932 = pi224 & ~n29929;
  assign n29933 = ~n29930 & n29932;
  assign n29934 = ~n29929 & n29931;
  assign n29935 = ~n2971 & ~n29877;
  assign n29936 = n2971 & ~n29879;
  assign n29937 = n2978 & ~n29936;
  assign n29938 = ~n29935 & n29937;
  assign n29939 = n7034 & n29885;
  assign n29940 = pi614 & n62807;
  assign n29941 = ~pi223 & ~n64043;
  assign n29942 = ~n29938 & n29941;
  assign n29943 = ~n64042 & n29942;
  assign n29944 = ~n29928 & ~n29943;
  assign n29945 = ~pi299 & ~n29944;
  assign n29946 = pi39 & ~n29945;
  assign n29947 = pi39 & ~n29921;
  assign n29948 = ~n29945 & n29947;
  assign n29949 = ~n29921 & n29946;
  assign n29950 = ~pi614 & n7285;
  assign n29951 = pi224 & ~n29950;
  assign n29952 = n7163 & n29951;
  assign n29953 = pi614 & n7285;
  assign n29954 = ~pi224 & n29953;
  assign n29955 = ~pi299 & ~n29954;
  assign n29956 = ~n29952 & n29955;
  assign n29957 = pi614 & n7290;
  assign n29958 = pi224 & ~n6936;
  assign n29959 = ~n29957 & ~n29958;
  assign n29960 = pi299 & n29959;
  assign n29961 = ~pi39 & ~n29960;
  assign n29962 = ~pi39 & ~n29956;
  assign n29963 = ~n29960 & n29962;
  assign n29964 = ~n29956 & n29961;
  assign n29965 = ~pi38 & ~n64045;
  assign n29966 = ~n64044 & n29965;
  assign n29967 = pi224 & ~n7357;
  assign n29968 = pi38 & ~n29967;
  assign n29969 = pi614 & n7359;
  assign n29970 = n7357 & n29834;
  assign n29971 = n29968 & ~n64046;
  assign n29972 = n62765 & ~n29971;
  assign n29973 = ~n29966 & n29972;
  assign n29974 = ~n29833 & ~n29973;
  assign n29975 = ~n8135 & ~n29974;
  assign n29976 = n8135 & n29831;
  assign n29977 = n8135 & ~n29831;
  assign n29978 = ~n8135 & n29974;
  assign n29979 = ~n29977 & ~n29978;
  assign n29980 = ~n29975 & ~n29976;
  assign n29981 = ~pi785 & n64047;
  assign n29982 = pi609 & ~n64047;
  assign n29983 = ~pi609 & ~n29831;
  assign n29984 = pi1155 & ~n29983;
  assign n29985 = ~n29982 & n29984;
  assign n29986 = ~pi609 & ~n64047;
  assign n29987 = pi609 & ~n29831;
  assign n29988 = ~pi1155 & ~n29987;
  assign n29989 = ~n29986 & n29988;
  assign n29990 = ~n29985 & ~n29989;
  assign n29991 = pi785 & ~n29990;
  assign n29992 = ~n29981 & ~n29991;
  assign n29993 = ~pi781 & ~n29992;
  assign n29994 = pi618 & n29992;
  assign n29995 = ~pi618 & ~n29831;
  assign n29996 = pi1154 & ~n29995;
  assign n29997 = ~n29994 & n29996;
  assign n29998 = ~pi618 & n29992;
  assign n29999 = pi618 & ~n29831;
  assign n30000 = ~pi1154 & ~n29999;
  assign n30001 = ~n29998 & n30000;
  assign n30002 = ~n29997 & ~n30001;
  assign n30003 = pi781 & ~n30002;
  assign n30004 = ~n29993 & ~n30003;
  assign n30005 = pi619 & n30004;
  assign n30006 = ~pi619 & ~n29831;
  assign n30007 = pi1159 & ~n30006;
  assign n30008 = ~n30005 & n30007;
  assign n30009 = ~pi619 & n30004;
  assign n30010 = pi619 & ~n29831;
  assign n30011 = ~pi1159 & ~n30010;
  assign n30012 = ~n30009 & n30011;
  assign n30013 = ~n30009 & ~n30010;
  assign n30014 = ~pi1159 & ~n30013;
  assign n30015 = ~n30005 & ~n30006;
  assign n30016 = pi1159 & ~n30015;
  assign n30017 = ~n30014 & ~n30016;
  assign n30018 = ~n30008 & ~n30012;
  assign n30019 = pi789 & ~n64048;
  assign n30020 = ~pi789 & n30004;
  assign n30021 = ~pi789 & ~n30004;
  assign n30022 = pi789 & n64048;
  assign n30023 = ~n30021 & ~n30022;
  assign n30024 = ~n30019 & ~n30020;
  assign n30025 = ~n8595 & n64049;
  assign n30026 = n8685 & n30025;
  assign n30027 = n16172 & n30026;
  assign n30028 = ~n29832 & ~n30027;
  assign n30029 = ~pi644 & ~n30028;
  assign n30030 = n16172 & ~n29831;
  assign n30031 = n16177 & n30026;
  assign n30032 = ~n30030 & ~n30031;
  assign n30033 = pi644 & ~n30032;
  assign n30034 = n29305 & ~n29831;
  assign n30035 = ~n10206 & ~n29831;
  assign n30036 = ~pi224 & ~n7849;
  assign n30037 = pi662 & pi680;
  assign n30038 = n7849 & ~n30037;
  assign n30039 = pi224 & n7826;
  assign n30040 = pi299 & ~n30039;
  assign n30041 = ~n30038 & n30040;
  assign n30042 = ~n30036 & n30040;
  assign n30043 = ~n30038 & n30042;
  assign n30044 = ~n30036 & n30041;
  assign n30045 = ~pi224 & ~n7840;
  assign n30046 = n7840 & ~n30037;
  assign n30047 = pi224 & n7820;
  assign n30048 = ~pi299 & ~n30047;
  assign n30049 = ~n30046 & n30048;
  assign n30050 = ~n30045 & n30048;
  assign n30051 = ~n30046 & n30050;
  assign n30052 = ~n30045 & n30049;
  assign n30053 = ~pi39 & ~n64051;
  assign n30054 = ~pi39 & ~n64050;
  assign n30055 = ~n64051 & n30054;
  assign n30056 = ~n64050 & n30053;
  assign n30057 = pi662 & n62828;
  assign n30058 = n7544 & n30037;
  assign n30059 = n29887 & ~n64053;
  assign n30060 = pi662 & ~n7937;
  assign n30061 = ~pi662 & ~n7104;
  assign n30062 = ~n30060 & ~n30061;
  assign n30063 = n62393 & n30062;
  assign n30064 = ~n2905 & ~n28534;
  assign n30065 = n62787 & ~n30064;
  assign n30066 = ~n62393 & n30065;
  assign n30067 = pi224 & ~n30066;
  assign n30068 = ~n30063 & n30067;
  assign n30069 = ~n8018 & n30037;
  assign n30070 = n62393 & ~n30069;
  assign n30071 = pi662 & n8013;
  assign n30072 = ~n62393 & ~n30071;
  assign n30073 = ~pi224 & ~n30072;
  assign n30074 = ~pi224 & ~n30070;
  assign n30075 = ~n30072 & n30074;
  assign n30076 = ~n30070 & n30073;
  assign n30077 = ~n7118 & ~n64054;
  assign n30078 = ~n30068 & n30077;
  assign n30079 = ~n30059 & ~n30078;
  assign n30080 = ~pi215 & ~n30079;
  assign n30081 = ~pi662 & ~n7002;
  assign n30082 = pi662 & ~n7964;
  assign n30083 = ~n30081 & ~n30082;
  assign n30084 = ~n62393 & n30083;
  assign n30085 = ~pi662 & ~n62784;
  assign n30086 = pi662 & ~n7959;
  assign n30087 = ~n30085 & ~n30086;
  assign n30088 = n62393 & n30087;
  assign n30089 = pi224 & ~n30088;
  assign n30090 = ~n30084 & n30089;
  assign n30091 = ~pi224 & pi662;
  assign n30092 = n8052 & n30091;
  assign n30093 = pi215 & ~n30092;
  assign n30094 = ~n30090 & n30093;
  assign n30095 = pi299 & ~n30094;
  assign n30096 = ~n30080 & n30095;
  assign n30097 = n2971 & n30062;
  assign n30098 = ~n2971 & n30065;
  assign n30099 = pi224 & ~n30098;
  assign n30100 = ~n30097 & n30099;
  assign n30101 = n2971 & ~n30069;
  assign n30102 = ~n2971 & ~n30071;
  assign n30103 = n2978 & ~n30102;
  assign n30104 = n2978 & ~n30101;
  assign n30105 = ~n30102 & n30104;
  assign n30106 = ~n30101 & n30103;
  assign n30107 = pi662 & n8012;
  assign n30108 = ~pi223 & ~n30107;
  assign n30109 = ~n64055 & n30108;
  assign n30110 = ~n30100 & n30109;
  assign n30111 = ~n2971 & n30083;
  assign n30112 = n2971 & n30087;
  assign n30113 = pi224 & ~n30112;
  assign n30114 = ~n30111 & n30113;
  assign n30115 = n8031 & n30091;
  assign n30116 = pi223 & ~n30115;
  assign n30117 = ~n30114 & n30116;
  assign n30118 = ~pi299 & ~n30117;
  assign n30119 = ~n30110 & n30118;
  assign n30120 = pi39 & ~n30119;
  assign n30121 = ~n30096 & n30120;
  assign n30122 = ~n64052 & ~n30121;
  assign n30123 = ~pi38 & ~n30122;
  assign n30124 = pi662 & n8084;
  assign n30125 = n29968 & ~n30124;
  assign n30126 = n62765 & ~n30125;
  assign n30127 = ~n30123 & n30126;
  assign n30128 = ~n29833 & ~n30127;
  assign n30129 = ~pi778 & ~n30128;
  assign n30130 = pi625 & n30128;
  assign n30131 = ~pi625 & ~n29831;
  assign n30132 = pi1153 & ~n30131;
  assign n30133 = ~n30130 & n30132;
  assign n30134 = ~pi625 & n30128;
  assign n30135 = pi625 & ~n29831;
  assign n30136 = ~pi1153 & ~n30135;
  assign n30137 = ~n30134 & n30136;
  assign n30138 = ~n30133 & ~n30137;
  assign n30139 = pi778 & ~n30138;
  assign n30140 = ~n30129 & ~n30139;
  assign n30141 = ~n62880 & ~n30140;
  assign n30142 = n62880 & n29831;
  assign n30143 = n62880 & ~n29831;
  assign n30144 = ~n62880 & n30140;
  assign n30145 = ~n30143 & ~n30144;
  assign n30146 = ~n30141 & ~n30142;
  assign n30147 = ~n62882 & n64056;
  assign n30148 = n62882 & n29831;
  assign n30149 = ~n62882 & ~n64056;
  assign n30150 = n62882 & ~n29831;
  assign n30151 = ~n30149 & ~n30150;
  assign n30152 = ~n30147 & ~n30148;
  assign n30153 = ~n8257 & ~n64057;
  assign n30154 = ~n8303 & n30153;
  assign n30155 = ~n30035 & ~n30154;
  assign n30156 = ~n62892 & ~n30155;
  assign n30157 = n62892 & ~n29831;
  assign n30158 = ~n62892 & n30155;
  assign n30159 = n62892 & n29831;
  assign n30160 = ~n30158 & ~n30159;
  assign n30161 = ~n30156 & ~n30157;
  assign n30162 = pi647 & n64058;
  assign n30163 = ~pi647 & ~n29831;
  assign n30164 = pi1157 & ~n30163;
  assign n30165 = ~n30162 & n30164;
  assign n30166 = ~pi647 & n64058;
  assign n30167 = pi647 & ~n29831;
  assign n30168 = ~pi1157 & ~n30167;
  assign n30169 = ~n30166 & n30168;
  assign n30170 = ~n30165 & ~n30169;
  assign n30171 = pi787 & ~n30170;
  assign n30172 = ~pi787 & ~n64058;
  assign n30173 = ~n63036 & ~n30172;
  assign n30174 = ~n30171 & n30173;
  assign n30175 = ~n30034 & ~n30174;
  assign n30176 = ~n30033 & n30175;
  assign n30177 = ~n30029 & n30176;
  assign n30178 = pi790 & ~n30177;
  assign n30179 = n8595 & ~n29831;
  assign n30180 = ~n30025 & ~n30179;
  assign n30181 = ~n63052 & n30180;
  assign n30182 = ~n8500 & n29831;
  assign n30183 = n8500 & n30155;
  assign n30184 = ~n30182 & ~n30183;
  assign n30185 = ~pi628 & ~n30155;
  assign n30186 = pi628 & ~n29831;
  assign n30187 = n8332 & ~n30186;
  assign n30188 = ~n30185 & n30187;
  assign n30189 = pi628 & ~n30155;
  assign n30190 = ~pi628 & ~n29831;
  assign n30191 = n8331 & ~n30190;
  assign n30192 = ~n30189 & n30191;
  assign n30193 = ~n30188 & ~n30192;
  assign n30194 = ~n8333 & ~n30184;
  assign n30195 = ~n30181 & n64059;
  assign n30196 = pi792 & ~n30195;
  assign n30197 = ~pi614 & ~n13901;
  assign n30198 = pi614 & ~n28891;
  assign n30199 = ~n30197 & ~n30198;
  assign n30200 = ~n6948 & n30199;
  assign n30201 = pi616 & ~n30200;
  assign n30202 = pi614 & ~n7712;
  assign n30203 = ~n7375 & ~n30202;
  assign n30204 = ~pi616 & ~n30203;
  assign n30205 = ~n30201 & ~n30204;
  assign n30206 = pi680 & ~n30205;
  assign n30207 = ~n29839 & ~n30206;
  assign n30208 = pi662 & ~n30207;
  assign n30209 = ~pi662 & ~n7007;
  assign n30210 = ~n29837 & n30209;
  assign n30211 = ~n29843 & ~n30210;
  assign n30212 = ~n30208 & n30211;
  assign n30213 = pi224 & ~n30212;
  assign n30214 = pi662 & ~n29885;
  assign n30215 = ~n28664 & n30214;
  assign n30216 = ~n62826 & n29850;
  assign n30217 = ~n28663 & ~n30216;
  assign n30218 = n30037 & ~n30217;
  assign n30219 = ~pi662 & ~n29879;
  assign n30220 = ~n30218 & ~n30219;
  assign n30221 = pi680 & ~n30217;
  assign n30222 = ~n28664 & ~n29885;
  assign n30223 = ~n30221 & ~n30222;
  assign n30224 = pi662 & ~n30223;
  assign n30225 = ~n30219 & ~n30224;
  assign n30226 = ~n30215 & n30220;
  assign n30227 = ~pi224 & n64060;
  assign n30228 = n62393 & ~n30227;
  assign n30229 = ~n30213 & n30228;
  assign n30230 = pi614 & ~n63970;
  assign n30231 = n28688 & n29850;
  assign n30232 = ~n30230 & ~n30231;
  assign n30233 = ~n63969 & n30232;
  assign n30234 = pi680 & ~n30233;
  assign n30235 = ~n29859 & ~n30234;
  assign n30236 = pi662 & ~n30235;
  assign n30237 = ~n64038 & n30209;
  assign n30238 = ~n29865 & ~n30237;
  assign n30239 = ~n30236 & n30238;
  assign n30240 = pi224 & ~n30239;
  assign n30241 = ~pi614 & n7537;
  assign n30242 = pi614 & ~n7639;
  assign n30243 = pi680 & ~n30242;
  assign n30244 = ~n30241 & n30243;
  assign n30245 = ~n29873 & ~n30244;
  assign n30246 = pi662 & ~n30245;
  assign n30247 = ~n29872 & n30209;
  assign n30248 = ~n29875 & ~n30247;
  assign n30249 = ~n30246 & n30248;
  assign n30250 = ~pi224 & n30249;
  assign n30251 = ~n62393 & ~n30250;
  assign n30252 = ~n30240 & n30251;
  assign n30253 = ~n30229 & ~n30252;
  assign n30254 = ~pi224 & ~n30249;
  assign n30255 = pi224 & n30239;
  assign n30256 = ~n62393 & ~n30255;
  assign n30257 = ~n62393 & ~n30254;
  assign n30258 = ~n30255 & n30257;
  assign n30259 = ~n30254 & n30256;
  assign n30260 = pi224 & n30212;
  assign n30261 = ~pi224 & ~n64060;
  assign n30262 = n62393 & ~n30261;
  assign n30263 = ~n30260 & n30262;
  assign n30264 = ~n7118 & ~n30263;
  assign n30265 = ~n64061 & n30264;
  assign n30266 = ~n7118 & ~n64061;
  assign n30267 = ~n30263 & n30266;
  assign n30268 = ~n7118 & ~n30253;
  assign n30269 = n62826 & n30037;
  assign n30270 = ~n29885 & ~n30269;
  assign n30271 = ~pi224 & ~n30270;
  assign n30272 = n30037 & n30199;
  assign n30273 = ~n29834 & ~n30037;
  assign n30274 = n6955 & n30273;
  assign n30275 = pi224 & ~n30274;
  assign n30276 = ~n30272 & n30275;
  assign n30277 = n29887 & ~n30276;
  assign n30278 = ~n30271 & n30277;
  assign n30279 = ~pi215 & ~n30278;
  assign n30280 = ~n64062 & n30279;
  assign n30281 = pi680 & ~n7577;
  assign n30282 = ~n29885 & ~n30281;
  assign n30283 = ~pi662 & ~n64040;
  assign n30284 = ~n30218 & ~n30283;
  assign n30285 = ~n30221 & ~n30282;
  assign n30286 = pi662 & ~n30285;
  assign n30287 = ~n30283 & ~n30286;
  assign n30288 = ~n30282 & n30284;
  assign n30289 = ~pi224 & ~n64063;
  assign n30290 = ~n7438 & ~n30202;
  assign n30291 = ~pi616 & ~n30290;
  assign n30292 = ~n30201 & ~n30291;
  assign n30293 = pi680 & ~n30292;
  assign n30294 = ~n29897 & ~n30293;
  assign n30295 = pi662 & ~n30294;
  assign n30296 = ~n29895 & n30209;
  assign n30297 = pi224 & ~n30296;
  assign n30298 = ~n29900 & n30297;
  assign n30299 = ~n29900 & ~n30296;
  assign n30300 = ~n30295 & n30299;
  assign n30301 = pi224 & n30300;
  assign n30302 = ~n30295 & n30298;
  assign n30303 = ~n30289 & ~n64064;
  assign n30304 = n62393 & ~n30303;
  assign n30305 = pi614 & ~n28754;
  assign n30306 = n7453 & ~n30305;
  assign n30307 = pi680 & ~n30306;
  assign n30308 = ~n29908 & ~n30307;
  assign n30309 = pi662 & ~n30308;
  assign n30310 = ~n29907 & n30209;
  assign n30311 = pi224 & ~n30310;
  assign n30312 = ~n29912 & n30311;
  assign n30313 = ~n29912 & ~n30310;
  assign n30314 = ~n30309 & n30313;
  assign n30315 = pi224 & n30314;
  assign n30316 = ~n30309 & n30312;
  assign n30317 = pi614 & ~n28768;
  assign n30318 = ~pi616 & n7586;
  assign n30319 = ~pi614 & n7584;
  assign n30320 = ~n30318 & n30319;
  assign n30321 = ~n30317 & ~n30320;
  assign n30322 = pi614 & n7323;
  assign n30323 = ~n6973 & n29885;
  assign n30324 = ~pi680 & ~n64066;
  assign n30325 = pi662 & ~n30324;
  assign n30326 = ~n30321 & n30325;
  assign n30327 = ~pi662 & ~n6973;
  assign n30328 = n64040 & n30327;
  assign n30329 = ~pi224 & ~n30328;
  assign n30330 = ~n6973 & n64040;
  assign n30331 = ~pi662 & n6973;
  assign n30332 = ~n30283 & ~n30331;
  assign n30333 = ~pi662 & ~n30330;
  assign n30334 = ~pi614 & n7597;
  assign n30335 = pi614 & n28768;
  assign n30336 = pi680 & ~n30335;
  assign n30337 = ~n30334 & n30336;
  assign n30338 = ~n7594 & n30337;
  assign n30339 = pi614 & ~pi680;
  assign n30340 = n7323 & n30339;
  assign n30341 = pi662 & ~n30340;
  assign n30342 = n7584 & ~n30318;
  assign n30343 = ~pi614 & ~n30342;
  assign n30344 = ~n30324 & ~n30335;
  assign n30345 = ~n30343 & n30344;
  assign n30346 = pi662 & ~n30345;
  assign n30347 = ~n30338 & n30341;
  assign n30348 = n64067 & ~n64068;
  assign n30349 = ~pi224 & ~n30348;
  assign n30350 = ~n30326 & n30329;
  assign n30351 = ~n64065 & ~n64069;
  assign n30352 = ~n62393 & ~n30351;
  assign n30353 = pi215 & ~n30352;
  assign n30354 = n62393 & ~n30300;
  assign n30355 = ~n62393 & ~n30314;
  assign n30356 = pi224 & ~n30355;
  assign n30357 = ~n30354 & n30356;
  assign n30358 = n62393 & n64063;
  assign n30359 = ~n62393 & n30348;
  assign n30360 = ~pi224 & ~n30359;
  assign n30361 = ~n30358 & n30360;
  assign n30362 = pi215 & ~n30361;
  assign n30363 = ~n30357 & n30362;
  assign n30364 = ~n30304 & n30353;
  assign n30365 = pi299 & ~n64070;
  assign n30366 = ~n30280 & n30365;
  assign n30367 = n2971 & ~n30289;
  assign n30368 = n2971 & n30303;
  assign n30369 = ~n64064 & n30367;
  assign n30370 = ~n2971 & ~n64069;
  assign n30371 = ~n2971 & n30351;
  assign n30372 = ~n64065 & n30370;
  assign n30373 = pi223 & ~n64072;
  assign n30374 = ~n64071 & n30373;
  assign n30375 = n2971 & ~n64060;
  assign n30376 = n2978 & ~n30375;
  assign n30377 = ~n2971 & ~n30249;
  assign n30378 = n30376 & ~n30377;
  assign n30379 = n30249 & n30376;
  assign n30380 = ~pi222 & n30271;
  assign n30381 = ~pi223 & ~n30380;
  assign n30382 = ~n64073 & n30381;
  assign n30383 = n2971 & n30212;
  assign n30384 = ~n2971 & n30239;
  assign n30385 = pi224 & ~n30384;
  assign n30386 = pi224 & ~n30383;
  assign n30387 = ~n30384 & n30386;
  assign n30388 = ~n30383 & n30385;
  assign n30389 = ~n2971 & n30240;
  assign n30390 = ~n30213 & ~n30376;
  assign n30391 = n2971 & ~n30390;
  assign n30392 = n30382 & ~n30391;
  assign n30393 = ~n30389 & n30392;
  assign n30394 = n30382 & ~n64074;
  assign n30395 = ~n30374 & ~n64075;
  assign n30396 = ~pi299 & ~n30395;
  assign n30397 = pi39 & ~n30396;
  assign n30398 = ~n30366 & n30397;
  assign n30399 = n7844 & n30037;
  assign n30400 = ~n29953 & ~n30399;
  assign n30401 = ~pi224 & ~n30400;
  assign n30402 = n7844 & ~n30037;
  assign n30403 = ~n28846 & n29951;
  assign n30404 = ~n30402 & n30403;
  assign n30405 = ~n30401 & ~n30404;
  assign n30406 = ~pi299 & ~n30405;
  assign n30407 = ~pi614 & n7290;
  assign n30408 = ~n28838 & ~n30407;
  assign n30409 = pi224 & ~n30408;
  assign n30410 = ~pi224 & ~n7852;
  assign n30411 = ~n29957 & n30410;
  assign n30412 = ~n30409 & ~n30411;
  assign n30413 = n30037 & ~n30412;
  assign n30414 = n29959 & ~n30037;
  assign n30415 = pi299 & ~n30414;
  assign n30416 = ~n30413 & n30415;
  assign n30417 = ~n30406 & ~n30416;
  assign n30418 = ~pi39 & ~n30417;
  assign n30419 = ~pi38 & ~n30418;
  assign n30420 = ~n30398 & n30419;
  assign n30421 = pi662 & n7408;
  assign n30422 = n7357 & n30421;
  assign n30423 = n29971 & ~n30422;
  assign n30424 = n62765 & ~n30423;
  assign n30425 = ~n30420 & n30424;
  assign n30426 = ~n29833 & ~n30425;
  assign n30427 = ~pi625 & n30426;
  assign n30428 = pi625 & n29974;
  assign n30429 = ~pi1153 & ~n30428;
  assign n30430 = ~n30427 & n30429;
  assign n30431 = ~pi608 & ~n30133;
  assign n30432 = ~n30430 & n30431;
  assign n30433 = pi625 & n30426;
  assign n30434 = ~pi625 & n29974;
  assign n30435 = pi1153 & ~n30434;
  assign n30436 = ~n30433 & n30435;
  assign n30437 = pi608 & ~n30137;
  assign n30438 = ~n30436 & n30437;
  assign n30439 = ~n30432 & ~n30438;
  assign n30440 = pi778 & ~n30439;
  assign n30441 = ~pi778 & n30426;
  assign n30442 = ~n30440 & ~n30441;
  assign n30443 = ~pi609 & ~n30442;
  assign n30444 = pi609 & n30140;
  assign n30445 = ~pi1155 & ~n30444;
  assign n30446 = ~n30443 & n30445;
  assign n30447 = ~pi660 & ~n29985;
  assign n30448 = ~n30446 & n30447;
  assign n30449 = pi609 & ~n30442;
  assign n30450 = ~pi609 & n30140;
  assign n30451 = pi1155 & ~n30450;
  assign n30452 = ~n30449 & n30451;
  assign n30453 = pi660 & ~n29989;
  assign n30454 = ~n30452 & n30453;
  assign n30455 = ~n30448 & ~n30454;
  assign n30456 = pi785 & ~n30455;
  assign n30457 = ~pi785 & ~n30442;
  assign n30458 = ~n30456 & ~n30457;
  assign n30459 = ~pi618 & ~n30458;
  assign n30460 = pi618 & ~n64056;
  assign n30461 = ~pi1154 & ~n30460;
  assign n30462 = ~n30459 & n30461;
  assign n30463 = ~pi627 & ~n29997;
  assign n30464 = ~n30462 & n30463;
  assign n30465 = pi618 & ~n30458;
  assign n30466 = ~pi618 & ~n64056;
  assign n30467 = pi1154 & ~n30466;
  assign n30468 = ~n30465 & n30467;
  assign n30469 = pi627 & ~n30001;
  assign n30470 = ~n30468 & n30469;
  assign n30471 = ~n30464 & ~n30470;
  assign n30472 = pi781 & ~n30471;
  assign n30473 = ~pi781 & ~n30458;
  assign n30474 = ~n30472 & ~n30473;
  assign n30475 = n63021 & n30474;
  assign n30476 = ~n62884 & n64048;
  assign n30477 = ~n11431 & n64057;
  assign n30478 = ~n30476 & ~n30477;
  assign n30479 = ~n30475 & n30478;
  assign n30480 = pi619 & ~n30474;
  assign n30481 = ~pi619 & ~n64057;
  assign n30482 = pi1159 & ~n30481;
  assign n30483 = ~n30480 & n30482;
  assign n30484 = pi648 & ~n30012;
  assign n30485 = ~n30483 & n30484;
  assign n30486 = ~pi619 & ~n30474;
  assign n30487 = pi619 & ~n64057;
  assign n30488 = ~pi1159 & ~n30487;
  assign n30489 = ~n30486 & n30488;
  assign n30490 = ~pi648 & ~n30008;
  assign n30491 = ~n30489 & n30490;
  assign n30492 = pi789 & ~n30491;
  assign n30493 = ~n30485 & n30492;
  assign n30494 = pi789 & ~n30485;
  assign n30495 = ~n30491 & n30494;
  assign n30496 = pi789 & ~n30479;
  assign n30497 = ~pi789 & n30474;
  assign n30498 = n62894 & ~n30497;
  assign n30499 = ~n64076 & n30498;
  assign n30500 = ~pi626 & ~n64049;
  assign n30501 = pi626 & n29831;
  assign n30502 = n8301 & ~n30501;
  assign n30503 = ~n30500 & n30502;
  assign n30504 = n8257 & ~n29831;
  assign n30505 = ~n30153 & ~n30504;
  assign n30506 = n8525 & ~n30505;
  assign n30507 = pi626 & ~n64049;
  assign n30508 = ~pi626 & n29831;
  assign n30509 = n8300 & ~n30508;
  assign n30510 = ~n30507 & n30509;
  assign n30511 = ~n30506 & ~n30510;
  assign n30512 = ~n30503 & ~n30506;
  assign n30513 = ~n30510 & n30512;
  assign n30514 = ~n30503 & n30511;
  assign n30515 = pi788 & ~n64077;
  assign n30516 = ~n63030 & ~n30515;
  assign n30517 = ~n30499 & n30516;
  assign n30518 = ~n30196 & ~n30517;
  assign n30519 = ~n8651 & ~n30518;
  assign n30520 = ~n8334 & ~n30180;
  assign n30521 = n8334 & ~n29831;
  assign n30522 = ~n8413 & ~n30521;
  assign n30523 = ~n8334 & n30180;
  assign n30524 = n8334 & n29831;
  assign n30525 = ~n30523 & ~n30524;
  assign n30526 = ~n8413 & ~n30525;
  assign n30527 = ~n30520 & n30522;
  assign n30528 = ~pi630 & n30165;
  assign n30529 = pi630 & n30169;
  assign n30530 = ~n30528 & ~n30529;
  assign n30531 = ~n64078 & n30530;
  assign n30532 = pi787 & ~n30531;
  assign n30533 = ~n11547 & ~n30532;
  assign n30534 = ~n30519 & n30533;
  assign n30535 = ~n30519 & ~n30532;
  assign n30536 = pi644 & n30535;
  assign n30537 = ~n30171 & ~n30172;
  assign n30538 = ~pi644 & n30537;
  assign n30539 = pi715 & ~n30538;
  assign n30540 = ~n30536 & n30539;
  assign n30541 = ~n11558 & ~n29831;
  assign n30542 = n8376 & ~n29831;
  assign n30543 = ~n8376 & n30525;
  assign n30544 = ~n30542 & ~n30543;
  assign n30545 = ~n30026 & ~n30541;
  assign n30546 = pi644 & ~n64079;
  assign n30547 = ~pi644 & ~n29831;
  assign n30548 = ~pi715 & ~n30547;
  assign n30549 = ~n30546 & n30548;
  assign n30550 = pi1160 & ~n30549;
  assign n30551 = ~n30540 & n30550;
  assign n30552 = ~pi644 & n30535;
  assign n30553 = pi644 & n30537;
  assign n30554 = ~pi715 & ~n30553;
  assign n30555 = ~n30552 & n30554;
  assign n30556 = ~pi644 & ~n64079;
  assign n30557 = pi644 & ~n29831;
  assign n30558 = pi715 & ~n30557;
  assign n30559 = ~n30556 & n30558;
  assign n30560 = ~pi1160 & ~n30559;
  assign n30561 = ~n30555 & n30560;
  assign n30562 = ~n30551 & ~n30561;
  assign n30563 = pi790 & ~n30562;
  assign n30564 = ~pi790 & n30535;
  assign n30565 = ~n30563 & ~n30564;
  assign n30566 = ~n30178 & ~n30534;
  assign n30567 = n62455 & ~n64080;
  assign n30568 = ~pi224 & ~n62455;
  assign po381 = ~n30567 & ~n30568;
  assign n30570 = pi57 & pi59;
  assign n30571 = ~pi87 & n2764;
  assign n30572 = ~pi92 & n2765;
  assign n30573 = n30571 & n30572;
  assign n30574 = n2806 & n6793;
  assign n30575 = n62373 & n6796;
  assign n30576 = n62373 & n6797;
  assign n30577 = ~pi39 & n62952;
  assign n30578 = ~pi87 & n62374;
  assign n30579 = n62373 & n6795;
  assign n30580 = n2765 & n30571;
  assign n30581 = n2580 & n64083;
  assign n30582 = n2764 & n62765;
  assign n30583 = n6792 & n64081;
  assign n30584 = ~pi55 & n6797;
  assign n30585 = ~pi55 & n64082;
  assign n30586 = n62373 & n30584;
  assign n30587 = n3470 & n64084;
  assign n30588 = n3471 & n64082;
  assign n30589 = n62380 & n64085;
  assign n30590 = ~n3472 & ~n30589;
  assign n30591 = ~n30570 & ~n30590;
  assign n30592 = ~pi54 & n6796;
  assign n30593 = n62373 & n30592;
  assign n30594 = ~pi54 & n64081;
  assign n30595 = n62373 & n62380;
  assign n30596 = n30592 & n30595;
  assign n30597 = n62380 & n64086;
  assign n30598 = pi74 & ~n64087;
  assign n30599 = n7356 & n62951;
  assign n30600 = pi75 & ~n30599;
  assign n30601 = n2766 & n6795;
  assign n30602 = n2765 & n9735;
  assign n30603 = n7356 & n64088;
  assign n30604 = pi92 & ~n30603;
  assign n30605 = ~n30600 & ~n30604;
  assign n30606 = pi38 & ~n7356;
  assign n30607 = pi145 & pi180;
  assign n30608 = pi181 & pi182;
  assign n30609 = n30607 & n30608;
  assign n30610 = pi32 & n6909;
  assign n30611 = ~pi95 & n30610;
  assign n30612 = ~pi198 & n30611;
  assign n30613 = pi95 & ~pi479;
  assign n30614 = n2795 & n30613;
  assign n30615 = ~pi51 & n62767;
  assign n30616 = n2694 & n62770;
  assign n30617 = n62357 & n64089;
  assign n30618 = pi72 & ~n30617;
  assign n30619 = n2751 & ~n30618;
  assign n30620 = pi70 & ~n62364;
  assign n30621 = ~pi51 & ~n30620;
  assign n30622 = ~pi96 & n30621;
  assign n30623 = n2787 & ~n30620;
  assign n30624 = pi841 & n2659;
  assign n30625 = pi93 & ~n30624;
  assign n30626 = ~pi35 & ~n30625;
  assign n30627 = pi90 & ~n62357;
  assign n30628 = ~pi91 & ~pi314;
  assign n30629 = pi46 & n2639;
  assign n30630 = n62389 & n30629;
  assign n30631 = ~pi60 & n2627;
  assign n30632 = ~pi60 & n62348;
  assign n30633 = n2625 & n30631;
  assign n30634 = n2587 & n64091;
  assign n30635 = ~pi60 & n62349;
  assign n30636 = n2630 & n30631;
  assign n30637 = pi53 & ~n64092;
  assign n30638 = pi60 & n62349;
  assign n30639 = ~pi53 & ~n30638;
  assign n30640 = pi50 & ~n2860;
  assign n30641 = ~pi60 & ~n30640;
  assign n30642 = pi77 & n2611;
  assign n30643 = pi77 & n2859;
  assign n30644 = n62358 & n30642;
  assign n30645 = ~pi50 & ~n64093;
  assign n30646 = pi69 & ~n2607;
  assign n30647 = pi83 & ~n62345;
  assign n30648 = ~pi103 & ~n30647;
  assign n30649 = ~n30646 & n30648;
  assign n30650 = n2596 & n2601;
  assign n30651 = ~pi84 & n30650;
  assign n30652 = ~pi68 & ~pi111;
  assign n30653 = pi82 & n30652;
  assign n30654 = ~pi68 & n30651;
  assign n30655 = pi82 & ~pi111;
  assign n30656 = n30654 & n30655;
  assign n30657 = n30651 & n30653;
  assign n30658 = pi66 & pi73;
  assign n30659 = ~n2596 & ~n2601;
  assign n30660 = ~n30658 & ~n30659;
  assign n30661 = pi85 & pi106;
  assign n30662 = n2589 & ~n30661;
  assign n30663 = pi61 & pi76;
  assign n30664 = n2590 & ~n30663;
  assign n30665 = ~n30662 & ~n30664;
  assign n30666 = ~pi48 & ~n30665;
  assign n30667 = ~n2591 & ~n30666;
  assign n30668 = pi89 & ~n2592;
  assign n30669 = ~pi49 & ~n30668;
  assign n30670 = ~n30667 & n30669;
  assign n30671 = ~n2593 & ~n30670;
  assign n30672 = pi104 & ~n2594;
  assign n30673 = ~pi45 & ~n30672;
  assign n30674 = ~n30671 & n30673;
  assign n30675 = ~n2595 & ~n30674;
  assign n30676 = ~n2596 & ~n30675;
  assign n30677 = pi85 & n30676;
  assign n30678 = n2601 & ~n30677;
  assign n30679 = n30660 & ~n30678;
  assign n30680 = n2597 & ~n30679;
  assign n30681 = pi84 & ~n30650;
  assign n30682 = pi68 & ~n30651;
  assign n30683 = ~n30681 & ~n30682;
  assign n30684 = ~n30680 & n30683;
  assign n30685 = n2598 & n30684;
  assign n30686 = ~n64094 & ~n30685;
  assign n30687 = n6806 & ~n30686;
  assign n30688 = pi67 & n62344;
  assign n30689 = n6810 & ~n30688;
  assign n30690 = ~n30687 & n30689;
  assign n30691 = n30649 & ~n30690;
  assign n30692 = ~pi71 & ~n30691;
  assign n30693 = pi71 & ~n2610;
  assign n30694 = ~pi65 & ~n30693;
  assign n30695 = ~pi64 & n2587;
  assign n30696 = n30694 & n30695;
  assign n30697 = ~n30692 & n30696;
  assign n30698 = ~pi81 & ~n30697;
  assign n30699 = ~pi83 & pi103;
  assign n30700 = pi103 & n6810;
  assign n30701 = n2607 & n30700;
  assign n30702 = n62345 & n30699;
  assign n30703 = n30696 & n64095;
  assign n30704 = n30698 & ~n30703;
  assign n30705 = pi81 & ~n2632;
  assign n30706 = ~pi102 & ~n30705;
  assign n30707 = n2612 & n30706;
  assign n30708 = ~n30704 & n30707;
  assign n30709 = n30645 & ~n30708;
  assign n30710 = n30641 & ~n30709;
  assign n30711 = n30639 & ~n30710;
  assign n30712 = ~n30637 & ~n30711;
  assign n30713 = ~pi86 & ~n30712;
  assign n30714 = pi86 & ~n2861;
  assign n30715 = ~pi94 & ~n30714;
  assign n30716 = n2643 & n30715;
  assign n30717 = ~n30713 & n30716;
  assign n30718 = ~n30630 & ~n30717;
  assign n30719 = n2870 & ~n30718;
  assign n30720 = n30628 & ~n30719;
  assign n30721 = pi91 & ~n2856;
  assign n30722 = ~pi58 & ~n30721;
  assign n30723 = ~pi91 & pi314;
  assign n30724 = ~n30698 & n30707;
  assign n30725 = n30645 & ~n30724;
  assign n30726 = n30641 & ~n30725;
  assign n30727 = n30639 & ~n30726;
  assign n30728 = ~n30637 & ~n30727;
  assign n30729 = ~pi86 & ~n30728;
  assign n30730 = n30716 & ~n30729;
  assign n30731 = ~n30630 & ~n30730;
  assign n30732 = n2870 & ~n30731;
  assign n30733 = n30723 & ~n30732;
  assign n30734 = n30722 & ~n30733;
  assign n30735 = ~n30720 & n30734;
  assign n30736 = ~pi90 & ~n30735;
  assign n30737 = ~n30627 & ~n30736;
  assign n30738 = ~pi93 & ~n30737;
  assign n30739 = n30626 & ~n30738;
  assign n30740 = ~pi70 & ~n30739;
  assign n30741 = n64090 & ~n30740;
  assign n30742 = ~pi72 & ~n30741;
  assign n30743 = n30619 & ~n30742;
  assign n30744 = ~n30614 & ~n30743;
  assign n30745 = ~n30612 & n30744;
  assign n30746 = n2814 & ~n30745;
  assign n30747 = n30609 & n30746;
  assign n30748 = pi109 & ~n2671;
  assign n30749 = n2866 & ~n30748;
  assign n30750 = ~pi109 & ~n30630;
  assign n30751 = ~n30717 & n30750;
  assign n30752 = n30749 & ~n30751;
  assign n30753 = n30628 & ~n30752;
  assign n30754 = ~n30730 & n30750;
  assign n30755 = n30749 & ~n30754;
  assign n30756 = n30723 & ~n30755;
  assign n30757 = n30722 & ~n30756;
  assign n30758 = ~n30753 & n30757;
  assign n30759 = ~pi90 & ~n30758;
  assign n30760 = ~n30627 & ~n30759;
  assign n30761 = ~pi93 & ~n30760;
  assign n30762 = n30626 & ~n30761;
  assign n30763 = ~pi70 & ~n30762;
  assign n30764 = n64090 & ~n30763;
  assign n30765 = ~pi72 & ~n30764;
  assign n30766 = n30619 & ~n30765;
  assign n30767 = ~n30614 & ~n30766;
  assign n30768 = ~n30612 & n30767;
  assign n30769 = ~n30609 & ~n30768;
  assign n30770 = ~n2814 & ~n30768;
  assign n30771 = ~pi299 & ~n30770;
  assign n30772 = ~n30769 & n30771;
  assign n30773 = ~n30747 & n30772;
  assign n30774 = pi160 & pi197;
  assign n30775 = ~pi210 & n30611;
  assign n30776 = n30744 & ~n30775;
  assign n30777 = n2814 & ~n30776;
  assign n30778 = n30774 & ~n30777;
  assign n30779 = n30767 & ~n30775;
  assign n30780 = ~n30774 & n30779;
  assign n30781 = ~n30778 & ~n30780;
  assign n30782 = ~n2814 & ~n30779;
  assign n30783 = pi158 & pi159;
  assign n30784 = pi299 & n30783;
  assign n30785 = ~n30782 & n30784;
  assign n30786 = ~n30781 & n30785;
  assign n30787 = pi299 & n30779;
  assign n30788 = ~n30783 & n30787;
  assign n30789 = pi232 & ~n30788;
  assign n30790 = ~n30786 & n30789;
  assign n30791 = ~n30773 & n30789;
  assign n30792 = ~n30786 & n30791;
  assign n30793 = ~n30773 & n30790;
  assign n30794 = ~pi299 & n30768;
  assign n30795 = ~pi232 & ~n30787;
  assign n30796 = ~n30794 & n30795;
  assign n30797 = ~pi39 & ~n30796;
  assign n30798 = ~n30773 & ~n30786;
  assign n30799 = pi232 & ~n30798;
  assign n30800 = ~pi232 & ~pi299;
  assign n30801 = n30768 & n30800;
  assign n30802 = pi232 & n30783;
  assign n30803 = pi299 & ~n30802;
  assign n30804 = n30779 & n30803;
  assign n30805 = ~n30787 & ~n30794;
  assign n30806 = ~n30789 & ~n30805;
  assign n30807 = ~n30801 & ~n30804;
  assign n30808 = ~n30799 & ~n64097;
  assign n30809 = ~pi39 & ~n30808;
  assign n30810 = ~n64096 & n30797;
  assign n30811 = n2939 & n62442;
  assign n30812 = ~pi1091 & n30811;
  assign n30813 = pi1091 & n2824;
  assign n30814 = n2582 & ~n30813;
  assign n30815 = n3322 & n30814;
  assign n30816 = n62442 & ~n30813;
  assign n30817 = ~n62395 & ~n64099;
  assign n30818 = pi1091 & ~n30817;
  assign n30819 = n2939 & n30818;
  assign n30820 = ~n30812 & ~n30819;
  assign n30821 = pi216 & ~n30820;
  assign n30822 = ~pi829 & ~n2824;
  assign n30823 = pi1091 & ~n30822;
  assign n30824 = n30811 & ~n30823;
  assign n30825 = ~pi216 & n30824;
  assign n30826 = ~pi216 & ~n30824;
  assign n30827 = pi216 & n30820;
  assign n30828 = ~n30826 & ~n30827;
  assign n30829 = ~n30821 & ~n30825;
  assign n30830 = n2960 & n64100;
  assign n30831 = pi299 & ~n2920;
  assign n30832 = n30830 & n30831;
  assign n30833 = ~pi224 & ~n30824;
  assign n30834 = pi224 & n30820;
  assign n30835 = pi224 & ~n30820;
  assign n30836 = ~pi224 & n30824;
  assign n30837 = ~n30835 & ~n30836;
  assign n30838 = ~n30833 & ~n30834;
  assign n30839 = pi222 & ~n2973;
  assign n30840 = n2979 & n30839;
  assign n30841 = ~pi299 & ~n2973;
  assign n30842 = n2980 & n30841;
  assign n30843 = ~n2973 & n62403;
  assign n30844 = n2980 & ~n30833;
  assign n30845 = n2980 & ~n64101;
  assign n30846 = ~n30834 & n30844;
  assign n30847 = n30841 & n64103;
  assign n30848 = ~n64101 & n64102;
  assign n30849 = pi39 & ~n64104;
  assign n30850 = ~n30832 & n30849;
  assign n30851 = ~n64098 & ~n30850;
  assign n30852 = ~pi38 & ~n30851;
  assign n30853 = ~n30606 & ~n30852;
  assign n30854 = ~pi100 & ~n30853;
  assign n30855 = ~pi38 & pi100;
  assign n30856 = n7356 & n30855;
  assign n30857 = ~pi252 & n62380;
  assign n30858 = ~pi142 & ~n2808;
  assign n30859 = ~pi299 & n30858;
  assign n30860 = ~pi146 & ~n2811;
  assign n30861 = pi299 & n30860;
  assign n30862 = pi146 & n2812;
  assign n30863 = pi142 & n2809;
  assign n30864 = ~n30862 & ~n30863;
  assign n30865 = ~n2813 & n30864;
  assign n30866 = ~n30859 & ~n30861;
  assign n30867 = n30857 & ~n64105;
  assign n30868 = ~pi683 & ~n2843;
  assign n30869 = ~pi250 & ~po740;
  assign n30870 = pi129 & pi250;
  assign n30871 = ~n30869 & ~n30870;
  assign n30872 = ~n30868 & ~n30871;
  assign n30873 = n64105 & ~n30872;
  assign n30874 = n2843 & n64105;
  assign n30875 = ~n30873 & ~n30874;
  assign n30876 = ~n30857 & ~n64105;
  assign n30877 = ~n2843 & n64105;
  assign n30878 = n30872 & n30877;
  assign n30879 = ~n30876 & ~n30878;
  assign n30880 = ~n30867 & n30875;
  assign n30881 = n30856 & ~n30878;
  assign n30882 = ~n30876 & n30881;
  assign n30883 = n30856 & n64106;
  assign n30884 = ~pi38 & n7356;
  assign n30885 = pi100 & ~n30884;
  assign n30886 = ~pi87 & ~n30885;
  assign n30887 = ~pi87 & ~n64107;
  assign n30888 = ~n30885 & n30887;
  assign n30889 = ~n64107 & n30886;
  assign n30890 = ~n30854 & n64108;
  assign n30891 = n6793 & ~n30890;
  assign n30892 = n30605 & ~n30891;
  assign n30893 = ~pi54 & ~n30892;
  assign n30894 = ~pi92 & n30603;
  assign n30895 = pi54 & ~n30894;
  assign n30896 = ~n30893 & ~n30895;
  assign n30897 = ~pi74 & ~n30896;
  assign n30898 = ~n30598 & ~n30897;
  assign n30899 = ~pi55 & ~n30898;
  assign n30900 = ~pi74 & n64087;
  assign n30901 = n6797 & n30595;
  assign n30902 = n62380 & n64082;
  assign n30903 = pi55 & ~n64109;
  assign n30904 = ~pi56 & ~n30903;
  assign n30905 = ~pi62 & n30904;
  assign n30906 = ~n30899 & n30905;
  assign n30907 = n3472 & ~n30906;
  assign po195 = n30591 & ~n30907;
  assign n30909 = ~pi954 & ~po195;
  assign n30910 = pi24 & pi954;
  assign po182 = ~n30909 & ~n30910;
  assign n30912 = ~pi31 & ~pi80;
  assign n30913 = pi818 & n30912;
  assign n30914 = ~n2580 & n3036;
  assign n30915 = ~n3318 & ~n30914;
  assign n30916 = ~pi120 & ~n2580;
  assign n30917 = ~pi1093 & n30916;
  assign n30918 = n30915 & ~n30917;
  assign n30919 = n62380 & n2846;
  assign n30920 = pi120 & ~n3036;
  assign n30921 = ~n2996 & n30920;
  assign n30922 = ~pi120 & pi1093;
  assign n30923 = pi120 & n2996;
  assign n30924 = n2996 & ~n30922;
  assign n30925 = ~pi120 & n30919;
  assign n30926 = ~n64110 & ~n30925;
  assign n30927 = n30919 & ~n30921;
  assign n30928 = n2998 & ~n64111;
  assign n30929 = ~pi1091 & n5791;
  assign n30930 = n30922 & ~n30929;
  assign n30931 = ~n30920 & ~n30930;
  assign n30932 = pi100 & ~n30931;
  assign n30933 = ~n30928 & n30932;
  assign n30934 = ~pi1093 & n2761;
  assign n30935 = pi120 & n30934;
  assign n30936 = ~pi39 & ~n30935;
  assign n30937 = pi97 & ~n62389;
  assign n30938 = ~pi108 & ~n30937;
  assign n30939 = ~pi110 & n30938;
  assign n30940 = n2636 & n2867;
  assign n30941 = ~n2693 & n30940;
  assign n30942 = n30939 & n30941;
  assign n30943 = ~n2858 & ~n30942;
  assign n30944 = n2586 & ~n30943;
  assign n30945 = n2676 & ~n30944;
  assign n30946 = n2662 & ~n30945;
  assign n30947 = ~pi51 & ~n30946;
  assign n30948 = ~n2725 & ~n30947;
  assign n30949 = ~pi96 & ~n30948;
  assign n30950 = n62392 & ~n30949;
  assign n30951 = n62368 & n2852;
  assign n30952 = ~pi829 & n30951;
  assign n30953 = ~pi122 & ~n30952;
  assign n30954 = ~n30950 & n30953;
  assign n30955 = pi122 & ~n2739;
  assign n30956 = ~n2824 & ~n30955;
  assign n30957 = ~n30954 & n30956;
  assign n30958 = n2924 & ~n30957;
  assign n30959 = n3032 & ~n30951;
  assign n30960 = ~n5791 & n30959;
  assign n30961 = ~n30958 & ~n30960;
  assign n30962 = n30936 & n30961;
  assign n30963 = n2953 & ~n30931;
  assign n30964 = ~n62397 & n30920;
  assign n30965 = pi1091 & pi1092;
  assign n30966 = n62398 & n30965;
  assign n30967 = n2929 & n62396;
  assign n30968 = n30930 & ~n64112;
  assign n30969 = ~n30964 & ~n30968;
  assign n30970 = ~n2953 & ~n30969;
  assign n30971 = ~n30963 & ~n30970;
  assign n30972 = ~n2971 & ~n30971;
  assign n30973 = ~n2909 & n30931;
  assign n30974 = n2909 & n30969;
  assign n30975 = ~n30973 & ~n30974;
  assign n30976 = n2971 & n30975;
  assign n30977 = n3076 & ~n30976;
  assign n30978 = n3076 & ~n30972;
  assign n30979 = ~n30976 & n30978;
  assign n30980 = ~n30972 & n30977;
  assign n30981 = ~n3076 & n30931;
  assign n30982 = ~pi299 & ~n30981;
  assign n30983 = ~n64113 & n30982;
  assign n30984 = ~n62393 & ~n30971;
  assign n30985 = n62393 & n30975;
  assign n30986 = n3056 & ~n30985;
  assign n30987 = n3056 & ~n30984;
  assign n30988 = ~n30985 & n30987;
  assign n30989 = ~n30984 & n30986;
  assign n30990 = ~n3056 & n30931;
  assign n30991 = pi299 & ~n30990;
  assign n30992 = ~n64114 & n30991;
  assign n30993 = pi39 & ~n30992;
  assign n30994 = pi39 & ~n30983;
  assign n30995 = ~n30992 & n30994;
  assign n30996 = ~n30983 & n30993;
  assign n30997 = ~n30962 & ~n64115;
  assign n30998 = ~pi38 & ~n30997;
  assign n30999 = ~pi120 & ~pi1093;
  assign n31000 = pi38 & n30999;
  assign n31001 = ~pi100 & ~n31000;
  assign n31002 = ~n3093 & n31001;
  assign n31003 = ~n30998 & n31002;
  assign n31004 = ~n30933 & ~n31003;
  assign n31005 = ~pi87 & ~n31004;
  assign n31006 = n3336 & ~n30999;
  assign n31007 = n3032 & ~n5791;
  assign n31008 = ~n3118 & n31007;
  assign n31009 = n3334 & ~n31008;
  assign n31010 = ~n62373 & n3036;
  assign n31011 = pi87 & ~n31010;
  assign n31012 = ~n31009 & n31011;
  assign n31013 = n31006 & n31012;
  assign n31014 = ~n31005 & ~n31013;
  assign n31015 = ~pi75 & ~n31014;
  assign n31016 = n2816 & n30931;
  assign n31017 = ~n2847 & n30930;
  assign n31018 = ~pi1091 & ~n3035;
  assign n31019 = ~n3025 & ~n31018;
  assign n31020 = pi120 & ~n31019;
  assign n31021 = ~n2816 & ~n31020;
  assign n31022 = ~n31017 & n31021;
  assign n31023 = ~n31016 & ~n31022;
  assign n31024 = n2806 & ~n31023;
  assign n31025 = ~n2806 & n30931;
  assign n31026 = pi75 & ~n31025;
  assign n31027 = ~n31024 & n31026;
  assign n31028 = n2580 & ~n31027;
  assign n31029 = ~n31015 & n31028;
  assign n31030 = n30918 & ~n31029;
  assign n31031 = ~n30958 & ~n30959;
  assign n31032 = n30936 & n31031;
  assign n31033 = ~pi299 & ~n30999;
  assign n31034 = ~n62537 & n31033;
  assign n31035 = pi299 & ~n30999;
  assign n31036 = ~n62538 & n31035;
  assign n31037 = pi39 & ~n31036;
  assign n31038 = pi39 & ~n31034;
  assign n31039 = ~n31036 & n31038;
  assign n31040 = ~n31034 & n31037;
  assign n31041 = ~n31032 & ~n64116;
  assign n31042 = ~pi38 & ~n31041;
  assign n31043 = n31001 & ~n31042;
  assign n31044 = pi100 & ~n30999;
  assign n31045 = ~n30928 & n31044;
  assign n31046 = ~n31043 & ~n31045;
  assign n31047 = ~pi87 & ~n31046;
  assign n31048 = ~n31006 & ~n31047;
  assign n31049 = ~pi75 & ~n31048;
  assign n31050 = n2850 & ~n30999;
  assign n31051 = n2580 & ~n31050;
  assign n31052 = ~n31049 & n31051;
  assign n31053 = n3318 & ~n30917;
  assign n31054 = ~n31052 & n31053;
  assign n31055 = ~n31030 & ~n31054;
  assign n31056 = n30913 & ~n31055;
  assign n31057 = n62455 & ~n31056;
  assign n31058 = ~n3318 & n30931;
  assign n31059 = pi120 & ~n31058;
  assign n31060 = n30913 & ~n30999;
  assign n31061 = ~n31058 & n31060;
  assign n31062 = ~n62455 & ~n31061;
  assign n31063 = ~n31059 & n31062;
  assign n31064 = ~n5530 & ~n31063;
  assign n31065 = pi951 & pi982;
  assign n31066 = pi1092 & n31065;
  assign n31067 = pi1093 & n31066;
  assign n31068 = ~pi120 & ~n31067;
  assign n31069 = ~n31058 & ~n31068;
  assign n31070 = n31062 & ~n31069;
  assign n31071 = n5530 & ~n31070;
  assign n31072 = ~n31064 & ~n31071;
  assign n31073 = ~n31057 & ~n31072;
  assign n31074 = pi120 & n2848;
  assign n31075 = ~pi1091 & n31067;
  assign n31076 = ~pi120 & ~n31075;
  assign n31077 = n2924 & n31066;
  assign n31078 = pi252 & n2751;
  assign n31079 = ~pi24 & ~pi90;
  assign n31080 = pi950 & n2581;
  assign n31081 = ~pi122 & n2921;
  assign n31082 = n31079 & n64117;
  assign n31083 = n31078 & n31082;
  assign n31084 = ~pi93 & ~pi122;
  assign n31085 = n2729 & n31084;
  assign n31086 = n2921 & n31079;
  assign n31087 = n31085 & n31086;
  assign n31088 = n62769 & n31082;
  assign n31089 = n6832 & n31079;
  assign n31090 = n64117 & n31089;
  assign n31091 = n62770 & n31090;
  assign n31092 = n2743 & n31087;
  assign n31093 = n31078 & n64118;
  assign n31094 = n62769 & n31083;
  assign n31095 = n2844 & n64119;
  assign n31096 = n62357 & n31095;
  assign n31097 = n31077 & ~n31096;
  assign n31098 = n31076 & ~n31097;
  assign n31099 = ~n31074 & ~n31098;
  assign n31100 = ~n2816 & ~n31099;
  assign n31101 = n2816 & n31068;
  assign n31102 = n2806 & ~n31101;
  assign n31103 = ~n31100 & n31102;
  assign n31104 = ~n2806 & ~n31068;
  assign n31105 = pi75 & ~n31104;
  assign n31106 = ~n31103 & n31105;
  assign n31107 = n2581 & n2844;
  assign n31108 = n3113 & n31107;
  assign n31109 = n31077 & ~n31108;
  assign n31110 = n31076 & ~n31109;
  assign n31111 = ~n64110 & ~n31110;
  assign n31112 = ~pi39 & n2997;
  assign n31113 = ~n31111 & n31112;
  assign n31114 = pi100 & ~n31113;
  assign n31115 = ~pi38 & ~n31114;
  assign n31116 = ~n2998 & n31068;
  assign n31117 = ~n31115 & ~n31116;
  assign n31118 = ~n30934 & n31031;
  assign n31119 = pi120 & n31118;
  assign n31120 = n62391 & ~n30949;
  assign n31121 = n2581 & n31066;
  assign n31122 = ~n31120 & n31121;
  assign n31123 = pi950 & n62367;
  assign n31124 = ~n2714 & n31123;
  assign n31125 = pi122 & n2887;
  assign n31126 = pi122 & n31065;
  assign n31127 = n2887 & n31126;
  assign n31128 = n31065 & n31125;
  assign n31129 = ~n31124 & n64120;
  assign n31130 = pi824 & n31124;
  assign n31131 = n31066 & ~n31130;
  assign n31132 = ~pi829 & n31131;
  assign n31133 = ~n31129 & ~n31132;
  assign n31134 = ~n31122 & n31133;
  assign n31135 = n2851 & ~n31134;
  assign n31136 = n2824 & n31067;
  assign n31137 = n3007 & n31066;
  assign n31138 = ~n31135 & ~n64121;
  assign n31139 = pi1091 & ~n31138;
  assign n31140 = n3032 & n31131;
  assign n31141 = n31075 & ~n31130;
  assign n31142 = ~pi120 & ~n64122;
  assign n31143 = ~n31139 & n31142;
  assign n31144 = ~pi39 & ~n31143;
  assign n31145 = ~pi39 & ~n31119;
  assign n31146 = ~n31143 & n31145;
  assign n31147 = ~n31119 & n31144;
  assign n31148 = pi39 & ~n31068;
  assign n31149 = ~n3076 & n31068;
  assign n31150 = ~pi299 & ~n31149;
  assign n31151 = ~n2954 & ~n31068;
  assign n31152 = ~n2971 & n31151;
  assign n31153 = ~n2950 & ~n31068;
  assign n31154 = n2971 & n31153;
  assign n31155 = n3076 & ~n31154;
  assign n31156 = n3076 & ~n31152;
  assign n31157 = ~n31154 & n31156;
  assign n31158 = ~n31152 & n31155;
  assign n31159 = n31150 & ~n64124;
  assign n31160 = ~n3056 & n31068;
  assign n31161 = pi299 & ~n31160;
  assign n31162 = ~n62393 & n31151;
  assign n31163 = n62393 & n31153;
  assign n31164 = n3056 & ~n31163;
  assign n31165 = n3056 & ~n31162;
  assign n31166 = ~n31163 & n31165;
  assign n31167 = ~n31162 & n31164;
  assign n31168 = n31161 & ~n64125;
  assign n31169 = ~n31159 & ~n31168;
  assign n31170 = pi39 & ~n31169;
  assign n31171 = n62539 & n31148;
  assign n31172 = ~n64123 & ~n64126;
  assign n31173 = n2766 & ~n31172;
  assign n31174 = ~n31117 & ~n31173;
  assign n31175 = ~pi87 & ~n31174;
  assign n31176 = ~n62373 & n31068;
  assign n31177 = pi87 & ~n31176;
  assign n31178 = n3113 & n6959;
  assign n31179 = n31077 & ~n31178;
  assign n31180 = ~n62420 & n31075;
  assign n31181 = ~n31179 & ~n31180;
  assign n31182 = ~pi120 & ~n31181;
  assign n31183 = ~n3332 & ~n3333;
  assign n31184 = pi120 & ~n31183;
  assign n31185 = n62373 & ~n31184;
  assign n31186 = ~n31182 & n31185;
  assign n31187 = n31177 & ~n31186;
  assign n31188 = ~pi75 & ~n31187;
  assign n31189 = ~n31175 & n31188;
  assign n31190 = ~n31106 & ~n31189;
  assign n31191 = n2580 & ~n31190;
  assign n31192 = n3318 & ~n31191;
  assign n31193 = ~n5791 & n31075;
  assign n31194 = ~n31109 & ~n31193;
  assign n31195 = ~pi120 & ~n31194;
  assign n31196 = ~n30921 & ~n31195;
  assign n31197 = n2997 & ~n31196;
  assign n31198 = ~n30931 & ~n31068;
  assign n31199 = ~n2997 & n31198;
  assign n31200 = n2764 & ~n31199;
  assign n31201 = ~n31197 & n31200;
  assign n31202 = ~n2764 & ~n31198;
  assign n31203 = pi100 & ~n31202;
  assign n31204 = ~n31201 & n31203;
  assign n31205 = ~n30934 & n30961;
  assign n31206 = pi120 & n31205;
  assign n31207 = n31007 & n31131;
  assign n31208 = ~pi120 & ~n31207;
  assign n31209 = ~n31139 & n31208;
  assign n31210 = ~pi39 & ~n31209;
  assign n31211 = ~n31206 & n31210;
  assign n31212 = ~n62398 & n31077;
  assign n31213 = ~n31193 & ~n31212;
  assign n31214 = ~pi120 & ~n31213;
  assign n31215 = ~n30964 & ~n31214;
  assign n31216 = ~n2953 & ~n31215;
  assign n31217 = n2953 & n31198;
  assign n31218 = ~n31216 & ~n31217;
  assign n31219 = ~n2971 & ~n31218;
  assign n31220 = n2909 & ~n31215;
  assign n31221 = ~n2909 & n31198;
  assign n31222 = ~n31220 & ~n31221;
  assign n31223 = n2971 & ~n31222;
  assign n31224 = n3076 & ~n31223;
  assign n31225 = n3076 & ~n31219;
  assign n31226 = ~n31223 & n31225;
  assign n31227 = ~n31219 & n31224;
  assign n31228 = ~n3076 & ~n31198;
  assign n31229 = ~pi299 & ~n31228;
  assign n31230 = ~n30981 & n31150;
  assign n31231 = ~n64127 & n64128;
  assign n31232 = ~n62393 & ~n31218;
  assign n31233 = n62393 & ~n31222;
  assign n31234 = n3056 & ~n31233;
  assign n31235 = n3056 & ~n31232;
  assign n31236 = ~n31233 & n31235;
  assign n31237 = ~n31232 & n31234;
  assign n31238 = pi299 & ~n3070;
  assign n31239 = ~n3070 & n31161;
  assign n31240 = ~n31160 & n31238;
  assign n31241 = ~n64129 & n64130;
  assign n31242 = ~n31231 & ~n31241;
  assign n31243 = pi39 & ~n31242;
  assign n31244 = ~pi38 & ~n31243;
  assign n31245 = ~n31206 & ~n31209;
  assign n31246 = ~pi39 & ~n31245;
  assign n31247 = pi39 & ~n31241;
  assign n31248 = pi39 & ~n31231;
  assign n31249 = ~n31241 & n31248;
  assign n31250 = ~n31231 & n31247;
  assign n31251 = ~n31246 & ~n64131;
  assign n31252 = ~pi38 & ~n31251;
  assign n31253 = ~n31211 & n31244;
  assign n31254 = pi38 & ~n31198;
  assign n31255 = ~pi100 & ~n31254;
  assign n31256 = ~n64132 & n31255;
  assign n31257 = ~n31204 & ~n31256;
  assign n31258 = ~pi87 & ~n31257;
  assign n31259 = ~n31009 & ~n31185;
  assign n31260 = ~n31179 & ~n31193;
  assign n31261 = n31182 & ~n31260;
  assign n31262 = ~n31259 & ~n31261;
  assign n31263 = ~n31010 & n31177;
  assign n31264 = ~n31262 & n31263;
  assign n31265 = ~n31258 & ~n31264;
  assign n31266 = ~pi75 & ~n31265;
  assign n31267 = n2816 & ~n31198;
  assign n31268 = ~n31097 & ~n31193;
  assign n31269 = ~pi120 & ~n31268;
  assign n31270 = n31021 & ~n31269;
  assign n31271 = ~n31267 & ~n31270;
  assign n31272 = n2806 & ~n31271;
  assign n31273 = ~n2806 & ~n31198;
  assign n31274 = pi75 & ~n31273;
  assign n31275 = ~n31272 & n31274;
  assign n31276 = n2580 & ~n31275;
  assign n31277 = ~n31266 & n31276;
  assign n31278 = n30918 & ~n31277;
  assign n31279 = ~n31192 & ~n31278;
  assign n31280 = n30916 & ~n31067;
  assign n31281 = n31071 & ~n31280;
  assign n31282 = ~n31279 & n31281;
  assign n31283 = ~pi39 & ~n31118;
  assign n31284 = n2990 & ~n31283;
  assign n31285 = ~pi100 & ~n31284;
  assign n31286 = ~n3003 & ~n31285;
  assign n31287 = ~pi87 & ~n31286;
  assign n31288 = ~n3336 & ~n31287;
  assign n31289 = ~pi75 & ~n31288;
  assign n31290 = ~n2850 & ~n31289;
  assign n31291 = n3318 & ~n30916;
  assign n31292 = ~n31290 & n31291;
  assign n31293 = n3003 & ~n3036;
  assign n31294 = ~pi39 & ~n31205;
  assign n31295 = ~n3048 & ~n31018;
  assign n31296 = ~n2953 & ~n31295;
  assign n31297 = n2953 & ~n3036;
  assign n31298 = ~n31296 & ~n31297;
  assign n31299 = ~n3050 & n31295;
  assign n31300 = ~n62393 & ~n64133;
  assign n31301 = ~n3057 & ~n31018;
  assign n31302 = ~n3057 & n31295;
  assign n31303 = n2909 & ~n31295;
  assign n31304 = ~n2909 & ~n3036;
  assign n31305 = ~n31303 & ~n31304;
  assign n31306 = ~n3048 & n31301;
  assign n31307 = n62393 & ~n64134;
  assign n31308 = n3056 & ~n31307;
  assign n31309 = n3056 & ~n31300;
  assign n31310 = ~n31307 & n31309;
  assign n31311 = ~n31300 & n31308;
  assign n31312 = n31238 & ~n64135;
  assign n31313 = ~n2971 & ~n64133;
  assign n31314 = n2971 & ~n64134;
  assign n31315 = n3076 & ~n31314;
  assign n31316 = n3076 & ~n31313;
  assign n31317 = ~n31314 & n31316;
  assign n31318 = ~n31313 & n31315;
  assign n31319 = ~pi299 & ~n3082;
  assign n31320 = ~n64136 & n31319;
  assign n31321 = ~n31312 & ~n31320;
  assign n31322 = pi39 & ~n31321;
  assign n31323 = ~pi38 & ~n31322;
  assign n31324 = ~n31294 & n31323;
  assign n31325 = ~pi100 & ~n3093;
  assign n31326 = ~n31324 & n31325;
  assign n31327 = ~n31293 & ~n31326;
  assign n31328 = ~pi87 & ~n31327;
  assign n31329 = ~n31012 & ~n31328;
  assign n31330 = ~pi75 & ~n31329;
  assign n31331 = n2817 & n31019;
  assign n31332 = ~n2817 & n3036;
  assign n31333 = pi75 & ~n31332;
  assign n31334 = ~n31331 & n31333;
  assign n31335 = ~n31330 & ~n31334;
  assign n31336 = n30915 & ~n31335;
  assign n31337 = ~n2580 & ~n31058;
  assign n31338 = ~n31336 & ~n31337;
  assign n31339 = ~n31292 & ~n31337;
  assign n31340 = ~n31336 & n31339;
  assign n31341 = ~n31292 & n31338;
  assign n31342 = pi120 & n31064;
  assign n31343 = ~n64137 & n31342;
  assign n31344 = ~n31282 & ~n31343;
  assign n31345 = ~n30913 & ~n31344;
  assign n31346 = ~n31073 & ~n31345;
  assign n31347 = ~pi149 & ~pi157;
  assign n31348 = pi197 & n31347;
  assign n31349 = ~pi197 & ~n31347;
  assign n31350 = ~n31348 & ~n31349;
  assign n31351 = pi162 & n2814;
  assign n31352 = n31350 & ~n31351;
  assign n31353 = n31348 & n31351;
  assign n31354 = n2814 & ~n31347;
  assign n31355 = ~pi162 & ~pi197;
  assign n31356 = n31354 & ~n31355;
  assign n31357 = n2814 & ~n31356;
  assign n31358 = ~n31353 & n31357;
  assign n31359 = ~n31350 & ~n31358;
  assign n31360 = ~n31352 & ~n31359;
  assign n31361 = pi232 & ~n2765;
  assign n31362 = pi232 & n31360;
  assign n31363 = ~n2765 & n31362;
  assign n31364 = n31360 & n31361;
  assign n31365 = pi167 & n2815;
  assign n31366 = n2765 & n2815;
  assign n31367 = pi167 & n31366;
  assign n31368 = n2765 & n31365;
  assign n31369 = ~n64138 & ~n64139;
  assign n31370 = ~pi74 & n31369;
  assign n31371 = pi148 & n31366;
  assign n31372 = pi74 & ~n31371;
  assign n31373 = ~n64138 & n31372;
  assign n31374 = ~n31370 & ~n31373;
  assign n31375 = ~n3472 & n31374;
  assign n31376 = ~pi54 & ~n64138;
  assign n31377 = pi38 & n31365;
  assign n31378 = n2765 & n31377;
  assign n31379 = pi38 & n64139;
  assign n31380 = n31376 & ~n64140;
  assign n31381 = ~pi74 & n31380;
  assign n31382 = n31374 & ~n31381;
  assign n31383 = ~n3470 & ~n31382;
  assign n31384 = n3472 & ~n31383;
  assign n31385 = ~pi40 & n2587;
  assign n31386 = ~pi38 & n31385;
  assign n31387 = n2765 & n31386;
  assign n31388 = n6792 & n31387;
  assign n31389 = ~n3470 & ~n31388;
  assign n31390 = n3472 & ~n31389;
  assign n31391 = ~n31384 & ~n31390;
  assign n31392 = pi299 & ~n31360;
  assign n31393 = ~pi178 & ~pi183;
  assign n31394 = pi140 & pi145;
  assign n31395 = n31393 & ~n31394;
  assign n31396 = ~pi140 & ~pi145;
  assign n31397 = n2814 & ~n31396;
  assign n31398 = n31395 & n31397;
  assign n31399 = n2814 & ~n31393;
  assign n31400 = ~n31394 & ~n31396;
  assign n31401 = n31399 & ~n31400;
  assign n31402 = ~pi299 & ~n31401;
  assign n31403 = ~pi299 & ~n31398;
  assign n31404 = ~n31401 & n31403;
  assign n31405 = ~n31398 & n31402;
  assign n31406 = pi232 & ~n64141;
  assign n31407 = ~n31392 & n31406;
  assign n31408 = pi100 & ~n31407;
  assign n31409 = pi75 & ~n31407;
  assign n31410 = ~n31408 & ~n31409;
  assign n31411 = pi141 & ~pi299;
  assign n31412 = pi148 & pi299;
  assign n31413 = ~n31411 & ~n31412;
  assign n31414 = n2815 & ~n31413;
  assign n31415 = n2765 & ~n31414;
  assign n31416 = n31410 & ~n31415;
  assign n31417 = pi74 & ~n31416;
  assign n31418 = ~pi55 & ~n31417;
  assign n31419 = pi188 & ~pi299;
  assign n31420 = pi167 & pi299;
  assign n31421 = ~pi167 & pi299;
  assign n31422 = ~pi188 & ~pi299;
  assign n31423 = ~n31421 & ~n31422;
  assign n31424 = ~n31419 & ~n31420;
  assign n31425 = n2815 & n64142;
  assign n31426 = ~pi100 & ~n31425;
  assign n31427 = ~pi75 & n31426;
  assign n31428 = n2765 & ~n31425;
  assign n31429 = n31410 & ~n64143;
  assign n31430 = pi54 & ~n31429;
  assign n31431 = pi95 & ~n31385;
  assign n31432 = ~n30613 & ~n31431;
  assign n31433 = ~pi40 & ~pi479;
  assign n31434 = n2682 & n62360;
  assign n31435 = ~pi53 & n31434;
  assign n31436 = n64091 & n31435;
  assign n31437 = ~pi58 & n31436;
  assign n31438 = n2695 & n31437;
  assign n31439 = ~pi32 & n62375;
  assign n31440 = n31438 & n31439;
  assign n31441 = n2587 & ~n31440;
  assign n31442 = n31433 & n31441;
  assign n31443 = ~n31432 & ~n31442;
  assign n31444 = pi32 & ~n31385;
  assign n31445 = n2587 & ~n2729;
  assign n31446 = n2587 & ~n31438;
  assign n31447 = pi70 & ~n31446;
  assign n31448 = n2587 & ~n31436;
  assign n31449 = pi58 & ~n31448;
  assign n31450 = pi50 & n2860;
  assign n31451 = ~pi60 & n31450;
  assign n31452 = n30639 & ~n31451;
  assign n31453 = pi53 & ~n64091;
  assign n31454 = ~n31452 & ~n31453;
  assign n31455 = ~pi111 & n2588;
  assign n31456 = ~pi68 & n2606;
  assign n31457 = ~pi36 & ~pi82;
  assign n31458 = ~pi82 & ~pi84;
  assign n31459 = ~pi36 & n31458;
  assign n31460 = ~pi84 & n31457;
  assign n31461 = n31456 & n64144;
  assign n31462 = n31455 & n64144;
  assign n31463 = n31456 & n31462;
  assign n31464 = n31455 & n31461;
  assign n31465 = ~pi66 & pi73;
  assign n31466 = n2620 & n31465;
  assign n31467 = n64145 & n31466;
  assign n31468 = ~pi36 & n31455;
  assign n31469 = ~pi36 & n31456;
  assign n31470 = n31455 & n31469;
  assign n31471 = n31456 & n31468;
  assign n31472 = pi73 & ~pi82;
  assign n31473 = n6804 & n31472;
  assign n31474 = n64146 & n31473;
  assign n31475 = n2624 & n31474;
  assign n31476 = n2624 & n31473;
  assign n31477 = n64146 & n31476;
  assign n31478 = n2627 & n31467;
  assign n31479 = n2596 & n64147;
  assign n31480 = n2637 & n31479;
  assign n31481 = n2587 & ~n31480;
  assign n31482 = ~n31454 & n31481;
  assign n31483 = n2682 & ~n31482;
  assign n31484 = ~n2587 & ~n2682;
  assign n31485 = n62360 & ~n31484;
  assign n31486 = ~n31483 & n31485;
  assign n31487 = n2587 & ~n62360;
  assign n31488 = ~pi58 & ~n31487;
  assign n31489 = ~n31486 & n31488;
  assign n31490 = ~n31449 & ~n31489;
  assign n31491 = ~pi90 & ~n31490;
  assign n31492 = ~pi841 & n31437;
  assign n31493 = n2587 & ~n31492;
  assign n31494 = pi90 & ~n31493;
  assign n31495 = n2719 & ~n31494;
  assign n31496 = ~n31491 & n31495;
  assign n31497 = n2587 & ~n2719;
  assign n31498 = ~pi70 & ~n31497;
  assign n31499 = ~n31496 & n31498;
  assign n31500 = ~n31447 & ~n31499;
  assign n31501 = ~pi51 & ~n31500;
  assign n31502 = pi51 & ~n2587;
  assign n31503 = n2729 & ~n31502;
  assign n31504 = ~n31501 & n31503;
  assign n31505 = ~n31445 & ~n31504;
  assign n31506 = ~pi40 & ~n31505;
  assign n31507 = ~pi32 & ~n31506;
  assign n31508 = ~n31444 & ~n31507;
  assign n31509 = ~pi95 & ~n31508;
  assign n31510 = ~n31443 & ~n31509;
  assign n31511 = ~pi198 & ~pi299;
  assign n31512 = ~pi210 & pi299;
  assign n31513 = pi210 & pi299;
  assign n31514 = pi198 & ~pi299;
  assign n31515 = ~n31513 & ~n31514;
  assign n31516 = ~n31511 & ~n31512;
  assign n31517 = n62768 & n31492;
  assign n31518 = n31385 & ~n31517;
  assign n31519 = pi32 & ~n31518;
  assign n31520 = ~n31507 & ~n31519;
  assign n31521 = ~pi95 & ~n31520;
  assign n31522 = n64148 & n31521;
  assign n31523 = n31510 & ~n31522;
  assign n31524 = ~pi232 & ~n31523;
  assign n31525 = ~pi198 & n31521;
  assign n31526 = n31510 & ~n31525;
  assign n31527 = ~n2814 & n31526;
  assign n31528 = ~pi40 & ~n2587;
  assign n31529 = pi32 & ~n31528;
  assign n31530 = ~n2587 & ~n2720;
  assign n31531 = n2695 & n31489;
  assign n31532 = ~n31530 & ~n31531;
  assign n31533 = ~pi70 & ~n31532;
  assign n31534 = ~n31447 & ~n31533;
  assign n31535 = ~pi51 & ~n31534;
  assign n31536 = n31503 & ~n31535;
  assign n31537 = ~pi40 & ~n31445;
  assign n31538 = ~n31536 & n31537;
  assign n31539 = ~pi32 & ~n31538;
  assign n31540 = ~n31529 & ~n31539;
  assign n31541 = ~n2730 & ~n31385;
  assign n31542 = ~n31540 & ~n31541;
  assign n31543 = ~pi95 & ~n31542;
  assign n31544 = ~n31443 & ~n31543;
  assign n31545 = n2814 & ~n31385;
  assign n31546 = ~n31431 & ~n31543;
  assign n31547 = pi95 & ~n31528;
  assign n31548 = ~pi40 & ~n31518;
  assign n31549 = pi32 & ~n31548;
  assign n31550 = ~n31539 & ~n31549;
  assign n31551 = ~pi95 & ~n31550;
  assign n31552 = ~n31547 & ~n31551;
  assign n31553 = n31546 & ~n31552;
  assign n31554 = ~pi198 & ~n31553;
  assign n31555 = n2814 & ~n31554;
  assign n31556 = ~n31545 & ~n31555;
  assign n31557 = n31544 & ~n31556;
  assign n31558 = ~n31527 & ~n31557;
  assign n31559 = ~pi142 & ~n31558;
  assign n31560 = pi142 & n31526;
  assign n31561 = ~pi140 & ~n31560;
  assign n31562 = ~n31559 & n31561;
  assign n31563 = ~pi32 & n62775;
  assign n31564 = n31479 & n31563;
  assign n31565 = n31385 & ~n31564;
  assign n31566 = ~pi95 & ~n31565;
  assign n31567 = n2814 & ~n31566;
  assign n31568 = ~n31443 & n31567;
  assign n31569 = ~n31527 & ~n31568;
  assign n31570 = ~pi142 & ~n31569;
  assign n31571 = ~n2814 & ~n31526;
  assign n31572 = ~pi40 & ~n31444;
  assign n31573 = n2587 & ~n62382;
  assign n31574 = ~pi32 & ~n31573;
  assign n31575 = pi93 & ~n2587;
  assign n31576 = n62382 & ~n31575;
  assign n31577 = n2587 & ~n31449;
  assign n31578 = ~pi90 & ~n31577;
  assign n31579 = ~n31494 & ~n31578;
  assign n31580 = n62356 & n31479;
  assign n31581 = ~pi90 & n31580;
  assign n31582 = n31579 & ~n31581;
  assign n31583 = ~pi93 & ~n31582;
  assign n31584 = n31576 & ~n31583;
  assign n31585 = n31574 & ~n31584;
  assign n31586 = n31572 & ~n31585;
  assign n31587 = ~pi95 & ~n31586;
  assign n31588 = ~n31443 & ~n31587;
  assign n31589 = n2814 & ~n31588;
  assign n31590 = pi142 & ~n31589;
  assign n31591 = ~n31571 & n31590;
  assign n31592 = pi140 & ~n31591;
  assign n31593 = ~n31570 & n31592;
  assign n31594 = ~n31562 & ~n31593;
  assign n31595 = ~pi181 & ~n31594;
  assign n31596 = n2814 & ~n31431;
  assign n31597 = ~n31566 & n31596;
  assign n31598 = ~n31527 & ~n31597;
  assign n31599 = ~pi142 & ~n31598;
  assign n31600 = ~n31587 & n31596;
  assign n31601 = ~n31527 & ~n31600;
  assign n31602 = pi142 & ~n31601;
  assign n31603 = pi140 & ~n31602;
  assign n31604 = pi140 & ~n31599;
  assign n31605 = ~n31602 & n31604;
  assign n31606 = ~n31599 & n31603;
  assign n31607 = n31546 & n31555;
  assign n31608 = ~n31527 & ~n31607;
  assign n31609 = ~pi142 & ~n31608;
  assign n31610 = ~pi40 & n2814;
  assign n31611 = ~n31431 & ~n31509;
  assign n31612 = ~n31525 & n31611;
  assign n31613 = n31610 & n31612;
  assign n31614 = ~n31527 & ~n31613;
  assign n31615 = pi142 & ~n31614;
  assign n31616 = ~pi140 & ~n31615;
  assign n31617 = ~n31609 & n31616;
  assign n31618 = ~n64149 & ~n31617;
  assign n31619 = pi181 & ~n31618;
  assign n31620 = pi144 & ~n31619;
  assign n31621 = ~n31595 & n31620;
  assign n31622 = ~pi93 & ~n31579;
  assign n31623 = n31576 & ~n31622;
  assign n31624 = n31574 & ~n31623;
  assign n31625 = n31572 & ~n31624;
  assign n31626 = ~pi95 & ~n31625;
  assign n31627 = n31596 & ~n31626;
  assign n31628 = ~n31527 & ~n31627;
  assign n31629 = pi142 & ~n31628;
  assign n31630 = ~n31545 & ~n31571;
  assign n31631 = ~pi142 & n31630;
  assign n31632 = pi140 & ~n31631;
  assign n31633 = pi140 & ~n31629;
  assign n31634 = ~n31631 & n31633;
  assign n31635 = ~n31629 & n31632;
  assign n31636 = n31434 & n31454;
  assign n31637 = n2587 & ~n31636;
  assign n31638 = ~pi58 & ~n31637;
  assign n31639 = n2695 & n31638;
  assign n31640 = ~n31530 & ~n31639;
  assign n31641 = ~pi70 & ~n31640;
  assign n31642 = ~n31447 & ~n31641;
  assign n31643 = ~pi51 & ~n31642;
  assign n31644 = n31503 & ~n31643;
  assign n31645 = ~n31445 & ~n31644;
  assign n31646 = ~pi40 & n31645;
  assign n31647 = ~pi32 & ~n31646;
  assign n31648 = ~n31529 & ~n31647;
  assign n31649 = ~pi95 & ~n31648;
  assign n31650 = pi198 & n31649;
  assign n31651 = ~n31549 & ~n31647;
  assign n31652 = ~pi95 & ~n31651;
  assign n31653 = ~pi198 & n31652;
  assign n31654 = ~n31547 & ~n31653;
  assign n31655 = ~n31547 & ~n31649;
  assign n31656 = pi198 & ~n31655;
  assign n31657 = ~n31547 & ~n31652;
  assign n31658 = ~pi198 & ~n31657;
  assign n31659 = ~n31656 & ~n31658;
  assign n31660 = ~n31650 & n31654;
  assign n31661 = n31610 & ~n64151;
  assign n31662 = ~n31527 & ~n31661;
  assign n31663 = ~pi142 & ~n31662;
  assign n31664 = ~n31449 & ~n31638;
  assign n31665 = ~pi90 & ~n31664;
  assign n31666 = n31495 & ~n31665;
  assign n31667 = n31498 & ~n31666;
  assign n31668 = ~n31447 & ~n31667;
  assign n31669 = ~pi51 & ~n31668;
  assign n31670 = n31503 & ~n31669;
  assign n31671 = ~n31445 & ~n31670;
  assign n31672 = ~pi40 & ~n31671;
  assign n31673 = ~pi32 & ~n31672;
  assign n31674 = ~n31444 & ~n31673;
  assign n31675 = ~pi95 & ~n31674;
  assign n31676 = n31596 & ~n31675;
  assign n31677 = ~n31519 & ~n31673;
  assign n31678 = ~pi95 & ~n31677;
  assign n31679 = ~pi198 & n31678;
  assign n31680 = n31676 & ~n31679;
  assign n31681 = ~n31527 & ~n31680;
  assign n31682 = pi142 & ~n31681;
  assign n31683 = ~pi140 & ~n31682;
  assign n31684 = ~pi140 & ~n31663;
  assign n31685 = ~n31682 & n31684;
  assign n31686 = ~n31663 & n31683;
  assign n31687 = ~n64150 & ~n64152;
  assign n31688 = pi181 & ~n31687;
  assign n31689 = ~pi40 & ~n31645;
  assign n31690 = ~pi32 & ~n31689;
  assign n31691 = ~n31444 & ~n31690;
  assign n31692 = ~pi95 & ~n31691;
  assign n31693 = ~n31443 & ~n31692;
  assign n31694 = ~n31519 & ~n31690;
  assign n31695 = ~pi95 & ~n31694;
  assign n31696 = ~pi198 & n31695;
  assign n31697 = n31693 & ~n31696;
  assign n31698 = n2814 & ~n31697;
  assign n31699 = ~n31571 & ~n31698;
  assign n31700 = ~pi142 & n31699;
  assign n31701 = ~n31443 & ~n31675;
  assign n31702 = ~n31679 & n31701;
  assign n31703 = n2814 & ~n31702;
  assign n31704 = pi142 & ~n31703;
  assign n31705 = ~n31571 & n31704;
  assign n31706 = ~pi140 & ~n31705;
  assign n31707 = ~n31700 & n31706;
  assign n31708 = ~pi95 & ~n31385;
  assign n31709 = ~n31443 & ~n31708;
  assign n31710 = n2814 & n31709;
  assign n31711 = ~n31527 & ~n31710;
  assign n31712 = ~pi142 & ~n31711;
  assign n31713 = ~n31443 & ~n31626;
  assign n31714 = n2814 & ~n31713;
  assign n31715 = pi142 & ~n31714;
  assign n31716 = ~n31571 & n31715;
  assign n31717 = pi140 & ~n31716;
  assign n31718 = ~n31712 & n31717;
  assign n31719 = ~n31707 & ~n31718;
  assign n31720 = ~pi181 & ~n31719;
  assign n31721 = ~pi144 & ~n31720;
  assign n31722 = ~n31688 & n31721;
  assign n31723 = ~pi299 & ~n31722;
  assign n31724 = ~pi181 & ~n31593;
  assign n31725 = ~n31562 & n31724;
  assign n31726 = pi181 & ~n31617;
  assign n31727 = pi181 & ~n64149;
  assign n31728 = ~n31617 & n31727;
  assign n31729 = ~n64149 & n31726;
  assign n31730 = pi144 & ~n64153;
  assign n31731 = ~n31725 & n31730;
  assign n31732 = pi181 & ~n64152;
  assign n31733 = ~n64150 & n31732;
  assign n31734 = ~pi140 & ~n31702;
  assign n31735 = pi140 & ~n31713;
  assign n31736 = pi142 & ~n31735;
  assign n31737 = ~n31734 & n31736;
  assign n31738 = ~pi140 & ~n31697;
  assign n31739 = pi140 & ~n31709;
  assign n31740 = ~pi142 & ~n31739;
  assign n31741 = ~n31738 & n31740;
  assign n31742 = n2814 & ~n31741;
  assign n31743 = ~pi140 & n31702;
  assign n31744 = pi140 & n31713;
  assign n31745 = pi142 & ~n31744;
  assign n31746 = ~n31743 & n31745;
  assign n31747 = ~pi140 & n31697;
  assign n31748 = pi140 & n31709;
  assign n31749 = ~pi142 & ~n31748;
  assign n31750 = ~n31747 & n31749;
  assign n31751 = ~n31746 & ~n31750;
  assign n31752 = n2814 & ~n31751;
  assign n31753 = ~n31737 & n31742;
  assign n31754 = ~pi181 & ~n31571;
  assign n31755 = ~n64154 & n31754;
  assign n31756 = ~pi144 & ~n31755;
  assign n31757 = ~n31733 & n31756;
  assign n31758 = ~n31731 & ~n31757;
  assign n31759 = ~pi299 & ~n31758;
  assign n31760 = ~n31621 & n31723;
  assign n31761 = pi159 & pi299;
  assign n31762 = ~pi210 & n31521;
  assign n31763 = n31510 & ~n31762;
  assign n31764 = ~n2814 & n31763;
  assign n31765 = ~n31600 & ~n31764;
  assign n31766 = pi146 & ~n31765;
  assign n31767 = ~n31597 & ~n31764;
  assign n31768 = ~pi146 & ~n31767;
  assign n31769 = pi161 & ~n31768;
  assign n31770 = pi161 & ~n31766;
  assign n31771 = ~n31768 & n31770;
  assign n31772 = ~n31766 & n31769;
  assign n31773 = ~n31627 & ~n31764;
  assign n31774 = pi146 & ~n31773;
  assign n31775 = ~n2814 & ~n31763;
  assign n31776 = ~n31545 & ~n31775;
  assign n31777 = ~pi146 & n31776;
  assign n31778 = ~pi161 & ~n31777;
  assign n31779 = ~pi161 & ~n31774;
  assign n31780 = ~n31777 & n31779;
  assign n31781 = ~n31774 & n31778;
  assign n31782 = ~n64156 & ~n64157;
  assign n31783 = n31761 & ~n31782;
  assign n31784 = ~pi159 & pi299;
  assign n31785 = ~n31568 & ~n31764;
  assign n31786 = ~pi146 & ~n31785;
  assign n31787 = ~n31589 & ~n31775;
  assign n31788 = pi146 & n31787;
  assign n31789 = pi161 & ~n31788;
  assign n31790 = pi161 & ~n31786;
  assign n31791 = ~n31788 & n31790;
  assign n31792 = ~n31786 & n31789;
  assign n31793 = ~n31714 & ~n31775;
  assign n31794 = pi146 & n31793;
  assign n31795 = ~n31710 & ~n31764;
  assign n31796 = ~pi146 & ~n31795;
  assign n31797 = ~pi161 & ~n31796;
  assign n31798 = ~pi161 & ~n31794;
  assign n31799 = ~n31796 & n31798;
  assign n31800 = ~n31794 & n31797;
  assign n31801 = ~n64158 & ~n64159;
  assign n31802 = n31784 & ~n31801;
  assign n31803 = ~n31783 & ~n31802;
  assign n31804 = pi162 & ~n31803;
  assign n31805 = ~pi210 & n31678;
  assign n31806 = n31676 & ~n31805;
  assign n31807 = ~n31764 & ~n31806;
  assign n31808 = pi146 & ~n31807;
  assign n31809 = ~n31431 & ~n31695;
  assign n31810 = ~pi210 & ~n31809;
  assign n31811 = n2814 & ~n31810;
  assign n31812 = ~n31431 & ~n31692;
  assign n31813 = n31811 & n31812;
  assign n31814 = ~n31764 & ~n31813;
  assign n31815 = ~pi146 & ~n31814;
  assign n31816 = ~pi161 & ~n31815;
  assign n31817 = ~pi161 & ~n31808;
  assign n31818 = ~n31815 & n31817;
  assign n31819 = ~n31808 & n31816;
  assign n31820 = ~pi210 & ~n31553;
  assign n31821 = n2814 & ~n31820;
  assign n31822 = n31546 & n31821;
  assign n31823 = ~n31764 & ~n31822;
  assign n31824 = ~pi146 & ~n31823;
  assign n31825 = n31611 & ~n31762;
  assign n31826 = n2814 & ~n31825;
  assign n31827 = ~n31775 & ~n31826;
  assign n31828 = pi146 & n31827;
  assign n31829 = pi161 & ~n31828;
  assign n31830 = ~n31824 & n31829;
  assign n31831 = ~n64160 & ~n31830;
  assign n31832 = n31761 & ~n31831;
  assign n31833 = ~n31545 & ~n31821;
  assign n31834 = n31544 & ~n31833;
  assign n31835 = pi161 & n31834;
  assign n31836 = ~n31545 & ~n31811;
  assign n31837 = n31693 & ~n31836;
  assign n31838 = ~pi161 & n31837;
  assign n31839 = ~pi146 & ~n31838;
  assign n31840 = ~n31835 & n31839;
  assign n31841 = pi161 & n31763;
  assign n31842 = n31701 & ~n31805;
  assign n31843 = n2814 & n31842;
  assign n31844 = ~pi161 & n31843;
  assign n31845 = pi146 & ~n31844;
  assign n31846 = ~n31841 & n31845;
  assign n31847 = ~n31840 & ~n31846;
  assign n31848 = ~n31764 & n31784;
  assign n31849 = ~n31847 & n31848;
  assign n31850 = ~n31832 & ~n31849;
  assign n31851 = ~pi162 & ~n31850;
  assign n31852 = pi162 & ~n31801;
  assign n31853 = pi161 & ~n31834;
  assign n31854 = ~pi161 & ~n31837;
  assign n31855 = ~pi146 & ~n31854;
  assign n31856 = ~n31853 & n31855;
  assign n31857 = ~pi161 & ~n31843;
  assign n31858 = pi161 & ~n31763;
  assign n31859 = pi146 & ~n31858;
  assign n31860 = pi146 & ~n31857;
  assign n31861 = ~n31858 & n31860;
  assign n31862 = ~n31857 & n31859;
  assign n31863 = ~pi162 & ~n31764;
  assign n31864 = ~n64161 & n31863;
  assign n31865 = ~n31856 & n31864;
  assign n31866 = ~n31852 & ~n31865;
  assign n31867 = n31784 & ~n31866;
  assign n31868 = ~pi162 & ~n64160;
  assign n31869 = ~pi162 & ~n31830;
  assign n31870 = ~n64160 & n31869;
  assign n31871 = ~n31830 & n31868;
  assign n31872 = pi162 & ~n64156;
  assign n31873 = pi162 & ~n64157;
  assign n31874 = ~n64156 & n31873;
  assign n31875 = ~n64157 & n31872;
  assign n31876 = n31761 & ~n64163;
  assign n31877 = n31761 & ~n64162;
  assign n31878 = ~n64163 & n31877;
  assign n31879 = ~n64162 & n31876;
  assign n31880 = ~n31867 & ~n64164;
  assign n31881 = ~n31804 & ~n31851;
  assign n31882 = ~n64155 & n64165;
  assign n31883 = pi232 & ~n31882;
  assign n31884 = ~n31524 & ~n31883;
  assign n31885 = n2764 & ~n31884;
  assign n31886 = pi216 & n2960;
  assign n31887 = ~pi95 & n31440;
  assign n31888 = n62395 & n6958;
  assign n31889 = pi1092 & n6958;
  assign n31890 = n3322 & ~n30823;
  assign n31891 = n31889 & n31890;
  assign n31892 = ~n31888 & ~n31891;
  assign n31893 = n31887 & ~n31892;
  assign n31894 = n2909 & n31893;
  assign n31895 = n31385 & ~n31894;
  assign n31896 = n2814 & n31893;
  assign n31897 = n31385 & ~n31896;
  assign n31898 = ~n62393 & ~n31897;
  assign n31899 = n31895 & ~n31898;
  assign n31900 = n31887 & n31888;
  assign n31901 = ~n2953 & n31900;
  assign n31902 = n31385 & ~n31901;
  assign n31903 = n2814 & n31902;
  assign n31904 = ~pi161 & n31903;
  assign n31905 = ~n31899 & ~n31904;
  assign n31906 = n31886 & ~n31905;
  assign n31907 = n31385 & ~n31886;
  assign n31908 = pi299 & ~n31907;
  assign n31909 = ~pi38 & ~pi155;
  assign n31910 = n31908 & n31909;
  assign n31911 = ~n31906 & n31910;
  assign n31912 = n31887 & n31891;
  assign n31913 = n31385 & ~n31912;
  assign n31914 = n2919 & ~n31913;
  assign n31915 = pi161 & n31914;
  assign n31916 = n31886 & n31895;
  assign n31917 = ~n31915 & n31916;
  assign n31918 = ~pi38 & pi155;
  assign n31919 = n31908 & n31918;
  assign n31920 = ~n31917 & n31919;
  assign n31921 = ~n31906 & n31909;
  assign n31922 = ~n31917 & n31918;
  assign n31923 = ~n31921 & ~n31922;
  assign n31924 = n31908 & ~n31923;
  assign n31925 = ~n31911 & ~n31920;
  assign n31926 = pi224 & n2980;
  assign n31927 = n31385 & ~n31926;
  assign n31928 = ~n31895 & ~n31927;
  assign n31929 = ~n2971 & ~n31897;
  assign n31930 = ~n31927 & n31929;
  assign n31931 = n31895 & ~n31929;
  assign n31932 = ~n31927 & ~n31931;
  assign n31933 = ~n31928 & ~n31930;
  assign n31934 = pi144 & ~n64167;
  assign n31935 = ~pi177 & ~pi299;
  assign n31936 = n2972 & n31900;
  assign n31937 = n31385 & n31926;
  assign n31938 = ~n31936 & n31937;
  assign n31939 = ~n31927 & ~n31938;
  assign n31940 = ~pi144 & ~n31928;
  assign n31941 = ~n31939 & n31940;
  assign n31942 = n31935 & ~n31941;
  assign n31943 = ~n31934 & n31942;
  assign n31944 = n2814 & n31926;
  assign n31945 = n31912 & n31944;
  assign n31946 = n31385 & ~n31945;
  assign n31947 = n2814 & n31912;
  assign n31948 = n31385 & ~n31947;
  assign n31949 = ~n2971 & ~n31948;
  assign n31950 = ~n31927 & n31949;
  assign n31951 = ~n2971 & ~n31946;
  assign n31952 = ~n31928 & ~n64168;
  assign n31953 = ~pi299 & ~n31952;
  assign n31954 = pi177 & ~n31940;
  assign n31955 = pi177 & ~pi299;
  assign n31956 = ~n31940 & n31955;
  assign n31957 = ~n31952 & n31956;
  assign n31958 = n31953 & n31954;
  assign n31959 = ~n31943 & ~n64169;
  assign n31960 = ~pi38 & ~n31959;
  assign n31961 = ~n64166 & ~n31960;
  assign n31962 = pi232 & ~n31961;
  assign n31963 = ~n31899 & n31908;
  assign n31964 = ~pi299 & n64167;
  assign n31965 = ~n31963 & ~n31964;
  assign n31966 = ~pi232 & ~n31965;
  assign n31967 = ~pi38 & n31966;
  assign n31968 = pi232 & ~n31959;
  assign n31969 = ~n31966 & ~n31968;
  assign n31970 = ~pi38 & ~n31969;
  assign n31971 = pi232 & n31908;
  assign n31972 = ~n31923 & n31971;
  assign n31973 = pi232 & n64166;
  assign n31974 = ~n31970 & ~n64170;
  assign n31975 = ~n31962 & ~n31967;
  assign n31976 = pi39 & ~n64171;
  assign n31977 = ~pi299 & n2815;
  assign n31978 = ~n7356 & n31977;
  assign n31979 = ~pi167 & ~n31978;
  assign n31980 = n2815 & ~n7356;
  assign n31981 = pi167 & ~n31980;
  assign n31982 = pi188 & ~n31981;
  assign n31983 = ~n31979 & n31982;
  assign n31984 = pi299 & ~n7356;
  assign n31985 = ~pi188 & n31365;
  assign n31986 = n31984 & n31985;
  assign n31987 = pi38 & ~n31986;
  assign n31988 = pi188 & n31978;
  assign n31989 = ~pi167 & ~n31988;
  assign n31990 = pi299 & n2815;
  assign n31991 = n2815 & n31984;
  assign n31992 = ~n7356 & n31990;
  assign n31993 = ~pi188 & ~n64172;
  assign n31994 = pi167 & pi188;
  assign n31995 = ~n31980 & n31994;
  assign n31996 = ~n31993 & ~n31995;
  assign n31997 = pi188 & ~n31979;
  assign n31998 = pi167 & n64172;
  assign n31999 = ~n31997 & ~n31998;
  assign n32000 = ~n31995 & ~n31999;
  assign n32001 = ~n31989 & n31996;
  assign n32002 = pi38 & ~n64173;
  assign n32003 = ~n31983 & n31987;
  assign n32004 = ~pi87 & ~n64174;
  assign n32005 = ~n31976 & n32004;
  assign n32006 = ~n31885 & n32005;
  assign n32007 = pi38 & n64142;
  assign n32008 = n2815 & n32007;
  assign n32009 = ~pi38 & ~n31385;
  assign n32010 = pi38 & ~n31425;
  assign n32011 = ~n32009 & ~n32010;
  assign n32012 = ~n31386 & ~n32008;
  assign n32013 = pi87 & n64175;
  assign n32014 = ~pi100 & ~n32013;
  assign n32015 = ~n32006 & n32014;
  assign n32016 = ~n31408 & ~n32015;
  assign n32017 = n6793 & ~n32016;
  assign n32018 = ~pi75 & pi92;
  assign n32019 = ~pi39 & ~pi95;
  assign n32020 = ~pi87 & n32019;
  assign n32021 = n2805 & n31887;
  assign n32022 = n31440 & n32020;
  assign n32023 = pi155 & pi299;
  assign n32024 = ~pi155 & pi299;
  assign n32025 = ~n31935 & ~n32024;
  assign n32026 = ~n31955 & ~n32023;
  assign n32027 = ~pi38 & ~n64177;
  assign n32028 = n2815 & ~n32027;
  assign n32029 = n64176 & ~n32028;
  assign n32030 = n64175 & ~n32029;
  assign n32031 = ~pi100 & ~n32030;
  assign n32032 = ~n31408 & ~n32031;
  assign n32033 = n32018 & ~n32032;
  assign n32034 = ~n31409 & ~n32033;
  assign n32035 = ~n32017 & n32034;
  assign n32036 = ~pi54 & ~n32035;
  assign n32037 = ~n31430 & ~n32036;
  assign n32038 = ~pi74 & ~n32037;
  assign n32039 = n31418 & ~n32038;
  assign n32040 = pi55 & ~n31373;
  assign n32041 = pi54 & n31369;
  assign n32042 = n31380 & ~n31387;
  assign n32043 = ~n2579 & ~n32042;
  assign n32044 = ~n2765 & n31360;
  assign n32045 = n31351 & n31387;
  assign n32046 = ~n32044 & ~n32045;
  assign n32047 = pi232 & ~n32046;
  assign n32048 = n31386 & ~n64176;
  assign n32049 = ~n31377 & ~n32048;
  assign n32050 = n2765 & ~n32049;
  assign n32051 = ~n32047 & ~n32050;
  assign n32052 = pi100 & ~n31362;
  assign n32053 = ~n31351 & n64176;
  assign n32054 = n31386 & ~n32053;
  assign n32055 = ~pi100 & ~n32054;
  assign n32056 = ~pi232 & n64176;
  assign n32057 = ~n32055 & ~n32056;
  assign n32058 = ~n31377 & ~n32057;
  assign n32059 = ~n32052 & ~n32058;
  assign n32060 = ~pi75 & ~n32059;
  assign n32061 = pi75 & ~n31362;
  assign n32062 = ~pi92 & ~n32061;
  assign n32063 = ~n32060 & n32062;
  assign n32064 = ~pi92 & ~n32051;
  assign n32065 = ~n32043 & ~n64178;
  assign n32066 = ~n32041 & ~n32065;
  assign n32067 = ~pi74 & ~n32066;
  assign n32068 = n32040 & ~n32067;
  assign n32069 = n3470 & ~n32068;
  assign n32070 = ~n32039 & n32069;
  assign n32071 = ~n31391 & ~n32070;
  assign n32072 = ~n31375 & ~n32071;
  assign n32073 = ~pi34 & n32072;
  assign n32074 = pi159 & n30614;
  assign n32075 = n2728 & n64090;
  assign n32076 = pi58 & n2658;
  assign n32077 = ~pi90 & ~n32076;
  assign n32078 = pi90 & ~n2674;
  assign n32079 = n2719 & ~n32078;
  assign n32080 = ~n32077 & ~n32078;
  assign n32081 = n2719 & n32080;
  assign n32082 = n2719 & ~n32077;
  assign n32083 = ~n32078 & n32082;
  assign n32084 = ~n32077 & n32079;
  assign n32085 = n2682 & ~n30637;
  assign n32086 = n2710 & n2719;
  assign n32087 = n32085 & n32086;
  assign n32088 = n2587 & n32087;
  assign n32089 = n31483 & n32088;
  assign n32090 = ~pi70 & ~n32089;
  assign n32091 = ~n64179 & n32090;
  assign n32092 = n32075 & ~n32091;
  assign n32093 = ~pi146 & n32092;
  assign n32094 = n32075 & ~n32090;
  assign n32095 = ~n30775 & ~n32094;
  assign n32096 = ~pi161 & n32095;
  assign n32097 = ~n32093 & n32096;
  assign n32098 = ~n31452 & n32087;
  assign n32099 = ~pi70 & ~n32098;
  assign n32100 = ~n64179 & n32099;
  assign n32101 = n32075 & ~n32100;
  assign n32102 = ~pi146 & n32101;
  assign n32103 = n32075 & ~n32099;
  assign n32104 = ~n30775 & ~n32103;
  assign n32105 = pi161 & n32104;
  assign n32106 = ~n32102 & n32105;
  assign n32107 = pi162 & ~n32106;
  assign n32108 = ~n32097 & n32107;
  assign n32109 = ~n32074 & ~n32108;
  assign n32110 = n2814 & ~n32109;
  assign n32111 = n2727 & n2814;
  assign n32112 = ~pi40 & n32111;
  assign n32113 = n62769 & ~n32078;
  assign n32114 = n2587 & n31580;
  assign n32115 = n32077 & ~n32114;
  assign n32116 = n32113 & ~n32115;
  assign n32117 = n32112 & n32116;
  assign n32118 = ~pi146 & ~n32117;
  assign n32119 = n62768 & n32114;
  assign n32120 = n2727 & n32119;
  assign n32121 = n31610 & n32120;
  assign n32122 = pi146 & ~n32121;
  assign n32123 = ~pi161 & ~n32122;
  assign n32124 = ~n32118 & n32123;
  assign n32125 = n62769 & n32080;
  assign n32126 = ~n32077 & n32113;
  assign n32127 = n32112 & n64180;
  assign n32128 = ~pi146 & pi161;
  assign n32129 = n32127 & n32128;
  assign n32130 = ~n32124 & ~n32129;
  assign n32131 = ~pi162 & ~n32130;
  assign n32132 = pi299 & ~n32131;
  assign n32133 = ~pi162 & ~n32074;
  assign n32134 = n2814 & ~n32133;
  assign n32135 = n2814 & n30614;
  assign n32136 = ~pi162 & n32135;
  assign n32137 = n31761 & ~n32136;
  assign n32138 = ~n31784 & ~n32137;
  assign n32139 = ~n31351 & ~n32138;
  assign n32140 = pi299 & ~n32134;
  assign n32141 = ~n32093 & n32095;
  assign n32142 = ~pi161 & ~n32141;
  assign n32143 = ~n32102 & n32104;
  assign n32144 = pi161 & ~n32143;
  assign n32145 = pi299 & ~n32074;
  assign n32146 = ~n32144 & n32145;
  assign n32147 = ~n32142 & n32146;
  assign n32148 = ~n64181 & ~n32147;
  assign n32149 = ~n32131 & ~n32148;
  assign n32150 = ~n32110 & n32132;
  assign n32151 = ~pi142 & n32092;
  assign n32152 = ~n30612 & ~n32094;
  assign n32153 = ~pi144 & n32152;
  assign n32154 = ~n32151 & n32153;
  assign n32155 = ~pi142 & n32101;
  assign n32156 = ~n30612 & ~n32103;
  assign n32157 = pi144 & n32156;
  assign n32158 = ~n32155 & n32157;
  assign n32159 = pi140 & n2814;
  assign n32160 = ~n32158 & n32159;
  assign n32161 = ~n32154 & n32160;
  assign n32162 = ~pi142 & ~n32117;
  assign n32163 = pi142 & ~n32121;
  assign n32164 = ~pi144 & ~n32163;
  assign n32165 = ~n32162 & n32164;
  assign n32166 = ~pi142 & pi144;
  assign n32167 = n32127 & n32166;
  assign n32168 = ~n32165 & ~n32167;
  assign n32169 = ~pi140 & ~n32168;
  assign n32170 = pi181 & n32135;
  assign n32171 = ~pi299 & ~n32170;
  assign n32172 = ~n32169 & n32171;
  assign n32173 = ~pi142 & n32117;
  assign n32174 = pi142 & n32121;
  assign n32175 = ~pi140 & ~n32174;
  assign n32176 = ~n32173 & n32175;
  assign n32177 = pi140 & n32152;
  assign n32178 = ~n32151 & n32177;
  assign n32179 = ~n32176 & ~n32178;
  assign n32180 = ~pi144 & ~n32179;
  assign n32181 = pi140 & ~n2814;
  assign n32182 = ~pi142 & n32127;
  assign n32183 = ~pi140 & ~n32182;
  assign n32184 = pi140 & ~n32155;
  assign n32185 = n32156 & n32184;
  assign n32186 = ~n32183 & ~n32185;
  assign n32187 = ~n32155 & n32156;
  assign n32188 = pi140 & ~n32187;
  assign n32189 = pi144 & ~n32188;
  assign n32190 = ~n32182 & n32189;
  assign n32191 = pi144 & ~n32186;
  assign n32192 = n2814 & ~n32189;
  assign n32193 = pi140 & ~n32192;
  assign n32194 = ~n64183 & ~n32193;
  assign n32195 = ~n32181 & ~n64183;
  assign n32196 = ~n32180 & n64184;
  assign n32197 = n32171 & ~n32196;
  assign n32198 = ~n32161 & n32172;
  assign n32199 = pi232 & ~n64185;
  assign n32200 = pi232 & ~n64182;
  assign n32201 = ~n64185 & n32200;
  assign n32202 = ~n64182 & n32199;
  assign n32203 = n2764 & ~n64186;
  assign n32204 = n2919 & ~n30820;
  assign n32205 = ~pi161 & ~n32204;
  assign n32206 = n2814 & n62397;
  assign n32207 = ~n62393 & n32206;
  assign n32208 = n2919 & n62397;
  assign n32209 = pi161 & ~n64187;
  assign n32210 = n31886 & ~n32209;
  assign n32211 = n31886 & ~n32205;
  assign n32212 = ~n32209 & n32211;
  assign n32213 = ~n32205 & n32210;
  assign n32214 = n31918 & ~n64188;
  assign n32215 = n2919 & n30824;
  assign n32216 = ~pi161 & n31886;
  assign n32217 = n32215 & n32216;
  assign n32218 = n31909 & ~n32217;
  assign n32219 = ~n32214 & ~n32218;
  assign n32220 = pi299 & ~n32219;
  assign n32221 = ~n2971 & n31926;
  assign n32222 = n2814 & n32221;
  assign n32223 = n2972 & n31926;
  assign n32224 = ~n30820 & n31926;
  assign n32225 = n2972 & n32224;
  assign n32226 = ~n30820 & n64189;
  assign n32227 = ~pi144 & n64190;
  assign n32228 = n62397 & n64189;
  assign n32229 = pi144 & n32228;
  assign n32230 = n31955 & ~n32229;
  assign n32231 = n31955 & ~n32227;
  assign n32232 = ~n32229 & n32231;
  assign n32233 = ~n32227 & n32230;
  assign n32234 = n2972 & n30824;
  assign n32235 = n31926 & n32234;
  assign n32236 = n30824 & n64189;
  assign n32237 = ~pi144 & n64192;
  assign n32238 = n31935 & ~n32237;
  assign n32239 = pi232 & ~n32238;
  assign n32240 = ~n64191 & n32239;
  assign n32241 = ~pi38 & ~n32240;
  assign n32242 = ~n32220 & ~n32241;
  assign n32243 = pi39 & ~n32242;
  assign n32244 = ~n64174 & ~n32243;
  assign n32245 = ~n32203 & n32244;
  assign n32246 = ~pi100 & ~n32245;
  assign n32247 = ~n31408 & ~n32246;
  assign n32248 = ~pi87 & ~n32247;
  assign n32249 = ~n2766 & ~n31426;
  assign n32250 = ~pi100 & ~n32008;
  assign n32251 = ~n31408 & n64193;
  assign n32252 = pi87 & ~n32251;
  assign n32253 = ~n32248 & ~n32252;
  assign n32254 = n6793 & ~n32253;
  assign n32255 = n2764 & n64177;
  assign n32256 = n62380 & n32255;
  assign n32257 = ~n32007 & ~n32256;
  assign n32258 = n2815 & ~n32257;
  assign n32259 = ~pi100 & ~n32258;
  assign n32260 = ~n31408 & ~n32259;
  assign n32261 = ~pi87 & ~n32260;
  assign n32262 = ~n32252 & ~n32261;
  assign n32263 = n32018 & ~n32262;
  assign n32264 = ~n31409 & ~n32263;
  assign n32265 = ~n32254 & n32264;
  assign n32266 = ~pi54 & ~n32265;
  assign n32267 = ~n31430 & ~n32266;
  assign n32268 = ~pi74 & ~n32267;
  assign n32269 = n31418 & ~n32268;
  assign n32270 = n62380 & n2814;
  assign n32271 = ~pi39 & pi232;
  assign n32272 = ~pi92 & pi162;
  assign n32273 = n9735 & n32272;
  assign n32274 = n32271 & n32272;
  assign n32275 = n9735 & n32274;
  assign n32276 = n32271 & n32273;
  assign n32277 = n32270 & n64194;
  assign n32278 = ~n31377 & ~n32277;
  assign n32279 = n2765 & ~n32278;
  assign n32280 = n31376 & ~n32279;
  assign n32281 = ~n32041 & ~n32280;
  assign n32282 = ~pi74 & ~n32281;
  assign n32283 = n32040 & ~n32282;
  assign n32284 = n3470 & ~n32283;
  assign n32285 = ~n32269 & n32284;
  assign n32286 = n31384 & ~n32285;
  assign n32287 = ~n31375 & ~n32286;
  assign n32288 = pi34 & n32287;
  assign n32289 = ~pi33 & ~pi954;
  assign n32290 = ~n32288 & ~n32289;
  assign n32291 = ~n32073 & n32290;
  assign n32292 = ~pi195 & ~pi196;
  assign n32293 = ~pi138 & n32292;
  assign n32294 = ~pi139 & n32293;
  assign n32295 = ~pi118 & n32294;
  assign n32296 = ~pi79 & n32295;
  assign n32297 = ~pi34 & ~n32296;
  assign n32298 = n32072 & ~n32297;
  assign n32299 = n32287 & n32297;
  assign n32300 = n32289 & ~n32299;
  assign n32301 = ~n32298 & n32300;
  assign po192 = ~n32291 & ~n32301;
  assign n32303 = pi163 & ~n31358;
  assign n32304 = ~pi163 & ~n31353;
  assign n32305 = ~n31356 & n32304;
  assign n32306 = ~n32303 & ~n32305;
  assign n32307 = pi232 & n32306;
  assign n32308 = pi75 & ~n32307;
  assign n32309 = pi100 & ~n32307;
  assign n32310 = ~n32308 & ~n32309;
  assign n32311 = pi147 & n2815;
  assign n32312 = n2765 & n32311;
  assign n32313 = n32310 & ~n32312;
  assign n32314 = ~n2765 & n32307;
  assign n32315 = pi74 & ~n32314;
  assign n32316 = ~n3472 & ~n32315;
  assign n32317 = n32313 & n32316;
  assign n32318 = pi299 & ~n32306;
  assign n32319 = ~n31395 & n31397;
  assign n32320 = pi184 & n2814;
  assign n32321 = ~n32319 & n32320;
  assign n32322 = ~pi184 & n32319;
  assign n32323 = ~pi299 & ~n32322;
  assign n32324 = ~n32319 & ~n32320;
  assign n32325 = pi184 & n32319;
  assign n32326 = ~n32324 & ~n32325;
  assign n32327 = ~pi299 & ~n32326;
  assign n32328 = ~pi299 & ~n32321;
  assign n32329 = ~n32322 & n32328;
  assign n32330 = ~n32321 & n32323;
  assign n32331 = pi232 & ~n64195;
  assign n32332 = ~n32318 & n32331;
  assign n32333 = ~n2765 & n32332;
  assign n32334 = pi74 & ~n32333;
  assign n32335 = ~pi55 & ~n32334;
  assign n32336 = ~pi187 & ~pi299;
  assign n32337 = ~pi147 & pi299;
  assign n32338 = ~n32336 & ~n32337;
  assign n32339 = n2815 & n32338;
  assign n32340 = n2765 & ~n32339;
  assign n32341 = pi54 & ~n32340;
  assign n32342 = ~n32333 & n32341;
  assign n32343 = ~pi187 & ~n64172;
  assign n32344 = pi187 & ~n31980;
  assign n32345 = pi147 & ~n32344;
  assign n32346 = ~n32343 & n32345;
  assign n32347 = ~pi147 & pi187;
  assign n32348 = n31978 & n32347;
  assign n32349 = ~n32346 & ~n32348;
  assign n32350 = pi38 & ~n32349;
  assign n32351 = ~pi40 & ~n31625;
  assign n32352 = ~pi95 & ~n32351;
  assign n32353 = ~pi40 & ~n31586;
  assign n32354 = pi166 & n32353;
  assign n32355 = n32352 & ~n32354;
  assign n32356 = n2814 & ~n31547;
  assign n32357 = ~n32355 & n32356;
  assign n32358 = ~pi153 & ~n32357;
  assign n32359 = ~pi40 & ~n31565;
  assign n32360 = ~pi95 & ~n32359;
  assign n32361 = pi166 & ~n32360;
  assign n32362 = n32356 & n32361;
  assign n32363 = ~pi166 & n2814;
  assign n32364 = n31528 & n32363;
  assign n32365 = pi153 & ~n32364;
  assign n32366 = ~n32362 & n32365;
  assign n32367 = pi160 & ~n32366;
  assign n32368 = ~n32358 & n32367;
  assign n32369 = ~pi153 & n32355;
  assign n32370 = ~n30613 & ~n31547;
  assign n32371 = n31433 & ~n31441;
  assign n32372 = ~n32370 & ~n32371;
  assign n32373 = n2751 & n62768;
  assign n32374 = n2694 & n2751;
  assign n32375 = n62382 & n32374;
  assign n32376 = n2728 & n64089;
  assign n32377 = n2751 & n32119;
  assign n32378 = n32114 & n64196;
  assign n32379 = ~n32360 & ~n64197;
  assign n32380 = pi153 & ~n32361;
  assign n32381 = ~n32379 & n32380;
  assign n32382 = ~pi160 & n2814;
  assign n32383 = ~n32381 & n32382;
  assign n32384 = ~n32372 & n32383;
  assign n32385 = ~n32369 & n32384;
  assign n32386 = pi163 & ~n32385;
  assign n32387 = ~n32368 & n32386;
  assign n32388 = ~pi40 & ~n31825;
  assign n32389 = ~pi95 & ~n32388;
  assign n32390 = ~n32372 & ~n32389;
  assign n32391 = pi166 & n32390;
  assign n32392 = ~pi40 & n31671;
  assign n32393 = ~pi32 & ~n32392;
  assign n32394 = ~n31529 & ~n32393;
  assign n32395 = ~pi95 & ~n32394;
  assign n32396 = ~n32372 & ~n32395;
  assign n32397 = pi210 & ~n32396;
  assign n32398 = ~n31549 & ~n32393;
  assign n32399 = ~pi95 & ~n32398;
  assign n32400 = ~n32372 & ~n32399;
  assign n32401 = ~pi210 & ~n32400;
  assign n32402 = n32363 & ~n32401;
  assign n32403 = n32363 & ~n32397;
  assign n32404 = ~n32401 & n32403;
  assign n32405 = ~n32397 & n32402;
  assign n32406 = ~pi153 & ~n64198;
  assign n32407 = ~n32391 & n32406;
  assign n32408 = ~pi210 & n31551;
  assign n32409 = pi166 & n2814;
  assign n32410 = ~pi95 & ~n31540;
  assign n32411 = pi210 & n32410;
  assign n32412 = n32409 & ~n32411;
  assign n32413 = ~n32408 & n32409;
  assign n32414 = ~n32411 & n32413;
  assign n32415 = ~n32408 & n32412;
  assign n32416 = pi210 & n31649;
  assign n32417 = ~pi210 & n31652;
  assign n32418 = n32363 & ~n32417;
  assign n32419 = ~n32416 & n32418;
  assign n32420 = ~n64199 & ~n32419;
  assign n32421 = ~n32372 & ~n32420;
  assign n32422 = ~n31652 & ~n32372;
  assign n32423 = ~pi210 & ~n32422;
  assign n32424 = ~n31649 & ~n32372;
  assign n32425 = pi210 & ~n32424;
  assign n32426 = n32363 & ~n32425;
  assign n32427 = n32363 & ~n32423;
  assign n32428 = ~n32425 & n32427;
  assign n32429 = ~n32423 & n32426;
  assign n32430 = ~n32372 & ~n32410;
  assign n32431 = pi210 & ~n32430;
  assign n32432 = ~n31551 & ~n32372;
  assign n32433 = ~pi210 & ~n32432;
  assign n32434 = n32409 & ~n32433;
  assign n32435 = n32409 & ~n32431;
  assign n32436 = ~n32433 & n32435;
  assign n32437 = ~n32431 & n32434;
  assign n32438 = pi153 & ~n64201;
  assign n32439 = ~n64200 & n32438;
  assign n32440 = pi153 & ~n64200;
  assign n32441 = ~n64201 & n32440;
  assign n32442 = pi153 & ~n32421;
  assign n32443 = ~pi160 & ~n64202;
  assign n32444 = ~n32407 & n32443;
  assign n32445 = n32388 & n32409;
  assign n32446 = ~n31547 & ~n32399;
  assign n32447 = ~pi210 & ~n32446;
  assign n32448 = ~n31547 & ~n32395;
  assign n32449 = pi210 & ~n32448;
  assign n32450 = n32363 & ~n32449;
  assign n32451 = n32363 & ~n32447;
  assign n32452 = ~n32449 & n32451;
  assign n32453 = ~n32447 & n32450;
  assign n32454 = ~pi153 & ~n64203;
  assign n32455 = ~n32445 & n32454;
  assign n32456 = ~n31547 & ~n32420;
  assign n32457 = ~pi210 & ~n31552;
  assign n32458 = ~n31547 & ~n32410;
  assign n32459 = pi210 & ~n32458;
  assign n32460 = n32409 & ~n32459;
  assign n32461 = n32409 & ~n32457;
  assign n32462 = ~n32459 & n32461;
  assign n32463 = ~n32457 & n32460;
  assign n32464 = pi210 & ~n31655;
  assign n32465 = ~pi210 & ~n31657;
  assign n32466 = n32363 & ~n32465;
  assign n32467 = n32363 & ~n32464;
  assign n32468 = ~n32465 & n32467;
  assign n32469 = ~n32464 & n32466;
  assign n32470 = pi153 & ~n64205;
  assign n32471 = ~n64204 & n32470;
  assign n32472 = pi153 & ~n64204;
  assign n32473 = ~n64205 & n32472;
  assign n32474 = pi153 & ~n32456;
  assign n32475 = pi160 & ~n64206;
  assign n32476 = ~n32455 & n32475;
  assign n32477 = ~pi163 & ~n32476;
  assign n32478 = ~n32444 & n32477;
  assign n32479 = ~n32387 & ~n32478;
  assign n32480 = ~n2814 & n32390;
  assign n32481 = pi299 & ~n32480;
  assign n32482 = ~n32479 & n32481;
  assign n32483 = ~pi40 & ~n31612;
  assign n32484 = ~pi95 & ~n32483;
  assign n32485 = ~n32372 & ~n32484;
  assign n32486 = ~n2814 & n32485;
  assign n32487 = ~pi175 & ~pi299;
  assign n32488 = pi189 & n32353;
  assign n32489 = n32352 & ~n32488;
  assign n32490 = ~pi182 & n32372;
  assign n32491 = pi182 & n31547;
  assign n32492 = n2814 & ~n32491;
  assign n32493 = n2814 & ~n32490;
  assign n32494 = ~n32491 & n32493;
  assign n32495 = ~n32490 & n32492;
  assign n32496 = ~n32489 & n64207;
  assign n32497 = pi184 & ~n32496;
  assign n32498 = pi189 & n2814;
  assign n32499 = n32483 & n32498;
  assign n32500 = pi198 & ~n32448;
  assign n32501 = ~pi189 & n2814;
  assign n32502 = ~pi198 & ~n32446;
  assign n32503 = n32501 & ~n32502;
  assign n32504 = ~n32500 & n32501;
  assign n32505 = ~n32502 & n32504;
  assign n32506 = ~n32500 & n32503;
  assign n32507 = pi182 & ~pi184;
  assign n32508 = ~n64208 & n32507;
  assign n32509 = ~n32499 & n32508;
  assign n32510 = ~n32497 & ~n32509;
  assign n32511 = n32487 & ~n32510;
  assign n32512 = ~pi198 & ~n31551;
  assign n32513 = pi198 & ~n32410;
  assign n32514 = ~n32512 & ~n32513;
  assign n32515 = pi189 & n64207;
  assign n32516 = ~n32514 & n32515;
  assign n32517 = pi95 & ~pi182;
  assign n32518 = ~n64151 & ~n32517;
  assign n32519 = ~pi189 & n32493;
  assign n32520 = ~n32372 & n32501;
  assign n32521 = ~n32518 & n32520;
  assign n32522 = ~n32518 & n32519;
  assign n32523 = n64151 & n32501;
  assign n32524 = ~pi198 & ~n31552;
  assign n32525 = pi198 & ~n32458;
  assign n32526 = n32498 & ~n32525;
  assign n32527 = n32498 & ~n32524;
  assign n32528 = ~n32525 & n32527;
  assign n32529 = ~n32524 & n32526;
  assign n32530 = pi182 & ~n64210;
  assign n32531 = pi182 & ~n32523;
  assign n32532 = ~n64210 & n32531;
  assign n32533 = ~n32523 & n32530;
  assign n32534 = ~pi198 & ~n32432;
  assign n32535 = pi198 & ~n32430;
  assign n32536 = n32498 & ~n32535;
  assign n32537 = n32498 & ~n32534;
  assign n32538 = ~n32535 & n32537;
  assign n32539 = ~n32534 & n32536;
  assign n32540 = ~pi182 & ~n64212;
  assign n32541 = ~n64211 & ~n32540;
  assign n32542 = ~n64209 & ~n32541;
  assign n32543 = ~n32516 & ~n64209;
  assign n32544 = ~pi184 & ~n64213;
  assign n32545 = pi175 & ~pi299;
  assign n32546 = ~pi95 & pi189;
  assign n32547 = n2587 & ~n32546;
  assign n32548 = n32359 & ~n32547;
  assign n32549 = ~n32517 & ~n32548;
  assign n32550 = n32320 & ~n32549;
  assign n32551 = ~n32490 & n32550;
  assign n32552 = n32545 & ~n32551;
  assign n32553 = ~n32544 & n32552;
  assign n32554 = ~n32511 & ~n32553;
  assign n32555 = ~n32486 & ~n32554;
  assign n32556 = n32485 & ~n32501;
  assign n32557 = ~pi198 & ~n32400;
  assign n32558 = pi198 & ~n32396;
  assign n32559 = n32501 & ~n32558;
  assign n32560 = n32501 & ~n32557;
  assign n32561 = ~n32558 & n32560;
  assign n32562 = ~n32557 & n32559;
  assign n32563 = ~pi182 & ~pi184;
  assign n32564 = n32487 & n32563;
  assign n32565 = ~n64214 & n32564;
  assign n32566 = ~n32556 & n32565;
  assign n32567 = ~n32555 & ~n32566;
  assign n32568 = ~n32482 & n32567;
  assign n32569 = pi232 & ~n32568;
  assign n32570 = pi299 & n32390;
  assign n32571 = ~pi299 & n32485;
  assign n32572 = ~pi232 & ~n32571;
  assign n32573 = ~pi232 & ~n32570;
  assign n32574 = ~n32571 & n32573;
  assign n32575 = ~n32570 & n32572;
  assign n32576 = ~pi39 & ~n64215;
  assign n32577 = ~n32569 & n32576;
  assign n32578 = ~n31528 & ~n31926;
  assign n32579 = ~pi40 & ~n31895;
  assign n32580 = ~pi189 & ~n32579;
  assign n32581 = n2587 & ~n31912;
  assign n32582 = n31610 & ~n32581;
  assign n32583 = n2953 & n31528;
  assign n32584 = n2587 & ~n31893;
  assign n32585 = ~pi40 & ~n32584;
  assign n32586 = n2909 & n32585;
  assign n32587 = ~n32583 & ~n32586;
  assign n32588 = ~n32582 & n32587;
  assign n32589 = pi189 & ~n2971;
  assign n32590 = n32588 & n32589;
  assign n32591 = ~n32580 & ~n32590;
  assign n32592 = pi179 & ~n32591;
  assign n32593 = n2971 & ~n32579;
  assign n32594 = n2587 & ~n31900;
  assign n32595 = n31610 & n31900;
  assign n32596 = ~n2587 & n31610;
  assign n32597 = ~n32595 & ~n32596;
  assign n32598 = n31610 & ~n32594;
  assign n32599 = n32587 & n64216;
  assign n32600 = ~pi189 & ~n32599;
  assign n32601 = ~n2953 & n32585;
  assign n32602 = ~n32583 & ~n32601;
  assign n32603 = pi189 & ~n32602;
  assign n32604 = ~pi179 & ~n2971;
  assign n32605 = ~n32603 & n32604;
  assign n32606 = ~n32600 & n32605;
  assign n32607 = ~n32593 & ~n32606;
  assign n32608 = ~n32592 & n32607;
  assign n32609 = n31926 & ~n32608;
  assign n32610 = ~n32578 & ~n32609;
  assign n32611 = ~pi299 & ~n32610;
  assign n32612 = n31528 & ~n31886;
  assign n32613 = pi299 & ~n32612;
  assign n32614 = pi166 & ~n62393;
  assign n32615 = n32588 & n32614;
  assign n32616 = ~n32579 & ~n32614;
  assign n32617 = n31886 & ~n32616;
  assign n32618 = ~n32615 & n32617;
  assign n32619 = n32613 & ~n32618;
  assign n32620 = ~n32611 & ~n32619;
  assign n32621 = pi156 & pi232;
  assign n32622 = ~n32620 & n32621;
  assign n32623 = ~n62393 & n32602;
  assign n32624 = n62393 & ~n32579;
  assign n32625 = ~n62393 & ~n32602;
  assign n32626 = n62393 & n32579;
  assign n32627 = ~n32625 & ~n32626;
  assign n32628 = ~n32623 & ~n32624;
  assign n32629 = ~pi166 & ~n62393;
  assign n32630 = n64217 & ~n32629;
  assign n32631 = n32599 & n32629;
  assign n32632 = n31886 & ~n32631;
  assign n32633 = ~n32630 & n32632;
  assign n32634 = n32613 & ~n32633;
  assign n32635 = ~n32611 & ~n32634;
  assign n32636 = ~pi156 & pi232;
  assign n32637 = ~n32635 & n32636;
  assign n32638 = ~n2971 & n32602;
  assign n32639 = ~n32593 & ~n32638;
  assign n32640 = n31926 & ~n32639;
  assign n32641 = ~pi299 & ~n32578;
  assign n32642 = ~n32640 & n32641;
  assign n32643 = n31908 & ~n64217;
  assign n32644 = ~pi232 & ~n32643;
  assign n32645 = ~n32642 & n32644;
  assign n32646 = pi39 & ~n32645;
  assign n32647 = ~n32637 & n32646;
  assign n32648 = ~n32622 & n32646;
  assign n32649 = ~n32637 & n32648;
  assign n32650 = ~n32622 & n32647;
  assign n32651 = ~pi38 & ~n64218;
  assign n32652 = ~n32577 & n32651;
  assign n32653 = ~n32350 & ~n32652;
  assign n32654 = n6791 & ~n32653;
  assign n32655 = pi100 & ~n32332;
  assign n32656 = pi38 & ~n32339;
  assign n32657 = ~pi100 & ~n32656;
  assign n32658 = ~pi38 & ~pi40;
  assign n32659 = pi87 & ~n2587;
  assign n32660 = n32658 & n32659;
  assign n32661 = n32657 & ~n32660;
  assign n32662 = pi87 & n32661;
  assign n32663 = ~n32655 & ~n32662;
  assign n32664 = ~n32654 & n32663;
  assign n32665 = n6793 & ~n32664;
  assign n32666 = pi75 & ~n32332;
  assign n32667 = pi39 & ~n31528;
  assign n32668 = n9735 & ~n32667;
  assign n32669 = n2587 & ~n31887;
  assign n32670 = ~pi40 & ~n32669;
  assign n32671 = ~pi179 & ~pi299;
  assign n32672 = ~pi156 & pi299;
  assign n32673 = ~n32671 & ~n32672;
  assign n32674 = n2815 & n32673;
  assign n32675 = n2587 & n32674;
  assign n32676 = n32670 & ~n32675;
  assign n32677 = ~pi39 & ~n32676;
  assign n32678 = n32668 & ~n32677;
  assign n32679 = n32661 & ~n32678;
  assign n32680 = ~n32655 & ~n32679;
  assign n32681 = n32018 & ~n32680;
  assign n32682 = ~n32666 & ~n32681;
  assign n32683 = ~n32665 & n32682;
  assign n32684 = ~pi54 & ~n32683;
  assign n32685 = ~n32342 & ~n32684;
  assign n32686 = ~pi74 & ~n32685;
  assign n32687 = n32335 & ~n32686;
  assign n32688 = pi55 & ~n32315;
  assign n32689 = pi54 & ~n32313;
  assign n32690 = pi163 & pi232;
  assign n32691 = ~n2814 & n31887;
  assign n32692 = n31385 & ~n32691;
  assign n32693 = n32690 & n32692;
  assign n32694 = n32670 & ~n32693;
  assign n32695 = ~pi39 & ~n32694;
  assign n32696 = n32668 & ~n32695;
  assign n32697 = pi38 & ~n32311;
  assign n32698 = ~pi100 & ~n32697;
  assign n32699 = ~n32660 & n32698;
  assign n32700 = ~n32696 & n32699;
  assign n32701 = ~n32309 & ~n32700;
  assign n32702 = n6793 & ~n32701;
  assign n32703 = n2766 & n31385;
  assign n32704 = ~n32658 & n32698;
  assign n32705 = ~n32309 & ~n32704;
  assign n32706 = ~n32703 & n32705;
  assign n32707 = n32018 & ~n32706;
  assign n32708 = ~n32308 & ~n32707;
  assign n32709 = ~n32702 & n32708;
  assign n32710 = ~pi54 & ~n32709;
  assign n32711 = ~n32689 & ~n32710;
  assign n32712 = ~pi74 & ~n32711;
  assign n32713 = n32688 & ~n32712;
  assign n32714 = n3470 & ~n32713;
  assign n32715 = ~n32687 & n32714;
  assign n32716 = ~n3470 & n31388;
  assign n32717 = ~pi75 & ~n32705;
  assign n32718 = ~n32308 & ~n32717;
  assign n32719 = ~pi54 & ~n32718;
  assign n32720 = ~n32689 & ~n32719;
  assign n32721 = ~pi74 & ~n32720;
  assign n32722 = ~n32315 & ~n32721;
  assign n32723 = ~n3470 & ~n32722;
  assign n32724 = n3472 & ~n32723;
  assign n32725 = ~n32716 & n32724;
  assign n32726 = ~n32715 & n32725;
  assign n32727 = ~n32317 & ~n32726;
  assign n32728 = ~pi79 & n32727;
  assign n32729 = pi153 & pi160;
  assign n32730 = ~n32095 & ~n32729;
  assign n32731 = ~pi32 & pi95;
  assign n32732 = ~pi479 & n32731;
  assign n32733 = n62383 & n32732;
  assign n32734 = n2814 & n32733;
  assign n32735 = ~n30611 & ~n32094;
  assign n32736 = ~pi210 & ~n32735;
  assign n32737 = ~n32734 & ~n32736;
  assign n32738 = pi160 & ~n32737;
  assign n32739 = ~n32092 & ~n32738;
  assign n32740 = pi160 & n32734;
  assign n32741 = ~pi153 & ~n32740;
  assign n32742 = ~n32739 & ~n32741;
  assign n32743 = ~n32730 & ~n32742;
  assign n32744 = ~n32363 & ~n32740;
  assign n32745 = pi153 & n32092;
  assign n32746 = n32095 & ~n32745;
  assign n32747 = n32363 & ~n32746;
  assign n32748 = ~pi160 & ~n32747;
  assign n32749 = ~n32092 & ~n32736;
  assign n32750 = pi153 & ~n32749;
  assign n32751 = ~pi153 & ~n32095;
  assign n32752 = pi160 & ~n32751;
  assign n32753 = ~n32750 & n32752;
  assign n32754 = n32363 & ~n32753;
  assign n32755 = ~n32734 & ~n32754;
  assign n32756 = ~n32748 & ~n32755;
  assign n32757 = ~n32743 & ~n32744;
  assign n32758 = pi153 & n32101;
  assign n32759 = n32104 & ~n32758;
  assign n32760 = n32409 & ~n32759;
  assign n32761 = ~pi40 & pi163;
  assign n32762 = ~n32760 & n32761;
  assign n32763 = ~n64219 & n32762;
  assign n32764 = pi153 & n32111;
  assign n32765 = n64180 & n32764;
  assign n32766 = n32120 & n32363;
  assign n32767 = ~pi40 & ~pi163;
  assign n32768 = ~n32766 & n32767;
  assign n32769 = ~n32740 & n32768;
  assign n32770 = ~n32765 & n32768;
  assign n32771 = ~n32740 & n32770;
  assign n32772 = ~n32765 & n32769;
  assign n32773 = pi299 & ~n64220;
  assign n32774 = ~pi40 & ~n32733;
  assign n32775 = n32095 & n32774;
  assign n32776 = n32363 & ~n32775;
  assign n32777 = n32104 & n32774;
  assign n32778 = n32409 & ~n32777;
  assign n32779 = ~pi153 & ~n32778;
  assign n32780 = ~n32776 & n32779;
  assign n32781 = ~n32092 & n32774;
  assign n32782 = ~n32736 & n32781;
  assign n32783 = n32363 & ~n32782;
  assign n32784 = ~n32101 & n32777;
  assign n32785 = n32409 & ~n32784;
  assign n32786 = pi153 & ~n32785;
  assign n32787 = ~n32783 & n32786;
  assign n32788 = ~n32780 & ~n32787;
  assign n32789 = pi40 & ~n2814;
  assign n32790 = pi163 & ~n32789;
  assign n32791 = ~n32788 & n32790;
  assign n32792 = pi160 & ~n32791;
  assign n32793 = ~n32747 & n32762;
  assign n32794 = ~pi160 & ~n32770;
  assign n32795 = ~n32793 & n32794;
  assign n32796 = ~n32792 & ~n32795;
  assign n32797 = ~n32734 & n32770;
  assign n32798 = pi299 & ~n32797;
  assign n32799 = ~n32796 & n32798;
  assign n32800 = ~n32763 & n32773;
  assign n32801 = pi184 & n32152;
  assign n32802 = ~pi184 & ~n32120;
  assign n32803 = ~pi189 & ~n32802;
  assign n32804 = ~n32801 & n32803;
  assign n32805 = pi182 & n32733;
  assign n32806 = pi184 & pi189;
  assign n32807 = ~n32156 & n32806;
  assign n32808 = ~n32805 & ~n32807;
  assign n32809 = ~n32804 & n32808;
  assign n32810 = n2814 & ~n32809;
  assign n32811 = ~pi40 & ~n32810;
  assign n32812 = n32487 & ~n32811;
  assign n32813 = ~pi189 & ~n32116;
  assign n32814 = pi189 & ~n64180;
  assign n32815 = n2727 & ~n32814;
  assign n32816 = n2727 & ~n32813;
  assign n32817 = ~n32814 & n32816;
  assign n32818 = ~n32813 & n32815;
  assign n32819 = ~n32805 & ~n64222;
  assign n32820 = n2814 & ~n32819;
  assign n32821 = ~pi184 & ~n32820;
  assign n32822 = ~pi198 & ~n32735;
  assign n32823 = ~n32092 & ~n32822;
  assign n32824 = n32501 & ~n32823;
  assign n32825 = ~pi182 & pi184;
  assign n32826 = ~n30612 & ~n32101;
  assign n32827 = n2814 & ~n32826;
  assign n32828 = pi189 & n32827;
  assign n32829 = n32825 & ~n32828;
  assign n32830 = ~n32824 & n32829;
  assign n32831 = ~n32821 & ~n32830;
  assign n32832 = ~pi40 & ~n32831;
  assign n32833 = n32781 & ~n32822;
  assign n32834 = n32501 & ~n32833;
  assign n32835 = n32774 & n32826;
  assign n32836 = n32498 & ~n32835;
  assign n32837 = pi182 & pi184;
  assign n32838 = ~n32789 & n32837;
  assign n32839 = ~n32836 & n32838;
  assign n32840 = ~n32834 & n32839;
  assign n32841 = n32545 & ~n32840;
  assign n32842 = ~pi189 & ~n32823;
  assign n32843 = pi189 & ~n32826;
  assign n32844 = ~n32842 & ~n32843;
  assign n32845 = pi184 & ~n32733;
  assign n32846 = n32844 & n32845;
  assign n32847 = ~pi184 & ~n32805;
  assign n32848 = ~n64222 & n32847;
  assign n32849 = n2814 & ~n32825;
  assign n32850 = ~n32848 & n32849;
  assign n32851 = ~n32846 & n32850;
  assign n32852 = n2814 & n32825;
  assign n32853 = ~n32844 & n32852;
  assign n32854 = ~pi40 & ~n32853;
  assign n32855 = ~n32851 & n32854;
  assign n32856 = n32545 & ~n32855;
  assign n32857 = ~n32832 & n32841;
  assign n32858 = ~n32812 & ~n64223;
  assign n32859 = ~n64221 & n32858;
  assign n32860 = ~pi39 & ~n32859;
  assign n32861 = n62383 & n32111;
  assign n32862 = ~pi189 & n31891;
  assign n32863 = pi179 & n31888;
  assign n32864 = ~n32862 & ~n32863;
  assign n32865 = n32221 & ~n32864;
  assign n32866 = n32861 & n32865;
  assign n32867 = ~pi40 & ~pi299;
  assign n32868 = ~n32866 & n32867;
  assign n32869 = pi156 & n31888;
  assign n32870 = ~pi166 & n31891;
  assign n32871 = ~n32869 & ~n32870;
  assign n32872 = ~n62393 & n31886;
  assign n32873 = ~n32871 & n32872;
  assign n32874 = n32861 & n32873;
  assign n32875 = ~pi40 & pi299;
  assign n32876 = ~n32874 & n32875;
  assign n32877 = pi39 & ~n32876;
  assign n32878 = pi39 & ~n32868;
  assign n32879 = ~n32876 & n32878;
  assign n32880 = ~n32868 & n32877;
  assign n32881 = pi232 & ~n64224;
  assign n32882 = ~n32860 & n32881;
  assign n32883 = ~pi40 & ~pi232;
  assign n32884 = ~pi38 & ~n32883;
  assign n32885 = ~n32882 & n32884;
  assign n32886 = ~n32350 & ~n32885;
  assign n32887 = n6791 & ~n32886;
  assign n32888 = pi87 & ~n32658;
  assign n32889 = n32657 & n32888;
  assign n32890 = ~n32655 & ~n32889;
  assign n32891 = ~n32887 & n32890;
  assign n32892 = n6793 & ~n32891;
  assign n32893 = n2727 & n2805;
  assign n32894 = n32674 & n32893;
  assign n32895 = n62383 & n32894;
  assign n32896 = n32658 & ~n32895;
  assign n32897 = n32657 & ~n32896;
  assign n32898 = ~n32655 & ~n32897;
  assign n32899 = n32018 & ~n32898;
  assign n32900 = ~n32666 & ~n32899;
  assign n32901 = ~n32892 & n32900;
  assign n32902 = ~pi54 & ~n32901;
  assign n32903 = ~n32342 & ~n32902;
  assign n32904 = ~pi74 & ~n32903;
  assign n32905 = n32335 & ~n32904;
  assign n32906 = ~pi92 & n2805;
  assign n32907 = n32690 & n32906;
  assign n32908 = n32861 & n32907;
  assign n32909 = n32658 & ~n32908;
  assign n32910 = ~pi75 & n32698;
  assign n32911 = ~n32909 & n32910;
  assign n32912 = n32310 & ~n32911;
  assign n32913 = ~pi54 & ~n32912;
  assign n32914 = ~n32689 & ~n32913;
  assign n32915 = ~pi74 & ~n32914;
  assign n32916 = n32688 & ~n32915;
  assign n32917 = n3470 & ~n32916;
  assign n32918 = ~n32905 & n32917;
  assign n32919 = n32724 & ~n32918;
  assign n32920 = ~n32317 & ~n32919;
  assign n32921 = pi79 & n32920;
  assign n32922 = ~pi34 & n32289;
  assign n32923 = ~n32921 & ~n32922;
  assign n32924 = ~n32728 & n32923;
  assign n32925 = ~pi79 & ~n32295;
  assign n32926 = n32727 & ~n32925;
  assign n32927 = n32920 & n32925;
  assign n32928 = n32922 & ~n32927;
  assign n32929 = ~n32926 & n32928;
  assign n32930 = ~n32924 & ~n32929;
  assign n32931 = pi163 & n2814;
  assign n32932 = ~n32306 & ~n32931;
  assign n32933 = ~pi150 & ~n32932;
  assign n32934 = pi150 & n31357;
  assign n32935 = n32304 & n32934;
  assign n32936 = ~n32933 & ~n32935;
  assign n32937 = pi232 & ~n32936;
  assign n32938 = ~n2765 & n32937;
  assign n32939 = n31361 & ~n32936;
  assign n32940 = pi165 & n2815;
  assign n32941 = ~pi74 & n2765;
  assign n32942 = ~n32940 & n32941;
  assign n32943 = ~n64225 & ~n32942;
  assign n32944 = pi74 & ~n64225;
  assign n32945 = ~n2765 & ~n32937;
  assign n32946 = n2765 & n32940;
  assign n32947 = ~n3472 & ~n32946;
  assign n32948 = n2765 & ~n32940;
  assign n32949 = ~n64225 & ~n32948;
  assign n32950 = ~n3472 & ~n32949;
  assign n32951 = ~n32945 & n32947;
  assign n32952 = ~n32944 & n64226;
  assign n32953 = ~n3472 & ~n32943;
  assign n32954 = ~pi74 & ~n64225;
  assign n32955 = ~pi38 & ~pi54;
  assign n32956 = ~n32940 & ~n32955;
  assign n32957 = n2765 & n32956;
  assign n32958 = n32954 & ~n32957;
  assign n32959 = ~n32944 & ~n32958;
  assign n32960 = ~n3470 & ~n32959;
  assign n32961 = n3472 & ~n32960;
  assign n32962 = ~n31390 & ~n32961;
  assign n32963 = pi299 & n32936;
  assign n32964 = ~pi184 & ~n32319;
  assign n32965 = pi185 & ~n32964;
  assign n32966 = ~pi185 & n32964;
  assign n32967 = n2814 & ~n32966;
  assign n32968 = n2814 & ~n32965;
  assign n32969 = ~n32966 & n32968;
  assign n32970 = ~n32965 & n32967;
  assign n32971 = ~pi299 & ~n64228;
  assign n32972 = pi232 & ~n32971;
  assign n32973 = ~n32963 & n32972;
  assign n32974 = ~n2765 & n32973;
  assign n32975 = pi74 & ~n32974;
  assign n32976 = ~pi55 & ~n32975;
  assign n32977 = ~pi143 & ~pi299;
  assign n32978 = ~pi165 & pi299;
  assign n32979 = ~n32977 & ~n32978;
  assign n32980 = n2815 & n32979;
  assign n32981 = n2765 & ~n32980;
  assign n32982 = pi54 & ~n32981;
  assign n32983 = ~n32974 & n32982;
  assign n32984 = ~pi143 & ~n64172;
  assign n32985 = pi143 & ~n31980;
  assign n32986 = pi165 & ~n32985;
  assign n32987 = ~n32984 & n32986;
  assign n32988 = pi143 & ~pi165;
  assign n32989 = n31978 & n32988;
  assign n32990 = pi38 & ~n32989;
  assign n32991 = ~n32987 & n32990;
  assign n32992 = n6791 & ~n32991;
  assign n32993 = ~n2814 & n31709;
  assign n32994 = pi151 & ~pi168;
  assign n32995 = ~n31843 & n32994;
  assign n32996 = pi168 & n31834;
  assign n32997 = ~pi168 & n31837;
  assign n32998 = ~pi151 & ~n32997;
  assign n32999 = ~n32996 & n32998;
  assign n33000 = ~n32995 & ~n32999;
  assign n33001 = ~n32993 & ~n33000;
  assign n33002 = ~n2814 & ~n31709;
  assign n33003 = n2814 & ~n31763;
  assign n33004 = ~n33002 & ~n33003;
  assign n33005 = pi151 & pi168;
  assign n33006 = ~n33004 & n33005;
  assign n33007 = pi150 & ~n33006;
  assign n33008 = ~n33001 & n33007;
  assign n33009 = ~n31589 & ~n33002;
  assign n33010 = pi168 & n33009;
  assign n33011 = ~n31714 & ~n33002;
  assign n33012 = ~pi168 & n33011;
  assign n33013 = pi151 & ~n33012;
  assign n33014 = ~n33010 & n33013;
  assign n33015 = pi168 & n31568;
  assign n33016 = pi168 & n2814;
  assign n33017 = n31709 & ~n33016;
  assign n33018 = ~pi151 & ~n33017;
  assign n33019 = ~pi151 & ~n33015;
  assign n33020 = ~n33017 & n33019;
  assign n33021 = ~n33015 & n33018;
  assign n33022 = ~pi150 & ~n64229;
  assign n33023 = ~n33014 & n33022;
  assign n33024 = pi299 & ~n33023;
  assign n33025 = ~n33008 & n33024;
  assign n33026 = ~n31557 & ~n32993;
  assign n33027 = ~pi173 & ~n33026;
  assign n33028 = n2814 & ~n31526;
  assign n33029 = pi173 & ~n33002;
  assign n33030 = ~n33028 & n33029;
  assign n33031 = pi185 & ~n33030;
  assign n33032 = ~n33027 & n33031;
  assign n33033 = pi173 & n33009;
  assign n33034 = ~n31568 & ~n32993;
  assign n33035 = ~pi173 & ~n33034;
  assign n33036 = ~pi185 & ~n33035;
  assign n33037 = pi173 & ~n33009;
  assign n33038 = ~pi173 & ~n31568;
  assign n33039 = ~n32993 & n33038;
  assign n33040 = ~n33037 & ~n33039;
  assign n33041 = ~pi185 & ~n33040;
  assign n33042 = ~n33033 & n33036;
  assign n33043 = pi190 & ~n64230;
  assign n33044 = ~n33032 & n33043;
  assign n33045 = pi173 & ~n31702;
  assign n33046 = ~pi173 & ~n31697;
  assign n33047 = n2814 & ~n33046;
  assign n33048 = ~pi173 & n31697;
  assign n33049 = pi173 & n31702;
  assign n33050 = ~n33048 & ~n33049;
  assign n33051 = n2814 & ~n33050;
  assign n33052 = ~n33045 & n33047;
  assign n33053 = pi185 & ~n32993;
  assign n33054 = ~n64231 & n33053;
  assign n33055 = pi173 & n33011;
  assign n33056 = ~pi173 & n31709;
  assign n33057 = ~pi185 & ~n33056;
  assign n33058 = ~n33055 & n33057;
  assign n33059 = ~pi190 & ~n33058;
  assign n33060 = ~n33054 & n33059;
  assign n33061 = ~pi299 & ~n33060;
  assign n33062 = ~n33044 & n33061;
  assign n33063 = pi232 & ~n33062;
  assign n33064 = ~n33025 & n33063;
  assign n33065 = ~pi232 & n31709;
  assign n33066 = ~pi39 & ~n33065;
  assign n33067 = ~n33064 & n33066;
  assign n33068 = pi178 & ~n31893;
  assign n33069 = ~pi178 & ~n31912;
  assign n33070 = pi190 & ~n33069;
  assign n33071 = ~n33068 & n33070;
  assign n33072 = pi178 & ~pi190;
  assign n33073 = n31900 & n33072;
  assign n33074 = ~n33071 & ~n33073;
  assign n33075 = pi222 & pi224;
  assign n33076 = pi224 & n62403;
  assign n33077 = n2979 & n33075;
  assign n33078 = ~pi299 & n64189;
  assign n33079 = n2972 & n64232;
  assign n33080 = ~n33074 & n64233;
  assign n33081 = pi168 & n31912;
  assign n33082 = pi157 & n31900;
  assign n33083 = ~n33081 & ~n33082;
  assign n33084 = pi216 & pi221;
  assign n33085 = pi299 & n31886;
  assign n33086 = n2959 & n33084;
  assign n33087 = n2919 & n64234;
  assign n33088 = ~n33083 & n33087;
  assign n33089 = pi232 & n31385;
  assign n33090 = ~n33088 & n33089;
  assign n33091 = ~pi178 & ~pi299;
  assign n33092 = n2919 & n31886;
  assign n33093 = n2814 & n32872;
  assign n33094 = ~n33083 & n64235;
  assign n33095 = pi299 & ~n33094;
  assign n33096 = ~n33091 & ~n33095;
  assign n33097 = n31385 & ~n33096;
  assign n33098 = pi178 & ~n31939;
  assign n33099 = ~pi190 & ~n33098;
  assign n33100 = ~pi299 & ~n33099;
  assign n33101 = ~n33097 & ~n33100;
  assign n33102 = n2971 & ~n31385;
  assign n33103 = n31926 & ~n33102;
  assign n33104 = ~pi178 & n33103;
  assign n33105 = ~n31949 & n33104;
  assign n33106 = pi178 & n33103;
  assign n33107 = ~n31929 & n33106;
  assign n33108 = ~pi299 & ~n31927;
  assign n33109 = pi190 & n33108;
  assign n33110 = ~n33107 & n33109;
  assign n33111 = ~n33105 & n33109;
  assign n33112 = ~n33107 & n33111;
  assign n33113 = ~n33105 & n33110;
  assign n33114 = pi232 & ~n64236;
  assign n33115 = ~n33101 & n33114;
  assign n33116 = ~n33080 & n33090;
  assign n33117 = ~pi232 & n31385;
  assign n33118 = pi39 & ~n33117;
  assign n33119 = ~n64237 & n33118;
  assign n33120 = ~pi38 & ~n33119;
  assign n33121 = ~n33067 & n33120;
  assign n33122 = n32992 & ~n33121;
  assign n33123 = pi100 & ~n32973;
  assign n33124 = pi38 & ~n32980;
  assign n33125 = ~pi100 & ~n33124;
  assign n33126 = pi87 & n33125;
  assign n33127 = n3011 & ~n33124;
  assign n33128 = ~n31386 & n64238;
  assign n33129 = ~n33123 & ~n33128;
  assign n33130 = ~n33122 & n33129;
  assign n33131 = n6793 & ~n33130;
  assign n33132 = pi75 & ~n32973;
  assign n33133 = ~pi157 & pi299;
  assign n33134 = ~n33091 & ~n33133;
  assign n33135 = n2815 & n33134;
  assign n33136 = n64176 & n33135;
  assign n33137 = n31386 & ~n33136;
  assign n33138 = n33125 & ~n33137;
  assign n33139 = ~n33123 & ~n33138;
  assign n33140 = n32018 & ~n33139;
  assign n33141 = ~n33132 & ~n33140;
  assign n33142 = ~n33131 & n33141;
  assign n33143 = ~pi54 & ~n33142;
  assign n33144 = ~n32983 & ~n33143;
  assign n33145 = ~pi74 & ~n33144;
  assign n33146 = n32976 & ~n33145;
  assign n33147 = pi55 & ~n32944;
  assign n33148 = n31385 & n32955;
  assign n33149 = ~pi92 & n64176;
  assign n33150 = pi150 & n2815;
  assign n33151 = n33149 & n33150;
  assign n33152 = n33148 & ~n33151;
  assign n33153 = ~n32956 & ~n33152;
  assign n33154 = n2765 & ~n33153;
  assign n33155 = n32954 & ~n33154;
  assign n33156 = n33147 & ~n33155;
  assign n33157 = n3470 & ~n33156;
  assign n33158 = ~n33146 & n33157;
  assign n33159 = ~n32962 & ~n33158;
  assign n33160 = ~n64227 & ~n33159;
  assign n33161 = pi118 & n33160;
  assign n33162 = ~pi79 & n32922;
  assign n33163 = n2909 & ~n30820;
  assign n33164 = ~pi178 & n30820;
  assign n33165 = pi178 & ~n30824;
  assign n33166 = ~pi190 & ~n33165;
  assign n33167 = ~n33164 & n33166;
  assign n33168 = ~pi178 & pi190;
  assign n33169 = n62397 & n33168;
  assign n33170 = ~n33167 & ~n33169;
  assign n33171 = n2972 & ~n33170;
  assign n33172 = ~pi178 & ~n2971;
  assign n33173 = n32206 & n33172;
  assign n33174 = ~n33163 & ~n33173;
  assign n33175 = pi190 & ~n33174;
  assign n33176 = pi178 & ~n32234;
  assign n33177 = ~n33163 & n33176;
  assign n33178 = ~n2973 & ~n30820;
  assign n33179 = ~pi178 & ~n33178;
  assign n33180 = ~pi190 & ~n33179;
  assign n33181 = ~pi190 & ~n33177;
  assign n33182 = ~n33179 & n33181;
  assign n33183 = ~n33177 & n33180;
  assign n33184 = ~n33175 & ~n64239;
  assign n33185 = ~n33163 & ~n33171;
  assign n33186 = n64232 & ~n64240;
  assign n33187 = ~pi168 & ~n32204;
  assign n33188 = pi168 & ~n64187;
  assign n33189 = ~pi157 & ~n33188;
  assign n33190 = ~n33187 & n33189;
  assign n33191 = pi157 & ~pi168;
  assign n33192 = n32215 & n33191;
  assign n33193 = ~n33163 & ~n33192;
  assign n33194 = ~pi157 & n64187;
  assign n33195 = pi168 & ~n33194;
  assign n33196 = pi157 & ~n32215;
  assign n33197 = ~pi157 & ~pi168;
  assign n33198 = ~n32204 & n33197;
  assign n33199 = ~n33196 & ~n33198;
  assign n33200 = ~n33195 & n33199;
  assign n33201 = ~n33163 & ~n33200;
  assign n33202 = ~n33190 & n33193;
  assign n33203 = n64234 & ~n64241;
  assign n33204 = pi232 & ~n33203;
  assign n33205 = pi232 & ~n33186;
  assign n33206 = ~n33203 & n33205;
  assign n33207 = ~n33186 & n33204;
  assign n33208 = n30831 & n31886;
  assign n33209 = pi216 & ~n2920;
  assign n33210 = n2961 & n33209;
  assign n33211 = ~n2920 & n64234;
  assign n33212 = pi224 & n30839;
  assign n33213 = ~n2973 & n33075;
  assign n33214 = n2979 & n64244;
  assign n33215 = pi224 & n64102;
  assign n33216 = ~n2973 & n64232;
  assign n33217 = ~n64243 & ~n64245;
  assign n33218 = ~n30820 & ~n33217;
  assign n33219 = n30841 & n32224;
  assign n33220 = ~n30820 & n64243;
  assign n33221 = ~pi232 & ~n33220;
  assign n33222 = ~n33219 & n33221;
  assign n33223 = ~pi232 & ~n33218;
  assign n33224 = pi39 & ~n64246;
  assign n33225 = ~n64242 & n33224;
  assign n33226 = n32119 & n32994;
  assign n33227 = ~pi168 & ~n32116;
  assign n33228 = pi168 & ~n64180;
  assign n33229 = ~pi151 & ~n33228;
  assign n33230 = ~pi151 & ~n33227;
  assign n33231 = ~n33228 & n33230;
  assign n33232 = ~n33227 & n33229;
  assign n33233 = ~n33226 & ~n64247;
  assign n33234 = n32112 & ~n33233;
  assign n33235 = pi150 & ~n33234;
  assign n33236 = ~pi151 & n32092;
  assign n33237 = n32095 & ~n33236;
  assign n33238 = ~pi168 & ~n33237;
  assign n33239 = ~pi151 & n32101;
  assign n33240 = n32104 & ~n33239;
  assign n33241 = n33016 & ~n33240;
  assign n33242 = ~pi150 & ~n33241;
  assign n33243 = ~n33238 & n33242;
  assign n33244 = ~n33235 & ~n33243;
  assign n33245 = ~n2814 & ~n32749;
  assign n33246 = pi299 & ~n33245;
  assign n33247 = ~n33244 & n33246;
  assign n33248 = pi173 & n64197;
  assign n33249 = ~pi173 & n2751;
  assign n33250 = n32116 & n33249;
  assign n33251 = ~n33248 & ~n33250;
  assign n33252 = ~pi190 & n2814;
  assign n33253 = ~n33251 & n33252;
  assign n33254 = ~pi173 & pi190;
  assign n33255 = n32127 & n33254;
  assign n33256 = pi185 & ~n33255;
  assign n33257 = ~n33253 & n33256;
  assign n33258 = ~pi173 & n32092;
  assign n33259 = n32152 & ~n33258;
  assign n33260 = ~pi190 & ~n33259;
  assign n33261 = pi173 & n32156;
  assign n33262 = pi190 & ~n33261;
  assign n33263 = pi190 & n32827;
  assign n33264 = ~n33261 & n33263;
  assign n33265 = n32827 & n33262;
  assign n33266 = ~pi185 & ~n64248;
  assign n33267 = n32827 & ~n33261;
  assign n33268 = pi190 & ~n33267;
  assign n33269 = ~pi190 & n32152;
  assign n33270 = ~n33258 & n33269;
  assign n33271 = ~n33268 & ~n33270;
  assign n33272 = ~pi185 & ~n33271;
  assign n33273 = ~n33260 & n33266;
  assign n33274 = ~n33257 & ~n64249;
  assign n33275 = ~n2814 & ~n32823;
  assign n33276 = ~pi299 & ~n33275;
  assign n33277 = ~n33274 & n33276;
  assign n33278 = ~n33247 & ~n33277;
  assign n33279 = pi232 & ~n33278;
  assign n33280 = n64148 & ~n32735;
  assign n33281 = ~pi232 & ~n32092;
  assign n33282 = ~n33280 & n33281;
  assign n33283 = ~pi39 & ~n33282;
  assign n33284 = ~n33279 & n33283;
  assign n33285 = ~n33225 & ~n33284;
  assign n33286 = ~pi38 & ~n33285;
  assign n33287 = n32992 & ~n33286;
  assign n33288 = ~n33123 & ~n64238;
  assign n33289 = ~n33287 & n33288;
  assign n33290 = n6793 & ~n33289;
  assign n33291 = n30571 & ~n33135;
  assign n33292 = n62380 & n33291;
  assign n33293 = n33125 & ~n33292;
  assign n33294 = ~n33123 & ~n33293;
  assign n33295 = n32018 & ~n33294;
  assign n33296 = ~n33132 & ~n33295;
  assign n33297 = ~n33290 & n33296;
  assign n33298 = ~pi54 & ~n33297;
  assign n33299 = ~n32983 & ~n33298;
  assign n33300 = ~pi74 & ~n33299;
  assign n33301 = n32976 & ~n33300;
  assign n33302 = pi54 & n32940;
  assign n33303 = n64081 & ~n33150;
  assign n33304 = ~n33302 & n33303;
  assign n33305 = n62380 & n33304;
  assign n33306 = n32958 & ~n33305;
  assign n33307 = n33147 & ~n33306;
  assign n33308 = n3470 & ~n33307;
  assign n33309 = ~n33301 & n33308;
  assign n33310 = n32961 & ~n33309;
  assign n33311 = ~n64227 & ~n33310;
  assign n33312 = ~pi118 & n33311;
  assign n33313 = ~n33162 & ~n33312;
  assign n33314 = ~n33161 & n33313;
  assign n33315 = ~pi118 & ~n32294;
  assign n33316 = n33160 & n33315;
  assign n33317 = n33311 & ~n33315;
  assign n33318 = n33162 & ~n33317;
  assign n33319 = ~n33316 & n33318;
  assign n33320 = ~n33314 & ~n33319;
  assign n33321 = ~pi34 & n32296;
  assign n33322 = ~pi33 & ~n33321;
  assign n33323 = pi149 & pi157;
  assign n33324 = n31354 & ~n33323;
  assign n33325 = pi232 & n33324;
  assign n33326 = pi75 & ~n33325;
  assign n33327 = pi100 & ~n33325;
  assign n33328 = ~n33326 & ~n33327;
  assign n33329 = ~n2765 & ~n33325;
  assign n33330 = pi169 & n2815;
  assign n33331 = pi169 & n31366;
  assign n33332 = n2765 & n33330;
  assign n33333 = n64250 & ~n64251;
  assign n33334 = pi74 & ~n33333;
  assign n33335 = pi164 & n2815;
  assign n33336 = pi164 & n31366;
  assign n33337 = n2765 & n33335;
  assign n33338 = n64250 & ~n64252;
  assign n33339 = ~pi74 & ~n33338;
  assign n33340 = ~n3472 & ~n33339;
  assign n33341 = ~n3472 & ~n33334;
  assign n33342 = ~n33339 & n33341;
  assign n33343 = ~n33334 & n33340;
  assign n33344 = pi178 & pi183;
  assign n33345 = n31399 & ~n33344;
  assign n33346 = ~pi299 & ~n33345;
  assign n33347 = pi299 & ~n33324;
  assign n33348 = pi232 & ~n33347;
  assign n33349 = pi232 & ~n33346;
  assign n33350 = ~n33347 & n33349;
  assign n33351 = ~n33346 & n33348;
  assign n33352 = pi100 & ~n64254;
  assign n33353 = pi75 & ~n64254;
  assign n33354 = ~n33352 & ~n33353;
  assign n33355 = pi191 & ~pi299;
  assign n33356 = pi169 & pi299;
  assign n33357 = ~n33355 & ~n33356;
  assign n33358 = n31366 & ~n33357;
  assign n33359 = n33354 & ~n33358;
  assign n33360 = pi74 & ~n33359;
  assign n33361 = ~pi55 & ~n33360;
  assign n33362 = ~pi186 & ~pi299;
  assign n33363 = ~pi164 & pi299;
  assign n33364 = ~n33362 & ~n33363;
  assign n33365 = n2815 & n33364;
  assign n33366 = n2765 & n33365;
  assign n33367 = n33354 & ~n33366;
  assign n33368 = pi54 & ~n33367;
  assign n33369 = ~pi186 & ~n64172;
  assign n33370 = pi186 & ~n31980;
  assign n33371 = pi164 & ~n33370;
  assign n33372 = ~n33369 & n33371;
  assign n33373 = ~pi164 & pi186;
  assign n33374 = n31978 & n33373;
  assign n33375 = ~n33372 & ~n33374;
  assign n33376 = pi38 & ~n33375;
  assign n33377 = ~pi152 & n31903;
  assign n33378 = ~pi154 & ~n31899;
  assign n33379 = ~pi154 & ~n33377;
  assign n33380 = ~n31899 & n33379;
  assign n33381 = ~n33377 & n33378;
  assign n33382 = pi152 & n31914;
  assign n33383 = n31895 & ~n33382;
  assign n33384 = pi154 & ~n33383;
  assign n33385 = n31886 & ~n33384;
  assign n33386 = ~n64255 & n33385;
  assign n33387 = n31908 & ~n33386;
  assign n33388 = ~pi176 & ~pi299;
  assign n33389 = n31939 & n33388;
  assign n33390 = ~pi174 & ~n31928;
  assign n33391 = ~pi299 & ~n33390;
  assign n33392 = ~n31952 & n33391;
  assign n33393 = pi174 & n64168;
  assign n33394 = ~n31928 & ~n33393;
  assign n33395 = ~pi299 & ~n33394;
  assign n33396 = n31953 & ~n33390;
  assign n33397 = ~n33389 & ~n64256;
  assign n33398 = ~n33387 & n33397;
  assign n33399 = pi232 & ~n33398;
  assign n33400 = pi39 & ~n31966;
  assign n33401 = ~pi176 & pi232;
  assign n33402 = ~n33387 & ~n64256;
  assign n33403 = ~pi299 & n31939;
  assign n33404 = n33402 & ~n33403;
  assign n33405 = n33401 & ~n33404;
  assign n33406 = pi176 & pi232;
  assign n33407 = ~n33402 & n33406;
  assign n33408 = n33400 & ~n33407;
  assign n33409 = ~n33405 & n33408;
  assign n33410 = ~n33399 & n33400;
  assign n33411 = pi183 & n31601;
  assign n33412 = ~pi183 & n31614;
  assign n33413 = pi174 & ~n33412;
  assign n33414 = pi183 & ~n31601;
  assign n33415 = ~pi183 & ~n31614;
  assign n33416 = ~n33414 & ~n33415;
  assign n33417 = pi174 & ~n33416;
  assign n33418 = ~n33411 & n33413;
  assign n33419 = ~pi183 & ~n31681;
  assign n33420 = pi183 & ~n31628;
  assign n33421 = ~n33419 & ~n33420;
  assign n33422 = ~pi174 & ~n33421;
  assign n33423 = pi180 & ~n33422;
  assign n33424 = pi180 & ~n64258;
  assign n33425 = ~n33422 & n33424;
  assign n33426 = ~n64258 & n33423;
  assign n33427 = ~pi95 & n33421;
  assign n33428 = ~pi174 & ~n31443;
  assign n33429 = ~n33427 & n33428;
  assign n33430 = pi183 & n2814;
  assign n33431 = ~n31526 & ~n33430;
  assign n33432 = pi183 & n31589;
  assign n33433 = pi174 & ~n33432;
  assign n33434 = ~n33431 & n33433;
  assign n33435 = ~pi180 & ~n33434;
  assign n33436 = ~n33429 & n33435;
  assign n33437 = ~n64259 & ~n33436;
  assign n33438 = ~pi193 & ~n33437;
  assign n33439 = ~pi183 & ~n31558;
  assign n33440 = pi183 & ~n31569;
  assign n33441 = ~pi180 & ~n33440;
  assign n33442 = ~n33439 & n33441;
  assign n33443 = ~pi183 & ~n31608;
  assign n33444 = pi183 & ~n31598;
  assign n33445 = pi180 & ~n33444;
  assign n33446 = ~n33443 & n33445;
  assign n33447 = pi174 & ~n33446;
  assign n33448 = ~n33442 & n33447;
  assign n33449 = pi183 & n31630;
  assign n33450 = ~pi183 & ~n31662;
  assign n33451 = pi180 & ~n33450;
  assign n33452 = ~n33449 & n33451;
  assign n33453 = ~pi183 & n31697;
  assign n33454 = pi183 & n31709;
  assign n33455 = ~n33453 & ~n33454;
  assign n33456 = n2814 & ~n33455;
  assign n33457 = ~pi180 & ~n31527;
  assign n33458 = ~n33456 & n33457;
  assign n33459 = ~pi174 & ~n33458;
  assign n33460 = ~n33452 & n33459;
  assign n33461 = pi193 & ~n33460;
  assign n33462 = pi174 & ~n33444;
  assign n33463 = ~n33443 & n33462;
  assign n33464 = ~pi174 & ~n33450;
  assign n33465 = ~pi174 & ~n33449;
  assign n33466 = ~n33450 & n33465;
  assign n33467 = ~n33449 & n33464;
  assign n33468 = pi180 & ~n64260;
  assign n33469 = pi180 & ~n33463;
  assign n33470 = ~n64260 & n33469;
  assign n33471 = ~n33463 & n33468;
  assign n33472 = pi174 & ~n33440;
  assign n33473 = ~n33439 & n33472;
  assign n33474 = ~pi174 & ~n31527;
  assign n33475 = ~pi183 & n31699;
  assign n33476 = pi183 & ~n31711;
  assign n33477 = ~pi174 & ~n33476;
  assign n33478 = ~n33475 & n33477;
  assign n33479 = ~pi174 & ~n33475;
  assign n33480 = ~n33476 & n33479;
  assign n33481 = ~n33456 & n33474;
  assign n33482 = ~pi180 & ~n64262;
  assign n33483 = ~n33473 & n33482;
  assign n33484 = pi193 & ~n33483;
  assign n33485 = ~n64261 & n33484;
  assign n33486 = pi193 & ~n64261;
  assign n33487 = ~n33483 & n33486;
  assign n33488 = ~n33448 & n33461;
  assign n33489 = ~n33438 & ~n64263;
  assign n33490 = ~pi193 & ~n33436;
  assign n33491 = ~n64259 & n33490;
  assign n33492 = ~n64261 & ~n33483;
  assign n33493 = pi193 & ~n33492;
  assign n33494 = ~pi299 & ~n33493;
  assign n33495 = ~n33491 & n33494;
  assign n33496 = ~pi299 & ~n33489;
  assign n33497 = pi158 & pi299;
  assign n33498 = ~pi152 & ~n31773;
  assign n33499 = pi152 & ~n31765;
  assign n33500 = ~pi172 & ~n33499;
  assign n33501 = ~pi172 & ~n33498;
  assign n33502 = ~n33499 & n33501;
  assign n33503 = ~n33498 & n33500;
  assign n33504 = ~pi152 & n31776;
  assign n33505 = pi152 & ~n31767;
  assign n33506 = pi172 & ~n33505;
  assign n33507 = pi172 & ~n33504;
  assign n33508 = ~n33505 & n33507;
  assign n33509 = ~n33504 & n33506;
  assign n33510 = ~n64265 & ~n64266;
  assign n33511 = n33497 & ~n33510;
  assign n33512 = ~pi158 & pi299;
  assign n33513 = ~pi152 & ~n31795;
  assign n33514 = pi152 & ~n31785;
  assign n33515 = pi172 & ~n33514;
  assign n33516 = pi172 & ~n33513;
  assign n33517 = ~n33514 & n33516;
  assign n33518 = ~n33513 & n33515;
  assign n33519 = pi152 & n31787;
  assign n33520 = ~pi152 & n31793;
  assign n33521 = ~pi172 & ~n33520;
  assign n33522 = ~pi172 & ~n33519;
  assign n33523 = ~n33520 & n33522;
  assign n33524 = ~n33519 & n33521;
  assign n33525 = ~n64267 & ~n64268;
  assign n33526 = n33512 & ~n33525;
  assign n33527 = ~n33511 & ~n33526;
  assign n33528 = pi149 & ~n33527;
  assign n33529 = pi152 & n31827;
  assign n33530 = ~pi152 & ~n31807;
  assign n33531 = ~pi172 & ~n33530;
  assign n33532 = ~pi172 & ~n33529;
  assign n33533 = ~n33530 & n33532;
  assign n33534 = ~n33529 & n33531;
  assign n33535 = pi152 & ~n31823;
  assign n33536 = ~pi152 & ~n31814;
  assign n33537 = pi172 & ~n33536;
  assign n33538 = ~n33535 & n33537;
  assign n33539 = ~n64269 & ~n33538;
  assign n33540 = n33497 & ~n33539;
  assign n33541 = pi152 & ~n31834;
  assign n33542 = ~pi152 & ~n31837;
  assign n33543 = pi172 & ~n33542;
  assign n33544 = ~n33541 & n33543;
  assign n33545 = ~n31764 & n33512;
  assign n33546 = ~pi152 & ~n31843;
  assign n33547 = pi152 & ~n31763;
  assign n33548 = ~pi172 & ~n33547;
  assign n33549 = ~pi172 & ~n33546;
  assign n33550 = ~n33547 & n33549;
  assign n33551 = ~n33546 & n33548;
  assign n33552 = n33545 & ~n64270;
  assign n33553 = pi152 & n31763;
  assign n33554 = ~pi152 & n31843;
  assign n33555 = ~pi172 & ~n33554;
  assign n33556 = ~n33553 & n33555;
  assign n33557 = pi152 & n31834;
  assign n33558 = ~pi152 & n31837;
  assign n33559 = pi172 & ~n33558;
  assign n33560 = ~n33557 & n33559;
  assign n33561 = ~n33556 & ~n33560;
  assign n33562 = n33545 & ~n33561;
  assign n33563 = ~n33544 & n33552;
  assign n33564 = ~n33540 & ~n64271;
  assign n33565 = ~pi149 & ~n33564;
  assign n33566 = ~pi149 & ~n64271;
  assign n33567 = ~n33540 & n33566;
  assign n33568 = pi149 & ~n33526;
  assign n33569 = pi149 & ~n33511;
  assign n33570 = ~n33526 & n33569;
  assign n33571 = ~n33511 & n33568;
  assign n33572 = ~n33567 & ~n64272;
  assign n33573 = ~n33528 & ~n33565;
  assign n33574 = ~n64264 & ~n64273;
  assign n33575 = pi232 & ~n33574;
  assign n33576 = ~pi39 & ~n31524;
  assign n33577 = ~n33575 & n33576;
  assign n33578 = ~n64257 & ~n33577;
  assign n33579 = ~pi38 & ~n33578;
  assign n33580 = ~n33376 & ~n33579;
  assign n33581 = ~pi100 & ~n33580;
  assign n33582 = ~pi87 & ~n33352;
  assign n33583 = ~n33581 & n33582;
  assign n33584 = pi38 & n33365;
  assign n33585 = ~pi100 & n33584;
  assign n33586 = ~n33352 & ~n33585;
  assign n33587 = pi87 & ~n32703;
  assign n33588 = n33586 & n33587;
  assign n33589 = n6793 & ~n33588;
  assign n33590 = ~n33583 & n33589;
  assign n33591 = ~pi154 & pi299;
  assign n33592 = ~n33388 & ~n33591;
  assign n33593 = pi232 & ~n33591;
  assign n33594 = n2814 & ~n33388;
  assign n33595 = n33593 & n33594;
  assign n33596 = n2815 & n33592;
  assign n33597 = n64176 & ~n64274;
  assign n33598 = n32703 & ~n33597;
  assign n33599 = n33586 & ~n33598;
  assign n33600 = n32018 & ~n33599;
  assign n33601 = ~n33353 & ~n33600;
  assign n33602 = ~n33590 & n33601;
  assign n33603 = ~pi54 & ~n33602;
  assign n33604 = ~n33368 & ~n33603;
  assign n33605 = ~pi74 & ~n33604;
  assign n33606 = n33361 & ~n33605;
  assign n33607 = pi55 & ~n33334;
  assign n33608 = pi54 & ~n33338;
  assign n33609 = ~pi92 & n64250;
  assign n33610 = pi38 & ~n33335;
  assign n33611 = n2765 & ~n32009;
  assign n33612 = ~pi100 & ~n32009;
  assign n33613 = ~n33610 & n33612;
  assign n33614 = ~pi75 & n33613;
  assign n33615 = ~n33610 & n33611;
  assign n33616 = pi149 & n2815;
  assign n33617 = ~pi38 & ~n33616;
  assign n33618 = n64176 & n33617;
  assign n33619 = n64275 & ~n33618;
  assign n33620 = ~pi92 & ~n33326;
  assign n33621 = n6791 & ~n33610;
  assign n33622 = ~pi39 & ~n33616;
  assign n33623 = n31887 & n33622;
  assign n33624 = n31385 & ~n33623;
  assign n33625 = ~pi38 & ~n33624;
  assign n33626 = n33621 & ~n33625;
  assign n33627 = pi87 & n33613;
  assign n33628 = ~n33327 & ~n33627;
  assign n33629 = ~n33626 & n33628;
  assign n33630 = ~pi75 & ~n33629;
  assign n33631 = n33620 & ~n33630;
  assign n33632 = n33609 & ~n33619;
  assign n33633 = pi92 & n64250;
  assign n33634 = ~n64275 & n33633;
  assign n33635 = ~pi54 & ~n33634;
  assign n33636 = ~n64276 & n33635;
  assign n33637 = n33149 & ~n33616;
  assign n33638 = n33148 & ~n33637;
  assign n33639 = ~n32955 & n33335;
  assign n33640 = ~n33638 & ~n33639;
  assign n33641 = n2765 & ~n33640;
  assign n33642 = n64250 & ~n33641;
  assign n33643 = ~n33608 & ~n33636;
  assign n33644 = ~pi74 & ~n64277;
  assign n33645 = n33607 & ~n33644;
  assign n33646 = n3470 & ~n33645;
  assign n33647 = ~n33606 & n33646;
  assign n33648 = pi164 & ~n32955;
  assign n33649 = n31366 & n33648;
  assign n33650 = pi38 & n33335;
  assign n33651 = pi38 & n64252;
  assign n33652 = n2765 & n33650;
  assign n33653 = n64250 & ~n64278;
  assign n33654 = ~n33608 & n33653;
  assign n33655 = n64250 & ~n33649;
  assign n33656 = ~pi74 & ~n64279;
  assign n33657 = ~n33334 & ~n33656;
  assign n33658 = ~n3470 & ~n33657;
  assign n33659 = n3472 & ~n33658;
  assign n33660 = ~n32716 & n33659;
  assign n33661 = ~n33647 & n33660;
  assign n33662 = ~n64253 & ~n33661;
  assign n33663 = ~n33322 & ~n33662;
  assign n33664 = pi39 & pi232;
  assign n33665 = pi154 & ~n32204;
  assign n33666 = ~pi154 & ~n32215;
  assign n33667 = ~pi152 & ~n33666;
  assign n33668 = ~n33665 & n33667;
  assign n33669 = pi152 & pi154;
  assign n33670 = n64187 & n33669;
  assign n33671 = ~n33668 & ~n33670;
  assign n33672 = n64234 & ~n33671;
  assign n33673 = ~pi174 & ~n64190;
  assign n33674 = pi174 & ~n32228;
  assign n33675 = pi176 & ~n33674;
  assign n33676 = ~n33673 & n33675;
  assign n33677 = ~pi174 & ~pi176;
  assign n33678 = n64192 & n33677;
  assign n33679 = ~n33676 & ~n33678;
  assign n33680 = ~pi299 & ~n33679;
  assign n33681 = ~n33672 & ~n33680;
  assign n33682 = ~pi174 & n64192;
  assign n33683 = ~pi299 & ~n33682;
  assign n33684 = n33401 & ~n33683;
  assign n33685 = ~pi174 & n64190;
  assign n33686 = pi174 & n32228;
  assign n33687 = ~pi299 & ~n33686;
  assign n33688 = ~n33685 & n33687;
  assign n33689 = n33406 & ~n33688;
  assign n33690 = ~n33684 & ~n33689;
  assign n33691 = n31886 & ~n33671;
  assign n33692 = pi299 & ~n33691;
  assign n33693 = pi39 & ~n33692;
  assign n33694 = ~n33690 & n33693;
  assign n33695 = pi176 & ~n33688;
  assign n33696 = ~pi176 & ~n33683;
  assign n33697 = ~n33695 & ~n33696;
  assign n33698 = n33664 & ~n33697;
  assign n33699 = pi39 & ~n33690;
  assign n33700 = ~n33692 & n64281;
  assign n33701 = n33664 & ~n33681;
  assign n33702 = ~n32823 & n33430;
  assign n33703 = ~pi183 & n32117;
  assign n33704 = pi193 & ~n33703;
  assign n33705 = ~n33702 & n33704;
  assign n33706 = ~n32152 & n33430;
  assign n33707 = ~pi183 & n32121;
  assign n33708 = ~pi193 & ~n33707;
  assign n33709 = ~n33706 & n33708;
  assign n33710 = ~pi174 & ~n33709;
  assign n33711 = ~n33705 & n33710;
  assign n33712 = pi183 & n32827;
  assign n33713 = ~pi183 & n32127;
  assign n33714 = pi193 & ~n33713;
  assign n33715 = ~n33712 & n33714;
  assign n33716 = ~n32156 & n33430;
  assign n33717 = ~pi193 & ~n33716;
  assign n33718 = pi174 & ~n33717;
  assign n33719 = pi183 & ~n32827;
  assign n33720 = ~pi183 & ~n32127;
  assign n33721 = pi193 & ~n33720;
  assign n33722 = ~n33719 & n33721;
  assign n33723 = ~pi193 & n33430;
  assign n33724 = ~n32156 & n33723;
  assign n33725 = ~n33722 & ~n33724;
  assign n33726 = pi174 & ~n33725;
  assign n33727 = ~n33715 & n33718;
  assign n33728 = pi180 & n32135;
  assign n33729 = ~pi299 & ~n33728;
  assign n33730 = ~n64282 & n33729;
  assign n33731 = ~pi174 & ~n33703;
  assign n33732 = ~n33702 & n33731;
  assign n33733 = pi174 & ~n33713;
  assign n33734 = ~n33712 & n33733;
  assign n33735 = ~n33732 & ~n33734;
  assign n33736 = pi193 & ~n33735;
  assign n33737 = ~pi174 & n32152;
  assign n33738 = pi174 & n32156;
  assign n33739 = n33430 & ~n33738;
  assign n33740 = ~n33737 & n33739;
  assign n33741 = ~pi174 & ~pi183;
  assign n33742 = n32121 & n33741;
  assign n33743 = ~pi193 & ~n33742;
  assign n33744 = ~n33740 & n33743;
  assign n33745 = ~n33736 & ~n33744;
  assign n33746 = n33729 & ~n33745;
  assign n33747 = ~n33711 & n33730;
  assign n33748 = pi172 & n32092;
  assign n33749 = ~pi152 & n32095;
  assign n33750 = ~n33748 & n33749;
  assign n33751 = pi149 & n2814;
  assign n33752 = pi172 & n32101;
  assign n33753 = pi152 & n32104;
  assign n33754 = pi152 & ~n33752;
  assign n33755 = n32104 & n33754;
  assign n33756 = ~n33752 & n33753;
  assign n33757 = n33751 & ~n64284;
  assign n33758 = n32104 & ~n33752;
  assign n33759 = pi152 & ~n33758;
  assign n33760 = n32095 & ~n33748;
  assign n33761 = ~pi152 & ~n33760;
  assign n33762 = ~n33759 & ~n33761;
  assign n33763 = n33751 & ~n33762;
  assign n33764 = ~n33750 & n33757;
  assign n33765 = ~pi152 & n32117;
  assign n33766 = pi172 & ~n32127;
  assign n33767 = ~n33765 & n33766;
  assign n33768 = ~pi152 & n32121;
  assign n33769 = ~pi172 & ~n33768;
  assign n33770 = ~pi149 & ~n33769;
  assign n33771 = ~n32127 & ~n33765;
  assign n33772 = pi172 & ~n33771;
  assign n33773 = ~pi152 & ~pi172;
  assign n33774 = n32121 & n33773;
  assign n33775 = ~n33772 & ~n33774;
  assign n33776 = ~pi149 & ~n33775;
  assign n33777 = ~n33767 & n33770;
  assign n33778 = pi158 & n32135;
  assign n33779 = pi299 & ~n33778;
  assign n33780 = ~n64286 & n33779;
  assign n33781 = ~n64285 & n33780;
  assign n33782 = n32271 & ~n33781;
  assign n33783 = n32271 & ~n64283;
  assign n33784 = ~n33781 & n33783;
  assign n33785 = ~n64283 & n33782;
  assign n33786 = ~n64280 & ~n64287;
  assign n33787 = ~pi38 & ~n33786;
  assign n33788 = ~pi87 & ~n33376;
  assign n33789 = ~n33787 & n33788;
  assign n33790 = pi87 & ~n33584;
  assign n33791 = ~pi100 & ~n33790;
  assign n33792 = ~n33789 & n33791;
  assign n33793 = ~n33352 & ~n33792;
  assign n33794 = n6793 & ~n33793;
  assign n33795 = n62951 & n64274;
  assign n33796 = n7356 & n33795;
  assign n33797 = n33586 & ~n33796;
  assign n33798 = n32018 & ~n33797;
  assign n33799 = ~n33353 & ~n33798;
  assign n33800 = ~n33794 & n33799;
  assign n33801 = ~pi54 & ~n33800;
  assign n33802 = ~n33368 & ~n33801;
  assign n33803 = ~pi74 & ~n33802;
  assign n33804 = n33361 & ~n33803;
  assign n33805 = pi149 & n2579;
  assign n33806 = n9735 & n33805;
  assign n33807 = n7356 & n33806;
  assign n33808 = ~n33648 & ~n33807;
  assign n33809 = n31366 & ~n33808;
  assign n33810 = n30571 & n33616;
  assign n33811 = n62380 & n33810;
  assign n33812 = ~n33650 & ~n33811;
  assign n33813 = n2765 & ~n33812;
  assign n33814 = n7356 & n33616;
  assign n33815 = ~pi38 & ~n33814;
  assign n33816 = n33621 & ~n33815;
  assign n33817 = pi38 & pi87;
  assign n33818 = ~pi100 & n33817;
  assign n33819 = n3011 & n33650;
  assign n33820 = n33335 & n33818;
  assign n33821 = ~n33327 & ~n64288;
  assign n33822 = ~n33816 & n33821;
  assign n33823 = ~pi75 & ~n33822;
  assign n33824 = n33620 & ~n33823;
  assign n33825 = n33609 & ~n33813;
  assign n33826 = n33633 & ~n64278;
  assign n33827 = pi92 & n33653;
  assign n33828 = ~pi54 & ~n64290;
  assign n33829 = ~n64289 & n33828;
  assign n33830 = ~n33608 & ~n33829;
  assign n33831 = n64250 & ~n33809;
  assign n33832 = ~pi74 & ~n64291;
  assign n33833 = n33607 & ~n33832;
  assign n33834 = n3470 & ~n33833;
  assign n33835 = ~n33804 & n33834;
  assign n33836 = n33659 & ~n33835;
  assign n33837 = ~n64253 & ~n33836;
  assign n33838 = n33322 & ~n33837;
  assign n33839 = ~pi954 & ~n33838;
  assign n33840 = ~n33663 & n33839;
  assign n33841 = ~pi33 & ~n33662;
  assign n33842 = pi33 & ~n33837;
  assign n33843 = pi954 & ~n33842;
  assign n33844 = ~n33841 & n33843;
  assign po191 = ~n33840 & ~n33844;
  assign n33846 = n3036 & n5427;
  assign n33847 = n2580 & n31335;
  assign n33848 = n30915 & ~n33847;
  assign n33849 = n2580 & n31290;
  assign n33850 = n3318 & ~n33849;
  assign n33851 = n62455 & ~n33850;
  assign n33852 = n62455 & ~n33848;
  assign n33853 = ~n33850 & n33852;
  assign n33854 = ~n33848 & n33851;
  assign n33855 = ~n33846 & ~n64292;
  assign n33856 = pi57 & ~n30591;
  assign n33857 = ~pi55 & ~n30598;
  assign n33858 = ~pi100 & ~n30606;
  assign n33859 = ~pi32 & ~n6864;
  assign n33860 = ~pi40 & ~n30618;
  assign n33861 = ~pi91 & n2743;
  assign n33862 = ~pi91 & n2715;
  assign n33863 = n2743 & n33862;
  assign n33864 = n2715 & n33861;
  assign n33865 = n2856 & n64293;
  assign n33866 = n2658 & n2783;
  assign n33867 = pi96 & n64294;
  assign n33868 = ~pi72 & ~n33867;
  assign n33869 = pi108 & ~n6854;
  assign n33870 = ~pi46 & ~n33869;
  assign n33871 = ~pi86 & pi94;
  assign n33872 = n2861 & n33871;
  assign n33873 = ~pi97 & ~n33872;
  assign n33874 = ~n6821 & ~n30705;
  assign n33875 = pi64 & ~n2630;
  assign n33876 = n2601 & ~n30676;
  assign n33877 = n30660 & ~n33876;
  assign n33878 = ~pi84 & ~n33877;
  assign n33879 = ~n30681 & ~n33878;
  assign n33880 = n30652 & ~n33879;
  assign n33881 = pi111 & ~n30654;
  assign n33882 = ~pi82 & ~n33881;
  assign n33883 = ~n30682 & n33882;
  assign n33884 = ~n33880 & n33883;
  assign n33885 = n6806 & ~n64094;
  assign n33886 = ~n33884 & n33885;
  assign n33887 = pi67 & ~n62344;
  assign n33888 = n2598 & n30654;
  assign n33889 = pi36 & ~n33888;
  assign n33890 = ~n33887 & ~n33889;
  assign n33891 = ~n33886 & n33890;
  assign n33892 = n6810 & ~n33891;
  assign n33893 = n30649 & ~n33892;
  assign n33894 = ~pi71 & ~n64095;
  assign n33895 = ~n33893 & n33894;
  assign n33896 = n30694 & ~n33895;
  assign n33897 = ~pi107 & ~n33896;
  assign n33898 = pi65 & ~pi71;
  assign n33899 = n2610 & n33898;
  assign n33900 = n33897 & ~n33899;
  assign n33901 = pi107 & ~n2625;
  assign n33902 = ~pi63 & ~n33901;
  assign n33903 = ~n33900 & n33902;
  assign n33904 = ~pi64 & ~n33903;
  assign n33905 = ~n33875 & ~n33904;
  assign n33906 = n2614 & ~n33905;
  assign n33907 = ~n33897 & n33902;
  assign n33908 = pi63 & ~pi107;
  assign n33909 = n2625 & n33908;
  assign n33910 = ~pi64 & ~n33909;
  assign n33911 = ~n33907 & n33910;
  assign n33912 = ~n33875 & ~n33911;
  assign n33913 = n33906 & ~n33912;
  assign n33914 = n33874 & ~n33913;
  assign n33915 = n2611 & ~n33914;
  assign n33916 = pi98 & ~n62358;
  assign n33917 = ~pi77 & ~n33916;
  assign n33918 = ~n6874 & n33917;
  assign n33919 = ~n33915 & n33918;
  assign n33920 = n2682 & n2683;
  assign n33921 = n33919 & n33920;
  assign n33922 = n33873 & ~n33921;
  assign n33923 = ~n30937 & ~n33922;
  assign n33924 = ~pi108 & ~n33923;
  assign n33925 = n33870 & ~n33924;
  assign n33926 = ~pi110 & n30750;
  assign n33927 = ~n33925 & n33926;
  assign n33928 = ~pi109 & n2671;
  assign n33929 = pi110 & ~n33928;
  assign n33930 = ~n30748 & ~n33929;
  assign n33931 = ~n33927 & n33930;
  assign n33932 = ~pi47 & ~n33931;
  assign n33933 = n6848 & ~n33932;
  assign n33934 = n32077 & ~n33933;
  assign n33935 = ~n30627 & ~n33934;
  assign n33936 = ~pi93 & ~n33935;
  assign n33937 = ~n2661 & ~n33936;
  assign n33938 = ~pi35 & ~n33937;
  assign n33939 = pi35 & ~n62363;
  assign n33940 = ~pi70 & ~n33939;
  assign n33941 = ~n33938 & n33940;
  assign n33942 = ~pi51 & ~n33941;
  assign n33943 = n2733 & ~n33942;
  assign n33944 = n33868 & ~n33943;
  assign n33945 = n33860 & ~n33944;
  assign n33946 = n33859 & ~n33945;
  assign n33947 = ~pi93 & n30624;
  assign n33948 = pi841 & n62363;
  assign n33949 = ~pi35 & ~pi40;
  assign n33950 = ~pi35 & n62376;
  assign n33951 = ~pi40 & n62382;
  assign n33952 = n62375 & n33949;
  assign n33953 = n64295 & n64296;
  assign n33954 = pi32 & ~n33953;
  assign n33955 = n64148 & ~n33954;
  assign n33956 = n2726 & n30617;
  assign n33957 = pi32 & ~n33956;
  assign n33958 = ~n64148 & ~n33957;
  assign n33959 = ~n33955 & ~n33958;
  assign n33960 = ~n33946 & ~n33959;
  assign n33961 = ~pi95 & ~n33960;
  assign n33962 = pi95 & ~n2795;
  assign n33963 = ~pi39 & ~n33962;
  assign n33964 = ~n33961 & n33963;
  assign n33965 = n31888 & n33084;
  assign n33966 = pi221 & n31888;
  assign n33967 = n33209 & n33966;
  assign n33968 = ~n2920 & n33084;
  assign n33969 = n31888 & n33968;
  assign n33970 = ~n2920 & n33965;
  assign n33971 = n62380 & ~n64297;
  assign n33972 = ~pi215 & ~n33971;
  assign n33973 = pi1093 & ~n2929;
  assign n33974 = pi824 & ~pi1091;
  assign n33975 = n33973 & ~n33974;
  assign n33976 = pi829 & ~n33973;
  assign n33977 = ~pi824 & ~n33976;
  assign n33978 = ~n6899 & ~n33977;
  assign n33979 = ~n2583 & ~n33975;
  assign n33980 = n31889 & n64298;
  assign n33981 = ~n2814 & ~n33980;
  assign n33982 = ~n2908 & ~n33981;
  assign n33983 = n62380 & ~n33982;
  assign n33984 = ~n2908 & n32270;
  assign n33985 = ~n33983 & ~n33984;
  assign n33986 = n62393 & ~n33985;
  assign n33987 = ~n2953 & n33980;
  assign n33988 = n62380 & ~n33987;
  assign n33989 = ~n62393 & n33988;
  assign n33990 = pi215 & ~n33989;
  assign n33991 = ~n33986 & n33990;
  assign n33992 = ~n33972 & ~n33991;
  assign n33993 = pi299 & ~n33992;
  assign n33994 = n2971 & n33985;
  assign n33995 = ~n2971 & ~n33988;
  assign n33996 = pi223 & ~n33995;
  assign n33997 = ~n33994 & n33996;
  assign n33998 = pi224 & n31888;
  assign n33999 = n30839 & n33998;
  assign n34000 = n31888 & n33075;
  assign n34001 = ~n2973 & n34000;
  assign n34002 = n31888 & n64244;
  assign n34003 = ~pi223 & ~n64299;
  assign n34004 = n62380 & n34003;
  assign n34005 = ~pi299 & ~n34004;
  assign n34006 = ~n33997 & n34005;
  assign n34007 = pi39 & ~n34006;
  assign n34008 = ~n33993 & n34007;
  assign n34009 = ~pi38 & ~n34008;
  assign n34010 = ~n33961 & ~n33962;
  assign n34011 = ~pi39 & ~n34010;
  assign n34012 = n2971 & ~n33985;
  assign n34013 = ~n2971 & n33988;
  assign n34014 = pi223 & ~n34013;
  assign n34015 = ~n34012 & n34014;
  assign n34016 = n62380 & ~n64299;
  assign n34017 = ~pi223 & ~n34016;
  assign n34018 = ~pi299 & ~n34017;
  assign n34019 = ~n33997 & ~n34004;
  assign n34020 = ~pi299 & ~n34019;
  assign n34021 = ~n34015 & n34018;
  assign n34022 = pi299 & ~n33972;
  assign n34023 = ~n33991 & n34022;
  assign n34024 = pi39 & ~n34023;
  assign n34025 = pi39 & ~n64300;
  assign n34026 = ~n34023 & n34025;
  assign n34027 = ~n64300 & n34024;
  assign n34028 = ~n34011 & ~n64301;
  assign n34029 = ~pi38 & ~n34028;
  assign n34030 = ~n33964 & n34009;
  assign n34031 = n33858 & ~n64302;
  assign n34032 = n30887 & ~n34031;
  assign n34033 = pi87 & ~n30595;
  assign n34034 = ~pi75 & ~n34033;
  assign n34035 = n2579 & n34034;
  assign n34036 = ~n34032 & n34035;
  assign n34037 = ~pi74 & ~n34036;
  assign n34038 = n33857 & ~n34037;
  assign n34039 = ~pi56 & ~n34038;
  assign n34040 = ~pi55 & ~pi74;
  assign n34041 = n30584 & n30595;
  assign n34042 = n64087 & n34040;
  assign n34043 = pi56 & ~n64303;
  assign n34044 = ~n34039 & ~n34043;
  assign n34045 = ~pi62 & ~n34044;
  assign n34046 = ~pi56 & n30584;
  assign n34047 = n30595 & n34046;
  assign n34048 = pi62 & ~n34047;
  assign n34049 = ~pi59 & ~n34048;
  assign n34050 = ~n34045 & n34049;
  assign n34051 = ~pi57 & ~n34050;
  assign po167 = ~n33856 & ~n34051;
  assign n34053 = ~pi228 & ~n3475;
  assign n34054 = pi57 & ~n34053;
  assign n34055 = ~n2814 & ~n2907;
  assign n34056 = ~pi907 & n2814;
  assign n34057 = ~n34055 & ~n34056;
  assign n34058 = pi30 & pi228;
  assign n34059 = ~pi228 & n62380;
  assign n34060 = n2764 & n34059;
  assign n34061 = n6791 & n34060;
  assign n34062 = ~pi100 & n34059;
  assign n34063 = n30571 & n34062;
  assign n34064 = ~pi228 & n30599;
  assign n34065 = n6794 & n64304;
  assign n34066 = ~pi54 & n6793;
  assign n34067 = n64304 & n34066;
  assign n34068 = n64086 & n34059;
  assign n34069 = ~pi74 & n64306;
  assign n34070 = ~pi228 & n64109;
  assign n34071 = ~n34058 & ~n34059;
  assign n34072 = ~pi228 & ~n64082;
  assign n34073 = ~n34071 & ~n34072;
  assign n34074 = ~n34058 & ~n64305;
  assign n34075 = n34057 & n64307;
  assign n34076 = n34054 & n34075;
  assign n34077 = ~pi602 & n2814;
  assign n34078 = ~n34055 & ~n34077;
  assign n34079 = ~pi228 & ~n30768;
  assign n34080 = ~n34058 & ~n34079;
  assign n34081 = n34078 & ~n34080;
  assign n34082 = ~pi299 & ~n34081;
  assign n34083 = ~pi299 & n30609;
  assign n34084 = ~n34082 & ~n34083;
  assign n34085 = n34058 & n34078;
  assign n34086 = ~n30746 & ~n30770;
  assign n34087 = ~pi228 & n34078;
  assign n34088 = ~n34086 & n34087;
  assign n34089 = ~n34085 & ~n34088;
  assign n34090 = n30609 & ~n34089;
  assign n34091 = ~n34084 & ~n34090;
  assign n34092 = n34057 & n34058;
  assign n34093 = pi299 & ~n34092;
  assign n34094 = n30774 & n30783;
  assign n34095 = ~n30777 & ~n30782;
  assign n34096 = n34057 & ~n34095;
  assign n34097 = n34094 & ~n34096;
  assign n34098 = ~n30779 & n34057;
  assign n34099 = ~n34094 & ~n34098;
  assign n34100 = ~pi228 & ~n34099;
  assign n34101 = ~n34097 & n34100;
  assign n34102 = n34093 & ~n34101;
  assign n34103 = pi232 & ~n34102;
  assign n34104 = pi232 & ~n34091;
  assign n34105 = ~n34102 & n34104;
  assign n34106 = ~n34091 & n34103;
  assign n34107 = ~pi228 & n34098;
  assign n34108 = n34093 & ~n34107;
  assign n34109 = ~pi232 & ~n34108;
  assign n34110 = ~n34082 & n34109;
  assign n34111 = ~n64308 & ~n34110;
  assign n34112 = ~pi39 & ~n34111;
  assign n34113 = ~pi228 & n64100;
  assign n34114 = ~n34058 & ~n34113;
  assign n34115 = n2960 & ~n34114;
  assign n34116 = ~n34058 & ~n34115;
  assign n34117 = n34057 & ~n34116;
  assign n34118 = pi299 & ~n34117;
  assign n34119 = ~pi228 & n64103;
  assign n34120 = ~n34058 & ~n34119;
  assign n34121 = n34078 & ~n34120;
  assign n34122 = ~pi299 & ~n34121;
  assign n34123 = pi39 & ~n34122;
  assign n34124 = ~n34118 & n34123;
  assign n34125 = ~pi38 & ~n34124;
  assign n34126 = ~n34112 & n34125;
  assign n34127 = pi299 & n34057;
  assign n34128 = ~pi299 & n34078;
  assign n34129 = ~n34127 & ~n34128;
  assign n34130 = ~pi39 & ~n34071;
  assign n34131 = ~n34129 & n34130;
  assign n34132 = n34058 & ~n34129;
  assign n34133 = pi38 & ~n34132;
  assign n34134 = ~n34131 & n34133;
  assign n34135 = ~n34126 & ~n34134;
  assign n34136 = ~pi100 & ~n34135;
  assign n34137 = n62380 & ~n30871;
  assign n34138 = pi683 & ~n2843;
  assign n34139 = n34137 & n34138;
  assign n34140 = ~n34055 & n34139;
  assign n34141 = n30858 & n34140;
  assign n34142 = pi252 & n32270;
  assign n34143 = ~n2907 & n34142;
  assign n34144 = n2821 & n2907;
  assign n34145 = ~n2907 & ~n34142;
  assign n34146 = ~n2821 & n2907;
  assign n34147 = ~n34145 & ~n34146;
  assign n34148 = ~n34143 & ~n34144;
  assign n34149 = pi252 & ~n30858;
  assign n34150 = n64309 & n34149;
  assign n34151 = ~n34141 & ~n34150;
  assign n34152 = ~pi228 & ~n34077;
  assign n34153 = ~n34151 & n34152;
  assign n34154 = ~pi299 & ~n34085;
  assign n34155 = ~n34153 & n34154;
  assign n34156 = ~n30860 & ~n64309;
  assign n34157 = n30860 & ~n34140;
  assign n34158 = ~pi228 & ~n34056;
  assign n34159 = ~n34157 & n34158;
  assign n34160 = ~n34156 & n34159;
  assign n34161 = n34093 & ~n34160;
  assign n34162 = n2764 & ~n34161;
  assign n34163 = ~n34155 & n34162;
  assign n34164 = ~n2764 & n34132;
  assign n34165 = pi100 & ~n34164;
  assign n34166 = ~n34163 & n34165;
  assign n34167 = ~pi87 & ~n34166;
  assign n34168 = ~n34136 & n34167;
  assign n34169 = pi87 & n34132;
  assign n34170 = ~pi75 & ~n34169;
  assign n34171 = ~n34168 & n34170;
  assign n34172 = ~n2806 & n34132;
  assign n34173 = n62951 & n34131;
  assign n34174 = ~n34172 & ~n34173;
  assign n34175 = pi75 & n34174;
  assign n34176 = ~pi92 & ~n34175;
  assign n34177 = ~n34171 & n34176;
  assign n34178 = ~pi75 & n34174;
  assign n34179 = pi75 & ~n34132;
  assign n34180 = pi92 & ~n34179;
  assign n34181 = ~n34178 & n34180;
  assign n34182 = ~pi54 & ~n34181;
  assign n34183 = ~n34177 & n34182;
  assign n34184 = n6793 & n34174;
  assign n34185 = ~n6793 & ~n34132;
  assign n34186 = ~n34184 & ~n34185;
  assign n34187 = pi54 & ~n34186;
  assign n34188 = ~pi74 & ~n34187;
  assign n34189 = ~n34183 & n34188;
  assign n34190 = ~pi54 & n34184;
  assign n34191 = ~n34066 & ~n34132;
  assign n34192 = pi74 & ~n34191;
  assign n34193 = ~n34190 & n34192;
  assign n34194 = ~pi55 & ~n34193;
  assign n34195 = ~n34189 & n34194;
  assign n34196 = pi55 & ~n34075;
  assign n34197 = n3470 & ~n34196;
  assign n34198 = ~n34195 & n34197;
  assign n34199 = ~n3470 & n34092;
  assign n34200 = ~pi59 & ~n34199;
  assign n34201 = ~n34198 & n34200;
  assign n34202 = ~pi228 & ~n3471;
  assign n34203 = n34075 & ~n34202;
  assign n34204 = pi59 & ~n34203;
  assign n34205 = ~pi57 & ~n34204;
  assign n34206 = ~n34201 & n34205;
  assign po171 = ~n34076 & ~n34206;
  assign n34208 = ~pi947 & n2814;
  assign n34209 = ~n2952 & ~n34208;
  assign n34210 = n64307 & n34209;
  assign n34211 = n34054 & n34210;
  assign n34212 = ~pi587 & n2814;
  assign n34213 = ~n2952 & ~n34212;
  assign n34214 = n34058 & n34213;
  assign n34215 = ~pi228 & n34213;
  assign n34216 = ~n34086 & n34215;
  assign n34217 = ~n34214 & ~n34216;
  assign n34218 = n30609 & ~n34217;
  assign n34219 = ~n34080 & n34213;
  assign n34220 = ~n30609 & n34219;
  assign n34221 = ~pi299 & ~n34220;
  assign n34222 = ~n34218 & n34221;
  assign n34223 = n34058 & n34209;
  assign n34224 = pi299 & ~n34223;
  assign n34225 = ~n34095 & n34209;
  assign n34226 = n34094 & ~n34225;
  assign n34227 = ~n30779 & n34209;
  assign n34228 = ~n34094 & ~n34227;
  assign n34229 = ~pi228 & ~n34228;
  assign n34230 = ~n34226 & n34229;
  assign n34231 = n34224 & ~n34230;
  assign n34232 = pi232 & ~n34231;
  assign n34233 = pi232 & ~n34222;
  assign n34234 = ~n34231 & n34233;
  assign n34235 = ~n34222 & n34232;
  assign n34236 = ~pi299 & ~n34219;
  assign n34237 = ~pi228 & n34227;
  assign n34238 = n34224 & ~n34237;
  assign n34239 = ~pi232 & ~n34238;
  assign n34240 = ~n34236 & n34239;
  assign n34241 = ~n64310 & ~n34240;
  assign n34242 = ~pi39 & ~n34241;
  assign n34243 = ~n2961 & ~n34224;
  assign n34244 = n34115 & n34209;
  assign n34245 = ~n34243 & ~n34244;
  assign n34246 = ~n34120 & n34213;
  assign n34247 = ~pi299 & ~n34246;
  assign n34248 = pi39 & ~n34247;
  assign n34249 = pi39 & ~n34245;
  assign n34250 = ~n34247 & n34249;
  assign n34251 = ~n34245 & n34248;
  assign n34252 = ~pi38 & ~n64311;
  assign n34253 = ~n34242 & n34252;
  assign n34254 = pi299 & ~n34209;
  assign n34255 = ~pi299 & ~n34213;
  assign n34256 = ~n34254 & ~n34255;
  assign n34257 = n34130 & n34256;
  assign n34258 = n34058 & n34256;
  assign n34259 = pi38 & ~n34258;
  assign n34260 = ~n34257 & n34259;
  assign n34261 = ~n34253 & ~n34260;
  assign n34262 = ~pi100 & ~n34261;
  assign n34263 = ~pi228 & n2808;
  assign n34264 = ~n2904 & ~n34142;
  assign n34265 = ~n2821 & n2904;
  assign n34266 = ~n2904 & n34142;
  assign n34267 = n2821 & n2904;
  assign n34268 = ~n34266 & ~n34267;
  assign n34269 = ~n34264 & ~n34265;
  assign n34270 = ~n34212 & ~n64312;
  assign n34271 = n34263 & ~n34270;
  assign n34272 = pi142 & n64312;
  assign n34273 = ~n2952 & n34139;
  assign n34274 = ~pi142 & ~n34273;
  assign n34275 = ~n2814 & n2904;
  assign n34276 = ~pi587 & ~n34275;
  assign n34277 = ~pi228 & ~n34276;
  assign n34278 = ~n34274 & n34277;
  assign n34279 = ~n34272 & n34278;
  assign n34280 = ~n34214 & ~n34263;
  assign n34281 = ~n34279 & n34280;
  assign n34282 = ~n34271 & ~n34281;
  assign n34283 = ~pi299 & ~n34282;
  assign n34284 = n30860 & ~n34208;
  assign n34285 = n34273 & n34284;
  assign n34286 = ~pi947 & ~n34275;
  assign n34287 = ~n30860 & ~n34286;
  assign n34288 = ~n64312 & n34287;
  assign n34289 = ~n34285 & ~n34288;
  assign n34290 = ~pi228 & ~n34289;
  assign n34291 = n34224 & ~n34290;
  assign n34292 = n2764 & ~n34291;
  assign n34293 = ~n34283 & n34292;
  assign n34294 = ~n2764 & n34258;
  assign n34295 = pi100 & ~n34294;
  assign n34296 = ~n34293 & n34295;
  assign n34297 = ~pi87 & ~n34296;
  assign n34298 = ~n34262 & n34297;
  assign n34299 = pi87 & n34258;
  assign n34300 = ~pi75 & ~n34299;
  assign n34301 = ~n34298 & n34300;
  assign n34302 = ~n2806 & n34258;
  assign n34303 = n62951 & n34257;
  assign n34304 = ~n34302 & ~n34303;
  assign n34305 = pi75 & n34304;
  assign n34306 = ~pi92 & ~n34305;
  assign n34307 = ~n34301 & n34306;
  assign n34308 = ~pi75 & n34304;
  assign n34309 = pi75 & ~n34258;
  assign n34310 = pi92 & ~n34309;
  assign n34311 = ~n34308 & n34310;
  assign n34312 = ~pi54 & ~n34311;
  assign n34313 = ~n34307 & n34312;
  assign n34314 = n6793 & n34304;
  assign n34315 = ~n6793 & ~n34258;
  assign n34316 = ~n34314 & ~n34315;
  assign n34317 = pi54 & ~n34316;
  assign n34318 = ~pi74 & ~n34317;
  assign n34319 = ~n34313 & n34318;
  assign n34320 = ~pi54 & n34314;
  assign n34321 = ~n34066 & ~n34258;
  assign n34322 = pi74 & ~n34321;
  assign n34323 = ~n34320 & n34322;
  assign n34324 = ~pi55 & ~n34323;
  assign n34325 = ~n34319 & n34324;
  assign n34326 = pi55 & ~n34210;
  assign n34327 = n3470 & ~n34326;
  assign n34328 = ~n34325 & n34327;
  assign n34329 = ~n3470 & n34223;
  assign n34330 = ~pi59 & ~n34329;
  assign n34331 = ~n34328 & n34330;
  assign n34332 = ~n34202 & n34210;
  assign n34333 = pi59 & ~n34332;
  assign n34334 = ~pi57 & ~n34333;
  assign n34335 = ~n34331 & n34334;
  assign po172 = ~n34211 & ~n34335;
  assign n34337 = pi30 & n2814;
  assign n34338 = pi228 & n34337;
  assign n34339 = pi970 & n34338;
  assign n34340 = ~pi228 & pi970;
  assign n34341 = n32270 & n34340;
  assign n34342 = n64082 & n34341;
  assign n34343 = n3475 & n34342;
  assign n34344 = ~n34339 & ~n34343;
  assign n34345 = pi57 & ~n34344;
  assign n34346 = pi299 & ~n34339;
  assign n34347 = n2814 & ~n30779;
  assign n34348 = n34340 & n34347;
  assign n34349 = n34346 & ~n34348;
  assign n34350 = ~n30784 & ~n34349;
  assign n34351 = n2814 & n30781;
  assign n34352 = n34340 & n34351;
  assign n34353 = ~n34339 & ~n34352;
  assign n34354 = n30783 & ~n34353;
  assign n34355 = ~n34350 & ~n34354;
  assign n34356 = n2814 & ~n34080;
  assign n34357 = ~n30609 & ~n34356;
  assign n34358 = ~pi228 & n30746;
  assign n34359 = ~n30769 & ~n34338;
  assign n34360 = ~n34358 & n34359;
  assign n34361 = ~n34357 & ~n34360;
  assign n34362 = pi967 & n34361;
  assign n34363 = ~pi299 & ~n34362;
  assign n34364 = pi232 & ~n34363;
  assign n34365 = ~n34355 & n34364;
  assign n34366 = pi967 & n34356;
  assign n34367 = ~pi299 & ~n34366;
  assign n34368 = ~pi232 & ~n34349;
  assign n34369 = ~n34367 & n34368;
  assign n34370 = ~n34365 & ~n34369;
  assign n34371 = ~pi39 & ~n34370;
  assign n34372 = pi299 & pi970;
  assign n34373 = n2814 & n30830;
  assign n34374 = ~pi228 & ~n34373;
  assign n34375 = n34372 & ~n34374;
  assign n34376 = ~pi299 & pi967;
  assign n34377 = n2814 & n64103;
  assign n34378 = ~pi228 & ~n34377;
  assign n34379 = n34376 & ~n34378;
  assign n34380 = ~n34375 & ~n34379;
  assign n34381 = pi228 & ~n34337;
  assign n34382 = pi39 & ~n34381;
  assign n34383 = ~n34380 & n34382;
  assign n34384 = ~pi38 & ~n34383;
  assign n34385 = ~n34371 & n34384;
  assign n34386 = ~pi228 & ~n32270;
  assign n34387 = ~n34381 & ~n34386;
  assign n34388 = pi967 & n34387;
  assign n34389 = ~pi299 & ~n34388;
  assign n34390 = ~n34341 & n34346;
  assign n34391 = ~pi39 & ~n34390;
  assign n34392 = ~n34389 & n34391;
  assign n34393 = ~n34372 & ~n34376;
  assign n34394 = n34338 & ~n34393;
  assign n34395 = pi39 & n34394;
  assign n34396 = pi38 & ~n34395;
  assign n34397 = ~n34392 & n34396;
  assign n34398 = ~n34385 & ~n34397;
  assign n34399 = ~pi100 & ~n34398;
  assign n34400 = n2814 & n34139;
  assign n34401 = n30858 & n34400;
  assign n34402 = ~n30858 & n34142;
  assign n34403 = ~pi228 & ~n34402;
  assign n34404 = ~pi228 & ~n34401;
  assign n34405 = ~n34402 & n34404;
  assign n34406 = ~n34401 & n34403;
  assign n34407 = ~n34381 & ~n64313;
  assign n34408 = pi967 & n34407;
  assign n34409 = ~pi299 & ~n34408;
  assign n34410 = n30860 & ~n34400;
  assign n34411 = ~n30860 & ~n34142;
  assign n34412 = ~pi228 & ~n34411;
  assign n34413 = ~pi228 & ~n34410;
  assign n34414 = ~n34411 & n34413;
  assign n34415 = ~n34410 & n34412;
  assign n34416 = pi970 & n64314;
  assign n34417 = n34346 & ~n34416;
  assign n34418 = n2764 & ~n34417;
  assign n34419 = ~n34409 & n34418;
  assign n34420 = ~n2764 & n34394;
  assign n34421 = pi100 & ~n34420;
  assign n34422 = ~n34419 & n34421;
  assign n34423 = ~pi87 & ~n34422;
  assign n34424 = ~n34399 & n34423;
  assign n34425 = pi87 & n34394;
  assign n34426 = ~pi75 & ~n34425;
  assign n34427 = ~n34424 & n34426;
  assign n34428 = ~n2806 & n34394;
  assign n34429 = n62951 & n34392;
  assign n34430 = ~n34428 & ~n34429;
  assign n34431 = pi75 & n34430;
  assign n34432 = ~pi92 & ~n34431;
  assign n34433 = ~n34427 & n34432;
  assign n34434 = ~pi75 & n34430;
  assign n34435 = pi75 & ~n34394;
  assign n34436 = pi92 & ~n34435;
  assign n34437 = ~n34434 & n34436;
  assign n34438 = ~pi54 & ~n34437;
  assign n34439 = ~n34433 & n34438;
  assign n34440 = n6793 & n34430;
  assign n34441 = ~n6793 & ~n34394;
  assign n34442 = ~n34440 & ~n34441;
  assign n34443 = pi54 & ~n34442;
  assign n34444 = ~pi74 & ~n34443;
  assign n34445 = ~n34439 & n34444;
  assign n34446 = ~pi54 & n34440;
  assign n34447 = ~n34066 & ~n34394;
  assign n34448 = pi74 & ~n34447;
  assign n34449 = ~n34446 & n34448;
  assign n34450 = ~pi55 & ~n34449;
  assign n34451 = ~n34445 & n34450;
  assign n34452 = pi55 & ~n34339;
  assign n34453 = ~n34342 & n34452;
  assign n34454 = n3470 & ~n34453;
  assign n34455 = ~n34451 & n34454;
  assign n34456 = ~n3470 & n34339;
  assign n34457 = ~pi59 & ~n34456;
  assign n34458 = ~n34455 & n34457;
  assign n34459 = n3471 & n34342;
  assign n34460 = pi59 & ~n34339;
  assign n34461 = ~n34459 & n34460;
  assign n34462 = ~pi57 & ~n34461;
  assign n34463 = ~n34458 & n34462;
  assign po173 = ~n34345 & ~n34463;
  assign n34465 = pi972 & n34338;
  assign n34466 = ~pi228 & pi972;
  assign n34467 = n32270 & n34466;
  assign n34468 = n64082 & n34467;
  assign n34469 = n3475 & n34468;
  assign n34470 = ~n34465 & ~n34469;
  assign n34471 = pi57 & ~n34470;
  assign n34472 = pi299 & ~n34465;
  assign n34473 = n34347 & n34466;
  assign n34474 = n34472 & ~n34473;
  assign n34475 = ~n30784 & ~n34474;
  assign n34476 = n34351 & n34466;
  assign n34477 = ~n34465 & ~n34476;
  assign n34478 = n30783 & ~n34477;
  assign n34479 = ~n34475 & ~n34478;
  assign n34480 = pi961 & n34361;
  assign n34481 = ~pi299 & ~n34480;
  assign n34482 = pi232 & ~n34481;
  assign n34483 = ~n34479 & n34482;
  assign n34484 = pi961 & n34356;
  assign n34485 = ~pi299 & ~n34484;
  assign n34486 = ~pi232 & ~n34474;
  assign n34487 = ~n34485 & n34486;
  assign n34488 = ~n34483 & ~n34487;
  assign n34489 = ~pi39 & ~n34488;
  assign n34490 = ~pi299 & pi961;
  assign n34491 = ~n34378 & n34490;
  assign n34492 = pi299 & pi972;
  assign n34493 = ~n34374 & n34492;
  assign n34494 = ~n34491 & ~n34493;
  assign n34495 = n34382 & ~n34494;
  assign n34496 = ~pi38 & ~n34495;
  assign n34497 = ~n34489 & n34496;
  assign n34498 = pi961 & n34387;
  assign n34499 = ~pi299 & ~n34498;
  assign n34500 = ~n34467 & n34472;
  assign n34501 = ~pi39 & ~n34500;
  assign n34502 = ~n34499 & n34501;
  assign n34503 = ~n34490 & ~n34492;
  assign n34504 = n34338 & ~n34503;
  assign n34505 = pi39 & n34504;
  assign n34506 = pi38 & ~n34505;
  assign n34507 = ~n34502 & n34506;
  assign n34508 = ~n34497 & ~n34507;
  assign n34509 = ~pi100 & ~n34508;
  assign n34510 = pi961 & n34407;
  assign n34511 = ~pi299 & ~n34510;
  assign n34512 = pi972 & n64314;
  assign n34513 = n34472 & ~n34512;
  assign n34514 = n2764 & ~n34513;
  assign n34515 = ~n34511 & n34514;
  assign n34516 = ~n2764 & n34504;
  assign n34517 = pi100 & ~n34516;
  assign n34518 = ~n34515 & n34517;
  assign n34519 = ~pi87 & ~n34518;
  assign n34520 = ~n34509 & n34519;
  assign n34521 = pi87 & n34504;
  assign n34522 = ~pi75 & ~n34521;
  assign n34523 = ~n34520 & n34522;
  assign n34524 = ~n2806 & n34504;
  assign n34525 = n62951 & n34502;
  assign n34526 = ~n34524 & ~n34525;
  assign n34527 = pi75 & n34526;
  assign n34528 = ~pi92 & ~n34527;
  assign n34529 = ~n34523 & n34528;
  assign n34530 = ~pi75 & n34526;
  assign n34531 = pi75 & ~n34504;
  assign n34532 = pi92 & ~n34531;
  assign n34533 = ~n34530 & n34532;
  assign n34534 = ~pi54 & ~n34533;
  assign n34535 = ~n34529 & n34534;
  assign n34536 = n6793 & n34526;
  assign n34537 = ~n6793 & ~n34504;
  assign n34538 = ~n34536 & ~n34537;
  assign n34539 = pi54 & ~n34538;
  assign n34540 = ~pi74 & ~n34539;
  assign n34541 = ~n34535 & n34540;
  assign n34542 = ~pi54 & n34536;
  assign n34543 = ~n34066 & ~n34504;
  assign n34544 = pi74 & ~n34543;
  assign n34545 = ~n34542 & n34544;
  assign n34546 = ~pi55 & ~n34545;
  assign n34547 = ~n34541 & n34546;
  assign n34548 = pi55 & ~n34465;
  assign n34549 = ~n34468 & n34548;
  assign n34550 = n3470 & ~n34549;
  assign n34551 = ~n34547 & n34550;
  assign n34552 = ~n3470 & n34465;
  assign n34553 = ~pi59 & ~n34552;
  assign n34554 = ~n34551 & n34553;
  assign n34555 = n3471 & n34468;
  assign n34556 = pi59 & ~n34465;
  assign n34557 = ~n34555 & n34556;
  assign n34558 = ~pi57 & ~n34557;
  assign n34559 = ~n34554 & n34558;
  assign po174 = ~n34471 & ~n34559;
  assign n34561 = pi960 & n34338;
  assign n34562 = ~pi228 & pi960;
  assign n34563 = n32270 & n34562;
  assign n34564 = n64082 & n34563;
  assign n34565 = n3475 & n34564;
  assign n34566 = ~n34561 & ~n34565;
  assign n34567 = pi57 & ~n34566;
  assign n34568 = pi299 & ~n34561;
  assign n34569 = n34347 & n34562;
  assign n34570 = n34568 & ~n34569;
  assign n34571 = ~n30784 & ~n34570;
  assign n34572 = n34351 & n34562;
  assign n34573 = ~n34561 & ~n34572;
  assign n34574 = n30783 & ~n34573;
  assign n34575 = ~n34571 & ~n34574;
  assign n34576 = pi977 & n34361;
  assign n34577 = ~pi299 & ~n34576;
  assign n34578 = pi232 & ~n34577;
  assign n34579 = ~n34575 & n34578;
  assign n34580 = pi977 & n34356;
  assign n34581 = ~pi299 & ~n34580;
  assign n34582 = ~pi232 & ~n34570;
  assign n34583 = ~n34581 & n34582;
  assign n34584 = ~n34579 & ~n34583;
  assign n34585 = ~pi39 & ~n34584;
  assign n34586 = ~pi299 & pi977;
  assign n34587 = ~n34378 & n34586;
  assign n34588 = pi299 & pi960;
  assign n34589 = ~n34374 & n34588;
  assign n34590 = ~n34587 & ~n34589;
  assign n34591 = n34382 & ~n34590;
  assign n34592 = ~pi38 & ~n34591;
  assign n34593 = ~n34585 & n34592;
  assign n34594 = pi977 & n34387;
  assign n34595 = ~pi299 & ~n34594;
  assign n34596 = ~n34563 & n34568;
  assign n34597 = ~pi39 & ~n34596;
  assign n34598 = ~n34595 & n34597;
  assign n34599 = ~n34586 & ~n34588;
  assign n34600 = n34338 & ~n34599;
  assign n34601 = pi39 & n34600;
  assign n34602 = pi38 & ~n34601;
  assign n34603 = ~n34598 & n34602;
  assign n34604 = ~n34593 & ~n34603;
  assign n34605 = ~pi100 & ~n34604;
  assign n34606 = pi977 & n34407;
  assign n34607 = ~pi299 & ~n34606;
  assign n34608 = pi960 & n64314;
  assign n34609 = n34568 & ~n34608;
  assign n34610 = n2764 & ~n34609;
  assign n34611 = ~n34607 & n34610;
  assign n34612 = ~n2764 & n34600;
  assign n34613 = pi100 & ~n34612;
  assign n34614 = ~n34611 & n34613;
  assign n34615 = ~pi87 & ~n34614;
  assign n34616 = ~n34605 & n34615;
  assign n34617 = pi87 & n34600;
  assign n34618 = ~pi75 & ~n34617;
  assign n34619 = ~n34616 & n34618;
  assign n34620 = ~n2806 & n34600;
  assign n34621 = n62951 & n34598;
  assign n34622 = ~n34620 & ~n34621;
  assign n34623 = pi75 & n34622;
  assign n34624 = ~pi92 & ~n34623;
  assign n34625 = ~n34619 & n34624;
  assign n34626 = ~pi75 & n34622;
  assign n34627 = pi75 & ~n34600;
  assign n34628 = pi92 & ~n34627;
  assign n34629 = ~n34626 & n34628;
  assign n34630 = ~pi54 & ~n34629;
  assign n34631 = ~n34625 & n34630;
  assign n34632 = n6793 & n34622;
  assign n34633 = ~n6793 & ~n34600;
  assign n34634 = ~n34632 & ~n34633;
  assign n34635 = pi54 & ~n34634;
  assign n34636 = ~pi74 & ~n34635;
  assign n34637 = ~n34631 & n34636;
  assign n34638 = ~pi54 & n34632;
  assign n34639 = ~n34066 & ~n34600;
  assign n34640 = pi74 & ~n34639;
  assign n34641 = ~n34638 & n34640;
  assign n34642 = ~pi55 & ~n34641;
  assign n34643 = ~n34637 & n34642;
  assign n34644 = pi55 & ~n34561;
  assign n34645 = ~n34564 & n34644;
  assign n34646 = n3470 & ~n34645;
  assign n34647 = ~n34643 & n34646;
  assign n34648 = ~n3470 & n34561;
  assign n34649 = ~pi59 & ~n34648;
  assign n34650 = ~n34647 & n34649;
  assign n34651 = n3471 & n34564;
  assign n34652 = pi59 & ~n34561;
  assign n34653 = ~n34651 & n34652;
  assign n34654 = ~pi57 & ~n34653;
  assign n34655 = ~n34650 & n34654;
  assign po175 = ~n34567 & ~n34655;
  assign n34657 = pi963 & n34338;
  assign n34658 = ~pi228 & pi963;
  assign n34659 = n32270 & n34658;
  assign n34660 = n64082 & n34659;
  assign n34661 = n3475 & n34660;
  assign n34662 = ~n34657 & ~n34661;
  assign n34663 = pi57 & ~n34662;
  assign n34664 = pi299 & ~n34657;
  assign n34665 = n34347 & n34658;
  assign n34666 = n34664 & ~n34665;
  assign n34667 = ~n30784 & ~n34666;
  assign n34668 = n34351 & n34658;
  assign n34669 = ~n34657 & ~n34668;
  assign n34670 = n30783 & ~n34669;
  assign n34671 = ~n34667 & ~n34670;
  assign n34672 = pi969 & n34361;
  assign n34673 = ~pi299 & ~n34672;
  assign n34674 = pi232 & ~n34673;
  assign n34675 = ~n34671 & n34674;
  assign n34676 = pi969 & n34356;
  assign n34677 = ~pi299 & ~n34676;
  assign n34678 = ~pi232 & ~n34666;
  assign n34679 = ~n34677 & n34678;
  assign n34680 = ~n34675 & ~n34679;
  assign n34681 = ~pi39 & ~n34680;
  assign n34682 = ~pi299 & pi969;
  assign n34683 = ~n34378 & n34682;
  assign n34684 = pi299 & pi963;
  assign n34685 = ~n34374 & n34684;
  assign n34686 = ~n34683 & ~n34685;
  assign n34687 = n34382 & ~n34686;
  assign n34688 = ~pi38 & ~n34687;
  assign n34689 = ~n34681 & n34688;
  assign n34690 = pi969 & n34387;
  assign n34691 = ~pi299 & ~n34690;
  assign n34692 = ~n34659 & n34664;
  assign n34693 = ~pi39 & ~n34692;
  assign n34694 = ~n34691 & n34693;
  assign n34695 = ~n34682 & ~n34684;
  assign n34696 = n34338 & ~n34695;
  assign n34697 = pi39 & n34696;
  assign n34698 = pi38 & ~n34697;
  assign n34699 = ~n34694 & n34698;
  assign n34700 = ~n34689 & ~n34699;
  assign n34701 = ~pi100 & ~n34700;
  assign n34702 = pi969 & n34407;
  assign n34703 = ~pi299 & ~n34702;
  assign n34704 = pi963 & n64314;
  assign n34705 = n34664 & ~n34704;
  assign n34706 = n2764 & ~n34705;
  assign n34707 = ~n34703 & n34706;
  assign n34708 = ~n2764 & n34696;
  assign n34709 = pi100 & ~n34708;
  assign n34710 = ~n34707 & n34709;
  assign n34711 = ~pi87 & ~n34710;
  assign n34712 = ~n34701 & n34711;
  assign n34713 = pi87 & n34696;
  assign n34714 = ~pi75 & ~n34713;
  assign n34715 = ~n34712 & n34714;
  assign n34716 = ~n2806 & n34696;
  assign n34717 = n62951 & n34694;
  assign n34718 = ~n34716 & ~n34717;
  assign n34719 = pi75 & n34718;
  assign n34720 = ~pi92 & ~n34719;
  assign n34721 = ~n34715 & n34720;
  assign n34722 = ~pi75 & n34718;
  assign n34723 = pi75 & ~n34696;
  assign n34724 = pi92 & ~n34723;
  assign n34725 = ~n34722 & n34724;
  assign n34726 = ~pi54 & ~n34725;
  assign n34727 = ~n34721 & n34726;
  assign n34728 = n6793 & n34718;
  assign n34729 = ~n6793 & ~n34696;
  assign n34730 = ~n34728 & ~n34729;
  assign n34731 = pi54 & ~n34730;
  assign n34732 = ~pi74 & ~n34731;
  assign n34733 = ~n34727 & n34732;
  assign n34734 = ~pi54 & n34728;
  assign n34735 = ~n34066 & ~n34696;
  assign n34736 = pi74 & ~n34735;
  assign n34737 = ~n34734 & n34736;
  assign n34738 = ~pi55 & ~n34737;
  assign n34739 = ~n34733 & n34738;
  assign n34740 = pi55 & ~n34657;
  assign n34741 = ~n34660 & n34740;
  assign n34742 = n3470 & ~n34741;
  assign n34743 = ~n34739 & n34742;
  assign n34744 = ~n3470 & n34657;
  assign n34745 = ~pi59 & ~n34744;
  assign n34746 = ~n34743 & n34745;
  assign n34747 = n3471 & n34660;
  assign n34748 = pi59 & ~n34657;
  assign n34749 = ~n34747 & n34748;
  assign n34750 = ~pi57 & ~n34749;
  assign n34751 = ~n34746 & n34750;
  assign po176 = ~n34663 & ~n34751;
  assign n34753 = pi975 & n34338;
  assign n34754 = ~pi228 & pi975;
  assign n34755 = n32270 & n34754;
  assign n34756 = n64082 & n34755;
  assign n34757 = n3475 & n34756;
  assign n34758 = ~n34753 & ~n34757;
  assign n34759 = pi57 & ~n34758;
  assign n34760 = pi299 & ~n34753;
  assign n34761 = n34347 & n34754;
  assign n34762 = n34760 & ~n34761;
  assign n34763 = ~n30784 & ~n34762;
  assign n34764 = n34351 & n34754;
  assign n34765 = ~n34753 & ~n34764;
  assign n34766 = n30783 & ~n34765;
  assign n34767 = ~n34763 & ~n34766;
  assign n34768 = pi971 & n34361;
  assign n34769 = ~pi299 & ~n34768;
  assign n34770 = pi232 & ~n34769;
  assign n34771 = ~n34767 & n34770;
  assign n34772 = pi971 & n34356;
  assign n34773 = ~pi299 & ~n34772;
  assign n34774 = ~pi232 & ~n34762;
  assign n34775 = ~n34773 & n34774;
  assign n34776 = ~n34771 & ~n34775;
  assign n34777 = ~pi39 & ~n34776;
  assign n34778 = ~pi299 & pi971;
  assign n34779 = ~n34378 & n34778;
  assign n34780 = pi299 & pi975;
  assign n34781 = ~n34374 & n34780;
  assign n34782 = ~n34779 & ~n34781;
  assign n34783 = n34382 & ~n34782;
  assign n34784 = ~pi38 & ~n34783;
  assign n34785 = ~n34777 & n34784;
  assign n34786 = pi971 & n34387;
  assign n34787 = ~pi299 & ~n34786;
  assign n34788 = ~n34755 & n34760;
  assign n34789 = ~pi39 & ~n34788;
  assign n34790 = ~n34787 & n34789;
  assign n34791 = ~n34778 & ~n34780;
  assign n34792 = n34338 & ~n34791;
  assign n34793 = pi39 & n34792;
  assign n34794 = pi38 & ~n34793;
  assign n34795 = ~n34790 & n34794;
  assign n34796 = ~n34785 & ~n34795;
  assign n34797 = ~pi100 & ~n34796;
  assign n34798 = pi971 & n34407;
  assign n34799 = ~pi299 & ~n34798;
  assign n34800 = pi975 & n64314;
  assign n34801 = n34760 & ~n34800;
  assign n34802 = n2764 & ~n34801;
  assign n34803 = ~n34799 & n34802;
  assign n34804 = ~n2764 & n34792;
  assign n34805 = pi100 & ~n34804;
  assign n34806 = ~n34803 & n34805;
  assign n34807 = ~pi87 & ~n34806;
  assign n34808 = ~n34797 & n34807;
  assign n34809 = pi87 & n34792;
  assign n34810 = ~pi75 & ~n34809;
  assign n34811 = ~n34808 & n34810;
  assign n34812 = ~n2806 & n34792;
  assign n34813 = n62951 & n34790;
  assign n34814 = ~n34812 & ~n34813;
  assign n34815 = pi75 & n34814;
  assign n34816 = ~pi92 & ~n34815;
  assign n34817 = ~n34811 & n34816;
  assign n34818 = ~pi75 & n34814;
  assign n34819 = pi75 & ~n34792;
  assign n34820 = pi92 & ~n34819;
  assign n34821 = ~n34818 & n34820;
  assign n34822 = ~pi54 & ~n34821;
  assign n34823 = ~n34817 & n34822;
  assign n34824 = n6793 & n34814;
  assign n34825 = ~n6793 & ~n34792;
  assign n34826 = ~n34824 & ~n34825;
  assign n34827 = pi54 & ~n34826;
  assign n34828 = ~pi74 & ~n34827;
  assign n34829 = ~n34823 & n34828;
  assign n34830 = ~pi54 & n34824;
  assign n34831 = ~n34066 & ~n34792;
  assign n34832 = pi74 & ~n34831;
  assign n34833 = ~n34830 & n34832;
  assign n34834 = ~pi55 & ~n34833;
  assign n34835 = ~n34829 & n34834;
  assign n34836 = pi55 & ~n34753;
  assign n34837 = ~n34756 & n34836;
  assign n34838 = n3470 & ~n34837;
  assign n34839 = ~n34835 & n34838;
  assign n34840 = ~n3470 & n34753;
  assign n34841 = ~pi59 & ~n34840;
  assign n34842 = ~n34839 & n34841;
  assign n34843 = n3471 & n34756;
  assign n34844 = pi59 & ~n34753;
  assign n34845 = ~n34843 & n34844;
  assign n34846 = ~pi57 & ~n34845;
  assign n34847 = ~n34842 & n34846;
  assign po177 = ~n34759 & ~n34847;
  assign n34849 = pi978 & n34338;
  assign n34850 = ~pi228 & pi978;
  assign n34851 = n64082 & n34850;
  assign n34852 = n32270 & n34851;
  assign n34853 = n3475 & n34852;
  assign n34854 = ~n34849 & ~n34853;
  assign n34855 = pi57 & ~n34854;
  assign n34856 = ~pi299 & pi974;
  assign n34857 = pi299 & pi978;
  assign n34858 = ~n34856 & ~n34857;
  assign n34859 = n34387 & ~n34858;
  assign n34860 = ~pi39 & n34859;
  assign n34861 = n34338 & ~n34858;
  assign n34862 = pi39 & n34861;
  assign n34863 = pi38 & ~n34862;
  assign n34864 = ~n34860 & n34863;
  assign n34865 = pi299 & ~n34849;
  assign n34866 = n34347 & n34850;
  assign n34867 = n34865 & ~n34866;
  assign n34868 = ~n30784 & ~n34867;
  assign n34869 = n34351 & n34850;
  assign n34870 = ~n34849 & ~n34869;
  assign n34871 = n30783 & ~n34870;
  assign n34872 = ~n34868 & ~n34871;
  assign n34873 = pi974 & n34361;
  assign n34874 = ~pi299 & ~n34873;
  assign n34875 = pi232 & ~n34874;
  assign n34876 = ~n34872 & n34875;
  assign n34877 = pi974 & n34356;
  assign n34878 = ~pi299 & ~n34877;
  assign n34879 = ~pi232 & ~n34867;
  assign n34880 = ~n34878 & n34879;
  assign n34881 = ~n34876 & ~n34880;
  assign n34882 = ~pi39 & ~n34881;
  assign n34883 = ~n34378 & n34856;
  assign n34884 = ~n34374 & n34857;
  assign n34885 = ~n34883 & ~n34884;
  assign n34886 = n34382 & ~n34885;
  assign n34887 = ~pi38 & ~n34886;
  assign n34888 = ~n34882 & n34887;
  assign n34889 = ~n34864 & ~n34888;
  assign n34890 = ~pi100 & ~n34889;
  assign n34891 = pi974 & n34407;
  assign n34892 = ~pi299 & ~n34891;
  assign n34893 = pi978 & n64314;
  assign n34894 = n34865 & ~n34893;
  assign n34895 = n2764 & ~n34894;
  assign n34896 = ~n34892 & n34895;
  assign n34897 = ~n2764 & n34861;
  assign n34898 = pi100 & ~n34897;
  assign n34899 = ~n34896 & n34898;
  assign n34900 = ~pi87 & ~n34899;
  assign n34901 = ~n34890 & n34900;
  assign n34902 = pi87 & n34861;
  assign n34903 = ~pi75 & ~n34902;
  assign n34904 = ~n34901 & n34903;
  assign n34905 = ~pi228 & ~n2806;
  assign n34906 = n34859 & ~n34905;
  assign n34907 = pi75 & ~n34906;
  assign n34908 = ~pi92 & ~n34907;
  assign n34909 = ~n34904 & n34908;
  assign n34910 = ~pi75 & ~n34906;
  assign n34911 = pi75 & ~n34861;
  assign n34912 = pi92 & ~n34911;
  assign n34913 = ~n34910 & n34912;
  assign n34914 = ~pi54 & ~n34913;
  assign n34915 = ~n34909 & n34914;
  assign n34916 = n6793 & ~n34906;
  assign n34917 = ~n6793 & ~n34861;
  assign n34918 = ~n34916 & ~n34917;
  assign n34919 = pi54 & ~n34918;
  assign n34920 = ~pi74 & ~n34919;
  assign n34921 = ~n34915 & n34920;
  assign n34922 = ~pi54 & n34916;
  assign n34923 = ~n34066 & ~n34861;
  assign n34924 = pi74 & ~n34923;
  assign n34925 = ~n34922 & n34924;
  assign n34926 = ~pi55 & ~n34925;
  assign n34927 = ~n34921 & n34926;
  assign n34928 = pi55 & ~n34849;
  assign n34929 = ~n34852 & n34928;
  assign n34930 = n3470 & ~n34929;
  assign n34931 = ~n34927 & n34930;
  assign n34932 = ~n3470 & n34849;
  assign n34933 = ~pi59 & ~n34932;
  assign n34934 = ~n34931 & n34933;
  assign n34935 = n3471 & n34852;
  assign n34936 = pi59 & ~n34849;
  assign n34937 = ~n34935 & n34936;
  assign n34938 = ~pi57 & ~n34937;
  assign n34939 = ~n34934 & n34938;
  assign po178 = ~n34855 & ~n34939;
  assign n34941 = ~pi110 & n31891;
  assign n34942 = ~n2920 & n34941;
  assign n34943 = ~n2920 & n2960;
  assign n34944 = n2960 & n34942;
  assign n34945 = n34941 & n34943;
  assign n34946 = pi299 & n64315;
  assign n34947 = n2961 & n34942;
  assign n34948 = n64102 & n34941;
  assign n34949 = pi39 & ~n34948;
  assign n34950 = ~n64316 & n34949;
  assign n34951 = n2664 & n33928;
  assign n34952 = pi72 & n64089;
  assign n34953 = n34951 & n34952;
  assign n34954 = ~pi50 & n62356;
  assign n34955 = n30707 & n34954;
  assign n34956 = ~pi111 & ~n30684;
  assign n34957 = ~pi36 & n33882;
  assign n34958 = ~n34956 & n34957;
  assign n34959 = n2606 & ~n34958;
  assign n34960 = ~n30646 & ~n33887;
  assign n34961 = ~n34959 & n34960;
  assign n34962 = ~pi83 & ~n34961;
  assign n34963 = n30648 & ~n34962;
  assign n34964 = ~pi71 & ~n34963;
  assign n34965 = n30696 & ~n34964;
  assign n34966 = ~pi81 & ~n34965;
  assign n34967 = n34955 & ~n34966;
  assign n34968 = ~pi90 & ~n34967;
  assign n34969 = n62770 & ~n34968;
  assign n34970 = pi90 & ~n34951;
  assign n34971 = n6832 & ~n34970;
  assign n34972 = n34969 & n34971;
  assign n34973 = ~n34953 & ~n34972;
  assign n34974 = ~n2816 & ~n2843;
  assign n34975 = n2852 & ~n6899;
  assign n34976 = n34974 & n34975;
  assign n34977 = n2751 & n34976;
  assign n34978 = ~n34973 & n34977;
  assign n34979 = ~pi93 & ~n30627;
  assign n34980 = n34969 & n34979;
  assign n34981 = ~pi72 & ~n34980;
  assign n34982 = n30619 & ~n34976;
  assign n34983 = ~n34981 & n34982;
  assign n34984 = ~n34978 & ~n34983;
  assign n34985 = n62952 & ~n34984;
  assign n34986 = pi110 & n34976;
  assign n34987 = ~pi39 & ~n34986;
  assign n34988 = ~n34985 & n34987;
  assign n34989 = ~n34950 & ~n34988;
  assign n34990 = n62455 & ~n34989;
  assign n34991 = pi39 & n2960;
  assign n34992 = n34942 & n34991;
  assign n34993 = n2811 & n2815;
  assign n34994 = ~pi39 & pi110;
  assign n34995 = n34975 & n34994;
  assign n34996 = ~n34993 & n34995;
  assign n34997 = ~n2843 & n34996;
  assign n34998 = ~n62455 & ~n34997;
  assign n34999 = ~n34992 & n34998;
  assign n35000 = pi39 & ~n64315;
  assign n35001 = pi110 & n34975;
  assign n35002 = ~n34993 & n35001;
  assign n35003 = ~n2843 & n35002;
  assign n35004 = ~pi39 & ~n35003;
  assign n35005 = ~n62455 & ~n35004;
  assign n35006 = ~n34992 & ~n34997;
  assign n35007 = ~n62455 & ~n35006;
  assign n35008 = ~n35000 & n35005;
  assign n35009 = n2751 & ~n34973;
  assign n35010 = ~pi110 & ~n35009;
  assign n35011 = n34976 & ~n35010;
  assign n35012 = ~pi39 & ~n34983;
  assign n35013 = ~n35011 & n35012;
  assign n35014 = ~n34950 & ~n35013;
  assign n35015 = n62952 & ~n35014;
  assign n35016 = ~n34950 & ~n34987;
  assign n35017 = ~n62952 & ~n35016;
  assign n35018 = n62455 & ~n35017;
  assign n35019 = ~n35015 & n35018;
  assign n35020 = ~n64317 & ~n35019;
  assign n35021 = ~n34990 & ~n34999;
  assign n35022 = n2765 & n32048;
  assign n35023 = n31387 & ~n64176;
  assign n35024 = pi92 & ~n64319;
  assign n35025 = n6792 & ~n35024;
  assign n35026 = ~pi75 & ~n33587;
  assign n35027 = pi299 & ~n31842;
  assign n35028 = ~pi299 & ~n31702;
  assign n35029 = ~pi232 & ~n35028;
  assign n35030 = ~pi232 & ~n35027;
  assign n35031 = ~n35028 & n35030;
  assign n35032 = ~n35027 & n35029;
  assign n35033 = ~pi39 & ~n64320;
  assign n35034 = pi148 & n2814;
  assign n35035 = ~n31842 & ~n35034;
  assign n35036 = pi148 & n33003;
  assign n35037 = ~n35035 & ~n35036;
  assign n35038 = pi299 & ~n35037;
  assign n35039 = ~n2814 & ~n31702;
  assign n35040 = ~n33028 & ~n35039;
  assign n35041 = ~pi299 & ~n35040;
  assign n35042 = pi141 & n35041;
  assign n35043 = n31411 & ~n35040;
  assign n35044 = ~pi141 & n35028;
  assign n35045 = pi232 & ~n35044;
  assign n35046 = ~n64321 & n35045;
  assign n35047 = ~n35038 & n35045;
  assign n35048 = ~n64321 & n35047;
  assign n35049 = ~n35038 & n35046;
  assign n35050 = n35033 & ~n64322;
  assign n35051 = ~n31902 & ~n32692;
  assign n35052 = n31938 & ~n35051;
  assign n35053 = n33108 & ~n35052;
  assign n35054 = ~n62393 & ~n31902;
  assign n35055 = n31886 & ~n35051;
  assign n35056 = ~n35054 & n35055;
  assign n35057 = n31908 & ~n35056;
  assign n35058 = ~n35053 & ~n35057;
  assign n35059 = ~pi232 & ~n35058;
  assign n35060 = ~n31898 & ~n35051;
  assign n35061 = ~n31907 & ~n35060;
  assign n35062 = pi148 & ~n35061;
  assign n35063 = ~n31412 & ~n35057;
  assign n35064 = ~n35062 & ~n35063;
  assign n35065 = pi141 & n31929;
  assign n35066 = n35052 & ~n35065;
  assign n35067 = ~pi141 & n35053;
  assign n35068 = ~n31929 & n35052;
  assign n35069 = n33108 & ~n35068;
  assign n35070 = pi141 & n35069;
  assign n35071 = ~n35067 & ~n35070;
  assign n35072 = n33108 & ~n35066;
  assign n35073 = ~n35064 & n64323;
  assign n35074 = pi232 & ~n35073;
  assign n35075 = ~n35059 & ~n35074;
  assign n35076 = pi39 & ~n35075;
  assign n35077 = n2766 & ~n35076;
  assign n35078 = ~n35050 & n35077;
  assign n35079 = ~pi87 & ~n35078;
  assign n35080 = n35026 & ~n35079;
  assign n35081 = ~pi92 & ~n35080;
  assign n35082 = n35025 & ~n35081;
  assign n35083 = ~pi55 & ~n35082;
  assign n35084 = n31388 & ~n33149;
  assign n35085 = pi55 & ~n35084;
  assign n35086 = ~n35083 & ~n35085;
  assign n35087 = n3470 & ~n35086;
  assign n35088 = n31390 & ~n35087;
  assign n35089 = pi138 & n35088;
  assign n35090 = ~n2909 & n31412;
  assign n35091 = n2909 & n30824;
  assign n35092 = n31926 & n35091;
  assign n35093 = n31411 & ~n35092;
  assign n35094 = ~n35090 & ~n35093;
  assign n35095 = pi232 & ~n35094;
  assign n35096 = ~n2973 & n30824;
  assign n35097 = n31926 & n35096;
  assign n35098 = ~pi299 & ~n35097;
  assign n35099 = ~n2920 & n30824;
  assign n35100 = n31886 & n35099;
  assign n35101 = pi299 & ~n35100;
  assign n35102 = ~n35098 & ~n35101;
  assign n35103 = pi232 & ~pi299;
  assign n35104 = pi141 & n35103;
  assign n35105 = ~n35102 & ~n35104;
  assign n35106 = ~pi232 & ~n35102;
  assign n35107 = ~n31411 & ~n35102;
  assign n35108 = n35094 & ~n35107;
  assign n35109 = pi232 & ~n35108;
  assign n35110 = ~n35106 & ~n35109;
  assign n35111 = ~n35095 & ~n35105;
  assign n35112 = pi39 & ~n64324;
  assign n35113 = n62455 & n6792;
  assign n35114 = ~pi38 & n63888;
  assign n35115 = n9738 & n35113;
  assign n35116 = ~n31414 & n64197;
  assign n35117 = ~pi39 & ~n35116;
  assign n35118 = n64325 & ~n35117;
  assign n35119 = ~n35112 & n35118;
  assign n35120 = ~pi138 & n35119;
  assign n35121 = ~pi118 & n33162;
  assign n35122 = ~pi139 & n35121;
  assign n35123 = ~n35120 & ~n35122;
  assign n35124 = ~n35089 & n35123;
  assign n35125 = ~pi138 & ~n32292;
  assign n35126 = n35088 & n35125;
  assign n35127 = n35119 & ~n35125;
  assign n35128 = n35122 & ~n35127;
  assign n35129 = ~n35126 & n35128;
  assign po295 = ~n35124 & ~n35129;
  assign n35131 = pi169 & n2814;
  assign n35132 = ~n31842 & ~n35131;
  assign n35133 = pi169 & n33003;
  assign n35134 = ~n35132 & ~n35133;
  assign n35135 = pi299 & ~n35134;
  assign n35136 = pi191 & n35041;
  assign n35137 = n33355 & ~n35040;
  assign n35138 = ~pi191 & n35028;
  assign n35139 = pi232 & ~n35138;
  assign n35140 = ~n64326 & n35139;
  assign n35141 = ~n35135 & n35139;
  assign n35142 = ~n64326 & n35141;
  assign n35143 = ~n35135 & n35140;
  assign n35144 = n35033 & ~n64327;
  assign n35145 = ~pi169 & n31902;
  assign n35146 = ~n35060 & ~n35145;
  assign n35147 = n31886 & ~n35146;
  assign n35148 = n31908 & ~n35147;
  assign n35149 = pi191 & n35069;
  assign n35150 = ~n35148 & ~n35149;
  assign n35151 = pi232 & ~n35150;
  assign n35152 = ~pi191 & n35053;
  assign n35153 = ~n35059 & ~n35152;
  assign n35154 = ~n35149 & ~n35152;
  assign n35155 = ~n35148 & ~n35152;
  assign n35156 = ~n35149 & n35155;
  assign n35157 = ~n35148 & n35154;
  assign n35158 = pi232 & ~n64328;
  assign n35159 = ~n35059 & ~n35158;
  assign n35160 = ~n35151 & n35153;
  assign n35161 = pi39 & ~n64329;
  assign n35162 = n2766 & ~n35161;
  assign n35163 = ~n35144 & n35162;
  assign n35164 = ~pi87 & ~n35163;
  assign n35165 = n35026 & ~n35164;
  assign n35166 = ~pi92 & ~n35165;
  assign n35167 = n35025 & ~n35166;
  assign n35168 = ~pi55 & ~n35167;
  assign n35169 = ~n35085 & ~n35168;
  assign n35170 = n3470 & ~n35169;
  assign n35171 = n31390 & ~n35170;
  assign n35172 = pi139 & n35171;
  assign n35173 = ~n2909 & n33356;
  assign n35174 = ~n35101 & ~n35173;
  assign n35175 = ~pi191 & ~pi299;
  assign n35176 = ~n35097 & n35175;
  assign n35177 = n33355 & ~n35092;
  assign n35178 = ~n35176 & ~n35177;
  assign n35179 = n35174 & n35178;
  assign n35180 = pi232 & ~n35179;
  assign n35181 = ~n35106 & ~n35180;
  assign n35182 = pi39 & ~n35181;
  assign n35183 = n2815 & ~n33357;
  assign n35184 = n64197 & ~n35183;
  assign n35185 = ~pi39 & ~n35184;
  assign n35186 = n64325 & ~n35185;
  assign n35187 = ~n35182 & n35186;
  assign n35188 = ~pi139 & n35187;
  assign n35189 = ~n35121 & ~n35188;
  assign n35190 = ~n35172 & n35189;
  assign n35191 = ~pi139 & ~n32293;
  assign n35192 = n35171 & n35191;
  assign n35193 = n35187 & ~n35191;
  assign n35194 = n35121 & ~n35193;
  assign n35195 = ~n35192 & n35194;
  assign po296 = ~n35190 & ~n35195;
  assign n35197 = pi171 & pi299;
  assign n35198 = ~n2909 & n35197;
  assign n35199 = ~n35101 & ~n35198;
  assign n35200 = ~pi192 & ~pi299;
  assign n35201 = ~n35097 & n35200;
  assign n35202 = pi192 & ~pi299;
  assign n35203 = ~n35092 & n35202;
  assign n35204 = ~n35201 & ~n35203;
  assign n35205 = n35199 & n35204;
  assign n35206 = pi232 & ~n35205;
  assign n35207 = ~n35106 & ~n35206;
  assign n35208 = pi39 & ~n35207;
  assign n35209 = ~n35197 & ~n35202;
  assign n35210 = n2815 & ~n35209;
  assign n35211 = n64197 & ~n35210;
  assign n35212 = ~pi39 & ~n35211;
  assign n35213 = ~pi138 & n35122;
  assign n35214 = ~pi196 & n35213;
  assign n35215 = pi195 & ~n35214;
  assign n35216 = n64325 & ~n35215;
  assign n35217 = ~n35212 & n35216;
  assign n35218 = ~n35208 & n35217;
  assign n35219 = pi171 & n2814;
  assign n35220 = ~n31842 & ~n35219;
  assign n35221 = pi171 & n33003;
  assign n35222 = ~n35220 & ~n35221;
  assign n35223 = pi299 & ~n35222;
  assign n35224 = pi192 & n35041;
  assign n35225 = ~n35040 & n35202;
  assign n35226 = ~pi192 & n35028;
  assign n35227 = pi232 & ~n35226;
  assign n35228 = ~n64330 & n35227;
  assign n35229 = ~n35223 & n35227;
  assign n35230 = ~n64330 & n35229;
  assign n35231 = ~n35223 & n35228;
  assign n35232 = n35033 & ~n64331;
  assign n35233 = ~pi171 & n31902;
  assign n35234 = ~n35060 & ~n35233;
  assign n35235 = n31886 & ~n35234;
  assign n35236 = n31908 & ~n35235;
  assign n35237 = pi192 & n35069;
  assign n35238 = ~n35236 & ~n35237;
  assign n35239 = pi232 & ~n35238;
  assign n35240 = ~pi192 & n35053;
  assign n35241 = ~n35059 & ~n35240;
  assign n35242 = ~n35237 & ~n35240;
  assign n35243 = ~n35236 & ~n35240;
  assign n35244 = ~n35237 & n35243;
  assign n35245 = ~n35236 & n35242;
  assign n35246 = pi232 & ~n64332;
  assign n35247 = ~n35059 & ~n35246;
  assign n35248 = ~n35239 & n35241;
  assign n35249 = pi39 & ~n64333;
  assign n35250 = n2766 & ~n35249;
  assign n35251 = ~n35232 & n35250;
  assign n35252 = ~pi87 & ~n35251;
  assign n35253 = n35026 & ~n35252;
  assign n35254 = ~pi92 & ~n35253;
  assign n35255 = n35025 & ~n35254;
  assign n35256 = ~pi55 & ~n35255;
  assign n35257 = ~n35085 & ~n35256;
  assign n35258 = n3470 & ~n35257;
  assign n35259 = n31390 & n35215;
  assign n35260 = ~n35258 & n35259;
  assign n35261 = ~n35218 & ~n35260;
  assign n35262 = ~pi170 & n31902;
  assign n35263 = ~n35060 & ~n35262;
  assign n35264 = n31886 & ~n35263;
  assign n35265 = n31908 & ~n35264;
  assign n35266 = ~n35053 & ~n35265;
  assign n35267 = pi232 & ~n35266;
  assign n35268 = ~n35059 & ~n35267;
  assign n35269 = pi39 & ~n35268;
  assign n35270 = ~pi38 & ~pi194;
  assign n35271 = ~n35269 & n35270;
  assign n35272 = n31702 & n35271;
  assign n35273 = pi232 & n35069;
  assign n35274 = n35268 & ~n35273;
  assign n35275 = pi39 & ~n35274;
  assign n35276 = ~pi38 & pi194;
  assign n35277 = ~n35275 & n35276;
  assign n35278 = n35040 & n35277;
  assign n35279 = ~n35272 & ~n35278;
  assign n35280 = n35103 & ~n35279;
  assign n35281 = ~n35271 & ~n35277;
  assign n35282 = pi170 & n33003;
  assign n35283 = pi232 & pi299;
  assign n35284 = pi170 & n2814;
  assign n35285 = ~n31842 & ~n35284;
  assign n35286 = n35283 & ~n35285;
  assign n35287 = ~n35282 & n35286;
  assign n35288 = n35033 & ~n35287;
  assign n35289 = ~n35281 & ~n35288;
  assign n35290 = ~n35033 & ~n35281;
  assign n35291 = ~n35041 & n35277;
  assign n35292 = ~n35028 & n35271;
  assign n35293 = ~n35291 & ~n35292;
  assign n35294 = ~n35282 & ~n35285;
  assign n35295 = pi299 & ~n35294;
  assign n35296 = pi232 & ~n35295;
  assign n35297 = ~n35293 & n35296;
  assign n35298 = ~n35290 & ~n35297;
  assign n35299 = ~n35280 & ~n35289;
  assign n35300 = ~pi100 & ~n64334;
  assign n35301 = ~pi87 & ~n35300;
  assign n35302 = n35026 & ~n35301;
  assign n35303 = ~pi92 & ~n35302;
  assign n35304 = n35025 & ~n35303;
  assign n35305 = ~pi55 & ~n35304;
  assign n35306 = ~n35085 & ~n35305;
  assign n35307 = n3470 & ~n35306;
  assign n35308 = n31390 & ~n35307;
  assign n35309 = pi196 & ~n35308;
  assign n35310 = ~pi170 & n32215;
  assign n35311 = ~n35091 & ~n35310;
  assign n35312 = n64234 & ~n35311;
  assign n35313 = ~pi299 & n35092;
  assign n35314 = n64232 & n35091;
  assign n35315 = pi232 & ~n64335;
  assign n35316 = ~n35312 & n35315;
  assign n35317 = ~n35106 & ~n35316;
  assign n35318 = pi299 & ~n35317;
  assign n35319 = ~n35098 & ~n35318;
  assign n35320 = pi39 & ~n35319;
  assign n35321 = n35283 & n35284;
  assign n35322 = n64197 & ~n35321;
  assign n35323 = ~pi39 & ~n35322;
  assign n35324 = ~pi38 & ~n35323;
  assign n35325 = ~n35320 & n35324;
  assign n35326 = ~pi194 & ~n35325;
  assign n35327 = pi39 & ~n35317;
  assign n35328 = pi170 & n2815;
  assign n35329 = ~n31977 & ~n35328;
  assign n35330 = n64197 & n35329;
  assign n35331 = ~pi39 & ~n35330;
  assign n35332 = ~pi38 & ~n35331;
  assign n35333 = ~n35327 & n35332;
  assign n35334 = pi194 & ~n35333;
  assign n35335 = n63888 & ~n35334;
  assign n35336 = ~n35326 & n35335;
  assign n35337 = ~pi196 & ~n35336;
  assign n35338 = ~n35213 & ~n35337;
  assign n35339 = ~n35309 & n35338;
  assign n35340 = pi195 & ~pi196;
  assign n35341 = ~n35308 & n35340;
  assign n35342 = ~n35336 & ~n35340;
  assign n35343 = n35213 & ~n35342;
  assign n35344 = ~n35341 & n35343;
  assign n35345 = ~n35339 & ~n35344;
  assign n35346 = pi128 & pi228;
  assign n35347 = ~n35113 & n35346;
  assign n35348 = n2979 & ~n7034;
  assign n35349 = n62402 & n35348;
  assign n35350 = n2959 & ~n7118;
  assign n35351 = n62400 & n35350;
  assign n35352 = ~n35349 & ~n35351;
  assign n35353 = pi39 & ~n35352;
  assign n35354 = pi93 & n2659;
  assign n35355 = n2683 & n64093;
  assign n35356 = ~pi86 & ~n35355;
  assign n35357 = ~pi83 & n33888;
  assign n35358 = n2587 & n2611;
  assign n35359 = ~pi65 & n2611;
  assign n35360 = ~pi65 & n2587;
  assign n35361 = n2611 & n35360;
  assign n35362 = n2587 & n35359;
  assign n35363 = n2621 & n64336;
  assign n35364 = n62346 & n35358;
  assign n35365 = ~pi69 & n64337;
  assign n35366 = ~pi67 & ~pi71;
  assign n35367 = pi36 & ~pi103;
  assign n35368 = n35366 & n35367;
  assign n35369 = n35365 & n35368;
  assign n35370 = n35357 & n35369;
  assign n35371 = n2684 & n35370;
  assign n35372 = n35356 & ~n35371;
  assign n35373 = n30715 & ~n35372;
  assign n35374 = ~pi97 & ~n35373;
  assign n35375 = ~pi46 & n62395;
  assign n35376 = n30938 & n35375;
  assign n35377 = ~n35374 & n35376;
  assign n35378 = n30716 & ~n35356;
  assign n35379 = ~n62395 & n35378;
  assign n35380 = pi299 & n34094;
  assign n35381 = ~n34083 & ~n35380;
  assign n35382 = n2815 & ~n35381;
  assign n35383 = pi109 & ~n35382;
  assign n35384 = ~n35379 & ~n35383;
  assign n35385 = ~n35377 & n35384;
  assign n35386 = ~n2870 & n35382;
  assign n35387 = ~n30749 & ~n35382;
  assign n35388 = ~n35386 & ~n35387;
  assign n35389 = ~n35385 & n35388;
  assign n35390 = ~pi91 & ~n35389;
  assign n35391 = n2715 & ~n30721;
  assign n35392 = ~n35390 & n35391;
  assign n35393 = ~n35354 & ~n35392;
  assign n35394 = ~pi32 & n32019;
  assign n35395 = ~pi39 & n62366;
  assign n35396 = n2726 & n35394;
  assign n35397 = ~pi39 & n2728;
  assign n35398 = ~pi96 & n64339;
  assign n35399 = n2730 & n35394;
  assign n35400 = n62366 & n2743;
  assign n35401 = ~pi39 & n35400;
  assign n35402 = n2743 & n64338;
  assign n35403 = ~n35393 & n64340;
  assign n35404 = ~n35353 & ~n35403;
  assign n35405 = ~pi38 & ~n35404;
  assign n35406 = ~pi228 & n35405;
  assign n35407 = ~n35346 & ~n35406;
  assign n35408 = ~pi100 & ~n35407;
  assign n35409 = ~n34060 & ~n35346;
  assign n35410 = pi100 & ~n35409;
  assign n35411 = ~pi87 & ~n35410;
  assign n35412 = ~n35408 & n35411;
  assign n35413 = pi87 & ~n35346;
  assign n35414 = ~pi75 & ~n35413;
  assign n35415 = ~n35412 & n35414;
  assign n35416 = ~n64304 & ~n35346;
  assign n35417 = pi75 & ~n35416;
  assign n35418 = ~pi92 & ~n35417;
  assign n35419 = ~n35415 & n35418;
  assign n35420 = n62373 & n34059;
  assign n35421 = n6795 & n35420;
  assign n35422 = ~pi75 & n64304;
  assign n35423 = n64083 & n34059;
  assign n35424 = pi92 & ~n35346;
  assign n35425 = ~n64341 & n35424;
  assign n35426 = n35113 & ~n35425;
  assign n35427 = ~n35419 & n35426;
  assign n35428 = ~n35347 & ~n35427;
  assign n35429 = pi743 & pi947;
  assign n35430 = pi907 & ~pi947;
  assign n35431 = pi735 & n35430;
  assign n35432 = ~n35429 & ~n35431;
  assign n35433 = n2923 & n35432;
  assign n35434 = ~pi146 & ~n2923;
  assign n35435 = pi832 & ~n35434;
  assign n35436 = ~n35433 & n35435;
  assign n35437 = n62787 & ~n35432;
  assign n35438 = pi146 & ~n62953;
  assign n35439 = pi146 & ~n62787;
  assign n35440 = ~n2916 & n35439;
  assign n35441 = pi146 & ~n7104;
  assign n35442 = n2916 & n35441;
  assign n35443 = pi735 & pi907;
  assign n35444 = n62787 & n35443;
  assign n35445 = ~pi947 & ~n35444;
  assign n35446 = ~n35442 & n35445;
  assign n35447 = pi743 & n62787;
  assign n35448 = pi947 & ~n35439;
  assign n35449 = ~n35447 & n35448;
  assign n35450 = ~n35446 & ~n35449;
  assign n35451 = ~n35440 & ~n35450;
  assign n35452 = ~n35437 & ~n35438;
  assign n35453 = ~n7118 & ~n64342;
  assign n35454 = n6951 & ~n35432;
  assign n35455 = pi146 & ~n6951;
  assign n35456 = ~pi146 & ~n6951;
  assign n35457 = n6951 & n35432;
  assign n35458 = ~n35456 & ~n35457;
  assign n35459 = ~n35454 & ~n35455;
  assign n35460 = n7118 & n64343;
  assign n35461 = ~pi215 & ~n35460;
  assign n35462 = ~n35453 & n35461;
  assign n35463 = pi146 & n7139;
  assign n35464 = n7002 & ~n35432;
  assign n35465 = pi215 & ~n35464;
  assign n35466 = ~n35463 & n35465;
  assign n35467 = pi299 & ~n35466;
  assign n35468 = ~n35462 & n35467;
  assign n35469 = n7104 & ~n35432;
  assign n35470 = n2971 & ~n35441;
  assign n35471 = ~n35469 & n35470;
  assign n35472 = ~n2971 & ~n35439;
  assign n35473 = ~n2971 & ~n35437;
  assign n35474 = ~n35439 & n35473;
  assign n35475 = ~n35437 & n35472;
  assign n35476 = ~n7034 & ~n64344;
  assign n35477 = ~n35437 & ~n35439;
  assign n35478 = ~n2971 & ~n35477;
  assign n35479 = n7104 & n35432;
  assign n35480 = ~pi146 & ~n7104;
  assign n35481 = n2971 & ~n35480;
  assign n35482 = ~n35479 & n35481;
  assign n35483 = ~n35471 & ~n64344;
  assign n35484 = ~n35478 & ~n35482;
  assign n35485 = ~n7034 & n64345;
  assign n35486 = ~n35471 & n35476;
  assign n35487 = n7034 & n64343;
  assign n35488 = ~pi223 & ~n35487;
  assign n35489 = ~n64346 & n35488;
  assign n35490 = pi146 & ~n7002;
  assign n35491 = ~n35464 & ~n35490;
  assign n35492 = ~n2971 & ~n35491;
  assign n35493 = n62784 & n35432;
  assign n35494 = ~pi146 & ~n62784;
  assign n35495 = n2971 & ~n35494;
  assign n35496 = n2971 & ~n35493;
  assign n35497 = ~n35494 & n35496;
  assign n35498 = ~n35493 & n35495;
  assign n35499 = pi223 & ~n64347;
  assign n35500 = ~n35492 & n35499;
  assign n35501 = ~pi299 & ~n35500;
  assign n35502 = ~n35489 & n35501;
  assign n35503 = pi39 & ~n35502;
  assign n35504 = ~n35489 & ~n35500;
  assign n35505 = ~n7034 & ~n64345;
  assign n35506 = n7034 & ~n64343;
  assign n35507 = ~pi223 & ~n35506;
  assign n35508 = ~n35505 & n35507;
  assign n35509 = ~n35492 & ~n64347;
  assign n35510 = pi223 & ~n35509;
  assign n35511 = ~pi299 & ~n35510;
  assign n35512 = ~n35508 & n35511;
  assign n35513 = ~pi299 & ~n35504;
  assign n35514 = ~n7118 & ~n35437;
  assign n35515 = ~n35438 & n35514;
  assign n35516 = n7118 & ~n64343;
  assign n35517 = ~pi215 & ~n35516;
  assign n35518 = ~n35515 & n35517;
  assign n35519 = ~n35463 & ~n35464;
  assign n35520 = pi215 & ~n35519;
  assign n35521 = pi299 & ~n35520;
  assign n35522 = ~n35462 & ~n35466;
  assign n35523 = pi299 & ~n35522;
  assign n35524 = ~n35518 & n35521;
  assign n35525 = ~n64348 & ~n64349;
  assign n35526 = pi39 & ~n35525;
  assign n35527 = ~n35468 & n35503;
  assign n35528 = n6936 & ~n35432;
  assign n35529 = pi146 & ~n6936;
  assign n35530 = pi299 & ~n35529;
  assign n35531 = ~n35528 & n35530;
  assign n35532 = n6940 & ~n35432;
  assign n35533 = pi146 & ~n6940;
  assign n35534 = ~pi299 & ~n35533;
  assign n35535 = ~n35532 & n35534;
  assign n35536 = ~n35531 & ~n35535;
  assign n35537 = ~pi146 & ~n6940;
  assign n35538 = n6940 & n35432;
  assign n35539 = ~pi299 & ~n35538;
  assign n35540 = ~pi299 & ~n35537;
  assign n35541 = ~n35538 & n35540;
  assign n35542 = ~n35537 & n35539;
  assign n35543 = ~pi146 & ~n6936;
  assign n35544 = n6936 & n35432;
  assign n35545 = pi299 & ~n35544;
  assign n35546 = pi299 & ~n35543;
  assign n35547 = ~n35544 & n35546;
  assign n35548 = ~n35543 & n35545;
  assign n35549 = ~pi39 & ~n64352;
  assign n35550 = ~n64351 & n35549;
  assign n35551 = ~pi39 & ~n64351;
  assign n35552 = ~n64352 & n35551;
  assign n35553 = ~pi39 & ~n35536;
  assign n35554 = ~pi38 & ~n64353;
  assign n35555 = ~n64350 & n35554;
  assign n35556 = ~pi146 & ~n7357;
  assign n35557 = n7357 & n35432;
  assign n35558 = n7356 & n35433;
  assign n35559 = pi38 & ~n64354;
  assign n35560 = pi38 & ~n35556;
  assign n35561 = ~n64354 & n35560;
  assign n35562 = ~n35556 & n35559;
  assign n35563 = n63888 & ~n64355;
  assign n35564 = ~n35555 & n35563;
  assign n35565 = ~pi146 & ~n63888;
  assign n35566 = ~pi832 & ~n35565;
  assign n35567 = ~n35564 & n35566;
  assign n35568 = ~n35436 & ~n35567;
  assign n35569 = ~pi770 & pi947;
  assign n35570 = pi726 & n35430;
  assign n35571 = ~n35569 & ~n35570;
  assign n35572 = n2923 & ~n35571;
  assign n35573 = ~pi147 & ~n2923;
  assign n35574 = pi832 & ~n35573;
  assign n35575 = ~n35572 & n35574;
  assign n35576 = pi215 & ~n7138;
  assign n35577 = n7126 & ~n35430;
  assign n35578 = pi947 & n62787;
  assign n35579 = ~n7122 & ~n35578;
  assign n35580 = ~n7118 & ~n35579;
  assign n35581 = ~pi215 & ~n35580;
  assign n35582 = ~n35577 & n35581;
  assign n35583 = ~n35576 & ~n35582;
  assign n35584 = pi299 & ~n35583;
  assign n35585 = ~n7110 & ~n62790;
  assign n35586 = n2915 & ~n35585;
  assign n35587 = ~pi223 & ~n35586;
  assign n35588 = ~pi947 & ~n62785;
  assign n35589 = pi223 & ~n35588;
  assign n35590 = ~n62785 & ~n35430;
  assign n35591 = pi223 & ~n35590;
  assign n35592 = ~n35589 & ~n35591;
  assign n35593 = ~n35587 & n35592;
  assign n35594 = ~pi299 & ~n35593;
  assign n35595 = pi299 & pi947;
  assign n35596 = ~n35594 & ~n35595;
  assign n35597 = ~n35584 & ~n35595;
  assign n35598 = ~n35594 & n35597;
  assign n35599 = ~n35584 & n35596;
  assign n35600 = pi39 & n64356;
  assign n35601 = ~n2915 & ~n62781;
  assign n35602 = ~pi39 & ~n35601;
  assign n35603 = ~n62781 & n35602;
  assign n35604 = ~n35600 & ~n35603;
  assign n35605 = ~pi147 & n35604;
  assign n35606 = pi215 & ~n7134;
  assign n35607 = ~n2915 & n6951;
  assign n35608 = ~n2915 & n7126;
  assign n35609 = n7118 & n35607;
  assign n35610 = ~pi215 & ~n64357;
  assign n35611 = n7118 & ~n35607;
  assign n35612 = ~n7129 & ~n35611;
  assign n35613 = ~pi215 & ~n35612;
  assign n35614 = ~n7125 & n35610;
  assign n35615 = ~n35606 & ~n64358;
  assign n35616 = pi299 & ~n35615;
  assign n35617 = ~n2915 & n7116;
  assign n35618 = ~pi299 & ~n35617;
  assign n35619 = ~pi299 & n7116;
  assign n35620 = ~n2915 & n35619;
  assign n35621 = ~pi299 & n35617;
  assign n35622 = pi299 & ~n64358;
  assign n35623 = pi299 & ~n35606;
  assign n35624 = ~n64358 & n35623;
  assign n35625 = ~n35606 & n35622;
  assign n35626 = ~n64359 & ~n64360;
  assign n35627 = ~n35616 & ~n35618;
  assign n35628 = pi39 & n64361;
  assign n35629 = ~n35602 & ~n35628;
  assign n35630 = pi147 & n35629;
  assign n35631 = ~pi38 & ~n35630;
  assign n35632 = ~n35605 & n35631;
  assign n35633 = n2915 & n7357;
  assign n35634 = ~pi147 & ~n35633;
  assign n35635 = ~n2915 & n7357;
  assign n35636 = pi38 & ~n35635;
  assign n35637 = ~n35634 & n35636;
  assign n35638 = ~pi770 & ~n35637;
  assign n35639 = ~n35632 & n35638;
  assign n35640 = pi215 & pi947;
  assign n35641 = n7002 & n35640;
  assign n35642 = ~n35583 & ~n35641;
  assign n35643 = pi299 & ~n35642;
  assign n35644 = ~pi299 & ~n35430;
  assign n35645 = ~n35430 & n35619;
  assign n35646 = n7116 & n35644;
  assign n35647 = ~n35643 & ~n64362;
  assign n35648 = pi39 & ~n35647;
  assign n35649 = ~n62781 & ~n35430;
  assign n35650 = ~pi39 & n35649;
  assign n35651 = ~n35648 & ~n35650;
  assign n35652 = ~pi147 & n35651;
  assign n35653 = n7002 & n35430;
  assign n35654 = pi215 & ~n35653;
  assign n35655 = n62787 & n35430;
  assign n35656 = ~n7118 & ~n35655;
  assign n35657 = pi907 & n6951;
  assign n35658 = ~pi947 & n35657;
  assign n35659 = n7118 & ~n35658;
  assign n35660 = ~n35656 & ~n35659;
  assign n35661 = ~pi215 & ~n35660;
  assign n35662 = ~n35654 & ~n35661;
  assign n35663 = pi299 & ~n35662;
  assign n35664 = n7116 & n35430;
  assign n35665 = ~pi299 & ~n35664;
  assign n35666 = ~n35663 & ~n35665;
  assign n35667 = pi39 & ~n35666;
  assign n35668 = ~n62781 & n35430;
  assign n35669 = ~pi39 & ~n35668;
  assign n35670 = ~n35667 & ~n35669;
  assign n35671 = pi147 & n35670;
  assign n35672 = ~pi38 & ~n35671;
  assign n35673 = ~n35652 & n35672;
  assign n35674 = ~pi147 & ~n7357;
  assign n35675 = n7357 & n35430;
  assign n35676 = pi38 & ~n35675;
  assign n35677 = ~n35674 & n35676;
  assign n35678 = pi770 & ~n35677;
  assign n35679 = ~n35673 & n35678;
  assign n35680 = pi726 & ~n35679;
  assign n35681 = pi726 & ~n35639;
  assign n35682 = ~n35679 & n35681;
  assign n35683 = ~n35639 & n35680;
  assign n35684 = pi947 & n7116;
  assign n35685 = pi947 & n35619;
  assign n35686 = ~pi299 & n35684;
  assign n35687 = ~pi947 & n7126;
  assign n35688 = ~n7122 & ~n35655;
  assign n35689 = ~n7118 & ~n35688;
  assign n35690 = ~pi215 & ~n35689;
  assign n35691 = ~n35687 & n35690;
  assign n35692 = n35576 & ~n35653;
  assign n35693 = ~n35691 & ~n35692;
  assign n35694 = pi299 & ~n35693;
  assign n35695 = ~n7117 & ~n35694;
  assign n35696 = ~n64364 & n35695;
  assign n35697 = pi39 & ~n35696;
  assign n35698 = ~pi947 & ~n62781;
  assign n35699 = ~pi39 & ~n35698;
  assign n35700 = ~pi38 & ~n35699;
  assign n35701 = ~n35697 & ~n35699;
  assign n35702 = ~pi38 & n35701;
  assign n35703 = ~n35697 & n35700;
  assign n35704 = pi38 & ~pi947;
  assign n35705 = n7357 & n35704;
  assign n35706 = ~n64365 & ~n35705;
  assign n35707 = ~pi770 & ~n35706;
  assign n35708 = ~pi147 & ~n21074;
  assign n35709 = ~pi770 & n35706;
  assign n35710 = ~n21080 & ~n35709;
  assign n35711 = ~pi147 & ~n35710;
  assign n35712 = ~n35707 & n35708;
  assign n35713 = ~n8089 & ~n35705;
  assign n35714 = pi947 & ~n62781;
  assign n35715 = ~pi39 & ~n35714;
  assign n35716 = ~pi299 & ~n35684;
  assign n35717 = pi299 & ~n35641;
  assign n35718 = ~n7118 & ~n35578;
  assign n35719 = pi947 & n6951;
  assign n35720 = n7118 & ~n35719;
  assign n35721 = ~pi215 & ~n35720;
  assign n35722 = ~n35718 & n35721;
  assign n35723 = n35717 & ~n35722;
  assign n35724 = ~n35716 & ~n35723;
  assign n35725 = pi39 & ~n35724;
  assign n35726 = ~n35715 & ~n35725;
  assign n35727 = ~pi38 & ~n35726;
  assign n35728 = n35713 & ~n35727;
  assign n35729 = pi147 & ~pi770;
  assign n35730 = n35728 & n35729;
  assign n35731 = ~pi726 & ~n35730;
  assign n35732 = ~n64366 & n35731;
  assign n35733 = n63888 & ~n35732;
  assign n35734 = n63888 & ~n64363;
  assign n35735 = ~n35732 & n35734;
  assign n35736 = ~n64363 & n35733;
  assign n35737 = ~pi147 & ~n63888;
  assign n35738 = ~pi832 & ~n35737;
  assign n35739 = ~n64367 & n35738;
  assign po304 = ~n35575 & ~n35739;
  assign n35741 = pi749 & pi947;
  assign n35742 = n2923 & ~n35741;
  assign n35743 = pi706 & n35430;
  assign n35744 = n35742 & ~n35743;
  assign n35745 = pi148 & ~n2923;
  assign n35746 = pi832 & ~n35745;
  assign n35747 = ~n35744 & n35746;
  assign n35748 = ~pi148 & n64356;
  assign n35749 = pi148 & n64361;
  assign n35750 = pi749 & ~n35749;
  assign n35751 = ~n35748 & n35750;
  assign n35752 = ~n31412 & ~n35647;
  assign n35753 = ~n7117 & ~n35663;
  assign n35754 = pi148 & ~n35753;
  assign n35755 = ~pi749 & ~n35754;
  assign n35756 = ~n35752 & n35755;
  assign n35757 = pi39 & ~n35756;
  assign n35758 = ~n35752 & ~n35754;
  assign n35759 = ~pi749 & ~n35758;
  assign n35760 = ~pi148 & ~n64356;
  assign n35761 = pi148 & ~n64361;
  assign n35762 = pi749 & ~n35761;
  assign n35763 = ~n35760 & n35762;
  assign n35764 = ~n35759 & ~n35763;
  assign n35765 = pi39 & ~n35764;
  assign n35766 = pi39 & ~n35751;
  assign n35767 = ~n35756 & n35766;
  assign n35768 = ~n35751 & n35757;
  assign n35769 = ~pi148 & n62781;
  assign n35770 = ~pi39 & ~n35769;
  assign n35771 = ~pi749 & pi947;
  assign n35772 = n35601 & ~n35771;
  assign n35773 = n35770 & ~n35772;
  assign n35774 = ~pi38 & ~n35773;
  assign n35775 = ~n64368 & n35774;
  assign n35776 = n35635 & ~n35771;
  assign n35777 = ~pi148 & ~n7357;
  assign n35778 = ~n35776 & ~n35777;
  assign n35779 = pi38 & ~n35778;
  assign n35780 = pi706 & ~n35779;
  assign n35781 = ~n35775 & n35780;
  assign n35782 = ~pi148 & ~n35693;
  assign n35783 = ~n35641 & ~n35722;
  assign n35784 = pi148 & ~n35783;
  assign n35785 = pi299 & ~n35784;
  assign n35786 = ~n35782 & n35785;
  assign n35787 = ~pi148 & ~n7116;
  assign n35788 = n35716 & ~n35787;
  assign n35789 = pi749 & ~n35788;
  assign n35790 = ~n35786 & n35789;
  assign n35791 = ~pi148 & ~pi749;
  assign n35792 = ~n7143 & n35791;
  assign n35793 = pi39 & ~n35792;
  assign n35794 = ~n35790 & n35793;
  assign n35795 = ~n62781 & n35741;
  assign n35796 = n35770 & ~n35795;
  assign n35797 = ~pi38 & ~n35796;
  assign n35798 = ~n35794 & n35797;
  assign n35799 = pi148 & ~n7357;
  assign n35800 = n7357 & ~n35741;
  assign n35801 = n7356 & n35742;
  assign n35802 = pi38 & ~n64369;
  assign n35803 = ~n35799 & n35802;
  assign n35804 = ~pi706 & ~n35803;
  assign n35805 = ~n35798 & n35804;
  assign n35806 = n27338 & ~n35805;
  assign n35807 = ~n35781 & n35806;
  assign n35808 = ~pi148 & ~n27338;
  assign n35809 = ~pi57 & ~n35808;
  assign n35810 = ~n35807 & n35809;
  assign n35811 = pi57 & pi148;
  assign n35812 = ~pi832 & ~n35811;
  assign n35813 = ~n35810 & n35812;
  assign n35814 = ~n35747 & ~n35813;
  assign n35815 = ~pi149 & n64356;
  assign n35816 = pi149 & n64361;
  assign n35817 = ~pi755 & ~n35816;
  assign n35818 = ~n35815 & n35817;
  assign n35819 = ~pi149 & n35643;
  assign n35820 = pi149 & ~n35753;
  assign n35821 = pi755 & ~n64362;
  assign n35822 = ~n35820 & n35821;
  assign n35823 = ~n35819 & n35822;
  assign n35824 = pi39 & ~n35823;
  assign n35825 = ~n64362 & ~n35820;
  assign n35826 = ~n35819 & n35825;
  assign n35827 = pi755 & ~n35826;
  assign n35828 = ~pi149 & ~n64356;
  assign n35829 = pi149 & ~n64361;
  assign n35830 = ~pi755 & ~n35829;
  assign n35831 = ~n35828 & n35830;
  assign n35832 = ~n35827 & ~n35831;
  assign n35833 = pi39 & ~n35832;
  assign n35834 = ~n35818 & n35824;
  assign n35835 = ~pi755 & pi947;
  assign n35836 = ~n62781 & n35835;
  assign n35837 = ~pi149 & n62781;
  assign n35838 = ~pi39 & ~n35837;
  assign n35839 = ~pi39 & ~n35836;
  assign n35840 = ~n35837 & n35839;
  assign n35841 = ~n35836 & n35838;
  assign n35842 = ~n35668 & n64371;
  assign n35843 = ~pi38 & ~n35842;
  assign n35844 = ~n64370 & n35843;
  assign n35845 = n7357 & ~n35835;
  assign n35846 = ~n35430 & n35845;
  assign n35847 = pi149 & ~n7357;
  assign n35848 = pi38 & ~n35847;
  assign n35849 = ~n35846 & n35848;
  assign n35850 = ~pi725 & ~n35849;
  assign n35851 = ~n35844 & n35850;
  assign n35852 = ~pi149 & ~n35693;
  assign n35853 = ~pi149 & pi299;
  assign n35854 = ~n35723 & ~n35853;
  assign n35855 = ~n35852 & ~n35854;
  assign n35856 = ~pi149 & ~n7116;
  assign n35857 = n35716 & ~n35856;
  assign n35858 = ~pi755 & ~n35857;
  assign n35859 = ~n35855 & n35858;
  assign n35860 = ~pi149 & pi755;
  assign n35861 = ~n7143 & n35860;
  assign n35862 = pi39 & ~n35861;
  assign n35863 = ~n35859 & n35862;
  assign n35864 = ~pi38 & ~n64371;
  assign n35865 = ~n35863 & n35864;
  assign n35866 = pi38 & ~n35845;
  assign n35867 = ~n35847 & n35866;
  assign n35868 = pi725 & ~n35867;
  assign n35869 = ~n35865 & n35868;
  assign n35870 = n63888 & ~n35869;
  assign n35871 = ~n35865 & ~n35867;
  assign n35872 = pi725 & ~n35871;
  assign n35873 = ~n64370 & ~n35842;
  assign n35874 = ~pi38 & ~n35873;
  assign n35875 = ~pi149 & ~n7357;
  assign n35876 = ~n2915 & n6955;
  assign n35877 = pi755 & pi947;
  assign n35878 = ~pi39 & ~n35877;
  assign n35879 = ~n35430 & ~n35835;
  assign n35880 = n7357 & ~n35879;
  assign n35881 = n35876 & n35878;
  assign n35882 = pi38 & ~n64372;
  assign n35883 = pi38 & ~n35875;
  assign n35884 = ~n64372 & n35883;
  assign n35885 = ~n35875 & n35882;
  assign n35886 = ~pi725 & ~n64373;
  assign n35887 = ~n35874 & n35886;
  assign n35888 = ~n35872 & ~n35887;
  assign n35889 = n63888 & ~n35888;
  assign n35890 = ~n35851 & n35870;
  assign n35891 = ~pi149 & ~n63888;
  assign n35892 = ~pi832 & ~n35891;
  assign n35893 = ~n64374 & n35892;
  assign n35894 = ~pi725 & n35430;
  assign n35895 = ~n35835 & ~n35894;
  assign n35896 = n2923 & ~n35895;
  assign n35897 = ~pi149 & ~n2923;
  assign n35898 = pi832 & ~n35897;
  assign n35899 = ~n35896 & n35898;
  assign po306 = ~n35893 & ~n35899;
  assign n35901 = ~pi751 & pi947;
  assign n35902 = ~pi701 & n35430;
  assign n35903 = ~n35901 & ~n35902;
  assign n35904 = pi701 & ~n35901;
  assign n35905 = ~n35430 & ~n35901;
  assign n35906 = n2923 & ~n35905;
  assign n35907 = ~n35904 & n35906;
  assign n35908 = n2923 & ~n35903;
  assign n35909 = ~pi150 & ~n2923;
  assign n35910 = pi832 & ~n35909;
  assign n35911 = ~n64375 & n35910;
  assign n35912 = ~pi150 & ~n64356;
  assign n35913 = pi150 & ~n64361;
  assign n35914 = ~pi751 & ~n35913;
  assign n35915 = ~n35912 & n35914;
  assign n35916 = ~pi150 & n35647;
  assign n35917 = pi150 & n35666;
  assign n35918 = pi751 & ~n35917;
  assign n35919 = ~n35916 & n35918;
  assign n35920 = pi39 & ~n35919;
  assign n35921 = ~pi150 & ~n35647;
  assign n35922 = pi150 & ~n35666;
  assign n35923 = pi751 & ~n35922;
  assign n35924 = ~n35921 & n35923;
  assign n35925 = ~pi150 & n64356;
  assign n35926 = pi150 & n64361;
  assign n35927 = ~pi751 & ~n35926;
  assign n35928 = ~n35925 & n35927;
  assign n35929 = ~n35924 & ~n35928;
  assign n35930 = pi39 & ~n35929;
  assign n35931 = ~n35915 & n35920;
  assign n35932 = n35649 & ~n35901;
  assign n35933 = pi150 & n62781;
  assign n35934 = ~pi39 & ~n35933;
  assign n35935 = ~n35932 & n35934;
  assign n35936 = ~pi38 & ~n35935;
  assign n35937 = ~n64376 & n35936;
  assign n35938 = ~pi150 & ~n7357;
  assign n35939 = pi751 & pi947;
  assign n35940 = ~pi39 & ~n35939;
  assign n35941 = n35876 & n35940;
  assign n35942 = n7357 & ~n35905;
  assign n35943 = n7356 & n35906;
  assign n35944 = pi38 & ~n64377;
  assign n35945 = pi150 & ~n7357;
  assign n35946 = n7357 & ~n35901;
  assign n35947 = ~n35430 & n35946;
  assign n35948 = ~n35945 & ~n35947;
  assign n35949 = pi38 & ~n35948;
  assign n35950 = pi38 & ~n35938;
  assign n35951 = ~n64377 & n35950;
  assign n35952 = ~n35938 & n35944;
  assign n35953 = ~pi701 & ~n64378;
  assign n35954 = ~n35937 & n35953;
  assign n35955 = ~pi150 & n35696;
  assign n35956 = pi150 & ~n35724;
  assign n35957 = ~pi751 & ~n35956;
  assign n35958 = ~n35955 & n35957;
  assign n35959 = ~pi150 & pi751;
  assign n35960 = ~n7143 & n35959;
  assign n35961 = ~n35958 & ~n35960;
  assign n35962 = pi39 & ~n35961;
  assign n35963 = ~n19832 & ~n35933;
  assign n35964 = n35699 & n35963;
  assign n35965 = ~pi38 & ~n35964;
  assign n35966 = ~n35962 & n35965;
  assign n35967 = ~n35945 & ~n35946;
  assign n35968 = pi38 & ~n35967;
  assign n35969 = pi701 & ~n35968;
  assign n35970 = ~n35966 & n35969;
  assign n35971 = ~n35954 & ~n35970;
  assign n35972 = n63888 & ~n35971;
  assign n35973 = ~pi150 & ~n63888;
  assign n35974 = ~pi832 & ~n35973;
  assign n35975 = ~n35972 & n35974;
  assign po307 = ~n35911 & ~n35975;
  assign n35977 = ~pi745 & pi947;
  assign n35978 = ~pi723 & n35430;
  assign n35979 = ~n35977 & ~n35978;
  assign n35980 = n2923 & ~n35979;
  assign n35981 = ~pi151 & ~n2923;
  assign n35982 = pi832 & ~n35981;
  assign n35983 = ~n35980 & n35982;
  assign n35984 = ~pi745 & ~n7117;
  assign n35985 = ~pi151 & ~n7143;
  assign n35986 = ~n35984 & n35985;
  assign n35987 = ~pi151 & ~n6951;
  assign n35988 = n35720 & ~n35987;
  assign n35989 = pi151 & ~n7118;
  assign n35990 = pi151 & n7129;
  assign n35991 = ~n7124 & n35989;
  assign n35992 = ~n7123 & ~n64379;
  assign n35993 = ~n35988 & n35992;
  assign n35994 = n35690 & n35993;
  assign n35995 = ~n7138 & ~n35653;
  assign n35996 = ~pi151 & n35995;
  assign n35997 = ~n7134 & ~n35996;
  assign n35998 = pi215 & ~n35997;
  assign n35999 = ~n35653 & n35998;
  assign n36000 = n35654 & ~n35997;
  assign n36001 = pi299 & ~n64380;
  assign n36002 = ~n35994 & n36001;
  assign n36003 = ~pi745 & ~n35716;
  assign n36004 = ~n36002 & n36003;
  assign n36005 = ~n35986 & ~n36004;
  assign n36006 = pi39 & ~n36005;
  assign n36007 = ~pi151 & n62781;
  assign n36008 = ~pi745 & n35714;
  assign n36009 = ~n36007 & ~n36008;
  assign n36010 = ~pi39 & ~n36009;
  assign n36011 = ~pi38 & ~n36010;
  assign n36012 = ~n36006 & n36011;
  assign n36013 = n7357 & ~n35977;
  assign n36014 = pi151 & ~n7357;
  assign n36015 = ~n36013 & ~n36014;
  assign n36016 = pi38 & ~n36015;
  assign n36017 = pi723 & ~n36016;
  assign n36018 = ~n36012 & n36017;
  assign n36019 = n35669 & n36009;
  assign n36020 = pi151 & ~n35617;
  assign n36021 = n35594 & ~n36020;
  assign n36022 = n35659 & ~n35987;
  assign n36023 = ~n35607 & n36022;
  assign n36024 = ~pi215 & ~n36023;
  assign n36025 = n35992 & n36024;
  assign n36026 = ~n35998 & ~n36025;
  assign n36027 = pi299 & ~n36026;
  assign n36028 = ~n36021 & ~n36027;
  assign n36029 = ~pi745 & ~n36028;
  assign n36030 = n35992 & ~n36022;
  assign n36031 = n35581 & n36030;
  assign n36032 = ~n35998 & ~n36031;
  assign n36033 = ~n35641 & ~n36032;
  assign n36034 = pi299 & ~n36033;
  assign n36035 = ~pi151 & ~n7116;
  assign n36036 = n35665 & ~n36035;
  assign n36037 = pi745 & ~n36036;
  assign n36038 = ~n36034 & n36037;
  assign n36039 = pi39 & ~n36038;
  assign n36040 = ~n36034 & ~n36036;
  assign n36041 = pi745 & ~n36040;
  assign n36042 = ~pi745 & ~n36027;
  assign n36043 = ~n36021 & n36042;
  assign n36044 = ~n36041 & ~n36043;
  assign n36045 = pi39 & ~n36044;
  assign n36046 = ~n36029 & n36039;
  assign n36047 = ~n36019 & ~n64381;
  assign n36048 = ~pi38 & ~n36047;
  assign n36049 = pi745 & pi947;
  assign n36050 = ~pi39 & ~n36049;
  assign n36051 = ~n35430 & ~n35977;
  assign n36052 = n7357 & ~n36051;
  assign n36053 = n35876 & n36050;
  assign n36054 = ~pi151 & ~n7357;
  assign n36055 = pi38 & ~n36054;
  assign n36056 = ~n35430 & n36013;
  assign n36057 = ~n36014 & ~n36056;
  assign n36058 = pi38 & ~n36057;
  assign n36059 = pi38 & ~n64382;
  assign n36060 = ~n36054 & n36059;
  assign n36061 = ~n64382 & n36055;
  assign n36062 = ~pi723 & ~n64383;
  assign n36063 = ~n36048 & n36062;
  assign n36064 = ~n36018 & ~n36063;
  assign n36065 = n63888 & ~n36064;
  assign n36066 = ~pi151 & ~n63888;
  assign n36067 = ~pi832 & ~n36066;
  assign n36068 = ~n36065 & n36067;
  assign po308 = ~n35983 & ~n36068;
  assign n36070 = ~pi152 & ~n62789;
  assign n36071 = ~pi947 & n62789;
  assign n36072 = ~n7034 & ~n36071;
  assign n36073 = ~n36070 & n36072;
  assign n36074 = ~n2915 & n62789;
  assign n36075 = ~n7034 & ~n36074;
  assign n36076 = ~n36073 & n36075;
  assign n36077 = pi152 & ~n6951;
  assign n36078 = ~n35607 & ~n36077;
  assign n36079 = n7034 & n36078;
  assign n36080 = ~pi223 & ~n36079;
  assign n36081 = ~n36076 & n36080;
  assign n36082 = ~pi152 & n62785;
  assign n36083 = n35591 & ~n36082;
  assign n36084 = ~pi299 & ~n36083;
  assign n36085 = n35589 & ~n36082;
  assign n36086 = ~pi299 & ~n36085;
  assign n36087 = ~n36083 & n36086;
  assign n36088 = n36084 & ~n36085;
  assign n36089 = ~n36081 & n64384;
  assign n36090 = n7118 & n36078;
  assign n36091 = ~pi215 & ~n36090;
  assign n36092 = pi152 & n35579;
  assign n36093 = n35656 & ~n36092;
  assign n36094 = ~n7124 & n36093;
  assign n36095 = n36091 & ~n36094;
  assign n36096 = ~pi152 & ~n7134;
  assign n36097 = n35576 & ~n36096;
  assign n36098 = pi299 & ~n36097;
  assign n36099 = ~n36095 & n36098;
  assign n36100 = pi759 & ~n36099;
  assign n36101 = pi759 & ~n36089;
  assign n36102 = ~n36099 & n36101;
  assign n36103 = ~n36089 & n36100;
  assign n36104 = ~n35658 & ~n36077;
  assign n36105 = n7034 & ~n36104;
  assign n36106 = n62789 & ~n35430;
  assign n36107 = ~n7034 & ~n36106;
  assign n36108 = ~n36070 & n36107;
  assign n36109 = ~n36105 & ~n36108;
  assign n36110 = ~pi223 & ~n36109;
  assign n36111 = n36084 & ~n36110;
  assign n36112 = ~n35577 & n36091;
  assign n36113 = ~n36093 & n36112;
  assign n36114 = ~n35430 & ~n35606;
  assign n36115 = n36097 & ~n36114;
  assign n36116 = pi299 & ~n36115;
  assign n36117 = ~n36113 & n36116;
  assign n36118 = ~pi759 & ~n36117;
  assign n36119 = ~n36111 & n36118;
  assign n36120 = pi39 & ~n36119;
  assign n36121 = ~n64385 & n36120;
  assign n36122 = pi759 & n35714;
  assign n36123 = pi152 & n62781;
  assign n36124 = ~pi39 & ~n36123;
  assign n36125 = pi759 & pi947;
  assign n36126 = ~pi39 & ~n36125;
  assign n36127 = ~n7145 & ~n36126;
  assign n36128 = ~n36123 & ~n36127;
  assign n36129 = ~n36122 & n36124;
  assign n36130 = ~n35668 & n64386;
  assign n36131 = ~pi38 & ~n36130;
  assign n36132 = ~n36121 & n36131;
  assign n36133 = n6955 & ~n35430;
  assign n36134 = n7357 & ~n36125;
  assign n36135 = ~n35430 & n36134;
  assign n36136 = n36126 & n36133;
  assign n36137 = ~pi152 & ~n7357;
  assign n36138 = pi38 & ~n36137;
  assign n36139 = pi38 & ~n64387;
  assign n36140 = ~n36137 & n36139;
  assign n36141 = ~n64387 & n36138;
  assign n36142 = pi696 & ~n64388;
  assign n36143 = ~n36132 & n36142;
  assign n36144 = ~n35689 & ~n36093;
  assign n36145 = ~n35578 & ~n36144;
  assign n36146 = ~n35719 & ~n36077;
  assign n36147 = n7118 & n36146;
  assign n36148 = ~pi215 & ~n36147;
  assign n36149 = ~n36145 & n36148;
  assign n36150 = pi152 & n35692;
  assign n36151 = n35717 & ~n36150;
  assign n36152 = ~n36149 & n36151;
  assign n36153 = n7034 & ~n36146;
  assign n36154 = ~n36073 & ~n36153;
  assign n36155 = ~pi223 & ~n36154;
  assign n36156 = n36086 & ~n36155;
  assign n36157 = pi759 & ~n36156;
  assign n36158 = ~n36152 & n36157;
  assign n36159 = pi152 & n12805;
  assign n36160 = pi39 & ~n36159;
  assign n36161 = ~n36158 & n36160;
  assign n36162 = ~pi38 & ~n64386;
  assign n36163 = ~n36161 & n36162;
  assign n36164 = pi38 & ~n36134;
  assign n36165 = ~n36137 & n36164;
  assign n36166 = ~pi696 & ~n36165;
  assign n36167 = ~n36163 & n36166;
  assign n36168 = ~n36143 & ~n36167;
  assign n36169 = n63888 & ~n36168;
  assign n36170 = ~pi152 & ~n63888;
  assign n36171 = ~pi832 & ~n36170;
  assign n36172 = ~n36169 & n36171;
  assign n36173 = pi696 & n35430;
  assign n36174 = n2923 & ~n36125;
  assign n36175 = ~n36173 & n36174;
  assign n36176 = ~pi152 & ~n2923;
  assign n36177 = pi832 & ~n36176;
  assign n36178 = ~n36175 & n36177;
  assign n36179 = ~n36172 & ~n36178;
  assign n36180 = pi153 & ~n7134;
  assign n36181 = n35576 & ~n36180;
  assign n36182 = pi153 & ~n7118;
  assign n36183 = pi153 & n7129;
  assign n36184 = ~n7124 & n36182;
  assign n36185 = ~n7123 & ~n64389;
  assign n36186 = ~pi153 & ~n6951;
  assign n36187 = n35720 & ~n36186;
  assign n36188 = ~n35657 & n36187;
  assign n36189 = ~pi215 & ~n36188;
  assign n36190 = n36185 & n36189;
  assign n36191 = ~n36181 & ~n36190;
  assign n36192 = pi299 & ~n36191;
  assign n36193 = pi153 & ~n35617;
  assign n36194 = n35594 & ~n36193;
  assign n36195 = ~n36192 & ~n36194;
  assign n36196 = pi766 & ~n36195;
  assign n36197 = n35659 & ~n36186;
  assign n36198 = ~n35580 & ~n36197;
  assign n36199 = n36185 & n36198;
  assign n36200 = ~pi215 & ~n36199;
  assign n36201 = n35606 & ~n36181;
  assign n36202 = ~n35641 & ~n36201;
  assign n36203 = ~n36200 & n36202;
  assign n36204 = pi299 & ~n36203;
  assign n36205 = ~pi153 & ~n7116;
  assign n36206 = n35665 & ~n36205;
  assign n36207 = ~pi766 & ~n36206;
  assign n36208 = ~n36204 & n36207;
  assign n36209 = pi39 & ~n36208;
  assign n36210 = ~n36204 & ~n36206;
  assign n36211 = ~pi766 & ~n36210;
  assign n36212 = pi766 & ~n36192;
  assign n36213 = ~n36194 & n36212;
  assign n36214 = ~n36211 & ~n36213;
  assign n36215 = pi39 & ~n36214;
  assign n36216 = ~n36196 & n36209;
  assign n36217 = ~pi153 & n62781;
  assign n36218 = ~n13676 & ~n35715;
  assign n36219 = ~n36217 & ~n36218;
  assign n36220 = ~n35668 & n36219;
  assign n36221 = ~pi38 & ~n36220;
  assign n36222 = ~n64390 & n36221;
  assign n36223 = pi766 & pi947;
  assign n36224 = n2923 & ~n36223;
  assign n36225 = n7357 & ~n36223;
  assign n36226 = n7356 & n36224;
  assign n36227 = ~n35430 & n64391;
  assign n36228 = pi153 & ~n7357;
  assign n36229 = pi38 & ~n36228;
  assign n36230 = ~n36227 & n36229;
  assign n36231 = pi700 & ~n36230;
  assign n36232 = ~n64390 & ~n36220;
  assign n36233 = ~pi38 & ~n36232;
  assign n36234 = ~pi153 & ~n7357;
  assign n36235 = ~pi766 & pi947;
  assign n36236 = ~pi39 & ~n36235;
  assign n36237 = ~n35430 & ~n36223;
  assign n36238 = n7357 & ~n36237;
  assign n36239 = n35876 & n36236;
  assign n36240 = pi38 & ~n64392;
  assign n36241 = pi38 & ~n36234;
  assign n36242 = ~n64392 & n36241;
  assign n36243 = ~n36234 & n36240;
  assign n36244 = ~n36233 & ~n64393;
  assign n36245 = pi700 & ~n36244;
  assign n36246 = ~n36222 & n36231;
  assign n36247 = n35716 & ~n36205;
  assign n36248 = n36185 & ~n36187;
  assign n36249 = n35690 & n36248;
  assign n36250 = n35692 & ~n36180;
  assign n36251 = ~n35653 & n36181;
  assign n36252 = pi299 & ~n64395;
  assign n36253 = ~n36249 & n36252;
  assign n36254 = pi766 & ~n36253;
  assign n36255 = ~n36247 & n36254;
  assign n36256 = ~pi153 & ~pi766;
  assign n36257 = ~n7143 & n36256;
  assign n36258 = pi39 & ~n36257;
  assign n36259 = ~n36255 & n36258;
  assign n36260 = ~pi38 & ~n36219;
  assign n36261 = ~n36259 & n36260;
  assign n36262 = pi38 & ~n64391;
  assign n36263 = ~n36228 & n36262;
  assign n36264 = ~pi700 & ~n36263;
  assign n36265 = ~n36261 & n36264;
  assign n36266 = n27338 & ~n36265;
  assign n36267 = ~n36261 & ~n36263;
  assign n36268 = ~pi700 & ~n36267;
  assign n36269 = pi700 & ~n64393;
  assign n36270 = ~n36233 & n36269;
  assign n36271 = ~n36268 & ~n36270;
  assign n36272 = n27338 & ~n36271;
  assign n36273 = ~n64394 & n36266;
  assign n36274 = ~pi153 & ~n27338;
  assign n36275 = ~pi57 & ~n36274;
  assign n36276 = ~n64396 & n36275;
  assign n36277 = pi57 & pi153;
  assign n36278 = ~pi832 & ~n36277;
  assign n36279 = ~n36276 & n36278;
  assign n36280 = pi700 & n35430;
  assign n36281 = ~pi700 & ~n36223;
  assign n36282 = ~n36237 & ~n36281;
  assign n36283 = n2923 & ~n36282;
  assign n36284 = n36224 & ~n36280;
  assign n36285 = pi153 & ~n2923;
  assign n36286 = pi832 & ~n36285;
  assign n36287 = ~n64397 & n36286;
  assign n36288 = ~n36279 & ~n36287;
  assign n36289 = ~pi742 & pi947;
  assign n36290 = ~pi704 & n35430;
  assign n36291 = ~n36289 & ~n36290;
  assign n36292 = n2923 & ~n36291;
  assign n36293 = ~pi154 & ~n2923;
  assign n36294 = pi832 & ~n36293;
  assign n36295 = ~n36292 & n36294;
  assign n36296 = ~pi154 & n62781;
  assign n36297 = n35669 & ~n36296;
  assign n36298 = ~n35601 & n36297;
  assign n36299 = ~pi154 & ~n64356;
  assign n36300 = pi154 & ~n64361;
  assign n36301 = pi39 & ~n36300;
  assign n36302 = ~n36299 & n36301;
  assign n36303 = ~n36298 & ~n36302;
  assign n36304 = ~pi38 & ~n36303;
  assign n36305 = ~pi154 & ~n7357;
  assign n36306 = n35636 & ~n36305;
  assign n36307 = ~pi742 & ~n36306;
  assign n36308 = ~n36304 & n36307;
  assign n36309 = ~pi154 & n35647;
  assign n36310 = pi154 & n35666;
  assign n36311 = pi39 & ~n36310;
  assign n36312 = ~n36309 & n36311;
  assign n36313 = ~n36297 & ~n36312;
  assign n36314 = ~pi38 & ~n36313;
  assign n36315 = n35676 & ~n36305;
  assign n36316 = pi742 & ~n36315;
  assign n36317 = ~n36314 & n36316;
  assign n36318 = ~pi704 & ~n36317;
  assign n36319 = ~pi704 & ~n36308;
  assign n36320 = ~n36317 & n36319;
  assign n36321 = ~n36308 & n36318;
  assign n36322 = n35715 & ~n36296;
  assign n36323 = ~pi154 & ~n35696;
  assign n36324 = pi154 & n35724;
  assign n36325 = pi39 & ~n36324;
  assign n36326 = ~n36323 & n36325;
  assign n36327 = ~n36322 & ~n36326;
  assign n36328 = ~pi38 & ~n36327;
  assign n36329 = ~n35713 & ~n36305;
  assign n36330 = ~pi742 & ~n36329;
  assign n36331 = ~n36328 & n36330;
  assign n36332 = ~pi154 & pi742;
  assign n36333 = ~n8091 & n36332;
  assign n36334 = pi704 & ~n36333;
  assign n36335 = ~n36331 & n36334;
  assign n36336 = n63888 & ~n36335;
  assign n36337 = ~n64398 & n36336;
  assign n36338 = ~pi154 & ~n63888;
  assign n36339 = ~pi832 & ~n36338;
  assign n36340 = ~n36337 & n36339;
  assign po311 = ~n36295 & ~n36340;
  assign n36342 = ~pi38 & ~n35670;
  assign n36343 = ~n35676 & ~n36342;
  assign n36344 = pi757 & n36343;
  assign n36345 = ~pi38 & ~n35629;
  assign n36346 = ~n35636 & ~n36345;
  assign n36347 = ~pi757 & n36346;
  assign n36348 = ~pi686 & ~n36347;
  assign n36349 = ~pi686 & ~n36344;
  assign n36350 = ~n36347 & n36349;
  assign n36351 = ~n36344 & n36348;
  assign n36352 = ~pi757 & n35728;
  assign n36353 = pi686 & ~n36352;
  assign n36354 = n63888 & ~n36353;
  assign n36355 = ~n64399 & n36354;
  assign n36356 = pi155 & ~n36355;
  assign n36357 = ~pi757 & n35706;
  assign n36358 = pi686 & ~n14957;
  assign n36359 = ~pi757 & ~n35706;
  assign n36360 = ~n14951 & ~n36359;
  assign n36361 = pi686 & ~n36360;
  assign n36362 = ~n36357 & n36358;
  assign n36363 = ~pi38 & ~n35651;
  assign n36364 = n10335 & ~n35430;
  assign n36365 = pi38 & ~n35430;
  assign n36366 = n7357 & n36365;
  assign n36367 = n10335 & n36133;
  assign n36368 = n7357 & n35676;
  assign n36369 = n6955 & n36364;
  assign n36370 = ~n36363 & ~n64401;
  assign n36371 = pi757 & n36370;
  assign n36372 = ~pi38 & ~n35604;
  assign n36373 = pi38 & n35633;
  assign n36374 = ~n36372 & ~n36373;
  assign n36375 = ~pi757 & n36374;
  assign n36376 = ~pi686 & ~n36375;
  assign n36377 = ~pi686 & ~n36371;
  assign n36378 = ~n36375 & n36377;
  assign n36379 = ~n36371 & n36376;
  assign n36380 = ~n64400 & ~n64402;
  assign n36381 = ~pi155 & n63888;
  assign n36382 = ~n36380 & n36381;
  assign n36383 = ~n36356 & ~n36382;
  assign n36384 = ~pi832 & ~n36383;
  assign n36385 = ~pi757 & pi947;
  assign n36386 = ~pi686 & n35430;
  assign n36387 = ~n36385 & ~n36386;
  assign n36388 = n2923 & ~n36387;
  assign n36389 = ~pi155 & ~n2923;
  assign n36390 = pi832 & ~n36389;
  assign n36391 = ~n36388 & n36390;
  assign po312 = ~n36384 & ~n36391;
  assign n36393 = ~pi741 & pi947;
  assign n36394 = ~pi724 & n35430;
  assign n36395 = ~n36393 & ~n36394;
  assign n36396 = n2923 & ~n36395;
  assign n36397 = ~pi156 & ~n2923;
  assign n36398 = pi832 & ~n36397;
  assign n36399 = ~n36396 & n36398;
  assign n36400 = pi741 & ~n36370;
  assign n36401 = ~pi741 & ~n36374;
  assign n36402 = ~pi724 & ~n36401;
  assign n36403 = ~pi724 & ~n36400;
  assign n36404 = ~n36401 & n36403;
  assign n36405 = ~n36400 & n36402;
  assign n36406 = ~pi741 & ~n35706;
  assign n36407 = pi724 & ~n16107;
  assign n36408 = ~n36406 & n36407;
  assign n36409 = n63888 & ~n36408;
  assign n36410 = ~n64403 & n36409;
  assign n36411 = ~pi156 & ~n36410;
  assign n36412 = pi741 & ~n36343;
  assign n36413 = ~pi741 & ~n36346;
  assign n36414 = ~pi724 & ~n36413;
  assign n36415 = ~pi724 & ~n36412;
  assign n36416 = ~n36413 & n36415;
  assign n36417 = ~n36412 & n36414;
  assign n36418 = pi724 & ~pi741;
  assign n36419 = n35728 & n36418;
  assign n36420 = ~n64404 & ~n36419;
  assign n36421 = pi156 & n63888;
  assign n36422 = ~n36420 & n36421;
  assign n36423 = ~pi832 & ~n36422;
  assign n36424 = ~n36411 & n36423;
  assign po313 = ~n36399 & ~n36424;
  assign n36426 = pi760 & ~n35647;
  assign n36427 = ~pi760 & n64356;
  assign n36428 = ~pi157 & ~n36427;
  assign n36429 = ~pi157 & ~n36426;
  assign n36430 = ~n36427 & n36429;
  assign n36431 = ~n36426 & n36428;
  assign n36432 = ~pi760 & n64361;
  assign n36433 = pi760 & ~n35666;
  assign n36434 = pi157 & ~n36433;
  assign n36435 = pi157 & ~n36432;
  assign n36436 = ~n36433 & n36435;
  assign n36437 = ~n36432 & n36434;
  assign n36438 = pi39 & ~n64406;
  assign n36439 = pi760 & n35666;
  assign n36440 = ~pi760 & ~n64361;
  assign n36441 = pi157 & ~n36440;
  assign n36442 = ~n36439 & n36441;
  assign n36443 = ~pi760 & ~n64356;
  assign n36444 = pi760 & n35647;
  assign n36445 = ~pi157 & ~n36444;
  assign n36446 = ~n36443 & n36445;
  assign n36447 = ~n36442 & ~n36446;
  assign n36448 = pi39 & ~n36447;
  assign n36449 = ~n64405 & n36438;
  assign n36450 = ~pi760 & pi947;
  assign n36451 = ~n62781 & n36450;
  assign n36452 = ~pi157 & n62781;
  assign n36453 = ~pi39 & ~n36452;
  assign n36454 = ~pi39 & ~n36451;
  assign n36455 = ~n36452 & n36454;
  assign n36456 = ~n36451 & n36453;
  assign n36457 = ~n35668 & n64408;
  assign n36458 = ~pi38 & ~n36457;
  assign n36459 = ~n64407 & n36458;
  assign n36460 = n7357 & ~n36450;
  assign n36461 = ~n35430 & n36460;
  assign n36462 = pi157 & ~n7357;
  assign n36463 = pi38 & ~n36462;
  assign n36464 = ~n36461 & n36463;
  assign n36465 = ~pi688 & ~n36464;
  assign n36466 = ~n36459 & n36465;
  assign n36467 = ~pi157 & ~n35693;
  assign n36468 = ~n33133 & ~n35723;
  assign n36469 = ~n36467 & ~n36468;
  assign n36470 = ~pi157 & ~n7116;
  assign n36471 = n35716 & ~n36470;
  assign n36472 = ~pi760 & ~n36471;
  assign n36473 = ~n36469 & n36472;
  assign n36474 = ~pi157 & pi760;
  assign n36475 = ~n7143 & n36474;
  assign n36476 = pi39 & ~n36475;
  assign n36477 = ~n36473 & n36476;
  assign n36478 = ~pi38 & ~n64408;
  assign n36479 = ~n36477 & n36478;
  assign n36480 = pi38 & ~n36460;
  assign n36481 = ~n36462 & n36480;
  assign n36482 = pi688 & ~n36481;
  assign n36483 = ~n36479 & n36482;
  assign n36484 = n63888 & ~n36483;
  assign n36485 = ~n36479 & ~n36481;
  assign n36486 = pi688 & ~n36485;
  assign n36487 = ~n64407 & ~n36457;
  assign n36488 = ~pi38 & ~n36487;
  assign n36489 = ~pi157 & ~n7357;
  assign n36490 = pi760 & pi947;
  assign n36491 = ~pi39 & ~n36490;
  assign n36492 = ~n35430 & ~n36450;
  assign n36493 = n7357 & ~n36492;
  assign n36494 = n35876 & n36491;
  assign n36495 = pi38 & ~n64409;
  assign n36496 = pi38 & ~n36489;
  assign n36497 = ~n64409 & n36496;
  assign n36498 = ~n36489 & n36495;
  assign n36499 = ~pi688 & ~n64410;
  assign n36500 = ~n36488 & n36499;
  assign n36501 = ~n36486 & ~n36500;
  assign n36502 = n63888 & ~n36501;
  assign n36503 = ~n36466 & n36484;
  assign n36504 = ~pi157 & ~n63888;
  assign n36505 = ~pi832 & ~n36504;
  assign n36506 = ~n64411 & n36505;
  assign n36507 = ~pi688 & n35430;
  assign n36508 = ~n36450 & ~n36507;
  assign n36509 = n2923 & ~n36508;
  assign n36510 = ~pi157 & ~n2923;
  assign n36511 = pi832 & ~n36510;
  assign n36512 = ~n36509 & n36511;
  assign po314 = ~n36506 & ~n36512;
  assign n36514 = ~pi753 & pi947;
  assign n36515 = ~pi702 & n35430;
  assign n36516 = ~n36514 & ~n36515;
  assign n36517 = pi702 & ~n36514;
  assign n36518 = ~n35430 & ~n36514;
  assign n36519 = n2923 & ~n36518;
  assign n36520 = ~n36517 & n36519;
  assign n36521 = n2923 & ~n36516;
  assign n36522 = ~pi158 & ~n2923;
  assign n36523 = pi832 & ~n36522;
  assign n36524 = ~n64412 & n36523;
  assign n36525 = ~pi158 & ~n64356;
  assign n36526 = pi158 & ~n64361;
  assign n36527 = ~pi753 & ~n36526;
  assign n36528 = ~n36525 & n36527;
  assign n36529 = ~pi158 & n35647;
  assign n36530 = pi158 & n35666;
  assign n36531 = pi753 & ~n36530;
  assign n36532 = ~n36529 & n36531;
  assign n36533 = pi39 & ~n36532;
  assign n36534 = ~pi158 & ~n35647;
  assign n36535 = pi158 & ~n35666;
  assign n36536 = pi753 & ~n36535;
  assign n36537 = ~n36534 & n36536;
  assign n36538 = ~pi158 & n64356;
  assign n36539 = pi158 & n64361;
  assign n36540 = ~pi753 & ~n36539;
  assign n36541 = ~n36538 & n36540;
  assign n36542 = ~n36537 & ~n36541;
  assign n36543 = pi39 & ~n36542;
  assign n36544 = ~n36528 & n36533;
  assign n36545 = n35649 & ~n36514;
  assign n36546 = pi158 & n62781;
  assign n36547 = ~pi39 & ~n36546;
  assign n36548 = ~n36545 & n36547;
  assign n36549 = ~pi38 & ~n36548;
  assign n36550 = ~n64413 & n36549;
  assign n36551 = ~pi158 & ~n7357;
  assign n36552 = pi753 & pi947;
  assign n36553 = ~pi39 & ~n36552;
  assign n36554 = n35876 & n36553;
  assign n36555 = n7357 & ~n36518;
  assign n36556 = n7356 & n36519;
  assign n36557 = pi38 & ~n64414;
  assign n36558 = pi158 & ~n7357;
  assign n36559 = n7357 & ~n36514;
  assign n36560 = ~n35430 & n36559;
  assign n36561 = ~n36558 & ~n36560;
  assign n36562 = pi38 & ~n36561;
  assign n36563 = pi38 & ~n36551;
  assign n36564 = ~n64414 & n36563;
  assign n36565 = ~n36551 & n36557;
  assign n36566 = ~pi702 & ~n64415;
  assign n36567 = ~n36550 & n36566;
  assign n36568 = ~pi158 & n35696;
  assign n36569 = pi158 & ~n35724;
  assign n36570 = ~pi753 & ~n36569;
  assign n36571 = ~n36568 & n36570;
  assign n36572 = ~pi158 & pi753;
  assign n36573 = ~n7143 & n36572;
  assign n36574 = ~n36571 & ~n36573;
  assign n36575 = pi39 & ~n36574;
  assign n36576 = ~n16863 & ~n36546;
  assign n36577 = n35699 & n36576;
  assign n36578 = ~pi38 & ~n36577;
  assign n36579 = ~n36575 & n36578;
  assign n36580 = ~n36558 & ~n36559;
  assign n36581 = pi38 & ~n36580;
  assign n36582 = pi702 & ~n36581;
  assign n36583 = ~n36579 & n36582;
  assign n36584 = ~n36567 & ~n36583;
  assign n36585 = n63888 & ~n36584;
  assign n36586 = ~pi158 & ~n63888;
  assign n36587 = ~pi832 & ~n36586;
  assign n36588 = ~n36585 & n36587;
  assign po315 = ~n36524 & ~n36588;
  assign n36590 = ~pi754 & pi947;
  assign n36591 = ~pi709 & n35430;
  assign n36592 = ~n36590 & ~n36591;
  assign n36593 = pi709 & ~n36590;
  assign n36594 = ~n35430 & ~n36590;
  assign n36595 = n2923 & ~n36594;
  assign n36596 = ~n36593 & n36595;
  assign n36597 = n2923 & ~n36592;
  assign n36598 = ~pi159 & ~n2923;
  assign n36599 = pi832 & ~n36598;
  assign n36600 = ~n64416 & n36599;
  assign n36601 = ~pi159 & ~n64356;
  assign n36602 = pi159 & ~n64361;
  assign n36603 = ~pi754 & ~n36602;
  assign n36604 = ~n36601 & n36603;
  assign n36605 = ~pi159 & n35647;
  assign n36606 = pi159 & n35666;
  assign n36607 = pi754 & ~n36606;
  assign n36608 = ~n36605 & n36607;
  assign n36609 = pi39 & ~n36608;
  assign n36610 = ~pi159 & ~n35647;
  assign n36611 = pi159 & ~n35666;
  assign n36612 = pi754 & ~n36611;
  assign n36613 = ~n36610 & n36612;
  assign n36614 = ~pi159 & n64356;
  assign n36615 = pi159 & n64361;
  assign n36616 = ~pi754 & ~n36615;
  assign n36617 = ~n36614 & n36616;
  assign n36618 = ~n36613 & ~n36617;
  assign n36619 = pi39 & ~n36618;
  assign n36620 = ~n36604 & n36609;
  assign n36621 = n35649 & ~n36590;
  assign n36622 = pi159 & n62781;
  assign n36623 = ~pi39 & ~n36622;
  assign n36624 = ~n36621 & n36623;
  assign n36625 = ~pi38 & ~n36624;
  assign n36626 = ~n64417 & n36625;
  assign n36627 = ~pi159 & ~n7357;
  assign n36628 = pi754 & pi947;
  assign n36629 = ~pi39 & ~n36628;
  assign n36630 = n35876 & n36629;
  assign n36631 = n7357 & ~n36594;
  assign n36632 = n7356 & n36595;
  assign n36633 = pi38 & ~n64418;
  assign n36634 = pi159 & ~n7357;
  assign n36635 = n7357 & ~n36590;
  assign n36636 = ~n35430 & n36635;
  assign n36637 = ~n36634 & ~n36636;
  assign n36638 = pi38 & ~n36637;
  assign n36639 = pi38 & ~n36627;
  assign n36640 = ~n64418 & n36639;
  assign n36641 = ~n36627 & n36633;
  assign n36642 = ~pi709 & ~n64419;
  assign n36643 = ~n36626 & n36642;
  assign n36644 = ~pi159 & n35696;
  assign n36645 = pi159 & ~n35724;
  assign n36646 = ~pi754 & ~n36645;
  assign n36647 = ~n36644 & n36646;
  assign n36648 = ~pi159 & pi754;
  assign n36649 = ~n7143 & n36648;
  assign n36650 = ~n36647 & ~n36649;
  assign n36651 = pi39 & ~n36650;
  assign n36652 = ~n17458 & ~n36622;
  assign n36653 = n35699 & n36652;
  assign n36654 = ~pi38 & ~n36653;
  assign n36655 = ~n36651 & n36654;
  assign n36656 = ~n36634 & ~n36635;
  assign n36657 = pi38 & ~n36656;
  assign n36658 = pi709 & ~n36657;
  assign n36659 = ~n36655 & n36658;
  assign n36660 = ~n36643 & ~n36659;
  assign n36661 = n63888 & ~n36660;
  assign n36662 = ~pi159 & ~n63888;
  assign n36663 = ~pi832 & ~n36662;
  assign n36664 = ~n36661 & n36663;
  assign po316 = ~n36600 & ~n36664;
  assign n36666 = ~pi756 & pi947;
  assign n36667 = ~pi734 & n35430;
  assign n36668 = ~n36666 & ~n36667;
  assign n36669 = n2923 & ~n36668;
  assign n36670 = ~pi160 & ~n2923;
  assign n36671 = pi832 & ~n36670;
  assign n36672 = ~n36669 & n36671;
  assign n36673 = ~pi160 & n64356;
  assign n36674 = pi160 & n64361;
  assign n36675 = ~pi756 & ~n36674;
  assign n36676 = ~n36673 & n36675;
  assign n36677 = ~pi160 & n35643;
  assign n36678 = pi160 & ~n35753;
  assign n36679 = pi756 & ~n64362;
  assign n36680 = ~n36678 & n36679;
  assign n36681 = ~n36677 & n36680;
  assign n36682 = pi39 & ~n36681;
  assign n36683 = ~n64362 & ~n36678;
  assign n36684 = ~n36677 & n36683;
  assign n36685 = pi756 & ~n36684;
  assign n36686 = ~pi160 & ~n64356;
  assign n36687 = pi160 & ~n64361;
  assign n36688 = ~pi756 & ~n36687;
  assign n36689 = ~n36686 & n36688;
  assign n36690 = ~n36685 & ~n36689;
  assign n36691 = pi39 & ~n36690;
  assign n36692 = ~n36676 & n36682;
  assign n36693 = ~n62781 & n36666;
  assign n36694 = ~pi160 & n62781;
  assign n36695 = ~pi39 & ~n36694;
  assign n36696 = ~pi39 & ~n36693;
  assign n36697 = ~n36694 & n36696;
  assign n36698 = ~n36693 & n36695;
  assign n36699 = ~n35668 & n64421;
  assign n36700 = ~pi38 & ~n36699;
  assign n36701 = ~n64420 & n36700;
  assign n36702 = n7357 & ~n36666;
  assign n36703 = ~n35430 & n36702;
  assign n36704 = pi160 & ~n7357;
  assign n36705 = pi38 & ~n36704;
  assign n36706 = ~n36703 & n36705;
  assign n36707 = ~pi734 & ~n36706;
  assign n36708 = ~n36701 & n36707;
  assign n36709 = ~pi160 & ~n35693;
  assign n36710 = pi160 & ~n35783;
  assign n36711 = pi299 & ~n36710;
  assign n36712 = ~n36709 & n36711;
  assign n36713 = ~pi160 & ~n7116;
  assign n36714 = n35716 & ~n36713;
  assign n36715 = ~pi756 & ~n36714;
  assign n36716 = ~n36712 & n36715;
  assign n36717 = ~pi160 & pi756;
  assign n36718 = ~n7143 & n36717;
  assign n36719 = pi39 & ~n36718;
  assign n36720 = ~n36716 & n36719;
  assign n36721 = ~pi38 & ~n64421;
  assign n36722 = ~n36720 & n36721;
  assign n36723 = pi38 & ~n36702;
  assign n36724 = ~n36704 & n36723;
  assign n36725 = pi734 & ~n36724;
  assign n36726 = ~n36722 & n36725;
  assign n36727 = n63888 & ~n36726;
  assign n36728 = ~n36722 & ~n36724;
  assign n36729 = pi734 & ~n36728;
  assign n36730 = ~n64420 & ~n36699;
  assign n36731 = ~pi38 & ~n36730;
  assign n36732 = ~pi160 & ~n7357;
  assign n36733 = pi756 & pi947;
  assign n36734 = ~pi39 & ~n36733;
  assign n36735 = ~n35430 & ~n36666;
  assign n36736 = n7357 & ~n36735;
  assign n36737 = n35876 & n36734;
  assign n36738 = pi38 & ~n64422;
  assign n36739 = pi38 & ~n36732;
  assign n36740 = ~n64422 & n36739;
  assign n36741 = ~n36732 & n36738;
  assign n36742 = ~pi734 & ~n64423;
  assign n36743 = ~n36731 & n36742;
  assign n36744 = ~n36729 & ~n36743;
  assign n36745 = n63888 & ~n36744;
  assign n36746 = ~n36708 & n36727;
  assign n36747 = ~pi160 & ~n63888;
  assign n36748 = ~pi832 & ~n36747;
  assign n36749 = ~n64424 & n36748;
  assign po317 = ~n36672 & ~n36749;
  assign n36751 = ~pi161 & ~n62789;
  assign n36752 = n36072 & ~n36751;
  assign n36753 = n36075 & ~n36752;
  assign n36754 = pi161 & ~n6951;
  assign n36755 = ~n35607 & ~n36754;
  assign n36756 = n7034 & n36755;
  assign n36757 = ~pi223 & ~n36756;
  assign n36758 = ~n36753 & n36757;
  assign n36759 = ~pi161 & n62785;
  assign n36760 = n35591 & ~n36759;
  assign n36761 = ~pi299 & ~n36760;
  assign n36762 = n35589 & ~n36759;
  assign n36763 = ~pi299 & ~n36762;
  assign n36764 = ~n36760 & n36763;
  assign n36765 = n36761 & ~n36762;
  assign n36766 = ~n36758 & n64425;
  assign n36767 = n7118 & n36755;
  assign n36768 = ~pi215 & ~n36767;
  assign n36769 = pi161 & n35579;
  assign n36770 = n35656 & ~n36769;
  assign n36771 = ~n7124 & n36770;
  assign n36772 = n36768 & ~n36771;
  assign n36773 = ~pi161 & ~n7134;
  assign n36774 = n35576 & ~n36773;
  assign n36775 = pi299 & ~n36774;
  assign n36776 = ~n36772 & n36775;
  assign n36777 = pi758 & ~n36776;
  assign n36778 = pi758 & ~n36766;
  assign n36779 = ~n36776 & n36778;
  assign n36780 = ~n36766 & n36777;
  assign n36781 = ~n35658 & ~n36754;
  assign n36782 = n7034 & ~n36781;
  assign n36783 = n36107 & ~n36751;
  assign n36784 = ~n36782 & ~n36783;
  assign n36785 = ~pi223 & ~n36784;
  assign n36786 = n36761 & ~n36785;
  assign n36787 = ~n35577 & n36768;
  assign n36788 = ~n36770 & n36787;
  assign n36789 = ~n36114 & n36774;
  assign n36790 = pi299 & ~n36789;
  assign n36791 = ~n36788 & n36790;
  assign n36792 = ~pi758 & ~n36791;
  assign n36793 = ~n36786 & n36792;
  assign n36794 = pi39 & ~n36793;
  assign n36795 = ~n64426 & n36794;
  assign n36796 = pi758 & pi947;
  assign n36797 = ~n62781 & n36796;
  assign n36798 = pi161 & n62781;
  assign n36799 = ~pi39 & ~n36798;
  assign n36800 = ~pi39 & ~n36797;
  assign n36801 = ~n36798 & n36800;
  assign n36802 = ~n36797 & n36799;
  assign n36803 = ~n35668 & n64427;
  assign n36804 = ~pi38 & ~n36803;
  assign n36805 = ~n36795 & n36804;
  assign n36806 = ~pi39 & ~n36796;
  assign n36807 = n7357 & ~n36796;
  assign n36808 = ~n35430 & n36807;
  assign n36809 = n36133 & n36806;
  assign n36810 = ~pi161 & ~n7357;
  assign n36811 = pi38 & ~n36810;
  assign n36812 = pi38 & ~n64428;
  assign n36813 = ~n36810 & n36812;
  assign n36814 = ~n64428 & n36811;
  assign n36815 = pi736 & ~n64429;
  assign n36816 = ~n36805 & n36815;
  assign n36817 = ~n35689 & ~n36770;
  assign n36818 = ~n35578 & ~n36817;
  assign n36819 = ~n35719 & ~n36754;
  assign n36820 = n7118 & n36819;
  assign n36821 = ~pi215 & ~n36820;
  assign n36822 = ~n36818 & n36821;
  assign n36823 = pi161 & n35692;
  assign n36824 = n35717 & ~n36823;
  assign n36825 = ~n36822 & n36824;
  assign n36826 = n7034 & ~n36819;
  assign n36827 = ~n36752 & ~n36826;
  assign n36828 = ~pi223 & ~n36827;
  assign n36829 = n36763 & ~n36828;
  assign n36830 = pi758 & ~n36829;
  assign n36831 = ~n36825 & n36830;
  assign n36832 = pi161 & n10925;
  assign n36833 = pi39 & ~n36832;
  assign n36834 = ~n36831 & n36833;
  assign n36835 = ~pi38 & ~n64427;
  assign n36836 = ~n36834 & n36835;
  assign n36837 = pi38 & ~n36807;
  assign n36838 = ~n36810 & n36837;
  assign n36839 = ~pi736 & ~n36838;
  assign n36840 = ~n36836 & n36839;
  assign n36841 = ~n36816 & ~n36840;
  assign n36842 = n63888 & ~n36841;
  assign n36843 = ~pi161 & ~n63888;
  assign n36844 = ~pi832 & ~n36843;
  assign n36845 = ~n36842 & n36844;
  assign n36846 = pi736 & n35430;
  assign n36847 = n2923 & ~n36796;
  assign n36848 = ~n36846 & n36847;
  assign n36849 = ~pi161 & ~n2923;
  assign n36850 = pi832 & ~n36849;
  assign n36851 = ~n36848 & n36850;
  assign n36852 = ~n36845 & ~n36851;
  assign n36853 = ~pi761 & pi947;
  assign n36854 = ~pi738 & n35430;
  assign n36855 = ~n36853 & ~n36854;
  assign n36856 = pi738 & ~n36853;
  assign n36857 = ~n35430 & ~n36853;
  assign n36858 = n2923 & ~n36857;
  assign n36859 = ~n36856 & n36858;
  assign n36860 = n2923 & ~n36855;
  assign n36861 = ~pi162 & ~n2923;
  assign n36862 = pi832 & ~n36861;
  assign n36863 = ~n64430 & n36862;
  assign n36864 = ~pi162 & n64356;
  assign n36865 = pi162 & n64361;
  assign n36866 = ~pi761 & ~n36865;
  assign n36867 = ~n36864 & n36866;
  assign n36868 = pi162 & pi299;
  assign n36869 = ~n35647 & ~n36868;
  assign n36870 = pi162 & ~n35753;
  assign n36871 = pi761 & ~n36870;
  assign n36872 = ~n36869 & n36871;
  assign n36873 = pi39 & ~n36872;
  assign n36874 = ~n36869 & ~n36870;
  assign n36875 = pi761 & ~n36874;
  assign n36876 = ~pi162 & ~n64356;
  assign n36877 = pi162 & ~n64361;
  assign n36878 = ~pi761 & ~n36877;
  assign n36879 = ~n36876 & n36878;
  assign n36880 = ~n36875 & ~n36879;
  assign n36881 = pi39 & ~n36880;
  assign n36882 = pi39 & ~n36867;
  assign n36883 = ~n36872 & n36882;
  assign n36884 = ~n36867 & n36873;
  assign n36885 = ~n62781 & n36853;
  assign n36886 = ~pi162 & n62781;
  assign n36887 = ~pi39 & ~n36886;
  assign n36888 = ~pi39 & ~n36885;
  assign n36889 = ~n36886 & n36888;
  assign n36890 = ~n36885 & n36887;
  assign n36891 = ~n35668 & n64432;
  assign n36892 = ~pi38 & ~n36891;
  assign n36893 = ~n64431 & n36892;
  assign n36894 = n7357 & ~n36853;
  assign n36895 = ~n35430 & n36894;
  assign n36896 = pi162 & ~n7357;
  assign n36897 = pi38 & ~n36896;
  assign n36898 = ~n36895 & n36897;
  assign n36899 = ~pi738 & ~n36898;
  assign n36900 = ~n36893 & n36899;
  assign n36901 = ~pi761 & n35695;
  assign n36902 = pi761 & n7143;
  assign n36903 = ~pi162 & ~n36902;
  assign n36904 = ~n36901 & n36903;
  assign n36905 = ~n35783 & n36868;
  assign n36906 = ~n64364 & ~n36905;
  assign n36907 = ~pi761 & ~n36906;
  assign n36908 = pi39 & ~n36907;
  assign n36909 = ~pi162 & ~n7143;
  assign n36910 = pi761 & ~n36909;
  assign n36911 = ~pi162 & ~n36901;
  assign n36912 = n36906 & ~n36911;
  assign n36913 = ~n36910 & ~n36912;
  assign n36914 = pi39 & ~n36913;
  assign n36915 = ~n36904 & n36908;
  assign n36916 = ~pi38 & ~n64432;
  assign n36917 = ~n64433 & n36916;
  assign n36918 = pi38 & ~n36894;
  assign n36919 = ~n36896 & n36918;
  assign n36920 = pi738 & ~n36919;
  assign n36921 = ~n36917 & n36920;
  assign n36922 = n63888 & ~n36921;
  assign n36923 = ~n36917 & ~n36919;
  assign n36924 = pi738 & ~n36923;
  assign n36925 = ~n64431 & ~n36891;
  assign n36926 = ~pi38 & ~n36925;
  assign n36927 = ~pi162 & ~n7357;
  assign n36928 = pi761 & pi947;
  assign n36929 = ~pi39 & ~n36928;
  assign n36930 = n35876 & n36929;
  assign n36931 = n7357 & ~n36857;
  assign n36932 = n7356 & n36858;
  assign n36933 = pi38 & ~n64434;
  assign n36934 = pi38 & ~n36927;
  assign n36935 = ~n64434 & n36934;
  assign n36936 = ~n36927 & n36933;
  assign n36937 = ~pi738 & ~n64435;
  assign n36938 = ~n36926 & n36937;
  assign n36939 = ~n36924 & ~n36938;
  assign n36940 = n63888 & ~n36939;
  assign n36941 = ~n36900 & n36922;
  assign n36942 = ~pi162 & ~n63888;
  assign n36943 = ~pi832 & ~n36942;
  assign n36944 = ~n64436 & n36943;
  assign po319 = ~n36863 & ~n36944;
  assign n36946 = ~pi163 & n64356;
  assign n36947 = pi163 & n64361;
  assign n36948 = ~pi777 & ~n36947;
  assign n36949 = ~n36946 & n36948;
  assign n36950 = ~pi163 & n35643;
  assign n36951 = pi163 & ~n35753;
  assign n36952 = pi777 & ~n64362;
  assign n36953 = ~n36951 & n36952;
  assign n36954 = ~n36950 & n36953;
  assign n36955 = pi39 & ~n36954;
  assign n36956 = ~n64362 & ~n36951;
  assign n36957 = ~n36950 & n36956;
  assign n36958 = pi777 & ~n36957;
  assign n36959 = ~pi163 & ~n64356;
  assign n36960 = pi163 & ~n64361;
  assign n36961 = ~pi777 & ~n36960;
  assign n36962 = ~n36959 & n36961;
  assign n36963 = ~n36958 & ~n36962;
  assign n36964 = pi39 & ~n36963;
  assign n36965 = ~n36949 & n36955;
  assign n36966 = ~pi777 & pi947;
  assign n36967 = ~n62781 & n36966;
  assign n36968 = ~pi163 & n62781;
  assign n36969 = ~pi39 & ~n36968;
  assign n36970 = ~pi39 & ~n36967;
  assign n36971 = ~n36968 & n36970;
  assign n36972 = ~n36967 & n36969;
  assign n36973 = ~n35668 & n64438;
  assign n36974 = ~pi38 & ~n36973;
  assign n36975 = ~n64437 & n36974;
  assign n36976 = n7357 & ~n36966;
  assign n36977 = ~n35430 & n36976;
  assign n36978 = pi163 & ~n7357;
  assign n36979 = pi38 & ~n36978;
  assign n36980 = ~n36977 & n36979;
  assign n36981 = ~pi737 & ~n36980;
  assign n36982 = ~n36975 & n36981;
  assign n36983 = ~pi163 & ~n35693;
  assign n36984 = ~pi163 & pi299;
  assign n36985 = ~n35723 & ~n36984;
  assign n36986 = ~n36983 & ~n36985;
  assign n36987 = ~pi163 & ~n7116;
  assign n36988 = n35716 & ~n36987;
  assign n36989 = ~pi777 & ~n36988;
  assign n36990 = ~n36986 & n36989;
  assign n36991 = ~pi163 & pi777;
  assign n36992 = ~n7143 & n36991;
  assign n36993 = pi39 & ~n36992;
  assign n36994 = ~n36990 & n36993;
  assign n36995 = ~pi38 & ~n64438;
  assign n36996 = ~n36994 & n36995;
  assign n36997 = pi38 & ~n36976;
  assign n36998 = ~n36978 & n36997;
  assign n36999 = pi737 & ~n36998;
  assign n37000 = ~n36996 & n36999;
  assign n37001 = n63888 & ~n37000;
  assign n37002 = ~n36996 & ~n36998;
  assign n37003 = pi737 & ~n37002;
  assign n37004 = ~n64437 & ~n36973;
  assign n37005 = ~pi38 & ~n37004;
  assign n37006 = ~pi163 & ~n7357;
  assign n37007 = pi777 & pi947;
  assign n37008 = ~pi39 & ~n37007;
  assign n37009 = ~n35430 & ~n36966;
  assign n37010 = n7357 & ~n37009;
  assign n37011 = n35876 & n37008;
  assign n37012 = pi38 & ~n64439;
  assign n37013 = pi38 & ~n37006;
  assign n37014 = ~n64439 & n37013;
  assign n37015 = ~n37006 & n37012;
  assign n37016 = ~pi737 & ~n64440;
  assign n37017 = ~n37005 & n37016;
  assign n37018 = ~n37003 & ~n37017;
  assign n37019 = n63888 & ~n37018;
  assign n37020 = ~n36982 & n37001;
  assign n37021 = ~pi163 & ~n63888;
  assign n37022 = ~pi832 & ~n37021;
  assign n37023 = ~n64441 & n37022;
  assign n37024 = ~pi737 & n35430;
  assign n37025 = ~n36966 & ~n37024;
  assign n37026 = n2923 & ~n37025;
  assign n37027 = ~pi163 & ~n2923;
  assign n37028 = pi832 & ~n37027;
  assign n37029 = ~n37026 & n37028;
  assign po320 = ~n37023 & ~n37029;
  assign n37031 = ~pi752 & pi947;
  assign n37032 = pi703 & n35430;
  assign n37033 = ~n37031 & ~n37032;
  assign n37034 = n2923 & ~n37033;
  assign n37035 = ~pi164 & ~n2923;
  assign n37036 = pi832 & ~n37035;
  assign n37037 = ~n37034 & n37036;
  assign n37038 = ~pi164 & n35604;
  assign n37039 = pi164 & n35629;
  assign n37040 = ~pi38 & ~n37039;
  assign n37041 = ~n37038 & n37040;
  assign n37042 = ~pi164 & ~n35633;
  assign n37043 = n35636 & ~n37042;
  assign n37044 = ~pi752 & ~n37043;
  assign n37045 = ~n37041 & n37044;
  assign n37046 = ~pi164 & n35651;
  assign n37047 = pi164 & n35670;
  assign n37048 = ~pi38 & ~n37047;
  assign n37049 = ~n37046 & n37048;
  assign n37050 = ~pi164 & ~n7357;
  assign n37051 = n35676 & ~n37050;
  assign n37052 = pi752 & ~n37051;
  assign n37053 = ~n37049 & n37052;
  assign n37054 = ~n37045 & ~n37053;
  assign n37055 = pi703 & ~n37054;
  assign n37056 = pi164 & ~n35705;
  assign n37057 = ~pi752 & ~n37056;
  assign n37058 = ~n35706 & n37057;
  assign n37059 = ~pi164 & ~n8091;
  assign n37060 = pi752 & ~n37059;
  assign n37061 = pi164 & ~n35728;
  assign n37062 = ~pi703 & ~n37061;
  assign n37063 = ~pi752 & n35728;
  assign n37064 = pi164 & ~n37063;
  assign n37065 = pi752 & n8091;
  assign n37066 = ~pi703 & ~n37065;
  assign n37067 = ~n37064 & n37066;
  assign n37068 = ~n37060 & n37062;
  assign n37069 = ~n37058 & n64442;
  assign n37070 = ~n37055 & ~n37069;
  assign n37071 = n63888 & ~n37070;
  assign n37072 = ~pi164 & ~n63888;
  assign n37073 = ~pi832 & ~n37072;
  assign n37074 = ~n37071 & n37073;
  assign po321 = ~n37037 & ~n37074;
  assign n37076 = ~pi774 & pi947;
  assign n37077 = pi687 & n35430;
  assign n37078 = ~n37076 & ~n37077;
  assign n37079 = n2923 & ~n37078;
  assign n37080 = ~pi165 & ~n2923;
  assign n37081 = pi832 & ~n37080;
  assign n37082 = ~n37079 & n37081;
  assign n37083 = ~pi165 & n35604;
  assign n37084 = pi165 & n35629;
  assign n37085 = ~pi38 & ~n37084;
  assign n37086 = ~n37083 & n37085;
  assign n37087 = ~pi165 & ~n35633;
  assign n37088 = n35636 & ~n37087;
  assign n37089 = ~pi774 & ~n37088;
  assign n37090 = ~n37086 & n37089;
  assign n37091 = ~pi165 & n35651;
  assign n37092 = pi165 & n35670;
  assign n37093 = ~pi38 & ~n37092;
  assign n37094 = ~n37091 & n37093;
  assign n37095 = ~pi165 & ~n7357;
  assign n37096 = n35676 & ~n37095;
  assign n37097 = pi774 & ~n37096;
  assign n37098 = ~n37094 & n37097;
  assign n37099 = ~n37090 & ~n37098;
  assign n37100 = pi687 & ~n37099;
  assign n37101 = pi165 & ~n35705;
  assign n37102 = ~pi774 & ~n37101;
  assign n37103 = ~n35706 & n37102;
  assign n37104 = ~pi165 & ~n8091;
  assign n37105 = pi774 & ~n37104;
  assign n37106 = pi165 & ~n35728;
  assign n37107 = ~pi687 & ~n37106;
  assign n37108 = ~pi774 & n35728;
  assign n37109 = pi165 & ~n37108;
  assign n37110 = pi774 & n8091;
  assign n37111 = ~pi687 & ~n37110;
  assign n37112 = ~n37109 & n37111;
  assign n37113 = ~n37105 & n37107;
  assign n37114 = ~n37103 & n64443;
  assign n37115 = ~n37100 & ~n37114;
  assign n37116 = n63888 & ~n37115;
  assign n37117 = ~pi165 & ~n63888;
  assign n37118 = ~pi832 & ~n37117;
  assign n37119 = ~n37116 & n37118;
  assign po322 = ~n37082 & ~n37119;
  assign n37121 = pi166 & ~n6951;
  assign n37122 = ~n35607 & ~n37121;
  assign n37123 = n7118 & n37122;
  assign n37124 = ~pi215 & ~n37123;
  assign n37125 = pi166 & n35579;
  assign n37126 = n35656 & ~n37125;
  assign n37127 = ~n7124 & n37126;
  assign n37128 = n37124 & ~n37127;
  assign n37129 = ~pi166 & ~n7134;
  assign n37130 = n35576 & ~n37129;
  assign n37131 = pi299 & ~n37130;
  assign n37132 = ~n37128 & n37131;
  assign n37133 = n7034 & n37122;
  assign n37134 = ~pi223 & ~n37133;
  assign n37135 = ~pi166 & ~n62789;
  assign n37136 = ~n36106 & ~n37135;
  assign n37137 = n36075 & ~n37136;
  assign n37138 = n37134 & ~n37137;
  assign n37139 = ~n2915 & ~n62785;
  assign n37140 = ~pi166 & ~n37139;
  assign n37141 = n35591 & ~n37140;
  assign n37142 = ~pi166 & n62785;
  assign n37143 = n35589 & ~n37142;
  assign n37144 = ~pi299 & ~n37143;
  assign n37145 = ~pi299 & ~n37141;
  assign n37146 = ~n37143 & n37145;
  assign n37147 = ~n37141 & n37144;
  assign n37148 = ~n37138 & n64444;
  assign n37149 = pi772 & ~n37148;
  assign n37150 = ~n37132 & n37149;
  assign n37151 = ~n7034 & ~n37136;
  assign n37152 = n7034 & n35719;
  assign n37153 = pi947 & n62790;
  assign n37154 = n37134 & ~n64445;
  assign n37155 = ~n37151 & n37154;
  assign n37156 = n37145 & ~n37155;
  assign n37157 = ~n35577 & n37124;
  assign n37158 = ~n37126 & n37157;
  assign n37159 = ~n36114 & n37130;
  assign n37160 = pi299 & ~n37159;
  assign n37161 = ~n37158 & n37160;
  assign n37162 = ~pi772 & ~n37161;
  assign n37163 = ~pi772 & ~n37156;
  assign n37164 = ~n37161 & n37163;
  assign n37165 = ~n37156 & n37162;
  assign n37166 = pi39 & ~n64446;
  assign n37167 = pi39 & ~n37150;
  assign n37168 = ~n64446 & n37167;
  assign n37169 = ~n37150 & n37166;
  assign n37170 = pi772 & pi947;
  assign n37171 = ~n62781 & n37170;
  assign n37172 = pi166 & n62781;
  assign n37173 = ~pi39 & ~n37172;
  assign n37174 = ~pi39 & ~n37170;
  assign n37175 = ~n7145 & ~n37174;
  assign n37176 = ~n37172 & ~n37175;
  assign n37177 = ~n37171 & n37173;
  assign n37178 = ~n35668 & n64448;
  assign n37179 = ~pi38 & ~n37178;
  assign n37180 = ~n64447 & n37179;
  assign n37181 = n2923 & ~n37170;
  assign n37182 = n7357 & ~n37170;
  assign n37183 = n7356 & n37181;
  assign n37184 = n36133 & n37174;
  assign n37185 = ~n35430 & n64449;
  assign n37186 = ~pi166 & ~n7357;
  assign n37187 = pi38 & ~n37186;
  assign n37188 = pi38 & ~n64450;
  assign n37189 = ~n37186 & n37188;
  assign n37190 = ~n64450 & n37187;
  assign n37191 = pi727 & ~n64451;
  assign n37192 = ~n37180 & n37191;
  assign n37193 = ~n35689 & ~n37126;
  assign n37194 = ~n35578 & ~n37193;
  assign n37195 = ~n35719 & ~n37121;
  assign n37196 = n7118 & n37195;
  assign n37197 = ~pi215 & ~n37196;
  assign n37198 = ~n37194 & n37197;
  assign n37199 = pi166 & n35692;
  assign n37200 = n35717 & ~n37199;
  assign n37201 = ~n37198 & n37200;
  assign n37202 = n7034 & ~n37195;
  assign n37203 = n36072 & ~n37135;
  assign n37204 = ~n37202 & ~n37203;
  assign n37205 = ~pi223 & ~n37204;
  assign n37206 = n37144 & ~n37205;
  assign n37207 = pi772 & ~n37206;
  assign n37208 = ~n37201 & n37207;
  assign n37209 = pi166 & n22049;
  assign n37210 = pi39 & ~n37209;
  assign n37211 = ~n37208 & n37210;
  assign n37212 = ~pi38 & ~n64448;
  assign n37213 = ~n37211 & n37212;
  assign n37214 = pi38 & ~n64449;
  assign n37215 = ~n37186 & n37214;
  assign n37216 = ~pi727 & ~n37215;
  assign n37217 = ~n37213 & n37216;
  assign n37218 = ~n37192 & ~n37217;
  assign n37219 = n63888 & ~n37218;
  assign n37220 = ~pi166 & ~n63888;
  assign n37221 = ~pi832 & ~n37220;
  assign n37222 = ~n37219 & n37221;
  assign n37223 = pi727 & n35430;
  assign n37224 = n37181 & ~n37223;
  assign n37225 = ~pi166 & ~n2923;
  assign n37226 = pi832 & ~n37225;
  assign n37227 = ~n37224 & n37226;
  assign n37228 = ~n37222 & ~n37227;
  assign n37229 = ~pi768 & pi947;
  assign n37230 = pi705 & n35430;
  assign n37231 = ~n37229 & ~n37230;
  assign n37232 = n2923 & ~n37231;
  assign n37233 = ~pi167 & ~n2923;
  assign n37234 = pi832 & ~n37233;
  assign n37235 = ~n37232 & n37234;
  assign n37236 = ~pi167 & n35651;
  assign n37237 = pi167 & n35670;
  assign n37238 = ~pi38 & ~n37237;
  assign n37239 = ~n37236 & n37238;
  assign n37240 = ~pi167 & ~n7357;
  assign n37241 = n35676 & ~n37240;
  assign n37242 = pi768 & ~n37241;
  assign n37243 = ~n37239 & n37242;
  assign n37244 = ~pi167 & n35604;
  assign n37245 = pi167 & n35629;
  assign n37246 = ~pi38 & ~n37245;
  assign n37247 = ~n37244 & n37246;
  assign n37248 = ~pi167 & ~n35633;
  assign n37249 = n35636 & ~n37248;
  assign n37250 = ~pi768 & ~n37249;
  assign n37251 = ~n37247 & n37250;
  assign n37252 = pi705 & ~n37251;
  assign n37253 = pi705 & ~n37243;
  assign n37254 = ~n37251 & n37253;
  assign n37255 = ~n37243 & n37252;
  assign n37256 = ~pi167 & ~n35701;
  assign n37257 = pi167 & n35726;
  assign n37258 = ~pi38 & ~n37257;
  assign n37259 = ~n37256 & n37258;
  assign n37260 = ~n35713 & ~n37240;
  assign n37261 = ~pi768 & ~n37260;
  assign n37262 = ~n37259 & n37261;
  assign n37263 = ~pi167 & pi768;
  assign n37264 = ~pi167 & n21727;
  assign n37265 = ~n8091 & n37263;
  assign n37266 = ~pi705 & ~n64453;
  assign n37267 = ~n37262 & n37266;
  assign n37268 = n63888 & ~n37267;
  assign n37269 = ~n37243 & ~n37251;
  assign n37270 = pi705 & ~n37269;
  assign n37271 = ~pi167 & n64365;
  assign n37272 = ~n37260 & ~n37271;
  assign n37273 = ~pi768 & ~n37272;
  assign n37274 = ~pi768 & ~n35727;
  assign n37275 = pi167 & ~n37274;
  assign n37276 = ~pi705 & ~n21721;
  assign n37277 = ~n37275 & n37276;
  assign n37278 = ~n37273 & n37277;
  assign n37279 = ~n37270 & ~n37278;
  assign n37280 = n63888 & ~n37279;
  assign n37281 = ~n64452 & n37268;
  assign n37282 = ~pi167 & ~n63888;
  assign n37283 = ~pi832 & ~n37282;
  assign n37284 = ~n64454 & n37283;
  assign po324 = ~n37235 & ~n37284;
  assign n37286 = pi168 & ~n7134;
  assign n37287 = n35576 & ~n37286;
  assign n37288 = pi168 & ~n7118;
  assign n37289 = pi168 & n7129;
  assign n37290 = ~n7124 & n37288;
  assign n37291 = ~n7123 & ~n64455;
  assign n37292 = ~pi168 & ~n6951;
  assign n37293 = n35720 & ~n37292;
  assign n37294 = ~n35657 & n37293;
  assign n37295 = ~pi215 & ~n37294;
  assign n37296 = n37291 & n37295;
  assign n37297 = ~n37287 & ~n37296;
  assign n37298 = pi299 & ~n37297;
  assign n37299 = pi168 & ~n35617;
  assign n37300 = n35594 & ~n37299;
  assign n37301 = ~n37298 & ~n37300;
  assign n37302 = pi763 & ~n37301;
  assign n37303 = n35659 & ~n37292;
  assign n37304 = ~n35580 & ~n37303;
  assign n37305 = n37291 & n37304;
  assign n37306 = ~pi215 & ~n37305;
  assign n37307 = n35606 & ~n37287;
  assign n37308 = ~n35641 & ~n37307;
  assign n37309 = ~n37306 & n37308;
  assign n37310 = pi299 & ~n37309;
  assign n37311 = ~pi168 & ~n7116;
  assign n37312 = n35665 & ~n37311;
  assign n37313 = ~pi763 & ~n37312;
  assign n37314 = ~n37310 & n37313;
  assign n37315 = pi39 & ~n37314;
  assign n37316 = ~n37310 & ~n37312;
  assign n37317 = ~pi763 & ~n37316;
  assign n37318 = pi763 & ~n37298;
  assign n37319 = ~n37300 & n37318;
  assign n37320 = ~n37317 & ~n37319;
  assign n37321 = pi39 & ~n37320;
  assign n37322 = ~n37302 & n37315;
  assign n37323 = ~pi168 & n62781;
  assign n37324 = ~n22932 & ~n35715;
  assign n37325 = ~n37323 & ~n37324;
  assign n37326 = ~n35668 & n37325;
  assign n37327 = ~pi38 & ~n37326;
  assign n37328 = ~n64456 & n37327;
  assign n37329 = pi763 & pi947;
  assign n37330 = n2923 & ~n37329;
  assign n37331 = n7357 & ~n37329;
  assign n37332 = n7356 & n37330;
  assign n37333 = ~n35430 & n64457;
  assign n37334 = pi168 & ~n7357;
  assign n37335 = pi38 & ~n37334;
  assign n37336 = ~n37333 & n37335;
  assign n37337 = pi699 & ~n37336;
  assign n37338 = ~n64456 & ~n37326;
  assign n37339 = ~pi38 & ~n37338;
  assign n37340 = ~pi168 & ~n7357;
  assign n37341 = ~pi763 & pi947;
  assign n37342 = ~pi39 & ~n37341;
  assign n37343 = ~n35430 & ~n37329;
  assign n37344 = n7357 & ~n37343;
  assign n37345 = n35876 & n37342;
  assign n37346 = pi38 & ~n64458;
  assign n37347 = pi38 & ~n37340;
  assign n37348 = ~n64458 & n37347;
  assign n37349 = ~n37340 & n37346;
  assign n37350 = ~n37339 & ~n64459;
  assign n37351 = pi699 & ~n37350;
  assign n37352 = ~n37328 & n37337;
  assign n37353 = n35716 & ~n37311;
  assign n37354 = n37291 & ~n37293;
  assign n37355 = n35690 & n37354;
  assign n37356 = n35692 & ~n37286;
  assign n37357 = ~n35653 & n37287;
  assign n37358 = pi299 & ~n64461;
  assign n37359 = ~n37355 & n37358;
  assign n37360 = pi763 & ~n37359;
  assign n37361 = ~n37353 & n37360;
  assign n37362 = ~pi168 & ~pi763;
  assign n37363 = ~n7143 & n37362;
  assign n37364 = pi39 & ~n37363;
  assign n37365 = ~n37361 & n37364;
  assign n37366 = ~pi38 & ~n37325;
  assign n37367 = ~n37365 & n37366;
  assign n37368 = pi38 & ~n64457;
  assign n37369 = ~n37334 & n37368;
  assign n37370 = ~pi699 & ~n37369;
  assign n37371 = ~n37367 & n37370;
  assign n37372 = n27338 & ~n37371;
  assign n37373 = ~n37367 & ~n37369;
  assign n37374 = ~pi699 & ~n37373;
  assign n37375 = pi699 & ~n64459;
  assign n37376 = ~n37339 & n37375;
  assign n37377 = ~n37374 & ~n37376;
  assign n37378 = n27338 & ~n37377;
  assign n37379 = ~n64460 & n37372;
  assign n37380 = ~pi168 & ~n27338;
  assign n37381 = ~pi57 & ~n37380;
  assign n37382 = ~n64462 & n37381;
  assign n37383 = pi57 & pi168;
  assign n37384 = ~pi832 & ~n37383;
  assign n37385 = ~n37382 & n37384;
  assign n37386 = pi699 & n35430;
  assign n37387 = ~pi699 & ~n37329;
  assign n37388 = ~n37343 & ~n37387;
  assign n37389 = n2923 & ~n37388;
  assign n37390 = n37330 & ~n37386;
  assign n37391 = pi168 & ~n2923;
  assign n37392 = pi832 & ~n37391;
  assign n37393 = ~n64463 & n37392;
  assign n37394 = ~n37385 & ~n37393;
  assign n37395 = pi169 & ~n7134;
  assign n37396 = n35576 & ~n37395;
  assign n37397 = pi169 & ~n7118;
  assign n37398 = pi169 & n7129;
  assign n37399 = ~n7124 & n37397;
  assign n37400 = ~n7123 & ~n64464;
  assign n37401 = ~pi169 & ~n6951;
  assign n37402 = n35720 & ~n37401;
  assign n37403 = ~n35657 & n37402;
  assign n37404 = ~pi215 & ~n37403;
  assign n37405 = n37400 & n37404;
  assign n37406 = ~n37396 & ~n37405;
  assign n37407 = pi299 & ~n37406;
  assign n37408 = pi169 & ~n35617;
  assign n37409 = n35594 & ~n37408;
  assign n37410 = ~n37407 & ~n37409;
  assign n37411 = pi746 & ~n37410;
  assign n37412 = n35659 & ~n37401;
  assign n37413 = ~n35580 & ~n37412;
  assign n37414 = n37400 & n37413;
  assign n37415 = ~pi215 & ~n37414;
  assign n37416 = n35606 & ~n37396;
  assign n37417 = ~n35641 & ~n37416;
  assign n37418 = ~n37415 & n37417;
  assign n37419 = pi299 & ~n37418;
  assign n37420 = ~pi169 & ~n7116;
  assign n37421 = n35665 & ~n37420;
  assign n37422 = ~pi746 & ~n37421;
  assign n37423 = ~n37419 & n37422;
  assign n37424 = pi39 & ~n37423;
  assign n37425 = ~n37419 & ~n37421;
  assign n37426 = ~pi746 & ~n37425;
  assign n37427 = pi746 & ~n37407;
  assign n37428 = ~n37409 & n37427;
  assign n37429 = ~n37426 & ~n37428;
  assign n37430 = pi39 & ~n37429;
  assign n37431 = ~n37411 & n37424;
  assign n37432 = ~pi169 & n62781;
  assign n37433 = ~n23535 & ~n35715;
  assign n37434 = ~n37432 & ~n37433;
  assign n37435 = ~n35668 & n37434;
  assign n37436 = ~pi38 & ~n37435;
  assign n37437 = ~n64465 & n37436;
  assign n37438 = pi746 & pi947;
  assign n37439 = n2923 & ~n37438;
  assign n37440 = n7357 & ~n37438;
  assign n37441 = n7356 & n37439;
  assign n37442 = ~n35430 & n64466;
  assign n37443 = pi169 & ~n7357;
  assign n37444 = pi38 & ~n37443;
  assign n37445 = ~n37442 & n37444;
  assign n37446 = pi729 & ~n37445;
  assign n37447 = ~n64465 & ~n37435;
  assign n37448 = ~pi38 & ~n37447;
  assign n37449 = ~pi169 & ~n7357;
  assign n37450 = ~pi746 & pi947;
  assign n37451 = ~pi39 & ~n37450;
  assign n37452 = ~n35430 & ~n37438;
  assign n37453 = n7357 & ~n37452;
  assign n37454 = n35876 & n37451;
  assign n37455 = pi38 & ~n64467;
  assign n37456 = pi38 & ~n37449;
  assign n37457 = ~n64467 & n37456;
  assign n37458 = ~n37449 & n37455;
  assign n37459 = ~n37448 & ~n64468;
  assign n37460 = pi729 & ~n37459;
  assign n37461 = ~n37437 & n37446;
  assign n37462 = n35716 & ~n37420;
  assign n37463 = n37400 & ~n37402;
  assign n37464 = n35690 & n37463;
  assign n37465 = n35692 & ~n37395;
  assign n37466 = ~n35653 & n37396;
  assign n37467 = pi299 & ~n64470;
  assign n37468 = ~n37464 & n37467;
  assign n37469 = pi746 & ~n37468;
  assign n37470 = ~n37462 & n37469;
  assign n37471 = ~pi169 & ~pi746;
  assign n37472 = ~n7143 & n37471;
  assign n37473 = pi39 & ~n37472;
  assign n37474 = ~n37470 & n37473;
  assign n37475 = ~pi38 & ~n37434;
  assign n37476 = ~n37474 & n37475;
  assign n37477 = pi38 & ~n64466;
  assign n37478 = ~n37443 & n37477;
  assign n37479 = ~pi729 & ~n37478;
  assign n37480 = ~n37476 & n37479;
  assign n37481 = n27338 & ~n37480;
  assign n37482 = ~n37476 & ~n37478;
  assign n37483 = ~pi729 & ~n37482;
  assign n37484 = pi729 & ~n64468;
  assign n37485 = ~n37448 & n37484;
  assign n37486 = ~n37483 & ~n37485;
  assign n37487 = n27338 & ~n37486;
  assign n37488 = ~n64469 & n37481;
  assign n37489 = ~pi169 & ~n27338;
  assign n37490 = ~pi57 & ~n37489;
  assign n37491 = ~n64471 & n37490;
  assign n37492 = pi57 & pi169;
  assign n37493 = ~pi832 & ~n37492;
  assign n37494 = ~n37491 & n37493;
  assign n37495 = pi729 & n35430;
  assign n37496 = ~pi729 & ~n37438;
  assign n37497 = ~n37452 & ~n37496;
  assign n37498 = n2923 & ~n37497;
  assign n37499 = n37439 & ~n37495;
  assign n37500 = pi169 & ~n2923;
  assign n37501 = pi832 & ~n37500;
  assign n37502 = ~n64472 & n37501;
  assign n37503 = ~n37494 & ~n37502;
  assign n37504 = pi730 & n35430;
  assign n37505 = pi748 & pi947;
  assign n37506 = n2923 & ~n37505;
  assign n37507 = ~n37504 & n37506;
  assign n37508 = pi170 & ~n2923;
  assign n37509 = pi832 & ~n37508;
  assign n37510 = ~n37507 & n37509;
  assign n37511 = pi170 & ~n7118;
  assign n37512 = pi170 & n7129;
  assign n37513 = ~n7124 & n37511;
  assign n37514 = ~n7123 & ~n64473;
  assign n37515 = ~pi170 & ~n6951;
  assign n37516 = n35659 & ~n37515;
  assign n37517 = ~n35580 & ~n37516;
  assign n37518 = n37514 & n37517;
  assign n37519 = ~pi215 & ~n37518;
  assign n37520 = pi170 & ~n7134;
  assign n37521 = n35576 & ~n37520;
  assign n37522 = n35606 & ~n37521;
  assign n37523 = ~n35641 & ~n37522;
  assign n37524 = ~n37519 & n37523;
  assign n37525 = pi299 & ~n37524;
  assign n37526 = ~pi170 & ~n7116;
  assign n37527 = ~pi299 & ~n37526;
  assign n37528 = ~n35664 & n37527;
  assign n37529 = ~n37525 & ~n37528;
  assign n37530 = pi39 & ~n37529;
  assign n37531 = ~pi170 & n62781;
  assign n37532 = n35669 & ~n37531;
  assign n37533 = ~n37530 & ~n37532;
  assign n37534 = ~pi38 & ~n37533;
  assign n37535 = ~pi170 & ~n7357;
  assign n37536 = n35676 & ~n37535;
  assign n37537 = ~pi748 & ~n37536;
  assign n37538 = ~n37534 & n37537;
  assign n37539 = n35602 & ~n37531;
  assign n37540 = pi170 & ~n35617;
  assign n37541 = n35594 & ~n37540;
  assign n37542 = n35720 & ~n37515;
  assign n37543 = ~n35657 & n37542;
  assign n37544 = ~pi215 & ~n37543;
  assign n37545 = n37514 & n37544;
  assign n37546 = ~n37521 & ~n37545;
  assign n37547 = pi299 & ~n37546;
  assign n37548 = pi39 & ~n37547;
  assign n37549 = ~n37541 & n37548;
  assign n37550 = ~n37539 & ~n37549;
  assign n37551 = ~pi38 & ~n37550;
  assign n37552 = n35636 & ~n37535;
  assign n37553 = pi748 & ~n37552;
  assign n37554 = ~n37551 & n37553;
  assign n37555 = pi730 & ~n37554;
  assign n37556 = ~n37538 & n37555;
  assign n37557 = n35715 & ~n37531;
  assign n37558 = n37514 & ~n37542;
  assign n37559 = n35690 & n37558;
  assign n37560 = ~n35653 & n37521;
  assign n37561 = n35692 & ~n37520;
  assign n37562 = pi299 & ~n64474;
  assign n37563 = ~n37559 & n37562;
  assign n37564 = ~n35684 & n37527;
  assign n37565 = ~n37563 & ~n37564;
  assign n37566 = pi39 & ~n37565;
  assign n37567 = ~n37557 & ~n37566;
  assign n37568 = ~pi38 & ~n37567;
  assign n37569 = ~n35713 & ~n37535;
  assign n37570 = pi748 & ~n37569;
  assign n37571 = ~n37568 & n37570;
  assign n37572 = ~pi170 & ~pi748;
  assign n37573 = ~n8091 & n37572;
  assign n37574 = ~pi730 & ~n37573;
  assign n37575 = ~n37571 & n37574;
  assign n37576 = n27338 & ~n37575;
  assign n37577 = ~n37556 & n37576;
  assign n37578 = ~pi170 & ~n27338;
  assign n37579 = ~pi57 & ~n37578;
  assign n37580 = ~n37577 & n37579;
  assign n37581 = pi57 & pi170;
  assign n37582 = ~pi832 & ~n37581;
  assign n37583 = ~n37580 & n37582;
  assign n37584 = ~n37510 & ~n37583;
  assign n37585 = pi171 & ~n7134;
  assign n37586 = n35576 & ~n37585;
  assign n37587 = pi171 & ~n7118;
  assign n37588 = pi171 & n7129;
  assign n37589 = ~n7124 & n37587;
  assign n37590 = ~n7123 & ~n64475;
  assign n37591 = ~pi171 & ~n6951;
  assign n37592 = n35720 & ~n37591;
  assign n37593 = ~n35657 & n37592;
  assign n37594 = ~pi215 & ~n37593;
  assign n37595 = n37590 & n37594;
  assign n37596 = ~n37586 & ~n37595;
  assign n37597 = pi299 & ~n37596;
  assign n37598 = pi171 & ~n35617;
  assign n37599 = n35594 & ~n37598;
  assign n37600 = ~n37597 & ~n37599;
  assign n37601 = pi764 & ~n37600;
  assign n37602 = n35659 & ~n37591;
  assign n37603 = ~n35580 & ~n37602;
  assign n37604 = n37590 & n37603;
  assign n37605 = ~pi215 & ~n37604;
  assign n37606 = n35606 & ~n37586;
  assign n37607 = ~n35641 & ~n37606;
  assign n37608 = ~n37605 & n37607;
  assign n37609 = pi299 & ~n37608;
  assign n37610 = ~pi171 & ~n7116;
  assign n37611 = n35665 & ~n37610;
  assign n37612 = ~pi764 & ~n37611;
  assign n37613 = ~n37609 & n37612;
  assign n37614 = pi39 & ~n37613;
  assign n37615 = ~n37609 & ~n37611;
  assign n37616 = ~pi764 & ~n37615;
  assign n37617 = pi764 & ~n37597;
  assign n37618 = ~n37599 & n37617;
  assign n37619 = ~n37616 & ~n37618;
  assign n37620 = pi39 & ~n37619;
  assign n37621 = ~n37601 & n37614;
  assign n37622 = ~pi171 & n62781;
  assign n37623 = ~n24138 & ~n35715;
  assign n37624 = ~n37622 & ~n37623;
  assign n37625 = ~n35668 & n37624;
  assign n37626 = ~pi38 & ~n37625;
  assign n37627 = ~n64476 & n37626;
  assign n37628 = pi764 & pi947;
  assign n37629 = n2923 & ~n37628;
  assign n37630 = n7357 & ~n37628;
  assign n37631 = n7356 & n37629;
  assign n37632 = ~n35430 & n64477;
  assign n37633 = pi171 & ~n7357;
  assign n37634 = pi38 & ~n37633;
  assign n37635 = ~n37632 & n37634;
  assign n37636 = pi691 & ~n37635;
  assign n37637 = ~n64476 & ~n37625;
  assign n37638 = ~pi38 & ~n37637;
  assign n37639 = ~pi171 & ~n7357;
  assign n37640 = ~pi764 & pi947;
  assign n37641 = ~pi39 & ~n37640;
  assign n37642 = ~n35430 & ~n37628;
  assign n37643 = n7357 & ~n37642;
  assign n37644 = n35876 & n37641;
  assign n37645 = pi38 & ~n64478;
  assign n37646 = pi38 & ~n37639;
  assign n37647 = ~n64478 & n37646;
  assign n37648 = ~n37639 & n37645;
  assign n37649 = ~n37638 & ~n64479;
  assign n37650 = pi691 & ~n37649;
  assign n37651 = ~n37627 & n37636;
  assign n37652 = n35716 & ~n37610;
  assign n37653 = n37590 & ~n37592;
  assign n37654 = n35690 & n37653;
  assign n37655 = n35692 & ~n37585;
  assign n37656 = ~n35653 & n37586;
  assign n37657 = pi299 & ~n64481;
  assign n37658 = ~n37654 & n37657;
  assign n37659 = pi764 & ~n37658;
  assign n37660 = ~n37652 & n37659;
  assign n37661 = ~pi171 & ~pi764;
  assign n37662 = ~n7143 & n37661;
  assign n37663 = pi39 & ~n37662;
  assign n37664 = ~n37660 & n37663;
  assign n37665 = ~pi38 & ~n37624;
  assign n37666 = ~n37664 & n37665;
  assign n37667 = pi38 & ~n64477;
  assign n37668 = ~n37633 & n37667;
  assign n37669 = ~pi691 & ~n37668;
  assign n37670 = ~n37666 & n37669;
  assign n37671 = n27338 & ~n37670;
  assign n37672 = ~n37666 & ~n37668;
  assign n37673 = ~pi691 & ~n37672;
  assign n37674 = pi691 & ~n64479;
  assign n37675 = ~n37638 & n37674;
  assign n37676 = ~n37673 & ~n37675;
  assign n37677 = n27338 & ~n37676;
  assign n37678 = ~n64480 & n37671;
  assign n37679 = ~pi171 & ~n27338;
  assign n37680 = ~pi57 & ~n37679;
  assign n37681 = ~n64482 & n37680;
  assign n37682 = pi57 & pi171;
  assign n37683 = ~pi832 & ~n37682;
  assign n37684 = ~n37681 & n37683;
  assign n37685 = pi691 & n35430;
  assign n37686 = ~pi691 & ~n37628;
  assign n37687 = ~n37642 & ~n37686;
  assign n37688 = n2923 & ~n37687;
  assign n37689 = n37629 & ~n37685;
  assign n37690 = pi171 & ~n2923;
  assign n37691 = pi832 & ~n37690;
  assign n37692 = ~n64483 & n37691;
  assign n37693 = ~n37684 & ~n37692;
  assign n37694 = pi172 & ~n7357;
  assign n37695 = pi739 & pi947;
  assign n37696 = n2923 & ~n37695;
  assign n37697 = n7357 & ~n37695;
  assign n37698 = n7356 & n37696;
  assign n37699 = pi38 & ~n64484;
  assign n37700 = ~n37694 & n37699;
  assign n37701 = ~pi172 & ~n7116;
  assign n37702 = n35716 & ~n37701;
  assign n37703 = pi172 & ~n7118;
  assign n37704 = pi172 & n7129;
  assign n37705 = ~n7124 & n37703;
  assign n37706 = ~n7123 & ~n64485;
  assign n37707 = ~pi172 & ~n6951;
  assign n37708 = n35720 & ~n37707;
  assign n37709 = n37706 & ~n37708;
  assign n37710 = n35690 & n37709;
  assign n37711 = pi172 & ~n7134;
  assign n37712 = n35576 & ~n37711;
  assign n37713 = n35692 & ~n37711;
  assign n37714 = ~n35653 & n37712;
  assign n37715 = pi299 & ~n64486;
  assign n37716 = ~n37710 & n37715;
  assign n37717 = pi739 & ~n37716;
  assign n37718 = ~n37702 & n37717;
  assign n37719 = ~pi172 & ~pi739;
  assign n37720 = ~n7143 & n37719;
  assign n37721 = pi39 & ~n37720;
  assign n37722 = ~n37718 & n37721;
  assign n37723 = ~n62781 & n37695;
  assign n37724 = ~pi172 & n62781;
  assign n37725 = ~pi39 & ~n37724;
  assign n37726 = ~pi39 & ~n37723;
  assign n37727 = ~n37724 & n37726;
  assign n37728 = ~n37723 & n37725;
  assign n37729 = ~pi38 & ~n64487;
  assign n37730 = ~n37722 & n37729;
  assign n37731 = ~n37700 & ~n37730;
  assign n37732 = ~pi690 & ~n37731;
  assign n37733 = ~n35668 & n64487;
  assign n37734 = ~n35657 & n37708;
  assign n37735 = ~pi215 & ~n37734;
  assign n37736 = n37706 & n37735;
  assign n37737 = ~n37712 & ~n37736;
  assign n37738 = pi299 & ~n37737;
  assign n37739 = pi172 & ~n35617;
  assign n37740 = n35594 & ~n37739;
  assign n37741 = ~n37738 & ~n37740;
  assign n37742 = pi739 & ~n37741;
  assign n37743 = n35659 & ~n37707;
  assign n37744 = ~n35580 & ~n37743;
  assign n37745 = n37706 & n37744;
  assign n37746 = ~pi215 & ~n37745;
  assign n37747 = n35606 & ~n37712;
  assign n37748 = ~n35641 & ~n37747;
  assign n37749 = ~n37746 & n37748;
  assign n37750 = pi299 & ~n37749;
  assign n37751 = n35665 & ~n37701;
  assign n37752 = ~pi739 & ~n37751;
  assign n37753 = ~n37750 & n37752;
  assign n37754 = pi39 & ~n37753;
  assign n37755 = ~n37750 & ~n37751;
  assign n37756 = ~pi739 & ~n37755;
  assign n37757 = pi739 & ~n37738;
  assign n37758 = ~n37740 & n37757;
  assign n37759 = ~n37756 & ~n37758;
  assign n37760 = pi39 & ~n37759;
  assign n37761 = ~n37742 & n37754;
  assign n37762 = ~n37733 & ~n64488;
  assign n37763 = ~pi38 & ~n37762;
  assign n37764 = ~n35430 & ~n37695;
  assign n37765 = ~pi739 & pi947;
  assign n37766 = ~pi39 & ~n37765;
  assign n37767 = n35876 & n37766;
  assign n37768 = n7357 & ~n37764;
  assign n37769 = ~pi172 & ~n7357;
  assign n37770 = pi38 & ~n37769;
  assign n37771 = pi38 & ~n64489;
  assign n37772 = ~n37769 & n37771;
  assign n37773 = ~n64489 & n37770;
  assign n37774 = pi690 & ~n64490;
  assign n37775 = ~n37763 & n37774;
  assign n37776 = ~n37732 & ~n37775;
  assign n37777 = ~n37763 & ~n64490;
  assign n37778 = pi690 & ~n37777;
  assign n37779 = ~pi690 & ~n37700;
  assign n37780 = ~n37730 & n37779;
  assign n37781 = n27338 & ~n37780;
  assign n37782 = ~n37778 & n37781;
  assign n37783 = n27338 & ~n37776;
  assign n37784 = ~pi172 & ~n27338;
  assign n37785 = ~pi57 & ~n37784;
  assign n37786 = ~n64491 & n37785;
  assign n37787 = pi57 & pi172;
  assign n37788 = ~pi832 & ~n37787;
  assign n37789 = ~n37786 & n37788;
  assign n37790 = pi690 & n35430;
  assign n37791 = ~pi690 & ~n37695;
  assign n37792 = ~n37764 & ~n37791;
  assign n37793 = n2923 & ~n37792;
  assign n37794 = n37696 & ~n37790;
  assign n37795 = pi172 & ~n2923;
  assign n37796 = pi832 & ~n37795;
  assign n37797 = ~n64492 & n37796;
  assign n37798 = ~n37789 & ~n37797;
  assign n37799 = ~pi197 & n64356;
  assign n37800 = pi197 & n64361;
  assign n37801 = ~pi767 & ~n37800;
  assign n37802 = ~n37799 & n37801;
  assign n37803 = ~pi197 & n35642;
  assign n37804 = pi197 & n35662;
  assign n37805 = pi299 & ~n37804;
  assign n37806 = ~n37803 & n37805;
  assign n37807 = ~pi197 & ~n7116;
  assign n37808 = n35665 & ~n37807;
  assign n37809 = pi767 & ~n37808;
  assign n37810 = ~n37806 & n37809;
  assign n37811 = pi39 & ~n37810;
  assign n37812 = ~n37802 & n37811;
  assign n37813 = ~pi767 & pi947;
  assign n37814 = ~n62781 & n37813;
  assign n37815 = ~pi197 & n62781;
  assign n37816 = ~pi39 & ~n37815;
  assign n37817 = ~pi39 & ~n37814;
  assign n37818 = ~n37815 & n37817;
  assign n37819 = ~n37814 & n37816;
  assign n37820 = ~n35668 & n64493;
  assign n37821 = ~pi38 & ~n37820;
  assign n37822 = ~n37812 & n37821;
  assign n37823 = n7357 & ~n37813;
  assign n37824 = ~n35430 & n37823;
  assign n37825 = pi197 & ~n7357;
  assign n37826 = pi38 & ~n37825;
  assign n37827 = ~n37824 & n37826;
  assign n37828 = ~pi698 & ~n37827;
  assign n37829 = ~n37822 & n37828;
  assign n37830 = ~pi197 & ~n35693;
  assign n37831 = pi197 & ~n35783;
  assign n37832 = pi299 & ~n37831;
  assign n37833 = ~n37830 & n37832;
  assign n37834 = n35716 & ~n37807;
  assign n37835 = ~pi767 & ~n37834;
  assign n37836 = ~n37833 & n37835;
  assign n37837 = ~pi197 & pi767;
  assign n37838 = ~n7143 & n37837;
  assign n37839 = pi39 & ~n37838;
  assign n37840 = ~n37836 & n37839;
  assign n37841 = ~pi38 & ~n64493;
  assign n37842 = ~n37840 & n37841;
  assign n37843 = pi38 & ~n37823;
  assign n37844 = ~n37825 & n37843;
  assign n37845 = pi698 & ~n37844;
  assign n37846 = ~n37842 & n37845;
  assign n37847 = n63888 & ~n37846;
  assign n37848 = ~n37842 & ~n37844;
  assign n37849 = pi698 & ~n37848;
  assign n37850 = ~n37812 & ~n37820;
  assign n37851 = ~pi38 & ~n37850;
  assign n37852 = ~pi197 & ~n7357;
  assign n37853 = pi767 & pi947;
  assign n37854 = ~pi39 & ~n37853;
  assign n37855 = ~n35430 & ~n37813;
  assign n37856 = n7357 & ~n37855;
  assign n37857 = n35876 & n37854;
  assign n37858 = pi38 & ~n64494;
  assign n37859 = pi38 & ~n37852;
  assign n37860 = ~n64494 & n37859;
  assign n37861 = ~n37852 & n37858;
  assign n37862 = ~pi698 & ~n64495;
  assign n37863 = ~n37851 & n37862;
  assign n37864 = ~n37849 & ~n37863;
  assign n37865 = n63888 & ~n37864;
  assign n37866 = ~n37829 & n37847;
  assign n37867 = ~pi197 & ~n63888;
  assign n37868 = ~pi832 & ~n37867;
  assign n37869 = ~n64496 & n37868;
  assign n37870 = ~pi698 & n35430;
  assign n37871 = ~n37813 & ~n37870;
  assign n37872 = n2923 & ~n37871;
  assign n37873 = ~pi197 & ~n2923;
  assign n37874 = pi832 & ~n37873;
  assign n37875 = ~n37872 & n37874;
  assign po354 = ~n37869 & ~n37875;
  assign n37877 = ~pi100 & ~n35405;
  assign n37878 = n30886 & ~n37877;
  assign n37879 = ~pi75 & ~n37878;
  assign n37880 = ~n30600 & ~n37879;
  assign n37881 = ~pi92 & ~n37880;
  assign n37882 = ~pi74 & n3471;
  assign n37883 = n3470 & n34040;
  assign n37884 = ~pi74 & n62455;
  assign n37885 = n3473 & n34040;
  assign n37886 = n3472 & n64497;
  assign n37887 = ~pi54 & ~n30604;
  assign n37888 = n64498 & n37887;
  assign n37889 = ~n30604 & n35113;
  assign po288 = ~n37881 & n64499;
  assign n37891 = n62765 & ~n36374;
  assign n37892 = pi606 & n37891;
  assign n37893 = n62765 & ~n36370;
  assign n37894 = ~pi606 & n37893;
  assign n37895 = pi643 & ~n37894;
  assign n37896 = pi643 & ~n37892;
  assign n37897 = ~n37894 & n37896;
  assign n37898 = ~n37892 & n37895;
  assign n37899 = n62765 & ~n35706;
  assign n37900 = pi606 & n37899;
  assign n37901 = ~pi606 & n8098;
  assign n37902 = n8091 & n26393;
  assign n37903 = ~pi643 & ~n64501;
  assign n37904 = ~n37900 & n37903;
  assign n37905 = n62455 & ~n37904;
  assign n37906 = ~n64500 & n37905;
  assign n37907 = pi211 & ~n37906;
  assign n37908 = n62765 & n36346;
  assign n37909 = pi606 & ~n37908;
  assign n37910 = n62765 & n36343;
  assign n37911 = ~pi606 & ~n37910;
  assign n37912 = pi643 & ~n37911;
  assign n37913 = pi643 & ~n37909;
  assign n37914 = ~n37911 & n37913;
  assign n37915 = ~n37909 & n37912;
  assign n37916 = n62765 & n35728;
  assign n37917 = pi606 & ~pi643;
  assign n37918 = n37916 & n37917;
  assign n37919 = ~n64502 & ~n37918;
  assign n37920 = ~pi211 & n62455;
  assign n37921 = ~n37919 & n37920;
  assign n37922 = ~n37907 & ~n37921;
  assign n37923 = pi607 & n37891;
  assign n37924 = ~pi607 & n37893;
  assign n37925 = pi638 & ~n37924;
  assign n37926 = pi638 & ~n37923;
  assign n37927 = ~n37924 & n37926;
  assign n37928 = ~n37923 & n37925;
  assign n37929 = pi607 & n37899;
  assign n37930 = ~pi607 & n8098;
  assign n37931 = ~pi638 & ~n37930;
  assign n37932 = ~n37929 & n37931;
  assign n37933 = n62455 & ~n37932;
  assign n37934 = ~n64503 & n37933;
  assign n37935 = ~pi212 & ~n37934;
  assign n37936 = ~pi607 & ~n37910;
  assign n37937 = pi607 & ~n37908;
  assign n37938 = pi638 & ~n37937;
  assign n37939 = pi638 & ~n37936;
  assign n37940 = ~n37937 & n37939;
  assign n37941 = ~n37936 & n37938;
  assign n37942 = pi607 & ~pi638;
  assign n37943 = n37916 & n37942;
  assign n37944 = ~n64504 & ~n37943;
  assign n37945 = pi212 & n62455;
  assign n37946 = ~n37944 & n37945;
  assign n37947 = ~n37935 & ~n37946;
  assign n37948 = pi213 & n62455;
  assign n37949 = ~pi622 & ~n37910;
  assign n37950 = pi622 & ~n37908;
  assign n37951 = pi639 & ~n37950;
  assign n37952 = pi639 & ~n37949;
  assign n37953 = ~n37950 & n37952;
  assign n37954 = ~n37949 & n37951;
  assign n37955 = pi622 & ~pi639;
  assign n37956 = n37916 & n37955;
  assign n37957 = ~n64505 & ~n37956;
  assign n37958 = n37948 & ~n37957;
  assign n37959 = pi639 & ~n37891;
  assign n37960 = ~pi639 & ~n37899;
  assign n37961 = pi622 & ~n37960;
  assign n37962 = pi622 & ~n37959;
  assign n37963 = ~n37960 & n37962;
  assign n37964 = ~n37959 & n37961;
  assign n37965 = pi639 & ~n37893;
  assign n37966 = ~pi639 & ~n8098;
  assign n37967 = ~pi622 & ~n37966;
  assign n37968 = ~n37965 & n37967;
  assign n37969 = ~n64506 & ~n37968;
  assign n37970 = pi639 & n37891;
  assign n37971 = ~pi639 & n37899;
  assign n37972 = pi622 & ~n37971;
  assign n37973 = pi622 & ~n37970;
  assign n37974 = ~n37971 & n37973;
  assign n37975 = ~n37970 & n37972;
  assign n37976 = pi639 & n37893;
  assign n37977 = ~pi639 & n8098;
  assign n37978 = ~pi622 & ~n37977;
  assign n37979 = ~n37976 & n37978;
  assign n37980 = n62455 & ~n37979;
  assign n37981 = ~n64507 & n37980;
  assign n37982 = n62455 & ~n37969;
  assign n37983 = ~pi213 & ~n64508;
  assign n37984 = ~n37958 & ~n37983;
  assign n37985 = pi623 & n37891;
  assign n37986 = ~pi623 & n37893;
  assign n37987 = pi710 & ~n37986;
  assign n37988 = pi710 & ~n37985;
  assign n37989 = ~n37986 & n37988;
  assign n37990 = ~n37985 & n37987;
  assign n37991 = pi623 & n37899;
  assign n37992 = ~pi623 & n8098;
  assign n37993 = ~pi710 & ~n37992;
  assign n37994 = ~n37991 & n37993;
  assign n37995 = n62455 & ~n37994;
  assign n37996 = ~n64509 & n37995;
  assign n37997 = ~pi214 & ~n37996;
  assign n37998 = ~pi623 & ~n37910;
  assign n37999 = pi623 & ~n37908;
  assign n38000 = pi710 & ~n37999;
  assign n38001 = pi710 & ~n37998;
  assign n38002 = ~n37999 & n38001;
  assign n38003 = ~n37998 & n38000;
  assign n38004 = pi623 & ~pi710;
  assign n38005 = n37916 & n38004;
  assign n38006 = ~n64510 & ~n38005;
  assign n38007 = pi214 & n62455;
  assign n38008 = ~n38006 & n38007;
  assign n38009 = ~n37997 & ~n38008;
  assign n38010 = ~pi219 & n62455;
  assign n38011 = ~pi617 & ~n37910;
  assign n38012 = pi617 & ~n37908;
  assign n38013 = pi637 & ~n38012;
  assign n38014 = pi637 & ~n38011;
  assign n38015 = ~n38012 & n38014;
  assign n38016 = ~n38011 & n38013;
  assign n38017 = pi617 & ~pi637;
  assign n38018 = n37916 & n38017;
  assign n38019 = ~n64511 & ~n38018;
  assign n38020 = n38010 & ~n38019;
  assign n38021 = ~pi617 & n37893;
  assign n38022 = pi617 & n37891;
  assign n38023 = pi637 & ~n38022;
  assign n38024 = pi637 & ~n38021;
  assign n38025 = ~n38022 & n38024;
  assign n38026 = ~n38021 & n38023;
  assign n38027 = pi617 & n37899;
  assign n38028 = ~pi617 & n8098;
  assign n38029 = ~pi637 & ~n38028;
  assign n38030 = ~n38027 & n38029;
  assign n38031 = n62455 & ~n38030;
  assign n38032 = ~pi617 & ~n37893;
  assign n38033 = pi617 & ~n37891;
  assign n38034 = pi637 & ~n38033;
  assign n38035 = ~n38032 & n38034;
  assign n38036 = pi617 & ~n37899;
  assign n38037 = ~pi617 & ~n8098;
  assign n38038 = ~pi637 & ~n38037;
  assign n38039 = ~n38036 & n38038;
  assign n38040 = ~n38035 & ~n38039;
  assign n38041 = n62455 & ~n38040;
  assign n38042 = ~n64512 & n38031;
  assign n38043 = pi219 & ~n64513;
  assign n38044 = ~n38020 & ~n38043;
  assign n38045 = pi210 & ~n6951;
  assign n38046 = n2908 & n38045;
  assign n38047 = pi210 & ~n2908;
  assign n38048 = ~n7076 & n38047;
  assign n38049 = ~n38046 & ~n38048;
  assign n38050 = ~pi907 & n38049;
  assign n38051 = ~n27801 & ~n38045;
  assign n38052 = ~n2909 & ~n38051;
  assign n38053 = pi907 & ~n38052;
  assign n38054 = pi210 & n7055;
  assign n38055 = pi634 & ~n7055;
  assign n38056 = ~n38054 & ~n38055;
  assign n38057 = n2909 & ~n38056;
  assign n38058 = n38053 & ~n38057;
  assign n38059 = ~pi947 & ~n38058;
  assign n38060 = ~n38050 & n38059;
  assign n38061 = ~n27593 & ~n38045;
  assign n38062 = n2908 & n38061;
  assign n38063 = pi947 & ~n38062;
  assign n38064 = pi633 & ~n7055;
  assign n38065 = ~n38054 & ~n38064;
  assign n38066 = ~n2814 & ~n38065;
  assign n38067 = ~n2908 & n38061;
  assign n38068 = ~n2909 & ~n38067;
  assign n38069 = ~n38066 & ~n38068;
  assign n38070 = n38063 & ~n38069;
  assign n38071 = n2971 & ~n38070;
  assign n38072 = ~n38060 & n38071;
  assign n38073 = n2953 & n38051;
  assign n38074 = pi907 & ~n38073;
  assign n38075 = ~n2953 & n38056;
  assign n38076 = n38074 & ~n38075;
  assign n38077 = pi210 & ~n62787;
  assign n38078 = ~pi907 & n38077;
  assign n38079 = ~n38076 & ~n38078;
  assign n38080 = ~pi947 & ~n38079;
  assign n38081 = n2953 & n38061;
  assign n38082 = pi947 & ~n38081;
  assign n38083 = ~n2953 & n38065;
  assign n38084 = n38082 & ~n38083;
  assign n38085 = ~n2971 & ~n38084;
  assign n38086 = ~n38080 & n38085;
  assign n38087 = ~n38072 & ~n38086;
  assign n38088 = ~n7034 & ~n38087;
  assign n38089 = pi634 & n35430;
  assign n38090 = pi633 & pi947;
  assign n38091 = ~n38089 & ~n38090;
  assign n38092 = n6951 & ~n38091;
  assign n38093 = ~n38045 & ~n38092;
  assign n38094 = n7034 & n38093;
  assign n38095 = ~pi223 & ~n38094;
  assign n38096 = ~n38088 & n38095;
  assign n38097 = ~n6979 & n38047;
  assign n38098 = ~n38046 & ~n38097;
  assign n38099 = ~pi907 & n38098;
  assign n38100 = pi210 & n6971;
  assign n38101 = ~n27811 & ~n38100;
  assign n38102 = n2909 & ~n38101;
  assign n38103 = n38053 & ~n38102;
  assign n38104 = ~pi947 & ~n38103;
  assign n38105 = ~n38099 & n38104;
  assign n38106 = pi633 & ~n6971;
  assign n38107 = ~n38100 & ~n38106;
  assign n38108 = ~n2814 & ~n38107;
  assign n38109 = ~n38068 & ~n38108;
  assign n38110 = n38063 & ~n38109;
  assign n38111 = n2971 & ~n38110;
  assign n38112 = ~n38105 & n38111;
  assign n38113 = ~n2953 & n38101;
  assign n38114 = n38074 & ~n38113;
  assign n38115 = n2953 & n6950;
  assign n38116 = n2923 & n38115;
  assign n38117 = n38100 & ~n38116;
  assign n38118 = ~n38114 & ~n38117;
  assign n38119 = ~pi947 & ~n38118;
  assign n38120 = ~n2953 & n38107;
  assign n38121 = n38082 & ~n38120;
  assign n38122 = ~n2971 & ~n38121;
  assign n38123 = ~n38119 & n38122;
  assign n38124 = pi223 & ~n38123;
  assign n38125 = pi223 & ~n38112;
  assign n38126 = ~n38123 & n38125;
  assign n38127 = ~n38112 & n38124;
  assign n38128 = ~pi299 & ~n64514;
  assign n38129 = ~n38096 & n38128;
  assign n38130 = ~n2914 & ~n38077;
  assign n38131 = n2914 & n38049;
  assign n38132 = ~pi907 & ~n38131;
  assign n38133 = ~n38130 & n38132;
  assign n38134 = ~n38076 & ~n38133;
  assign n38135 = ~pi947 & ~n38134;
  assign n38136 = ~n7118 & ~n38084;
  assign n38137 = ~n38135 & n38136;
  assign n38138 = n7118 & n38093;
  assign n38139 = ~pi215 & ~n38138;
  assign n38140 = ~n38137 & n38139;
  assign n38141 = n2914 & n38098;
  assign n38142 = ~n2914 & ~n38117;
  assign n38143 = ~pi907 & ~n38142;
  assign n38144 = ~n38141 & n38143;
  assign n38145 = ~n38114 & ~n38144;
  assign n38146 = ~pi947 & ~n38145;
  assign n38147 = ~n38121 & ~n38146;
  assign n38148 = pi215 & ~n38147;
  assign n38149 = pi299 & ~n38148;
  assign n38150 = ~n38140 & n38149;
  assign n38151 = pi39 & ~n38150;
  assign n38152 = ~n38129 & n38151;
  assign n38153 = n6940 & ~n38091;
  assign n38154 = pi210 & ~n6940;
  assign n38155 = ~pi299 & ~n38154;
  assign n38156 = ~pi299 & ~n38153;
  assign n38157 = ~n38154 & n38156;
  assign n38158 = ~n38153 & n38155;
  assign n38159 = ~n6906 & ~n38091;
  assign n38160 = pi299 & ~n6935;
  assign n38161 = pi299 & ~n38159;
  assign n38162 = ~n6935 & n38161;
  assign n38163 = ~n38159 & n38160;
  assign n38164 = ~pi39 & ~n64516;
  assign n38165 = ~n64515 & n38164;
  assign n38166 = ~pi38 & ~n38165;
  assign n38167 = ~n38152 & n38166;
  assign n38168 = n7357 & ~n38091;
  assign n38169 = pi210 & ~n7357;
  assign n38170 = pi38 & ~n38169;
  assign n38171 = pi38 & ~n38168;
  assign n38172 = ~n38169 & n38171;
  assign n38173 = ~n38168 & n38170;
  assign n38174 = ~n38167 & ~n64517;
  assign n38175 = n63888 & ~n38174;
  assign n38176 = ~pi210 & ~n63888;
  assign po367 = ~n38175 & ~n38176;
  assign n38178 = ~pi51 & pi70;
  assign n38179 = n62364 & n38178;
  assign n38180 = ~pi96 & n38179;
  assign n38181 = pi24 & n64339;
  assign n38182 = pi24 & n35394;
  assign n38183 = n2748 & n38179;
  assign n38184 = n2726 & n38180;
  assign n38185 = n38182 & n64518;
  assign n38186 = n38180 & n38181;
  assign n38187 = pi198 & pi589;
  assign n38188 = n2979 & n7034;
  assign n38189 = ~pi223 & n7034;
  assign n38190 = n30841 & n38189;
  assign n38191 = ~n2973 & n38188;
  assign n38192 = n38187 & n64520;
  assign n38193 = pi210 & pi589;
  assign n38194 = ~pi221 & n2959;
  assign n38195 = ~pi216 & n64521;
  assign n38196 = n2959 & n7118;
  assign n38197 = ~n2920 & n2959;
  assign n38198 = n7118 & n38197;
  assign n38199 = ~pi215 & n7118;
  assign n38200 = n30831 & n38199;
  assign n38201 = ~n2920 & n64522;
  assign n38202 = n38193 & n64523;
  assign n38203 = ~n38192 & ~n38202;
  assign n38204 = ~pi593 & n2938;
  assign n38205 = ~n30817 & n38204;
  assign n38206 = ~n38203 & n38205;
  assign n38207 = ~pi287 & ~n38206;
  assign n38208 = pi39 & ~n38207;
  assign n38209 = n62380 & n38208;
  assign n38210 = ~n64519 & ~n38209;
  assign po228 = n64325 & ~n38210;
  assign n38212 = ~n38193 & n64523;
  assign n38213 = ~n2973 & n2979;
  assign n38214 = n7034 & ~n38187;
  assign n38215 = n38213 & n38214;
  assign n38216 = ~n38187 & n64520;
  assign n38217 = ~n38212 & ~n64524;
  assign n38218 = ~n30820 & ~n38217;
  assign n38219 = ~n38187 & n38188;
  assign n38220 = n33178 & n38219;
  assign n38221 = ~n30820 & n38212;
  assign n38222 = pi39 & ~n38221;
  assign n38223 = ~n38220 & n38222;
  assign n38224 = pi39 & ~n38218;
  assign n38225 = pi24 & n30617;
  assign n38226 = n2726 & n32731;
  assign n38227 = n38225 & n38226;
  assign n38228 = ~pi71 & n2587;
  assign n38229 = ~pi104 & n2591;
  assign n38230 = n38228 & n38229;
  assign n38231 = ~pi49 & ~pi66;
  assign n38232 = ~pi45 & ~pi73;
  assign n38233 = n38231 & n38232;
  assign n38234 = ~pi48 & ~pi65;
  assign n38235 = pi89 & n38234;
  assign n38236 = n38233 & n38235;
  assign n38237 = pi89 & n31458;
  assign n38238 = n38234 & n38237;
  assign n38239 = n38233 & n38238;
  assign n38240 = n64146 & n38239;
  assign n38241 = n64145 & n38236;
  assign n38242 = n38230 & n64526;
  assign n38243 = n2670 & n38242;
  assign n38244 = ~pi332 & n64196;
  assign n38245 = ~pi841 & n2694;
  assign n38246 = n38244 & n38245;
  assign n38247 = n38243 & n38245;
  assign n38248 = n38244 & n38247;
  assign n38249 = n38243 & n38246;
  assign n38250 = ~pi39 & ~n64527;
  assign n38251 = ~n38227 & n38250;
  assign n38252 = n64325 & ~n38251;
  assign po253 = ~n64525 & n38252;
  assign n38254 = pi39 & pi593;
  assign n38255 = ~n38203 & n38254;
  assign n38256 = ~n30820 & n38255;
  assign n38257 = n2874 & n64293;
  assign n38258 = n2783 & n62390;
  assign n38259 = pi829 & ~pi1093;
  assign n38260 = n2582 & n38259;
  assign n38261 = ~n62395 & ~n38260;
  assign n38262 = pi479 & n38261;
  assign n38263 = ~n64148 & n38262;
  assign n38264 = ~po740 & ~n38263;
  assign n38265 = n64338 & ~n38264;
  assign n38266 = n64528 & n38265;
  assign n38267 = ~n38256 & ~n38266;
  assign po255 = n64325 & ~n38267;
  assign n38269 = pi215 & ~n63888;
  assign n38270 = pi681 & pi907;
  assign n38271 = n36071 & ~n38270;
  assign n38272 = ~pi642 & n62787;
  assign n38273 = ~n2971 & ~n38272;
  assign n38274 = n7078 & n7186;
  assign n38275 = ~n7077 & n7190;
  assign n38276 = ~pi642 & n29114;
  assign n38277 = n6951 & n29529;
  assign n38278 = ~n2907 & ~n64530;
  assign n38279 = ~n64529 & n38278;
  assign n38280 = n2907 & ~n29122;
  assign n38281 = ~n38279 & ~n38280;
  assign n38282 = ~n64529 & ~n64530;
  assign n38283 = ~n2907 & ~n38282;
  assign n38284 = n2907 & n29122;
  assign n38285 = n2971 & ~n38284;
  assign n38286 = ~n38283 & n38285;
  assign n38287 = n2971 & ~n38281;
  assign n38288 = pi947 & ~n64531;
  assign n38289 = n2971 & ~n38280;
  assign n38290 = ~n38279 & n38289;
  assign n38291 = ~n2971 & n38272;
  assign n38292 = ~n38290 & ~n38291;
  assign n38293 = pi947 & ~n38292;
  assign n38294 = pi947 & ~n38273;
  assign n38295 = ~n64531 & n38294;
  assign n38296 = ~n38273 & n38288;
  assign n38297 = ~n7034 & ~n64532;
  assign n38298 = ~n38271 & n38297;
  assign n38299 = ~n6951 & n7034;
  assign n38300 = ~pi947 & n38270;
  assign n38301 = pi642 & pi947;
  assign n38302 = ~n38300 & ~n38301;
  assign n38303 = n7034 & ~n38302;
  assign n38304 = ~pi223 & ~n38303;
  assign n38305 = n6951 & n38302;
  assign n38306 = n7034 & ~n38305;
  assign n38307 = ~pi223 & ~n38306;
  assign n38308 = ~n38299 & n38304;
  assign n38309 = ~n38298 & n64533;
  assign n38310 = ~n2907 & ~n6992;
  assign n38311 = n7008 & n7012;
  assign n38312 = n2907 & ~n6979;
  assign n38313 = ~pi642 & ~n64534;
  assign n38314 = ~pi642 & n62784;
  assign n38315 = ~n38310 & n38313;
  assign n38316 = n2971 & ~n64535;
  assign n38317 = ~n2907 & ~n62783;
  assign n38318 = ~pi642 & ~n28374;
  assign n38319 = ~n38317 & n38318;
  assign n38320 = ~n2971 & ~n38319;
  assign n38321 = pi947 & ~n38320;
  assign n38322 = ~n38316 & n38321;
  assign n38323 = ~n35588 & ~n38322;
  assign n38324 = pi223 & ~n38300;
  assign n38325 = ~n38323 & n38324;
  assign n38326 = ~pi299 & ~n38325;
  assign n38327 = ~n38309 & n38326;
  assign n38328 = ~pi947 & n35995;
  assign n38329 = pi947 & ~n38319;
  assign n38330 = ~n38300 & ~n38329;
  assign n38331 = ~n38328 & n38330;
  assign n38332 = pi299 & ~n38331;
  assign n38333 = ~n38327 & ~n38332;
  assign n38334 = pi215 & ~n38333;
  assign n38335 = n7084 & n38300;
  assign n38336 = pi642 & ~n7008;
  assign n38337 = n6951 & n38336;
  assign n38338 = pi642 & n7008;
  assign n38339 = ~n7017 & n38338;
  assign n38340 = ~n7095 & n38339;
  assign n38341 = ~n38337 & ~n38340;
  assign n38342 = pi947 & ~n38341;
  assign n38343 = n2971 & ~n38342;
  assign n38344 = ~n38335 & n38343;
  assign n38345 = ~n62786 & n38270;
  assign n38346 = ~pi947 & ~n38345;
  assign n38347 = ~n2907 & n7057;
  assign n38348 = ~n7065 & ~n38347;
  assign n38349 = n38338 & n38348;
  assign n38350 = ~n7057 & n38336;
  assign n38351 = pi947 & ~n38350;
  assign n38352 = ~n38349 & n38351;
  assign n38353 = ~n38346 & ~n38352;
  assign n38354 = ~n2971 & ~n38353;
  assign n38355 = ~n7034 & ~n38354;
  assign n38356 = ~n38344 & n38355;
  assign n38357 = n62790 & ~n38302;
  assign n38358 = n6951 & n38303;
  assign n38359 = ~pi223 & ~n64536;
  assign n38360 = ~n38356 & n38359;
  assign n38361 = n2971 & ~n6992;
  assign n38362 = n38270 & ~n38361;
  assign n38363 = ~pi947 & ~n38362;
  assign n38364 = pi947 & ~n6973;
  assign n38365 = ~n62783 & ~n38364;
  assign n38366 = ~n2971 & n38365;
  assign n38367 = ~n7012 & n38339;
  assign n38368 = pi947 & ~n38337;
  assign n38369 = ~n38367 & n38368;
  assign n38370 = ~n38366 & ~n38369;
  assign n38371 = ~n38363 & n38370;
  assign n38372 = pi223 & ~n38371;
  assign n38373 = ~n38360 & ~n38372;
  assign n38374 = ~pi299 & ~n38373;
  assign n38375 = ~n7118 & n38353;
  assign n38376 = n7126 & ~n38302;
  assign n38377 = pi299 & ~n38376;
  assign n38378 = ~n38375 & n38377;
  assign n38379 = ~pi215 & ~n38378;
  assign n38380 = ~n38374 & n38379;
  assign n38381 = ~n38334 & ~n38380;
  assign n38382 = pi39 & ~n38381;
  assign n38383 = n6936 & n38302;
  assign n38384 = ~pi215 & ~n6936;
  assign n38385 = pi299 & ~n38384;
  assign n38386 = ~n38383 & n38385;
  assign n38387 = n6940 & n38302;
  assign n38388 = ~pi215 & ~n6940;
  assign n38389 = ~pi299 & ~n38388;
  assign n38390 = ~n38387 & n38389;
  assign n38391 = ~n38386 & ~n38390;
  assign n38392 = n6940 & ~n38302;
  assign n38393 = pi215 & ~n6940;
  assign n38394 = ~pi299 & ~n38393;
  assign n38395 = ~pi299 & ~n38392;
  assign n38396 = ~n38393 & n38395;
  assign n38397 = ~n38392 & n38394;
  assign n38398 = pi215 & ~n6936;
  assign n38399 = n6936 & ~n38302;
  assign n38400 = pi299 & ~n38399;
  assign n38401 = pi299 & ~n38398;
  assign n38402 = ~n38399 & n38401;
  assign n38403 = ~n38398 & n38400;
  assign n38404 = ~pi39 & ~n64538;
  assign n38405 = ~n64537 & n38404;
  assign n38406 = ~pi39 & ~n64537;
  assign n38407 = ~n64538 & n38406;
  assign n38408 = ~pi39 & ~n38391;
  assign n38409 = ~pi38 & ~n64539;
  assign n38410 = ~n38382 & n38409;
  assign n38411 = n7357 & ~n38302;
  assign n38412 = pi215 & ~n7357;
  assign n38413 = pi38 & ~n38412;
  assign n38414 = pi38 & ~n38411;
  assign n38415 = ~n38412 & n38414;
  assign n38416 = ~n38411 & n38413;
  assign n38417 = n63888 & ~n64540;
  assign n38418 = ~n38410 & n38417;
  assign n38419 = ~n38269 & ~n38418;
  assign n38420 = pi216 & ~n7357;
  assign n38421 = pi662 & pi907;
  assign n38422 = ~pi947 & n38421;
  assign n38423 = pi614 & pi947;
  assign n38424 = ~n38422 & ~n38423;
  assign n38425 = n7357 & ~n38424;
  assign n38426 = pi38 & ~n38425;
  assign n38427 = pi38 & ~n38420;
  assign n38428 = ~n38425 & n38427;
  assign n38429 = ~n38420 & n38426;
  assign n38430 = ~n7012 & n7097;
  assign n38431 = pi947 & ~n7100;
  assign n38432 = ~n38430 & n38431;
  assign n38433 = ~n38364 & ~n38422;
  assign n38434 = ~n38432 & ~n38433;
  assign n38435 = n62783 & n38421;
  assign n38436 = ~pi947 & ~n38435;
  assign n38437 = pi947 & n6973;
  assign n38438 = ~n38432 & ~n38437;
  assign n38439 = ~n38436 & n38438;
  assign n38440 = ~n38365 & n38434;
  assign n38441 = ~pi216 & ~n64542;
  assign n38442 = n7087 & ~n64041;
  assign n38443 = n62783 & n7087;
  assign n38444 = n2907 & n29909;
  assign n38445 = ~n64543 & ~n38444;
  assign n38446 = pi947 & n38445;
  assign n38447 = pi216 & ~n38422;
  assign n38448 = ~n38446 & n38447;
  assign n38449 = ~n38328 & n38448;
  assign n38450 = ~n38441 & ~n38449;
  assign n38451 = pi215 & ~n38450;
  assign n38452 = ~pi947 & n35688;
  assign n38453 = pi947 & ~n62787;
  assign n38454 = ~pi614 & n62787;
  assign n38455 = pi947 & ~n38454;
  assign n38456 = ~n38422 & ~n38455;
  assign n38457 = n38424 & ~n38453;
  assign n38458 = ~n38452 & n64544;
  assign n38459 = n62953 & n38424;
  assign n38460 = pi216 & ~n64545;
  assign n38461 = n38348 & n38423;
  assign n38462 = ~n62786 & n38422;
  assign n38463 = ~n38461 & ~n38462;
  assign n38464 = n2958 & ~n38463;
  assign n38465 = n7126 & ~n38424;
  assign n38466 = ~pi215 & ~n38465;
  assign n38467 = ~n38464 & n38466;
  assign n38468 = pi216 & ~n62953;
  assign n38469 = n38424 & ~n38468;
  assign n38470 = ~pi216 & ~n7126;
  assign n38471 = ~n38469 & ~n38470;
  assign n38472 = ~pi215 & ~n38464;
  assign n38473 = ~n38471 & n38472;
  assign n38474 = ~n38460 & n38467;
  assign n38475 = ~n38451 & ~n64546;
  assign n38476 = ~n38464 & ~n38465;
  assign n38477 = ~n38460 & n38476;
  assign n38478 = ~pi215 & ~n38477;
  assign n38479 = pi215 & ~n38441;
  assign n38480 = ~n38449 & n38479;
  assign n38481 = pi299 & ~n38480;
  assign n38482 = ~n38478 & n38481;
  assign n38483 = pi299 & ~n38475;
  assign n38484 = pi947 & ~n7094;
  assign n38485 = ~pi947 & ~n38421;
  assign n38486 = ~pi947 & n7104;
  assign n38487 = ~n38421 & n38486;
  assign n38488 = n7104 & n38485;
  assign n38489 = ~n38484 & ~n64548;
  assign n38490 = n2971 & ~n38489;
  assign n38491 = ~pi947 & ~n62787;
  assign n38492 = ~n2971 & ~n38491;
  assign n38493 = n64544 & n38492;
  assign n38494 = ~n2971 & ~n38422;
  assign n38495 = ~n38455 & n38494;
  assign n38496 = ~n38491 & n38495;
  assign n38497 = n7073 & n38424;
  assign n38498 = ~n7034 & ~n64549;
  assign n38499 = ~n38490 & n38498;
  assign n38500 = n7034 & ~n38424;
  assign n38501 = ~pi223 & ~n38500;
  assign n38502 = n6951 & n38424;
  assign n38503 = n7034 & ~n38502;
  assign n38504 = ~pi223 & ~n38503;
  assign n38505 = ~n38299 & n38501;
  assign n38506 = ~n38499 & n64550;
  assign n38507 = ~pi616 & n6981;
  assign n38508 = ~n2907 & ~n7021;
  assign n38509 = ~n38507 & n38508;
  assign n38510 = ~pi614 & ~n64534;
  assign n38511 = ~pi616 & ~n6981;
  assign n38512 = ~n2907 & ~n6988;
  assign n38513 = ~n38511 & n38512;
  assign n38514 = ~n7004 & ~n38513;
  assign n38515 = ~pi614 & ~n38514;
  assign n38516 = ~n38509 & n38510;
  assign n38517 = n2971 & ~n64551;
  assign n38518 = ~n2971 & n38445;
  assign n38519 = pi947 & ~n38518;
  assign n38520 = ~n38517 & n38519;
  assign n38521 = ~n35588 & ~n38520;
  assign n38522 = pi223 & ~n38422;
  assign n38523 = ~n38521 & n38522;
  assign n38524 = pi216 & ~n38523;
  assign n38525 = ~n38506 & n38524;
  assign n38526 = n7084 & n38422;
  assign n38527 = pi947 & ~n7101;
  assign n38528 = n2971 & ~n38527;
  assign n38529 = ~n38526 & n38528;
  assign n38530 = ~n2971 & n38463;
  assign n38531 = ~n7034 & ~n38530;
  assign n38532 = ~n38529 & n38531;
  assign n38533 = n62790 & ~n38424;
  assign n38534 = n6951 & n38500;
  assign n38535 = ~pi223 & ~n64552;
  assign n38536 = ~n38532 & n38535;
  assign n38537 = ~n38361 & n38421;
  assign n38538 = ~pi947 & ~n38537;
  assign n38539 = ~n38366 & ~n38432;
  assign n38540 = ~n38538 & n38539;
  assign n38541 = pi223 & ~n38540;
  assign n38542 = ~pi216 & ~n38541;
  assign n38543 = ~n38536 & n38542;
  assign n38544 = ~pi299 & ~n38543;
  assign n38545 = ~n38525 & n38544;
  assign n38546 = pi39 & ~n38545;
  assign n38547 = ~n64547 & n38546;
  assign n38548 = n6936 & n38424;
  assign n38549 = ~pi216 & ~n6936;
  assign n38550 = pi299 & ~n38549;
  assign n38551 = ~n38548 & n38550;
  assign n38552 = n6940 & n38424;
  assign n38553 = ~pi216 & ~n6940;
  assign n38554 = ~pi299 & ~n38553;
  assign n38555 = ~n38552 & n38554;
  assign n38556 = ~n38551 & ~n38555;
  assign n38557 = n6940 & ~n38424;
  assign n38558 = pi216 & ~n6940;
  assign n38559 = ~pi299 & ~n38558;
  assign n38560 = ~pi299 & ~n38557;
  assign n38561 = ~n38558 & n38560;
  assign n38562 = ~n38557 & n38559;
  assign n38563 = pi216 & ~n6936;
  assign n38564 = n6936 & ~n38424;
  assign n38565 = pi299 & ~n38564;
  assign n38566 = pi299 & ~n38563;
  assign n38567 = ~n38564 & n38566;
  assign n38568 = ~n38563 & n38565;
  assign n38569 = ~pi39 & ~n64554;
  assign n38570 = ~n64553 & n38569;
  assign n38571 = ~pi39 & ~n64553;
  assign n38572 = ~n64554 & n38571;
  assign n38573 = ~pi39 & ~n38556;
  assign n38574 = ~pi38 & ~n64555;
  assign n38575 = ~n38547 & n38574;
  assign n38576 = ~n64541 & ~n38575;
  assign n38577 = n63888 & ~n38576;
  assign n38578 = ~pi216 & ~n63888;
  assign po373 = ~n38577 & ~n38578;
  assign n38580 = n7009 & n7082;
  assign n38581 = n7094 & ~n7098;
  assign n38582 = n7013 & ~n38581;
  assign n38583 = ~n38580 & ~n38582;
  assign n38584 = pi947 & ~n38583;
  assign n38585 = n2971 & ~n38486;
  assign n38586 = ~n38584 & n38585;
  assign n38587 = pi661 & pi907;
  assign n38588 = ~pi947 & n38587;
  assign n38589 = n7009 & ~n28303;
  assign n38590 = ~n38272 & ~n38349;
  assign n38591 = n7013 & ~n38590;
  assign n38592 = pi947 & ~n38591;
  assign n38593 = ~n38589 & ~n38591;
  assign n38594 = pi947 & n38593;
  assign n38595 = ~n38589 & n38592;
  assign n38596 = ~n38491 & ~n64556;
  assign n38597 = ~n2971 & ~n38596;
  assign n38598 = ~n38588 & ~n38597;
  assign n38599 = n62789 & ~n38587;
  assign n38600 = ~pi947 & ~n38599;
  assign n38601 = n2971 & ~n38583;
  assign n38602 = ~n2971 & ~n38593;
  assign n38603 = pi947 & ~n38602;
  assign n38604 = ~n38601 & n38603;
  assign n38605 = ~n38600 & ~n38604;
  assign n38606 = ~n38586 & n38598;
  assign n38607 = ~n7034 & ~n64557;
  assign n38608 = pi616 & pi947;
  assign n38609 = ~n38588 & ~n38608;
  assign n38610 = n6951 & ~n38609;
  assign n38611 = n7034 & n38610;
  assign n38612 = n62790 & ~n38609;
  assign n38613 = ~pi223 & ~n64558;
  assign n38614 = ~n38299 & n38613;
  assign n38615 = ~n7034 & ~n38604;
  assign n38616 = ~n38600 & n38615;
  assign n38617 = ~n62790 & ~n38616;
  assign n38618 = n38613 & ~n38617;
  assign n38619 = ~n38607 & n38614;
  assign n38620 = ~pi947 & ~n7002;
  assign n38621 = ~n6973 & ~n6982;
  assign n38622 = ~n2907 & ~n38621;
  assign n38623 = ~pi616 & ~n28374;
  assign n38624 = ~n38622 & n38623;
  assign n38625 = pi947 & ~n38624;
  assign n38626 = ~n38620 & ~n38625;
  assign n38627 = ~n2971 & ~n38626;
  assign n38628 = ~pi947 & n62784;
  assign n38629 = pi947 & ~n7016;
  assign n38630 = n2971 & ~n38629;
  assign n38631 = ~n38628 & n38630;
  assign n38632 = pi223 & ~n38588;
  assign n38633 = ~n38631 & n38632;
  assign n38634 = ~n38627 & n38633;
  assign n38635 = pi221 & ~n38634;
  assign n38636 = ~n64559 & n38635;
  assign n38637 = n7084 & n38588;
  assign n38638 = n7019 & ~n7095;
  assign n38639 = ~n7022 & ~n38638;
  assign n38640 = pi947 & ~n38639;
  assign n38641 = n2971 & ~n38640;
  assign n38642 = ~n38637 & n38641;
  assign n38643 = n38348 & n38608;
  assign n38644 = ~n62786 & n38588;
  assign n38645 = ~n38643 & ~n38644;
  assign n38646 = ~n2971 & n38645;
  assign n38647 = ~n7034 & ~n38646;
  assign n38648 = ~n38642 & n38647;
  assign n38649 = n38613 & ~n38648;
  assign n38650 = pi947 & ~n7023;
  assign n38651 = ~n38588 & ~n38650;
  assign n38652 = ~n38366 & ~n38651;
  assign n38653 = ~n38361 & n38652;
  assign n38654 = pi223 & ~n38653;
  assign n38655 = ~pi221 & ~n38654;
  assign n38656 = ~n38649 & n38655;
  assign n38657 = ~pi299 & ~n38656;
  assign n38658 = ~n38636 & n38657;
  assign n38659 = ~pi947 & ~n38587;
  assign n38660 = ~n35688 & n38659;
  assign n38661 = ~n35688 & ~n38587;
  assign n38662 = ~pi947 & ~n64560;
  assign n38663 = pi221 & ~n64556;
  assign n38664 = pi947 & ~n38593;
  assign n38665 = ~n64560 & ~n38664;
  assign n38666 = pi221 & ~n38665;
  assign n38667 = ~n38662 & n38663;
  assign n38668 = pi216 & ~n38645;
  assign n38669 = ~pi216 & ~n38609;
  assign n38670 = ~pi216 & n38610;
  assign n38671 = n6951 & n38669;
  assign n38672 = ~pi221 & ~n64562;
  assign n38673 = ~n38668 & n38672;
  assign n38674 = ~pi215 & ~n38673;
  assign n38675 = ~n64561 & n38674;
  assign n38676 = pi221 & ~n38588;
  assign n38677 = ~n38625 & n38676;
  assign n38678 = ~n38328 & n38677;
  assign n38679 = ~n38365 & ~n38651;
  assign n38680 = ~pi221 & ~n38679;
  assign n38681 = pi215 & ~n38680;
  assign n38682 = ~n38678 & n38681;
  assign n38683 = pi299 & ~n38682;
  assign n38684 = ~n38675 & n38683;
  assign n38685 = pi39 & ~n38684;
  assign n38686 = pi39 & ~n38658;
  assign n38687 = ~n38684 & n38686;
  assign n38688 = ~n38658 & n38685;
  assign n38689 = n6936 & n38609;
  assign n38690 = ~pi221 & ~n6936;
  assign n38691 = pi299 & ~n38690;
  assign n38692 = ~n38689 & n38691;
  assign n38693 = n6940 & n38609;
  assign n38694 = ~pi221 & ~n6940;
  assign n38695 = ~pi299 & ~n38694;
  assign n38696 = ~n38693 & n38695;
  assign n38697 = ~n38692 & ~n38696;
  assign n38698 = n6940 & ~n38609;
  assign n38699 = pi221 & ~n6940;
  assign n38700 = ~pi299 & ~n38699;
  assign n38701 = ~pi299 & ~n38698;
  assign n38702 = ~n38699 & n38701;
  assign n38703 = ~n38698 & n38700;
  assign n38704 = pi221 & ~n6936;
  assign n38705 = n6936 & ~n38609;
  assign n38706 = pi299 & ~n38705;
  assign n38707 = pi299 & ~n38704;
  assign n38708 = ~n38705 & n38707;
  assign n38709 = ~n38704 & n38706;
  assign n38710 = ~pi39 & ~n64565;
  assign n38711 = ~n64564 & n38710;
  assign n38712 = ~pi39 & ~n64564;
  assign n38713 = ~n64565 & n38712;
  assign n38714 = ~pi39 & ~n38697;
  assign n38715 = ~pi38 & ~n64566;
  assign n38716 = ~n64563 & n38715;
  assign n38717 = pi221 & ~n7357;
  assign n38718 = n7357 & ~n38609;
  assign n38719 = pi38 & ~n38718;
  assign n38720 = pi38 & ~n38717;
  assign n38721 = ~n38718 & n38720;
  assign n38722 = ~n38717 & n38719;
  assign n38723 = ~n38716 & ~n64567;
  assign n38724 = n63888 & ~n38723;
  assign n38725 = ~pi221 & ~n63888;
  assign po378 = ~n38724 & ~n38725;
  assign n38727 = n63888 & ~n30606;
  assign n38728 = pi829 & pi1091;
  assign n38729 = n6924 & n38728;
  assign n38730 = ~n62778 & ~n64148;
  assign n38731 = ~n38729 & n38730;
  assign n38732 = ~n2852 & n6868;
  assign n38733 = ~n6894 & n64148;
  assign n38734 = ~n38732 & n38733;
  assign n38735 = ~n30813 & ~n38734;
  assign n38736 = ~n38731 & n38735;
  assign n38737 = ~pi824 & ~n38728;
  assign n38738 = n2582 & ~n38737;
  assign n38739 = ~n64148 & ~n38738;
  assign n38740 = n6868 & n38739;
  assign n38741 = n6868 & n30813;
  assign n38742 = pi1093 & ~n38741;
  assign n38743 = ~n38740 & n38742;
  assign n38744 = ~n6894 & ~n38732;
  assign n38745 = ~n30813 & ~n38744;
  assign n38746 = n64148 & ~n38745;
  assign n38747 = n6868 & ~n38738;
  assign n38748 = ~n30813 & ~n38731;
  assign n38749 = ~n38747 & ~n38748;
  assign n38750 = ~n38746 & ~n38749;
  assign n38751 = n38742 & ~n38750;
  assign n38752 = n6925 & n38728;
  assign n38753 = ~pi824 & ~n38752;
  assign n38754 = pi824 & ~n6916;
  assign n38755 = ~n30813 & ~n38754;
  assign n38756 = ~n30813 & ~n38753;
  assign n38757 = ~n38754 & n38756;
  assign n38758 = ~n38753 & n38755;
  assign n38759 = ~n6868 & ~n64569;
  assign n38760 = ~n30813 & n64148;
  assign n38761 = n38728 & n38753;
  assign n38762 = ~n38754 & ~n38761;
  assign n38763 = n30814 & ~n38762;
  assign n38764 = ~n38760 & ~n38763;
  assign n38765 = ~n38759 & n38764;
  assign n38766 = ~n38759 & ~n38760;
  assign n38767 = ~n38744 & n38760;
  assign n38768 = pi1093 & ~n38767;
  assign n38769 = ~n64570 & n38768;
  assign n38770 = ~n38736 & n38743;
  assign n38771 = ~n2584 & n6868;
  assign n38772 = n62382 & n62771;
  assign n38773 = n62768 & n6848;
  assign n38774 = ~n6853 & n64571;
  assign n38775 = ~pi40 & ~n38774;
  assign n38776 = n6802 & ~n38775;
  assign n38777 = pi252 & ~n38776;
  assign n38778 = n2584 & ~n6841;
  assign n38779 = ~n38777 & n38778;
  assign n38780 = ~pi1093 & ~n38779;
  assign n38781 = ~n38771 & n38780;
  assign n38782 = ~pi39 & ~n38781;
  assign n38783 = ~n64568 & n38782;
  assign n38784 = ~n2909 & n6950;
  assign n38785 = ~n2583 & n2851;
  assign n38786 = n6947 & ~n38785;
  assign n38787 = n7040 & n38785;
  assign n38788 = pi1091 & ~n38787;
  assign n38789 = pi1091 & ~n38786;
  assign n38790 = ~n38787 & n38789;
  assign n38791 = ~n38786 & n38788;
  assign n38792 = ~n3322 & n6947;
  assign n38793 = n3322 & n7040;
  assign n38794 = ~pi1091 & ~n38793;
  assign n38795 = ~pi1091 & ~n38792;
  assign n38796 = ~n38793 & n38795;
  assign n38797 = ~n38792 & n38794;
  assign n38798 = ~n64572 & ~n64573;
  assign n38799 = ~pi120 & ~n38798;
  assign n38800 = ~n6949 & ~n38799;
  assign n38801 = n2909 & n38800;
  assign n38802 = ~n38784 & ~n38801;
  assign n38803 = n2971 & n38802;
  assign n38804 = ~n2953 & n38800;
  assign n38805 = ~n38115 & ~n38804;
  assign n38806 = ~n2971 & n38805;
  assign n38807 = ~n7034 & ~n38806;
  assign n38808 = ~n7034 & ~n38803;
  assign n38809 = ~n38806 & n38808;
  assign n38810 = ~n38803 & n38807;
  assign n38811 = ~pi223 & ~n7111;
  assign n38812 = ~n64574 & n38811;
  assign n38813 = pi120 & n33980;
  assign n38814 = n6950 & ~n38813;
  assign n38815 = ~n38115 & ~n38814;
  assign n38816 = ~n2971 & ~n38815;
  assign n38817 = ~n38784 & ~n38814;
  assign n38818 = n2971 & ~n38817;
  assign n38819 = pi223 & ~n38818;
  assign n38820 = pi223 & ~n38816;
  assign n38821 = ~n38818 & n38820;
  assign n38822 = ~n38816 & n38819;
  assign n38823 = ~pi299 & ~n64575;
  assign n38824 = ~n38812 & n38823;
  assign n38825 = n62393 & n38802;
  assign n38826 = ~n62393 & n38805;
  assign n38827 = ~n7118 & ~n38826;
  assign n38828 = ~n7118 & ~n38825;
  assign n38829 = ~n38826 & n38828;
  assign n38830 = ~n38825 & n38827;
  assign n38831 = ~pi215 & ~n7315;
  assign n38832 = ~n64576 & n38831;
  assign n38833 = ~n62393 & ~n38815;
  assign n38834 = n62393 & ~n38817;
  assign n38835 = pi215 & ~n38834;
  assign n38836 = pi215 & ~n38833;
  assign n38837 = ~n38834 & n38836;
  assign n38838 = ~n38833 & n38835;
  assign n38839 = pi299 & ~n64577;
  assign n38840 = ~n38832 & n38839;
  assign n38841 = ~n38824 & ~n38840;
  assign n38842 = pi39 & ~n38841;
  assign n38843 = ~pi38 & ~n38842;
  assign n38844 = ~pi38 & ~n38783;
  assign n38845 = ~n38842 & n38844;
  assign n38846 = ~n38783 & n38843;
  assign po387 = n38727 & ~n64578;
  assign n38848 = ~n7039 & n64298;
  assign n38849 = pi1093 & n38848;
  assign n38850 = n2933 & n2937;
  assign n38851 = ~n38849 & n38850;
  assign n38852 = ~pi223 & n38851;
  assign n38853 = ~n2953 & n38848;
  assign n38854 = n38850 & ~n38853;
  assign n38855 = ~n2971 & n38854;
  assign n38856 = n2909 & n38848;
  assign n38857 = n38850 & ~n38856;
  assign n38858 = n2971 & n38857;
  assign n38859 = ~pi299 & ~n38858;
  assign n38860 = ~pi299 & ~n38855;
  assign n38861 = ~n38858 & n38860;
  assign n38862 = ~n38855 & n38859;
  assign n38863 = ~n38852 & n64579;
  assign n38864 = ~pi215 & n38851;
  assign n38865 = ~n62393 & n38854;
  assign n38866 = n62393 & n38857;
  assign n38867 = pi299 & ~n38866;
  assign n38868 = pi299 & ~n38865;
  assign n38869 = ~n38866 & n38868;
  assign n38870 = ~n38865 & n38867;
  assign n38871 = ~n38864 & n64580;
  assign n38872 = pi786 & ~pi1082;
  assign n38873 = ~n38871 & ~n38872;
  assign n38874 = ~n38863 & ~n38872;
  assign n38875 = ~n38871 & n38874;
  assign n38876 = ~n38863 & n38873;
  assign n38877 = ~n38197 & ~n38213;
  assign n38878 = po740 & n38872;
  assign n38879 = ~n38877 & n38878;
  assign n38880 = n2939 & n38879;
  assign n38881 = ~n64581 & ~n38880;
  assign n38882 = pi39 & ~n38881;
  assign n38883 = n30610 & ~n64148;
  assign n38884 = ~pi89 & ~pi102;
  assign n38885 = n2687 & n38884;
  assign n38886 = n2611 & n6806;
  assign n38887 = n38885 & n38886;
  assign n38888 = n31455 & n38887;
  assign n38889 = ~pi65 & ~pi69;
  assign n38890 = n6805 & n38889;
  assign n38891 = pi48 & ~pi49;
  assign n38892 = ~pi68 & ~pi82;
  assign n38893 = n38891 & n38892;
  assign n38894 = n38232 & n38893;
  assign n38895 = n38890 & n38894;
  assign n38896 = n38888 & n38895;
  assign n38897 = n38230 & n38896;
  assign n38898 = ~pi47 & ~pi841;
  assign n38899 = n38897 & n38898;
  assign n38900 = ~n6845 & ~n38899;
  assign n38901 = ~pi986 & ~po740;
  assign n38902 = pi252 & ~n38901;
  assign n38903 = pi314 & ~n38902;
  assign n38904 = n62353 & n2663;
  assign n38905 = ~n38903 & n38904;
  assign n38906 = ~n38900 & n38905;
  assign n38907 = n2641 & n33870;
  assign n38908 = n2642 & ~n33869;
  assign n38909 = ~pi841 & n2637;
  assign n38910 = n2682 & n38909;
  assign n38911 = ~pi97 & n38910;
  assign n38912 = n38897 & n38911;
  assign n38913 = n64582 & n38912;
  assign n38914 = ~pi47 & ~n6858;
  assign n38915 = ~n38913 & n38914;
  assign n38916 = n6848 & n38903;
  assign n38917 = ~n38915 & n38916;
  assign n38918 = ~n38906 & ~n38917;
  assign n38919 = n2694 & ~n38918;
  assign n38920 = ~pi35 & ~n38919;
  assign n38921 = ~pi32 & n6844;
  assign n38922 = n2750 & n6843;
  assign n38923 = ~n38920 & n64583;
  assign n38924 = ~n38883 & ~n38923;
  assign n38925 = n32019 & ~n38924;
  assign n38926 = ~n38882 & ~n38925;
  assign po197 = n64325 & ~n38926;
  assign n38928 = pi39 & ~n35102;
  assign n38929 = ~pi314 & pi1050;
  assign n38930 = n64197 & n38929;
  assign n38931 = ~pi39 & ~n38930;
  assign n38932 = n64325 & ~n38931;
  assign n38933 = pi39 & n35102;
  assign n38934 = ~pi39 & n38929;
  assign n38935 = n64197 & n38934;
  assign n38936 = ~n38933 & ~n38935;
  assign n38937 = n64325 & ~n38936;
  assign n38938 = ~n38928 & n38932;
  assign n38939 = pi72 & n38225;
  assign n38940 = n2685 & n62361;
  assign n38941 = pi88 & n38940;
  assign n38942 = n62768 & n64099;
  assign n38943 = n38941 & n38942;
  assign n38944 = n6873 & n38941;
  assign n38945 = n38942 & n38944;
  assign n38946 = n6873 & n38943;
  assign n38947 = ~n38939 & ~n64585;
  assign n38948 = n2751 & ~n38947;
  assign n38949 = ~pi39 & ~n38948;
  assign n38950 = n62401 & n35099;
  assign n38951 = n62404 & n35096;
  assign n38952 = pi39 & ~n38951;
  assign n38953 = pi39 & ~n38950;
  assign n38954 = ~n38951 & n38953;
  assign n38955 = ~n38950 & n38952;
  assign n38956 = n64325 & ~n64586;
  assign po230 = ~n38949 & n38956;
  assign n38958 = ~pi100 & n27583;
  assign n38959 = n6796 & n38958;
  assign n38960 = ~n33217 & n38959;
  assign n38961 = n62400 & n64234;
  assign n38962 = n62402 & n64232;
  assign n38963 = ~n38961 & ~n38962;
  assign n38964 = n38959 & ~n38963;
  assign n38965 = n62397 & n38960;
  assign n38966 = pi92 & n62380;
  assign n38967 = n64083 & n38929;
  assign n38968 = n38966 & n38967;
  assign n38969 = ~n64587 & ~n38968;
  assign po250 = n35113 & ~n38969;
  assign n38971 = ~pi39 & pi228;
  assign n38972 = ~n64520 & ~n64523;
  assign n38973 = pi39 & ~n38972;
  assign n38974 = n30819 & n38973;
  assign n38975 = ~pi96 & ~n64528;
  assign n38976 = pi96 & ~n64294;
  assign n38977 = n2726 & ~n38976;
  assign n38978 = ~n2924 & ~n38260;
  assign n38979 = n35394 & ~n38978;
  assign n38980 = n38977 & n38979;
  assign n38981 = ~n38975 & n38980;
  assign n38982 = ~n38974 & ~n38981;
  assign n38983 = n64325 & ~n38982;
  assign n38984 = ~n38971 & ~n38983;
  assign n38985 = pi207 & pi208;
  assign n38986 = pi42 & ~pi72;
  assign n38987 = ~pi39 & ~n38986;
  assign n38988 = ~pi72 & pi199;
  assign n38989 = ~pi232 & ~n38988;
  assign n38990 = ~pi299 & ~n38989;
  assign n38991 = ~pi72 & ~n32501;
  assign n38992 = pi199 & n38991;
  assign n38993 = pi232 & ~n38992;
  assign n38994 = n38990 & ~n38993;
  assign n38995 = ~pi72 & pi200;
  assign n38996 = ~pi232 & ~n38995;
  assign n38997 = ~pi299 & ~n38996;
  assign n38998 = pi200 & n38991;
  assign n38999 = pi232 & ~n38998;
  assign n39000 = n38997 & ~n38999;
  assign n39001 = pi39 & ~n39000;
  assign n39002 = ~n38994 & n39001;
  assign n39003 = ~n38987 & ~n39002;
  assign n39004 = ~n2580 & n39003;
  assign n39005 = n38985 & ~n39004;
  assign n39006 = ~pi115 & n2929;
  assign n39007 = n38986 & ~n39006;
  assign n39008 = n2997 & ~n39007;
  assign n39009 = pi114 & ~n38986;
  assign n39010 = n39006 & ~n39009;
  assign n39011 = n2825 & n2827;
  assign n39012 = ~pi44 & n62380;
  assign n39013 = ~pi101 & n39012;
  assign n39014 = n2993 & n39013;
  assign n39015 = n2825 & n39013;
  assign n39016 = n2827 & n39015;
  assign n39017 = n2993 & n39016;
  assign n39018 = n39011 & n39014;
  assign n39019 = ~pi114 & ~n2838;
  assign n39020 = n64588 & n39019;
  assign n39021 = n62385 & n39020;
  assign n39022 = ~pi42 & n39020;
  assign n39023 = n62385 & n39022;
  assign n39024 = ~pi42 & n39021;
  assign n39025 = ~pi24 & n30617;
  assign n39026 = n2993 & n31078;
  assign n39027 = n39025 & n39026;
  assign n39028 = ~pi44 & n39027;
  assign n39029 = n2826 & n39028;
  assign n39030 = ~pi113 & n39029;
  assign n39031 = ~pi116 & n39030;
  assign n39032 = n38986 & ~n39031;
  assign n39033 = ~pi114 & ~n39032;
  assign n39034 = ~n64589 & n39033;
  assign n39035 = n39010 & ~n39034;
  assign n39036 = n39008 & ~n39035;
  assign n39037 = ~n2997 & ~n38986;
  assign n39038 = n62951 & ~n39037;
  assign n39039 = ~n39036 & n39038;
  assign n39040 = ~n62951 & n38986;
  assign n39041 = ~pi39 & ~n39040;
  assign n39042 = ~n39039 & n39041;
  assign n39043 = pi75 & ~n39042;
  assign n39044 = n2751 & n30617;
  assign n39045 = ~pi44 & n39044;
  assign n39046 = pi228 & n2826;
  assign n39047 = n2826 & n39045;
  assign n39048 = pi228 & n39047;
  assign n39049 = n39045 & n39046;
  assign n39050 = pi228 & n2827;
  assign n39051 = n39047 & n39050;
  assign n39052 = n2827 & n39047;
  assign n39053 = pi228 & n39052;
  assign n39054 = n2827 & n64590;
  assign n39055 = ~pi115 & n64591;
  assign n39056 = ~pi114 & n39055;
  assign n39057 = n2829 & n64591;
  assign n39058 = n2839 & n64590;
  assign n39059 = n38986 & ~n64592;
  assign n39060 = pi228 & n62386;
  assign n39061 = pi228 & n2825;
  assign n39062 = pi228 & n39015;
  assign n39063 = n39013 & n39061;
  assign n39064 = ~pi113 & n64593;
  assign n39065 = pi228 & n39016;
  assign n39066 = ~pi116 & n39064;
  assign n39067 = n62386 & n64594;
  assign n39068 = ~pi115 & n64594;
  assign n39069 = ~pi114 & n39068;
  assign n39070 = ~pi42 & n39069;
  assign n39071 = n39016 & n39060;
  assign n39072 = n62373 & ~n64595;
  assign n39073 = n62373 & ~n39059;
  assign n39074 = ~n64595 & n39073;
  assign n39075 = ~n39059 & n39072;
  assign n39076 = ~n2766 & n38987;
  assign n39077 = pi87 & ~n39076;
  assign n39078 = ~n64596 & n39077;
  assign n39079 = ~pi75 & n39078;
  assign n39080 = ~n39043 & ~n39079;
  assign n39081 = ~pi166 & n2815;
  assign n39082 = pi232 & n32363;
  assign n39083 = ~pi72 & ~n64597;
  assign n39084 = pi299 & n39083;
  assign n39085 = pi39 & ~n39084;
  assign n39086 = ~n38994 & n39085;
  assign n39087 = n39001 & n39086;
  assign n39088 = ~n39080 & ~n39087;
  assign n39089 = pi42 & ~pi114;
  assign n39090 = pi72 & pi116;
  assign n39091 = pi72 & pi113;
  assign n39092 = pi72 & ~n2825;
  assign n39093 = ~pi72 & pi101;
  assign n39094 = ~pi41 & ~n39093;
  assign n39095 = pi44 & pi72;
  assign n39096 = n2755 & ~n2758;
  assign n39097 = ~pi72 & ~n62368;
  assign n39098 = ~n2742 & n39097;
  assign n39099 = ~pi1093 & ~n39098;
  assign n39100 = ~pi1093 & ~n39096;
  assign n39101 = ~n39098 & n39100;
  assign n39102 = ~n39096 & n39099;
  assign n39103 = n62368 & ~n2742;
  assign n39104 = ~pi122 & n30950;
  assign n39105 = n62371 & ~n30949;
  assign n39106 = ~n39103 & ~n64599;
  assign n39107 = ~pi72 & n39106;
  assign n39108 = pi1093 & ~n39107;
  assign n39109 = ~n64598 & ~n39108;
  assign n39110 = ~pi44 & ~n39109;
  assign n39111 = ~n39095 & ~n39110;
  assign n39112 = ~pi101 & n39111;
  assign n39113 = n39094 & ~n39112;
  assign n39114 = ~pi99 & n39113;
  assign n39115 = ~n39092 & ~n39114;
  assign n39116 = ~pi113 & ~n39115;
  assign n39117 = ~n39091 & ~n39116;
  assign n39118 = ~pi116 & ~n39117;
  assign n39119 = ~n39090 & ~n39118;
  assign n39120 = n39089 & ~n39119;
  assign n39121 = ~pi1093 & ~n39103;
  assign n39122 = ~pi1093 & ~n62372;
  assign n39123 = ~n39103 & n39122;
  assign n39124 = ~n62372 & n39121;
  assign n39125 = ~pi44 & ~n64600;
  assign n39126 = pi1093 & n39106;
  assign n39127 = n39125 & ~n39126;
  assign n39128 = ~pi101 & n39127;
  assign n39129 = n2825 & n39128;
  assign n39130 = n2826 & n39127;
  assign n39131 = n2827 & n64601;
  assign n39132 = n39011 & n39128;
  assign n39133 = ~pi42 & ~n64602;
  assign n39134 = ~n39009 & ~n39133;
  assign n39135 = ~n39120 & n39134;
  assign n39136 = n39006 & ~n39135;
  assign n39137 = n39097 & ~n64598;
  assign n39138 = ~pi44 & ~n39137;
  assign n39139 = ~n39095 & ~n39138;
  assign n39140 = ~pi101 & n39139;
  assign n39141 = n39094 & ~n39140;
  assign n39142 = ~pi99 & n39141;
  assign n39143 = ~n39092 & ~n39142;
  assign n39144 = ~pi113 & ~n39143;
  assign n39145 = ~n39091 & ~n39144;
  assign n39146 = ~pi116 & ~n39145;
  assign n39147 = ~n39090 & ~n39146;
  assign n39148 = pi42 & n39147;
  assign n39149 = pi1093 & ~n62368;
  assign n39150 = n39125 & ~n39149;
  assign n39151 = ~pi101 & n39150;
  assign n39152 = n2825 & n39151;
  assign n39153 = n2826 & n39150;
  assign n39154 = n2827 & n64603;
  assign n39155 = n39011 & n39151;
  assign n39156 = ~pi42 & n64604;
  assign n39157 = ~pi114 & ~n39156;
  assign n39158 = ~n39148 & n39157;
  assign n39159 = ~n39009 & ~n39158;
  assign n39160 = ~pi115 & ~n2929;
  assign n39161 = ~n39159 & n39160;
  assign n39162 = pi115 & ~n38986;
  assign n39163 = pi228 & ~n39162;
  assign n39164 = ~n39161 & n39163;
  assign n39165 = ~n39136 & n39164;
  assign n39166 = pi110 & n34951;
  assign n39167 = ~pi480 & pi949;
  assign n39168 = n64089 & n39167;
  assign n39169 = pi901 & ~pi959;
  assign n39170 = ~pi250 & pi252;
  assign n39171 = n39169 & n39170;
  assign n39172 = n2751 & ~n39171;
  assign n39173 = n39168 & n39172;
  assign n39174 = n39166 & n39173;
  assign n39175 = n62361 & n33872;
  assign n39176 = n64089 & ~n39167;
  assign n39177 = n64089 & n39175;
  assign n39178 = ~n39167 & n39177;
  assign n39179 = n39175 & n39176;
  assign n39180 = n2698 & n33872;
  assign n39181 = ~pi110 & ~n39180;
  assign n39182 = n2663 & ~n33929;
  assign n39183 = ~pi47 & n39168;
  assign n39184 = n39182 & n39183;
  assign n39185 = ~n39181 & n39184;
  assign n39186 = ~n64605 & ~n39185;
  assign n39187 = ~pi250 & n39169;
  assign n39188 = n31078 & n39187;
  assign n39189 = ~n39186 & n39188;
  assign n39190 = ~n39174 & ~n39189;
  assign n39191 = ~pi44 & ~n39190;
  assign n39192 = n39169 & ~n64605;
  assign n39193 = n39169 & ~n39185;
  assign n39194 = ~n64605 & n39193;
  assign n39195 = ~n39185 & n39192;
  assign n39196 = n39166 & n39168;
  assign n39197 = ~n39169 & ~n39196;
  assign n39198 = n2751 & n39170;
  assign n39199 = ~n39197 & n39198;
  assign n39200 = ~n64606 & n39199;
  assign n39201 = n2751 & ~n39170;
  assign n39202 = n39196 & n39201;
  assign n39203 = ~pi72 & ~n39202;
  assign n39204 = ~n39200 & n39203;
  assign n39205 = ~pi44 & ~n39204;
  assign n39206 = ~n39095 & ~n39205;
  assign n39207 = ~pi72 & ~n39191;
  assign n39208 = ~pi101 & n64607;
  assign n39209 = n39094 & ~n39208;
  assign n39210 = ~pi99 & n39209;
  assign n39211 = ~n39092 & ~n39210;
  assign n39212 = ~pi113 & ~n39211;
  assign n39213 = ~n39091 & ~n39212;
  assign n39214 = ~pi116 & ~n39213;
  assign n39215 = ~n39090 & ~n39214;
  assign n39216 = n39089 & ~n39215;
  assign n39217 = ~pi72 & n39200;
  assign n39218 = n64196 & n39166;
  assign n39219 = n39167 & ~n39170;
  assign n39220 = n2728 & ~n39170;
  assign n39221 = n39196 & n39220;
  assign n39222 = n39218 & n39219;
  assign n39223 = ~n39217 & ~n64608;
  assign n39224 = ~pi44 & ~n39223;
  assign n39225 = ~pi72 & n39191;
  assign n39226 = ~pi101 & n64609;
  assign n39227 = n2825 & n39226;
  assign n39228 = ~pi113 & n39227;
  assign n39229 = ~pi116 & n39228;
  assign n39230 = n2827 & n39227;
  assign n39231 = ~pi42 & ~n64610;
  assign n39232 = ~n39009 & ~n39231;
  assign n39233 = ~n39216 & n39232;
  assign n39234 = ~pi115 & ~n39233;
  assign n39235 = ~pi228 & ~n39162;
  assign n39236 = ~n39234 & n39235;
  assign n39237 = ~pi39 & ~n39236;
  assign n39238 = ~n39165 & n39237;
  assign n39239 = pi287 & n62380;
  assign n39240 = n2814 & n39239;
  assign n39241 = ~pi189 & n39240;
  assign n39242 = ~n38991 & ~n39241;
  assign n39243 = pi199 & ~n39242;
  assign n39244 = pi200 & ~n39242;
  assign n39245 = pi232 & ~n39244;
  assign n39246 = ~pi299 & n39245;
  assign n39247 = n35103 & ~n39244;
  assign n39248 = pi232 & ~n39243;
  assign n39249 = ~n39244 & n39248;
  assign n39250 = ~n39243 & n39245;
  assign n39251 = ~pi299 & n64612;
  assign n39252 = ~n39243 & n64611;
  assign n39253 = n32363 & n39239;
  assign n39254 = n35283 & ~n39083;
  assign n39255 = ~n39253 & n39254;
  assign n39256 = pi72 & ~pi232;
  assign n39257 = pi299 & ~n39256;
  assign n39258 = n38989 & ~n39257;
  assign n39259 = ~n38995 & n39258;
  assign n39260 = ~n39255 & ~n39259;
  assign n39261 = ~n64613 & n39260;
  assign n39262 = pi39 & ~n39261;
  assign n39263 = ~n39238 & ~n39262;
  assign n39264 = n2766 & ~n39263;
  assign n39265 = n2993 & n39044;
  assign n39266 = n2993 & n39045;
  assign n39267 = ~pi44 & n39265;
  assign n39268 = n2993 & n39047;
  assign n39269 = n2826 & n64614;
  assign n39270 = ~pi113 & n64615;
  assign n39271 = ~pi116 & n39270;
  assign n39272 = n2827 & n64615;
  assign n39273 = ~pi72 & ~n2993;
  assign n39274 = ~pi72 & ~n39052;
  assign n39275 = ~n39273 & ~n39274;
  assign n39276 = ~pi72 & ~n64616;
  assign n39277 = pi42 & ~n64617;
  assign n39278 = ~pi114 & ~n39022;
  assign n39279 = ~pi114 & ~n39277;
  assign n39280 = ~n39022 & n39279;
  assign n39281 = ~n39277 & n39278;
  assign n39282 = n39010 & ~n64618;
  assign n39283 = n39008 & ~n39282;
  assign n39284 = ~n39037 & ~n39283;
  assign n39285 = ~pi39 & ~n39284;
  assign n39286 = ~n39087 & ~n39285;
  assign n39287 = n30855 & ~n39286;
  assign n39288 = ~n38987 & ~n39086;
  assign n39289 = pi38 & ~n39288;
  assign n39290 = ~n39003 & n39289;
  assign n39291 = ~pi87 & ~n39289;
  assign n39292 = pi38 & ~n39003;
  assign n39293 = ~pi87 & ~n39292;
  assign n39294 = ~n39291 & ~n39293;
  assign n39295 = ~pi75 & ~n39294;
  assign n39296 = n6795 & ~n39290;
  assign n39297 = ~n39287 & n64619;
  assign n39298 = ~n39264 & n39297;
  assign n39299 = ~n39088 & ~n39298;
  assign n39300 = ~n39287 & ~n39294;
  assign n39301 = ~n39264 & n39300;
  assign n39302 = n39077 & ~n39087;
  assign n39303 = n39078 & ~n39087;
  assign n39304 = ~n64596 & n39302;
  assign n39305 = ~pi75 & ~n64620;
  assign n39306 = ~n39301 & n39305;
  assign n39307 = ~n39042 & ~n39087;
  assign n39308 = pi75 & ~n39307;
  assign n39309 = n2580 & ~n39308;
  assign n39310 = ~n39306 & n39309;
  assign n39311 = n2580 & ~n39299;
  assign n39312 = n39005 & ~n64621;
  assign n39313 = ~pi299 & n39248;
  assign n39314 = n35103 & ~n39243;
  assign n39315 = ~n39255 & ~n39258;
  assign n39316 = ~n64622 & n39315;
  assign n39317 = pi39 & ~n39316;
  assign n39318 = ~n39238 & ~n39317;
  assign n39319 = n2766 & ~n39318;
  assign n39320 = ~n39086 & ~n39285;
  assign n39321 = n30855 & ~n39320;
  assign n39322 = n39291 & ~n39321;
  assign n39323 = ~n39319 & n39322;
  assign n39324 = n39078 & ~n39086;
  assign n39325 = ~pi75 & ~n39324;
  assign n39326 = ~n39323 & n39325;
  assign n39327 = ~n39042 & ~n39086;
  assign n39328 = pi75 & ~n39327;
  assign n39329 = n2580 & ~n39328;
  assign n39330 = ~n39326 & n39329;
  assign n39331 = ~n39323 & ~n39324;
  assign n39332 = ~pi75 & ~n39331;
  assign n39333 = n39043 & ~n39086;
  assign n39334 = ~n38985 & ~n39333;
  assign n39335 = ~n39332 & n39334;
  assign n39336 = ~n2580 & ~n38985;
  assign n39337 = ~n39335 & ~n39336;
  assign n39338 = ~n38985 & ~n39330;
  assign n39339 = ~n39312 & ~n39336;
  assign n39340 = ~n39335 & n39339;
  assign n39341 = ~n39312 & n64623;
  assign n39342 = pi212 & pi214;
  assign n39343 = pi211 & pi214;
  assign n39344 = pi212 & n39343;
  assign n39345 = pi211 & n39342;
  assign n39346 = ~pi219 & ~n64625;
  assign n39347 = ~n2580 & n39288;
  assign n39348 = ~n39346 & ~n39347;
  assign n39349 = ~n64624 & n39348;
  assign n39350 = ~n39002 & ~n39080;
  assign n39351 = ~n38990 & ~n38997;
  assign n39352 = ~n64612 & ~n39351;
  assign n39353 = pi39 & ~n39352;
  assign n39354 = ~n39238 & ~n39353;
  assign n39355 = n2766 & ~n39354;
  assign n39356 = ~n39002 & ~n39285;
  assign n39357 = n30855 & ~n39356;
  assign n39358 = n6795 & ~n39292;
  assign n39359 = ~n39357 & n39358;
  assign n39360 = ~n39355 & n39359;
  assign n39361 = n39293 & ~n39357;
  assign n39362 = ~n39355 & n39361;
  assign n39363 = ~n39002 & n39078;
  assign n39364 = ~n39362 & ~n39363;
  assign n39365 = ~pi75 & ~n39364;
  assign n39366 = ~n39002 & n39043;
  assign n39367 = ~n39365 & ~n39366;
  assign n39368 = ~n39350 & ~n39360;
  assign n39369 = ~pi75 & ~n39363;
  assign n39370 = ~n39362 & n39369;
  assign n39371 = ~n39002 & ~n39042;
  assign n39372 = pi75 & ~n39371;
  assign n39373 = n2580 & ~n39372;
  assign n39374 = ~n39370 & n39373;
  assign n39375 = n2580 & ~n64626;
  assign n39376 = n39005 & ~n64627;
  assign n39377 = pi39 & ~n38994;
  assign n39378 = ~n39080 & ~n39377;
  assign n39379 = n38990 & ~n39248;
  assign n39380 = pi39 & ~n39379;
  assign n39381 = ~n39238 & ~n39380;
  assign n39382 = n2766 & ~n39381;
  assign n39383 = ~n39285 & ~n39377;
  assign n39384 = n30855 & ~n39383;
  assign n39385 = ~n38987 & ~n39377;
  assign n39386 = pi38 & ~n39385;
  assign n39387 = n6795 & ~n39386;
  assign n39388 = ~n39384 & n39387;
  assign n39389 = ~n39382 & n39388;
  assign n39390 = ~pi87 & ~n39386;
  assign n39391 = ~n39384 & n39390;
  assign n39392 = ~n39382 & n39391;
  assign n39393 = n39078 & ~n39377;
  assign n39394 = ~n39392 & ~n39393;
  assign n39395 = ~pi75 & ~n39394;
  assign n39396 = n39043 & ~n39377;
  assign n39397 = ~n39395 & ~n39396;
  assign n39398 = ~n39378 & ~n39389;
  assign n39399 = ~pi75 & ~n39393;
  assign n39400 = ~n39392 & n39399;
  assign n39401 = ~n39042 & ~n39377;
  assign n39402 = pi75 & ~n39401;
  assign n39403 = n2580 & ~n39402;
  assign n39404 = ~n39400 & n39403;
  assign n39405 = n2580 & ~n64628;
  assign n39406 = ~n2580 & n39385;
  assign n39407 = ~n38985 & ~n39406;
  assign n39408 = ~n64629 & n39407;
  assign n39409 = ~n39376 & ~n39408;
  assign n39410 = n39346 & ~n39409;
  assign n39411 = n62455 & ~n39410;
  assign n39412 = n62455 & ~n39349;
  assign n39413 = ~n39410 & n39412;
  assign n39414 = ~n39349 & n39411;
  assign n39415 = n39083 & ~n39346;
  assign n39416 = pi39 & ~n39415;
  assign n39417 = ~n62455 & ~n38987;
  assign n39418 = ~n39416 & n39417;
  assign n39419 = ~n64630 & ~n39418;
  assign n39420 = pi211 & ~n39342;
  assign n39421 = ~pi211 & ~pi219;
  assign n39422 = n39342 & n39421;
  assign n39423 = ~pi211 & pi219;
  assign n39424 = ~pi211 & ~n39342;
  assign n39425 = ~n64625 & ~n39424;
  assign n39426 = ~n39423 & n39425;
  assign n39427 = n39342 & ~n39421;
  assign n39428 = ~n39424 & ~n39427;
  assign n39429 = ~n39420 & ~n39422;
  assign n39430 = ~n2929 & ~n64603;
  assign n39431 = n2929 & ~n64601;
  assign n39432 = ~n39430 & ~n39431;
  assign n39433 = pi228 & ~n39432;
  assign n39434 = ~pi228 & ~n39227;
  assign n39435 = n2827 & ~n39434;
  assign n39436 = n2929 & n64602;
  assign n39437 = ~n2929 & n64604;
  assign n39438 = pi228 & ~n39437;
  assign n39439 = n2827 & n39432;
  assign n39440 = pi228 & ~n39439;
  assign n39441 = ~n39436 & n39438;
  assign n39442 = ~pi228 & ~n64610;
  assign n39443 = ~n64632 & ~n39442;
  assign n39444 = ~n39433 & n39435;
  assign n39445 = ~pi43 & ~n64633;
  assign n39446 = pi43 & ~pi72;
  assign n39447 = ~n62386 & ~n39446;
  assign n39448 = n62386 & ~n39445;
  assign n39449 = ~n39446 & ~n39448;
  assign n39450 = ~n39445 & ~n39447;
  assign n39451 = ~pi228 & ~n39215;
  assign n39452 = n2929 & ~n39119;
  assign n39453 = ~n2929 & ~n39147;
  assign n39454 = ~n39452 & ~n39453;
  assign n39455 = pi228 & ~n39454;
  assign n39456 = ~n39451 & ~n39455;
  assign n39457 = pi43 & n62386;
  assign n39458 = ~n39456 & n39457;
  assign n39459 = ~n64634 & ~n39458;
  assign n39460 = ~pi39 & ~n39459;
  assign n39461 = n38997 & ~n39245;
  assign n39462 = pi39 & ~n39461;
  assign n39463 = ~n39460 & ~n39462;
  assign n39464 = n2766 & ~n39463;
  assign n39465 = ~n2997 & ~n39446;
  assign n39466 = n62386 & n2929;
  assign n39467 = n39446 & ~n39466;
  assign n39468 = n2997 & ~n39467;
  assign n39469 = ~pi43 & pi52;
  assign n39470 = n64588 & n39469;
  assign n39471 = pi43 & ~n64617;
  assign n39472 = ~n39470 & ~n39471;
  assign n39473 = n39466 & ~n39472;
  assign n39474 = n39468 & ~n39473;
  assign n39475 = ~n39465 & ~n39474;
  assign n39476 = ~pi39 & ~n39475;
  assign n39477 = ~n39001 & ~n39476;
  assign n39478 = n30855 & ~n39477;
  assign n39479 = ~pi39 & ~n39446;
  assign n39480 = ~n39001 & ~n39479;
  assign n39481 = pi38 & ~n39480;
  assign n39482 = ~pi87 & ~n39481;
  assign n39483 = ~n39478 & n39482;
  assign n39484 = ~n39464 & n39483;
  assign n39485 = ~pi43 & n39060;
  assign n39486 = pi228 & n62387;
  assign n39487 = n39016 & n64635;
  assign n39488 = n2766 & n2830;
  assign n39489 = n39069 & n39488;
  assign n39490 = n2766 & n39487;
  assign n39491 = n2766 & n62386;
  assign n39492 = n2766 & n39055;
  assign n39493 = n2831 & n39492;
  assign n39494 = n64591 & n39491;
  assign n39495 = n39446 & ~n64637;
  assign n39496 = ~pi39 & ~n39495;
  assign n39497 = ~n64636 & n39496;
  assign n39498 = ~pi43 & ~n39016;
  assign n39499 = pi43 & ~n39274;
  assign n39500 = n39060 & ~n39499;
  assign n39501 = ~n39498 & n39500;
  assign n39502 = ~n39060 & n39446;
  assign n39503 = n62373 & ~n39502;
  assign n39504 = ~n39501 & n39503;
  assign n39505 = ~n2766 & n39479;
  assign n39506 = pi87 & ~n39505;
  assign n39507 = ~n39504 & n39506;
  assign n39508 = pi87 & ~n39497;
  assign n39509 = ~n39001 & n64638;
  assign n39510 = ~pi75 & ~n39509;
  assign n39511 = ~n39484 & n39510;
  assign n39512 = ~pi72 & ~n39031;
  assign n39513 = pi43 & n39512;
  assign n39514 = ~n39031 & n39446;
  assign n39515 = n62385 & n64588;
  assign n39516 = n39469 & n39515;
  assign n39517 = n62385 & n39470;
  assign n39518 = ~n64639 & ~n64640;
  assign n39519 = n39466 & ~n39518;
  assign n39520 = n39468 & ~n39519;
  assign n39521 = n62951 & ~n39465;
  assign n39522 = ~n39520 & n39521;
  assign n39523 = ~n62951 & n39446;
  assign n39524 = ~pi39 & ~n39523;
  assign n39525 = ~n39465 & ~n39520;
  assign n39526 = ~pi39 & ~n39525;
  assign n39527 = n62951 & ~n39526;
  assign n39528 = ~n62951 & ~n39479;
  assign n39529 = ~n39527 & ~n39528;
  assign n39530 = ~n39522 & n39524;
  assign n39531 = ~n39001 & ~n64641;
  assign n39532 = pi75 & ~n39531;
  assign n39533 = n2580 & ~n39532;
  assign n39534 = ~n39511 & n39533;
  assign n39535 = ~n2580 & n39480;
  assign n39536 = ~n38985 & ~n39535;
  assign n39537 = ~n39534 & n39536;
  assign n39538 = ~pi199 & ~pi200;
  assign n39539 = ~pi299 & ~n39538;
  assign n39540 = ~pi72 & ~n39539;
  assign n39541 = ~pi232 & ~n39540;
  assign n39542 = ~pi299 & ~n39541;
  assign n39543 = ~n39242 & n39538;
  assign n39544 = pi232 & ~n39543;
  assign n39545 = n39542 & ~n39544;
  assign n39546 = pi39 & ~n39545;
  assign n39547 = ~n39460 & ~n39546;
  assign n39548 = n2766 & ~n39547;
  assign n39549 = n38991 & n39538;
  assign n39550 = pi232 & ~n39549;
  assign n39551 = n39542 & ~n39550;
  assign n39552 = pi39 & ~n39551;
  assign n39553 = ~n39476 & ~n39552;
  assign n39554 = n30855 & ~n39553;
  assign n39555 = ~n39479 & ~n39552;
  assign n39556 = pi38 & ~n39555;
  assign n39557 = ~pi87 & ~n39556;
  assign n39558 = ~n39554 & n39557;
  assign n39559 = ~n39548 & n39558;
  assign n39560 = ~n62373 & ~n39555;
  assign n39561 = n64638 & ~n39560;
  assign n39562 = ~pi75 & ~n39561;
  assign n39563 = ~n39559 & n39562;
  assign n39564 = ~n64641 & ~n39552;
  assign n39565 = pi75 & ~n39564;
  assign n39566 = n2580 & ~n39565;
  assign n39567 = ~n39563 & n39566;
  assign n39568 = ~n2580 & n39555;
  assign n39569 = n38985 & ~n39568;
  assign n39570 = ~n39567 & n39569;
  assign n39571 = ~n39537 & ~n39570;
  assign n39572 = ~n64631 & ~n39571;
  assign n39573 = n38996 & ~n39257;
  assign n39574 = ~n39255 & ~n39573;
  assign n39575 = ~n64611 & n39574;
  assign n39576 = pi39 & ~n39575;
  assign n39577 = ~n39460 & ~n39576;
  assign n39578 = n2766 & ~n39577;
  assign n39579 = ~n39000 & n39085;
  assign n39580 = ~n39476 & ~n39579;
  assign n39581 = n30855 & ~n39580;
  assign n39582 = ~n39479 & ~n39579;
  assign n39583 = pi38 & ~n39582;
  assign n39584 = ~pi87 & ~n39583;
  assign n39585 = ~n39581 & n39584;
  assign n39586 = ~n39578 & n39585;
  assign n39587 = n64638 & ~n39579;
  assign n39588 = ~pi75 & ~n39587;
  assign n39589 = ~n39586 & n39588;
  assign n39590 = ~n64641 & ~n39579;
  assign n39591 = pi75 & ~n39590;
  assign n39592 = n2580 & ~n39591;
  assign n39593 = ~n39589 & n39592;
  assign n39594 = ~n2580 & n39582;
  assign n39595 = ~n38985 & ~n39594;
  assign n39596 = ~n39593 & n39595;
  assign n39597 = n35103 & ~n39543;
  assign n39598 = ~n39255 & ~n39541;
  assign n39599 = ~n39597 & n39598;
  assign n39600 = pi39 & ~n39599;
  assign n39601 = ~n39460 & ~n39600;
  assign n39602 = n2766 & ~n39601;
  assign n39603 = ~n39084 & n39552;
  assign n39604 = ~n39476 & ~n39603;
  assign n39605 = n30855 & ~n39604;
  assign n39606 = ~n39479 & ~n39603;
  assign n39607 = pi38 & ~n39606;
  assign n39608 = ~pi87 & ~n39607;
  assign n39609 = ~n39605 & n39608;
  assign n39610 = ~n39602 & n39609;
  assign n39611 = n64638 & ~n39603;
  assign n39612 = ~pi75 & ~n39611;
  assign n39613 = ~n39610 & n39612;
  assign n39614 = ~n64641 & ~n39603;
  assign n39615 = pi75 & ~n39614;
  assign n39616 = n2580 & ~n39615;
  assign n39617 = ~n39613 & n39616;
  assign n39618 = ~n2580 & n39606;
  assign n39619 = n38985 & ~n39618;
  assign n39620 = ~n39617 & n39619;
  assign n39621 = ~n39596 & ~n39620;
  assign n39622 = n64631 & ~n39621;
  assign n39623 = n62455 & ~n39622;
  assign n39624 = n62455 & ~n39572;
  assign n39625 = ~n39622 & n39624;
  assign n39626 = ~n39572 & n39623;
  assign n39627 = n39083 & n64631;
  assign n39628 = pi39 & ~n39627;
  assign n39629 = ~n62455 & ~n39479;
  assign n39630 = ~n39628 & n39629;
  assign n39631 = ~n64642 & ~n39630;
  assign n39632 = pi52 & n39454;
  assign n39633 = n2828 & n39432;
  assign n39634 = n62387 & ~n39633;
  assign n39635 = pi52 & n39119;
  assign n39636 = ~pi52 & n64602;
  assign n39637 = n39006 & ~n39636;
  assign n39638 = ~n39635 & n39637;
  assign n39639 = pi52 & n39147;
  assign n39640 = ~pi52 & n64604;
  assign n39641 = n39160 & ~n39640;
  assign n39642 = ~n39639 & n39641;
  assign n39643 = ~n39638 & ~n39642;
  assign n39644 = n2835 & ~n39643;
  assign n39645 = ~n39632 & n39634;
  assign n39646 = pi52 & ~pi72;
  assign n39647 = ~n62387 & ~n39646;
  assign n39648 = pi228 & ~n39647;
  assign n39649 = ~n64643 & n39648;
  assign n39650 = pi52 & n39215;
  assign n39651 = ~pi52 & n64610;
  assign n39652 = n2828 & n39227;
  assign n39653 = n62387 & ~n64644;
  assign n39654 = ~n39650 & n39653;
  assign n39655 = ~pi228 & ~n39647;
  assign n39656 = ~n39654 & n39655;
  assign n39657 = ~pi39 & ~n39656;
  assign n39658 = ~n39649 & n39657;
  assign n39659 = ~n39600 & ~n39658;
  assign n39660 = n2766 & ~n39659;
  assign n39661 = ~pi39 & ~n39646;
  assign n39662 = ~n39085 & ~n39661;
  assign n39663 = ~n39552 & ~n39661;
  assign n39664 = pi38 & ~n39663;
  assign n39665 = ~n39662 & n39664;
  assign n39666 = n2929 & n2997;
  assign n39667 = n2997 & n39006;
  assign n39668 = n2835 & n39667;
  assign n39669 = n62387 & n39666;
  assign n39670 = n2993 & n64645;
  assign n39671 = n64616 & n64645;
  assign n39672 = n39052 & n39670;
  assign n39673 = n39646 & ~n64646;
  assign n39674 = ~pi39 & ~n39673;
  assign n39675 = ~n39603 & ~n39674;
  assign n39676 = n30855 & ~n39675;
  assign n39677 = ~n39665 & ~n39676;
  assign n39678 = ~n39660 & n39677;
  assign n39679 = ~pi87 & ~n39678;
  assign n39680 = n2835 & n39055;
  assign n39681 = n2830 & n64592;
  assign n39682 = n39646 & ~n64647;
  assign n39683 = n2838 & n39069;
  assign n39684 = ~pi52 & n39487;
  assign n39685 = ~pi52 & n39016;
  assign n39686 = pi52 & n39274;
  assign n39687 = ~n39685 & ~n39686;
  assign n39688 = n64635 & ~n39687;
  assign n39689 = ~n64635 & n39646;
  assign n39690 = ~n39688 & ~n39689;
  assign n39691 = ~n39682 & ~n64648;
  assign n39692 = ~pi39 & n64649;
  assign n39693 = n2766 & ~n39603;
  assign n39694 = ~n39692 & n39693;
  assign n39695 = ~n2766 & n39662;
  assign n39696 = pi87 & ~n39695;
  assign n39697 = ~n2766 & n39663;
  assign n39698 = n39696 & ~n39697;
  assign n39699 = ~n39694 & n39698;
  assign n39700 = ~n38985 & ~n39699;
  assign n39701 = ~n39679 & n39700;
  assign n39702 = ~pi39 & pi100;
  assign n39703 = pi100 & n2764;
  assign n39704 = ~pi38 & n39702;
  assign n39705 = n64646 & n64650;
  assign n39706 = ~n39255 & n39257;
  assign n39707 = pi39 & ~n39706;
  assign n39708 = n2766 & ~n39707;
  assign n39709 = ~n39658 & n39708;
  assign n39710 = ~n39695 & ~n39709;
  assign n39711 = ~n39658 & ~n39707;
  assign n39712 = n2766 & ~n39711;
  assign n39713 = pi38 & ~n39662;
  assign n39714 = ~n39085 & ~n39674;
  assign n39715 = n30855 & ~n39714;
  assign n39716 = ~n39713 & ~n39715;
  assign n39717 = ~n39712 & n39716;
  assign n39718 = ~n39705 & ~n39710;
  assign n39719 = ~pi87 & ~n64651;
  assign n39720 = n2766 & ~n39085;
  assign n39721 = ~n39692 & n39720;
  assign n39722 = n39696 & ~n39721;
  assign n39723 = n38985 & ~n39722;
  assign n39724 = ~n39719 & n39723;
  assign n39725 = ~pi75 & ~n39724;
  assign n39726 = ~n39701 & n39725;
  assign n39727 = n62951 & n64645;
  assign n39728 = n39031 & n64645;
  assign n39729 = n62951 & n39728;
  assign n39730 = n39031 & n39727;
  assign n39731 = n39646 & ~n64652;
  assign n39732 = ~pi39 & n39646;
  assign n39733 = ~n64652 & n39732;
  assign n39734 = ~pi39 & ~n39733;
  assign n39735 = ~pi39 & ~n39731;
  assign n39736 = ~n38985 & n39551;
  assign n39737 = n39085 & ~n39736;
  assign n39738 = ~n64653 & ~n39737;
  assign n39739 = pi75 & ~n39738;
  assign n39740 = n2580 & ~n39739;
  assign n39741 = ~n39701 & ~n39724;
  assign n39742 = ~pi75 & ~n39741;
  assign n39743 = ~n38985 & n39603;
  assign n39744 = n38985 & n39085;
  assign n39745 = pi75 & ~n39744;
  assign n39746 = ~n39743 & n39745;
  assign n39747 = pi75 & ~n39737;
  assign n39748 = ~n64653 & n64654;
  assign n39749 = ~n39742 & ~n39748;
  assign n39750 = n2580 & ~n39749;
  assign n39751 = ~n39726 & n39740;
  assign n39752 = ~pi219 & n39424;
  assign n39753 = ~n39342 & n39421;
  assign n39754 = ~n2580 & n39662;
  assign n39755 = n64656 & ~n39754;
  assign n39756 = ~n64655 & n39755;
  assign n39757 = n2766 & n64649;
  assign n39758 = pi87 & ~n38958;
  assign n39759 = ~n2766 & ~n39732;
  assign n39760 = n39758 & ~n39759;
  assign n39761 = pi38 & ~n39732;
  assign n39762 = ~pi38 & n64649;
  assign n39763 = ~n39761 & ~n39762;
  assign n39764 = ~pi100 & ~n39763;
  assign n39765 = pi100 & ~n39732;
  assign n39766 = n39758 & ~n39765;
  assign n39767 = ~n39764 & n39766;
  assign n39768 = ~n39757 & n39760;
  assign n39769 = ~pi100 & n39658;
  assign n39770 = pi100 & ~n39673;
  assign n39771 = ~pi39 & ~n39770;
  assign n39772 = ~n39769 & n39771;
  assign n39773 = ~pi38 & ~n39772;
  assign n39774 = ~pi87 & ~n39761;
  assign n39775 = ~n39773 & n39774;
  assign n39776 = ~n64657 & ~n39775;
  assign n39777 = ~pi75 & ~n39776;
  assign n39778 = pi75 & n39732;
  assign n39779 = ~pi39 & pi75;
  assign n39780 = n39731 & n39779;
  assign n39781 = pi75 & n39733;
  assign n39782 = ~n64652 & n39778;
  assign n39783 = n2580 & ~n64658;
  assign n39784 = ~n39777 & n39783;
  assign n39785 = ~n2580 & ~n39732;
  assign n39786 = n38985 & ~n39785;
  assign n39787 = ~n39784 & n39786;
  assign n39788 = ~n39546 & ~n39658;
  assign n39789 = n2766 & ~n39788;
  assign n39790 = ~n39552 & ~n39674;
  assign n39791 = n30855 & ~n39790;
  assign n39792 = ~pi87 & ~n39664;
  assign n39793 = ~n39791 & n39792;
  assign n39794 = ~n39789 & n39793;
  assign n39795 = n2766 & ~n39552;
  assign n39796 = ~n39692 & n39795;
  assign n39797 = ~n39697 & ~n39796;
  assign n39798 = pi87 & ~n39797;
  assign n39799 = ~pi75 & ~n39798;
  assign n39800 = ~n39794 & n39799;
  assign n39801 = n2580 & ~n38985;
  assign n39802 = n39646 & ~n39728;
  assign n39803 = ~pi39 & ~n39802;
  assign n39804 = ~pi87 & n39795;
  assign n39805 = n62951 & ~n39552;
  assign n39806 = ~n39803 & n64659;
  assign n39807 = ~n62951 & n39663;
  assign n39808 = pi75 & ~n39807;
  assign n39809 = ~n39806 & n39808;
  assign n39810 = n39801 & ~n39809;
  assign n39811 = ~n39794 & ~n39798;
  assign n39812 = ~pi75 & ~n39811;
  assign n39813 = pi75 & ~n39552;
  assign n39814 = ~n64653 & n39813;
  assign n39815 = ~n39812 & ~n39814;
  assign n39816 = n39801 & ~n39815;
  assign n39817 = ~n39800 & n39810;
  assign n39818 = ~n64656 & ~n64660;
  assign n39819 = ~n39787 & n39818;
  assign n39820 = ~n39756 & ~n39819;
  assign n39821 = n39336 & n39663;
  assign n39822 = n62455 & ~n39821;
  assign n39823 = ~n39787 & ~n64660;
  assign n39824 = ~n64656 & ~n39823;
  assign n39825 = n2580 & ~n39748;
  assign n39826 = ~n39742 & n39825;
  assign n39827 = ~n2580 & ~n39662;
  assign n39828 = n64656 & ~n39827;
  assign n39829 = ~n39826 & n39828;
  assign n39830 = n39822 & ~n39829;
  assign n39831 = ~n39824 & n39830;
  assign n39832 = ~n39820 & n39822;
  assign n39833 = pi39 & n64656;
  assign n39834 = n39083 & n39833;
  assign n39835 = ~n62455 & ~n39732;
  assign n39836 = ~n39834 & n39835;
  assign po210 = ~n64661 & ~n39836;
  assign n39838 = n63888 & n27583;
  assign n39839 = pi216 & ~pi221;
  assign n39840 = n2959 & n39839;
  assign n39841 = n35099 & n39840;
  assign n39842 = n2979 & n28811;
  assign n39843 = n35096 & n39842;
  assign n39844 = ~n39841 & ~n39843;
  assign po226 = n39838 & ~n39844;
  assign n39846 = n35370 & n38940;
  assign n39847 = ~pi58 & n2857;
  assign n39848 = ~n39846 & ~n39847;
  assign n39849 = n62395 & n64196;
  assign n39850 = ~n39848 & n39849;
  assign n39851 = pi24 & n2783;
  assign n39852 = n62366 & ~n62395;
  assign n39853 = pi24 & ~n62395;
  assign n39854 = n62379 & n39853;
  assign n39855 = pi24 & n2715;
  assign n39856 = ~n62395 & n39855;
  assign n39857 = n35400 & n39856;
  assign n39858 = n39851 & n39852;
  assign n39859 = n2857 & n64662;
  assign n39860 = ~pi39 & ~n39859;
  assign n39861 = ~n39850 & n39860;
  assign n39862 = n63888 & ~n39861;
  assign po249 = n2990 & n39862;
  assign n39864 = n64089 & n30722;
  assign n39865 = ~pi82 & n2593;
  assign n39866 = ~pi84 & pi104;
  assign n39867 = n30652 & n39866;
  assign n39868 = n38233 & n39867;
  assign n39869 = n39865 & n39868;
  assign n39870 = ~pi36 & ~n39869;
  assign n39871 = n62347 & n6810;
  assign n39872 = n2621 & n6811;
  assign n39873 = ~pi67 & ~pi103;
  assign n39874 = n2587 & n39873;
  assign n39875 = ~pi98 & n39874;
  assign n39876 = n64663 & n39875;
  assign n39877 = ~n39870 & n39876;
  assign n39878 = ~pi36 & n39877;
  assign n39879 = ~pi88 & ~n39878;
  assign n39880 = n6875 & ~n39879;
  assign n39881 = n2655 & n6921;
  assign n39882 = n39880 & n39881;
  assign n39883 = ~pi91 & ~n6846;
  assign n39884 = ~n33889 & n39877;
  assign n39885 = ~pi88 & ~n39884;
  assign n39886 = n2655 & ~n39885;
  assign n39887 = n6875 & n39886;
  assign n39888 = ~n2582 & n39887;
  assign n39889 = n39883 & ~n39888;
  assign n39890 = ~n39882 & n39883;
  assign n39891 = ~n39888 & n39890;
  assign n39892 = ~n39882 & n39889;
  assign n39893 = n39864 & ~n64664;
  assign n39894 = ~pi72 & ~n39893;
  assign n39895 = n30619 & ~n39894;
  assign n39896 = n33976 & ~n39895;
  assign n39897 = n2852 & n64089;
  assign n39898 = n30619 & n39897;
  assign n39899 = ~n39848 & n39897;
  assign n39900 = n30619 & n39899;
  assign n39901 = ~n39848 & n39898;
  assign n39902 = ~n30823 & ~n64665;
  assign n39903 = pi1093 & ~n39902;
  assign n39904 = n39864 & n39887;
  assign n39905 = ~n2852 & n39904;
  assign n39906 = n39864 & ~n39883;
  assign n39907 = ~pi72 & ~n39906;
  assign n39908 = ~n38259 & n39907;
  assign n39909 = ~n38259 & ~n39905;
  assign n39910 = n39907 & n39909;
  assign n39911 = ~n39905 & n39908;
  assign n39912 = n30619 & ~n64666;
  assign n39913 = ~n39903 & ~n39912;
  assign n39914 = ~n39904 & n39907;
  assign n39915 = n30619 & ~n39914;
  assign n39916 = n6899 & ~n39915;
  assign n39917 = ~n39913 & ~n39916;
  assign n39918 = ~n39896 & n39917;
  assign n39919 = ~pi39 & ~n39918;
  assign n39920 = n38956 & ~n39919;
  assign n39921 = n30874 & n34137;
  assign n39922 = pi137 & n39921;
  assign n39923 = pi129 & n62380;
  assign n39924 = ~pi137 & pi252;
  assign n39925 = pi683 & n34975;
  assign n39926 = pi252 & ~n39925;
  assign n39927 = pi252 & ~n2843;
  assign n39928 = ~n39925 & n39927;
  assign n39929 = ~n2843 & n39926;
  assign n39930 = ~n64105 & ~n64667;
  assign n39931 = ~n2816 & ~n39930;
  assign n39932 = ~n39924 & ~n39931;
  assign n39933 = ~n64105 & ~n34974;
  assign n39934 = ~n64105 & ~n39933;
  assign n39935 = ~n64105 & n34974;
  assign n39936 = ~n64667 & n64668;
  assign n39937 = ~n39932 & ~n39936;
  assign n39938 = n39923 & ~n39937;
  assign n39939 = ~n39922 & ~n39938;
  assign n39940 = n64650 & ~n39939;
  assign n39941 = ~pi90 & n32076;
  assign n39942 = ~pi93 & ~n39941;
  assign n39943 = ~n2661 & ~n39942;
  assign n39944 = ~pi35 & ~n39943;
  assign n39945 = pi35 & ~n64295;
  assign n39946 = n62376 & ~n39945;
  assign n39947 = ~n39944 & n39946;
  assign n39948 = ~pi32 & n39947;
  assign n39949 = n31079 & n64296;
  assign n39950 = pi32 & ~pi93;
  assign n39951 = n39949 & n39950;
  assign n39952 = n2674 & n39951;
  assign n39953 = ~n39948 & ~n39952;
  assign n39954 = ~pi95 & n64148;
  assign n39955 = ~n39953 & n39954;
  assign n39956 = ~n64148 & ~n39944;
  assign n39957 = n2929 & n2993;
  assign n39958 = ~pi122 & n62395;
  assign n39959 = ~n3318 & n64669;
  assign n39960 = ~pi122 & ~po740;
  assign n39961 = n3318 & n39960;
  assign n39962 = ~n3318 & ~n64669;
  assign n39963 = n3318 & ~n39960;
  assign n39964 = ~n39962 & ~n39963;
  assign n39965 = ~n39959 & ~n39961;
  assign n39966 = ~n39956 & ~n64670;
  assign n39967 = pi76 & ~pi84;
  assign n39968 = n2598 & n39967;
  assign n39969 = n6809 & n38231;
  assign n39970 = ~pi73 & pi76;
  assign n39971 = n30652 & n39970;
  assign n39972 = n31458 & n38231;
  assign n39973 = n39971 & n39972;
  assign n39974 = n39968 & n39969;
  assign n39975 = n2587 & n2616;
  assign n39976 = n38885 & n39975;
  assign n39977 = n64671 & n39976;
  assign n39978 = ~pi45 & ~pi48;
  assign n39979 = ~pi61 & ~pi104;
  assign n39980 = n39978 & n39979;
  assign n39981 = n6811 & n39980;
  assign n39982 = ~pi103 & n2590;
  assign n39983 = n38886 & n39982;
  assign n39984 = n39981 & n39983;
  assign n39985 = n39977 & n39984;
  assign n39986 = n2638 & n39985;
  assign n39987 = n62355 & n2694;
  assign n39988 = n62355 & n39986;
  assign n39989 = n62356 & n39985;
  assign n39990 = n2694 & n64672;
  assign n39991 = n39986 & n39987;
  assign n39992 = n39944 & ~n64673;
  assign n39993 = ~pi137 & n64148;
  assign n39994 = n2727 & ~n39993;
  assign n39995 = n39946 & n39994;
  assign n39996 = ~n39992 & n39995;
  assign n39997 = ~n3318 & ~n39993;
  assign n39998 = n64669 & n39997;
  assign n39999 = n3318 & ~n39993;
  assign n40000 = n39960 & n39999;
  assign n40001 = ~n39998 & ~n40000;
  assign n40002 = n39944 & ~n64670;
  assign n40003 = ~n64148 & ~n40002;
  assign n40004 = pi137 & n64670;
  assign n40005 = ~n40003 & ~n40004;
  assign n40006 = ~n39956 & n40001;
  assign n40007 = n2727 & n39946;
  assign n40008 = ~n39992 & n40007;
  assign n40009 = ~n64674 & n40008;
  assign n40010 = ~n39966 & n39996;
  assign n40011 = ~n6864 & ~n39947;
  assign n40012 = pi1082 & n2727;
  assign n40013 = ~n40011 & n40012;
  assign n40014 = ~pi38 & ~n40013;
  assign n40015 = ~pi38 & ~n64675;
  assign n40016 = ~n40013 & n40015;
  assign n40017 = ~n64675 & n40014;
  assign n40018 = ~n39955 & n64676;
  assign n40019 = pi38 & ~n62384;
  assign n40020 = ~pi39 & ~pi100;
  assign n40021 = ~n40019 & n40020;
  assign n40022 = ~n40018 & n40021;
  assign n40023 = ~n39940 & ~n40022;
  assign n40024 = n6795 & ~n40023;
  assign n40025 = pi75 & ~pi100;
  assign n40026 = n30571 & n40025;
  assign n40027 = ~pi24 & n40026;
  assign n40028 = pi252 & ~n34974;
  assign n40029 = pi137 & n38261;
  assign n40030 = ~n30877 & n40029;
  assign n40031 = ~n40028 & ~n40030;
  assign n40032 = n40027 & ~n40031;
  assign n40033 = n40026 & ~n40031;
  assign n40034 = n62384 & n40033;
  assign n40035 = n62380 & n40032;
  assign n40036 = ~n40024 & ~n64677;
  assign n40037 = ~pi92 & ~n40036;
  assign n40038 = ~pi54 & ~n40037;
  assign n40039 = ~pi24 & n30894;
  assign n40040 = pi54 & ~n40039;
  assign n40041 = n64497 & ~n40040;
  assign n40042 = ~n40038 & n40041;
  assign n40043 = ~pi59 & ~n40042;
  assign n40044 = n3470 & n64082;
  assign n40045 = n62384 & n40044;
  assign n40046 = ~pi55 & n40045;
  assign n40047 = pi59 & ~n40046;
  assign n40048 = ~pi57 & ~n40047;
  assign po193 = ~n40043 & n40048;
  assign n40050 = n62400 & n39840;
  assign n40051 = n62402 & n39842;
  assign n40052 = ~n40050 & ~n40051;
  assign po244 = n39838 & ~n40052;
  assign n40054 = ~pi979 & ~pi984;
  assign n40055 = pi1001 & n40054;
  assign n40056 = n6957 & n40055;
  assign n40057 = ~n2583 & n40056;
  assign n40058 = n2933 & n40057;
  assign n40059 = ~pi252 & ~n40058;
  assign n40060 = pi1092 & ~pi1093;
  assign n40061 = ~n40059 & n40060;
  assign n40062 = n30820 & ~n40061;
  assign n40063 = ~n2953 & ~n40062;
  assign n40064 = pi252 & pi1092;
  assign n40065 = ~pi1093 & n40064;
  assign n40066 = n2953 & n40065;
  assign n40067 = ~n40063 & ~n40066;
  assign n40068 = ~n2971 & ~n40067;
  assign n40069 = ~n2909 & n40065;
  assign n40070 = n2909 & ~n40062;
  assign n40071 = ~n40069 & ~n40070;
  assign n40072 = n2971 & ~n40071;
  assign n40073 = ~pi299 & ~n40072;
  assign n40074 = ~pi299 & ~n40068;
  assign n40075 = ~n40072 & n40074;
  assign n40076 = ~n40068 & n40073;
  assign n40077 = n62393 & ~n40071;
  assign n40078 = ~n62393 & ~n40067;
  assign n40079 = pi299 & ~n40078;
  assign n40080 = pi299 & ~n40077;
  assign n40081 = ~n40078 & n40080;
  assign n40082 = ~n40077 & n40079;
  assign n40083 = n39838 & ~n64679;
  assign n40084 = n39838 & ~n64678;
  assign n40085 = ~n64679 & n40084;
  assign n40086 = ~n64678 & n40083;
  assign n40087 = ~n39838 & n40065;
  assign n40088 = ~n5530 & ~n40087;
  assign n40089 = ~n64680 & n40088;
  assign n40090 = ~n30831 & ~n30841;
  assign n40091 = n27583 & n40056;
  assign n40092 = n27338 & n40091;
  assign n40093 = n64298 & n40092;
  assign n40094 = ~n40090 & n40093;
  assign n40095 = n2933 & n40094;
  assign n40096 = ~pi252 & ~n40095;
  assign n40097 = ~pi57 & pi1092;
  assign n40098 = ~n40096 & n40097;
  assign n40099 = pi57 & n40064;
  assign n40100 = n5530 & ~n40099;
  assign n40101 = ~n40098 & n40100;
  assign po409 = ~n40089 & ~n40101;
  assign n40103 = n2579 & n64498;
  assign n40104 = ~n64105 & n40028;
  assign n40105 = n39923 & n40104;
  assign n40106 = ~n39921 & ~n40105;
  assign n40107 = ~pi137 & n64650;
  assign n40108 = ~pi137 & n39921;
  assign n40109 = ~n64105 & n39924;
  assign n40110 = n39924 & n39933;
  assign n40111 = ~n34974 & n40109;
  assign n40112 = n39923 & n64681;
  assign n40113 = ~n40108 & ~n40112;
  assign n40114 = n64650 & ~n40113;
  assign n40115 = ~n40106 & n40107;
  assign n40116 = ~n3318 & n38261;
  assign n40117 = ~pi137 & ~n40116;
  assign n40118 = n2638 & n31450;
  assign n40119 = ~pi93 & n62355;
  assign n40120 = n40118 & n40119;
  assign n40121 = n39949 & n40120;
  assign n40122 = ~n40117 & ~n40121;
  assign n40123 = ~pi24 & n31450;
  assign n40124 = ~n39985 & ~n40123;
  assign n40125 = ~pi40 & n62775;
  assign n40126 = ~n31450 & ~n39985;
  assign n40127 = n62356 & ~n40126;
  assign n40128 = ~pi24 & ~n40127;
  assign n40129 = pi24 & ~n64672;
  assign n40130 = ~pi40 & n62768;
  assign n40131 = n2695 & n62376;
  assign n40132 = ~n40129 & n64683;
  assign n40133 = ~n40128 & n40132;
  assign n40134 = ~n40124 & n40125;
  assign n40135 = n40117 & ~n64684;
  assign n40136 = ~pi32 & ~n40135;
  assign n40137 = ~pi32 & ~n40122;
  assign n40138 = ~n40135 & n40137;
  assign n40139 = ~n40117 & n40121;
  assign n40140 = ~pi137 & n2695;
  assign n40141 = n62376 & n40140;
  assign n40142 = ~n40116 & n40141;
  assign n40143 = ~n40129 & n40142;
  assign n40144 = ~n40128 & n40143;
  assign n40145 = ~n40139 & ~n40144;
  assign n40146 = ~pi32 & ~n40145;
  assign n40147 = ~n40122 & n40136;
  assign n40148 = ~pi24 & ~pi841;
  assign n40149 = pi32 & ~n40148;
  assign n40150 = n33956 & n40149;
  assign n40151 = ~n64685 & ~n40150;
  assign n40152 = n64148 & ~n40151;
  assign n40153 = ~pi32 & ~n40121;
  assign n40154 = ~n64148 & ~n33954;
  assign n40155 = ~n40153 & n40154;
  assign n40156 = ~n40152 & ~n40155;
  assign n40157 = ~pi95 & n62373;
  assign n40158 = ~n40156 & n40157;
  assign n40159 = ~n64682 & ~n40158;
  assign n40160 = n6795 & ~n40159;
  assign n40161 = n62384 & n38261;
  assign n40162 = ~pi137 & n40026;
  assign n40163 = ~n30877 & n40162;
  assign n40164 = ~n40028 & n40163;
  assign n40165 = n40161 & n40164;
  assign n40166 = ~n40160 & ~n40165;
  assign po190 = n40103 & ~n40166;
  assign n40168 = pi39 & n38872;
  assign n40169 = n64325 & n40168;
  assign n40170 = n38872 & n39838;
  assign n40171 = ~n64580 & n64686;
  assign n40172 = ~n64579 & n64686;
  assign n40173 = ~n64580 & n40172;
  assign n40174 = ~n64579 & n40171;
  assign n40175 = ~n30598 & ~n30903;
  assign n40176 = pi93 & ~n2659;
  assign n40177 = ~n33939 & ~n40176;
  assign n40178 = pi58 & ~n2658;
  assign n40179 = ~n30627 & ~n40178;
  assign n40180 = n2586 & ~n2857;
  assign n40181 = ~pi91 & ~n33929;
  assign n40182 = n6849 & ~n33929;
  assign n40183 = ~n6847 & n40181;
  assign n40184 = ~pi81 & ~n33912;
  assign n40185 = n30706 & ~n40184;
  assign n40186 = n2611 & ~n40185;
  assign n40187 = n33918 & ~n40186;
  assign n40188 = n30645 & ~n40187;
  assign n40189 = n30641 & ~n40188;
  assign n40190 = n30639 & ~n40189;
  assign n40191 = ~n30637 & ~n40190;
  assign n40192 = ~pi86 & ~n40191;
  assign n40193 = n30715 & ~n40192;
  assign n40194 = n33873 & ~n40193;
  assign n40195 = ~n30937 & ~n40194;
  assign n40196 = ~pi108 & ~n40195;
  assign n40197 = n33870 & ~n40196;
  assign n40198 = n30750 & ~n40197;
  assign n40199 = ~n30748 & ~n40198;
  assign n40200 = n2866 & ~n40199;
  assign n40201 = n64688 & ~n40200;
  assign n40202 = n40180 & ~n40201;
  assign n40203 = n40179 & ~n40202;
  assign n40204 = n2719 & ~n40203;
  assign n40205 = n40177 & ~n40204;
  assign n40206 = ~pi70 & ~n40205;
  assign n40207 = ~n30620 & ~n40206;
  assign n40208 = ~pi51 & ~n40207;
  assign n40209 = n2733 & ~n40208;
  assign n40210 = n33868 & ~n40209;
  assign n40211 = n33860 & ~n40210;
  assign n40212 = ~pi1082 & n6864;
  assign n40213 = ~pi32 & ~n40212;
  assign n40214 = ~n40211 & n40213;
  assign n40215 = ~n33957 & ~n40214;
  assign n40216 = ~pi95 & ~n40215;
  assign n40217 = ~n33962 & ~n40216;
  assign n40218 = ~pi39 & ~n40217;
  assign n40219 = pi39 & ~n62380;
  assign n40220 = n2582 & n64298;
  assign n40221 = n2938 & n40220;
  assign n40222 = ~n40090 & n40221;
  assign n40223 = n6956 & n40168;
  assign n40224 = ~n40222 & n40223;
  assign n40225 = ~n40219 & ~n40224;
  assign n40226 = ~n40218 & n40225;
  assign n40227 = ~pi38 & ~n40226;
  assign n40228 = n33858 & ~n40227;
  assign n40229 = ~pi87 & ~n30856;
  assign n40230 = ~n40228 & n40229;
  assign n40231 = ~n34033 & ~n40230;
  assign n40232 = n6793 & ~n40231;
  assign n40233 = n30605 & ~n40232;
  assign n40234 = ~pi54 & ~n40233;
  assign n40235 = ~n30895 & ~n40234;
  assign n40236 = n34040 & ~n40235;
  assign n40237 = n40175 & ~n40236;
  assign n40238 = ~pi56 & ~n40237;
  assign n40239 = ~n34043 & ~n40238;
  assign n40240 = ~pi62 & ~n40239;
  assign n40241 = ~n34048 & ~n40240;
  assign n40242 = n3472 & ~n40241;
  assign po389 = n30591 & ~n40242;
  assign n40244 = ~pi41 & ~pi72;
  assign n40245 = ~n2997 & ~n40244;
  assign n40246 = ~n2929 & n40244;
  assign n40247 = n2997 & ~n40246;
  assign n40248 = n62385 & n39014;
  assign n40249 = pi41 & ~n40248;
  assign n40250 = ~pi41 & pi72;
  assign n40251 = n2929 & ~n40250;
  assign n40252 = ~pi99 & n62388;
  assign n40253 = n39028 & n39094;
  assign n40254 = ~n40252 & n40253;
  assign n40255 = n40251 & ~n40254;
  assign n40256 = ~n40249 & n40255;
  assign n40257 = n40247 & ~n40256;
  assign n40258 = ~n40245 & ~n40257;
  assign n40259 = ~pi39 & ~n40258;
  assign n40260 = pi161 & n32363;
  assign n40261 = ~pi152 & n40260;
  assign n40262 = ~n2809 & ~n40261;
  assign n40263 = pi144 & n32501;
  assign n40264 = ~pi174 & n40263;
  assign n40265 = ~pi299 & ~n40264;
  assign n40266 = pi232 & ~n40265;
  assign n40267 = pi232 & ~n40262;
  assign n40268 = ~n40265 & n40267;
  assign n40269 = ~n40262 & n40266;
  assign n40270 = ~pi72 & ~n64689;
  assign n40271 = pi39 & ~n40270;
  assign n40272 = n62951 & ~n40271;
  assign n40273 = ~n40259 & n40272;
  assign n40274 = ~pi39 & ~n40244;
  assign n40275 = ~n40271 & ~n40274;
  assign n40276 = ~n62951 & n40275;
  assign n40277 = pi75 & ~n40276;
  assign n40278 = ~n40273 & n40277;
  assign n40279 = pi41 & ~n39128;
  assign n40280 = n2929 & ~n39113;
  assign n40281 = ~n40279 & n40280;
  assign n40282 = pi41 & ~n39151;
  assign n40283 = ~n2929 & ~n40282;
  assign n40284 = ~n2929 & ~n39141;
  assign n40285 = ~n40282 & n40284;
  assign n40286 = ~n39141 & n40283;
  assign n40287 = pi228 & ~n64690;
  assign n40288 = ~n40281 & n40287;
  assign n40289 = pi41 & ~n39226;
  assign n40290 = ~n39209 & ~n40289;
  assign n40291 = ~pi228 & ~n40290;
  assign n40292 = ~pi39 & ~n40291;
  assign n40293 = ~n40288 & n40292;
  assign n40294 = n39239 & n64689;
  assign n40295 = ~n40270 & ~n40294;
  assign n40296 = pi39 & ~n40295;
  assign n40297 = n2766 & ~n40296;
  assign n40298 = ~n40293 & n40297;
  assign n40299 = n39045 & n39094;
  assign n40300 = ~n40250 & ~n40299;
  assign n40301 = ~n39273 & ~n40300;
  assign n40302 = ~n40252 & n40301;
  assign n40303 = n2929 & ~n40252;
  assign n40304 = ~n40251 & ~n40303;
  assign n40305 = pi41 & ~n39014;
  assign n40306 = ~n40304 & ~n40305;
  assign n40307 = ~n40302 & ~n40304;
  assign n40308 = ~n40305 & n40307;
  assign n40309 = ~n40302 & n40306;
  assign n40310 = n40247 & ~n64691;
  assign n40311 = ~n40245 & ~n40310;
  assign n40312 = ~pi39 & ~n40311;
  assign n40313 = ~n40271 & ~n40312;
  assign n40314 = n30855 & ~n40313;
  assign n40315 = pi38 & ~n40275;
  assign n40316 = ~pi87 & ~n40315;
  assign n40317 = ~n40314 & n40316;
  assign n40318 = ~n40298 & n40317;
  assign n40319 = pi41 & ~n39013;
  assign n40320 = pi228 & n40300;
  assign n40321 = ~n40319 & n40320;
  assign n40322 = ~pi228 & n40244;
  assign n40323 = n62373 & ~n40322;
  assign n40324 = ~n40321 & n40323;
  assign n40325 = ~n2766 & n40274;
  assign n40326 = pi87 & ~n40325;
  assign n40327 = ~n40271 & n40326;
  assign n40328 = ~n40324 & n40327;
  assign n40329 = ~pi75 & ~n40328;
  assign n40330 = ~n40318 & n40329;
  assign n40331 = ~n40278 & ~n40330;
  assign n40332 = n2580 & ~n40331;
  assign n40333 = ~n2580 & ~n40275;
  assign n40334 = n62455 & ~n40333;
  assign n40335 = ~n40332 & n40334;
  assign n40336 = n33664 & n40261;
  assign n40337 = ~pi72 & ~n40274;
  assign n40338 = ~n62455 & n40337;
  assign n40339 = ~n40336 & n40338;
  assign po199 = ~n40335 & ~n40339;
  assign n40341 = pi44 & ~pi72;
  assign n40342 = ~n2997 & ~n40341;
  assign n40343 = ~pi39 & ~n40342;
  assign n40344 = ~n2929 & n40341;
  assign n40345 = n2997 & ~n40344;
  assign n40346 = n2845 & ~n39095;
  assign n40347 = n2993 & n39012;
  assign n40348 = n62385 & n40347;
  assign n40349 = pi44 & ~n39027;
  assign n40350 = ~n40348 & ~n40349;
  assign n40351 = n40346 & ~n40350;
  assign n40352 = n40345 & ~n40351;
  assign n40353 = n40343 & ~n40352;
  assign n40354 = ~pi72 & n2816;
  assign n40355 = pi39 & n2816;
  assign n40356 = ~pi72 & n40355;
  assign n40357 = pi39 & n40354;
  assign n40358 = ~n40353 & ~n64692;
  assign n40359 = n62951 & ~n40358;
  assign n40360 = pi39 & ~n40354;
  assign n40361 = ~pi39 & ~n40341;
  assign n40362 = ~n40360 & ~n40361;
  assign n40363 = ~n62951 & n40362;
  assign n40364 = pi75 & ~n40363;
  assign n40365 = ~n40359 & n40364;
  assign n40366 = pi44 & n39137;
  assign n40367 = ~n2929 & ~n39150;
  assign n40368 = ~n40366 & n40367;
  assign n40369 = pi44 & n39109;
  assign n40370 = n2929 & ~n39127;
  assign n40371 = ~n40369 & n40370;
  assign n40372 = ~n40368 & ~n40371;
  assign n40373 = pi228 & ~n40372;
  assign n40374 = pi44 & n39204;
  assign n40375 = n39190 & n40341;
  assign n40376 = ~pi228 & ~n64693;
  assign n40377 = ~n64609 & n40376;
  assign n40378 = ~pi39 & ~n40377;
  assign n40379 = ~n40373 & n40378;
  assign n40380 = pi287 & n39044;
  assign n40381 = ~pi72 & ~n40380;
  assign n40382 = n40355 & n40381;
  assign n40383 = n64692 & ~n40380;
  assign n40384 = n2766 & ~n64694;
  assign n40385 = ~n40379 & n40384;
  assign n40386 = pi44 & ~n39265;
  assign n40387 = ~n40347 & ~n40386;
  assign n40388 = n40346 & ~n40387;
  assign n40389 = n40345 & ~n40388;
  assign n40390 = n40343 & ~n40389;
  assign n40391 = n30855 & ~n64692;
  assign n40392 = ~n40390 & n40391;
  assign n40393 = pi38 & ~n40362;
  assign n40394 = ~pi87 & ~n40393;
  assign n40395 = ~n40392 & n40394;
  assign n40396 = ~n40385 & n40395;
  assign n40397 = pi228 & n2766;
  assign n40398 = n39044 & n40397;
  assign n40399 = n40341 & ~n40398;
  assign n40400 = n39012 & n40397;
  assign n40401 = ~pi39 & ~n40400;
  assign n40402 = ~pi39 & ~n40399;
  assign n40403 = ~n40400 & n40402;
  assign n40404 = ~n40399 & n40401;
  assign n40405 = pi87 & ~n40360;
  assign n40406 = ~n64695 & n40405;
  assign n40407 = ~pi75 & ~n40406;
  assign n40408 = ~n40396 & n40407;
  assign n40409 = ~n40365 & ~n40408;
  assign n40410 = n2580 & ~n40409;
  assign n40411 = ~n2580 & ~n40362;
  assign n40412 = n62455 & ~n40411;
  assign n40413 = ~n40410 & n40412;
  assign n40414 = ~pi72 & n34993;
  assign n40415 = pi39 & ~n40414;
  assign n40416 = ~n62455 & ~n40361;
  assign n40417 = ~n40415 & n40416;
  assign n40418 = ~n40413 & ~n40417;
  assign n40419 = ~pi72 & pi99;
  assign n40420 = ~n2997 & ~n40419;
  assign n40421 = ~n2929 & n40419;
  assign n40422 = n2997 & ~n40421;
  assign n40423 = ~n40253 & n40419;
  assign n40424 = n2826 & n40348;
  assign n40425 = ~n40423 & ~n40424;
  assign n40426 = n40303 & ~n40425;
  assign n40427 = n40422 & ~n40426;
  assign n40428 = ~n40420 & ~n40427;
  assign n40429 = ~pi39 & ~n40428;
  assign n40430 = ~pi72 & pi152;
  assign n40431 = n40260 & n40430;
  assign n40432 = pi299 & n40431;
  assign n40433 = ~pi72 & pi174;
  assign n40434 = ~pi299 & n40433;
  assign n40435 = n40263 & n40434;
  assign n40436 = ~n40432 & ~n40435;
  assign n40437 = pi232 & ~n40436;
  assign n40438 = pi39 & ~n40437;
  assign n40439 = n62951 & ~n40438;
  assign n40440 = ~n40429 & n40439;
  assign n40441 = ~pi39 & ~n40419;
  assign n40442 = ~n40438 & ~n40441;
  assign n40443 = ~n62951 & n40442;
  assign n40444 = pi75 & ~n40443;
  assign n40445 = ~n40440 & n40444;
  assign n40446 = pi41 & pi72;
  assign n40447 = pi99 & ~n40446;
  assign n40448 = ~n39113 & n40447;
  assign n40449 = n39431 & ~n40448;
  assign n40450 = ~n39141 & n40447;
  assign n40451 = n39430 & ~n40450;
  assign n40452 = ~n40449 & ~n40451;
  assign n40453 = pi228 & ~n40452;
  assign n40454 = ~n39209 & n40447;
  assign n40455 = n39434 & ~n40454;
  assign n40456 = ~pi39 & ~n40455;
  assign n40457 = ~n40453 & n40456;
  assign n40458 = n33664 & ~n40436;
  assign n40459 = ~n40380 & n40458;
  assign n40460 = n2766 & ~n40459;
  assign n40461 = ~n40457 & n40460;
  assign n40462 = ~n40301 & n40419;
  assign n40463 = n2825 & n39014;
  assign n40464 = ~n40462 & ~n40463;
  assign n40465 = n40303 & ~n40464;
  assign n40466 = n40422 & ~n40465;
  assign n40467 = ~n40420 & ~n40466;
  assign n40468 = ~pi39 & ~n40467;
  assign n40469 = ~n40438 & ~n40468;
  assign n40470 = n30855 & ~n40469;
  assign n40471 = pi38 & ~n40442;
  assign n40472 = ~pi87 & ~n40471;
  assign n40473 = ~n40470 & n40472;
  assign n40474 = ~n40461 & n40473;
  assign n40475 = pi228 & n40299;
  assign n40476 = n40419 & ~n40475;
  assign n40477 = n62373 & ~n64593;
  assign n40478 = n62373 & ~n40476;
  assign n40479 = ~n64593 & n40478;
  assign n40480 = ~n40476 & n40477;
  assign n40481 = ~n62373 & ~n40442;
  assign n40482 = pi87 & ~n40481;
  assign n40483 = ~n64696 & n40482;
  assign n40484 = ~pi75 & ~n40483;
  assign n40485 = ~n40474 & n40484;
  assign n40486 = ~n40445 & ~n40485;
  assign n40487 = n2580 & ~n40486;
  assign n40488 = ~n2580 & ~n40442;
  assign n40489 = n62455 & ~n40488;
  assign n40490 = ~n40487 & n40489;
  assign n40491 = pi232 & n40431;
  assign n40492 = pi39 & ~n40491;
  assign n40493 = ~n62455 & ~n40441;
  assign n40494 = ~n40492 & n40493;
  assign n40495 = ~n40490 & ~n40494;
  assign n40496 = ~n2997 & ~n39093;
  assign n40497 = ~n2929 & n39093;
  assign n40498 = n2997 & ~n40497;
  assign n40499 = ~n2842 & n2929;
  assign n40500 = ~n39028 & n39093;
  assign n40501 = ~n40248 & ~n40500;
  assign n40502 = n40499 & ~n40501;
  assign n40503 = n40498 & ~n40502;
  assign n40504 = ~n40496 & ~n40503;
  assign n40505 = ~pi39 & ~n40504;
  assign n40506 = ~pi161 & ~pi166;
  assign n40507 = pi152 & n40506;
  assign n40508 = n2814 & n40507;
  assign n40509 = ~pi72 & n40508;
  assign n40510 = pi299 & ~n40509;
  assign n40511 = ~pi144 & pi174;
  assign n40512 = ~pi72 & n40511;
  assign n40513 = n32501 & n40511;
  assign n40514 = ~pi72 & n40513;
  assign n40515 = n32501 & n40512;
  assign n40516 = ~pi299 & ~n64697;
  assign n40517 = pi232 & ~n40516;
  assign n40518 = pi232 & ~n40510;
  assign n40519 = ~n40516 & n40518;
  assign n40520 = ~n40510 & n40517;
  assign n40521 = pi39 & ~n64698;
  assign n40522 = n62951 & ~n40521;
  assign n40523 = ~n40505 & n40522;
  assign n40524 = ~pi39 & ~n39093;
  assign n40525 = ~n40521 & ~n40524;
  assign n40526 = ~n62951 & n40525;
  assign n40527 = pi75 & ~n40526;
  assign n40528 = ~n40523 & n40527;
  assign n40529 = pi101 & n39139;
  assign n40530 = ~n2929 & ~n39151;
  assign n40531 = ~n40529 & n40530;
  assign n40532 = pi101 & n39111;
  assign n40533 = n2929 & ~n39128;
  assign n40534 = ~n40532 & n40533;
  assign n40535 = ~n40531 & ~n40534;
  assign n40536 = pi228 & ~n40535;
  assign n40537 = pi101 & n64607;
  assign n40538 = ~pi228 & ~n39226;
  assign n40539 = ~n40537 & n40538;
  assign n40540 = ~pi39 & ~n40539;
  assign n40541 = ~n40536 & n40540;
  assign n40542 = pi299 & n40508;
  assign n40543 = ~pi299 & n40511;
  assign n40544 = n32501 & n40543;
  assign n40545 = ~n40542 & ~n40544;
  assign n40546 = ~pi72 & n33664;
  assign n40547 = ~n40545 & n40546;
  assign n40548 = n40381 & n40513;
  assign n40549 = ~pi299 & ~n40548;
  assign n40550 = n40381 & n40508;
  assign n40551 = pi299 & ~n40550;
  assign n40552 = n33664 & ~n40551;
  assign n40553 = ~n40549 & n40552;
  assign n40554 = n33664 & ~n40549;
  assign n40555 = ~n40551 & n40554;
  assign n40556 = ~n40380 & n40547;
  assign n40557 = n2766 & ~n64699;
  assign n40558 = ~n40541 & n40557;
  assign n40559 = n39093 & ~n64614;
  assign n40560 = ~n39014 & ~n40559;
  assign n40561 = n40499 & ~n40560;
  assign n40562 = n40498 & ~n40561;
  assign n40563 = ~n40496 & ~n40562;
  assign n40564 = ~pi39 & ~n40563;
  assign n40565 = ~n40521 & ~n40564;
  assign n40566 = n30855 & ~n40565;
  assign n40567 = pi38 & ~n40525;
  assign n40568 = ~pi87 & ~n40567;
  assign n40569 = ~n40566 & n40568;
  assign n40570 = ~n40558 & n40569;
  assign n40571 = ~pi101 & n40400;
  assign n40572 = n39045 & n40397;
  assign n40573 = n39093 & ~n40572;
  assign n40574 = ~pi39 & ~n40573;
  assign n40575 = ~n40571 & n40574;
  assign n40576 = pi87 & ~n40521;
  assign n40577 = ~n40575 & n40576;
  assign n40578 = ~pi75 & ~n40577;
  assign n40579 = ~n40570 & n40578;
  assign n40580 = ~n40528 & ~n40579;
  assign n40581 = n2580 & ~n40580;
  assign n40582 = ~n2580 & ~n40525;
  assign n40583 = n62455 & ~n40582;
  assign n40584 = ~n40581 & n40583;
  assign n40585 = pi232 & n40509;
  assign n40586 = pi39 & ~n40585;
  assign n40587 = ~n62455 & ~n40524;
  assign n40588 = ~n40586 & n40587;
  assign n40589 = ~n40584 & ~n40588;
  assign n40590 = pi252 & n2883;
  assign n40591 = n62361 & n64196;
  assign n40592 = n2728 & n39177;
  assign n40593 = n33872 & n40591;
  assign n40594 = ~n40590 & n64700;
  assign n40595 = ~pi137 & n40594;
  assign n40596 = ~pi137 & n2929;
  assign n40597 = ~n62355 & ~n39175;
  assign n40598 = ~pi94 & ~n39986;
  assign n40599 = n64196 & ~n40598;
  assign n40600 = ~n40597 & n40599;
  assign n40601 = ~n2883 & ~n40600;
  assign n40602 = ~pi252 & n40600;
  assign n40603 = n2720 & n2751;
  assign n40604 = n62354 & n40603;
  assign n40605 = n62375 & n40604;
  assign n40606 = n2751 & n62775;
  assign n40607 = n62354 & n62379;
  assign n40608 = n39985 & n64701;
  assign n40609 = pi252 & n40608;
  assign n40610 = n2883 & ~n40609;
  assign n40611 = ~n40602 & n40610;
  assign n40612 = ~n40601 & ~n40611;
  assign n40613 = pi122 & ~n40612;
  assign n40614 = n2852 & n40601;
  assign n40615 = ~n2584 & ~n64700;
  assign n40616 = ~n40611 & ~n40615;
  assign n40617 = ~n40614 & n40616;
  assign n40618 = ~pi122 & ~n40617;
  assign n40619 = ~n40613 & ~n40618;
  assign n40620 = ~pi1093 & ~n40619;
  assign n40621 = ~pi122 & ~n40594;
  assign n40622 = ~n40613 & ~n40621;
  assign n40623 = pi1093 & ~n40622;
  assign n40624 = ~n40620 & ~n40623;
  assign n40625 = n2929 & ~n40624;
  assign n40626 = ~n40596 & ~n40625;
  assign n40627 = ~n40595 & ~n40626;
  assign n40628 = ~pi122 & n64700;
  assign n40629 = pi1093 & ~n40600;
  assign n40630 = ~n3028 & ~n40629;
  assign n40631 = ~n40628 & ~n40630;
  assign n40632 = ~n40620 & ~n40631;
  assign n40633 = ~n2929 & ~n40632;
  assign n40634 = ~pi137 & ~n2929;
  assign n40635 = ~n40633 & ~n40634;
  assign n40636 = n2921 & n40065;
  assign n40637 = ~pi137 & ~n40636;
  assign n40638 = n64700 & n40637;
  assign n40639 = ~n40635 & ~n40638;
  assign n40640 = ~n40627 & ~n40639;
  assign n40641 = n2843 & ~n40640;
  assign n40642 = ~n39960 & n40608;
  assign n40643 = ~n2843 & ~n40642;
  assign n40644 = ~pi137 & ~n2843;
  assign n40645 = ~n40643 & ~n40644;
  assign n40646 = ~n40641 & n40645;
  assign n40647 = ~pi210 & ~n40646;
  assign n40648 = ~n40625 & ~n40633;
  assign n40649 = n2843 & ~n40648;
  assign n40650 = ~n40643 & ~n40649;
  assign n40651 = pi210 & ~n40650;
  assign n40652 = ~n40647 & ~n40651;
  assign n40653 = n2810 & n32363;
  assign n40654 = ~n40652 & ~n40653;
  assign n40655 = ~pi210 & n40640;
  assign n40656 = pi210 & n40648;
  assign n40657 = n40653 & ~n40656;
  assign n40658 = pi210 & ~n40648;
  assign n40659 = ~pi210 & ~n40640;
  assign n40660 = ~n40658 & ~n40659;
  assign n40661 = n40653 & ~n40660;
  assign n40662 = ~n40655 & n40657;
  assign n40663 = pi299 & ~n64702;
  assign n40664 = ~n40654 & n40663;
  assign n40665 = ~pi198 & ~n40646;
  assign n40666 = pi198 & ~n40650;
  assign n40667 = ~n40665 & ~n40666;
  assign n40668 = n2808 & n2814;
  assign n40669 = ~n40667 & ~n40668;
  assign n40670 = ~pi198 & n40640;
  assign n40671 = pi198 & n40648;
  assign n40672 = n40668 & ~n40671;
  assign n40673 = pi198 & ~n40648;
  assign n40674 = ~pi198 & ~n40640;
  assign n40675 = ~n40673 & ~n40674;
  assign n40676 = n40668 & ~n40675;
  assign n40677 = ~n40670 & n40672;
  assign n40678 = ~pi299 & ~n64703;
  assign n40679 = ~n40669 & n40678;
  assign n40680 = ~n40664 & ~n40679;
  assign n40681 = pi232 & ~n40680;
  assign n40682 = ~pi299 & ~n40667;
  assign n40683 = pi299 & ~n40652;
  assign n40684 = ~pi232 & ~n40683;
  assign n40685 = ~pi232 & ~n40682;
  assign n40686 = ~n40683 & n40685;
  assign n40687 = ~n40682 & n40684;
  assign n40688 = n3318 & ~n64704;
  assign n40689 = ~n40681 & n40688;
  assign n40690 = n62455 & n64082;
  assign n40691 = n62455 & n64086;
  assign n40692 = ~pi74 & n40691;
  assign n40693 = n6793 & n35113;
  assign n40694 = n34066 & n64498;
  assign n40695 = n62455 & n6794;
  assign n40696 = n2806 & n64706;
  assign n40697 = n64083 & n35113;
  assign n40698 = ~pi92 & n40697;
  assign n40699 = n64081 & n35113;
  assign n40700 = n2764 & n63888;
  assign n40701 = n2883 & ~n64700;
  assign n40702 = ~n40590 & ~n40701;
  assign n40703 = ~n40590 & ~n40601;
  assign n40704 = ~n40701 & n40703;
  assign n40705 = ~n40601 & n40702;
  assign n40706 = n3028 & ~n64707;
  assign n40707 = ~n40613 & ~n40706;
  assign n40708 = n2929 & ~n40707;
  assign n40709 = ~n2929 & n40629;
  assign n40710 = ~pi1093 & ~n40612;
  assign n40711 = ~n40709 & ~n40710;
  assign n40712 = ~n40708 & n40711;
  assign n40713 = n2843 & n40712;
  assign n40714 = ~n2843 & n40608;
  assign n40715 = ~n64669 & n40714;
  assign n40716 = ~n40713 & ~n40715;
  assign n40717 = pi210 & ~n40716;
  assign n40718 = pi137 & n40710;
  assign n40719 = ~pi137 & ~n64707;
  assign n40720 = ~pi1093 & n40719;
  assign n40721 = ~n40629 & ~n40720;
  assign n40722 = ~n40629 & ~n40718;
  assign n40723 = ~n40720 & n40722;
  assign n40724 = ~n40718 & n40721;
  assign n40725 = n2843 & n64708;
  assign n40726 = ~n40714 & ~n40725;
  assign n40727 = n38260 & n40644;
  assign n40728 = ~n2929 & ~n40727;
  assign n40729 = ~n40726 & n40728;
  assign n40730 = pi137 & ~n40707;
  assign n40731 = ~n40718 & ~n40719;
  assign n40732 = ~n40730 & n40731;
  assign n40733 = n2843 & ~n40732;
  assign n40734 = pi137 & ~n3028;
  assign n40735 = n2883 & ~n40734;
  assign n40736 = n40608 & ~n40735;
  assign n40737 = ~n2843 & ~n40736;
  assign n40738 = n2929 & ~n40737;
  assign n40739 = ~n40733 & n40738;
  assign n40740 = ~n40729 & ~n40739;
  assign n40741 = ~pi210 & ~n40740;
  assign n40742 = ~n40717 & ~n40741;
  assign n40743 = ~n40653 & ~n40742;
  assign n40744 = ~n2929 & n64708;
  assign n40745 = n2929 & n40732;
  assign n40746 = ~n40744 & ~n40745;
  assign n40747 = ~pi210 & n40746;
  assign n40748 = pi210 & ~n40712;
  assign n40749 = n40653 & ~n40748;
  assign n40750 = ~pi210 & ~n40746;
  assign n40751 = pi210 & n40712;
  assign n40752 = ~n40750 & ~n40751;
  assign n40753 = n40653 & ~n40752;
  assign n40754 = ~n40747 & n40749;
  assign n40755 = pi299 & ~n64709;
  assign n40756 = ~n40743 & n40755;
  assign n40757 = pi198 & ~n40716;
  assign n40758 = ~pi198 & ~n40740;
  assign n40759 = ~n40757 & ~n40758;
  assign n40760 = ~n40668 & ~n40759;
  assign n40761 = ~pi198 & n40746;
  assign n40762 = pi198 & ~n40712;
  assign n40763 = n40668 & ~n40762;
  assign n40764 = ~pi198 & ~n40746;
  assign n40765 = pi198 & n40712;
  assign n40766 = ~n40764 & ~n40765;
  assign n40767 = n40668 & ~n40766;
  assign n40768 = ~n40761 & n40763;
  assign n40769 = ~pi299 & ~n64710;
  assign n40770 = ~n40760 & n40769;
  assign n40771 = ~n40756 & ~n40770;
  assign n40772 = pi232 & ~n40771;
  assign n40773 = pi299 & ~n40742;
  assign n40774 = ~pi299 & ~n40759;
  assign n40775 = ~pi232 & ~n40774;
  assign n40776 = ~pi232 & ~n40773;
  assign n40777 = ~n40774 & n40776;
  assign n40778 = ~n40773 & n40775;
  assign n40779 = ~n40772 & ~n64711;
  assign n40780 = ~n3318 & ~n40779;
  assign n40781 = n64705 & ~n40780;
  assign n40782 = ~n40681 & ~n64704;
  assign n40783 = n3318 & ~n40782;
  assign n40784 = ~n3318 & ~n64711;
  assign n40785 = ~n40772 & n40784;
  assign n40786 = ~n40783 & ~n40785;
  assign n40787 = n64705 & ~n40786;
  assign n40788 = ~n40689 & n40781;
  assign n40789 = ~pi99 & ~n40284;
  assign n40790 = ~n40280 & n40789;
  assign n40791 = pi113 & ~n39092;
  assign n40792 = ~n40790 & n40791;
  assign n40793 = ~pi113 & n39432;
  assign n40794 = pi228 & ~n40793;
  assign n40795 = ~n40792 & n40794;
  assign n40796 = pi113 & n39211;
  assign n40797 = ~pi228 & ~n39228;
  assign n40798 = ~n40796 & n40797;
  assign n40799 = ~pi39 & ~n40798;
  assign n40800 = ~n40795 & n40799;
  assign n40801 = n2766 & ~n40800;
  assign n40802 = ~pi72 & pi113;
  assign n40803 = ~pi39 & n40802;
  assign n40804 = pi38 & ~n40803;
  assign n40805 = ~n62388 & ~n64615;
  assign n40806 = n39666 & ~n40805;
  assign n40807 = n40802 & ~n40806;
  assign n40808 = ~n62388 & n39666;
  assign n40809 = ~pi113 & n40808;
  assign n40810 = n40463 & n40809;
  assign n40811 = ~n40807 & ~n40810;
  assign n40812 = ~pi39 & ~n40811;
  assign n40813 = n30855 & ~n40812;
  assign n40814 = ~n40804 & ~n40813;
  assign n40815 = ~n40801 & n40814;
  assign n40816 = ~pi87 & ~n40815;
  assign n40817 = ~n64590 & n40802;
  assign n40818 = ~n39064 & ~n40817;
  assign n40819 = n62373 & ~n40818;
  assign n40820 = ~n2766 & n40803;
  assign n40821 = pi87 & ~n40820;
  assign n40822 = ~n40819 & n40821;
  assign n40823 = ~n40816 & ~n40822;
  assign n40824 = ~pi75 & ~n40823;
  assign n40825 = n62385 & n40810;
  assign n40826 = ~n62388 & ~n39029;
  assign n40827 = n39666 & ~n40826;
  assign n40828 = n40802 & ~n40827;
  assign n40829 = ~n40825 & ~n40828;
  assign n40830 = n2806 & ~n40829;
  assign n40831 = ~n62951 & n40803;
  assign n40832 = pi75 & ~n40831;
  assign n40833 = ~n40830 & n40832;
  assign n40834 = ~n40824 & ~n40833;
  assign n40835 = n40103 & ~n40834;
  assign n40836 = ~n40103 & ~n40803;
  assign po271 = ~n40835 & ~n40836;
  assign n40838 = ~pi72 & pi114;
  assign n40839 = pi114 & n39512;
  assign n40840 = ~n39031 & n40838;
  assign n40841 = ~n39021 & n39667;
  assign n40842 = n39667 & ~n64713;
  assign n40843 = ~n39021 & n40842;
  assign n40844 = ~n64713 & n40841;
  assign n40845 = ~n39667 & ~n40838;
  assign n40846 = n2806 & ~n40845;
  assign n40847 = n39031 & n39666;
  assign n40848 = ~pi115 & n40847;
  assign n40849 = n40838 & ~n40848;
  assign n40850 = n39021 & n39667;
  assign n40851 = ~n40849 & ~n40850;
  assign n40852 = n2806 & ~n40851;
  assign n40853 = ~n64714 & n40846;
  assign n40854 = ~pi39 & n40838;
  assign n40855 = ~n62951 & n40854;
  assign n40856 = pi75 & ~n40855;
  assign n40857 = ~n64715 & n40856;
  assign n40858 = pi114 & n39456;
  assign n40859 = ~pi114 & n64633;
  assign n40860 = ~pi115 & ~n40859;
  assign n40861 = pi114 & ~n39456;
  assign n40862 = ~pi114 & ~n64633;
  assign n40863 = ~n40861 & ~n40862;
  assign n40864 = ~pi115 & ~n40863;
  assign n40865 = ~n40858 & n40860;
  assign n40866 = pi115 & ~n40838;
  assign n40867 = ~pi39 & ~n40866;
  assign n40868 = ~n64716 & n40867;
  assign n40869 = n2766 & ~n40868;
  assign n40870 = pi114 & ~n64617;
  assign n40871 = ~n39020 & n39667;
  assign n40872 = n39667 & ~n40870;
  assign n40873 = ~n39020 & n40872;
  assign n40874 = ~n40870 & n40871;
  assign n40875 = ~pi39 & ~n40845;
  assign n40876 = ~n64717 & n40875;
  assign n40877 = n30855 & ~n40876;
  assign n40878 = pi38 & ~n40854;
  assign n40879 = ~pi87 & ~n40878;
  assign n40880 = ~n40877 & n40879;
  assign n40881 = ~n40869 & n40880;
  assign n40882 = ~n39492 & n40838;
  assign n40883 = ~n39069 & ~n40882;
  assign n40884 = ~n2766 & ~n40854;
  assign n40885 = n39758 & ~n40884;
  assign n40886 = ~n39055 & n40838;
  assign n40887 = n2766 & ~n40886;
  assign n40888 = ~n39069 & n40887;
  assign n40889 = n40885 & ~n40888;
  assign n40890 = ~n40883 & n40885;
  assign n40891 = ~pi75 & ~n64718;
  assign n40892 = ~n40881 & n40891;
  assign n40893 = ~n40857 & ~n40892;
  assign n40894 = n40103 & ~n40893;
  assign n40895 = ~n40103 & ~n40854;
  assign po272 = ~n40894 & ~n40895;
  assign n40897 = ~pi72 & pi115;
  assign n40898 = ~n40847 & n40897;
  assign n40899 = ~pi52 & n2835;
  assign n40900 = ~pi114 & n2838;
  assign n40901 = ~pi115 & ~n64719;
  assign n40902 = n64588 & n40901;
  assign n40903 = n62385 & n39666;
  assign n40904 = n40902 & n40903;
  assign n40905 = ~n40898 & ~n40904;
  assign n40906 = n62385 & n40902;
  assign n40907 = pi115 & n39512;
  assign n40908 = n39666 & ~n40907;
  assign n40909 = ~n40906 & n40908;
  assign n40910 = ~n39666 & ~n40897;
  assign n40911 = n2806 & ~n40910;
  assign n40912 = ~n40909 & n40911;
  assign n40913 = n2806 & ~n40905;
  assign n40914 = ~pi39 & n40897;
  assign n40915 = ~n62951 & n40914;
  assign n40916 = pi75 & ~n40915;
  assign n40917 = ~n64720 & n40916;
  assign n40918 = pi115 & ~n39456;
  assign n40919 = ~pi115 & ~n64633;
  assign n40920 = ~pi39 & ~n40919;
  assign n40921 = ~n40918 & n40920;
  assign n40922 = n2766 & ~n40921;
  assign n40923 = pi115 & ~n64617;
  assign n40924 = n39666 & ~n40902;
  assign n40925 = n39666 & ~n40923;
  assign n40926 = ~n40902 & n40925;
  assign n40927 = ~n40923 & n40924;
  assign n40928 = ~pi39 & ~n40910;
  assign n40929 = ~n64721 & n40928;
  assign n40930 = n30855 & ~n40929;
  assign n40931 = pi38 & ~n40914;
  assign n40932 = ~pi87 & ~n40931;
  assign n40933 = ~n40930 & n40932;
  assign n40934 = ~n40922 & n40933;
  assign n40935 = ~n64591 & n40897;
  assign n40936 = n2766 & ~n40935;
  assign n40937 = ~n39068 & n40936;
  assign n40938 = ~n2766 & ~n40914;
  assign n40939 = n39758 & ~n40938;
  assign n40940 = ~n40937 & n40939;
  assign n40941 = ~pi75 & ~n40940;
  assign n40942 = ~n40934 & n40941;
  assign n40943 = ~n40917 & ~n40942;
  assign n40944 = n40103 & ~n40943;
  assign n40945 = ~n40103 & ~n40914;
  assign po273 = ~n40944 & ~n40945;
  assign n40947 = n2929 & ~n39117;
  assign n40948 = ~n2929 & ~n39145;
  assign n40949 = pi116 & ~n40948;
  assign n40950 = ~n40947 & n40949;
  assign n40951 = pi116 & n39145;
  assign n40952 = ~n2929 & ~n40951;
  assign n40953 = pi116 & ~n40947;
  assign n40954 = ~n64602 & ~n40953;
  assign n40955 = ~n40952 & ~n40954;
  assign n40956 = n39438 & ~n40955;
  assign n40957 = n64632 & ~n40950;
  assign n40958 = pi116 & n39213;
  assign n40959 = n39442 & ~n40958;
  assign n40960 = ~pi39 & ~n40959;
  assign n40961 = ~n64722 & n40960;
  assign n40962 = n2766 & ~n40961;
  assign n40963 = ~pi72 & pi116;
  assign n40964 = ~n39666 & n40963;
  assign n40965 = ~n39270 & n40963;
  assign n40966 = ~n64588 & ~n40965;
  assign n40967 = n40808 & ~n40966;
  assign n40968 = ~n40964 & ~n40967;
  assign n40969 = ~pi39 & ~n40968;
  assign n40970 = n30855 & ~n40969;
  assign n40971 = ~pi39 & n40963;
  assign n40972 = pi38 & ~n40971;
  assign n40973 = ~pi87 & ~n40972;
  assign n40974 = ~n40970 & n40973;
  assign n40975 = ~n40962 & n40974;
  assign n40976 = ~pi38 & ~pi113;
  assign n40977 = n64590 & n40976;
  assign n40978 = n40963 & ~n40977;
  assign n40979 = ~n64594 & ~n40978;
  assign n40980 = ~pi113 & n64590;
  assign n40981 = n40963 & ~n40980;
  assign n40982 = ~pi38 & ~n40981;
  assign n40983 = ~pi38 & ~n64594;
  assign n40984 = ~n40981 & n40983;
  assign n40985 = ~n64594 & n40982;
  assign n40986 = ~n40972 & ~n64723;
  assign n40987 = ~n40972 & ~n40979;
  assign n40988 = ~pi100 & ~n64724;
  assign n40989 = pi100 & ~n40971;
  assign n40990 = n39758 & ~n40989;
  assign n40991 = ~n40988 & n40990;
  assign n40992 = ~pi75 & ~n40991;
  assign n40993 = ~n40975 & n40992;
  assign n40994 = ~n39030 & n40963;
  assign n40995 = ~n39515 & ~n40994;
  assign n40996 = n40808 & ~n40995;
  assign n40997 = ~n40964 & ~n40996;
  assign n40998 = n2806 & ~n40997;
  assign n40999 = ~n62951 & n40971;
  assign n41000 = pi75 & ~n40999;
  assign n41001 = ~n40998 & n41000;
  assign n41002 = ~n40993 & ~n41001;
  assign n41003 = n40103 & ~n41002;
  assign n41004 = ~n40103 & ~n40971;
  assign po274 = ~n41003 & ~n41004;
  assign n41006 = ~pi332 & ~pi1144;
  assign n41007 = pi215 & ~n41006;
  assign n41008 = pi265 & ~pi332;
  assign n41009 = pi216 & ~n41008;
  assign n41010 = pi105 & pi228;
  assign n41011 = pi234 & n30613;
  assign n41012 = ~pi332 & ~n41011;
  assign n41013 = n41010 & n41012;
  assign n41014 = pi153 & ~pi332;
  assign n41015 = ~n41010 & n41014;
  assign n41016 = ~pi216 & ~n41015;
  assign n41017 = ~n41013 & n41016;
  assign n41018 = ~n41009 & ~n41017;
  assign n41019 = ~pi221 & ~n41018;
  assign n41020 = ~pi216 & pi833;
  assign n41021 = pi929 & n41020;
  assign n41022 = pi1144 & ~n41020;
  assign n41023 = ~pi332 & ~n41022;
  assign n41024 = ~pi332 & ~n41021;
  assign n41025 = ~n41022 & n41024;
  assign n41026 = ~n41021 & n41023;
  assign n41027 = pi221 & ~n64725;
  assign n41028 = ~n41019 & ~n41027;
  assign n41029 = ~pi215 & ~n41028;
  assign n41030 = ~n41007 & ~n41029;
  assign n41031 = ~n62380 & ~n30613;
  assign n41032 = pi234 & ~n41031;
  assign n41033 = ~pi234 & n62380;
  assign n41034 = ~n41032 & ~n41033;
  assign n41035 = pi137 & ~n41034;
  assign n41036 = n41012 & ~n41035;
  assign n41037 = ~pi215 & ~pi221;
  assign n41038 = n41016 & n41037;
  assign n41039 = ~n41036 & n41038;
  assign n41040 = n64085 & n41039;
  assign n41041 = ~pi59 & n41040;
  assign n41042 = n41030 & ~n41041;
  assign n41043 = pi57 & ~n41042;
  assign n41044 = ~pi105 & ~pi153;
  assign n41045 = pi228 & ~pi332;
  assign n41046 = ~n41044 & n41045;
  assign n41047 = ~n30613 & ~n33962;
  assign n41048 = n2772 & n64295;
  assign n41049 = pi225 & n2771;
  assign n41050 = pi225 & n33949;
  assign n41051 = n2771 & n41050;
  assign n41052 = n33949 & n41049;
  assign n41053 = n41048 & n64726;
  assign n41054 = pi32 & ~n41053;
  assign n41055 = n2733 & ~n38178;
  assign n41056 = pi35 & n62363;
  assign n41057 = ~pi225 & n41056;
  assign n41058 = ~n33939 & ~n41057;
  assign n41059 = ~pi35 & ~n35354;
  assign n41060 = n34979 & ~n40178;
  assign n41061 = n30645 & ~n33919;
  assign n41062 = n30641 & ~n41061;
  assign n41063 = n30639 & ~n41062;
  assign n41064 = ~n30637 & ~n41063;
  assign n41065 = ~pi86 & ~n41064;
  assign n41066 = n30715 & ~n41065;
  assign n41067 = n33873 & ~n41066;
  assign n41068 = ~n30937 & ~n41067;
  assign n41069 = ~pi108 & ~n41068;
  assign n41070 = n33870 & ~n41069;
  assign n41071 = n30750 & ~n41070;
  assign n41072 = ~n30748 & ~n41071;
  assign n41073 = n2866 & ~n41072;
  assign n41074 = n64688 & ~n41073;
  assign n41075 = n40180 & ~n41074;
  assign n41076 = n41060 & ~n41075;
  assign n41077 = n41059 & ~n41076;
  assign n41078 = n41058 & ~n41077;
  assign n41079 = ~pi51 & ~n41078;
  assign n41080 = n41055 & ~n41079;
  assign n41081 = ~pi72 & ~n41080;
  assign n41082 = n33860 & ~n41081;
  assign n41083 = n33859 & ~n41082;
  assign n41084 = ~n41054 & ~n41083;
  assign n41085 = ~pi95 & ~n41084;
  assign n41086 = n41047 & ~n41085;
  assign n41087 = pi137 & ~n41086;
  assign n41088 = ~pi70 & ~n41057;
  assign n41089 = ~pi51 & n41088;
  assign n41090 = ~n33939 & n41089;
  assign n41091 = ~n30639 & n32085;
  assign n41092 = n2694 & n62361;
  assign n41093 = n41091 & n41092;
  assign n41094 = ~pi35 & ~n41093;
  assign n41095 = n41090 & ~n41094;
  assign n41096 = n2730 & n41095;
  assign n41097 = ~pi32 & ~n41096;
  assign n41098 = ~pi95 & ~n41054;
  assign n41099 = ~n41097 & n41098;
  assign n41100 = ~pi137 & ~n41099;
  assign n41101 = n30860 & n41100;
  assign n41102 = ~pi97 & ~n41091;
  assign n41103 = n2715 & n30940;
  assign n41104 = ~n41102 & n41103;
  assign n41105 = n30939 & n41103;
  assign n41106 = ~n41102 & n41105;
  assign n41107 = n30939 & n41104;
  assign n41108 = ~pi35 & ~n64727;
  assign n41109 = n62395 & n41108;
  assign n41110 = ~n62395 & n41094;
  assign n41111 = n2730 & n41090;
  assign n41112 = n62376 & n41058;
  assign n41113 = ~n41110 & n64728;
  assign n41114 = ~n62395 & ~n41094;
  assign n41115 = n62395 & ~n41108;
  assign n41116 = ~n41114 & ~n41115;
  assign n41117 = n64728 & ~n41116;
  assign n41118 = ~n41109 & n41113;
  assign n41119 = ~pi32 & ~n64729;
  assign n41120 = n41098 & ~n41119;
  assign n41121 = ~pi137 & ~n41120;
  assign n41122 = ~n30860 & n41121;
  assign n41123 = ~n41101 & ~n41122;
  assign n41124 = ~n41087 & n41123;
  assign n41125 = ~pi234 & ~n41124;
  assign n41126 = n2772 & n33949;
  assign n41127 = ~pi51 & n2726;
  assign n41128 = ~pi40 & n2772;
  assign n41129 = n62364 & n64730;
  assign n41130 = n62363 & n41126;
  assign n41131 = n33867 & n64731;
  assign n41132 = n41083 & ~n41131;
  assign n41133 = ~n41054 & ~n41132;
  assign n41134 = ~pi95 & ~n41133;
  assign n41135 = pi479 & n33962;
  assign n41136 = ~n41134 & ~n41135;
  assign n41137 = pi137 & ~n41136;
  assign n41138 = pi95 & pi479;
  assign n41139 = ~pi96 & ~n41095;
  assign n41140 = n38977 & ~n41139;
  assign n41141 = ~pi32 & ~n41140;
  assign n41142 = ~n41054 & ~n41141;
  assign n41143 = ~pi95 & ~n41142;
  assign n41144 = ~n41138 & ~n41143;
  assign n41145 = ~pi137 & ~n41144;
  assign n41146 = ~n41137 & ~n41145;
  assign n41147 = n30860 & n41146;
  assign n41148 = n41090 & ~n41108;
  assign n41149 = ~pi96 & ~n41148;
  assign n41150 = n38977 & ~n41149;
  assign n41151 = ~pi32 & ~n41150;
  assign n41152 = ~n41054 & ~n41151;
  assign n41153 = ~pi95 & ~n41152;
  assign n41154 = ~n41138 & ~n41153;
  assign n41155 = n62395 & n41154;
  assign n41156 = ~n62395 & n41144;
  assign n41157 = ~pi137 & ~n41156;
  assign n41158 = ~n41155 & n41157;
  assign n41159 = ~n2929 & n41146;
  assign n41160 = n2930 & ~n41138;
  assign n41161 = ~n41153 & n41160;
  assign n41162 = ~n2930 & n41144;
  assign n41163 = ~pi137 & ~n41162;
  assign n41164 = ~pi137 & ~n41161;
  assign n41165 = ~n41162 & n41164;
  assign n41166 = ~n41161 & n41163;
  assign n41167 = n2929 & ~n64732;
  assign n41168 = ~n41137 & n41167;
  assign n41169 = ~n41159 & ~n41168;
  assign n41170 = ~n41137 & ~n41158;
  assign n41171 = ~n30860 & ~n64733;
  assign n41172 = pi234 & ~n41171;
  assign n41173 = ~n41147 & n41172;
  assign n41174 = ~n41125 & ~n41173;
  assign n41175 = ~pi210 & ~n41174;
  assign n41176 = pi225 & n33956;
  assign n41177 = pi32 & ~n41176;
  assign n41178 = ~pi95 & ~n41177;
  assign n41179 = ~n41141 & n41178;
  assign n41180 = ~n30613 & ~n41179;
  assign n41181 = ~pi137 & n41180;
  assign n41182 = ~n41132 & ~n41177;
  assign n41183 = ~pi95 & ~n41182;
  assign n41184 = ~n41135 & ~n41183;
  assign n41185 = pi137 & ~n41184;
  assign n41186 = ~n41181 & ~n41185;
  assign n41187 = pi234 & n41186;
  assign n41188 = ~n41097 & n41178;
  assign n41189 = ~pi137 & ~n41188;
  assign n41190 = ~n41083 & ~n41177;
  assign n41191 = ~pi95 & ~n41190;
  assign n41192 = n41047 & ~n41191;
  assign n41193 = pi137 & ~n41192;
  assign n41194 = ~n41189 & ~n41193;
  assign n41195 = ~pi234 & n41194;
  assign n41196 = pi210 & ~n41195;
  assign n41197 = ~n41187 & n41196;
  assign n41198 = pi105 & ~n41197;
  assign n41199 = ~pi210 & ~n41146;
  assign n41200 = pi210 & ~n41186;
  assign n41201 = pi234 & ~n41200;
  assign n41202 = ~n41199 & n41201;
  assign n41203 = ~n41087 & ~n41100;
  assign n41204 = ~pi210 & ~n41203;
  assign n41205 = pi210 & ~n41194;
  assign n41206 = ~pi234 & ~n41205;
  assign n41207 = ~n41204 & n41206;
  assign n41208 = n30860 & ~n41207;
  assign n41209 = ~n41202 & n41208;
  assign n41210 = ~pi210 & n64733;
  assign n41211 = ~n41200 & ~n41210;
  assign n41212 = n41201 & ~n41210;
  assign n41213 = pi234 & n41211;
  assign n41214 = ~n41087 & ~n41121;
  assign n41215 = ~pi210 & ~n41214;
  assign n41216 = ~n41205 & ~n41215;
  assign n41217 = n41206 & ~n41215;
  assign n41218 = ~pi234 & n41216;
  assign n41219 = ~n30860 & ~n64735;
  assign n41220 = ~n64734 & n41219;
  assign n41221 = pi105 & ~n41220;
  assign n41222 = ~n41209 & n41221;
  assign n41223 = ~n41175 & n41198;
  assign n41224 = n41046 & ~n64736;
  assign n41225 = ~pi109 & ~n41070;
  assign n41226 = ~n30748 & ~n41225;
  assign n41227 = n2866 & ~n41226;
  assign n41228 = n64688 & ~n41227;
  assign n41229 = n40180 & ~n41228;
  assign n41230 = n41060 & ~n41229;
  assign n41231 = n41059 & ~n41230;
  assign n41232 = n41058 & ~n41231;
  assign n41233 = ~pi51 & ~n41232;
  assign n41234 = n41055 & ~n41233;
  assign n41235 = ~pi72 & ~n41234;
  assign n41236 = n33860 & ~n41235;
  assign n41237 = n33859 & ~n41236;
  assign n41238 = ~n41131 & n41237;
  assign n41239 = ~n41054 & ~n41238;
  assign n41240 = ~pi95 & pi137;
  assign n41241 = ~n41239 & n41240;
  assign n41242 = n2929 & ~n30860;
  assign n41243 = n2930 & n41242;
  assign n41244 = n62395 & ~n30860;
  assign n41245 = n41154 & n64737;
  assign n41246 = n41144 & ~n64737;
  assign n41247 = ~pi137 & ~n41246;
  assign n41248 = ~n41245 & n41247;
  assign n41249 = ~n33962 & ~n41248;
  assign n41250 = ~pi95 & ~n41239;
  assign n41251 = ~n33962 & ~n41250;
  assign n41252 = pi137 & ~n41251;
  assign n41253 = ~n41162 & n41242;
  assign n41254 = ~n33962 & n41144;
  assign n41255 = ~n41253 & n41254;
  assign n41256 = ~n33962 & n41242;
  assign n41257 = n41161 & n41256;
  assign n41258 = ~pi137 & ~n41257;
  assign n41259 = ~n41255 & n41258;
  assign n41260 = ~n41252 & ~n41259;
  assign n41261 = ~n41241 & n41249;
  assign n41262 = ~pi210 & ~n64738;
  assign n41263 = pi234 & ~n41262;
  assign n41264 = pi210 & ~n41189;
  assign n41265 = n41176 & n41264;
  assign n41266 = n41054 & ~n41265;
  assign n41267 = ~n41237 & ~n41266;
  assign n41268 = ~pi95 & ~n41267;
  assign n41269 = n41047 & ~n41268;
  assign n41270 = pi137 & ~n41269;
  assign n41271 = ~pi210 & ~pi234;
  assign n41272 = ~n41101 & n41271;
  assign n41273 = ~n41122 & n41272;
  assign n41274 = ~n41264 & ~n41273;
  assign n41275 = ~n41054 & ~n41237;
  assign n41276 = ~pi95 & ~n41275;
  assign n41277 = n41047 & ~n41276;
  assign n41278 = pi137 & ~n41277;
  assign n41279 = n41273 & ~n41278;
  assign n41280 = ~n41177 & ~n41237;
  assign n41281 = ~pi95 & ~n41280;
  assign n41282 = n41047 & ~n41281;
  assign n41283 = pi137 & ~n41282;
  assign n41284 = n41264 & ~n41283;
  assign n41285 = ~n41279 & ~n41284;
  assign n41286 = ~n41270 & ~n41274;
  assign n41287 = ~n41263 & n64739;
  assign n41288 = ~n41177 & ~n41238;
  assign n41289 = ~pi95 & ~n41288;
  assign n41290 = pi137 & ~n33962;
  assign n41291 = ~n41289 & n41290;
  assign n41292 = ~pi137 & ~n33962;
  assign n41293 = ~n41180 & n41292;
  assign n41294 = pi210 & pi234;
  assign n41295 = ~n41293 & n41294;
  assign n41296 = ~n41291 & n41295;
  assign n41297 = ~n41287 & ~n41296;
  assign n41298 = n41014 & ~n41297;
  assign n41299 = pi225 & pi841;
  assign n41300 = n33956 & ~n41299;
  assign n41301 = pi32 & ~n41300;
  assign n41302 = ~pi95 & ~n41301;
  assign n41303 = n2730 & ~n41088;
  assign n41304 = n2726 & n64090;
  assign n41305 = ~n41088 & n41304;
  assign n41306 = n30621 & n41303;
  assign n41307 = ~pi32 & ~n64740;
  assign n41308 = n41302 & ~n41307;
  assign n41309 = pi137 & ~n41308;
  assign n41310 = ~pi35 & ~n40176;
  assign n41311 = ~pi53 & n41062;
  assign n41312 = ~pi86 & ~n41311;
  assign n41313 = n30715 & ~n41312;
  assign n41314 = n33873 & ~n41313;
  assign n41315 = ~n30937 & ~n41314;
  assign n41316 = ~pi108 & ~n41315;
  assign n41317 = n33870 & ~n41316;
  assign n41318 = ~pi109 & ~n41317;
  assign n41319 = ~n30748 & ~n41318;
  assign n41320 = n2866 & ~n41319;
  assign n41321 = n64688 & ~n41320;
  assign n41322 = n40180 & ~n41321;
  assign n41323 = n40179 & ~n41322;
  assign n41324 = ~pi93 & ~n41323;
  assign n41325 = n41310 & ~n41324;
  assign n41326 = n41089 & ~n41325;
  assign n41327 = n2733 & ~n30620;
  assign n41328 = ~n41326 & n41327;
  assign n41329 = ~pi72 & ~n41328;
  assign n41330 = n33860 & ~n41329;
  assign n41331 = n33859 & ~n41330;
  assign n41332 = ~n62395 & n41331;
  assign n41333 = n62395 & n33859;
  assign n41334 = ~pi97 & ~n41314;
  assign n41335 = ~pi108 & ~n41334;
  assign n41336 = n33870 & ~n41335;
  assign n41337 = ~pi109 & ~n41336;
  assign n41338 = ~n30748 & ~n41337;
  assign n41339 = n2866 & ~n41338;
  assign n41340 = n64688 & ~n41339;
  assign n41341 = n40180 & ~n41340;
  assign n41342 = n40179 & ~n41341;
  assign n41343 = ~pi93 & ~n41342;
  assign n41344 = n41310 & ~n41343;
  assign n41345 = n41089 & ~n41344;
  assign n41346 = n41327 & ~n41345;
  assign n41347 = ~pi72 & ~n41346;
  assign n41348 = n33860 & ~n41347;
  assign n41349 = n41333 & ~n41348;
  assign n41350 = ~n41301 & ~n41349;
  assign n41351 = ~n41332 & n41350;
  assign n41352 = ~pi95 & ~n41351;
  assign n41353 = n41047 & ~n41352;
  assign n41354 = ~pi137 & ~n41353;
  assign n41355 = ~n41309 & ~n41354;
  assign n41356 = ~pi210 & ~n41355;
  assign n41357 = pi146 & n41356;
  assign n41358 = pi234 & ~pi332;
  assign n41359 = ~pi225 & n33956;
  assign n41360 = pi32 & ~n41359;
  assign n41361 = ~n41331 & ~n41360;
  assign n41362 = ~pi95 & ~n41361;
  assign n41363 = ~pi137 & n41047;
  assign n41364 = ~n41362 & n41363;
  assign n41365 = ~pi95 & ~n41360;
  assign n41366 = pi137 & n41365;
  assign n41367 = ~n41307 & n41366;
  assign n41368 = pi210 & ~n41367;
  assign n41369 = ~n41364 & n41368;
  assign n41370 = n41358 & ~n41369;
  assign n41371 = ~pi146 & ~pi210;
  assign n41372 = ~n41301 & ~n41331;
  assign n41373 = ~pi95 & ~n41372;
  assign n41374 = n41047 & ~n41373;
  assign n41375 = ~pi137 & ~n41374;
  assign n41376 = ~n41309 & ~n41375;
  assign n41377 = n41371 & ~n41376;
  assign n41378 = n41370 & ~n41377;
  assign n41379 = ~n41357 & n41378;
  assign n41380 = n33868 & ~n41328;
  assign n41381 = n33860 & ~n41380;
  assign n41382 = n33859 & ~n41381;
  assign n41383 = ~n62395 & n41382;
  assign n41384 = n33868 & ~n41346;
  assign n41385 = n33860 & ~n41384;
  assign n41386 = n41333 & ~n41385;
  assign n41387 = ~n41301 & ~n41386;
  assign n41388 = ~n41383 & n41387;
  assign n41389 = ~pi95 & ~n41388;
  assign n41390 = ~n33962 & ~n41389;
  assign n41391 = ~pi137 & ~n41390;
  assign n41392 = ~pi72 & n2750;
  assign n41393 = n33867 & n41392;
  assign n41394 = n41307 & ~n41393;
  assign n41395 = n41302 & ~n41394;
  assign n41396 = pi137 & ~n30614;
  assign n41397 = ~n41395 & n41396;
  assign n41398 = ~n41391 & ~n41397;
  assign n41399 = ~pi210 & ~n41398;
  assign n41400 = pi146 & n41399;
  assign n41401 = ~pi234 & ~pi332;
  assign n41402 = ~n41360 & ~n41382;
  assign n41403 = ~pi95 & ~n41402;
  assign n41404 = n41292 & ~n41403;
  assign n41405 = n41365 & ~n41394;
  assign n41406 = ~n30614 & ~n41405;
  assign n41407 = pi137 & ~n41406;
  assign n41408 = pi210 & ~n41407;
  assign n41409 = ~n41404 & n41408;
  assign n41410 = n41401 & ~n41409;
  assign n41411 = ~n41301 & ~n41382;
  assign n41412 = ~pi95 & ~n41411;
  assign n41413 = ~n33962 & ~n41412;
  assign n41414 = ~pi137 & ~n41413;
  assign n41415 = ~n41397 & ~n41414;
  assign n41416 = n41371 & ~n41415;
  assign n41417 = n41410 & ~n41416;
  assign n41418 = ~n41400 & n41417;
  assign n41419 = ~n2811 & ~n41418;
  assign n41420 = ~n2811 & ~n41379;
  assign n41421 = ~n41418 & n41420;
  assign n41422 = ~n41379 & n41419;
  assign n41423 = ~n41399 & n41410;
  assign n41424 = ~n41356 & n41370;
  assign n41425 = n2811 & ~n41424;
  assign n41426 = n2811 & ~n41423;
  assign n41427 = ~n41424 & n41426;
  assign n41428 = ~n41423 & n41425;
  assign n41429 = ~pi153 & ~n64742;
  assign n41430 = ~n64741 & n41429;
  assign n41431 = ~n41298 & ~n41430;
  assign n41432 = ~pi228 & ~n41431;
  assign n41433 = ~pi216 & ~n41432;
  assign n41434 = ~pi105 & ~n41014;
  assign n41435 = ~pi332 & ~n64735;
  assign n41436 = ~n64734 & n41435;
  assign n41437 = n2811 & ~n41436;
  assign n41438 = pi146 & n41211;
  assign n41439 = ~pi146 & ~n41200;
  assign n41440 = ~n41199 & n41439;
  assign n41441 = n41358 & ~n41440;
  assign n41442 = ~n41438 & n41441;
  assign n41443 = pi146 & n41216;
  assign n41444 = ~pi146 & ~n41205;
  assign n41445 = ~n41204 & n41444;
  assign n41446 = n41401 & ~n41445;
  assign n41447 = n41401 & ~n41443;
  assign n41448 = ~n41445 & n41447;
  assign n41449 = ~n41443 & n41446;
  assign n41450 = ~n2811 & ~n64743;
  assign n41451 = ~n41442 & n41450;
  assign n41452 = ~n41437 & ~n41451;
  assign n41453 = pi105 & ~n41452;
  assign n41454 = ~n41434 & ~n41453;
  assign n41455 = pi228 & ~n41454;
  assign n41456 = ~pi228 & ~n41298;
  assign n41457 = ~pi228 & ~n41430;
  assign n41458 = ~n41298 & n41457;
  assign n41459 = ~n41430 & n41456;
  assign n41460 = ~n41455 & ~n64744;
  assign n41461 = ~pi216 & ~n41460;
  assign n41462 = ~n41224 & n41433;
  assign n41463 = ~n41009 & ~n64745;
  assign n41464 = ~pi221 & ~n41463;
  assign n41465 = ~n41027 & ~n41464;
  assign n41466 = ~pi215 & ~n41465;
  assign n41467 = pi299 & ~n41007;
  assign n41468 = ~n41466 & n41467;
  assign n41469 = ~pi224 & pi833;
  assign n41470 = pi222 & ~n41469;
  assign n41471 = ~pi223 & ~n41470;
  assign n41472 = n41006 & ~n41471;
  assign n41473 = pi224 & ~n41008;
  assign n41474 = ~pi222 & ~n41473;
  assign n41475 = ~pi332 & ~pi929;
  assign n41476 = n41469 & n41475;
  assign n41477 = ~n41474 & ~n41476;
  assign n41478 = ~pi223 & ~n41477;
  assign n41479 = ~n41472 & ~n41478;
  assign n41480 = ~pi299 & ~n41479;
  assign n41481 = ~pi223 & n2808;
  assign n41482 = pi198 & ~n41186;
  assign n41483 = ~pi198 & n64733;
  assign n41484 = ~n41482 & ~n41483;
  assign n41485 = pi234 & n41484;
  assign n41486 = pi198 & ~n41194;
  assign n41487 = ~pi198 & ~n41214;
  assign n41488 = ~n41486 & ~n41487;
  assign n41489 = ~pi234 & n41488;
  assign n41490 = ~pi332 & ~n41489;
  assign n41491 = ~n41485 & n41490;
  assign n41492 = n41481 & ~n41491;
  assign n41493 = ~pi198 & ~n41146;
  assign n41494 = ~pi142 & ~n41482;
  assign n41495 = ~n41493 & n41494;
  assign n41496 = pi142 & n41484;
  assign n41497 = n41358 & ~n41496;
  assign n41498 = n41358 & ~n41495;
  assign n41499 = ~n41496 & n41498;
  assign n41500 = ~n41495 & n41497;
  assign n41501 = ~pi223 & ~n2808;
  assign n41502 = ~pi198 & ~n41203;
  assign n41503 = ~pi142 & ~n41486;
  assign n41504 = ~pi142 & ~n41502;
  assign n41505 = ~n41486 & n41504;
  assign n41506 = ~n41502 & n41503;
  assign n41507 = pi142 & n41488;
  assign n41508 = n41401 & ~n41507;
  assign n41509 = n41401 & ~n64747;
  assign n41510 = ~n41507 & n41509;
  assign n41511 = ~n64747 & n41508;
  assign n41512 = n41501 & ~n64748;
  assign n41513 = ~n64746 & n41512;
  assign n41514 = ~n41492 & ~n41513;
  assign n41515 = n7034 & ~n41514;
  assign n41516 = n41480 & ~n41515;
  assign n41517 = ~pi39 & ~n41516;
  assign n41518 = ~n41468 & n41517;
  assign n41519 = n38189 & ~n41036;
  assign n41520 = ~n41479 & ~n41519;
  assign n41521 = ~pi299 & ~n41520;
  assign n41522 = pi105 & ~n41036;
  assign n41523 = pi228 & ~n41434;
  assign n41524 = ~n41522 & n41523;
  assign n41525 = ~pi137 & n62380;
  assign n41526 = ~pi153 & ~n41525;
  assign n41527 = ~pi228 & ~pi332;
  assign n41528 = pi137 & n62380;
  assign n41529 = n41527 & ~n41528;
  assign n41530 = ~n41526 & n41529;
  assign n41531 = ~pi216 & ~n41530;
  assign n41532 = ~n41434 & ~n41522;
  assign n41533 = pi228 & ~n41532;
  assign n41534 = ~pi137 & ~pi153;
  assign n41535 = ~pi332 & n41534;
  assign n41536 = ~pi332 & n62380;
  assign n41537 = n41534 & n41536;
  assign n41538 = n62380 & n41535;
  assign n41539 = n41014 & ~n41528;
  assign n41540 = ~pi228 & ~n41539;
  assign n41541 = ~n64749 & n41540;
  assign n41542 = ~n41533 & ~n41541;
  assign n41543 = ~pi216 & ~n41542;
  assign n41544 = ~n41524 & n41531;
  assign n41545 = ~n41009 & ~n64750;
  assign n41546 = ~pi221 & ~n41545;
  assign n41547 = ~n41027 & ~n41546;
  assign n41548 = ~pi215 & ~n41547;
  assign n41549 = ~n41007 & ~n41548;
  assign n41550 = pi299 & ~n41549;
  assign n41551 = ~n41521 & ~n41550;
  assign n41552 = pi39 & ~n41551;
  assign n41553 = ~pi38 & ~n41552;
  assign n41554 = ~n41518 & n41553;
  assign n41555 = n41030 & ~n41039;
  assign n41556 = pi299 & ~n41555;
  assign n41557 = ~n41521 & ~n41556;
  assign n41558 = ~pi39 & ~n41557;
  assign n41559 = n38189 & ~n41012;
  assign n41560 = n41480 & ~n41559;
  assign n41561 = pi299 & n41030;
  assign n41562 = ~n41560 & ~n41561;
  assign n41563 = pi39 & n41562;
  assign n41564 = pi38 & ~n41563;
  assign n41565 = ~n41558 & n41564;
  assign n41566 = ~pi100 & ~n41565;
  assign n41567 = ~n41554 & n41566;
  assign n41568 = ~pi210 & ~n30860;
  assign n41569 = pi95 & pi234;
  assign n41570 = ~pi137 & ~n41569;
  assign n41571 = ~pi137 & ~n41568;
  assign n41572 = ~n41569 & n41571;
  assign n41573 = ~n41568 & n41570;
  assign n41574 = pi105 & ~n64751;
  assign n41575 = ~n41034 & n41574;
  assign n41576 = ~n41034 & ~n64751;
  assign n41577 = ~pi332 & ~n41576;
  assign n41578 = pi105 & ~n41577;
  assign n41579 = n41523 & ~n41578;
  assign n41580 = n41046 & ~n41575;
  assign n41581 = ~pi153 & pi252;
  assign n41582 = ~pi137 & pi210;
  assign n41583 = ~pi252 & ~n41582;
  assign n41584 = n62380 & n41583;
  assign n41585 = ~n41581 & ~n41584;
  assign n41586 = ~n30860 & ~n41585;
  assign n41587 = n30860 & n41528;
  assign n41588 = n41527 & ~n41587;
  assign n41589 = ~n41526 & n41588;
  assign n41590 = ~pi252 & ~n30860;
  assign n41591 = n62380 & n41590;
  assign n41592 = pi153 & ~n41587;
  assign n41593 = ~n41591 & n41592;
  assign n41594 = pi252 & ~n30860;
  assign n41595 = n41571 & ~n41594;
  assign n41596 = n62380 & n41595;
  assign n41597 = ~n41593 & ~n41596;
  assign n41598 = n41527 & ~n41597;
  assign n41599 = ~n30860 & n41583;
  assign n41600 = n41536 & n41599;
  assign n41601 = n41014 & ~n41587;
  assign n41602 = ~n41600 & n41601;
  assign n41603 = ~n41568 & ~n41594;
  assign n41604 = n64749 & n41603;
  assign n41605 = ~n41602 & ~n41604;
  assign n41606 = ~pi228 & ~n41605;
  assign n41607 = ~n41586 & n41589;
  assign n41608 = ~pi216 & ~n64753;
  assign n41609 = ~n64752 & n41608;
  assign n41610 = ~n41009 & ~n41609;
  assign n41611 = ~pi221 & ~n41610;
  assign n41612 = ~n41027 & ~n41611;
  assign n41613 = ~pi215 & ~n41612;
  assign n41614 = ~n41007 & ~n41613;
  assign n41615 = pi299 & ~n41614;
  assign n41616 = pi142 & ~pi198;
  assign n41617 = ~pi137 & ~n41616;
  assign n41618 = ~n41034 & ~n41617;
  assign n41619 = n41012 & ~n41618;
  assign n41620 = n41501 & ~n41619;
  assign n41621 = ~pi137 & pi198;
  assign n41622 = ~pi95 & n41621;
  assign n41623 = ~n41031 & ~n41622;
  assign n41624 = n41358 & ~n41623;
  assign n41625 = n62380 & ~n41621;
  assign n41626 = n41401 & ~n41625;
  assign n41627 = n41481 & ~n41626;
  assign n41628 = ~n41624 & n41627;
  assign n41629 = ~n41620 & ~n41628;
  assign n41630 = n7034 & ~n41629;
  assign n41631 = ~n41479 & ~n41630;
  assign n41632 = ~pi299 & ~n41631;
  assign n41633 = n2764 & ~n41632;
  assign n41634 = ~n41615 & n41633;
  assign n41635 = ~n2764 & ~n41562;
  assign n41636 = pi100 & ~n41635;
  assign n41637 = ~n41634 & n41636;
  assign n41638 = ~pi87 & ~n41637;
  assign n41639 = ~n41567 & n41638;
  assign n41640 = ~n62373 & ~n41562;
  assign n41641 = n62373 & n41551;
  assign n41642 = ~n41640 & ~n41641;
  assign n41643 = pi87 & ~n41642;
  assign n41644 = ~pi75 & ~n41643;
  assign n41645 = ~n41639 & n41644;
  assign n41646 = n41016 & ~n64752;
  assign n41647 = ~n41009 & ~n41646;
  assign n41648 = ~pi221 & ~n41647;
  assign n41649 = ~n41027 & ~n41648;
  assign n41650 = ~pi215 & ~n41649;
  assign n41651 = ~n41007 & ~n41650;
  assign n41652 = pi299 & ~n41651;
  assign n41653 = n2806 & ~n41632;
  assign n41654 = ~n41652 & n41653;
  assign n41655 = ~n2806 & ~n41562;
  assign n41656 = pi75 & ~n41655;
  assign n41657 = ~n41654 & n41656;
  assign n41658 = ~n41645 & ~n41657;
  assign n41659 = ~pi92 & ~n41658;
  assign n41660 = n6795 & ~n41642;
  assign n41661 = ~n6795 & ~n41562;
  assign n41662 = pi92 & ~n41661;
  assign n41663 = ~n41660 & n41662;
  assign n41664 = ~pi54 & ~n41663;
  assign n41665 = ~n41659 & n41664;
  assign n41666 = ~n64081 & n41562;
  assign n41667 = n9738 & n41558;
  assign n41668 = ~n41666 & ~n41667;
  assign n41669 = pi54 & n41668;
  assign n41670 = ~pi74 & ~n41669;
  assign n41671 = ~n41665 & n41670;
  assign n41672 = ~pi54 & n41668;
  assign n41673 = pi54 & ~n41562;
  assign n41674 = pi74 & ~n41673;
  assign n41675 = ~n41672 & n41674;
  assign n41676 = ~n41671 & ~n41675;
  assign n41677 = ~pi55 & ~n41676;
  assign n41678 = ~pi332 & n41034;
  assign n41679 = pi105 & ~n41678;
  assign n41680 = n41523 & ~n41679;
  assign n41681 = ~pi228 & n41014;
  assign n41682 = ~n62380 & n41681;
  assign n41683 = ~pi216 & ~n41682;
  assign n41684 = ~n41680 & n41683;
  assign n41685 = ~n41009 & ~n41684;
  assign n41686 = ~pi221 & ~n41685;
  assign n41687 = ~n41027 & ~n41686;
  assign n41688 = ~pi215 & ~n41687;
  assign n41689 = n64082 & ~n41007;
  assign n41690 = ~n41688 & n41689;
  assign n41691 = ~n64082 & n41030;
  assign n41692 = pi55 & ~n41691;
  assign n41693 = ~n41690 & n41692;
  assign n41694 = ~pi56 & ~n41693;
  assign n41695 = ~n41677 & n41694;
  assign n41696 = ~n64084 & n41030;
  assign n41697 = n64084 & n41549;
  assign n41698 = ~n41696 & ~n41697;
  assign n41699 = pi56 & ~n41698;
  assign n41700 = ~pi62 & ~n41699;
  assign n41701 = ~n41695 & n41700;
  assign n41702 = ~pi56 & ~n41698;
  assign n41703 = pi56 & n41030;
  assign n41704 = pi62 & ~n41703;
  assign n41705 = ~n41702 & n41704;
  assign n41706 = ~pi59 & ~n41705;
  assign n41707 = ~n41701 & n41706;
  assign n41708 = pi59 & n41030;
  assign n41709 = ~n41040 & n41708;
  assign n41710 = ~pi57 & ~n41709;
  assign n41711 = ~n41707 & n41710;
  assign n41712 = ~n41043 & ~n41711;
  assign n41713 = n30877 & n40026;
  assign n41714 = n40161 & n41713;
  assign n41715 = pi24 & n62355;
  assign n41716 = ~n39175 & ~n41715;
  assign n41717 = pi24 & ~pi94;
  assign n41718 = ~n40118 & n41717;
  assign n41719 = pi252 & n38261;
  assign n41720 = ~pi252 & ~n34974;
  assign n41721 = pi252 & ~n38261;
  assign n41722 = ~pi252 & n34974;
  assign n41723 = ~n41721 & ~n41722;
  assign n41724 = ~n41719 & ~n41720;
  assign n41725 = n64196 & ~n64754;
  assign n41726 = ~n41718 & n41725;
  assign n41727 = ~n41716 & n41726;
  assign n41728 = pi24 & ~pi90;
  assign n41729 = n35400 & n41728;
  assign n41730 = n64754 & n41729;
  assign n41731 = n40120 & n41730;
  assign n41732 = ~n41727 & ~n41731;
  assign n41733 = ~pi100 & ~n41732;
  assign n41734 = pi100 & n64105;
  assign n41735 = n34139 & n41734;
  assign n41736 = ~n41733 & ~n41735;
  assign n41737 = ~pi75 & n30571;
  assign n41738 = n2764 & n6795;
  assign n41739 = ~n41736 & n64755;
  assign n41740 = ~n41714 & ~n41739;
  assign po208 = n40103 & ~n41740;
  assign n41742 = n2815 & n30864;
  assign n41743 = n64667 & ~n41742;
  assign n41744 = pi129 & ~n41743;
  assign n41745 = ~n64105 & ~n41744;
  assign n41746 = ~n2815 & n64667;
  assign n41747 = pi129 & ~n41746;
  assign n41748 = n2813 & ~n41747;
  assign n41749 = pi129 & ~n64667;
  assign n41750 = ~n30864 & ~n41749;
  assign n41751 = ~n30873 & ~n41750;
  assign n41752 = ~n41748 & n41751;
  assign n41753 = ~n30873 & ~n41745;
  assign n41754 = ~pi75 & n2805;
  assign n41755 = n30855 & n41754;
  assign n41756 = ~n64756 & n41755;
  assign n41757 = ~n38261 & n40027;
  assign n41758 = ~n40028 & n41757;
  assign n41759 = ~n41756 & ~n41758;
  assign n41760 = n40103 & ~n41759;
  assign po258 = n62380 & n41760;
  assign n41762 = pi51 & n2814;
  assign n41763 = ~pi146 & n41762;
  assign n41764 = pi161 & ~n41763;
  assign n41765 = n2597 & n35366;
  assign n41766 = ~pi51 & n41765;
  assign n41767 = n2814 & ~n41766;
  assign n41768 = pi51 & pi146;
  assign n41769 = n41767 & ~n41768;
  assign n41770 = ~n41764 & ~n41768;
  assign n41771 = n41767 & n41770;
  assign n41772 = ~n41764 & n41769;
  assign n41773 = ~pi87 & ~n64757;
  assign n41774 = pi87 & ~n32931;
  assign n41775 = pi232 & ~n41774;
  assign n41776 = ~n41773 & n41775;
  assign n41777 = ~pi134 & ~pi135;
  assign n41778 = ~pi136 & n41777;
  assign n41779 = ~pi130 & n41778;
  assign n41780 = ~pi132 & n41779;
  assign n41781 = ~pi126 & n41780;
  assign n41782 = ~pi121 & n41781;
  assign n41783 = ~pi125 & ~pi133;
  assign n41784 = pi121 & ~n41783;
  assign n41785 = ~pi121 & n41783;
  assign n41786 = ~n41784 & ~n41785;
  assign n41787 = ~n41782 & ~n41786;
  assign n41788 = ~pi87 & n41766;
  assign n41789 = ~n41787 & n41788;
  assign n41790 = ~n62455 & ~n41789;
  assign n41791 = ~n62455 & ~n41776;
  assign n41792 = ~n41789 & n41791;
  assign n41793 = ~n41776 & n41790;
  assign n41794 = pi299 & ~n64757;
  assign n41795 = ~pi142 & n41762;
  assign n41796 = pi144 & ~n41795;
  assign n41797 = pi51 & pi142;
  assign n41798 = n41767 & ~n41797;
  assign n41799 = ~n41796 & n41798;
  assign n41800 = ~pi299 & ~n41799;
  assign n41801 = pi232 & ~n41800;
  assign n41802 = pi232 & ~n41794;
  assign n41803 = ~n41800 & n41802;
  assign n41804 = ~n41794 & n41801;
  assign n41805 = pi38 & ~n64759;
  assign n41806 = ~pi100 & ~n41805;
  assign n41807 = pi38 & ~n41766;
  assign n41808 = ~pi100 & ~n41807;
  assign n41809 = ~n41806 & ~n41808;
  assign n41810 = n2599 & n30650;
  assign n41811 = n2588 & n2683;
  assign n41812 = n35365 & n41811;
  assign n41813 = n41810 & n41812;
  assign n41814 = pi77 & ~pi86;
  assign n41815 = n2588 & n35365;
  assign n41816 = n41810 & n41815;
  assign n41817 = ~pi50 & pi77;
  assign n41818 = n2638 & n41817;
  assign n41819 = n41816 & n41818;
  assign n41820 = n41813 & n41814;
  assign n41821 = ~pi24 & pi314;
  assign n41822 = n62767 & n41821;
  assign n41823 = ~pi24 & n62361;
  assign n41824 = ~pi94 & n41823;
  assign n41825 = ~pi24 & n62355;
  assign n41826 = pi314 & n62767;
  assign n41827 = n64761 & n41826;
  assign n41828 = n62355 & n41822;
  assign n41829 = n64760 & n64762;
  assign n41830 = n2728 & n41829;
  assign n41831 = ~n62767 & n41765;
  assign n41832 = ~pi51 & ~n41831;
  assign n41833 = n2684 & n41816;
  assign n41834 = ~pi77 & n41813;
  assign n41835 = pi86 & n64763;
  assign n41836 = ~n64760 & ~n41835;
  assign n41837 = n41715 & ~n41836;
  assign n41838 = pi86 & n62355;
  assign n41839 = ~pi24 & n41838;
  assign n41840 = n64761 & n41835;
  assign n41841 = n64763 & n41839;
  assign n41842 = n41765 & ~n64764;
  assign n41843 = ~n41837 & n41842;
  assign n41844 = n41832 & ~n41843;
  assign n41845 = n2728 & n41844;
  assign n41846 = n41766 & ~n41845;
  assign n41847 = ~pi58 & n62767;
  assign n41848 = n31434 & n41847;
  assign n41849 = n64763 & n41848;
  assign n41850 = pi72 & n2751;
  assign n41851 = n41849 & n41850;
  assign n41852 = n41846 & ~n41851;
  assign n41853 = ~n41830 & n41852;
  assign n41854 = ~n2814 & ~n41853;
  assign n41855 = n2861 & n41838;
  assign n41856 = ~pi24 & ~n41855;
  assign n41857 = n2665 & n35378;
  assign n41858 = pi24 & ~n41857;
  assign n41859 = ~n41856 & ~n41858;
  assign n41860 = ~pi314 & ~n41859;
  assign n41861 = pi314 & ~n41857;
  assign n41862 = ~n41860 & ~n41861;
  assign n41863 = n2695 & n62378;
  assign n41864 = n2696 & n62366;
  assign n41865 = n41862 & n64765;
  assign n41866 = ~pi51 & ~n41865;
  assign n41867 = pi72 & n39044;
  assign n41868 = n41866 & ~n41867;
  assign n41869 = n2814 & ~n41868;
  assign n41870 = ~n41854 & ~n41869;
  assign n41871 = pi142 & n41870;
  assign n41872 = ~n2814 & n41853;
  assign n41873 = n64089 & n41862;
  assign n41874 = ~pi72 & ~n41873;
  assign n41875 = n30619 & ~n41874;
  assign n41876 = n2814 & ~n41875;
  assign n41877 = ~n41872 & ~n41876;
  assign n41878 = ~pi142 & ~n41877;
  assign n41879 = ~pi144 & ~n41878;
  assign n41880 = ~pi144 & ~n41871;
  assign n41881 = ~n41878 & n41880;
  assign n41882 = ~n41871 & n41879;
  assign n41883 = n41796 & ~n41853;
  assign n41884 = ~pi180 & ~n41883;
  assign n41885 = ~n64766 & n41884;
  assign n41886 = n64089 & n41859;
  assign n41887 = ~pi72 & ~n41886;
  assign n41888 = n30619 & ~n41887;
  assign n41889 = n2814 & ~n41888;
  assign n41890 = ~n41872 & ~n41889;
  assign n41891 = ~pi142 & ~n41890;
  assign n41892 = n2728 & n2814;
  assign n41893 = n2726 & n32111;
  assign n41894 = n41886 & n64767;
  assign n41895 = ~n41762 & ~n41867;
  assign n41896 = n2814 & ~n41895;
  assign n41897 = ~n41894 & ~n41896;
  assign n41898 = ~n41854 & n41897;
  assign n41899 = pi142 & n41898;
  assign n41900 = ~pi144 & ~n41899;
  assign n41901 = ~n41891 & n41900;
  assign n41902 = ~pi51 & ~n41765;
  assign n41903 = n2814 & n41902;
  assign n41904 = ~n64767 & ~n41903;
  assign n41905 = n2728 & ~n41844;
  assign n41906 = ~n41904 & ~n41905;
  assign n41907 = pi142 & ~n41906;
  assign n41908 = n2814 & ~n41846;
  assign n41909 = ~pi142 & ~n41908;
  assign n41910 = ~n41907 & ~n41909;
  assign n41911 = n41766 & ~n41830;
  assign n41912 = ~n41845 & n41911;
  assign n41913 = ~n2814 & ~n41912;
  assign n41914 = ~n41767 & ~n41913;
  assign n41915 = ~n41910 & ~n41914;
  assign n41916 = ~pi51 & n2814;
  assign n41917 = ~n41852 & n41916;
  assign n41918 = ~n41854 & ~n41917;
  assign n41919 = ~n41915 & n41918;
  assign n41920 = pi144 & ~n41919;
  assign n41921 = pi180 & ~n41920;
  assign n41922 = ~n41901 & n41921;
  assign n41923 = ~pi179 & ~n41922;
  assign n41924 = ~n64766 & ~n41883;
  assign n41925 = ~pi180 & ~n41924;
  assign n41926 = ~pi142 & n41890;
  assign n41927 = pi142 & ~n41898;
  assign n41928 = ~pi144 & ~n41927;
  assign n41929 = ~n41926 & n41928;
  assign n41930 = pi144 & n41918;
  assign n41931 = ~n41915 & n41930;
  assign n41932 = pi180 & ~n41931;
  assign n41933 = ~n41929 & n41932;
  assign n41934 = ~n41925 & ~n41933;
  assign n41935 = ~pi179 & ~n41934;
  assign n41936 = ~n41885 & n41923;
  assign n41937 = n64093 & n34954;
  assign n41938 = ~pi24 & ~pi51;
  assign n41939 = n41826 & n41938;
  assign n41940 = ~pi51 & n41822;
  assign n41941 = n64089 & n41821;
  assign n41942 = n41937 & n64769;
  assign n41943 = n64767 & n41942;
  assign n41944 = ~n41854 & ~n41896;
  assign n41945 = ~n41943 & n41944;
  assign n41946 = pi142 & n41945;
  assign n41947 = ~pi72 & ~n41942;
  assign n41948 = n30619 & ~n41947;
  assign n41949 = n2814 & ~n41948;
  assign n41950 = ~n41872 & ~n41949;
  assign n41951 = ~pi142 & ~n41950;
  assign n41952 = ~pi144 & ~n41951;
  assign n41953 = ~n41946 & n41952;
  assign n41954 = ~n41851 & n41914;
  assign n41955 = ~n41830 & n41954;
  assign n41956 = n41796 & ~n41955;
  assign n41957 = ~pi180 & ~n41956;
  assign n41958 = ~n41953 & n41957;
  assign n41959 = ~pi144 & n41944;
  assign n41960 = pi144 & n41954;
  assign n41961 = ~n41795 & ~n41960;
  assign n41962 = pi144 & ~n41954;
  assign n41963 = ~pi144 & ~n41944;
  assign n41964 = ~n41962 & ~n41963;
  assign n41965 = ~n41795 & ~n41964;
  assign n41966 = ~n41959 & n41961;
  assign n41967 = pi180 & ~n64770;
  assign n41968 = pi179 & ~n41967;
  assign n41969 = pi179 & ~n41958;
  assign n41970 = ~n41967 & n41969;
  assign n41971 = ~n41958 & n41968;
  assign n41972 = ~n64768 & ~n64771;
  assign n41973 = ~pi299 & ~n41972;
  assign n41974 = ~pi161 & ~n41763;
  assign n41975 = ~n41944 & n41974;
  assign n41976 = pi146 & n41954;
  assign n41977 = n41765 & ~n41851;
  assign n41978 = n41916 & ~n41977;
  assign n41979 = ~pi146 & ~n41978;
  assign n41980 = ~n41854 & n41979;
  assign n41981 = pi161 & ~n41980;
  assign n41982 = pi161 & ~n41976;
  assign n41983 = ~n41980 & n41982;
  assign n41984 = ~n41976 & n41981;
  assign n41985 = ~n41975 & ~n64772;
  assign n41986 = n33497 & ~n41985;
  assign n41987 = pi146 & n41945;
  assign n41988 = ~pi146 & ~n41950;
  assign n41989 = ~pi161 & ~n41988;
  assign n41990 = ~n41987 & n41989;
  assign n41991 = n41916 & n41977;
  assign n41992 = ~n41830 & n41991;
  assign n41993 = ~n41762 & ~n41992;
  assign n41994 = pi146 & ~n41766;
  assign n41995 = ~n41993 & ~n41994;
  assign n41996 = pi161 & ~n41995;
  assign n41997 = ~n41872 & n41996;
  assign n41998 = ~n41990 & ~n41997;
  assign n41999 = n33512 & ~n41998;
  assign n42000 = ~n41986 & ~n41999;
  assign n42001 = pi156 & ~n42000;
  assign n42002 = pi146 & n41870;
  assign n42003 = ~pi146 & ~n41877;
  assign n42004 = n33512 & ~n42003;
  assign n42005 = n33512 & ~n42002;
  assign n42006 = ~n42003 & n42005;
  assign n42007 = ~n42002 & n42004;
  assign n42008 = ~pi146 & ~n41890;
  assign n42009 = pi146 & n41898;
  assign n42010 = n33497 & ~n42009;
  assign n42011 = ~n42008 & n42010;
  assign n42012 = ~pi161 & ~n42011;
  assign n42013 = ~n64773 & n42012;
  assign n42014 = pi146 & ~n41906;
  assign n42015 = ~pi146 & ~n41908;
  assign n42016 = ~n42014 & ~n42015;
  assign n42017 = ~n41914 & ~n42016;
  assign n42018 = n41918 & ~n42017;
  assign n42019 = n33497 & ~n42018;
  assign n42020 = n33512 & ~n41763;
  assign n42021 = ~n41853 & n42020;
  assign n42022 = pi161 & ~n42021;
  assign n42023 = ~n42019 & n42022;
  assign n42024 = ~pi156 & ~n42023;
  assign n42025 = ~n42013 & n42024;
  assign n42026 = ~n42001 & ~n42025;
  assign n42027 = ~n41973 & n42026;
  assign n42028 = n32271 & ~n42027;
  assign n42029 = n2728 & n41849;
  assign n42030 = n41766 & ~n42029;
  assign n42031 = ~n41763 & ~n42030;
  assign n42032 = pi161 & ~n42031;
  assign n42033 = ~n2814 & ~n42030;
  assign n42034 = n62364 & n62378;
  assign n42035 = n62365 & n62366;
  assign n42036 = ~pi51 & ~n64774;
  assign n42037 = n2814 & ~n42036;
  assign n42038 = ~n42033 & ~n42037;
  assign n42039 = pi146 & ~n42038;
  assign n42040 = ~n32270 & ~n42033;
  assign n42041 = ~pi146 & ~n42040;
  assign n42042 = ~pi161 & ~n42041;
  assign n42043 = ~pi161 & ~n42039;
  assign n42044 = ~n42041 & n42043;
  assign n42045 = ~n42039 & n42042;
  assign n42046 = ~n42032 & ~n64775;
  assign n42047 = n2960 & ~n42046;
  assign n42048 = ~n31886 & ~n42047;
  assign n42049 = ~pi287 & n2814;
  assign n42050 = ~pi51 & n42049;
  assign n42051 = ~n42038 & ~n42050;
  assign n42052 = n41974 & n42051;
  assign n42053 = n42029 & ~n42049;
  assign n42054 = n41766 & ~n42053;
  assign n42055 = n41764 & ~n42054;
  assign n42056 = ~n42052 & ~n42055;
  assign n42057 = pi216 & ~n42056;
  assign n42058 = ~n42048 & ~n42057;
  assign n42059 = ~n41766 & ~n64757;
  assign n42060 = ~n2960 & ~n42059;
  assign n42061 = n31761 & ~n42060;
  assign n42062 = ~n42058 & n42061;
  assign n42063 = ~pi51 & ~n42030;
  assign n42064 = ~pi287 & ~n42063;
  assign n42065 = ~n41903 & ~n42049;
  assign n42066 = ~n42064 & ~n42065;
  assign n42067 = ~n41798 & ~n42066;
  assign n42068 = n31926 & ~n42067;
  assign n42069 = pi181 & n41765;
  assign n42070 = n42068 & n42069;
  assign n42071 = ~n41766 & ~n41795;
  assign n42072 = ~n2980 & ~n42071;
  assign n42073 = pi144 & ~n42072;
  assign n42074 = pi51 & ~n2814;
  assign n42075 = ~n42063 & ~n42074;
  assign n42076 = n2980 & ~n41797;
  assign n42077 = n42075 & n42076;
  assign n42078 = n42073 & ~n42077;
  assign n42079 = ~n42070 & n42078;
  assign n42080 = pi142 & n42038;
  assign n42081 = pi181 & pi224;
  assign n42082 = ~pi142 & n42040;
  assign n42083 = ~n42081 & ~n42082;
  assign n42084 = ~n42080 & n42083;
  assign n42085 = ~n41795 & n42081;
  assign n42086 = n42051 & n42085;
  assign n42087 = n2980 & ~n42086;
  assign n42088 = ~n42084 & n42087;
  assign n42089 = ~n2980 & n41903;
  assign n42090 = ~n42072 & ~n42089;
  assign n42091 = ~n42073 & n42090;
  assign n42092 = ~n42088 & n42091;
  assign n42093 = ~n42079 & ~n42092;
  assign n42094 = pi142 & ~n42038;
  assign n42095 = ~pi142 & ~n42040;
  assign n42096 = n2980 & ~n42095;
  assign n42097 = n2980 & ~n42094;
  assign n42098 = ~n42095 & n42097;
  assign n42099 = ~n42094 & n42096;
  assign n42100 = ~n31926 & ~n64776;
  assign n42101 = pi224 & ~n41795;
  assign n42102 = n42051 & n42101;
  assign n42103 = ~n42100 & ~n42102;
  assign n42104 = n42091 & ~n42103;
  assign n42105 = n41765 & n42068;
  assign n42106 = n42078 & ~n42105;
  assign n42107 = pi181 & ~n42106;
  assign n42108 = ~n42104 & n42107;
  assign n42109 = n42091 & ~n64776;
  assign n42110 = ~pi181 & ~n42078;
  assign n42111 = ~n42109 & n42110;
  assign n42112 = ~pi299 & ~n42111;
  assign n42113 = ~n42108 & n42112;
  assign n42114 = ~pi299 & ~n42093;
  assign n42115 = n31784 & ~n42060;
  assign n42116 = ~n42047 & n42115;
  assign n42117 = pi232 & ~n42116;
  assign n42118 = ~n64777 & n42117;
  assign n42119 = ~n42062 & n42117;
  assign n42120 = ~n64777 & n42119;
  assign n42121 = ~n42062 & n42118;
  assign n42122 = ~n2961 & ~n62403;
  assign n42123 = n42029 & ~n42122;
  assign n42124 = ~pi232 & n41766;
  assign n42125 = ~n42123 & n42124;
  assign n42126 = pi39 & ~n42125;
  assign n42127 = ~n64778 & n42126;
  assign n42128 = ~pi39 & ~pi232;
  assign n42129 = ~n41853 & n42128;
  assign n42130 = ~n42127 & ~n42129;
  assign n42131 = ~n42028 & n42130;
  assign n42132 = ~pi38 & ~n42131;
  assign n42133 = ~n41809 & ~n42132;
  assign n42134 = pi100 & n64759;
  assign n42135 = pi100 & n41766;
  assign n42136 = n6797 & ~n42135;
  assign n42137 = ~n42134 & n42136;
  assign n42138 = ~n42133 & n42137;
  assign n42139 = ~pi87 & ~n6794;
  assign n42140 = ~n41766 & n42139;
  assign n42141 = ~n64759 & n42140;
  assign n42142 = ~pi184 & ~pi299;
  assign n42143 = ~n36984 & ~n42142;
  assign n42144 = n2815 & n42143;
  assign n42145 = pi87 & ~n42144;
  assign n42146 = ~n41787 & ~n42145;
  assign n42147 = ~n42141 & n42146;
  assign n42148 = ~n42138 & n42147;
  assign n42149 = n2814 & ~n41866;
  assign n42150 = ~n41797 & n42149;
  assign n42151 = pi144 & ~n42150;
  assign n42152 = n41765 & ~n41829;
  assign n42153 = n62767 & n42152;
  assign n42154 = n41843 & n42153;
  assign n42155 = n41832 & ~n42154;
  assign n42156 = n2728 & ~n42155;
  assign n42157 = ~n41904 & ~n42156;
  assign n42158 = pi142 & n42157;
  assign n42159 = n2814 & ~n41912;
  assign n42160 = ~pi142 & n42159;
  assign n42161 = ~pi144 & ~n42160;
  assign n42162 = ~pi144 & ~n42158;
  assign n42163 = ~n42160 & n42162;
  assign n42164 = ~n42158 & n42161;
  assign n42165 = pi180 & ~n64779;
  assign n42166 = ~n42151 & n42165;
  assign n42167 = n41796 & ~n41894;
  assign n42168 = ~pi144 & ~n41910;
  assign n42169 = ~pi180 & ~n42168;
  assign n42170 = ~n42167 & n42169;
  assign n42171 = pi179 & ~n42170;
  assign n42172 = ~n42166 & n42171;
  assign n42173 = n41796 & ~n41943;
  assign n42174 = ~pi51 & ~n42152;
  assign n42175 = n2728 & ~n42174;
  assign n42176 = ~n41904 & ~n42175;
  assign n42177 = pi142 & n42176;
  assign n42178 = n2814 & ~n41911;
  assign n42179 = ~pi142 & n42178;
  assign n42180 = ~pi144 & ~n42179;
  assign n42181 = ~n42177 & n42180;
  assign n42182 = pi180 & ~n42181;
  assign n42183 = ~n42173 & n42182;
  assign n42184 = ~pi180 & n41799;
  assign n42185 = ~pi179 & ~n42184;
  assign n42186 = ~n42183 & n42185;
  assign n42187 = ~n42172 & ~n42186;
  assign n42188 = ~pi299 & ~n42187;
  assign n42189 = ~n41768 & n42149;
  assign n42190 = pi161 & ~n42189;
  assign n42191 = ~pi146 & n42159;
  assign n42192 = pi146 & n42157;
  assign n42193 = ~pi161 & ~n42192;
  assign n42194 = ~pi161 & ~n42191;
  assign n42195 = ~n42192 & n42194;
  assign n42196 = ~n42191 & n42193;
  assign n42197 = ~n42190 & ~n64780;
  assign n42198 = n33497 & ~n42197;
  assign n42199 = n41764 & ~n41894;
  assign n42200 = ~pi161 & ~n42016;
  assign n42201 = ~n42199 & ~n42200;
  assign n42202 = n33512 & ~n42201;
  assign n42203 = pi232 & ~n42202;
  assign n42204 = ~n42198 & n42203;
  assign n42205 = pi156 & ~n42204;
  assign n42206 = ~pi39 & ~n42205;
  assign n42207 = ~pi39 & ~n42188;
  assign n42208 = ~n42205 & n42207;
  assign n42209 = ~n42188 & n42206;
  assign n42210 = ~pi144 & ~n41798;
  assign n42211 = ~n42068 & n42210;
  assign n42212 = n31926 & n42049;
  assign n42213 = ~n41797 & n42212;
  assign n42214 = n64774 & n42049;
  assign n42215 = n31926 & ~n41797;
  assign n42216 = n42214 & n42215;
  assign n42217 = ~pi142 & ~n64774;
  assign n42218 = pi142 & ~n62380;
  assign n42219 = n42212 & ~n42218;
  assign n42220 = ~n42217 & n42219;
  assign n42221 = n42212 & ~n42217;
  assign n42222 = ~n42218 & n42221;
  assign n42223 = n64774 & n42213;
  assign n42224 = n41796 & ~n64782;
  assign n42225 = pi181 & ~n42224;
  assign n42226 = pi181 & ~n42211;
  assign n42227 = ~n42224 & n42226;
  assign n42228 = ~n42211 & n42225;
  assign n42229 = ~pi181 & n41799;
  assign n42230 = ~pi299 & ~n42229;
  assign n42231 = ~n64783 & n42230;
  assign n42232 = n2814 & n2933;
  assign n42233 = n41764 & ~n42232;
  assign n42234 = pi159 & n31886;
  assign n42235 = n41974 & ~n42066;
  assign n42236 = n42234 & ~n42235;
  assign n42237 = ~n42233 & n42236;
  assign n42238 = n64757 & ~n42234;
  assign n42239 = pi299 & ~n42238;
  assign n42240 = ~n42237 & n42239;
  assign n42241 = n31886 & ~n42235;
  assign n42242 = ~n42233 & n42241;
  assign n42243 = ~n31886 & n64757;
  assign n42244 = n31761 & ~n42243;
  assign n42245 = ~n42242 & n42244;
  assign n42246 = ~pi159 & n41794;
  assign n42247 = n33664 & ~n42246;
  assign n42248 = ~n42245 & n42247;
  assign n42249 = n33664 & ~n42240;
  assign n42250 = ~n42231 & n64784;
  assign n42251 = ~pi38 & ~n42250;
  assign n42252 = ~n64781 & n42251;
  assign n42253 = n41764 & ~n41943;
  assign n42254 = pi146 & n42176;
  assign n42255 = ~pi146 & n42178;
  assign n42256 = ~pi161 & ~n42255;
  assign n42257 = ~n42254 & n42256;
  assign n42258 = ~n42253 & ~n42257;
  assign n42259 = n33497 & ~n42258;
  assign n42260 = ~pi158 & n41794;
  assign n42261 = pi232 & ~n42260;
  assign n42262 = ~n42259 & n42261;
  assign n42263 = ~pi156 & n2764;
  assign n42264 = ~n42262 & n42263;
  assign n42265 = n41806 & ~n42264;
  assign n42266 = ~n42252 & n42265;
  assign n42267 = n6797 & ~n42134;
  assign n42268 = ~n42266 & n42267;
  assign n42269 = ~n64759 & n42139;
  assign n42270 = n41787 & ~n42145;
  assign n42271 = ~n42269 & n42270;
  assign n42272 = ~n42268 & n42271;
  assign n42273 = n62455 & ~n42272;
  assign n42274 = ~n42148 & n42273;
  assign n42275 = ~n64758 & ~n42274;
  assign n42276 = ~pi125 & n41782;
  assign n42277 = pi125 & pi133;
  assign n42278 = ~n41783 & ~n42277;
  assign n42279 = ~n42276 & ~n42278;
  assign n42280 = n41766 & ~n42279;
  assign n42281 = pi172 & n41762;
  assign n42282 = ~pi152 & n41903;
  assign n42283 = ~n42281 & ~n42282;
  assign n42284 = pi232 & ~n42283;
  assign n42285 = ~n42280 & ~n42284;
  assign n42286 = ~pi87 & ~n42285;
  assign n42287 = pi87 & n2815;
  assign n42288 = pi162 & n42287;
  assign n42289 = ~n62455 & ~n42288;
  assign n42290 = ~n42286 & n42289;
  assign n42291 = ~pi152 & n2814;
  assign n42292 = n41867 & ~n42291;
  assign n42293 = ~pi152 & n41978;
  assign n42294 = ~pi197 & ~n42293;
  assign n42295 = ~n42292 & n42294;
  assign n42296 = ~n2814 & n41867;
  assign n42297 = ~n41916 & ~n42296;
  assign n42298 = ~n41992 & ~n42297;
  assign n42299 = ~pi152 & pi197;
  assign n42300 = ~n42298 & n42299;
  assign n42301 = ~n42295 & ~n42300;
  assign n42302 = ~n42281 & ~n42301;
  assign n42303 = ~n2814 & ~n41867;
  assign n42304 = ~n41949 & ~n42303;
  assign n42305 = ~pi172 & n42304;
  assign n42306 = ~n41762 & ~n41943;
  assign n42307 = ~n41867 & n42306;
  assign n42308 = n41895 & ~n41943;
  assign n42309 = pi172 & ~n64785;
  assign n42310 = pi152 & pi197;
  assign n42311 = ~n42309 & n42310;
  assign n42312 = ~n42305 & n42311;
  assign n42313 = ~n42302 & ~n42312;
  assign n42314 = n31909 & ~n42313;
  assign n42315 = ~n41876 & ~n42303;
  assign n42316 = ~pi172 & n42315;
  assign n42317 = ~n41868 & ~n42303;
  assign n42318 = pi172 & n42317;
  assign n42319 = pi152 & ~n42318;
  assign n42320 = ~n42316 & n42319;
  assign n42321 = n2814 & n41853;
  assign n42322 = ~n42297 & ~n42321;
  assign n42323 = ~pi152 & ~n42281;
  assign n42324 = ~n42322 & n42323;
  assign n42325 = pi197 & ~n42324;
  assign n42326 = ~n42281 & ~n42322;
  assign n42327 = ~pi152 & ~n42326;
  assign n42328 = ~pi172 & ~n42315;
  assign n42329 = pi172 & ~n42317;
  assign n42330 = pi152 & ~n42329;
  assign n42331 = ~n42328 & n42330;
  assign n42332 = ~n42327 & ~n42331;
  assign n42333 = pi197 & ~n42332;
  assign n42334 = ~n42320 & n42325;
  assign n42335 = ~n41889 & ~n42303;
  assign n42336 = pi152 & n42335;
  assign n42337 = ~n41917 & ~n42296;
  assign n42338 = ~pi152 & ~n42337;
  assign n42339 = ~pi172 & ~n42338;
  assign n42340 = ~n42336 & n42339;
  assign n42341 = ~n41894 & n41895;
  assign n42342 = pi152 & ~n42341;
  assign n42343 = n41852 & n41991;
  assign n42344 = n41846 & n41991;
  assign n42345 = ~n42303 & ~n64787;
  assign n42346 = ~pi152 & n42345;
  assign n42347 = pi172 & ~n42346;
  assign n42348 = ~n42342 & n42347;
  assign n42349 = ~pi197 & ~n42348;
  assign n42350 = ~n42340 & n42349;
  assign n42351 = n31918 & ~n42350;
  assign n42352 = ~n64786 & n42351;
  assign n42353 = ~n42314 & ~n42352;
  assign n42354 = pi299 & ~n42353;
  assign n42355 = pi145 & n42304;
  assign n42356 = ~pi145 & n41867;
  assign n42357 = pi174 & ~n42356;
  assign n42358 = ~n42355 & n42357;
  assign n42359 = pi145 & n42298;
  assign n42360 = ~n41978 & ~n42296;
  assign n42361 = ~pi145 & ~n42360;
  assign n42362 = ~pi174 & ~n42361;
  assign n42363 = ~n42359 & n42362;
  assign n42364 = ~n42358 & ~n42363;
  assign n42365 = ~pi193 & ~n42364;
  assign n42366 = ~pi145 & n41943;
  assign n42367 = pi174 & ~n64785;
  assign n42368 = ~n42306 & ~n42366;
  assign n42369 = ~n41867 & ~n42368;
  assign n42370 = pi174 & ~n42369;
  assign n42371 = ~n42366 & n42367;
  assign n42372 = ~n41762 & ~n41830;
  assign n42373 = pi145 & ~n42372;
  assign n42374 = n41991 & ~n42373;
  assign n42375 = ~pi174 & ~n42374;
  assign n42376 = ~n42303 & n42375;
  assign n42377 = pi193 & ~n42376;
  assign n42378 = ~n64788 & n42377;
  assign n42379 = ~n42365 & ~n42378;
  assign n42380 = n31935 & ~n42379;
  assign n42381 = pi145 & n42315;
  assign n42382 = ~pi145 & n42335;
  assign n42383 = ~pi193 & ~n42382;
  assign n42384 = ~n42381 & n42383;
  assign n42385 = pi145 & n42317;
  assign n42386 = ~pi145 & ~n42341;
  assign n42387 = pi193 & ~n42386;
  assign n42388 = ~n42385 & n42387;
  assign n42389 = pi174 & ~n42388;
  assign n42390 = pi145 & ~n42317;
  assign n42391 = ~pi145 & n42341;
  assign n42392 = pi193 & ~n42391;
  assign n42393 = ~n42390 & n42392;
  assign n42394 = pi145 & ~n42315;
  assign n42395 = ~pi145 & ~n42335;
  assign n42396 = ~pi193 & ~n42395;
  assign n42397 = ~n42394 & n42396;
  assign n42398 = ~n42393 & ~n42397;
  assign n42399 = pi174 & ~n42398;
  assign n42400 = ~n42384 & n42389;
  assign n42401 = pi193 & n41762;
  assign n42402 = pi145 & ~n42401;
  assign n42403 = ~n42322 & n42402;
  assign n42404 = ~pi193 & ~n42337;
  assign n42405 = pi193 & n42345;
  assign n42406 = ~pi145 & ~n42405;
  assign n42407 = ~pi145 & ~n42404;
  assign n42408 = ~n42405 & n42407;
  assign n42409 = ~n42404 & n42406;
  assign n42410 = ~pi174 & ~n64790;
  assign n42411 = ~pi174 & ~n42403;
  assign n42412 = ~n64790 & n42411;
  assign n42413 = ~n42403 & n42410;
  assign n42414 = n31955 & ~n64791;
  assign n42415 = ~n64789 & n42414;
  assign n42416 = ~n42380 & ~n42415;
  assign n42417 = ~pi38 & ~n42416;
  assign n42418 = ~n42354 & ~n42417;
  assign n42419 = n32271 & ~n42418;
  assign n42420 = ~pi299 & ~n3076;
  assign n42421 = pi299 & ~n3056;
  assign n42422 = ~n42420 & ~n42421;
  assign n42423 = ~n62401 & ~n62404;
  assign n42424 = n62380 & n64792;
  assign n42425 = ~pi232 & ~n42424;
  assign n42426 = pi39 & ~n42425;
  assign n42427 = ~n41762 & ~n42214;
  assign n42428 = pi224 & n42427;
  assign n42429 = n2980 & ~n42428;
  assign n42430 = n62380 & ~n2814;
  assign n42431 = ~n42037 & ~n42430;
  assign n42432 = ~n42036 & ~n42074;
  assign n42433 = n3076 & n64793;
  assign n42434 = n42429 & ~n42433;
  assign n42435 = ~n41762 & ~n42434;
  assign n42436 = pi174 & ~n42435;
  assign n42437 = n2814 & ~n42030;
  assign n42438 = ~n42430 & ~n42437;
  assign n42439 = n3076 & n42438;
  assign n42440 = n42029 & n42049;
  assign n42441 = pi224 & ~n42440;
  assign n42442 = n2980 & ~n42441;
  assign n42443 = ~n41767 & ~n42442;
  assign n42444 = ~n42439 & ~n42443;
  assign n42445 = ~pi174 & n42444;
  assign n42446 = pi193 & ~n42445;
  assign n42447 = ~n42436 & n42446;
  assign n42448 = n2814 & n42063;
  assign n42449 = ~n42430 & ~n42448;
  assign n42450 = ~pi224 & n42449;
  assign n42451 = pi224 & ~n42066;
  assign n42452 = n2980 & ~n42451;
  assign n42453 = ~n42450 & n42452;
  assign n42454 = ~n42089 & ~n42453;
  assign n42455 = ~pi174 & ~n42454;
  assign n42456 = ~n3076 & ~n42212;
  assign n42457 = n62380 & ~n42456;
  assign n42458 = pi174 & n42457;
  assign n42459 = ~pi193 & ~n42458;
  assign n42460 = ~n42455 & n42459;
  assign n42461 = pi180 & ~n42460;
  assign n42462 = ~n42447 & n42461;
  assign n42463 = ~n3076 & ~n41767;
  assign n42464 = ~n42449 & ~n42463;
  assign n42465 = ~pi174 & n42464;
  assign n42466 = n3076 & n64774;
  assign n42467 = ~pi51 & n42466;
  assign n42468 = n62380 & n3076;
  assign n42469 = pi174 & n64794;
  assign n42470 = ~n42401 & ~n42469;
  assign n42471 = ~n42401 & ~n42465;
  assign n42472 = ~n42469 & n42471;
  assign n42473 = ~n42465 & n42470;
  assign n42474 = ~pi180 & ~n64795;
  assign n42475 = ~pi299 & ~n42474;
  assign n42476 = ~n42462 & n42475;
  assign n42477 = ~n3056 & n42283;
  assign n42478 = pi152 & n64793;
  assign n42479 = ~pi152 & n42438;
  assign n42480 = pi51 & ~pi172;
  assign n42481 = ~n42479 & ~n42480;
  assign n42482 = ~n42478 & ~n42480;
  assign n42483 = ~n42479 & n42482;
  assign n42484 = ~pi152 & ~n42438;
  assign n42485 = pi152 & ~n64793;
  assign n42486 = ~n42484 & ~n42485;
  assign n42487 = ~n42480 & ~n42486;
  assign n42488 = ~n42478 & n42481;
  assign n42489 = ~pi216 & ~n64796;
  assign n42490 = n2960 & n42489;
  assign n42491 = ~n42477 & ~n42490;
  assign n42492 = n33512 & ~n42491;
  assign n42493 = pi152 & ~n42232;
  assign n42494 = ~pi152 & ~n42066;
  assign n42495 = ~pi172 & ~n42494;
  assign n42496 = ~n42493 & n42495;
  assign n42497 = pi152 & n42427;
  assign n42498 = ~n41767 & ~n42440;
  assign n42499 = ~pi152 & n42498;
  assign n42500 = pi172 & ~n42499;
  assign n42501 = ~n42497 & n42500;
  assign n42502 = pi216 & ~n42501;
  assign n42503 = pi152 & ~n42427;
  assign n42504 = ~pi152 & ~n42498;
  assign n42505 = pi172 & ~n42504;
  assign n42506 = ~n42503 & n42505;
  assign n42507 = pi152 & n42232;
  assign n42508 = ~pi152 & n42066;
  assign n42509 = ~pi172 & ~n42508;
  assign n42510 = ~n42507 & n42509;
  assign n42511 = ~n42506 & ~n42510;
  assign n42512 = pi216 & ~n42511;
  assign n42513 = pi216 & ~n42496;
  assign n42514 = ~n42501 & n42513;
  assign n42515 = ~n42496 & n42502;
  assign n42516 = n2960 & ~n42489;
  assign n42517 = n2960 & ~n64797;
  assign n42518 = ~n42489 & n42517;
  assign n42519 = ~n64797 & n42516;
  assign n42520 = ~n2960 & ~n42283;
  assign n42521 = n33497 & ~n42520;
  assign n42522 = ~n64798 & n42521;
  assign n42523 = ~n42492 & ~n42522;
  assign n42524 = ~n42476 & ~n42522;
  assign n42525 = ~n42492 & n42524;
  assign n42526 = ~n42476 & n42523;
  assign n42527 = pi232 & ~n64799;
  assign n42528 = n42426 & ~n42527;
  assign n42529 = ~pi232 & ~n41867;
  assign n42530 = ~pi39 & ~n42529;
  assign n42531 = ~pi38 & ~n42530;
  assign n42532 = ~n42528 & n42531;
  assign n42533 = pi299 & n42283;
  assign n42534 = ~pi174 & n41903;
  assign n42535 = ~pi299 & ~n42401;
  assign n42536 = ~n42534 & n42535;
  assign n42537 = pi232 & ~n42536;
  assign n42538 = ~n42533 & n42537;
  assign n42539 = pi38 & ~n42538;
  assign n42540 = ~pi100 & ~n42539;
  assign n42541 = ~n42532 & n42540;
  assign n42542 = ~n42419 & n42541;
  assign n42543 = pi100 & n42538;
  assign n42544 = n6797 & ~n42543;
  assign n42545 = ~n42542 & n42544;
  assign n42546 = n42139 & ~n42538;
  assign n42547 = pi140 & ~pi299;
  assign n42548 = ~n36868 & ~n42547;
  assign n42549 = n2815 & ~n42548;
  assign n42550 = pi87 & ~n42549;
  assign n42551 = n42279 & ~n42550;
  assign n42552 = ~n42546 & n42551;
  assign n42553 = ~n42545 & n42552;
  assign n42554 = ~pi232 & ~n41912;
  assign n42555 = ~pi39 & ~n42554;
  assign n42556 = n31926 & n42029;
  assign n42557 = n41766 & ~n42556;
  assign n42558 = ~pi299 & ~n42557;
  assign n42559 = n31886 & n42029;
  assign n42560 = n41766 & ~n42559;
  assign n42561 = pi299 & ~n42560;
  assign n42562 = ~n42558 & ~n42561;
  assign n42563 = ~pi232 & ~n42562;
  assign n42564 = pi39 & ~n42563;
  assign n42565 = ~n41766 & n42283;
  assign n42566 = ~n31886 & ~n42565;
  assign n42567 = n42051 & n42323;
  assign n42568 = pi152 & ~n42281;
  assign n42569 = ~n42054 & n42568;
  assign n42570 = n31886 & ~n42569;
  assign n42571 = ~pi152 & ~n42051;
  assign n42572 = pi152 & n42054;
  assign n42573 = ~n42281 & ~n42572;
  assign n42574 = ~n42571 & n42573;
  assign n42575 = n31886 & ~n42574;
  assign n42576 = ~n42567 & n42570;
  assign n42577 = n33497 & ~n64800;
  assign n42578 = ~n42030 & ~n42291;
  assign n42579 = ~pi152 & n42037;
  assign n42580 = ~n42578 & ~n42579;
  assign n42581 = ~pi172 & ~n42580;
  assign n42582 = ~pi152 & n42040;
  assign n42583 = pi152 & n42075;
  assign n42584 = pi172 & ~n42583;
  assign n42585 = ~n42582 & n42584;
  assign n42586 = n31886 & ~n42585;
  assign n42587 = n31886 & ~n42581;
  assign n42588 = ~n42585 & n42587;
  assign n42589 = ~n42581 & n42586;
  assign n42590 = n33512 & ~n64801;
  assign n42591 = ~n42577 & ~n42590;
  assign n42592 = ~n42566 & ~n42591;
  assign n42593 = ~n2814 & ~n41765;
  assign n42594 = ~n31926 & ~n42593;
  assign n42595 = ~n42074 & n42594;
  assign n42596 = n31926 & n42040;
  assign n42597 = ~n42595 & ~n42596;
  assign n42598 = ~pi174 & n42597;
  assign n42599 = ~n41762 & ~n42557;
  assign n42600 = pi174 & n42599;
  assign n42601 = ~pi180 & ~n42600;
  assign n42602 = ~n42598 & n42601;
  assign n42603 = n31926 & ~n42033;
  assign n42604 = ~n39240 & n42603;
  assign n42605 = ~n42595 & ~n42604;
  assign n42606 = ~pi174 & n42605;
  assign n42607 = ~pi51 & ~n42054;
  assign n42608 = n2814 & ~n42607;
  assign n42609 = ~n42557 & ~n42608;
  assign n42610 = pi174 & n42609;
  assign n42611 = pi180 & ~n42610;
  assign n42612 = ~n42606 & n42611;
  assign n42613 = ~n42602 & ~n42612;
  assign n42614 = ~pi174 & ~n42597;
  assign n42615 = pi174 & ~n42599;
  assign n42616 = ~pi180 & ~n42615;
  assign n42617 = ~n42614 & n42616;
  assign n42618 = ~pi174 & ~n42605;
  assign n42619 = pi174 & ~n42609;
  assign n42620 = pi180 & ~n42619;
  assign n42621 = ~n42618 & n42620;
  assign n42622 = pi193 & ~n42621;
  assign n42623 = ~n42617 & n42622;
  assign n42624 = pi193 & ~n42613;
  assign n42625 = ~pi51 & n42594;
  assign n42626 = n31926 & n42038;
  assign n42627 = ~n42625 & ~n42626;
  assign n42628 = pi180 & n42050;
  assign n42629 = ~pi174 & ~n42628;
  assign n42630 = n42627 & n42629;
  assign n42631 = pi180 & n42054;
  assign n42632 = pi174 & ~n42557;
  assign n42633 = ~n42631 & n42632;
  assign n42634 = ~pi193 & ~n42633;
  assign n42635 = ~n42630 & n42634;
  assign n42636 = ~pi299 & ~n42635;
  assign n42637 = ~n64802 & n42636;
  assign n42638 = ~n42592 & ~n42637;
  assign n42639 = pi232 & ~n42638;
  assign n42640 = n42564 & ~n42639;
  assign n42641 = ~n42555 & ~n42640;
  assign n42642 = ~n41762 & ~n41913;
  assign n42643 = ~pi174 & ~n42366;
  assign n42644 = pi145 & n41765;
  assign n42645 = ~n42643 & ~n42644;
  assign n42646 = n42642 & ~n42645;
  assign n42647 = ~n41913 & ~n42178;
  assign n42648 = pi174 & n42647;
  assign n42649 = ~n42646 & ~n42648;
  assign n42650 = ~pi193 & ~n42649;
  assign n42651 = pi145 & ~n41903;
  assign n42652 = ~pi145 & pi174;
  assign n42653 = ~n42176 & n42652;
  assign n42654 = ~n42651 & ~n42653;
  assign n42655 = ~n42643 & n42654;
  assign n42656 = pi193 & ~n41913;
  assign n42657 = ~n42655 & n42656;
  assign n42658 = n31955 & ~n42657;
  assign n42659 = ~n42650 & n42658;
  assign n42660 = n41873 & n64767;
  assign n42661 = ~n41913 & ~n42660;
  assign n42662 = ~pi145 & n42661;
  assign n42663 = ~n41894 & ~n41913;
  assign n42664 = pi145 & n42663;
  assign n42665 = ~pi174 & ~n42664;
  assign n42666 = ~n42662 & n42665;
  assign n42667 = ~pi145 & ~n41911;
  assign n42668 = ~n2814 & ~n41911;
  assign n42669 = ~n41767 & ~n42668;
  assign n42670 = ~n41845 & n42669;
  assign n42671 = ~n42667 & n42670;
  assign n42672 = n2728 & n42671;
  assign n42673 = ~n41913 & ~n42157;
  assign n42674 = pi174 & ~n42673;
  assign n42675 = pi174 & ~n42672;
  assign n42676 = ~n42673 & n42675;
  assign n42677 = ~n42672 & n42674;
  assign n42678 = pi193 & ~n64803;
  assign n42679 = ~n42666 & n42678;
  assign n42680 = ~pi145 & ~n41913;
  assign n42681 = ~n42149 & n42680;
  assign n42682 = ~pi51 & n42664;
  assign n42683 = ~pi174 & ~n42682;
  assign n42684 = ~n42681 & n42683;
  assign n42685 = pi174 & ~n42671;
  assign n42686 = ~pi193 & ~n42685;
  assign n42687 = ~n42684 & n42686;
  assign n42688 = n31935 & ~n42687;
  assign n42689 = n31935 & ~n42679;
  assign n42690 = ~n42687 & n42689;
  assign n42691 = ~n42679 & n42688;
  assign n42692 = ~n42659 & ~n64804;
  assign n42693 = n32271 & ~n42692;
  assign n42694 = ~n42641 & ~n42693;
  assign n42695 = ~pi38 & ~n42694;
  assign n42696 = ~n41808 & ~n42540;
  assign n42697 = pi152 & n42647;
  assign n42698 = ~pi152 & ~n41762;
  assign n42699 = ~pi172 & ~n42698;
  assign n42700 = ~n42697 & n42699;
  assign n42701 = ~n41913 & ~n41943;
  assign n42702 = ~pi152 & ~n42701;
  assign n42703 = ~n41913 & ~n42176;
  assign n42704 = pi152 & pi172;
  assign n42705 = ~n42703 & n42704;
  assign n42706 = ~n42702 & ~n42705;
  assign n42707 = ~pi172 & ~n42647;
  assign n42708 = pi172 & ~n42703;
  assign n42709 = pi152 & ~n42708;
  assign n42710 = ~n42707 & n42709;
  assign n42711 = ~pi172 & n41762;
  assign n42712 = ~pi152 & ~n42711;
  assign n42713 = n42701 & n42712;
  assign n42714 = ~n42710 & ~n42713;
  assign n42715 = ~n42700 & n42706;
  assign n42716 = ~pi152 & n42701;
  assign n42717 = ~n41762 & n42716;
  assign n42718 = ~pi172 & ~n42697;
  assign n42719 = ~n42717 & n42718;
  assign n42720 = pi152 & n42703;
  assign n42721 = pi172 & ~n42720;
  assign n42722 = ~n42716 & n42721;
  assign n42723 = ~pi197 & ~n42722;
  assign n42724 = ~n42719 & n42723;
  assign n42725 = ~pi197 & ~n64805;
  assign n42726 = ~pi172 & ~n42282;
  assign n42727 = ~n41914 & n42726;
  assign n42728 = pi152 & n41903;
  assign n42729 = ~n41913 & ~n42728;
  assign n42730 = pi172 & ~n42729;
  assign n42731 = pi197 & ~n42730;
  assign n42732 = pi197 & ~n42727;
  assign n42733 = ~n42730 & n42732;
  assign n42734 = ~n42727 & n42731;
  assign n42735 = pi299 & n31918;
  assign n42736 = ~n64807 & n42735;
  assign n42737 = ~n42727 & ~n42730;
  assign n42738 = pi197 & ~n42737;
  assign n42739 = ~pi197 & n64805;
  assign n42740 = ~n42738 & ~n42739;
  assign n42741 = n42735 & ~n42740;
  assign n42742 = ~n64806 & n42736;
  assign n42743 = ~pi152 & n42149;
  assign n42744 = ~n41912 & ~n42291;
  assign n42745 = ~pi172 & ~n42744;
  assign n42746 = ~n42743 & n42745;
  assign n42747 = ~pi152 & ~n42661;
  assign n42748 = pi152 & ~n42673;
  assign n42749 = pi172 & ~n42748;
  assign n42750 = ~n42747 & n42749;
  assign n42751 = ~n42746 & ~n42750;
  assign n42752 = ~n42743 & ~n42744;
  assign n42753 = ~pi172 & ~n42752;
  assign n42754 = ~pi152 & n42661;
  assign n42755 = pi152 & n42673;
  assign n42756 = pi172 & ~n42755;
  assign n42757 = ~n42754 & n42756;
  assign n42758 = ~pi197 & ~n42757;
  assign n42759 = ~n42753 & n42758;
  assign n42760 = ~pi197 & ~n42751;
  assign n42761 = ~pi152 & ~n42663;
  assign n42762 = ~n41906 & ~n41913;
  assign n42763 = pi172 & n42762;
  assign n42764 = ~pi172 & n42670;
  assign n42765 = pi152 & ~n42764;
  assign n42766 = pi172 & ~n42762;
  assign n42767 = ~pi172 & ~n42670;
  assign n42768 = ~n42766 & ~n42767;
  assign n42769 = pi152 & ~n42768;
  assign n42770 = ~n42763 & n42765;
  assign n42771 = pi197 & ~n42711;
  assign n42772 = ~n64810 & n42771;
  assign n42773 = ~n42761 & n42772;
  assign n42774 = pi299 & n31909;
  assign n42775 = ~n42773 & n42774;
  assign n42776 = ~n64809 & n42775;
  assign n42777 = ~n64808 & ~n42776;
  assign n42778 = n32271 & ~n42777;
  assign n42779 = ~n42696 & ~n42778;
  assign n42780 = ~pi38 & ~n42692;
  assign n42781 = n42777 & ~n42780;
  assign n42782 = n32271 & ~n42781;
  assign n42783 = ~pi38 & ~n42555;
  assign n42784 = ~n42640 & n42783;
  assign n42785 = ~n42696 & ~n42784;
  assign n42786 = ~n42782 & n42785;
  assign n42787 = ~n42695 & n42779;
  assign n42788 = ~n42135 & n42544;
  assign n42789 = n42136 & ~n42543;
  assign n42790 = ~n64811 & n64812;
  assign n42791 = n42140 & ~n42538;
  assign n42792 = ~n42279 & ~n42550;
  assign n42793 = ~n42791 & n42792;
  assign n42794 = ~n42790 & n42793;
  assign n42795 = n62455 & ~n42794;
  assign n42796 = ~n42553 & n42795;
  assign n42797 = ~n42290 & ~n42796;
  assign n42798 = ~pi189 & n42322;
  assign n42799 = pi189 & n42315;
  assign n42800 = ~n42798 & ~n42799;
  assign n42801 = pi178 & ~n42800;
  assign n42802 = pi189 & ~n42304;
  assign n42803 = ~pi189 & ~n42298;
  assign n42804 = ~pi178 & ~n42803;
  assign n42805 = ~pi178 & ~n42802;
  assign n42806 = ~n42803 & n42805;
  assign n42807 = ~n42802 & n42804;
  assign n42808 = ~n42801 & ~n64813;
  assign n42809 = pi181 & ~n42808;
  assign n42810 = pi189 & n42335;
  assign n42811 = ~pi189 & ~n42337;
  assign n42812 = pi178 & ~n42811;
  assign n42813 = ~n42810 & n42812;
  assign n42814 = ~pi189 & ~n42360;
  assign n42815 = pi189 & n41867;
  assign n42816 = ~pi178 & ~n42815;
  assign n42817 = ~n41762 & n42816;
  assign n42818 = ~n42814 & n42817;
  assign n42819 = ~pi181 & ~n42818;
  assign n42820 = n42360 & n42816;
  assign n42821 = n42819 & ~n42820;
  assign n42822 = ~n42813 & n42821;
  assign n42823 = n32487 & ~n42822;
  assign n42824 = ~n42809 & n42823;
  assign n42825 = ~pi153 & ~n42315;
  assign n42826 = pi153 & ~n42317;
  assign n42827 = pi157 & ~n42826;
  assign n42828 = ~n42825 & n42827;
  assign n42829 = ~pi153 & ~n42304;
  assign n42830 = pi153 & n64785;
  assign n42831 = ~pi157 & ~n42830;
  assign n42832 = ~n42829 & n42831;
  assign n42833 = pi166 & ~n42832;
  assign n42834 = ~pi153 & n42315;
  assign n42835 = pi153 & n42317;
  assign n42836 = pi157 & ~n42835;
  assign n42837 = ~n42834 & n42836;
  assign n42838 = ~pi153 & n42304;
  assign n42839 = pi153 & ~n64785;
  assign n42840 = ~pi157 & ~n42839;
  assign n42841 = ~n42838 & n42840;
  assign n42842 = ~n42837 & ~n42841;
  assign n42843 = pi166 & ~n42842;
  assign n42844 = ~n42828 & n42833;
  assign n42845 = pi157 & n42322;
  assign n42846 = ~pi157 & n42298;
  assign n42847 = pi153 & n41762;
  assign n42848 = ~pi166 & ~n42847;
  assign n42849 = ~n42846 & n42848;
  assign n42850 = ~n42845 & n42848;
  assign n42851 = ~n42846 & n42850;
  assign n42852 = ~n42845 & n42849;
  assign n42853 = ~n64814 & ~n64815;
  assign n42854 = n31761 & ~n42853;
  assign n42855 = pi166 & ~n42341;
  assign n42856 = ~pi166 & n42345;
  assign n42857 = pi153 & ~n42856;
  assign n42858 = ~n42855 & n42857;
  assign n42859 = pi166 & n42335;
  assign n42860 = ~pi166 & ~n42337;
  assign n42861 = ~pi153 & ~n42860;
  assign n42862 = ~n42859 & n42861;
  assign n42863 = ~n42858 & ~n42862;
  assign n42864 = pi157 & ~n42863;
  assign n42865 = ~pi166 & ~n42360;
  assign n42866 = pi166 & n41867;
  assign n42867 = ~pi157 & ~n42847;
  assign n42868 = ~n42866 & n42867;
  assign n42869 = ~n42865 & n42868;
  assign n42870 = ~n42864 & ~n42869;
  assign n42871 = n31784 & ~n42870;
  assign n42872 = ~pi189 & n42642;
  assign n42873 = n42317 & ~n42872;
  assign n42874 = pi178 & ~n42798;
  assign n42875 = ~n42873 & n42874;
  assign n42876 = pi189 & n64785;
  assign n42877 = ~n41762 & n42803;
  assign n42878 = ~n42876 & ~n42877;
  assign n42879 = ~pi178 & ~n42878;
  assign n42880 = pi181 & ~n42879;
  assign n42881 = ~n42875 & n42880;
  assign n42882 = pi189 & ~n42341;
  assign n42883 = ~pi189 & n42345;
  assign n42884 = pi178 & ~n42883;
  assign n42885 = ~n42882 & n42884;
  assign n42886 = n42819 & ~n42885;
  assign n42887 = n32545 & ~n42886;
  assign n42888 = ~n42881 & n42887;
  assign n42889 = ~n42871 & ~n42888;
  assign n42890 = ~n42854 & n42889;
  assign n42891 = ~n42824 & n42889;
  assign n42892 = ~n42854 & n42891;
  assign n42893 = ~n42824 & n42890;
  assign n42894 = pi232 & ~n64816;
  assign n42895 = n42530 & ~n42894;
  assign n42896 = ~pi126 & n41785;
  assign n42897 = pi126 & ~n41785;
  assign n42898 = ~n42896 & ~n42897;
  assign n42899 = ~n41781 & ~n42898;
  assign n42900 = ~pi189 & n42464;
  assign n42901 = pi189 & n64794;
  assign n42902 = ~pi182 & ~n42901;
  assign n42903 = ~pi182 & ~n42900;
  assign n42904 = ~n42901 & n42903;
  assign n42905 = ~n42900 & n42902;
  assign n42906 = ~n41762 & n64817;
  assign n42907 = pi189 & ~n42435;
  assign n42908 = ~pi189 & n42444;
  assign n42909 = pi182 & ~n42908;
  assign n42910 = ~n42907 & n42909;
  assign n42911 = ~n42906 & ~n42910;
  assign n42912 = n32545 & ~n42911;
  assign n42913 = ~pi189 & ~n42454;
  assign n42914 = pi189 & n42457;
  assign n42915 = pi182 & ~n42914;
  assign n42916 = ~n42913 & n42915;
  assign n42917 = ~n64817 & ~n42916;
  assign n42918 = n32487 & ~n42917;
  assign n42919 = pi166 & n42232;
  assign n42920 = n2933 & n32409;
  assign n42921 = ~pi166 & n42066;
  assign n42922 = ~pi153 & ~n42921;
  assign n42923 = ~n64818 & n42922;
  assign n42924 = pi166 & ~n42427;
  assign n42925 = ~pi166 & ~n42498;
  assign n42926 = pi153 & ~n42925;
  assign n42927 = ~n42924 & n42926;
  assign n42928 = pi160 & ~n42927;
  assign n42929 = pi166 & n42427;
  assign n42930 = ~pi166 & n42498;
  assign n42931 = pi153 & ~n42930;
  assign n42932 = ~n42929 & n42931;
  assign n42933 = pi166 & ~n42232;
  assign n42934 = ~pi166 & ~n42066;
  assign n42935 = ~pi153 & ~n42934;
  assign n42936 = ~n42933 & n42935;
  assign n42937 = ~n42932 & ~n42936;
  assign n42938 = pi160 & ~n42937;
  assign n42939 = pi160 & ~n42923;
  assign n42940 = ~n42927 & n42939;
  assign n42941 = ~n42923 & n42928;
  assign n42942 = pi216 & ~n64819;
  assign n42943 = pi166 & n64793;
  assign n42944 = ~pi166 & n42438;
  assign n42945 = pi51 & ~pi153;
  assign n42946 = ~n42944 & ~n42945;
  assign n42947 = ~n42943 & ~n42945;
  assign n42948 = ~n42944 & n42947;
  assign n42949 = ~pi166 & ~n42438;
  assign n42950 = pi166 & ~n64793;
  assign n42951 = ~n42949 & ~n42950;
  assign n42952 = ~n42945 & ~n42951;
  assign n42953 = ~n42943 & n42946;
  assign n42954 = ~pi216 & ~n64820;
  assign n42955 = n2960 & ~n42954;
  assign n42956 = n2960 & ~n42942;
  assign n42957 = ~n42954 & n42956;
  assign n42958 = ~n42942 & n42955;
  assign n42959 = ~pi51 & ~n41903;
  assign n42960 = ~n32363 & ~n41765;
  assign n42961 = ~pi51 & ~n42960;
  assign n42962 = ~n42847 & ~n42961;
  assign n42963 = ~n42959 & ~n42962;
  assign n42964 = ~pi160 & pi216;
  assign n42965 = n2960 & ~n42964;
  assign n42966 = n42963 & ~n42965;
  assign n42967 = pi299 & ~n42966;
  assign n42968 = ~n64821 & n42967;
  assign n42969 = ~n42918 & ~n42968;
  assign n42970 = ~n42912 & ~n42918;
  assign n42971 = ~n42968 & n42970;
  assign n42972 = ~n42912 & n42969;
  assign n42973 = pi232 & ~n64822;
  assign n42974 = n42426 & ~n42973;
  assign n42975 = n42899 & ~n42974;
  assign n42976 = ~n42895 & n42975;
  assign n42977 = ~n32363 & ~n41912;
  assign n42978 = ~pi166 & n42149;
  assign n42979 = ~n42977 & ~n42978;
  assign n42980 = ~pi153 & ~n42979;
  assign n42981 = ~pi166 & n42661;
  assign n42982 = pi166 & n42673;
  assign n42983 = pi153 & ~n42982;
  assign n42984 = ~n42981 & n42983;
  assign n42985 = ~pi157 & ~n42984;
  assign n42986 = ~pi166 & ~n42661;
  assign n42987 = pi166 & ~n42673;
  assign n42988 = pi153 & ~n42987;
  assign n42989 = ~n42986 & n42988;
  assign n42990 = ~pi153 & ~n42977;
  assign n42991 = ~n42978 & n42990;
  assign n42992 = ~n42989 & ~n42991;
  assign n42993 = ~pi157 & ~n42992;
  assign n42994 = ~n42980 & n42985;
  assign n42995 = pi166 & ~n42647;
  assign n42996 = pi51 & n32363;
  assign n42997 = ~n42995 & ~n42996;
  assign n42998 = ~pi153 & ~n42997;
  assign n42999 = ~pi166 & ~n42701;
  assign n43000 = pi153 & pi166;
  assign n43001 = ~n42703 & n43000;
  assign n43002 = pi157 & ~n43001;
  assign n43003 = ~n42999 & n43002;
  assign n43004 = ~n42998 & n43002;
  assign n43005 = ~n42999 & n43004;
  assign n43006 = ~n42998 & n43003;
  assign n43007 = n31784 & ~n64824;
  assign n43008 = ~n64823 & n43007;
  assign n43009 = ~n32501 & ~n41912;
  assign n43010 = ~pi189 & n42149;
  assign n43011 = ~n43009 & ~n43010;
  assign n43012 = ~pi178 & ~n43011;
  assign n43013 = pi189 & n42647;
  assign n43014 = pi178 & ~n42872;
  assign n43015 = ~pi189 & n42701;
  assign n43016 = pi178 & ~n43015;
  assign n43017 = ~n43014 & ~n43016;
  assign n43018 = ~n43013 & ~n43017;
  assign n43019 = ~pi181 & ~n43018;
  assign n43020 = ~n43012 & n43019;
  assign n43021 = ~n41894 & n42872;
  assign n43022 = pi189 & n42670;
  assign n43023 = ~pi178 & ~n43022;
  assign n43024 = ~n43021 & n43023;
  assign n43025 = pi189 & n41914;
  assign n43026 = n43014 & ~n43025;
  assign n43027 = pi181 & ~n43026;
  assign n43028 = ~n43024 & n43027;
  assign n43029 = n32487 & ~n43028;
  assign n43030 = ~n43020 & n43029;
  assign n43031 = ~pi189 & n42661;
  assign n43032 = pi189 & n42673;
  assign n43033 = ~pi178 & ~n43032;
  assign n43034 = ~n43031 & n43033;
  assign n43035 = pi189 & n42703;
  assign n43036 = n43016 & ~n43035;
  assign n43037 = ~pi181 & ~n43036;
  assign n43038 = ~n43034 & n43037;
  assign n43039 = ~pi189 & ~n41894;
  assign n43040 = pi189 & ~n41906;
  assign n43041 = ~pi178 & ~n43040;
  assign n43042 = ~n43039 & n43041;
  assign n43043 = pi178 & n32498;
  assign n43044 = n41902 & n43043;
  assign n43045 = pi181 & ~n43044;
  assign n43046 = ~n41913 & n43045;
  assign n43047 = ~n43042 & n43046;
  assign n43048 = n32545 & ~n43047;
  assign n43049 = ~n43038 & n43048;
  assign n43050 = ~pi166 & ~n42663;
  assign n43051 = ~n42762 & n43000;
  assign n43052 = pi166 & ~n42670;
  assign n43053 = ~n42996 & ~n43052;
  assign n43054 = ~pi153 & ~n43053;
  assign n43055 = ~pi157 & ~n43054;
  assign n43056 = ~pi157 & ~n43051;
  assign n43057 = ~n43054 & n43056;
  assign n43058 = ~n43051 & n43055;
  assign n43059 = ~n43050 & n64825;
  assign n43060 = ~pi153 & ~n42963;
  assign n43061 = ~n41914 & n43060;
  assign n43062 = pi166 & n41903;
  assign n43063 = n32409 & n41902;
  assign n43064 = ~n41913 & ~n64826;
  assign n43065 = pi153 & ~n43064;
  assign n43066 = pi157 & ~n43065;
  assign n43067 = pi157 & ~n43061;
  assign n43068 = ~n43065 & n43067;
  assign n43069 = ~n43061 & n43066;
  assign n43070 = n31761 & ~n64827;
  assign n43071 = ~n43059 & n43070;
  assign n43072 = ~n43049 & ~n43071;
  assign n43073 = ~n43030 & n43072;
  assign n43074 = ~n43008 & n43072;
  assign n43075 = ~n43030 & n43074;
  assign n43076 = ~n43008 & n43073;
  assign n43077 = pi232 & ~n64828;
  assign n43078 = n42555 & ~n43077;
  assign n43079 = ~pi166 & ~n42051;
  assign n43080 = pi166 & n42054;
  assign n43081 = pi160 & ~n42847;
  assign n43082 = ~n43080 & n43081;
  assign n43083 = ~pi166 & n42051;
  assign n43084 = pi166 & ~n42054;
  assign n43085 = ~n43083 & ~n43084;
  assign n43086 = n43081 & ~n43085;
  assign n43087 = ~n43079 & n43082;
  assign n43088 = ~pi166 & ~n42040;
  assign n43089 = pi166 & ~n42075;
  assign n43090 = pi153 & ~n43089;
  assign n43091 = ~n43088 & n43090;
  assign n43092 = ~pi166 & n42037;
  assign n43093 = ~n32363 & ~n42030;
  assign n43094 = ~pi153 & ~n43093;
  assign n43095 = ~n43092 & n43094;
  assign n43096 = ~pi160 & ~n43095;
  assign n43097 = ~n43092 & ~n43093;
  assign n43098 = ~pi153 & ~n43097;
  assign n43099 = ~pi166 & n42040;
  assign n43100 = pi166 & n42075;
  assign n43101 = pi153 & ~n43100;
  assign n43102 = ~n43099 & n43101;
  assign n43103 = ~n43098 & ~n43102;
  assign n43104 = ~pi160 & ~n43103;
  assign n43105 = ~n43091 & n43096;
  assign n43106 = n31886 & ~n64830;
  assign n43107 = n31886 & ~n64829;
  assign n43108 = ~n64830 & n43107;
  assign n43109 = ~n64829 & n43106;
  assign n43110 = ~n31886 & ~n42962;
  assign n43111 = pi299 & ~n43110;
  assign n43112 = ~n64831 & n43111;
  assign n43113 = ~pi189 & ~n42597;
  assign n43114 = pi189 & ~n42599;
  assign n43115 = ~pi182 & ~n43114;
  assign n43116 = ~n43113 & n43115;
  assign n43117 = ~pi189 & ~n42605;
  assign n43118 = pi189 & ~n42609;
  assign n43119 = pi182 & ~n43118;
  assign n43120 = ~n43117 & n43119;
  assign n43121 = ~n43116 & ~n43120;
  assign n43122 = n32545 & ~n43121;
  assign n43123 = pi182 & n42054;
  assign n43124 = pi189 & ~n42557;
  assign n43125 = ~n43123 & n43124;
  assign n43126 = pi182 & n42050;
  assign n43127 = ~pi189 & ~n43126;
  assign n43128 = n42627 & n43127;
  assign n43129 = ~n43125 & ~n43128;
  assign n43130 = n32487 & ~n43129;
  assign n43131 = ~n43122 & ~n43130;
  assign n43132 = ~n43112 & n43131;
  assign n43133 = pi232 & ~n43132;
  assign n43134 = n42564 & ~n43133;
  assign n43135 = ~n42899 & ~n43134;
  assign n43136 = ~n43078 & n43135;
  assign n43137 = n2766 & ~n43136;
  assign n43138 = ~n42976 & n43137;
  assign n43139 = pi299 & ~n42963;
  assign n43140 = ~pi189 & n41903;
  assign n43141 = n32501 & n41902;
  assign n43142 = pi175 & n41762;
  assign n43143 = ~pi299 & ~n43142;
  assign n43144 = ~n64832 & n43143;
  assign n43145 = pi232 & ~n43144;
  assign n43146 = ~n43139 & n43145;
  assign n43147 = ~n2766 & n43146;
  assign n43148 = ~n2766 & n41766;
  assign n43149 = ~n42899 & n43148;
  assign n43150 = n6797 & ~n43149;
  assign n43151 = n41766 & ~n42899;
  assign n43152 = ~n43146 & ~n43151;
  assign n43153 = ~n2766 & ~n43152;
  assign n43154 = n6797 & ~n43153;
  assign n43155 = ~n43147 & n43150;
  assign n43156 = ~n43138 & n64833;
  assign n43157 = ~pi150 & pi299;
  assign n43158 = ~pi185 & ~pi299;
  assign n43159 = ~n43157 & ~n43158;
  assign n43160 = n2815 & n43159;
  assign n43161 = pi87 & ~n43160;
  assign n43162 = n42139 & n43152;
  assign n43163 = n42139 & ~n43146;
  assign n43164 = ~n43161 & ~n43163;
  assign n43165 = n41788 & ~n42899;
  assign n43166 = ~n43164 & ~n43165;
  assign n43167 = ~n43161 & ~n43162;
  assign n43168 = n62455 & ~n64834;
  assign n43169 = ~n43156 & n43168;
  assign n43170 = pi232 & ~n42959;
  assign n43171 = n42899 & ~n43170;
  assign n43172 = ~pi232 & ~n41766;
  assign n43173 = ~n42962 & ~n43172;
  assign n43174 = ~n43171 & n43173;
  assign n43175 = ~pi87 & ~n43174;
  assign n43176 = pi87 & ~n33150;
  assign n43177 = ~n62455 & ~n43176;
  assign n43178 = ~n43175 & n43177;
  assign n43179 = ~n43156 & ~n64834;
  assign n43180 = n62455 & ~n43179;
  assign n43181 = ~pi232 & ~n43151;
  assign n43182 = n42899 & n42959;
  assign n43183 = ~pi87 & ~n42962;
  assign n43184 = ~n43182 & n43183;
  assign n43185 = pi232 & ~n43182;
  assign n43186 = ~n43151 & ~n43185;
  assign n43187 = n43183 & ~n43186;
  assign n43188 = ~n43181 & n43184;
  assign n43189 = pi87 & n33150;
  assign n43190 = ~n62455 & ~n43189;
  assign n43191 = ~n64835 & n43190;
  assign n43192 = ~n43180 & ~n43191;
  assign n43193 = ~n43169 & ~n43178;
  assign n43194 = n3318 & ~n34974;
  assign n43195 = n34975 & ~n43194;
  assign n43196 = n64196 & ~n43195;
  assign n43197 = n39218 & ~n43195;
  assign n43198 = n39166 & n43196;
  assign n43199 = ~pi94 & n6803;
  assign n43200 = n2698 & n43199;
  assign n43201 = n2688 & n5549;
  assign n43202 = n39878 & n64838;
  assign n43203 = n2852 & n64196;
  assign n43204 = n62651 & n43203;
  assign n43205 = n43202 & n43204;
  assign n43206 = n34974 & n43205;
  assign n43207 = ~pi110 & ~n43202;
  assign n43208 = ~pi47 & ~n34974;
  assign n43209 = n43203 & n43208;
  assign n43210 = ~n43207 & n43209;
  assign n43211 = n39182 & n43210;
  assign n43212 = ~n43206 & ~n43211;
  assign n43213 = ~n3318 & ~n6899;
  assign n43214 = ~pi47 & n43203;
  assign n43215 = ~n43207 & n43214;
  assign n43216 = n39182 & n43215;
  assign n43217 = ~n34974 & ~n43216;
  assign n43218 = n34974 & ~n43205;
  assign n43219 = n43213 & ~n43218;
  assign n43220 = ~n43217 & n43219;
  assign n43221 = n2843 & ~n43216;
  assign n43222 = ~n2843 & ~n43205;
  assign n43223 = ~n2816 & ~n6899;
  assign n43224 = ~n43222 & n43223;
  assign n43225 = ~n43221 & n43224;
  assign n43226 = n2816 & ~n6899;
  assign n43227 = n43216 & n43226;
  assign n43228 = ~n43225 & ~n43227;
  assign n43229 = ~n3318 & ~n43228;
  assign n43230 = ~n43212 & n43213;
  assign n43231 = ~n64837 & ~n64839;
  assign po262 = n64705 & ~n43231;
  assign n43233 = pi51 & ~pi151;
  assign n43234 = ~n33016 & ~n41762;
  assign n43235 = ~n43233 & ~n43234;
  assign n43236 = n41767 & n43235;
  assign n43237 = pi232 & n43236;
  assign n43238 = ~pi132 & n42896;
  assign n43239 = pi132 & ~n42896;
  assign n43240 = ~n43238 & ~n43239;
  assign n43241 = ~n41780 & ~n43240;
  assign n43242 = n41766 & ~n43241;
  assign n43243 = ~n43237 & ~n43242;
  assign n43244 = ~pi87 & ~n43243;
  assign n43245 = pi164 & n42287;
  assign n43246 = ~n62455 & ~n43245;
  assign n43247 = ~n43244 & n43246;
  assign n43248 = pi299 & ~n43236;
  assign n43249 = pi190 & n41903;
  assign n43250 = pi173 & n41762;
  assign n43251 = ~pi299 & ~n43250;
  assign n43252 = ~n43249 & n43251;
  assign n43253 = pi232 & ~n43252;
  assign n43254 = pi232 & ~n43248;
  assign n43255 = ~n43252 & n43254;
  assign n43256 = ~n43248 & n43253;
  assign n43257 = ~n2766 & n64840;
  assign n43258 = n6797 & ~n43257;
  assign n43259 = pi183 & n42434;
  assign n43260 = ~pi183 & n64794;
  assign n43261 = ~n41762 & ~n43260;
  assign n43262 = ~n43259 & n43261;
  assign n43263 = pi183 & n42435;
  assign n43264 = ~pi183 & ~n41762;
  assign n43265 = ~n64794 & n43264;
  assign n43266 = pi173 & ~n43265;
  assign n43267 = ~n43263 & n43266;
  assign n43268 = pi173 & ~n43262;
  assign n43269 = ~pi190 & ~pi299;
  assign n43270 = ~pi183 & ~n3076;
  assign n43271 = ~pi173 & ~n43270;
  assign n43272 = n42457 & n43271;
  assign n43273 = n43269 & ~n43272;
  assign n43274 = ~n64841 & n43273;
  assign n43275 = pi190 & ~pi299;
  assign n43276 = pi183 & ~n42454;
  assign n43277 = ~pi183 & ~n42449;
  assign n43278 = ~pi173 & ~n43277;
  assign n43279 = ~n43276 & n43278;
  assign n43280 = ~pi183 & n42463;
  assign n43281 = ~pi183 & ~n42439;
  assign n43282 = pi173 & ~n42444;
  assign n43283 = ~n43281 & n43282;
  assign n43284 = ~n43280 & ~n43283;
  assign n43285 = ~n43279 & n43284;
  assign n43286 = n43275 & ~n43285;
  assign n43287 = ~pi168 & ~n42427;
  assign n43288 = pi168 & ~n42498;
  assign n43289 = pi151 & ~n43288;
  assign n43290 = ~n43287 & n43289;
  assign n43291 = pi168 & n42066;
  assign n43292 = ~pi168 & n42232;
  assign n43293 = ~pi151 & ~n43292;
  assign n43294 = ~pi151 & ~n43291;
  assign n43295 = ~n43292 & n43294;
  assign n43296 = ~n43291 & n43293;
  assign n43297 = pi149 & ~n64842;
  assign n43298 = pi149 & ~n43290;
  assign n43299 = ~n64842 & n43298;
  assign n43300 = ~n43290 & n43297;
  assign n43301 = pi216 & ~n64843;
  assign n43302 = ~pi168 & n64793;
  assign n43303 = pi168 & n42438;
  assign n43304 = ~n43233 & ~n43303;
  assign n43305 = ~n43233 & ~n43302;
  assign n43306 = ~n43303 & n43305;
  assign n43307 = pi168 & ~n42438;
  assign n43308 = ~pi168 & ~n64793;
  assign n43309 = ~n43307 & ~n43308;
  assign n43310 = ~n43233 & ~n43309;
  assign n43311 = ~n43302 & n43304;
  assign n43312 = ~pi216 & ~n64844;
  assign n43313 = n2960 & ~n43312;
  assign n43314 = n2960 & ~n43301;
  assign n43315 = ~n43312 & n43314;
  assign n43316 = ~n43301 & n43313;
  assign n43317 = ~pi149 & pi216;
  assign n43318 = n2960 & ~n43317;
  assign n43319 = n43236 & ~n43318;
  assign n43320 = pi299 & ~n43319;
  assign n43321 = ~n64845 & n43320;
  assign n43322 = ~n43286 & ~n43321;
  assign n43323 = ~n43274 & ~n43286;
  assign n43324 = ~n43321 & n43323;
  assign n43325 = ~n43274 & n43322;
  assign n43326 = pi232 & ~n64846;
  assign n43327 = n42426 & ~n43326;
  assign n43328 = ~n2814 & n41888;
  assign n43329 = pi182 & n41830;
  assign n43330 = n41852 & ~n43329;
  assign n43331 = pi51 & ~pi173;
  assign n43332 = n2814 & ~n43331;
  assign n43333 = ~n43330 & n43332;
  assign n43334 = n43275 & ~n43333;
  assign n43335 = pi173 & n41868;
  assign n43336 = ~pi173 & ~n41875;
  assign n43337 = pi182 & n2814;
  assign n43338 = ~n43336 & n43337;
  assign n43339 = ~n43335 & n43338;
  assign n43340 = pi173 & n41897;
  assign n43341 = ~pi173 & ~n41888;
  assign n43342 = ~pi182 & ~n43341;
  assign n43343 = ~n43340 & n43342;
  assign n43344 = n43269 & ~n43343;
  assign n43345 = ~n43339 & n43344;
  assign n43346 = ~n43334 & ~n43345;
  assign n43347 = ~n43328 & ~n43346;
  assign n43348 = pi151 & n41868;
  assign n43349 = ~pi151 & ~n41875;
  assign n43350 = ~pi168 & ~n43349;
  assign n43351 = ~pi168 & ~n43348;
  assign n43352 = ~n43349 & n43351;
  assign n43353 = ~n43348 & n43350;
  assign n43354 = pi168 & ~n43233;
  assign n43355 = ~n41853 & n43354;
  assign n43356 = n2814 & ~n43355;
  assign n43357 = ~n64847 & n43356;
  assign n43358 = ~n2814 & ~n41888;
  assign n43359 = pi160 & ~n43358;
  assign n43360 = ~pi151 & n41875;
  assign n43361 = pi151 & ~n41868;
  assign n43362 = ~pi168 & ~n43361;
  assign n43363 = ~n43360 & n43362;
  assign n43364 = ~n41853 & ~n43233;
  assign n43365 = pi168 & ~n43364;
  assign n43366 = n2814 & ~n43365;
  assign n43367 = ~n43363 & n43366;
  assign n43368 = ~n43328 & ~n43367;
  assign n43369 = pi160 & ~n43368;
  assign n43370 = ~n43357 & n43359;
  assign n43371 = n41897 & ~n43328;
  assign n43372 = ~pi168 & ~n43371;
  assign n43373 = pi168 & ~n64787;
  assign n43374 = ~n43358 & n43373;
  assign n43375 = pi151 & ~n43374;
  assign n43376 = ~n43372 & n43375;
  assign n43377 = ~n33016 & n41888;
  assign n43378 = pi168 & n41917;
  assign n43379 = ~pi151 & ~n43378;
  assign n43380 = ~n43377 & n43379;
  assign n43381 = ~pi160 & ~n43380;
  assign n43382 = ~n43376 & n43381;
  assign n43383 = pi299 & ~n43382;
  assign n43384 = ~n64848 & n43383;
  assign n43385 = ~n43347 & ~n43384;
  assign n43386 = pi232 & ~n43385;
  assign n43387 = ~pi232 & ~n41888;
  assign n43388 = ~pi39 & ~n43387;
  assign n43389 = pi182 & ~n43358;
  assign n43390 = ~n41876 & n43389;
  assign n43391 = ~pi182 & n41888;
  assign n43392 = ~pi173 & ~n43391;
  assign n43393 = ~n43390 & n43392;
  assign n43394 = ~n41869 & ~n43328;
  assign n43395 = pi182 & ~n43394;
  assign n43396 = ~pi182 & ~n43371;
  assign n43397 = pi173 & ~n43396;
  assign n43398 = ~n43395 & n43397;
  assign n43399 = ~n43393 & ~n43398;
  assign n43400 = n43269 & ~n43399;
  assign n43401 = ~n43328 & n43334;
  assign n43402 = pi232 & ~n43401;
  assign n43403 = ~n43400 & n43402;
  assign n43404 = ~n43384 & n43402;
  assign n43405 = ~n43400 & n43404;
  assign n43406 = ~n43384 & n43403;
  assign n43407 = ~pi232 & n41888;
  assign n43408 = ~n64849 & ~n43407;
  assign n43409 = ~pi39 & ~n43408;
  assign n43410 = ~n43386 & n43388;
  assign n43411 = ~n43327 & ~n64850;
  assign n43412 = n2766 & ~n43411;
  assign n43413 = n43258 & ~n43412;
  assign n43414 = n42139 & ~n64840;
  assign n43415 = pi87 & ~n33365;
  assign n43416 = n43241 & ~n43415;
  assign n43417 = ~n43414 & n43416;
  assign n43418 = ~n43413 & n43417;
  assign n43419 = ~n41766 & n43248;
  assign n43420 = ~n64234 & ~n43419;
  assign n43421 = ~n42427 & ~n43233;
  assign n43422 = ~n42038 & ~n43421;
  assign n43423 = pi168 & ~n43422;
  assign n43424 = ~n42054 & ~n43235;
  assign n43425 = ~pi168 & ~n43424;
  assign n43426 = pi149 & ~n43425;
  assign n43427 = ~pi168 & ~n43235;
  assign n43428 = ~n42054 & n43427;
  assign n43429 = pi168 & ~n42038;
  assign n43430 = ~n43421 & n43429;
  assign n43431 = ~n43428 & ~n43430;
  assign n43432 = pi149 & ~n43431;
  assign n43433 = ~n43423 & n43426;
  assign n43434 = pi168 & ~n42040;
  assign n43435 = ~pi168 & ~n42075;
  assign n43436 = pi151 & ~n43435;
  assign n43437 = ~n43434 & n43436;
  assign n43438 = pi168 & n42037;
  assign n43439 = ~n33016 & ~n42030;
  assign n43440 = ~pi151 & ~n43439;
  assign n43441 = ~n43438 & n43440;
  assign n43442 = ~pi149 & ~n43441;
  assign n43443 = ~n43438 & ~n43439;
  assign n43444 = ~pi151 & ~n43443;
  assign n43445 = pi168 & n42040;
  assign n43446 = ~pi168 & n42075;
  assign n43447 = pi151 & ~n43446;
  assign n43448 = ~n43445 & n43447;
  assign n43449 = ~n43444 & ~n43448;
  assign n43450 = ~pi149 & ~n43449;
  assign n43451 = ~n43437 & n43442;
  assign n43452 = n31886 & ~n64852;
  assign n43453 = n31886 & ~n64851;
  assign n43454 = ~n64852 & n43453;
  assign n43455 = ~n64851 & n43452;
  assign n43456 = ~n43420 & ~n64853;
  assign n43457 = ~pi183 & ~n42597;
  assign n43458 = pi183 & ~n42605;
  assign n43459 = pi173 & ~n43458;
  assign n43460 = ~n43457 & n43459;
  assign n43461 = pi183 & n42050;
  assign n43462 = ~pi173 & ~n43461;
  assign n43463 = n42627 & n43462;
  assign n43464 = ~n43460 & ~n43463;
  assign n43465 = n43275 & ~n43464;
  assign n43466 = pi183 & n42054;
  assign n43467 = ~n43250 & n43269;
  assign n43468 = ~n42557 & n43467;
  assign n43469 = ~n43466 & n43468;
  assign n43470 = ~n43465 & ~n43469;
  assign n43471 = ~n43456 & ~n43469;
  assign n43472 = ~n43465 & n43471;
  assign n43473 = ~n43456 & n43470;
  assign n43474 = pi232 & ~n64854;
  assign n43475 = ~n42563 & ~n43474;
  assign n43476 = pi39 & ~n43475;
  assign n43477 = pi151 & n42176;
  assign n43478 = ~pi151 & ~n41911;
  assign n43479 = ~pi168 & ~n43478;
  assign n43480 = ~n43477 & n43479;
  assign n43481 = ~pi151 & n41762;
  assign n43482 = pi168 & ~n43481;
  assign n43483 = ~n41943 & n43482;
  assign n43484 = ~n43480 & ~n43483;
  assign n43485 = ~pi160 & ~n42668;
  assign n43486 = ~n43484 & n43485;
  assign n43487 = ~pi151 & ~n43236;
  assign n43488 = ~n42669 & n43487;
  assign n43489 = ~pi168 & n41903;
  assign n43490 = ~n42668 & ~n43489;
  assign n43491 = pi151 & ~n43490;
  assign n43492 = pi160 & ~n43491;
  assign n43493 = pi160 & ~n43488;
  assign n43494 = ~n43491 & n43493;
  assign n43495 = ~n43488 & n43492;
  assign n43496 = pi299 & ~n64855;
  assign n43497 = ~n43486 & n43496;
  assign n43498 = ~pi182 & n41943;
  assign n43499 = ~n42668 & ~n43331;
  assign n43500 = ~n43498 & n43499;
  assign n43501 = n43275 & ~n43500;
  assign n43502 = pi182 & n42669;
  assign n43503 = ~n41911 & n43467;
  assign n43504 = ~n43502 & n43503;
  assign n43505 = pi232 & ~n43504;
  assign n43506 = ~n43501 & n43505;
  assign n43507 = ~n43497 & n43506;
  assign n43508 = ~pi232 & n41911;
  assign n43509 = ~pi39 & ~n43508;
  assign n43510 = ~n43507 & n43509;
  assign n43511 = n2766 & ~n43510;
  assign n43512 = ~n43476 & n43511;
  assign n43513 = n6797 & ~n43148;
  assign n43514 = ~n43148 & n43258;
  assign n43515 = ~n43257 & n43513;
  assign n43516 = ~n43512 & n64856;
  assign n43517 = n42140 & ~n64840;
  assign n43518 = ~n43241 & ~n43415;
  assign n43519 = ~n43517 & n43518;
  assign n43520 = ~n43516 & n43519;
  assign n43521 = n62455 & ~n43520;
  assign n43522 = ~n43418 & n43521;
  assign n43523 = ~n43247 & ~n43522;
  assign n43524 = n2587 & n2613;
  assign n43525 = ~pi102 & ~pi104;
  assign n43526 = ~pi111 & n43525;
  assign n43527 = ~pi45 & pi49;
  assign n43528 = n43526 & n43527;
  assign n43529 = n43524 & n43528;
  assign n43530 = n6813 & n43528;
  assign n43531 = n43524 & n43530;
  assign n43532 = n6813 & n43529;
  assign n43533 = n39865 & n64857;
  assign n43534 = n38910 & n43533;
  assign n43535 = ~n33872 & ~n43534;
  assign n43536 = n62356 & n6829;
  assign n43537 = n43533 & n43536;
  assign n43538 = n62378 & n38245;
  assign n43539 = n43537 & n43538;
  assign n43540 = n34974 & n41719;
  assign n43541 = ~n43539 & ~n43540;
  assign n43542 = n40591 & ~n43541;
  assign n43543 = ~n43535 & n43542;
  assign n43544 = ~n38261 & ~n43539;
  assign n43545 = pi252 & n40591;
  assign n43546 = ~n43535 & n43545;
  assign n43547 = n2929 & n43539;
  assign n43548 = pi1093 & ~n43547;
  assign n43549 = n2883 & ~n43548;
  assign n43550 = ~pi252 & n43539;
  assign n43551 = ~n43549 & ~n43550;
  assign n43552 = ~n43546 & n43551;
  assign n43553 = ~n43546 & ~n43549;
  assign n43554 = n38261 & ~n43553;
  assign n43555 = ~n43539 & ~n43554;
  assign n43556 = ~n43544 & ~n43552;
  assign n43557 = n34974 & n64858;
  assign n43558 = ~n34974 & ~n43539;
  assign n43559 = n64705 & ~n43558;
  assign n43560 = ~n43557 & n43559;
  assign n43561 = n64705 & n43543;
  assign n43562 = n64084 & n39923;
  assign n43563 = ~n3470 & ~n43562;
  assign n43564 = pi129 & n7356;
  assign n43565 = pi38 & ~n43564;
  assign n43566 = ~n6801 & ~n33957;
  assign n43567 = n33874 & ~n33906;
  assign n43568 = n2611 & ~n43567;
  assign n43569 = n33918 & ~n43568;
  assign n43570 = n30645 & ~n43569;
  assign n43571 = n30641 & ~n43570;
  assign n43572 = n30639 & ~n43571;
  assign n43573 = ~n30637 & ~n43572;
  assign n43574 = ~pi86 & ~n43573;
  assign n43575 = n30715 & ~n43574;
  assign n43576 = pi250 & ~n2816;
  assign n43577 = pi252 & n34974;
  assign n43578 = pi250 & n43577;
  assign n43579 = n39927 & n43576;
  assign n43580 = ~pi127 & ~n64860;
  assign n43581 = po740 & n64860;
  assign n43582 = ~n43580 & ~n43581;
  assign n43583 = n33872 & n43582;
  assign n43584 = ~pi97 & ~n43583;
  assign n43585 = ~n43575 & n43584;
  assign n43586 = ~n30937 & ~n43585;
  assign n43587 = ~pi108 & ~n43586;
  assign n43588 = n33870 & ~n43587;
  assign n43589 = n30750 & ~n43588;
  assign n43590 = ~n30748 & ~n43589;
  assign n43591 = n2866 & ~n43590;
  assign n43592 = ~pi97 & ~n43575;
  assign n43593 = ~n30937 & ~n43592;
  assign n43594 = ~pi108 & ~n43593;
  assign n43595 = n33870 & ~n43594;
  assign n43596 = n30750 & ~n43595;
  assign n43597 = ~n30748 & ~n43596;
  assign n43598 = n2866 & ~n43597;
  assign n43599 = n64688 & ~n43598;
  assign n43600 = po740 & n43599;
  assign n43601 = n33873 & ~n43575;
  assign n43602 = ~n30937 & ~n43601;
  assign n43603 = ~pi108 & ~n43602;
  assign n43604 = n33870 & ~n43603;
  assign n43605 = n30750 & ~n43604;
  assign n43606 = ~n30748 & ~n43605;
  assign n43607 = n2866 & ~n43606;
  assign n43608 = n64688 & ~n43607;
  assign n43609 = ~po740 & n43608;
  assign n43610 = n64860 & ~n43609;
  assign n43611 = n64860 & ~n43600;
  assign n43612 = ~n43609 & n43611;
  assign n43613 = ~n43600 & n43610;
  assign n43614 = ~pi127 & n43599;
  assign n43615 = pi127 & n43608;
  assign n43616 = ~n64860 & ~n43615;
  assign n43617 = ~n64860 & ~n43614;
  assign n43618 = ~n43615 & n43617;
  assign n43619 = ~n43614 & n43616;
  assign n43620 = ~n64861 & ~n64862;
  assign n43621 = n64688 & ~n43591;
  assign n43622 = n40180 & ~n64863;
  assign n43623 = n40179 & ~n43622;
  assign n43624 = n2719 & ~n43623;
  assign n43625 = n40177 & ~n43624;
  assign n43626 = ~pi70 & ~n43625;
  assign n43627 = ~n30620 & ~n43626;
  assign n43628 = ~pi51 & ~n43627;
  assign n43629 = n2733 & ~n43628;
  assign n43630 = n33868 & ~n43629;
  assign n43631 = ~n30618 & ~n43630;
  assign n43632 = n2750 & ~n43631;
  assign n43633 = n43566 & ~n43632;
  assign n43634 = ~pi95 & ~n43633;
  assign n43635 = ~pi39 & pi129;
  assign n43636 = pi129 & n33963;
  assign n43637 = ~n33962 & n43635;
  assign n43638 = ~n43634 & n64864;
  assign n43639 = pi39 & n39923;
  assign n43640 = ~pi38 & ~n43639;
  assign n43641 = ~n43638 & n43640;
  assign n43642 = ~n43565 & ~n43641;
  assign n43643 = n6791 & ~n43642;
  assign n43644 = ~n62373 & ~n30571;
  assign n43645 = n39923 & ~n43644;
  assign n43646 = ~n6791 & ~n43645;
  assign n43647 = ~pi75 & ~n43646;
  assign n43648 = ~n43643 & n43647;
  assign n43649 = pi129 & n30599;
  assign n43650 = pi75 & n43649;
  assign n43651 = ~pi92 & ~n43650;
  assign n43652 = ~n43648 & n43651;
  assign n43653 = pi92 & ~pi129;
  assign n43654 = n37887 & ~n43653;
  assign n43655 = ~n43652 & n43654;
  assign n43656 = pi54 & n64081;
  assign n43657 = n39923 & n43656;
  assign n43658 = ~pi74 & ~n43657;
  assign n43659 = ~n43655 & n43658;
  assign n43660 = n34066 & n43649;
  assign n43661 = pi74 & ~n43660;
  assign n43662 = ~pi55 & ~n43661;
  assign n43663 = ~n43659 & n43662;
  assign n43664 = pi55 & n6794;
  assign n43665 = n43649 & n43664;
  assign n43666 = ~n43663 & ~n43665;
  assign n43667 = ~pi56 & ~n43666;
  assign n43668 = pi56 & ~pi62;
  assign n43669 = ~pi56 & pi62;
  assign n43670 = ~n43668 & ~n43669;
  assign n43671 = ~n43667 & n43670;
  assign n43672 = ~n43563 & ~n43671;
  assign n43673 = n3472 & ~n43672;
  assign n43674 = n3470 & n43562;
  assign n43675 = n64085 & n39923;
  assign n43676 = ~n3472 & ~n64865;
  assign n43677 = ~n30570 & ~n43676;
  assign po284 = ~n43673 & n43677;
  assign n43679 = n2751 & n64705;
  assign n43680 = n62768 & n43679;
  assign n43681 = n64196 & n64705;
  assign n43682 = n62347 & n43524;
  assign n43683 = n2588 & n43682;
  assign n43684 = ~pi69 & n43683;
  assign n43685 = n6806 & n43684;
  assign n43686 = ~pi82 & ~pi109;
  assign n43687 = pi111 & n43686;
  assign n43688 = n62651 & n43687;
  assign n43689 = n62352 & n43688;
  assign n43690 = n43685 & n43689;
  assign n43691 = n30654 & n43690;
  assign n43692 = pi314 & n43691;
  assign n43693 = n34976 & n39166;
  assign n43694 = ~n43692 & ~n43693;
  assign po268 = n64866 & ~n43694;
  assign n43696 = ~pi70 & n41231;
  assign n43697 = ~n30620 & ~n33939;
  assign n43698 = ~n43696 & n43697;
  assign n43699 = ~pi51 & ~n43698;
  assign n43700 = n2733 & ~n43699;
  assign n43701 = n33868 & ~n43700;
  assign n43702 = ~n30618 & ~n43701;
  assign n43703 = n2750 & ~n43702;
  assign n43704 = n43566 & ~n43703;
  assign n43705 = ~pi95 & ~n43704;
  assign n43706 = ~n33962 & ~n43705;
  assign n43707 = ~pi39 & ~n43706;
  assign n43708 = ~n40219 & ~n43707;
  assign n43709 = ~pi38 & ~n43708;
  assign n43710 = n33858 & ~n43709;
  assign n43711 = n30856 & ~n30871;
  assign n43712 = n34137 & n64650;
  assign n43713 = ~pi87 & ~n64867;
  assign n43714 = ~n43710 & n43713;
  assign n43715 = n34034 & ~n43714;
  assign n43716 = ~pi250 & n43577;
  assign n43717 = n34974 & n39170;
  assign n43718 = po740 & n64868;
  assign n43719 = ~pi129 & ~n64868;
  assign n43720 = n40026 & ~n43719;
  assign n43721 = n40026 & ~n43718;
  assign n43722 = ~n43719 & n43721;
  assign n43723 = ~n43718 & n43720;
  assign n43724 = n62380 & n64869;
  assign n43725 = n2579 & ~n43724;
  assign n43726 = ~n43715 & n43725;
  assign n43727 = ~n30604 & ~n30895;
  assign n43728 = ~n43726 & n43727;
  assign n43729 = n34040 & ~n43728;
  assign n43730 = n40175 & ~n43729;
  assign n43731 = ~pi56 & ~n43730;
  assign n43732 = ~n34043 & ~n43731;
  assign n43733 = ~pi62 & ~n43732;
  assign n43734 = ~n34048 & ~n43733;
  assign n43735 = n3472 & ~n43734;
  assign po286 = n30591 & ~n43735;
  assign n43737 = ~pi51 & ~n42562;
  assign n43738 = ~pi232 & ~n43737;
  assign n43739 = n27583 & ~n43738;
  assign n43740 = ~pi51 & ~n42038;
  assign n43741 = ~n42049 & n43740;
  assign n43742 = pi169 & ~n43741;
  assign n43743 = pi162 & n31886;
  assign n43744 = ~pi169 & ~n42607;
  assign n43745 = n43743 & ~n43744;
  assign n43746 = ~n43742 & n43745;
  assign n43747 = ~n35131 & ~n42063;
  assign n43748 = ~n62380 & n35131;
  assign n43749 = ~pi162 & n31886;
  assign n43750 = ~n43748 & n43749;
  assign n43751 = ~n43747 & n43749;
  assign n43752 = ~n43748 & n43751;
  assign n43753 = ~n43747 & n43750;
  assign n43754 = ~n31886 & n41902;
  assign n43755 = ~n35131 & n43754;
  assign n43756 = pi299 & ~n43755;
  assign n43757 = ~n64870 & n43756;
  assign n43758 = ~n43746 & n43757;
  assign n43759 = ~pi51 & n42627;
  assign n43760 = pi140 & n42049;
  assign n43761 = n43759 & ~n43760;
  assign n43762 = n33355 & ~n43761;
  assign n43763 = ~pi51 & ~n42557;
  assign n43764 = pi140 & n42608;
  assign n43765 = n43763 & ~n43764;
  assign n43766 = n35175 & ~n43765;
  assign n43767 = ~n43762 & ~n43766;
  assign n43768 = ~n43758 & ~n43766;
  assign n43769 = ~n43762 & n43768;
  assign n43770 = ~n43758 & n43767;
  assign n43771 = pi232 & ~n64871;
  assign n43772 = n43739 & ~n43771;
  assign n43773 = ~n35183 & n41902;
  assign n43774 = ~n27583 & n43773;
  assign n43775 = ~pi100 & ~n43774;
  assign n43776 = ~n43772 & n43775;
  assign n43777 = ~n42959 & ~n43773;
  assign n43778 = pi100 & n43777;
  assign n43779 = n6797 & ~n43778;
  assign n43780 = ~n42135 & n43779;
  assign n43781 = ~n43776 & n43780;
  assign n43782 = pi87 & ~n31425;
  assign n43783 = n42139 & ~n43777;
  assign n43784 = ~n43782 & ~n43783;
  assign n43785 = ~n41788 & ~n43784;
  assign n43786 = pi130 & ~n43238;
  assign n43787 = ~pi130 & n43238;
  assign n43788 = ~n43786 & ~n43787;
  assign n43789 = ~n41779 & ~n43788;
  assign n43790 = ~n43785 & ~n43789;
  assign n43791 = ~n43781 & n43790;
  assign n43792 = n64774 & n64792;
  assign n43793 = ~pi51 & ~n43792;
  assign n43794 = ~pi232 & ~n43793;
  assign n43795 = pi39 & ~n43794;
  assign n43796 = ~n2980 & ~n42959;
  assign n43797 = ~n2814 & ~n42036;
  assign n43798 = ~n42437 & ~n43797;
  assign n43799 = ~pi224 & n43798;
  assign n43800 = ~n42074 & n42498;
  assign n43801 = pi224 & n43800;
  assign n43802 = n2980 & ~n43801;
  assign n43803 = pi224 & ~n43800;
  assign n43804 = ~pi224 & ~n43798;
  assign n43805 = ~n43803 & ~n43804;
  assign n43806 = n2980 & ~n43805;
  assign n43807 = ~n43799 & n43802;
  assign n43808 = ~n43796 & ~n64872;
  assign n43809 = pi140 & n43808;
  assign n43810 = n3076 & ~n43798;
  assign n43811 = ~n3076 & ~n42959;
  assign n43812 = ~n3076 & n42959;
  assign n43813 = n2980 & n43799;
  assign n43814 = ~n43812 & ~n43813;
  assign n43815 = ~n43810 & ~n43811;
  assign n43816 = ~pi140 & ~n64873;
  assign n43817 = n33355 & ~n43816;
  assign n43818 = ~n43809 & n43817;
  assign n43819 = ~n35131 & ~n42036;
  assign n43820 = pi169 & n42437;
  assign n43821 = ~n43819 & ~n43820;
  assign n43822 = ~pi216 & ~n43821;
  assign n43823 = ~pi51 & ~n42214;
  assign n43824 = ~pi169 & n43823;
  assign n43825 = pi169 & n43800;
  assign n43826 = pi162 & pi216;
  assign n43827 = ~n43825 & n43826;
  assign n43828 = ~n43824 & n43827;
  assign n43829 = ~n43822 & ~n43828;
  assign n43830 = n2960 & ~n43829;
  assign n43831 = pi169 & n41903;
  assign n43832 = ~pi51 & ~n43831;
  assign n43833 = ~n3056 & ~n43743;
  assign n43834 = ~n43832 & n43833;
  assign n43835 = ~n43830 & ~n43834;
  assign n43836 = pi299 & ~n43835;
  assign n43837 = n64774 & n42429;
  assign n43838 = ~pi51 & ~n43837;
  assign n43839 = pi140 & n43838;
  assign n43840 = ~pi51 & ~n42466;
  assign n43841 = ~pi140 & n43840;
  assign n43842 = n35175 & ~n43841;
  assign n43843 = ~n43839 & n43842;
  assign n43844 = ~n43836 & ~n43843;
  assign n43845 = ~n43818 & n43844;
  assign n43846 = pi232 & ~n43845;
  assign n43847 = n43795 & ~n43846;
  assign n43848 = ~pi232 & ~n41868;
  assign n43849 = ~pi39 & ~n43848;
  assign n43850 = ~n2814 & n41868;
  assign n43851 = ~n42321 & ~n43850;
  assign n43852 = ~n33357 & ~n43851;
  assign n43853 = n33357 & n41868;
  assign n43854 = pi232 & ~n43853;
  assign n43855 = ~n43852 & n43854;
  assign n43856 = n43849 & ~n43855;
  assign n43857 = ~n43847 & ~n43856;
  assign n43858 = ~pi38 & ~n43857;
  assign n43859 = pi38 & ~n43777;
  assign n43860 = ~pi100 & ~n43859;
  assign n43861 = ~n43858 & n43860;
  assign n43862 = n43779 & ~n43861;
  assign n43863 = n43784 & n43789;
  assign n43864 = ~n43862 & n43863;
  assign n43865 = ~n43791 & ~n43864;
  assign n43866 = n62455 & ~n43865;
  assign n43867 = ~pi51 & ~pi87;
  assign n43868 = ~n43831 & n43867;
  assign n43869 = n43789 & n43868;
  assign n43870 = ~pi87 & n41902;
  assign n43871 = ~n41765 & n43867;
  assign n43872 = ~pi87 & ~n33330;
  assign n43873 = n41902 & n43872;
  assign n43874 = ~n33330 & n64874;
  assign n43875 = pi87 & ~n31365;
  assign n43876 = ~n62455 & ~n43875;
  assign n43877 = ~n64875 & n43876;
  assign n43878 = ~n43869 & n43877;
  assign po287 = ~n43866 & ~n43878;
  assign n43880 = n2766 & n6794;
  assign n43881 = pi197 & n42049;
  assign n43882 = ~n2958 & ~n43881;
  assign n43883 = n2961 & ~n43882;
  assign n43884 = ~pi145 & ~n3076;
  assign n43885 = ~pi299 & ~n43884;
  assign n43886 = ~n42456 & n43885;
  assign n43887 = ~n43883 & ~n43886;
  assign n43888 = n62380 & ~n43887;
  assign n43889 = pi232 & ~n43888;
  assign n43890 = n42426 & ~n43889;
  assign n43891 = n64274 & ~n41875;
  assign n43892 = ~n64274 & ~n41948;
  assign n43893 = ~pi39 & ~n43892;
  assign n43894 = ~n43891 & n43893;
  assign n43895 = ~n43890 & ~n43894;
  assign n43896 = ~n2814 & ~n41948;
  assign n43897 = ~n41876 & ~n43896;
  assign n43898 = pi154 & pi232;
  assign n43899 = pi299 & n43898;
  assign n43900 = n43897 & n43899;
  assign n43901 = n41948 & ~n43899;
  assign n43902 = ~pi39 & ~pi176;
  assign n43903 = ~n43901 & n43902;
  assign n43904 = ~n43900 & n43903;
  assign n43905 = n33593 & n43897;
  assign n43906 = ~n33593 & n41948;
  assign n43907 = ~pi39 & pi176;
  assign n43908 = ~n43906 & n43907;
  assign n43909 = ~n43905 & n43908;
  assign n43910 = ~n42425 & ~n43889;
  assign n43911 = pi39 & ~n43910;
  assign n43912 = n43880 & ~n43911;
  assign n43913 = ~n43909 & n43912;
  assign n43914 = ~n43904 & n43913;
  assign n43915 = ~n43904 & n43912;
  assign n43916 = ~n43909 & n43915;
  assign n43917 = n43880 & ~n43895;
  assign n43918 = ~pi133 & ~n42276;
  assign n43919 = ~pi87 & n43918;
  assign n43920 = ~n64876 & n43919;
  assign n43921 = pi145 & n42054;
  assign n43922 = n42558 & ~n43921;
  assign n43923 = n42559 & ~n43881;
  assign n43924 = n41766 & ~n43923;
  assign n43925 = pi299 & ~n43924;
  assign n43926 = ~n43922 & ~n43925;
  assign n43927 = pi232 & ~n43926;
  assign n43928 = n42564 & ~n43927;
  assign n43929 = ~n64274 & n41845;
  assign n43930 = ~pi39 & n41766;
  assign n43931 = ~n43929 & n43930;
  assign n43932 = ~pi38 & ~n43931;
  assign n43933 = ~n43928 & n43932;
  assign n43934 = n41808 & ~n43933;
  assign n43935 = n42136 & ~n43934;
  assign n43936 = ~n42140 & ~n43935;
  assign n43937 = ~n43918 & ~n43936;
  assign n43938 = ~pi183 & ~pi299;
  assign n43939 = ~n35853 & ~n43938;
  assign n43940 = n2815 & n43939;
  assign n43941 = pi87 & ~n43940;
  assign n43942 = ~n43937 & ~n43941;
  assign n43943 = ~n43920 & n43942;
  assign n43944 = n62455 & ~n43943;
  assign n43945 = n41788 & ~n43918;
  assign n43946 = pi87 & n33616;
  assign n43947 = pi149 & n42287;
  assign n43948 = ~n62455 & ~n64877;
  assign n43949 = ~n43945 & n43948;
  assign n43950 = ~n43944 & ~n43949;
  assign n43951 = ~pi136 & n43787;
  assign n43952 = ~pi135 & n43951;
  assign n43953 = pi134 & ~n43952;
  assign n43954 = n41765 & ~n43953;
  assign n43955 = ~n62455 & n43867;
  assign n43956 = n35219 & ~n41765;
  assign n43957 = pi232 & n43956;
  assign n43958 = n43955 & ~n43957;
  assign n43959 = ~n43954 & n43958;
  assign n43960 = ~n35210 & n41902;
  assign n43961 = ~n42959 & ~n43960;
  assign n43962 = ~n2766 & n43961;
  assign n43963 = n6797 & ~n43962;
  assign n43964 = pi232 & ~n35209;
  assign n43965 = n43851 & n43964;
  assign n43966 = ~n41868 & ~n43964;
  assign n43967 = ~pi39 & ~n43966;
  assign n43968 = ~n43965 & n43967;
  assign n43969 = ~pi51 & ~n43956;
  assign n43970 = ~pi164 & pi216;
  assign n43971 = n2960 & ~n43970;
  assign n43972 = ~n43969 & ~n43971;
  assign n43973 = ~n35219 & ~n42036;
  assign n43974 = pi171 & n42437;
  assign n43975 = ~n43973 & ~n43974;
  assign n43976 = ~pi216 & ~n43975;
  assign n43977 = ~pi171 & n43823;
  assign n43978 = pi171 & n43800;
  assign n43979 = pi164 & pi216;
  assign n43980 = ~n43978 & n43979;
  assign n43981 = ~n43977 & n43980;
  assign n43982 = ~n43976 & ~n43981;
  assign n43983 = n2960 & ~n43982;
  assign n43984 = ~n43972 & ~n43983;
  assign n43985 = pi299 & ~n43984;
  assign n43986 = n35200 & ~n43838;
  assign n43987 = n35202 & ~n43808;
  assign n43988 = pi186 & ~n43987;
  assign n43989 = pi186 & ~n43986;
  assign n43990 = ~n43987 & n43989;
  assign n43991 = ~n43986 & n43988;
  assign n43992 = n35202 & n64873;
  assign n43993 = pi39 & pi186;
  assign n43994 = n35200 & ~n43840;
  assign n43995 = ~n43993 & ~n43994;
  assign n43996 = ~n43992 & n43995;
  assign n43997 = ~n64878 & ~n43996;
  assign n43998 = ~n43985 & ~n43997;
  assign n43999 = pi232 & ~n43998;
  assign n44000 = n43795 & ~n43999;
  assign n44001 = n2766 & ~n44000;
  assign n44002 = n2766 & ~n43968;
  assign n44003 = ~n44000 & n44002;
  assign n44004 = ~n43968 & n44001;
  assign n44005 = n43963 & ~n64879;
  assign n44006 = n42139 & ~n43961;
  assign n44007 = n43953 & ~n44006;
  assign n44008 = ~n44005 & n44007;
  assign n44009 = ~n42049 & n43759;
  assign n44010 = n35202 & ~n44009;
  assign n44011 = ~n42608 & n43763;
  assign n44012 = n35200 & ~n44011;
  assign n44013 = ~n44010 & ~n44012;
  assign n44014 = ~n35219 & n43754;
  assign n44015 = pi299 & ~n44014;
  assign n44016 = pi171 & ~n62380;
  assign n44017 = n2814 & n44016;
  assign n44018 = ~n35219 & ~n42063;
  assign n44019 = n31886 & ~n44018;
  assign n44020 = ~n44017 & n44019;
  assign n44021 = n44015 & ~n44020;
  assign n44022 = n44013 & ~n44021;
  assign n44023 = pi232 & ~n44022;
  assign n44024 = ~n43738 & ~n44023;
  assign n44025 = n43993 & ~n44024;
  assign n44026 = n35202 & ~n43759;
  assign n44027 = n35200 & ~n43763;
  assign n44028 = ~n44026 & ~n44027;
  assign n44029 = ~n44021 & n44028;
  assign n44030 = pi232 & ~n44029;
  assign n44031 = ~n43738 & ~n44030;
  assign n44032 = pi39 & ~pi186;
  assign n44033 = ~n44031 & n44032;
  assign n44034 = ~pi39 & ~n43960;
  assign n44035 = ~pi164 & ~n44034;
  assign n44036 = ~n44033 & n44035;
  assign n44037 = ~n44025 & n44036;
  assign n44038 = n43993 & ~n44013;
  assign n44039 = ~n44028 & n44032;
  assign n44040 = ~n44038 & ~n44039;
  assign n44041 = pi232 & ~n44040;
  assign n44042 = pi164 & ~n44034;
  assign n44043 = pi171 & ~n43741;
  assign n44044 = ~pi171 & ~n42607;
  assign n44045 = n31886 & ~n44044;
  assign n44046 = ~n44043 & n44045;
  assign n44047 = pi232 & n44015;
  assign n44048 = ~n44046 & n44047;
  assign n44049 = ~n43738 & ~n44048;
  assign n44050 = pi39 & ~n44049;
  assign n44051 = n44042 & ~n44050;
  assign n44052 = pi186 & n44013;
  assign n44053 = ~pi186 & n44028;
  assign n44054 = pi232 & ~n44053;
  assign n44055 = ~n44052 & n44054;
  assign n44056 = n44049 & ~n44055;
  assign n44057 = pi39 & ~n44056;
  assign n44058 = n44042 & ~n44057;
  assign n44059 = n44015 & ~n44046;
  assign n44060 = n44013 & ~n44059;
  assign n44061 = pi232 & ~n44060;
  assign n44062 = ~n43738 & ~n44061;
  assign n44063 = n43993 & ~n44062;
  assign n44064 = n44028 & ~n44059;
  assign n44065 = pi232 & ~n44064;
  assign n44066 = ~n43738 & ~n44065;
  assign n44067 = n44032 & ~n44066;
  assign n44068 = n44042 & ~n44067;
  assign n44069 = ~n44063 & n44068;
  assign n44070 = ~n44041 & n44051;
  assign n44071 = n2766 & ~n64880;
  assign n44072 = n2766 & ~n44037;
  assign n44073 = ~n64880 & n44072;
  assign n44074 = ~n44037 & n44071;
  assign n44075 = ~n43148 & n43963;
  assign n44076 = ~n64881 & n44075;
  assign n44077 = n42139 & n43960;
  assign n44078 = ~n43953 & ~n44077;
  assign n44079 = ~n44076 & n44078;
  assign n44080 = n62455 & ~n44079;
  assign n44081 = n62455 & ~n44008;
  assign n44082 = ~n44079 & n44081;
  assign n44083 = ~n44008 & n44080;
  assign n44084 = ~n43959 & ~n64882;
  assign n44085 = ~n35284 & ~n42036;
  assign n44086 = pi170 & n42437;
  assign n44087 = n3056 & ~n44086;
  assign n44088 = ~n44085 & n44087;
  assign n44089 = ~n31886 & ~n44088;
  assign n44090 = ~pi170 & n43823;
  assign n44091 = pi170 & n43800;
  assign n44092 = pi216 & ~n44091;
  assign n44093 = ~n44090 & n44092;
  assign n44094 = ~n44089 & ~n44093;
  assign n44095 = pi150 & pi299;
  assign n44096 = n35284 & ~n41765;
  assign n44097 = ~pi51 & ~n44096;
  assign n44098 = ~n2960 & n44097;
  assign n44099 = n44095 & ~n44098;
  assign n44100 = ~n44094 & n44099;
  assign n44101 = ~n3056 & n44097;
  assign n44102 = n43157 & ~n44101;
  assign n44103 = ~n44088 & n44102;
  assign n44104 = ~n44100 & ~n44103;
  assign n44105 = pi185 & n43838;
  assign n44106 = ~pi185 & n43840;
  assign n44107 = ~pi299 & ~n44106;
  assign n44108 = ~n44105 & n44107;
  assign n44109 = n44104 & ~n44108;
  assign n44110 = pi232 & ~n44109;
  assign n44111 = n43795 & ~n44110;
  assign n44112 = ~pi299 & ~n41868;
  assign n44113 = pi170 & ~n43851;
  assign n44114 = ~pi170 & n41868;
  assign n44115 = n35283 & ~n44114;
  assign n44116 = ~n44113 & n44115;
  assign n44117 = n43849 & ~n44116;
  assign n44118 = ~n44112 & n44117;
  assign n44119 = ~n44111 & ~n44118;
  assign n44120 = ~pi38 & ~n44119;
  assign n44121 = ~n35321 & n41902;
  assign n44122 = ~n42959 & ~n44121;
  assign n44123 = pi38 & ~n44122;
  assign n44124 = ~pi194 & ~n44123;
  assign n44125 = ~n44120 & n44124;
  assign n44126 = pi185 & n43808;
  assign n44127 = ~pi185 & ~n64873;
  assign n44128 = ~pi299 & ~n44127;
  assign n44129 = ~pi299 & ~n44126;
  assign n44130 = ~n44127 & n44129;
  assign n44131 = ~n44126 & n44128;
  assign n44132 = n44104 & ~n64883;
  assign n44133 = pi232 & ~n44132;
  assign n44134 = n43795 & ~n44133;
  assign n44135 = n35103 & n43851;
  assign n44136 = n44117 & ~n44135;
  assign n44137 = ~n44134 & ~n44136;
  assign n44138 = ~pi38 & ~n44137;
  assign n44139 = n35329 & n41902;
  assign n44140 = ~n42959 & ~n44139;
  assign n44141 = pi38 & ~n44140;
  assign n44142 = pi194 & ~n44141;
  assign n44143 = ~n44138 & n44142;
  assign n44144 = ~n44125 & ~n44143;
  assign n44145 = ~pi100 & ~n44144;
  assign n44146 = pi194 & n31977;
  assign n44147 = n44121 & ~n44146;
  assign n44148 = ~n42959 & ~n44147;
  assign n44149 = pi100 & n44148;
  assign n44150 = n6797 & ~n44149;
  assign n44151 = ~n44145 & n44150;
  assign n44152 = pi135 & ~n43951;
  assign n44153 = pi134 & n43952;
  assign n44154 = ~n44152 & ~n44153;
  assign n44155 = n42139 & ~n44148;
  assign n44156 = ~n44154 & ~n44155;
  assign n44157 = ~n44151 & n44156;
  assign n44158 = pi185 & n42608;
  assign n44159 = n43763 & ~n44158;
  assign n44160 = ~n27583 & n44121;
  assign n44161 = ~pi194 & ~n44160;
  assign n44162 = ~n44159 & n44161;
  assign n44163 = ~n27583 & n44139;
  assign n44164 = pi194 & ~n44163;
  assign n44165 = pi185 & n42049;
  assign n44166 = n43759 & ~n44165;
  assign n44167 = ~pi185 & n43759;
  assign n44168 = ~n44009 & n44164;
  assign n44169 = ~n44167 & n44168;
  assign n44170 = n44164 & ~n44166;
  assign n44171 = ~n44162 & ~n64884;
  assign n44172 = ~pi299 & ~n44171;
  assign n44173 = pi170 & ~n43741;
  assign n44174 = ~pi170 & ~n42607;
  assign n44175 = n31886 & ~n44174;
  assign n44176 = ~n44173 & n44175;
  assign n44177 = n44095 & ~n44176;
  assign n44178 = pi170 & ~n62380;
  assign n44179 = n2814 & n44178;
  assign n44180 = ~n35284 & ~n42063;
  assign n44181 = n31886 & ~n44180;
  assign n44182 = ~n44179 & n44181;
  assign n44183 = n43157 & ~n44182;
  assign n44184 = ~n44177 & ~n44183;
  assign n44185 = ~n35284 & n43754;
  assign n44186 = ~n44161 & ~n44164;
  assign n44187 = ~n44185 & ~n44186;
  assign n44188 = ~n44184 & n44187;
  assign n44189 = ~n44172 & ~n44188;
  assign n44190 = pi232 & ~n44189;
  assign n44191 = ~n43739 & ~n44186;
  assign n44192 = ~n44190 & ~n44191;
  assign n44193 = ~pi100 & ~n44192;
  assign n44194 = ~n42135 & n44150;
  assign n44195 = n42136 & ~n44149;
  assign n44196 = ~n44193 & n64885;
  assign n44197 = n42139 & n44147;
  assign n44198 = n44154 & ~n44197;
  assign n44199 = ~n44196 & n44198;
  assign n44200 = n62455 & ~n44199;
  assign n44201 = ~n44157 & n44200;
  assign n44202 = n41765 & n44154;
  assign n44203 = n35328 & ~n41765;
  assign n44204 = pi232 & n44096;
  assign n44205 = n43955 & ~n64886;
  assign n44206 = ~n44202 & n44205;
  assign n44207 = ~n44201 & ~n44206;
  assign n44208 = pi136 & ~n43787;
  assign n44209 = ~n43951 & ~n44208;
  assign n44210 = ~n41778 & ~n44209;
  assign n44211 = ~n41902 & n44210;
  assign n44212 = pi148 & n2815;
  assign n44213 = ~n41765 & ~n44212;
  assign n44214 = ~n44211 & ~n44213;
  assign n44215 = n43955 & ~n44214;
  assign n44216 = ~n31413 & ~n43851;
  assign n44217 = n31413 & n41868;
  assign n44218 = pi232 & ~n44217;
  assign n44219 = ~n44216 & n44218;
  assign n44220 = n43849 & ~n44219;
  assign n44221 = pi184 & n43808;
  assign n44222 = ~pi184 & ~n64873;
  assign n44223 = n31411 & ~n44222;
  assign n44224 = ~n44221 & n44223;
  assign n44225 = pi184 & n43838;
  assign n44226 = ~pi141 & ~pi299;
  assign n44227 = ~pi184 & n43840;
  assign n44228 = n44226 & ~n44227;
  assign n44229 = ~n44225 & n44228;
  assign n44230 = n3056 & ~n43798;
  assign n44231 = pi163 & n2960;
  assign n44232 = ~n43800 & n44231;
  assign n44233 = ~n3056 & ~n44231;
  assign n44234 = ~n42959 & n44233;
  assign n44235 = pi148 & ~n44234;
  assign n44236 = n43800 & n44231;
  assign n44237 = ~n2960 & n42959;
  assign n44238 = ~n3056 & ~n42959;
  assign n44239 = ~pi163 & ~n44238;
  assign n44240 = ~n44237 & ~n44239;
  assign n44241 = ~n44236 & n44240;
  assign n44242 = pi148 & ~n44241;
  assign n44243 = ~n44232 & n44235;
  assign n44244 = ~n44230 & n64887;
  assign n44245 = ~pi287 & n32931;
  assign n44246 = pi216 & ~n44245;
  assign n44247 = n2960 & ~n44246;
  assign n44248 = n64774 & n44247;
  assign n44249 = ~pi51 & ~pi148;
  assign n44250 = ~n44248 & n44249;
  assign n44251 = pi299 & ~n44250;
  assign n44252 = ~n44244 & n44251;
  assign n44253 = ~n44229 & ~n44252;
  assign n44254 = ~n44224 & n44253;
  assign n44255 = pi232 & ~n44254;
  assign n44256 = n43795 & ~n44255;
  assign n44257 = n2766 & ~n44256;
  assign n44258 = ~n44220 & n44257;
  assign n44259 = n31414 & ~n41765;
  assign n44260 = ~pi51 & ~n44259;
  assign n44261 = ~n2766 & ~n44260;
  assign n44262 = n6797 & ~n44261;
  assign n44263 = ~n44258 & n44262;
  assign n44264 = n42139 & n44260;
  assign n44265 = n44210 & ~n44264;
  assign n44266 = ~n44263 & n44265;
  assign n44267 = ~n38958 & ~n41765;
  assign n44268 = n44260 & n44267;
  assign n44269 = ~pi51 & n42559;
  assign n44270 = ~pi148 & ~n44269;
  assign n44271 = ~n44245 & ~n44270;
  assign n44272 = ~pi148 & n41902;
  assign n44273 = ~n44271 & ~n44272;
  assign n44274 = n31886 & n43740;
  assign n44275 = ~n2814 & n43754;
  assign n44276 = pi148 & ~n44275;
  assign n44277 = ~n44274 & n44276;
  assign n44278 = ~n44273 & ~n44277;
  assign n44279 = pi299 & ~n44278;
  assign n44280 = pi184 & n42049;
  assign n44281 = n43759 & ~n44280;
  assign n44282 = n31411 & ~n44281;
  assign n44283 = pi184 & n42608;
  assign n44284 = n43763 & ~n44283;
  assign n44285 = n44226 & ~n44284;
  assign n44286 = ~n44282 & ~n44285;
  assign n44287 = ~n44279 & ~n44285;
  assign n44288 = ~n44282 & n44287;
  assign n44289 = ~n44279 & n44286;
  assign n44290 = pi232 & ~n64888;
  assign n44291 = ~pi100 & n43739;
  assign n44292 = ~n44290 & n44291;
  assign n44293 = ~n44268 & ~n44292;
  assign n44294 = n6797 & ~n44293;
  assign n44295 = ~n41765 & n44264;
  assign n44296 = ~n44210 & ~n44295;
  assign n44297 = ~n44294 & n44296;
  assign n44298 = n62455 & ~n44297;
  assign n44299 = ~n44266 & n44298;
  assign n44300 = ~n44215 & ~n44299;
  assign n44301 = pi215 & pi1142;
  assign n44302 = pi299 & ~n44301;
  assign n44303 = ~pi932 & n41020;
  assign n44304 = ~pi1142 & ~n41020;
  assign n44305 = pi221 & ~n44304;
  assign n44306 = pi221 & ~n44303;
  assign n44307 = ~n44304 & n44306;
  assign n44308 = ~n44303 & n44305;
  assign n44309 = pi216 & pi277;
  assign n44310 = ~pi221 & ~n44309;
  assign n44311 = ~pi72 & ~n43700;
  assign n44312 = ~n30618 & ~n44311;
  assign n44313 = n2750 & ~n44312;
  assign n44314 = n43566 & ~n44313;
  assign n44315 = ~pi95 & ~n44314;
  assign n44316 = n41047 & ~n44315;
  assign n44317 = ~pi262 & n44316;
  assign n44318 = pi172 & ~n44317;
  assign n44319 = pi262 & n43705;
  assign n44320 = n2728 & n33867;
  assign n44321 = ~n30613 & ~n44320;
  assign n44322 = ~pi262 & n44321;
  assign n44323 = ~pi172 & ~n33962;
  assign n44324 = ~n44322 & n44323;
  assign n44325 = ~n44319 & n44324;
  assign n44326 = ~pi228 & ~n44325;
  assign n44327 = ~n33962 & ~n44321;
  assign n44328 = ~pi262 & n44327;
  assign n44329 = ~pi172 & ~n44328;
  assign n44330 = pi172 & ~pi262;
  assign n44331 = n44316 & n44330;
  assign n44332 = ~n44329 & ~n44331;
  assign n44333 = pi262 & n43706;
  assign n44334 = ~pi228 & ~n44333;
  assign n44335 = ~n44332 & n44334;
  assign n44336 = ~n44318 & n44326;
  assign n44337 = pi105 & ~n44321;
  assign n44338 = pi262 & ~n30613;
  assign n44339 = pi105 & n44338;
  assign n44340 = ~n44320 & n44339;
  assign n44341 = ~pi105 & pi172;
  assign n44342 = pi228 & ~n44341;
  assign n44343 = ~n44340 & n44342;
  assign n44344 = ~n44337 & n44343;
  assign n44345 = ~pi216 & ~n44344;
  assign n44346 = ~n64890 & n44345;
  assign n44347 = n44310 & ~n44346;
  assign n44348 = ~n64889 & ~n44347;
  assign n44349 = ~pi215 & ~n44348;
  assign n44350 = n44302 & ~n44349;
  assign n44351 = pi223 & pi1142;
  assign n44352 = ~pi299 & ~n44351;
  assign n44353 = ~pi932 & n41469;
  assign n44354 = ~pi1142 & ~n41469;
  assign n44355 = pi222 & ~n44354;
  assign n44356 = pi222 & ~n44353;
  assign n44357 = ~n44354 & n44356;
  assign n44358 = ~n44353 & n44355;
  assign n44359 = pi224 & pi277;
  assign n44360 = ~pi222 & ~n44359;
  assign n44361 = ~pi224 & ~n44322;
  assign n44362 = n44360 & ~n44361;
  assign n44363 = ~n64891 & ~n44362;
  assign n44364 = n44352 & n44363;
  assign n44365 = ~n44321 & n44360;
  assign n44366 = n44363 & ~n44365;
  assign n44367 = ~pi223 & ~n44366;
  assign n44368 = n44352 & ~n44367;
  assign n44369 = ~pi39 & ~n44368;
  assign n44370 = ~n44364 & n44369;
  assign n44371 = ~n44350 & n44370;
  assign n44372 = n30613 & n38189;
  assign n44373 = ~pi224 & n44338;
  assign n44374 = n44360 & ~n44373;
  assign n44375 = ~n64891 & ~n44374;
  assign n44376 = ~pi223 & ~n44375;
  assign n44377 = ~n44351 & ~n44376;
  assign n44378 = ~pi299 & ~n44377;
  assign n44379 = ~n44372 & n44378;
  assign n44380 = ~pi262 & n62380;
  assign n44381 = pi172 & ~pi228;
  assign n44382 = ~n34059 & ~n44381;
  assign n44383 = ~n44380 & ~n44382;
  assign n44384 = n30613 & n41010;
  assign n44385 = ~n44339 & ~n44341;
  assign n44386 = pi228 & ~n44385;
  assign n44387 = ~n44384 & ~n44386;
  assign n44388 = ~n44383 & n44387;
  assign n44389 = ~pi216 & ~n44388;
  assign n44390 = n44310 & ~n44389;
  assign n44391 = ~n64889 & ~n44390;
  assign n44392 = ~pi215 & ~n44391;
  assign n44393 = ~n44301 & ~n44392;
  assign n44394 = pi299 & ~n44393;
  assign n44395 = ~n44379 & ~n44394;
  assign n44396 = pi39 & ~n44395;
  assign n44397 = ~pi38 & ~n44396;
  assign n44398 = ~n44371 & n44397;
  assign n44399 = n38199 & n44384;
  assign n44400 = ~n44381 & ~n44386;
  assign n44401 = ~pi216 & ~n44400;
  assign n44402 = n44310 & ~n44401;
  assign n44403 = ~n64889 & ~n44402;
  assign n44404 = ~pi215 & ~n44403;
  assign n44405 = ~n44301 & ~n44404;
  assign n44406 = ~n44399 & ~n44405;
  assign n44407 = pi299 & n44406;
  assign n44408 = ~n44379 & ~n44407;
  assign n44409 = pi38 & n44408;
  assign n44410 = ~pi100 & ~n44409;
  assign n44411 = ~n44398 & n44410;
  assign n44412 = pi146 & pi252;
  assign n44413 = pi146 & ~n30857;
  assign n44414 = ~pi146 & ~n62380;
  assign n44415 = ~n44413 & ~n44414;
  assign n44416 = n62380 & ~n44412;
  assign n44417 = pi152 & ~n64892;
  assign n44418 = ~n40506 & n64892;
  assign n44419 = n30857 & n40506;
  assign n44420 = ~pi152 & ~n44419;
  assign n44421 = ~n44418 & n44420;
  assign n44422 = ~n44417 & ~n44421;
  assign n44423 = ~pi262 & n44422;
  assign n44424 = ~pi228 & n44422;
  assign n44425 = ~n44381 & ~n44424;
  assign n44426 = ~n44423 & ~n44425;
  assign n44427 = n44387 & ~n44426;
  assign n44428 = ~pi216 & ~n44427;
  assign n44429 = n44310 & ~n44428;
  assign n44430 = ~n64889 & ~n44429;
  assign n44431 = ~pi215 & ~n44430;
  assign n44432 = ~n44301 & ~n44431;
  assign n44433 = pi299 & ~n44432;
  assign n44434 = n2764 & ~n44379;
  assign n44435 = ~n44433 & n44434;
  assign n44436 = ~n2764 & n44408;
  assign n44437 = pi100 & ~n44436;
  assign n44438 = ~n44435 & n44437;
  assign n44439 = ~n44411 & ~n44438;
  assign n44440 = ~pi87 & ~n44439;
  assign n44441 = ~n62373 & n44408;
  assign n44442 = n62373 & n44395;
  assign n44443 = ~n44441 & ~n44442;
  assign n44444 = pi87 & n44443;
  assign n44445 = ~pi75 & ~n44444;
  assign n44446 = ~n44440 & n44445;
  assign n44447 = pi75 & n44408;
  assign n44448 = ~pi92 & ~n44447;
  assign n44449 = ~n44446 & n44448;
  assign n44450 = n6795 & ~n44443;
  assign n44451 = ~n6795 & n44408;
  assign n44452 = pi92 & ~n44451;
  assign n44453 = ~n44450 & n44452;
  assign n44454 = n6792 & ~n44453;
  assign n44455 = ~n44449 & n44454;
  assign n44456 = ~n6792 & n44408;
  assign n44457 = ~pi55 & ~n44456;
  assign n44458 = ~n44455 & n44457;
  assign n44459 = n64082 & n44393;
  assign n44460 = ~n64082 & ~n44406;
  assign n44461 = pi55 & ~n44460;
  assign n44462 = ~n44459 & n44461;
  assign n44463 = ~pi56 & ~n44462;
  assign n44464 = ~n44458 & n44463;
  assign n44465 = n64084 & ~n44393;
  assign n44466 = ~n64084 & n44406;
  assign n44467 = pi56 & ~n44466;
  assign n44468 = ~n64084 & ~n44406;
  assign n44469 = ~pi55 & n44459;
  assign n44470 = ~n44468 & ~n44469;
  assign n44471 = pi56 & ~n44470;
  assign n44472 = ~n44465 & n44467;
  assign n44473 = ~pi62 & ~n64893;
  assign n44474 = ~n44464 & n44473;
  assign n44475 = n62373 & n34046;
  assign n44476 = n44393 & n44475;
  assign n44477 = ~n44406 & ~n44475;
  assign n44478 = pi62 & ~n44477;
  assign n44479 = ~n44476 & n44478;
  assign n44480 = n3472 & ~n44479;
  assign n44481 = ~n44474 & n44480;
  assign n44482 = ~n3472 & ~n44406;
  assign n44483 = ~pi249 & ~n44482;
  assign n44484 = ~n44481 & n44483;
  assign n44485 = pi262 & n44316;
  assign n44486 = ~pi172 & ~n44485;
  assign n44487 = ~pi262 & ~n43706;
  assign n44488 = pi262 & ~n44327;
  assign n44489 = pi172 & ~n44488;
  assign n44490 = ~n44487 & n44489;
  assign n44491 = ~n44486 & ~n44490;
  assign n44492 = ~pi228 & ~n44491;
  assign n44493 = ~pi216 & ~n44343;
  assign n44494 = ~n44492 & n44493;
  assign n44495 = n44310 & ~n44494;
  assign n44496 = ~n64889 & ~n44495;
  assign n44497 = ~pi215 & ~n44496;
  assign n44498 = n44302 & ~n44497;
  assign n44499 = n44369 & ~n44498;
  assign n44500 = ~n44383 & ~n44386;
  assign n44501 = ~pi216 & ~n44500;
  assign n44502 = n44310 & ~n44501;
  assign n44503 = ~n64889 & ~n44502;
  assign n44504 = ~pi215 & ~n44503;
  assign n44505 = ~n44301 & ~n44504;
  assign n44506 = pi299 & ~n44505;
  assign n44507 = ~n44378 & ~n44506;
  assign n44508 = pi39 & ~n44507;
  assign n44509 = ~pi38 & ~n44508;
  assign n44510 = ~n44499 & n44509;
  assign n44511 = pi299 & ~n44405;
  assign n44512 = ~n44378 & ~n44511;
  assign n44513 = pi38 & n44512;
  assign n44514 = ~pi100 & ~n44513;
  assign n44515 = ~n44510 & n44514;
  assign n44516 = ~n44386 & ~n44426;
  assign n44517 = ~pi216 & ~n44516;
  assign n44518 = n44310 & ~n44517;
  assign n44519 = ~n64889 & ~n44518;
  assign n44520 = ~pi215 & ~n44519;
  assign n44521 = ~n44301 & ~n44520;
  assign n44522 = pi299 & ~n44521;
  assign n44523 = n2764 & ~n44378;
  assign n44524 = ~n44522 & n44523;
  assign n44525 = ~n2764 & n44512;
  assign n44526 = pi100 & ~n44525;
  assign n44527 = ~n44524 & n44526;
  assign n44528 = ~n44515 & ~n44527;
  assign n44529 = ~pi87 & ~n44528;
  assign n44530 = ~n62373 & n44512;
  assign n44531 = n62373 & n44507;
  assign n44532 = ~n44530 & ~n44531;
  assign n44533 = pi87 & n44532;
  assign n44534 = ~pi75 & ~n44533;
  assign n44535 = ~n44529 & n44534;
  assign n44536 = pi75 & n44512;
  assign n44537 = ~pi92 & ~n44536;
  assign n44538 = ~n44535 & n44537;
  assign n44539 = n6795 & ~n44532;
  assign n44540 = ~n6795 & n44512;
  assign n44541 = pi92 & ~n44540;
  assign n44542 = ~n44539 & n44541;
  assign n44543 = n6792 & ~n44542;
  assign n44544 = ~n44538 & n44543;
  assign n44545 = ~n6792 & n44512;
  assign n44546 = ~pi55 & ~n44545;
  assign n44547 = ~n44544 & n44546;
  assign n44548 = n64082 & n44505;
  assign n44549 = ~n64082 & n44405;
  assign n44550 = pi55 & ~n44549;
  assign n44551 = ~n44548 & n44550;
  assign n44552 = ~pi56 & ~n44551;
  assign n44553 = ~n44547 & n44552;
  assign n44554 = n64084 & ~n44505;
  assign n44555 = ~n64084 & ~n44405;
  assign n44556 = pi56 & ~n44555;
  assign n44557 = ~n64084 & n44405;
  assign n44558 = ~pi55 & n44548;
  assign n44559 = ~n44557 & ~n44558;
  assign n44560 = pi56 & ~n44559;
  assign n44561 = ~n44554 & n44556;
  assign n44562 = ~pi62 & ~n64894;
  assign n44563 = ~n44553 & n44562;
  assign n44564 = n44475 & n44505;
  assign n44565 = n44405 & ~n44475;
  assign n44566 = pi62 & ~n44565;
  assign n44567 = ~n44564 & n44566;
  assign n44568 = n3472 & ~n44567;
  assign n44569 = ~n44563 & n44568;
  assign n44570 = ~n3472 & n44405;
  assign n44571 = pi249 & ~n44570;
  assign n44572 = ~n44569 & n44571;
  assign n44573 = ~n44484 & ~n44572;
  assign n44574 = pi223 & pi1141;
  assign n44575 = ~pi299 & ~n44574;
  assign n44576 = ~pi935 & n41469;
  assign n44577 = ~pi1141 & ~n41469;
  assign n44578 = pi222 & ~n44577;
  assign n44579 = pi222 & ~n44576;
  assign n44580 = ~n44577 & n44579;
  assign n44581 = ~n44576 & n44578;
  assign n44582 = pi224 & pi270;
  assign n44583 = ~pi222 & ~n44582;
  assign n44584 = pi861 & n44321;
  assign n44585 = ~pi224 & ~n44584;
  assign n44586 = n44583 & ~n44585;
  assign n44587 = ~n64895 & ~n44586;
  assign n44588 = ~n44321 & n44583;
  assign n44589 = n44587 & ~n44588;
  assign n44590 = ~pi223 & ~n44589;
  assign n44591 = n44575 & ~n44590;
  assign n44592 = ~pi39 & ~n44591;
  assign n44593 = pi215 & pi1141;
  assign n44594 = pi299 & ~n44593;
  assign n44595 = ~pi935 & n41020;
  assign n44596 = ~pi1141 & ~n41020;
  assign n44597 = pi221 & ~n44596;
  assign n44598 = pi221 & ~n44595;
  assign n44599 = ~n44596 & n44598;
  assign n44600 = ~n44595 & n44597;
  assign n44601 = pi216 & pi270;
  assign n44602 = ~pi221 & ~n44601;
  assign n44603 = ~pi861 & n44316;
  assign n44604 = ~pi171 & ~n44603;
  assign n44605 = pi861 & ~n43706;
  assign n44606 = ~pi861 & ~n44327;
  assign n44607 = pi171 & ~n44606;
  assign n44608 = ~n44605 & n44607;
  assign n44609 = ~n44604 & ~n44608;
  assign n44610 = ~pi228 & ~n44609;
  assign n44611 = n41010 & ~n44321;
  assign n44612 = pi861 & ~n30613;
  assign n44613 = pi105 & ~n44612;
  assign n44614 = ~pi105 & pi171;
  assign n44615 = pi228 & ~n44614;
  assign n44616 = ~n44613 & n44615;
  assign n44617 = ~pi216 & ~n44616;
  assign n44618 = ~n44611 & n44617;
  assign n44619 = ~n44610 & n44618;
  assign n44620 = n44602 & ~n44619;
  assign n44621 = ~n64896 & ~n44620;
  assign n44622 = ~pi215 & ~n44621;
  assign n44623 = n44594 & ~n44622;
  assign n44624 = n44592 & ~n44623;
  assign n44625 = ~pi299 & n44372;
  assign n44626 = n30613 & n38188;
  assign n44627 = ~pi224 & ~n44612;
  assign n44628 = n44583 & ~n44627;
  assign n44629 = ~n64895 & ~n44628;
  assign n44630 = ~pi223 & ~n44629;
  assign n44631 = ~n44574 & ~n44630;
  assign n44632 = ~pi299 & ~n44631;
  assign n44633 = ~n64897 & ~n44632;
  assign n44634 = ~pi861 & n62380;
  assign n44635 = ~pi228 & ~n44634;
  assign n44636 = ~pi228 & ~n44016;
  assign n44637 = ~n44634 & n44636;
  assign n44638 = ~n44016 & n44635;
  assign n44639 = ~n44384 & n44617;
  assign n44640 = ~n64898 & n44639;
  assign n44641 = n44602 & ~n44640;
  assign n44642 = ~n64896 & ~n44641;
  assign n44643 = ~pi215 & ~n44642;
  assign n44644 = ~n44593 & ~n44643;
  assign n44645 = pi299 & ~n44644;
  assign n44646 = n44633 & ~n44645;
  assign n44647 = pi39 & ~n44646;
  assign n44648 = ~pi38 & ~n44647;
  assign n44649 = ~n44624 & n44648;
  assign n44650 = ~pi171 & ~pi228;
  assign n44651 = n44617 & ~n44650;
  assign n44652 = n44602 & ~n44651;
  assign n44653 = ~n64896 & ~n44652;
  assign n44654 = ~pi215 & ~n44653;
  assign n44655 = ~n44593 & ~n44654;
  assign n44656 = n41037 & n44384;
  assign n44657 = ~n44601 & n44656;
  assign n44658 = n44655 & ~n44657;
  assign n44659 = pi299 & ~n44658;
  assign n44660 = n44633 & ~n44659;
  assign n44661 = pi38 & n44660;
  assign n44662 = ~pi100 & ~n44661;
  assign n44663 = ~n44649 & n44662;
  assign n44664 = pi171 & ~n44422;
  assign n44665 = ~pi861 & n44422;
  assign n44666 = ~pi228 & ~n44665;
  assign n44667 = ~pi228 & ~n44664;
  assign n44668 = ~n44665 & n44667;
  assign n44669 = ~n44664 & n44666;
  assign n44670 = n44639 & ~n64899;
  assign n44671 = n44602 & ~n44670;
  assign n44672 = ~n64896 & ~n44671;
  assign n44673 = ~pi215 & ~n44672;
  assign n44674 = ~n44593 & ~n44673;
  assign n44675 = pi299 & ~n44674;
  assign n44676 = n2764 & n44633;
  assign n44677 = ~n44675 & n44676;
  assign n44678 = ~n2764 & n44660;
  assign n44679 = pi100 & ~n44678;
  assign n44680 = ~n44677 & n44679;
  assign n44681 = ~n44663 & ~n44680;
  assign n44682 = ~pi87 & ~n44681;
  assign n44683 = ~n62373 & n44660;
  assign n44684 = n62373 & n44646;
  assign n44685 = ~n44683 & ~n44684;
  assign n44686 = pi87 & n44685;
  assign n44687 = ~pi75 & ~n44686;
  assign n44688 = ~n44682 & n44687;
  assign n44689 = pi75 & n44660;
  assign n44690 = ~pi92 & ~n44689;
  assign n44691 = ~n44688 & n44690;
  assign n44692 = n6795 & ~n44685;
  assign n44693 = ~n6795 & n44660;
  assign n44694 = pi92 & ~n44693;
  assign n44695 = ~n44692 & n44694;
  assign n44696 = n6792 & ~n44695;
  assign n44697 = ~n44691 & n44696;
  assign n44698 = ~n6792 & n44660;
  assign n44699 = ~pi55 & ~n44698;
  assign n44700 = ~n44697 & n44699;
  assign n44701 = n64082 & n44644;
  assign n44702 = ~n64082 & n44658;
  assign n44703 = pi55 & ~n44702;
  assign n44704 = ~n44701 & n44703;
  assign n44705 = ~pi56 & ~n44704;
  assign n44706 = ~n44700 & n44705;
  assign n44707 = n64084 & ~n44644;
  assign n44708 = ~n64084 & ~n44658;
  assign n44709 = pi56 & ~n44708;
  assign n44710 = ~pi55 & n44701;
  assign n44711 = ~n64084 & n44658;
  assign n44712 = ~n44710 & ~n44711;
  assign n44713 = pi56 & ~n44712;
  assign n44714 = ~n44707 & n44709;
  assign n44715 = ~pi62 & ~n64900;
  assign n44716 = ~n44706 & n44715;
  assign n44717 = n44475 & n44644;
  assign n44718 = ~n44475 & n44658;
  assign n44719 = pi62 & ~n44718;
  assign n44720 = ~n44717 & n44719;
  assign n44721 = pi241 & n3472;
  assign n44722 = ~n44720 & n44721;
  assign n44723 = ~n44716 & n44722;
  assign n44724 = ~pi861 & n43705;
  assign n44725 = ~n33962 & ~n44584;
  assign n44726 = ~n44724 & n44725;
  assign n44727 = pi861 & n44327;
  assign n44728 = ~pi171 & ~n44727;
  assign n44729 = ~pi861 & n43706;
  assign n44730 = n44728 & ~n44729;
  assign n44731 = ~pi171 & ~n44726;
  assign n44732 = pi171 & pi861;
  assign n44733 = n44316 & n44732;
  assign n44734 = pi171 & n44316;
  assign n44735 = ~n44728 & ~n44734;
  assign n44736 = pi861 & ~n44735;
  assign n44737 = ~n43706 & n44728;
  assign n44738 = ~n44736 & ~n44737;
  assign n44739 = ~n64901 & ~n44733;
  assign n44740 = ~pi228 & ~n64902;
  assign n44741 = ~n44337 & n44616;
  assign n44742 = ~pi216 & ~n44741;
  assign n44743 = ~n44740 & n44742;
  assign n44744 = n44602 & ~n44743;
  assign n44745 = ~n64896 & ~n44744;
  assign n44746 = ~pi215 & ~n44745;
  assign n44747 = n44594 & ~n44746;
  assign n44748 = n44575 & n44587;
  assign n44749 = n44592 & ~n44748;
  assign n44750 = ~n44747 & n44749;
  assign n44751 = n44617 & ~n64898;
  assign n44752 = n44602 & ~n44751;
  assign n44753 = ~n64896 & ~n44752;
  assign n44754 = ~pi215 & ~n44753;
  assign n44755 = ~n44593 & ~n44754;
  assign n44756 = pi299 & ~n44755;
  assign n44757 = ~n44632 & ~n44756;
  assign n44758 = pi39 & ~n44757;
  assign n44759 = ~pi38 & ~n44758;
  assign n44760 = ~n44750 & n44759;
  assign n44761 = pi299 & ~n44655;
  assign n44762 = ~n44632 & ~n44761;
  assign n44763 = pi38 & n44762;
  assign n44764 = ~pi100 & ~n44763;
  assign n44765 = ~n44760 & n44764;
  assign n44766 = n44617 & ~n64899;
  assign n44767 = n44602 & ~n44766;
  assign n44768 = ~n64896 & ~n44767;
  assign n44769 = ~pi215 & ~n44768;
  assign n44770 = ~n44593 & ~n44769;
  assign n44771 = pi299 & ~n44770;
  assign n44772 = n2764 & ~n44632;
  assign n44773 = ~n44771 & n44772;
  assign n44774 = ~n2764 & n44762;
  assign n44775 = pi100 & ~n44774;
  assign n44776 = ~n44773 & n44775;
  assign n44777 = ~n44765 & ~n44776;
  assign n44778 = ~pi87 & ~n44777;
  assign n44779 = ~n62373 & n44762;
  assign n44780 = n62373 & n44757;
  assign n44781 = ~n44779 & ~n44780;
  assign n44782 = pi87 & n44781;
  assign n44783 = ~pi75 & ~n44782;
  assign n44784 = ~n44778 & n44783;
  assign n44785 = pi75 & n44762;
  assign n44786 = ~pi92 & ~n44785;
  assign n44787 = ~n44784 & n44786;
  assign n44788 = n6795 & ~n44781;
  assign n44789 = ~n6795 & n44762;
  assign n44790 = pi92 & ~n44789;
  assign n44791 = ~n44788 & n44790;
  assign n44792 = n6792 & ~n44791;
  assign n44793 = ~n44787 & n44792;
  assign n44794 = ~n6792 & n44762;
  assign n44795 = ~pi55 & ~n44794;
  assign n44796 = ~n44793 & n44795;
  assign n44797 = n64082 & n44755;
  assign n44798 = ~n64082 & n44655;
  assign n44799 = pi55 & ~n44798;
  assign n44800 = ~n44797 & n44799;
  assign n44801 = ~pi56 & ~n44800;
  assign n44802 = ~n44796 & n44801;
  assign n44803 = n64084 & ~n44755;
  assign n44804 = ~n64084 & ~n44655;
  assign n44805 = pi56 & ~n44804;
  assign n44806 = ~n64084 & n44655;
  assign n44807 = ~pi55 & n44797;
  assign n44808 = ~n44806 & ~n44807;
  assign n44809 = pi56 & ~n44808;
  assign n44810 = ~n44803 & n44805;
  assign n44811 = ~pi62 & ~n64903;
  assign n44812 = ~n44802 & n44811;
  assign n44813 = n44475 & n44755;
  assign n44814 = ~n44475 & n44655;
  assign n44815 = pi62 & ~n44814;
  assign n44816 = ~n44813 & n44815;
  assign n44817 = ~pi241 & n3472;
  assign n44818 = ~n44816 & n44817;
  assign n44819 = ~n44812 & n44818;
  assign n44820 = pi241 & n44657;
  assign n44821 = ~n3472 & ~n44820;
  assign n44822 = n44655 & n44821;
  assign n44823 = ~n44819 & ~n44822;
  assign n44824 = ~n44723 & ~n44822;
  assign n44825 = ~n44819 & n44824;
  assign n44826 = ~n44723 & n44823;
  assign n44827 = pi223 & pi1140;
  assign n44828 = ~pi299 & ~n44827;
  assign n44829 = ~pi921 & n41469;
  assign n44830 = ~pi1140 & ~n41469;
  assign n44831 = pi222 & ~n44830;
  assign n44832 = pi222 & ~n44829;
  assign n44833 = ~n44830 & n44832;
  assign n44834 = ~n44829 & n44831;
  assign n44835 = pi224 & pi282;
  assign n44836 = ~pi222 & ~n44835;
  assign n44837 = pi869 & n44321;
  assign n44838 = ~pi224 & ~n44837;
  assign n44839 = n44836 & ~n44838;
  assign n44840 = ~n64905 & ~n44839;
  assign n44841 = ~n44321 & n44836;
  assign n44842 = n44840 & ~n44841;
  assign n44843 = ~pi223 & ~n44842;
  assign n44844 = n44828 & ~n44843;
  assign n44845 = ~pi39 & ~n44844;
  assign n44846 = pi215 & pi1140;
  assign n44847 = pi299 & ~n44846;
  assign n44848 = ~pi921 & n41020;
  assign n44849 = ~pi1140 & ~n41020;
  assign n44850 = pi221 & ~n44849;
  assign n44851 = pi221 & ~n44848;
  assign n44852 = ~n44849 & n44851;
  assign n44853 = ~n44848 & n44850;
  assign n44854 = pi216 & pi282;
  assign n44855 = ~pi221 & ~n44854;
  assign n44856 = ~pi869 & n44316;
  assign n44857 = ~pi170 & ~n44856;
  assign n44858 = pi869 & ~n43706;
  assign n44859 = ~pi869 & ~n44327;
  assign n44860 = pi170 & ~n44859;
  assign n44861 = ~n44858 & n44860;
  assign n44862 = ~n44857 & ~n44861;
  assign n44863 = ~pi228 & ~n44862;
  assign n44864 = pi869 & ~n30613;
  assign n44865 = pi105 & ~n44864;
  assign n44866 = ~pi105 & pi170;
  assign n44867 = pi228 & ~n44866;
  assign n44868 = ~n44865 & n44867;
  assign n44869 = ~pi216 & ~n44868;
  assign n44870 = ~n44611 & n44869;
  assign n44871 = ~n44863 & n44870;
  assign n44872 = n44855 & ~n44871;
  assign n44873 = ~n64906 & ~n44872;
  assign n44874 = ~pi215 & ~n44873;
  assign n44875 = n44847 & ~n44874;
  assign n44876 = n44845 & ~n44875;
  assign n44877 = ~pi224 & ~n44864;
  assign n44878 = n44836 & ~n44877;
  assign n44879 = ~n64905 & ~n44878;
  assign n44880 = ~pi223 & ~n44879;
  assign n44881 = ~n44827 & ~n44880;
  assign n44882 = ~pi299 & ~n44881;
  assign n44883 = ~n64897 & ~n44882;
  assign n44884 = ~pi869 & n62380;
  assign n44885 = ~pi228 & ~n44884;
  assign n44886 = ~pi228 & ~n44178;
  assign n44887 = ~n44884 & n44886;
  assign n44888 = ~n44178 & n44885;
  assign n44889 = ~n44384 & n44869;
  assign n44890 = ~n64907 & n44889;
  assign n44891 = n44855 & ~n44890;
  assign n44892 = ~n64906 & ~n44891;
  assign n44893 = ~pi215 & ~n44892;
  assign n44894 = ~n44846 & ~n44893;
  assign n44895 = pi299 & ~n44894;
  assign n44896 = n44883 & ~n44895;
  assign n44897 = pi39 & ~n44896;
  assign n44898 = ~pi38 & ~n44897;
  assign n44899 = ~n44876 & n44898;
  assign n44900 = ~pi170 & ~pi228;
  assign n44901 = n44869 & ~n44900;
  assign n44902 = n44855 & ~n44901;
  assign n44903 = ~n64906 & ~n44902;
  assign n44904 = ~pi215 & ~n44903;
  assign n44905 = ~n44846 & ~n44904;
  assign n44906 = n44656 & ~n44854;
  assign n44907 = n44905 & ~n44906;
  assign n44908 = pi299 & ~n44907;
  assign n44909 = n44883 & ~n44908;
  assign n44910 = pi38 & n44909;
  assign n44911 = ~pi100 & ~n44910;
  assign n44912 = ~n44899 & n44911;
  assign n44913 = pi170 & ~n44422;
  assign n44914 = ~pi869 & n44422;
  assign n44915 = ~pi228 & ~n44914;
  assign n44916 = ~pi228 & ~n44913;
  assign n44917 = ~n44914 & n44916;
  assign n44918 = ~n44913 & n44915;
  assign n44919 = n44889 & ~n64908;
  assign n44920 = n44855 & ~n44919;
  assign n44921 = ~n64906 & ~n44920;
  assign n44922 = ~pi215 & ~n44921;
  assign n44923 = ~n44846 & ~n44922;
  assign n44924 = pi299 & ~n44923;
  assign n44925 = n2764 & n44883;
  assign n44926 = ~n44924 & n44925;
  assign n44927 = ~n2764 & n44909;
  assign n44928 = pi100 & ~n44927;
  assign n44929 = ~n44926 & n44928;
  assign n44930 = ~n44912 & ~n44929;
  assign n44931 = ~pi87 & ~n44930;
  assign n44932 = ~n62373 & n44909;
  assign n44933 = n62373 & n44896;
  assign n44934 = ~n44932 & ~n44933;
  assign n44935 = pi87 & n44934;
  assign n44936 = ~pi75 & ~n44935;
  assign n44937 = ~n44931 & n44936;
  assign n44938 = pi75 & n44909;
  assign n44939 = ~pi92 & ~n44938;
  assign n44940 = ~n44937 & n44939;
  assign n44941 = n6795 & ~n44934;
  assign n44942 = ~n6795 & n44909;
  assign n44943 = pi92 & ~n44942;
  assign n44944 = ~n44941 & n44943;
  assign n44945 = n6792 & ~n44944;
  assign n44946 = ~n44940 & n44945;
  assign n44947 = ~n6792 & n44909;
  assign n44948 = ~pi55 & ~n44947;
  assign n44949 = ~n44946 & n44948;
  assign n44950 = n64082 & n44894;
  assign n44951 = ~n64082 & n44907;
  assign n44952 = pi55 & ~n44951;
  assign n44953 = ~n44950 & n44952;
  assign n44954 = ~pi56 & ~n44953;
  assign n44955 = ~n44949 & n44954;
  assign n44956 = n64084 & ~n44894;
  assign n44957 = ~n64084 & ~n44907;
  assign n44958 = pi56 & ~n44957;
  assign n44959 = ~pi55 & n44950;
  assign n44960 = ~n64084 & n44907;
  assign n44961 = ~n44959 & ~n44960;
  assign n44962 = pi56 & ~n44961;
  assign n44963 = ~n44956 & n44958;
  assign n44964 = ~pi62 & ~n64909;
  assign n44965 = ~n44955 & n44964;
  assign n44966 = n44475 & n44894;
  assign n44967 = ~n44475 & n44907;
  assign n44968 = pi62 & ~n44967;
  assign n44969 = ~n44966 & n44968;
  assign n44970 = pi248 & n3472;
  assign n44971 = ~n44969 & n44970;
  assign n44972 = ~n44965 & n44971;
  assign n44973 = ~pi869 & n43705;
  assign n44974 = ~n33962 & ~n44837;
  assign n44975 = ~n44973 & n44974;
  assign n44976 = pi869 & n44327;
  assign n44977 = ~pi170 & ~n44976;
  assign n44978 = ~pi869 & n43706;
  assign n44979 = n44977 & ~n44978;
  assign n44980 = ~pi170 & ~n44975;
  assign n44981 = pi170 & pi869;
  assign n44982 = n44316 & n44981;
  assign n44983 = pi170 & n44316;
  assign n44984 = ~n44977 & ~n44983;
  assign n44985 = pi869 & ~n44984;
  assign n44986 = ~n43706 & n44977;
  assign n44987 = ~n44985 & ~n44986;
  assign n44988 = ~n64910 & ~n44982;
  assign n44989 = ~pi228 & ~n64911;
  assign n44990 = ~n44337 & n44868;
  assign n44991 = ~pi216 & ~n44990;
  assign n44992 = ~n44989 & n44991;
  assign n44993 = n44855 & ~n44992;
  assign n44994 = ~n64906 & ~n44993;
  assign n44995 = ~pi215 & ~n44994;
  assign n44996 = n44847 & ~n44995;
  assign n44997 = n44828 & n44840;
  assign n44998 = n44845 & ~n44997;
  assign n44999 = ~n44996 & n44998;
  assign n45000 = n44869 & ~n64907;
  assign n45001 = n44855 & ~n45000;
  assign n45002 = ~n64906 & ~n45001;
  assign n45003 = ~pi215 & ~n45002;
  assign n45004 = ~n44846 & ~n45003;
  assign n45005 = pi299 & ~n45004;
  assign n45006 = ~n44882 & ~n45005;
  assign n45007 = pi39 & ~n45006;
  assign n45008 = ~pi38 & ~n45007;
  assign n45009 = ~n44999 & n45008;
  assign n45010 = pi299 & ~n44905;
  assign n45011 = ~n44882 & ~n45010;
  assign n45012 = pi38 & n45011;
  assign n45013 = ~pi100 & ~n45012;
  assign n45014 = ~n45009 & n45013;
  assign n45015 = n44869 & ~n64908;
  assign n45016 = n44855 & ~n45015;
  assign n45017 = ~n64906 & ~n45016;
  assign n45018 = ~pi215 & ~n45017;
  assign n45019 = ~n44846 & ~n45018;
  assign n45020 = pi299 & ~n45019;
  assign n45021 = n2764 & ~n44882;
  assign n45022 = ~n45020 & n45021;
  assign n45023 = ~n2764 & n45011;
  assign n45024 = pi100 & ~n45023;
  assign n45025 = ~n45022 & n45024;
  assign n45026 = ~n45014 & ~n45025;
  assign n45027 = ~pi87 & ~n45026;
  assign n45028 = ~n62373 & n45011;
  assign n45029 = n62373 & n45006;
  assign n45030 = ~n45028 & ~n45029;
  assign n45031 = pi87 & n45030;
  assign n45032 = ~pi75 & ~n45031;
  assign n45033 = ~n45027 & n45032;
  assign n45034 = pi75 & n45011;
  assign n45035 = ~pi92 & ~n45034;
  assign n45036 = ~n45033 & n45035;
  assign n45037 = n6795 & ~n45030;
  assign n45038 = ~n6795 & n45011;
  assign n45039 = pi92 & ~n45038;
  assign n45040 = ~n45037 & n45039;
  assign n45041 = n6792 & ~n45040;
  assign n45042 = ~n45036 & n45041;
  assign n45043 = ~n6792 & n45011;
  assign n45044 = ~pi55 & ~n45043;
  assign n45045 = ~n45042 & n45044;
  assign n45046 = n64082 & n45004;
  assign n45047 = ~n64082 & n44905;
  assign n45048 = pi55 & ~n45047;
  assign n45049 = ~n45046 & n45048;
  assign n45050 = ~pi56 & ~n45049;
  assign n45051 = ~n45045 & n45050;
  assign n45052 = n64084 & ~n45004;
  assign n45053 = ~n64084 & ~n44905;
  assign n45054 = pi56 & ~n45053;
  assign n45055 = ~n64084 & n44905;
  assign n45056 = ~pi55 & n45046;
  assign n45057 = ~n45055 & ~n45056;
  assign n45058 = pi56 & ~n45057;
  assign n45059 = ~n45052 & n45054;
  assign n45060 = ~pi62 & ~n64912;
  assign n45061 = ~n45051 & n45060;
  assign n45062 = n44475 & n45004;
  assign n45063 = ~n44475 & n44905;
  assign n45064 = pi62 & ~n45063;
  assign n45065 = ~n45062 & n45064;
  assign n45066 = ~pi248 & n3472;
  assign n45067 = ~n45065 & n45066;
  assign n45068 = ~n45061 & n45067;
  assign n45069 = pi248 & n44906;
  assign n45070 = ~n3472 & ~n45069;
  assign n45071 = n44905 & n45070;
  assign n45072 = ~n45068 & ~n45071;
  assign n45073 = ~n44972 & ~n45071;
  assign n45074 = ~n45068 & n45073;
  assign n45075 = ~n44972 & n45072;
  assign n45076 = pi216 & ~pi1139;
  assign n45077 = pi833 & pi920;
  assign n45078 = ~pi833 & pi1139;
  assign n45079 = ~pi216 & ~n45078;
  assign n45080 = ~pi216 & ~n45077;
  assign n45081 = ~n45078 & n45080;
  assign n45082 = ~n45077 & n45079;
  assign n45083 = pi221 & ~n64914;
  assign n45084 = ~n45076 & n45083;
  assign n45085 = pi216 & pi281;
  assign n45086 = ~pi221 & ~n45085;
  assign n45087 = ~pi216 & ~pi862;
  assign n45088 = ~n30613 & n41010;
  assign n45089 = ~n34059 & ~n45088;
  assign n45090 = n45087 & ~n45089;
  assign n45091 = n45086 & ~n45090;
  assign n45092 = ~n45084 & ~n45091;
  assign n45093 = ~n44424 & ~n45088;
  assign n45094 = n45086 & n45093;
  assign n45095 = n45092 & ~n45094;
  assign n45096 = pi148 & ~pi215;
  assign n45097 = ~pi216 & ~n45084;
  assign n45098 = ~pi216 & ~n45083;
  assign n45099 = n45093 & n64915;
  assign n45100 = n45096 & ~n45099;
  assign n45101 = ~n45095 & n45100;
  assign n45102 = pi215 & pi1139;
  assign n45103 = ~pi148 & ~pi215;
  assign n45104 = ~n34059 & ~n41010;
  assign n45105 = pi862 & ~n44384;
  assign n45106 = ~pi216 & ~n45105;
  assign n45107 = ~n45104 & n45106;
  assign n45108 = n45086 & ~n45107;
  assign n45109 = ~n45084 & ~n45108;
  assign n45110 = ~n41010 & ~n44424;
  assign n45111 = n45086 & n45110;
  assign n45112 = n45109 & ~n45111;
  assign n45113 = n45103 & ~n45112;
  assign n45114 = ~n45102 & ~n45113;
  assign n45115 = ~n45101 & ~n45102;
  assign n45116 = ~n45113 & n45115;
  assign n45117 = ~n45101 & n45114;
  assign n45118 = pi299 & ~n64916;
  assign n45119 = ~pi920 & n41469;
  assign n45120 = ~pi1139 & ~n41469;
  assign n45121 = pi222 & ~n45120;
  assign n45122 = pi222 & ~n45119;
  assign n45123 = ~n45120 & n45122;
  assign n45124 = ~n45119 & n45121;
  assign n45125 = pi223 & pi1139;
  assign n45126 = ~pi224 & ~n45125;
  assign n45127 = ~n64917 & n45126;
  assign n45128 = n30613 & n45127;
  assign n45129 = ~pi862 & n45127;
  assign n45130 = pi224 & pi281;
  assign n45131 = ~pi222 & ~n45130;
  assign n45132 = ~n64917 & ~n45131;
  assign n45133 = ~pi223 & ~n45132;
  assign n45134 = ~n45125 & ~n45133;
  assign n45135 = ~pi299 & ~n45134;
  assign n45136 = ~n45129 & n45135;
  assign n45137 = ~n45128 & n45136;
  assign n45138 = n2764 & ~n45137;
  assign n45139 = ~n45118 & n45138;
  assign n45140 = n45087 & n45088;
  assign n45141 = n45086 & ~n45140;
  assign n45142 = ~n45084 & ~n45141;
  assign n45143 = pi148 & ~n41010;
  assign n45144 = n64915 & n45143;
  assign n45145 = ~pi215 & ~n45144;
  assign n45146 = ~n45142 & n45145;
  assign n45147 = ~n45102 & ~n45146;
  assign n45148 = ~n44399 & ~n45147;
  assign n45149 = pi299 & n45148;
  assign n45150 = ~n45137 & ~n45149;
  assign n45151 = ~n2764 & n45150;
  assign n45152 = pi100 & ~n45151;
  assign n45153 = ~n45139 & n45152;
  assign n45154 = ~pi228 & n43706;
  assign n45155 = ~n41010 & ~n45154;
  assign n45156 = ~pi862 & n45155;
  assign n45157 = pi228 & ~n44337;
  assign n45158 = ~pi228 & ~n44327;
  assign n45159 = ~n45157 & ~n45158;
  assign n45160 = pi862 & ~n45159;
  assign n45161 = ~pi216 & ~n45160;
  assign n45162 = ~n45156 & n45161;
  assign n45163 = n45086 & ~n45162;
  assign n45164 = ~n45084 & ~n45163;
  assign n45165 = n45103 & ~n45164;
  assign n45166 = ~pi228 & n44316;
  assign n45167 = n41010 & n44321;
  assign n45168 = ~n45166 & ~n45167;
  assign n45169 = n45087 & ~n45168;
  assign n45170 = n45086 & ~n45169;
  assign n45171 = ~n45084 & ~n45170;
  assign n45172 = n64915 & n45168;
  assign n45173 = n45096 & ~n45172;
  assign n45174 = ~n45171 & n45173;
  assign n45175 = pi299 & ~n45102;
  assign n45176 = ~n45174 & n45175;
  assign n45177 = ~n45165 & n45176;
  assign n45178 = ~n44321 & n45127;
  assign n45179 = ~n45129 & ~n45134;
  assign n45180 = ~n45178 & n45179;
  assign n45181 = ~pi299 & ~n45180;
  assign n45182 = ~pi39 & ~n45181;
  assign n45183 = ~n45177 & n45182;
  assign n45184 = n45103 & ~n45109;
  assign n45185 = n45089 & n64915;
  assign n45186 = n45096 & ~n45185;
  assign n45187 = ~n45092 & n45096;
  assign n45188 = ~n45185 & n45187;
  assign n45189 = ~n45092 & n45186;
  assign n45190 = ~n45102 & ~n64918;
  assign n45191 = ~n45184 & n45190;
  assign n45192 = pi299 & ~n45191;
  assign n45193 = ~n45137 & ~n45192;
  assign n45194 = pi39 & ~n45193;
  assign n45195 = ~pi38 & ~n45194;
  assign n45196 = ~n45183 & n45195;
  assign n45197 = pi38 & n45150;
  assign n45198 = ~pi100 & ~n45197;
  assign n45199 = ~n45196 & n45198;
  assign n45200 = ~n45153 & ~n45199;
  assign n45201 = ~pi87 & ~n45200;
  assign n45202 = ~n62373 & n45150;
  assign n45203 = n62373 & n45193;
  assign n45204 = ~n45202 & ~n45203;
  assign n45205 = pi87 & n45204;
  assign n45206 = ~pi75 & ~n45205;
  assign n45207 = ~n45201 & n45206;
  assign n45208 = pi75 & n45150;
  assign n45209 = ~pi92 & ~n45208;
  assign n45210 = ~n45207 & n45209;
  assign n45211 = n6795 & ~n45204;
  assign n45212 = ~n6795 & n45150;
  assign n45213 = pi92 & ~n45212;
  assign n45214 = ~n45211 & n45213;
  assign n45215 = n6792 & ~n45214;
  assign n45216 = ~n45210 & n45215;
  assign n45217 = ~n6792 & n45150;
  assign n45218 = ~pi55 & ~n45217;
  assign n45219 = ~n45216 & n45218;
  assign n45220 = n64082 & n45191;
  assign n45221 = ~n64082 & ~n45148;
  assign n45222 = pi55 & ~n45221;
  assign n45223 = ~n45220 & n45222;
  assign n45224 = ~pi56 & ~n45223;
  assign n45225 = ~n45219 & n45224;
  assign n45226 = n64084 & ~n45191;
  assign n45227 = ~n64084 & n45148;
  assign n45228 = pi56 & ~n45227;
  assign n45229 = ~n64084 & ~n45148;
  assign n45230 = ~pi55 & n45220;
  assign n45231 = ~n45229 & ~n45230;
  assign n45232 = pi56 & ~n45231;
  assign n45233 = ~n45226 & n45228;
  assign n45234 = ~pi62 & ~n64919;
  assign n45235 = ~n45225 & n45234;
  assign n45236 = n44475 & n45191;
  assign n45237 = ~n44475 & ~n45148;
  assign n45238 = pi62 & ~n45237;
  assign n45239 = ~n45236 & n45238;
  assign n45240 = n3472 & ~n45239;
  assign n45241 = ~n45235 & n45240;
  assign n45242 = ~n3472 & ~n45148;
  assign n45243 = ~pi247 & ~n45242;
  assign n45244 = ~n45241 & n45243;
  assign n45245 = ~n45095 & n45103;
  assign n45246 = n64915 & n45110;
  assign n45247 = n45187 & ~n45246;
  assign n45248 = ~n45102 & ~n45247;
  assign n45249 = ~n45245 & n45248;
  assign n45250 = pi299 & ~n45249;
  assign n45251 = ~n64897 & ~n45136;
  assign n45252 = n2764 & n45251;
  assign n45253 = ~n45250 & n45252;
  assign n45254 = pi299 & ~n45147;
  assign n45255 = n45251 & ~n45254;
  assign n45256 = ~n2764 & n45255;
  assign n45257 = pi100 & ~n45256;
  assign n45258 = ~n45253 & n45257;
  assign n45259 = n44321 & n45129;
  assign n45260 = n45135 & ~n45259;
  assign n45261 = pi862 & ~n45155;
  assign n45262 = ~pi862 & n45159;
  assign n45263 = ~pi216 & ~n45262;
  assign n45264 = ~n45261 & n45263;
  assign n45265 = n45086 & ~n45264;
  assign n45266 = ~n45084 & ~n45265;
  assign n45267 = n45096 & ~n45266;
  assign n45268 = n45103 & ~n45171;
  assign n45269 = ~n45102 & ~n45268;
  assign n45270 = ~n45267 & n45269;
  assign n45271 = pi299 & ~n45270;
  assign n45272 = ~n45260 & ~n45271;
  assign n45273 = ~pi39 & ~n45272;
  assign n45274 = ~n45092 & n45145;
  assign n45275 = n45190 & ~n45274;
  assign n45276 = pi299 & ~n45275;
  assign n45277 = n45251 & ~n45276;
  assign n45278 = pi39 & ~n45277;
  assign n45279 = ~pi38 & ~n45278;
  assign n45280 = ~n45273 & n45279;
  assign n45281 = pi38 & n45255;
  assign n45282 = ~pi100 & ~n45281;
  assign n45283 = ~n45280 & n45282;
  assign n45284 = ~n45258 & ~n45283;
  assign n45285 = ~pi87 & ~n45284;
  assign n45286 = ~n62373 & n45255;
  assign n45287 = n62373 & n45277;
  assign n45288 = ~n45286 & ~n45287;
  assign n45289 = pi87 & n45288;
  assign n45290 = ~pi75 & ~n45289;
  assign n45291 = ~n45285 & n45290;
  assign n45292 = pi75 & n45255;
  assign n45293 = ~pi92 & ~n45292;
  assign n45294 = ~n45291 & n45293;
  assign n45295 = n6795 & ~n45288;
  assign n45296 = ~n6795 & n45255;
  assign n45297 = pi92 & ~n45296;
  assign n45298 = ~n45295 & n45297;
  assign n45299 = n6792 & ~n45298;
  assign n45300 = ~n45294 & n45299;
  assign n45301 = ~n6792 & n45255;
  assign n45302 = ~pi55 & ~n45301;
  assign n45303 = ~n45300 & n45302;
  assign n45304 = n64082 & n45275;
  assign n45305 = ~n64082 & n45147;
  assign n45306 = pi55 & ~n45305;
  assign n45307 = ~n45304 & n45306;
  assign n45308 = ~pi56 & ~n45307;
  assign n45309 = ~n45303 & n45308;
  assign n45310 = n64084 & ~n45275;
  assign n45311 = ~n64084 & ~n45147;
  assign n45312 = pi56 & ~n45311;
  assign n45313 = ~n64084 & n45147;
  assign n45314 = ~pi55 & n45304;
  assign n45315 = ~n45313 & ~n45314;
  assign n45316 = pi56 & ~n45315;
  assign n45317 = ~n45310 & n45312;
  assign n45318 = ~pi62 & ~n64920;
  assign n45319 = ~n45309 & n45318;
  assign n45320 = n44475 & n45275;
  assign n45321 = ~n44475 & n45147;
  assign n45322 = pi62 & ~n45321;
  assign n45323 = ~n45320 & n45322;
  assign n45324 = n3472 & ~n45323;
  assign n45325 = ~n45319 & n45324;
  assign n45326 = ~n3472 & n45147;
  assign n45327 = pi247 & ~n45326;
  assign n45328 = ~n45325 & n45327;
  assign n45329 = ~n45244 & ~n45328;
  assign n45330 = pi223 & pi1138;
  assign n45331 = ~pi299 & ~n45330;
  assign n45332 = ~pi940 & n41469;
  assign n45333 = ~pi1138 & ~n41469;
  assign n45334 = pi222 & ~n45333;
  assign n45335 = pi222 & ~n45332;
  assign n45336 = ~n45333 & n45335;
  assign n45337 = ~n45332 & n45334;
  assign n45338 = pi224 & pi269;
  assign n45339 = ~pi222 & ~n45338;
  assign n45340 = pi877 & n44321;
  assign n45341 = ~pi224 & ~n45340;
  assign n45342 = n45339 & ~n45341;
  assign n45343 = ~n64921 & ~n45342;
  assign n45344 = ~n44321 & n45339;
  assign n45345 = n45343 & ~n45344;
  assign n45346 = ~pi223 & ~n45345;
  assign n45347 = n45331 & ~n45346;
  assign n45348 = ~pi39 & ~n45347;
  assign n45349 = pi215 & pi1138;
  assign n45350 = pi299 & ~n45349;
  assign n45351 = ~pi940 & n41020;
  assign n45352 = ~pi1138 & ~n41020;
  assign n45353 = pi221 & ~n45352;
  assign n45354 = pi221 & ~n45351;
  assign n45355 = ~n45352 & n45354;
  assign n45356 = ~n45351 & n45353;
  assign n45357 = pi216 & pi269;
  assign n45358 = ~pi221 & ~n45357;
  assign n45359 = ~pi877 & n44316;
  assign n45360 = ~pi169 & ~n45359;
  assign n45361 = pi877 & ~n43706;
  assign n45362 = ~pi877 & ~n44327;
  assign n45363 = pi169 & ~n45362;
  assign n45364 = ~n45361 & n45363;
  assign n45365 = ~n45360 & ~n45364;
  assign n45366 = ~pi228 & ~n45365;
  assign n45367 = pi877 & ~n30613;
  assign n45368 = pi105 & ~n45367;
  assign n45369 = ~pi105 & pi169;
  assign n45370 = pi228 & ~n45369;
  assign n45371 = ~n45368 & n45370;
  assign n45372 = ~pi216 & ~n45371;
  assign n45373 = ~n44611 & n45372;
  assign n45374 = ~n45366 & n45373;
  assign n45375 = n45358 & ~n45374;
  assign n45376 = ~n64922 & ~n45375;
  assign n45377 = ~pi215 & ~n45376;
  assign n45378 = n45350 & ~n45377;
  assign n45379 = n45348 & ~n45378;
  assign n45380 = ~pi224 & ~n45367;
  assign n45381 = n45339 & ~n45380;
  assign n45382 = ~n64921 & ~n45381;
  assign n45383 = ~pi223 & ~n45382;
  assign n45384 = ~n45330 & ~n45383;
  assign n45385 = ~pi299 & ~n45384;
  assign n45386 = ~n64897 & ~n45385;
  assign n45387 = pi169 & ~n62380;
  assign n45388 = ~pi877 & n62380;
  assign n45389 = ~pi228 & ~n45388;
  assign n45390 = ~pi228 & ~n45387;
  assign n45391 = ~n45388 & n45390;
  assign n45392 = ~n45387 & n45389;
  assign n45393 = ~n44384 & n45372;
  assign n45394 = ~n64923 & n45393;
  assign n45395 = n45358 & ~n45394;
  assign n45396 = ~n64922 & ~n45395;
  assign n45397 = ~pi215 & ~n45396;
  assign n45398 = ~n45349 & ~n45397;
  assign n45399 = pi299 & ~n45398;
  assign n45400 = n45386 & ~n45399;
  assign n45401 = pi39 & ~n45400;
  assign n45402 = ~pi38 & ~n45401;
  assign n45403 = ~n45379 & n45402;
  assign n45404 = ~pi169 & ~pi228;
  assign n45405 = n45372 & ~n45404;
  assign n45406 = n45358 & ~n45405;
  assign n45407 = ~n64922 & ~n45406;
  assign n45408 = ~pi215 & ~n45407;
  assign n45409 = ~n45349 & ~n45408;
  assign n45410 = n44656 & ~n45357;
  assign n45411 = n45409 & ~n45410;
  assign n45412 = pi299 & ~n45411;
  assign n45413 = n45386 & ~n45412;
  assign n45414 = pi38 & n45413;
  assign n45415 = ~pi100 & ~n45414;
  assign n45416 = ~n45403 & n45415;
  assign n45417 = pi169 & ~n44422;
  assign n45418 = ~pi877 & n44422;
  assign n45419 = ~pi228 & ~n45418;
  assign n45420 = ~pi228 & ~n45417;
  assign n45421 = ~n45418 & n45420;
  assign n45422 = ~n45417 & n45419;
  assign n45423 = n45393 & ~n64924;
  assign n45424 = n45358 & ~n45423;
  assign n45425 = ~n64922 & ~n45424;
  assign n45426 = ~pi215 & ~n45425;
  assign n45427 = ~n45349 & ~n45426;
  assign n45428 = pi299 & ~n45427;
  assign n45429 = n2764 & n45386;
  assign n45430 = ~n45428 & n45429;
  assign n45431 = ~n2764 & n45413;
  assign n45432 = pi100 & ~n45431;
  assign n45433 = ~n45430 & n45432;
  assign n45434 = ~n45416 & ~n45433;
  assign n45435 = ~pi87 & ~n45434;
  assign n45436 = ~n62373 & n45413;
  assign n45437 = n62373 & n45400;
  assign n45438 = ~n45436 & ~n45437;
  assign n45439 = pi87 & n45438;
  assign n45440 = ~pi75 & ~n45439;
  assign n45441 = ~n45435 & n45440;
  assign n45442 = pi75 & n45413;
  assign n45443 = ~pi92 & ~n45442;
  assign n45444 = ~n45441 & n45443;
  assign n45445 = n6795 & ~n45438;
  assign n45446 = ~n6795 & n45413;
  assign n45447 = pi92 & ~n45446;
  assign n45448 = ~n45445 & n45447;
  assign n45449 = n6792 & ~n45448;
  assign n45450 = ~n45444 & n45449;
  assign n45451 = ~n6792 & n45413;
  assign n45452 = ~pi55 & ~n45451;
  assign n45453 = ~n45450 & n45452;
  assign n45454 = n64082 & n45398;
  assign n45455 = ~n64082 & n45411;
  assign n45456 = pi55 & ~n45455;
  assign n45457 = ~n45454 & n45456;
  assign n45458 = ~pi56 & ~n45457;
  assign n45459 = ~n45453 & n45458;
  assign n45460 = n64084 & ~n45398;
  assign n45461 = ~n64084 & ~n45411;
  assign n45462 = pi56 & ~n45461;
  assign n45463 = ~pi55 & n45454;
  assign n45464 = ~n64084 & n45411;
  assign n45465 = ~n45463 & ~n45464;
  assign n45466 = pi56 & ~n45465;
  assign n45467 = ~n45460 & n45462;
  assign n45468 = ~pi62 & ~n64925;
  assign n45469 = ~n45459 & n45468;
  assign n45470 = n44475 & n45398;
  assign n45471 = ~n44475 & n45411;
  assign n45472 = pi62 & ~n45471;
  assign n45473 = ~n45470 & n45472;
  assign n45474 = pi246 & n3472;
  assign n45475 = ~n45473 & n45474;
  assign n45476 = ~n45469 & n45475;
  assign n45477 = ~pi877 & n43705;
  assign n45478 = ~n33962 & ~n45340;
  assign n45479 = ~n45477 & n45478;
  assign n45480 = pi877 & n44327;
  assign n45481 = ~pi169 & ~n45480;
  assign n45482 = ~pi877 & n43706;
  assign n45483 = n45481 & ~n45482;
  assign n45484 = ~pi169 & ~n45479;
  assign n45485 = pi169 & pi877;
  assign n45486 = n44316 & n45485;
  assign n45487 = pi169 & n44316;
  assign n45488 = ~n45481 & ~n45487;
  assign n45489 = pi877 & ~n45488;
  assign n45490 = ~n43706 & n45481;
  assign n45491 = ~n45489 & ~n45490;
  assign n45492 = ~n64926 & ~n45486;
  assign n45493 = ~pi228 & ~n64927;
  assign n45494 = ~n44337 & n45371;
  assign n45495 = ~pi216 & ~n45494;
  assign n45496 = ~n45493 & n45495;
  assign n45497 = n45358 & ~n45496;
  assign n45498 = ~n64922 & ~n45497;
  assign n45499 = ~pi215 & ~n45498;
  assign n45500 = n45350 & ~n45499;
  assign n45501 = n45331 & n45343;
  assign n45502 = n45348 & ~n45501;
  assign n45503 = ~n45500 & n45502;
  assign n45504 = n45372 & ~n64923;
  assign n45505 = n45358 & ~n45504;
  assign n45506 = ~n64922 & ~n45505;
  assign n45507 = ~pi215 & ~n45506;
  assign n45508 = ~n45349 & ~n45507;
  assign n45509 = pi299 & ~n45508;
  assign n45510 = ~n45385 & ~n45509;
  assign n45511 = pi39 & ~n45510;
  assign n45512 = ~pi38 & ~n45511;
  assign n45513 = ~n45503 & n45512;
  assign n45514 = pi299 & ~n45409;
  assign n45515 = ~n45385 & ~n45514;
  assign n45516 = pi38 & n45515;
  assign n45517 = ~pi100 & ~n45516;
  assign n45518 = ~n45513 & n45517;
  assign n45519 = n45372 & ~n64924;
  assign n45520 = n45358 & ~n45519;
  assign n45521 = ~n64922 & ~n45520;
  assign n45522 = ~pi215 & ~n45521;
  assign n45523 = ~n45349 & ~n45522;
  assign n45524 = pi299 & ~n45523;
  assign n45525 = n2764 & ~n45385;
  assign n45526 = ~n45524 & n45525;
  assign n45527 = ~n2764 & n45515;
  assign n45528 = pi100 & ~n45527;
  assign n45529 = ~n45526 & n45528;
  assign n45530 = ~n45518 & ~n45529;
  assign n45531 = ~pi87 & ~n45530;
  assign n45532 = ~n62373 & n45515;
  assign n45533 = n62373 & n45510;
  assign n45534 = ~n45532 & ~n45533;
  assign n45535 = pi87 & n45534;
  assign n45536 = ~pi75 & ~n45535;
  assign n45537 = ~n45531 & n45536;
  assign n45538 = pi75 & n45515;
  assign n45539 = ~pi92 & ~n45538;
  assign n45540 = ~n45537 & n45539;
  assign n45541 = n6795 & ~n45534;
  assign n45542 = ~n6795 & n45515;
  assign n45543 = pi92 & ~n45542;
  assign n45544 = ~n45541 & n45543;
  assign n45545 = n6792 & ~n45544;
  assign n45546 = ~n45540 & n45545;
  assign n45547 = ~n6792 & n45515;
  assign n45548 = ~pi55 & ~n45547;
  assign n45549 = ~n45546 & n45548;
  assign n45550 = n64082 & n45508;
  assign n45551 = ~n64082 & n45409;
  assign n45552 = pi55 & ~n45551;
  assign n45553 = ~n45550 & n45552;
  assign n45554 = ~pi56 & ~n45553;
  assign n45555 = ~n45549 & n45554;
  assign n45556 = n64084 & ~n45508;
  assign n45557 = ~n64084 & ~n45409;
  assign n45558 = pi56 & ~n45557;
  assign n45559 = ~n64084 & n45409;
  assign n45560 = ~pi55 & n45550;
  assign n45561 = ~n45559 & ~n45560;
  assign n45562 = pi56 & ~n45561;
  assign n45563 = ~n45556 & n45558;
  assign n45564 = ~pi62 & ~n64928;
  assign n45565 = ~n45555 & n45564;
  assign n45566 = n44475 & n45508;
  assign n45567 = ~n44475 & n45409;
  assign n45568 = pi62 & ~n45567;
  assign n45569 = ~n45566 & n45568;
  assign n45570 = ~pi246 & n3472;
  assign n45571 = ~n45569 & n45570;
  assign n45572 = ~n45565 & n45571;
  assign n45573 = pi246 & n45410;
  assign n45574 = ~n3472 & ~n45573;
  assign n45575 = n45409 & n45574;
  assign n45576 = ~n45572 & ~n45575;
  assign n45577 = ~n45476 & ~n45575;
  assign n45578 = ~n45572 & n45577;
  assign n45579 = ~n45476 & n45576;
  assign n45580 = pi223 & pi1137;
  assign n45581 = ~pi299 & ~n45580;
  assign n45582 = ~pi933 & n41469;
  assign n45583 = ~pi1137 & ~n41469;
  assign n45584 = pi222 & ~n45583;
  assign n45585 = pi222 & ~n45582;
  assign n45586 = ~n45583 & n45585;
  assign n45587 = ~n45582 & n45584;
  assign n45588 = pi224 & pi280;
  assign n45589 = ~pi222 & ~n45588;
  assign n45590 = pi878 & n44321;
  assign n45591 = ~pi224 & ~n45590;
  assign n45592 = n45589 & ~n45591;
  assign n45593 = ~n64930 & ~n45592;
  assign n45594 = ~n44321 & n45589;
  assign n45595 = n45593 & ~n45594;
  assign n45596 = ~pi223 & ~n45595;
  assign n45597 = n45581 & ~n45596;
  assign n45598 = ~pi39 & ~n45597;
  assign n45599 = pi215 & pi1137;
  assign n45600 = pi299 & ~n45599;
  assign n45601 = ~pi933 & n41020;
  assign n45602 = ~pi1137 & ~n41020;
  assign n45603 = pi221 & ~n45602;
  assign n45604 = pi221 & ~n45601;
  assign n45605 = ~n45602 & n45604;
  assign n45606 = ~n45601 & n45603;
  assign n45607 = pi216 & pi280;
  assign n45608 = ~pi221 & ~n45607;
  assign n45609 = ~pi878 & n44316;
  assign n45610 = ~pi168 & ~n45609;
  assign n45611 = pi878 & ~n43706;
  assign n45612 = ~pi878 & ~n44327;
  assign n45613 = pi168 & ~n45612;
  assign n45614 = ~n45611 & n45613;
  assign n45615 = ~n45610 & ~n45614;
  assign n45616 = ~pi228 & ~n45615;
  assign n45617 = pi878 & ~n30613;
  assign n45618 = pi105 & ~n45617;
  assign n45619 = ~pi105 & pi168;
  assign n45620 = pi228 & ~n45619;
  assign n45621 = ~n45618 & n45620;
  assign n45622 = ~pi216 & ~n45621;
  assign n45623 = ~n44611 & n45622;
  assign n45624 = ~n45616 & n45623;
  assign n45625 = n45608 & ~n45624;
  assign n45626 = ~n64931 & ~n45625;
  assign n45627 = ~pi215 & ~n45626;
  assign n45628 = n45600 & ~n45627;
  assign n45629 = n45598 & ~n45628;
  assign n45630 = ~pi224 & ~n45617;
  assign n45631 = n45589 & ~n45630;
  assign n45632 = ~n64930 & ~n45631;
  assign n45633 = ~pi223 & ~n45632;
  assign n45634 = ~n45580 & ~n45633;
  assign n45635 = ~pi299 & ~n45634;
  assign n45636 = ~n64897 & ~n45635;
  assign n45637 = pi168 & ~n62380;
  assign n45638 = ~pi878 & n62380;
  assign n45639 = ~pi228 & ~n45638;
  assign n45640 = ~pi228 & ~n45637;
  assign n45641 = ~n45638 & n45640;
  assign n45642 = ~n45637 & n45639;
  assign n45643 = ~n44384 & n45622;
  assign n45644 = ~n64932 & n45643;
  assign n45645 = n45608 & ~n45644;
  assign n45646 = ~n64931 & ~n45645;
  assign n45647 = ~pi215 & ~n45646;
  assign n45648 = ~n45599 & ~n45647;
  assign n45649 = pi299 & ~n45648;
  assign n45650 = n45636 & ~n45649;
  assign n45651 = pi39 & ~n45650;
  assign n45652 = ~pi38 & ~n45651;
  assign n45653 = ~n45629 & n45652;
  assign n45654 = ~pi168 & ~pi228;
  assign n45655 = n45622 & ~n45654;
  assign n45656 = n45608 & ~n45655;
  assign n45657 = ~n64931 & ~n45656;
  assign n45658 = ~pi215 & ~n45657;
  assign n45659 = ~n45599 & ~n45658;
  assign n45660 = n44656 & ~n45607;
  assign n45661 = n45659 & ~n45660;
  assign n45662 = pi299 & ~n45661;
  assign n45663 = n45636 & ~n45662;
  assign n45664 = pi38 & n45663;
  assign n45665 = ~pi100 & ~n45664;
  assign n45666 = ~n45653 & n45665;
  assign n45667 = pi168 & ~n44422;
  assign n45668 = ~pi878 & n44422;
  assign n45669 = ~pi228 & ~n45668;
  assign n45670 = ~pi228 & ~n45667;
  assign n45671 = ~n45668 & n45670;
  assign n45672 = ~n45667 & n45669;
  assign n45673 = n45643 & ~n64933;
  assign n45674 = n45608 & ~n45673;
  assign n45675 = ~n64931 & ~n45674;
  assign n45676 = ~pi215 & ~n45675;
  assign n45677 = ~n45599 & ~n45676;
  assign n45678 = pi299 & ~n45677;
  assign n45679 = n2764 & n45636;
  assign n45680 = ~n45678 & n45679;
  assign n45681 = ~n2764 & n45663;
  assign n45682 = pi100 & ~n45681;
  assign n45683 = ~n45680 & n45682;
  assign n45684 = ~n45666 & ~n45683;
  assign n45685 = ~pi87 & ~n45684;
  assign n45686 = ~n62373 & n45663;
  assign n45687 = n62373 & n45650;
  assign n45688 = ~n45686 & ~n45687;
  assign n45689 = pi87 & n45688;
  assign n45690 = ~pi75 & ~n45689;
  assign n45691 = ~n45685 & n45690;
  assign n45692 = pi75 & n45663;
  assign n45693 = ~pi92 & ~n45692;
  assign n45694 = ~n45691 & n45693;
  assign n45695 = n6795 & ~n45688;
  assign n45696 = ~n6795 & n45663;
  assign n45697 = pi92 & ~n45696;
  assign n45698 = ~n45695 & n45697;
  assign n45699 = n6792 & ~n45698;
  assign n45700 = ~n45694 & n45699;
  assign n45701 = ~n6792 & n45663;
  assign n45702 = ~pi55 & ~n45701;
  assign n45703 = ~n45700 & n45702;
  assign n45704 = n64082 & n45648;
  assign n45705 = ~n64082 & n45661;
  assign n45706 = pi55 & ~n45705;
  assign n45707 = ~n45704 & n45706;
  assign n45708 = ~pi56 & ~n45707;
  assign n45709 = ~n45703 & n45708;
  assign n45710 = n64084 & ~n45648;
  assign n45711 = ~n64084 & ~n45661;
  assign n45712 = pi56 & ~n45711;
  assign n45713 = ~pi55 & n45704;
  assign n45714 = ~n64084 & n45661;
  assign n45715 = ~n45713 & ~n45714;
  assign n45716 = pi56 & ~n45715;
  assign n45717 = ~n45710 & n45712;
  assign n45718 = ~pi62 & ~n64934;
  assign n45719 = ~n45709 & n45718;
  assign n45720 = n44475 & n45648;
  assign n45721 = ~n44475 & n45661;
  assign n45722 = pi62 & ~n45721;
  assign n45723 = ~n45720 & n45722;
  assign n45724 = pi240 & n3472;
  assign n45725 = ~n45723 & n45724;
  assign n45726 = ~n45719 & n45725;
  assign n45727 = ~pi878 & n43705;
  assign n45728 = ~n33962 & ~n45590;
  assign n45729 = ~n45727 & n45728;
  assign n45730 = pi878 & n44327;
  assign n45731 = ~pi168 & ~n45730;
  assign n45732 = ~pi878 & n43706;
  assign n45733 = n45731 & ~n45732;
  assign n45734 = ~pi168 & ~n45729;
  assign n45735 = pi168 & pi878;
  assign n45736 = n44316 & n45735;
  assign n45737 = pi168 & n44316;
  assign n45738 = ~n45731 & ~n45737;
  assign n45739 = pi878 & ~n45738;
  assign n45740 = ~n43706 & n45731;
  assign n45741 = ~n45739 & ~n45740;
  assign n45742 = ~n64935 & ~n45736;
  assign n45743 = ~pi228 & ~n64936;
  assign n45744 = ~n44337 & n45621;
  assign n45745 = ~pi216 & ~n45744;
  assign n45746 = ~n45743 & n45745;
  assign n45747 = n45608 & ~n45746;
  assign n45748 = ~n64931 & ~n45747;
  assign n45749 = ~pi215 & ~n45748;
  assign n45750 = n45600 & ~n45749;
  assign n45751 = n45581 & n45593;
  assign n45752 = n45598 & ~n45751;
  assign n45753 = ~n45750 & n45752;
  assign n45754 = n45622 & ~n64932;
  assign n45755 = n45608 & ~n45754;
  assign n45756 = ~n64931 & ~n45755;
  assign n45757 = ~pi215 & ~n45756;
  assign n45758 = ~n45599 & ~n45757;
  assign n45759 = pi299 & ~n45758;
  assign n45760 = ~n45635 & ~n45759;
  assign n45761 = pi39 & ~n45760;
  assign n45762 = ~pi38 & ~n45761;
  assign n45763 = ~n45753 & n45762;
  assign n45764 = pi299 & ~n45659;
  assign n45765 = ~n45635 & ~n45764;
  assign n45766 = pi38 & n45765;
  assign n45767 = ~pi100 & ~n45766;
  assign n45768 = ~n45763 & n45767;
  assign n45769 = n45622 & ~n64933;
  assign n45770 = n45608 & ~n45769;
  assign n45771 = ~n64931 & ~n45770;
  assign n45772 = ~pi215 & ~n45771;
  assign n45773 = ~n45599 & ~n45772;
  assign n45774 = pi299 & ~n45773;
  assign n45775 = n2764 & ~n45635;
  assign n45776 = ~n45774 & n45775;
  assign n45777 = ~n2764 & n45765;
  assign n45778 = pi100 & ~n45777;
  assign n45779 = ~n45776 & n45778;
  assign n45780 = ~n45768 & ~n45779;
  assign n45781 = ~pi87 & ~n45780;
  assign n45782 = ~n62373 & n45765;
  assign n45783 = n62373 & n45760;
  assign n45784 = ~n45782 & ~n45783;
  assign n45785 = pi87 & n45784;
  assign n45786 = ~pi75 & ~n45785;
  assign n45787 = ~n45781 & n45786;
  assign n45788 = pi75 & n45765;
  assign n45789 = ~pi92 & ~n45788;
  assign n45790 = ~n45787 & n45789;
  assign n45791 = n6795 & ~n45784;
  assign n45792 = ~n6795 & n45765;
  assign n45793 = pi92 & ~n45792;
  assign n45794 = ~n45791 & n45793;
  assign n45795 = n6792 & ~n45794;
  assign n45796 = ~n45790 & n45795;
  assign n45797 = ~n6792 & n45765;
  assign n45798 = ~pi55 & ~n45797;
  assign n45799 = ~n45796 & n45798;
  assign n45800 = n64082 & n45758;
  assign n45801 = ~n64082 & n45659;
  assign n45802 = pi55 & ~n45801;
  assign n45803 = ~n45800 & n45802;
  assign n45804 = ~pi56 & ~n45803;
  assign n45805 = ~n45799 & n45804;
  assign n45806 = n64084 & ~n45758;
  assign n45807 = ~n64084 & ~n45659;
  assign n45808 = pi56 & ~n45807;
  assign n45809 = ~n64084 & n45659;
  assign n45810 = ~pi55 & n45800;
  assign n45811 = ~n45809 & ~n45810;
  assign n45812 = pi56 & ~n45811;
  assign n45813 = ~n45806 & n45808;
  assign n45814 = ~pi62 & ~n64937;
  assign n45815 = ~n45805 & n45814;
  assign n45816 = n44475 & n45758;
  assign n45817 = ~n44475 & n45659;
  assign n45818 = pi62 & ~n45817;
  assign n45819 = ~n45816 & n45818;
  assign n45820 = ~pi240 & n3472;
  assign n45821 = ~n45819 & n45820;
  assign n45822 = ~n45815 & n45821;
  assign n45823 = pi240 & n45660;
  assign n45824 = ~n3472 & ~n45823;
  assign n45825 = n45659 & n45824;
  assign n45826 = ~n45822 & ~n45825;
  assign n45827 = ~n45726 & ~n45825;
  assign n45828 = ~n45822 & n45827;
  assign n45829 = ~n45726 & n45826;
  assign n45830 = ~n64105 & n64148;
  assign n45831 = ~pi137 & ~n45830;
  assign n45832 = n30856 & ~n45831;
  assign n45833 = n33868 & ~n38180;
  assign n45834 = ~n41080 & n45833;
  assign n45835 = n33860 & ~n45834;
  assign n45836 = n33859 & ~n45835;
  assign n45837 = ~n41054 & ~n45836;
  assign n45838 = ~pi95 & ~n45837;
  assign n45839 = ~n33962 & ~n45838;
  assign n45840 = pi137 & ~n45839;
  assign n45841 = ~n64518 & n41097;
  assign n45842 = n41098 & ~n45841;
  assign n45843 = ~pi137 & ~n45842;
  assign n45844 = ~n45840 & ~n45843;
  assign n45845 = pi332 & ~n45844;
  assign n45846 = ~n33962 & ~n41134;
  assign n45847 = pi137 & ~n45846;
  assign n45848 = ~n41100 & ~n45847;
  assign n45849 = ~pi332 & ~n45848;
  assign n45850 = ~n45845 & ~n45849;
  assign n45851 = n30860 & n45850;
  assign n45852 = pi1093 & ~n45842;
  assign n45853 = n2883 & n41098;
  assign n45854 = n2748 & ~n41139;
  assign n45855 = ~pi32 & ~n45854;
  assign n45856 = n45853 & ~n45855;
  assign n45857 = ~pi1093 & ~n45856;
  assign n45858 = ~n2883 & n45842;
  assign n45859 = n64518 & n45853;
  assign n45860 = ~n45858 & ~n45859;
  assign n45861 = n45857 & n45860;
  assign n45862 = ~n45852 & ~n45861;
  assign n45863 = n40634 & ~n45862;
  assign n45864 = ~n2883 & n41099;
  assign n45865 = n45857 & ~n45864;
  assign n45866 = n2748 & ~n41149;
  assign n45867 = ~pi32 & ~n45866;
  assign n45868 = n45853 & ~n45867;
  assign n45869 = pi1093 & ~n45864;
  assign n45870 = ~n45868 & n45869;
  assign n45871 = ~n45865 & ~n45870;
  assign n45872 = n40596 & ~n45871;
  assign n45873 = n45860 & n45872;
  assign n45874 = ~n45863 & ~n45873;
  assign n45875 = ~n45840 & n45874;
  assign n45876 = pi332 & ~n45875;
  assign n45877 = pi1093 & ~n41099;
  assign n45878 = ~n45865 & ~n45877;
  assign n45879 = n40634 & ~n45878;
  assign n45880 = ~n45872 & ~n45879;
  assign n45881 = ~n45847 & n45880;
  assign n45882 = ~pi332 & ~n45881;
  assign n45883 = ~n45876 & ~n45882;
  assign n45884 = ~n30860 & n45883;
  assign n45885 = ~pi210 & ~n45884;
  assign n45886 = ~pi210 & ~n45851;
  assign n45887 = ~n45884 & n45886;
  assign n45888 = ~n45851 & n45885;
  assign n45889 = ~n33962 & ~n41183;
  assign n45890 = pi137 & ~n45889;
  assign n45891 = ~n41189 & ~n45890;
  assign n45892 = ~pi332 & ~n45891;
  assign n45893 = ~n41177 & ~n45836;
  assign n45894 = ~pi95 & ~n45893;
  assign n45895 = n41290 & ~n45894;
  assign n45896 = ~pi137 & n41178;
  assign n45897 = ~n45841 & n45896;
  assign n45898 = pi332 & ~n45897;
  assign n45899 = ~n45895 & n45898;
  assign n45900 = ~n45892 & ~n45899;
  assign n45901 = pi210 & ~n45900;
  assign n45902 = pi299 & ~n45901;
  assign n45903 = ~n64939 & n45902;
  assign n45904 = ~n30858 & n45883;
  assign n45905 = n30858 & n45850;
  assign n45906 = ~pi198 & ~n45905;
  assign n45907 = ~pi198 & ~n45904;
  assign n45908 = ~n45905 & n45907;
  assign n45909 = ~n45904 & n45906;
  assign n45910 = pi198 & ~n45900;
  assign n45911 = ~pi299 & ~n45910;
  assign n45912 = ~n64940 & n45911;
  assign n45913 = ~n45903 & ~n45912;
  assign n45914 = ~pi39 & ~n45913;
  assign n45915 = pi39 & n41528;
  assign n45916 = ~pi38 & ~n45915;
  assign n45917 = ~n45914 & n45916;
  assign n45918 = pi38 & ~pi137;
  assign n45919 = n33858 & ~n45918;
  assign n45920 = ~n45917 & n45919;
  assign n45921 = ~n45832 & ~n45920;
  assign n45922 = ~pi87 & ~n45921;
  assign n45923 = n62373 & n41528;
  assign n45924 = pi87 & n45923;
  assign n45925 = ~pi75 & ~n45924;
  assign n45926 = ~n45922 & n45925;
  assign n45927 = n30599 & ~n45831;
  assign n45928 = pi75 & ~n45927;
  assign n45929 = ~pi92 & ~n45928;
  assign n45930 = ~n45926 & n45929;
  assign n45931 = pi92 & n64083;
  assign n45932 = pi92 & n6795;
  assign n45933 = n45923 & n45932;
  assign n45934 = n41528 & n45931;
  assign n45935 = ~pi54 & ~n64941;
  assign n45936 = ~n45930 & n45935;
  assign n45937 = n6796 & n45923;
  assign n45938 = pi54 & ~n45937;
  assign n45939 = ~pi74 & ~n45938;
  assign n45940 = ~n45936 & n45939;
  assign n45941 = pi74 & n30592;
  assign n45942 = ~pi54 & pi74;
  assign n45943 = n45937 & n45942;
  assign n45944 = n45923 & n45941;
  assign n45945 = ~pi55 & ~n64942;
  assign n45946 = ~n45940 & n45945;
  assign n45947 = n30904 & ~n45946;
  assign n45948 = pi56 & n30584;
  assign n45949 = n45923 & n45948;
  assign n45950 = ~n45947 & ~n45949;
  assign n45951 = ~pi62 & ~n45950;
  assign n45952 = n34046 & n45923;
  assign n45953 = pi62 & n45952;
  assign n45954 = n3472 & ~n45953;
  assign n45955 = ~n45951 & n45954;
  assign n45956 = ~pi62 & n45952;
  assign n45957 = ~n3472 & ~n45956;
  assign n45958 = ~n30570 & ~n45957;
  assign po382 = ~n45955 & n45958;
  assign n45960 = ~pi939 & n41469;
  assign n45961 = ~pi1146 & ~n41469;
  assign n45962 = pi222 & ~n45961;
  assign n45963 = pi222 & ~n45960;
  assign n45964 = ~n45961 & n45963;
  assign n45965 = ~n45960 & n45962;
  assign n45966 = pi276 & n28811;
  assign n45967 = ~pi223 & ~n45966;
  assign n45968 = ~pi223 & ~n64943;
  assign n45969 = ~n45966 & n45968;
  assign n45970 = ~n64943 & n45967;
  assign n45971 = pi223 & ~pi1146;
  assign n45972 = ~pi299 & ~n45971;
  assign n45973 = ~n64944 & n45972;
  assign n45974 = ~pi939 & n41020;
  assign n45975 = ~pi1146 & ~n41020;
  assign n45976 = pi221 & ~n45975;
  assign n45977 = pi221 & ~n45974;
  assign n45978 = ~n45975 & n45977;
  assign n45979 = ~n45974 & n45976;
  assign n45980 = pi215 & pi1146;
  assign n45981 = ~pi216 & ~pi228;
  assign n45982 = ~n45980 & n45981;
  assign n45983 = ~n64945 & ~n45980;
  assign n45984 = n45981 & n45983;
  assign n45985 = ~n64945 & n45982;
  assign n45986 = ~pi216 & n34059;
  assign n45987 = n45983 & n45986;
  assign n45988 = n62380 & n64946;
  assign n45989 = pi276 & n39839;
  assign n45990 = ~pi216 & ~n41010;
  assign n45991 = ~n45989 & ~n45990;
  assign n45992 = ~pi221 & ~n45991;
  assign n45993 = ~n64945 & ~n45992;
  assign n45994 = ~pi215 & ~n45993;
  assign n45995 = ~n45980 & ~n45994;
  assign n45996 = pi299 & ~n45995;
  assign n45997 = ~n64947 & n45996;
  assign n45998 = ~n45973 & ~n45997;
  assign n45999 = ~pi154 & ~n45998;
  assign n46000 = ~n64945 & ~n45989;
  assign n46001 = ~pi215 & ~n46000;
  assign n46002 = ~n45980 & ~n46001;
  assign n46003 = pi299 & ~n46002;
  assign n46004 = ~n45973 & ~n46003;
  assign n46005 = pi154 & ~n46004;
  assign n46006 = n62373 & ~n46005;
  assign n46007 = ~n45999 & n46006;
  assign n46008 = pi154 & ~n46002;
  assign n46009 = ~pi154 & ~n45995;
  assign n46010 = ~n46008 & ~n46009;
  assign n46011 = pi299 & ~n46010;
  assign n46012 = ~n45973 & ~n46011;
  assign n46013 = ~n62373 & n46012;
  assign n46014 = ~n46007 & ~n46013;
  assign n46015 = pi87 & ~n46014;
  assign n46016 = n43708 & n64946;
  assign n46017 = n45996 & ~n46016;
  assign n46018 = ~n45973 & ~n46017;
  assign n46019 = ~pi154 & ~n46018;
  assign n46020 = ~pi38 & ~n46005;
  assign n46021 = ~n46019 & n46020;
  assign n46022 = pi38 & n46012;
  assign n46023 = ~pi100 & ~n46022;
  assign n46024 = ~n46021 & n46023;
  assign n46025 = n2764 & n33591;
  assign n46026 = ~pi38 & ~pi216;
  assign n46027 = ~pi228 & n46026;
  assign n46028 = ~pi39 & n33591;
  assign n46029 = n46027 & n46028;
  assign n46030 = n45983 & n46029;
  assign n46031 = n64946 & n46025;
  assign n46032 = n44422 & n64948;
  assign n46033 = pi100 & ~n46012;
  assign n46034 = ~n46032 & n46033;
  assign n46035 = ~pi87 & ~n46034;
  assign n46036 = ~n46024 & n46035;
  assign n46037 = ~n46015 & ~n46036;
  assign n46038 = ~pi75 & ~n46037;
  assign n46039 = pi75 & n46012;
  assign n46040 = ~pi92 & ~n46039;
  assign n46041 = ~n46038 & n46040;
  assign n46042 = n6795 & n46007;
  assign n46043 = ~n64083 & n46012;
  assign n46044 = pi92 & ~n46043;
  assign n46045 = ~n46042 & n46044;
  assign n46046 = n6792 & ~n46045;
  assign n46047 = ~n46041 & n46046;
  assign n46048 = ~n6792 & n46012;
  assign n46049 = ~pi55 & ~n46048;
  assign n46050 = ~n46047 & n46049;
  assign n46051 = n64082 & n64947;
  assign n46052 = pi55 & ~n46010;
  assign n46053 = ~n46051 & n46052;
  assign n46054 = ~pi56 & ~n46053;
  assign n46055 = ~n46050 & n46054;
  assign n46056 = n64084 & ~n46010;
  assign n46057 = ~n64947 & n46056;
  assign n46058 = ~n64084 & ~n46010;
  assign n46059 = pi56 & ~n46058;
  assign n46060 = ~n46057 & n46059;
  assign n46061 = ~pi62 & ~n46060;
  assign n46062 = ~n46055 & n46061;
  assign n46063 = ~n44475 & ~n46010;
  assign n46064 = ~n46057 & ~n46063;
  assign n46065 = pi62 & ~n46064;
  assign n46066 = n3472 & ~n46065;
  assign n46067 = ~n46062 & n46066;
  assign n46068 = ~n3472 & n46010;
  assign n46069 = ~pi239 & ~n46068;
  assign n46070 = ~n46067 & n46069;
  assign n46071 = ~pi154 & ~n45168;
  assign n46072 = pi154 & ~n45159;
  assign n46073 = n38199 & ~n46072;
  assign n46074 = ~n46071 & n46073;
  assign n46075 = n46002 & ~n46074;
  assign n46076 = pi299 & ~n46075;
  assign n46077 = ~pi224 & n44321;
  assign n46078 = pi224 & ~pi276;
  assign n46079 = ~pi222 & ~n46078;
  assign n46080 = ~n46077 & n46079;
  assign n46081 = n45968 & ~n46080;
  assign n46082 = n45972 & ~n46081;
  assign n46083 = ~pi39 & ~n46082;
  assign n46084 = ~n45971 & ~n46081;
  assign n46085 = ~pi299 & ~n46084;
  assign n46086 = pi299 & n46002;
  assign n46087 = ~n46074 & n46086;
  assign n46088 = ~n46085 & ~n46087;
  assign n46089 = ~pi39 & ~n46088;
  assign n46090 = ~n46076 & n46083;
  assign n46091 = ~n44399 & n46002;
  assign n46092 = pi154 & ~n46091;
  assign n46093 = ~pi215 & ~n46091;
  assign n46094 = ~n46009 & ~n46093;
  assign n46095 = ~n46009 & ~n46092;
  assign n46096 = ~n46093 & n46095;
  assign n46097 = ~n46092 & n46094;
  assign n46098 = pi299 & ~n64950;
  assign n46099 = ~n64897 & ~n45973;
  assign n46100 = ~n46098 & n46099;
  assign n46101 = ~n64947 & ~n64950;
  assign n46102 = pi299 & ~n46101;
  assign n46103 = ~n46100 & ~n46102;
  assign n46104 = pi39 & ~n46103;
  assign n46105 = n2766 & ~n46104;
  assign n46106 = ~n64949 & n46105;
  assign n46107 = pi100 & n46032;
  assign n46108 = ~n2766 & ~n46100;
  assign n46109 = ~n46107 & n46108;
  assign n46110 = ~n46106 & ~n46109;
  assign n46111 = ~pi87 & ~n46110;
  assign n46112 = n62373 & n46102;
  assign n46113 = pi87 & ~n46100;
  assign n46114 = ~n46112 & n46113;
  assign n46115 = ~pi75 & ~n46114;
  assign n46116 = ~n46111 & n46115;
  assign n46117 = pi75 & n46100;
  assign n46118 = ~pi92 & ~n46117;
  assign n46119 = ~n46116 & n46118;
  assign n46120 = n6795 & n46112;
  assign n46121 = n64083 & n46102;
  assign n46122 = pi92 & ~n46100;
  assign n46123 = ~n64951 & n46122;
  assign n46124 = n6792 & ~n46123;
  assign n46125 = ~n46119 & n46124;
  assign n46126 = ~n6792 & n46100;
  assign n46127 = ~pi55 & ~n46126;
  assign n46128 = ~n46125 & n46127;
  assign n46129 = pi55 & ~n64950;
  assign n46130 = ~n46051 & n46129;
  assign n46131 = ~pi56 & ~n46130;
  assign n46132 = ~n46128 & n46131;
  assign n46133 = ~n64084 & ~n64950;
  assign n46134 = pi56 & ~n46133;
  assign n46135 = n64084 & n46101;
  assign n46136 = n46134 & ~n46135;
  assign n46137 = ~n46101 & n46134;
  assign n46138 = ~pi62 & ~n64952;
  assign n46139 = ~n46132 & n46138;
  assign n46140 = n44475 & n64947;
  assign n46141 = pi62 & ~n64950;
  assign n46142 = ~n44475 & ~n64950;
  assign n46143 = ~pi56 & n46135;
  assign n46144 = ~n46142 & ~n46143;
  assign n46145 = pi62 & ~n46144;
  assign n46146 = ~n46140 & n46141;
  assign n46147 = n3472 & ~n64953;
  assign n46148 = ~n46139 & n46147;
  assign n46149 = ~n3472 & n64950;
  assign n46150 = pi239 & ~n46149;
  assign n46151 = ~n46148 & n46150;
  assign n46152 = ~n46070 & ~n46151;
  assign n46153 = ~pi927 & n41020;
  assign n46154 = ~pi1145 & ~n41020;
  assign n46155 = pi221 & ~n46154;
  assign n46156 = pi221 & ~n46153;
  assign n46157 = ~n46154 & n46156;
  assign n46158 = ~n46153 & n46155;
  assign n46159 = pi216 & pi274;
  assign n46160 = ~pi221 & ~n46159;
  assign n46161 = ~pi151 & n45168;
  assign n46162 = pi151 & n45159;
  assign n46163 = ~pi216 & ~n46162;
  assign n46164 = ~n46161 & n46163;
  assign n46165 = n46160 & ~n46164;
  assign n46166 = ~n64954 & ~n46165;
  assign n46167 = ~pi215 & ~n46166;
  assign n46168 = pi215 & pi1145;
  assign n46169 = pi299 & ~n46168;
  assign n46170 = ~n46167 & n46169;
  assign n46171 = ~pi927 & n41469;
  assign n46172 = ~pi1145 & ~n41469;
  assign n46173 = pi222 & ~n46172;
  assign n46174 = pi222 & ~n46171;
  assign n46175 = ~n46172 & n46174;
  assign n46176 = ~n46171 & n46173;
  assign n46177 = pi224 & pi274;
  assign n46178 = ~pi222 & ~n46177;
  assign n46179 = ~n46077 & n46178;
  assign n46180 = ~n64955 & ~n46179;
  assign n46181 = ~pi223 & ~n46180;
  assign n46182 = pi223 & pi1145;
  assign n46183 = ~pi299 & ~n46182;
  assign n46184 = ~n46181 & n46183;
  assign n46185 = ~pi39 & ~n46184;
  assign n46186 = ~n46170 & n46185;
  assign n46187 = n28811 & ~n46177;
  assign n46188 = ~n64955 & ~n46187;
  assign n46189 = ~pi223 & ~n46188;
  assign n46190 = ~n46182 & ~n46189;
  assign n46191 = ~pi299 & ~n46190;
  assign n46192 = ~n64897 & ~n46191;
  assign n46193 = ~pi151 & ~n41010;
  assign n46194 = ~n44384 & ~n46193;
  assign n46195 = ~pi151 & n34059;
  assign n46196 = ~n46194 & ~n46195;
  assign n46197 = ~pi216 & ~n46196;
  assign n46198 = n46160 & ~n46197;
  assign n46199 = ~n64954 & ~n46198;
  assign n46200 = ~pi215 & ~n46199;
  assign n46201 = ~n46168 & ~n46200;
  assign n46202 = pi299 & ~n46201;
  assign n46203 = n46192 & ~n46202;
  assign n46204 = pi39 & ~n46203;
  assign n46205 = ~pi38 & ~n46204;
  assign n46206 = ~n46186 & n46205;
  assign n46207 = ~pi216 & ~n46193;
  assign n46208 = n46160 & ~n46207;
  assign n46209 = ~n64954 & ~n46208;
  assign n46210 = ~pi215 & ~n46209;
  assign n46211 = ~n46168 & ~n46210;
  assign n46212 = n44656 & ~n46159;
  assign n46213 = n46211 & ~n46212;
  assign n46214 = pi299 & ~n46213;
  assign n46215 = n46192 & ~n46214;
  assign n46216 = pi38 & n46215;
  assign n46217 = ~pi100 & ~n46216;
  assign n46218 = ~n46206 & n46217;
  assign n46219 = ~pi151 & n45093;
  assign n46220 = n46197 & ~n46219;
  assign n46221 = n46160 & ~n46220;
  assign n46222 = ~n64954 & ~n46221;
  assign n46223 = ~pi215 & ~n46222;
  assign n46224 = ~n46168 & ~n46223;
  assign n46225 = pi299 & ~n46224;
  assign n46226 = n2764 & n46192;
  assign n46227 = ~n46225 & n46226;
  assign n46228 = ~n2764 & n46215;
  assign n46229 = pi100 & ~n46228;
  assign n46230 = ~n46227 & n46229;
  assign n46231 = ~n46218 & ~n46230;
  assign n46232 = ~pi87 & ~n46231;
  assign n46233 = ~n62373 & n46215;
  assign n46234 = n62373 & n46203;
  assign n46235 = ~n46233 & ~n46234;
  assign n46236 = pi87 & n46235;
  assign n46237 = ~pi75 & ~n46236;
  assign n46238 = ~n46232 & n46237;
  assign n46239 = pi75 & n46215;
  assign n46240 = ~pi92 & ~n46239;
  assign n46241 = ~n46238 & n46240;
  assign n46242 = n6795 & ~n46235;
  assign n46243 = ~n6795 & n46215;
  assign n46244 = pi92 & ~n46243;
  assign n46245 = ~n46242 & n46244;
  assign n46246 = n6792 & ~n46245;
  assign n46247 = ~n46241 & n46246;
  assign n46248 = ~n6792 & n46215;
  assign n46249 = ~pi55 & ~n46248;
  assign n46250 = ~n46247 & n46249;
  assign n46251 = n64082 & n46201;
  assign n46252 = ~n64082 & n46213;
  assign n46253 = pi55 & ~n46252;
  assign n46254 = ~n46251 & n46253;
  assign n46255 = ~pi56 & ~n46254;
  assign n46256 = ~n46250 & n46255;
  assign n46257 = n64084 & ~n46201;
  assign n46258 = ~n64084 & ~n46213;
  assign n46259 = pi56 & ~n46258;
  assign n46260 = ~n64084 & n46213;
  assign n46261 = ~pi55 & n46251;
  assign n46262 = ~n46260 & ~n46261;
  assign n46263 = pi56 & ~n46262;
  assign n46264 = ~n46257 & n46259;
  assign n46265 = ~pi62 & ~n64956;
  assign n46266 = ~n46256 & n46265;
  assign n46267 = n44475 & n46201;
  assign n46268 = ~n44475 & n46213;
  assign n46269 = pi62 & ~n46268;
  assign n46270 = ~n46267 & n46269;
  assign n46271 = pi235 & n3472;
  assign n46272 = ~n46270 & n46271;
  assign n46273 = ~n46266 & n46272;
  assign n46274 = pi299 & ~n46211;
  assign n46275 = ~pi87 & ~n43708;
  assign n46276 = pi87 & ~n7356;
  assign n46277 = ~pi100 & ~n46276;
  assign n46278 = ~n46275 & n46277;
  assign n46279 = pi100 & n2805;
  assign n46280 = n44422 & n46279;
  assign n46281 = ~n46278 & ~n46280;
  assign n46282 = n45981 & ~n46168;
  assign n46283 = ~n64954 & n46282;
  assign n46284 = ~n64954 & ~n46168;
  assign n46285 = n46027 & n46284;
  assign n46286 = ~pi38 & n46283;
  assign n46287 = ~n46281 & n64957;
  assign n46288 = n46274 & ~n46287;
  assign n46289 = ~pi75 & ~n46191;
  assign n46290 = n45986 & n46284;
  assign n46291 = n62380 & n46283;
  assign n46292 = n46274 & ~n64958;
  assign n46293 = n62373 & ~n46191;
  assign n46294 = ~n46292 & n46293;
  assign n46295 = ~n46191 & ~n46274;
  assign n46296 = ~n62373 & n46295;
  assign n46297 = ~n46294 & ~n46296;
  assign n46298 = pi87 & ~n46297;
  assign n46299 = ~pi100 & n43708;
  assign n46300 = n39702 & n44422;
  assign n46301 = ~n46299 & ~n46300;
  assign n46302 = n64957 & ~n46301;
  assign n46303 = n46274 & ~n46302;
  assign n46304 = ~pi87 & ~n46191;
  assign n46305 = ~n46303 & n46304;
  assign n46306 = ~n46298 & ~n46305;
  assign n46307 = ~pi75 & ~n46306;
  assign n46308 = ~n46288 & n46289;
  assign n46309 = pi75 & n46295;
  assign n46310 = ~pi92 & ~n46309;
  assign n46311 = ~n64959 & n46310;
  assign n46312 = n64083 & ~n46191;
  assign n46313 = n64958 & n46312;
  assign n46314 = pi92 & ~n46295;
  assign n46315 = n6795 & n46294;
  assign n46316 = ~n64083 & n46295;
  assign n46317 = pi92 & ~n46316;
  assign n46318 = ~n46315 & n46317;
  assign n46319 = ~n46313 & n46314;
  assign n46320 = n6792 & ~n64960;
  assign n46321 = ~n46311 & n46320;
  assign n46322 = ~n6792 & n46295;
  assign n46323 = ~pi55 & ~n46322;
  assign n46324 = ~n46321 & n46323;
  assign n46325 = n64082 & n64958;
  assign n46326 = pi55 & ~n46211;
  assign n46327 = ~n46325 & n46326;
  assign n46328 = ~pi56 & ~n46327;
  assign n46329 = ~n46324 & n46328;
  assign n46330 = ~pi55 & n46325;
  assign n46331 = n64084 & n64958;
  assign n46332 = ~n46211 & ~n64961;
  assign n46333 = pi56 & ~n46332;
  assign n46334 = ~pi62 & ~n46333;
  assign n46335 = ~n46329 & n46334;
  assign n46336 = ~pi56 & n64961;
  assign n46337 = n44475 & n64958;
  assign n46338 = pi62 & ~n46211;
  assign n46339 = ~n64962 & n46338;
  assign n46340 = ~pi235 & n3472;
  assign n46341 = ~n46339 & n46340;
  assign n46342 = ~n46335 & n46341;
  assign n46343 = pi235 & n46212;
  assign n46344 = ~n3472 & ~n46343;
  assign n46345 = n46211 & n46344;
  assign n46346 = ~n46342 & ~n46345;
  assign po155 = ~n46273 & n46346;
  assign n46348 = pi223 & pi1143;
  assign n46349 = ~pi299 & ~n46348;
  assign n46350 = ~pi944 & n41469;
  assign n46351 = ~pi1143 & ~n41469;
  assign n46352 = pi222 & ~n46351;
  assign n46353 = pi222 & ~n46350;
  assign n46354 = ~n46351 & n46353;
  assign n46355 = ~n46350 & n46352;
  assign n46356 = pi224 & pi264;
  assign n46357 = ~pi222 & ~n46356;
  assign n46358 = ~pi284 & n44321;
  assign n46359 = ~pi224 & ~n46358;
  assign n46360 = n46357 & ~n46359;
  assign n46361 = ~n64963 & ~n46360;
  assign n46362 = ~n44321 & n46357;
  assign n46363 = n46361 & ~n46362;
  assign n46364 = ~pi223 & ~n46363;
  assign n46365 = n46349 & ~n46364;
  assign n46366 = ~pi39 & ~n46365;
  assign n46367 = pi215 & pi1143;
  assign n46368 = pi299 & ~n46367;
  assign n46369 = ~pi944 & n41020;
  assign n46370 = ~pi1143 & ~n41020;
  assign n46371 = pi221 & ~n46370;
  assign n46372 = pi221 & ~n46369;
  assign n46373 = ~n46370 & n46372;
  assign n46374 = ~n46369 & n46371;
  assign n46375 = pi216 & pi264;
  assign n46376 = ~pi221 & ~n46375;
  assign n46377 = pi284 & ~n30613;
  assign n46378 = pi105 & ~n46377;
  assign n46379 = ~pi105 & pi146;
  assign n46380 = pi228 & ~n46379;
  assign n46381 = ~n46378 & n46380;
  assign n46382 = ~n44337 & n46381;
  assign n46383 = pi146 & ~n44316;
  assign n46384 = ~pi146 & n44327;
  assign n46385 = pi284 & ~n46384;
  assign n46386 = ~n46383 & n46385;
  assign n46387 = ~pi146 & ~pi284;
  assign n46388 = ~n43706 & n46387;
  assign n46389 = ~n46386 & ~n46388;
  assign n46390 = ~pi228 & ~n46389;
  assign n46391 = ~n46382 & ~n46390;
  assign n46392 = ~pi216 & ~n46391;
  assign n46393 = n46376 & ~n46392;
  assign n46394 = ~n64964 & ~n46393;
  assign n46395 = ~pi215 & ~n46394;
  assign n46396 = n46368 & ~n46395;
  assign n46397 = n46366 & ~n46396;
  assign n46398 = ~pi224 & n46377;
  assign n46399 = n46357 & ~n46398;
  assign n46400 = ~n64963 & ~n46399;
  assign n46401 = ~pi223 & ~n46400;
  assign n46402 = ~n46348 & ~n46401;
  assign n46403 = ~pi299 & ~n46402;
  assign n46404 = ~pi284 & n62380;
  assign n46405 = pi146 & ~n62380;
  assign n46406 = ~pi228 & ~n46405;
  assign n46407 = pi284 & n62380;
  assign n46408 = ~n44414 & ~n46407;
  assign n46409 = ~pi228 & ~n46408;
  assign n46410 = ~n46404 & n46406;
  assign n46411 = ~n46381 & ~n64965;
  assign n46412 = ~pi216 & ~n46411;
  assign n46413 = n46376 & ~n46412;
  assign n46414 = ~n64964 & ~n46413;
  assign n46415 = ~pi215 & ~n46414;
  assign n46416 = ~n46367 & ~n46415;
  assign n46417 = pi299 & ~n46416;
  assign n46418 = ~n46403 & ~n46417;
  assign n46419 = pi39 & ~n46418;
  assign n46420 = ~pi38 & ~n46419;
  assign n46421 = ~n46397 & n46420;
  assign n46422 = ~n44384 & ~n46381;
  assign n46423 = ~pi146 & ~pi228;
  assign n46424 = n46422 & ~n46423;
  assign n46425 = ~pi216 & ~n46424;
  assign n46426 = n46376 & ~n46425;
  assign n46427 = ~n64964 & ~n46426;
  assign n46428 = ~pi215 & ~n46427;
  assign n46429 = ~n46367 & ~n46428;
  assign n46430 = n44656 & ~n46375;
  assign n46431 = n46429 & ~n46430;
  assign n46432 = pi299 & ~n46431;
  assign n46433 = ~n46403 & ~n46432;
  assign n46434 = pi38 & n46433;
  assign n46435 = ~pi100 & ~n46434;
  assign n46436 = ~n46421 & n46435;
  assign n46437 = pi252 & n2811;
  assign n46438 = ~pi284 & ~n46437;
  assign n46439 = n46404 & ~n46437;
  assign n46440 = n62380 & n46438;
  assign n46441 = ~pi228 & ~n64966;
  assign n46442 = ~pi228 & ~n44413;
  assign n46443 = ~n64966 & n46442;
  assign n46444 = ~n44413 & n46441;
  assign n46445 = ~n46381 & ~n64967;
  assign n46446 = ~pi216 & ~n46445;
  assign n46447 = n46376 & ~n46446;
  assign n46448 = ~n64964 & ~n46447;
  assign n46449 = ~pi215 & ~n46448;
  assign n46450 = ~n46367 & ~n46449;
  assign n46451 = pi299 & ~n46450;
  assign n46452 = n2764 & ~n46403;
  assign n46453 = ~n46451 & n46452;
  assign n46454 = ~n2764 & n46433;
  assign n46455 = pi100 & ~n46454;
  assign n46456 = ~n46453 & n46455;
  assign n46457 = ~n46436 & ~n46456;
  assign n46458 = ~pi87 & ~n46457;
  assign n46459 = ~n62373 & n46433;
  assign n46460 = n62373 & n46418;
  assign n46461 = ~n46459 & ~n46460;
  assign n46462 = pi87 & n46461;
  assign n46463 = ~pi75 & ~n46462;
  assign n46464 = ~n46458 & n46463;
  assign n46465 = pi75 & n46433;
  assign n46466 = ~pi92 & ~n46465;
  assign n46467 = ~n46464 & n46466;
  assign n46468 = n6795 & ~n46461;
  assign n46469 = ~n6795 & n46433;
  assign n46470 = pi92 & ~n46469;
  assign n46471 = ~n46468 & n46470;
  assign n46472 = n6792 & ~n46471;
  assign n46473 = ~n46467 & n46472;
  assign n46474 = ~n6792 & n46433;
  assign n46475 = ~pi55 & ~n46474;
  assign n46476 = ~n46473 & n46475;
  assign n46477 = n64082 & n46416;
  assign n46478 = ~n64082 & n46431;
  assign n46479 = pi55 & ~n46478;
  assign n46480 = ~n46477 & n46479;
  assign n46481 = ~pi56 & ~n46480;
  assign n46482 = ~n46476 & n46481;
  assign n46483 = n64084 & ~n46416;
  assign n46484 = ~n64084 & ~n46431;
  assign n46485 = pi56 & ~n46484;
  assign n46486 = ~pi55 & n46477;
  assign n46487 = ~n64084 & n46431;
  assign n46488 = ~n46486 & ~n46487;
  assign n46489 = pi56 & ~n46488;
  assign n46490 = ~n46483 & n46485;
  assign n46491 = ~pi62 & ~n64968;
  assign n46492 = ~n46482 & n46491;
  assign n46493 = n44475 & n46416;
  assign n46494 = ~n44475 & n46431;
  assign n46495 = pi62 & ~n46494;
  assign n46496 = ~n46493 & n46495;
  assign n46497 = pi238 & n3472;
  assign n46498 = ~n46496 & n46497;
  assign n46499 = ~n46492 & n46498;
  assign n46500 = ~pi146 & ~n44316;
  assign n46501 = pi146 & n44327;
  assign n46502 = ~pi284 & ~n46501;
  assign n46503 = ~n46500 & n46502;
  assign n46504 = pi146 & pi284;
  assign n46505 = ~n43706 & n46504;
  assign n46506 = ~pi228 & ~n46505;
  assign n46507 = pi146 & ~n43706;
  assign n46508 = pi284 & ~n46507;
  assign n46509 = ~pi146 & n44316;
  assign n46510 = pi146 & ~n44327;
  assign n46511 = ~pi284 & ~n46510;
  assign n46512 = ~n46509 & n46511;
  assign n46513 = ~n46502 & ~n46505;
  assign n46514 = ~n46500 & ~n46513;
  assign n46515 = ~n46508 & ~n46512;
  assign n46516 = ~pi228 & ~n64969;
  assign n46517 = ~n46503 & n46506;
  assign n46518 = ~n44611 & ~n46381;
  assign n46519 = ~n64970 & n46518;
  assign n46520 = ~pi216 & ~n46519;
  assign n46521 = n46376 & ~n46520;
  assign n46522 = ~n64964 & ~n46521;
  assign n46523 = ~pi215 & ~n46522;
  assign n46524 = n46368 & ~n46523;
  assign n46525 = n46349 & n46361;
  assign n46526 = n46366 & ~n46525;
  assign n46527 = ~n46524 & n46526;
  assign n46528 = ~n44372 & n46403;
  assign n46529 = ~n64965 & n46422;
  assign n46530 = ~pi216 & ~n46529;
  assign n46531 = n46376 & ~n46530;
  assign n46532 = ~n64964 & ~n46531;
  assign n46533 = ~pi215 & ~n46532;
  assign n46534 = ~n46367 & ~n46533;
  assign n46535 = pi299 & ~n46534;
  assign n46536 = ~n46528 & ~n46535;
  assign n46537 = pi39 & ~n46536;
  assign n46538 = ~pi38 & ~n46537;
  assign n46539 = ~n46527 & n46538;
  assign n46540 = pi299 & ~n46429;
  assign n46541 = ~n46528 & ~n46540;
  assign n46542 = pi38 & n46541;
  assign n46543 = ~pi100 & ~n46542;
  assign n46544 = ~n46539 & n46543;
  assign n46545 = n46422 & ~n64967;
  assign n46546 = ~pi216 & ~n46545;
  assign n46547 = n46376 & ~n46546;
  assign n46548 = ~n64964 & ~n46547;
  assign n46549 = ~pi215 & ~n46548;
  assign n46550 = ~n46367 & ~n46549;
  assign n46551 = pi299 & ~n46550;
  assign n46552 = n2764 & ~n46528;
  assign n46553 = ~n46551 & n46552;
  assign n46554 = ~n2764 & n46541;
  assign n46555 = pi100 & ~n46554;
  assign n46556 = ~n46553 & n46555;
  assign n46557 = ~n46544 & ~n46556;
  assign n46558 = ~pi87 & ~n46557;
  assign n46559 = ~n62373 & n46541;
  assign n46560 = n62373 & n46536;
  assign n46561 = ~n46559 & ~n46560;
  assign n46562 = pi87 & n46561;
  assign n46563 = ~pi75 & ~n46562;
  assign n46564 = ~n46558 & n46563;
  assign n46565 = pi75 & n46541;
  assign n46566 = ~pi92 & ~n46565;
  assign n46567 = ~n46564 & n46566;
  assign n46568 = n6795 & ~n46561;
  assign n46569 = ~n6795 & n46541;
  assign n46570 = pi92 & ~n46569;
  assign n46571 = ~n46568 & n46570;
  assign n46572 = n6792 & ~n46571;
  assign n46573 = ~n46567 & n46572;
  assign n46574 = ~n6792 & n46541;
  assign n46575 = ~pi55 & ~n46574;
  assign n46576 = ~n46573 & n46575;
  assign n46577 = n64082 & n46534;
  assign n46578 = ~n64082 & n46429;
  assign n46579 = pi55 & ~n46578;
  assign n46580 = ~n46577 & n46579;
  assign n46581 = ~pi56 & ~n46580;
  assign n46582 = ~n46576 & n46581;
  assign n46583 = n64084 & ~n46534;
  assign n46584 = ~n64084 & ~n46429;
  assign n46585 = pi56 & ~n46584;
  assign n46586 = ~n64084 & n46429;
  assign n46587 = ~pi55 & n46577;
  assign n46588 = ~n46586 & ~n46587;
  assign n46589 = pi56 & ~n46588;
  assign n46590 = ~n46583 & n46585;
  assign n46591 = ~pi62 & ~n64971;
  assign n46592 = ~n46582 & n46591;
  assign n46593 = n44475 & n46534;
  assign n46594 = ~n44475 & n46429;
  assign n46595 = pi62 & ~n46594;
  assign n46596 = ~n46593 & n46595;
  assign n46597 = ~pi238 & n3472;
  assign n46598 = ~n46596 & n46597;
  assign n46599 = ~n46592 & n46598;
  assign n46600 = pi238 & n46430;
  assign n46601 = ~n3472 & ~n46600;
  assign n46602 = n46429 & n46601;
  assign n46603 = ~n46599 & ~n46602;
  assign n46604 = ~n46499 & ~n46602;
  assign n46605 = ~n46599 & n46604;
  assign n46606 = ~n46499 & n46603;
  assign n46607 = ~pi928 & n41020;
  assign n46608 = ~pi1136 & ~n41020;
  assign n46609 = pi221 & ~n46608;
  assign n46610 = pi221 & ~n46607;
  assign n46611 = ~n46608 & n46610;
  assign n46612 = ~n46607 & n46609;
  assign n46613 = pi216 & pi266;
  assign n46614 = ~pi166 & ~n44316;
  assign n46615 = pi166 & n44327;
  assign n46616 = pi875 & ~n46615;
  assign n46617 = ~n46614 & n46616;
  assign n46618 = pi166 & ~pi875;
  assign n46619 = ~n43706 & n46618;
  assign n46620 = ~pi228 & ~n46619;
  assign n46621 = ~n46617 & n46620;
  assign n46622 = pi875 & ~n30613;
  assign n46623 = pi105 & ~n46622;
  assign n46624 = ~pi105 & ~pi166;
  assign n46625 = ~n46623 & ~n46624;
  assign n46626 = n45157 & ~n46625;
  assign n46627 = ~pi216 & ~n46626;
  assign n46628 = ~n44611 & n46627;
  assign n46629 = ~n46617 & ~n46619;
  assign n46630 = ~pi228 & ~n46629;
  assign n46631 = ~n45157 & ~n46630;
  assign n46632 = n46627 & ~n46631;
  assign n46633 = ~n46621 & n46628;
  assign n46634 = ~n46613 & ~n64974;
  assign n46635 = ~pi221 & ~n46634;
  assign n46636 = ~n64973 & ~n46635;
  assign n46637 = ~pi215 & ~n46636;
  assign n46638 = pi215 & pi1136;
  assign n46639 = pi299 & ~n46638;
  assign n46640 = ~n46637 & n46639;
  assign n46641 = ~pi224 & ~pi875;
  assign n46642 = ~n30613 & n46641;
  assign n46643 = pi224 & ~pi266;
  assign n46644 = ~pi222 & ~n46643;
  assign n46645 = ~n46642 & n46644;
  assign n46646 = n7034 & ~n44321;
  assign n46647 = n46645 & ~n46646;
  assign n46648 = ~pi928 & n41469;
  assign n46649 = ~pi1136 & ~n41469;
  assign n46650 = pi222 & ~n46649;
  assign n46651 = pi222 & ~n46648;
  assign n46652 = ~n46649 & n46651;
  assign n46653 = ~n46648 & n46650;
  assign n46654 = pi223 & pi1136;
  assign n46655 = ~pi299 & ~n46654;
  assign n46656 = ~n64975 & n46655;
  assign n46657 = ~n46647 & n46656;
  assign n46658 = ~n46645 & ~n64975;
  assign n46659 = ~n46646 & n46658;
  assign n46660 = ~pi223 & ~n46659;
  assign n46661 = n46655 & ~n46660;
  assign n46662 = ~pi39 & ~n46661;
  assign n46663 = ~n46657 & n46662;
  assign n46664 = ~n46640 & n46663;
  assign n46665 = ~pi223 & ~n46658;
  assign n46666 = ~n46654 & ~n46665;
  assign n46667 = ~pi299 & ~n46666;
  assign n46668 = n38189 & ~n46622;
  assign n46669 = n46667 & ~n46668;
  assign n46670 = pi228 & n46625;
  assign n46671 = ~pi875 & n62380;
  assign n46672 = ~pi166 & ~n62380;
  assign n46673 = ~pi228 & ~n46672;
  assign n46674 = ~pi228 & ~n46671;
  assign n46675 = ~n46672 & n46674;
  assign n46676 = ~n46671 & n46673;
  assign n46677 = ~n46670 & ~n64976;
  assign n46678 = ~pi216 & ~n46677;
  assign n46679 = ~n46613 & ~n46678;
  assign n46680 = ~pi221 & ~n46679;
  assign n46681 = ~n64973 & ~n46680;
  assign n46682 = ~pi215 & ~n46681;
  assign n46683 = ~n46638 & ~n46682;
  assign n46684 = pi299 & ~n46683;
  assign n46685 = ~n46669 & ~n46684;
  assign n46686 = pi39 & ~n46685;
  assign n46687 = ~pi38 & ~n46686;
  assign n46688 = ~n46664 & n46687;
  assign n46689 = pi166 & ~pi228;
  assign n46690 = ~n46670 & ~n46689;
  assign n46691 = ~pi216 & ~n46690;
  assign n46692 = ~n46613 & ~n46691;
  assign n46693 = ~pi221 & ~n46692;
  assign n46694 = ~n64973 & ~n46693;
  assign n46695 = ~pi215 & ~n46694;
  assign n46696 = ~n46638 & ~n46695;
  assign n46697 = pi299 & ~n46696;
  assign n46698 = ~n46669 & ~n46697;
  assign n46699 = pi38 & n46698;
  assign n46700 = ~pi100 & ~n46699;
  assign n46701 = ~n46688 & n46700;
  assign n46702 = ~pi875 & n64892;
  assign n46703 = pi166 & ~n46702;
  assign n46704 = ~n2810 & ~n64892;
  assign n46705 = n2810 & ~n30857;
  assign n46706 = pi875 & ~n46705;
  assign n46707 = ~n46704 & n46706;
  assign n46708 = ~n46703 & ~n46707;
  assign n46709 = ~pi228 & ~n46708;
  assign n46710 = ~n46670 & ~n46709;
  assign n46711 = ~pi216 & ~n46710;
  assign n46712 = ~n46613 & ~n46711;
  assign n46713 = ~pi221 & ~n46712;
  assign n46714 = ~n64973 & ~n46713;
  assign n46715 = ~pi215 & ~n46714;
  assign n46716 = ~n46638 & ~n46715;
  assign n46717 = pi299 & ~n46716;
  assign n46718 = n2764 & ~n46669;
  assign n46719 = ~n46717 & n46718;
  assign n46720 = ~n2764 & n46698;
  assign n46721 = pi100 & ~n46720;
  assign n46722 = ~n46719 & n46721;
  assign n46723 = ~n46701 & ~n46722;
  assign n46724 = ~pi87 & ~n46723;
  assign n46725 = ~n62373 & n46698;
  assign n46726 = n62373 & n46685;
  assign n46727 = ~n46725 & ~n46726;
  assign n46728 = pi87 & n46727;
  assign n46729 = ~pi75 & ~n46728;
  assign n46730 = ~n46724 & n46729;
  assign n46731 = pi75 & n46698;
  assign n46732 = ~pi92 & ~n46731;
  assign n46733 = ~n46730 & n46732;
  assign n46734 = n6795 & ~n46727;
  assign n46735 = ~n6795 & n46698;
  assign n46736 = pi92 & ~n46735;
  assign n46737 = ~n46734 & n46736;
  assign n46738 = n6792 & ~n46737;
  assign n46739 = ~n46733 & n46738;
  assign n46740 = ~n6792 & n46698;
  assign n46741 = ~pi55 & ~n46740;
  assign n46742 = ~n46739 & n46741;
  assign n46743 = n64082 & n46683;
  assign n46744 = ~n64082 & n46696;
  assign n46745 = pi55 & ~n46744;
  assign n46746 = ~n46743 & n46745;
  assign n46747 = ~pi56 & ~n46746;
  assign n46748 = ~n46742 & n46747;
  assign n46749 = n64084 & ~n46683;
  assign n46750 = ~n64084 & ~n46696;
  assign n46751 = pi56 & ~n46750;
  assign n46752 = ~n64084 & n46696;
  assign n46753 = ~pi55 & n46743;
  assign n46754 = ~n46752 & ~n46753;
  assign n46755 = pi56 & ~n46754;
  assign n46756 = ~n46749 & n46751;
  assign n46757 = ~pi62 & ~n64977;
  assign n46758 = ~n46748 & n46757;
  assign n46759 = n44475 & n46683;
  assign n46760 = ~n44475 & n46696;
  assign n46761 = pi62 & ~n46760;
  assign n46762 = ~n46759 & n46761;
  assign n46763 = n3472 & ~n46762;
  assign n46764 = ~n46758 & n46763;
  assign n46765 = ~n3472 & n46696;
  assign n46766 = ~pi245 & ~n46765;
  assign n46767 = ~n46764 & n46766;
  assign n46768 = ~pi166 & ~n43706;
  assign n46769 = pi875 & ~n46768;
  assign n46770 = pi166 & n44316;
  assign n46771 = ~pi166 & ~n44327;
  assign n46772 = ~pi875 & ~n46771;
  assign n46773 = ~n46770 & n46772;
  assign n46774 = ~pi228 & ~n46773;
  assign n46775 = ~pi228 & ~n46769;
  assign n46776 = ~n46773 & n46775;
  assign n46777 = ~n46769 & n46774;
  assign n46778 = n46627 & ~n64978;
  assign n46779 = ~n46613 & ~n46778;
  assign n46780 = ~pi221 & ~n46779;
  assign n46781 = ~n64973 & ~n46780;
  assign n46782 = ~pi215 & ~n46781;
  assign n46783 = n46639 & ~n46782;
  assign n46784 = n46662 & ~n46783;
  assign n46785 = ~n44384 & ~n46670;
  assign n46786 = ~n64976 & n46785;
  assign n46787 = ~pi216 & ~n46786;
  assign n46788 = ~n46613 & ~n46787;
  assign n46789 = ~pi221 & ~n46788;
  assign n46790 = ~n64973 & ~n46789;
  assign n46791 = ~pi215 & ~n46790;
  assign n46792 = ~n46638 & ~n46791;
  assign n46793 = pi299 & ~n46792;
  assign n46794 = ~n46667 & ~n46793;
  assign n46795 = pi39 & ~n46794;
  assign n46796 = ~pi38 & ~n46795;
  assign n46797 = ~n46784 & n46796;
  assign n46798 = ~n44399 & n46696;
  assign n46799 = pi299 & ~n46798;
  assign n46800 = ~n46667 & ~n46799;
  assign n46801 = pi38 & n46800;
  assign n46802 = ~pi100 & ~n46801;
  assign n46803 = ~n46797 & n46802;
  assign n46804 = ~n46709 & n46785;
  assign n46805 = ~pi216 & ~n46804;
  assign n46806 = ~n46613 & ~n46805;
  assign n46807 = ~pi221 & ~n46806;
  assign n46808 = ~n64973 & ~n46807;
  assign n46809 = ~pi215 & ~n46808;
  assign n46810 = ~n46638 & ~n46809;
  assign n46811 = pi299 & ~n46810;
  assign n46812 = n2764 & ~n46667;
  assign n46813 = ~n46811 & n46812;
  assign n46814 = ~n2764 & n46800;
  assign n46815 = pi100 & ~n46814;
  assign n46816 = ~n46813 & n46815;
  assign n46817 = ~n46803 & ~n46816;
  assign n46818 = ~pi87 & ~n46817;
  assign n46819 = ~n62373 & n46800;
  assign n46820 = n62373 & n46794;
  assign n46821 = ~n46819 & ~n46820;
  assign n46822 = pi87 & n46821;
  assign n46823 = ~pi75 & ~n46822;
  assign n46824 = ~n46818 & n46823;
  assign n46825 = pi75 & n46800;
  assign n46826 = ~pi92 & ~n46825;
  assign n46827 = ~n46824 & n46826;
  assign n46828 = n6795 & ~n46821;
  assign n46829 = ~n6795 & n46800;
  assign n46830 = pi92 & ~n46829;
  assign n46831 = ~n46828 & n46830;
  assign n46832 = n6792 & ~n46831;
  assign n46833 = ~n46827 & n46832;
  assign n46834 = ~n6792 & n46800;
  assign n46835 = ~pi55 & ~n46834;
  assign n46836 = ~n46833 & n46835;
  assign n46837 = n64082 & n46792;
  assign n46838 = ~n64082 & n46798;
  assign n46839 = pi55 & ~n46838;
  assign n46840 = ~n46837 & n46839;
  assign n46841 = ~pi56 & ~n46840;
  assign n46842 = ~n46836 & n46841;
  assign n46843 = n64084 & ~n46792;
  assign n46844 = ~n64084 & ~n46798;
  assign n46845 = pi56 & ~n46844;
  assign n46846 = ~pi55 & n46837;
  assign n46847 = ~n64084 & n46798;
  assign n46848 = ~n46846 & ~n46847;
  assign n46849 = pi56 & ~n46848;
  assign n46850 = ~n46843 & n46845;
  assign n46851 = ~pi62 & ~n64979;
  assign n46852 = ~n46842 & n46851;
  assign n46853 = n44475 & n46792;
  assign n46854 = ~n44475 & n46798;
  assign n46855 = pi62 & ~n46854;
  assign n46856 = ~n46853 & n46855;
  assign n46857 = n3472 & ~n46856;
  assign n46858 = ~n46852 & n46857;
  assign n46859 = ~n3472 & n46798;
  assign n46860 = pi245 & ~n46859;
  assign n46861 = ~n46858 & n46860;
  assign n46862 = ~n46767 & ~n46861;
  assign n46863 = ~pi938 & n41020;
  assign n46864 = ~pi1135 & ~n41020;
  assign n46865 = pi221 & ~n46864;
  assign n46866 = pi221 & ~n46863;
  assign n46867 = ~n46864 & n46866;
  assign n46868 = ~n46863 & n46865;
  assign n46869 = pi216 & pi279;
  assign n46870 = ~pi161 & ~n44316;
  assign n46871 = pi161 & n44327;
  assign n46872 = pi879 & ~n46871;
  assign n46873 = ~n46870 & n46872;
  assign n46874 = pi161 & ~pi879;
  assign n46875 = ~n43706 & n46874;
  assign n46876 = ~pi228 & ~n46875;
  assign n46877 = ~n46873 & n46876;
  assign n46878 = pi879 & ~n30613;
  assign n46879 = pi105 & ~n46878;
  assign n46880 = ~pi105 & ~pi161;
  assign n46881 = ~n46879 & ~n46880;
  assign n46882 = n45157 & ~n46881;
  assign n46883 = ~pi216 & ~n46882;
  assign n46884 = ~n44611 & n46883;
  assign n46885 = ~n46873 & ~n46875;
  assign n46886 = ~pi228 & ~n46885;
  assign n46887 = ~n45157 & ~n46886;
  assign n46888 = n46883 & ~n46887;
  assign n46889 = ~n46877 & n46884;
  assign n46890 = ~n46869 & ~n64981;
  assign n46891 = ~pi221 & ~n46890;
  assign n46892 = ~n64980 & ~n46891;
  assign n46893 = ~pi215 & ~n46892;
  assign n46894 = pi215 & pi1135;
  assign n46895 = pi299 & ~n46894;
  assign n46896 = ~n46893 & n46895;
  assign n46897 = pi223 & pi1135;
  assign n46898 = ~pi299 & ~n46897;
  assign n46899 = ~pi938 & n41469;
  assign n46900 = ~pi1135 & ~n41469;
  assign n46901 = pi222 & ~n46900;
  assign n46902 = pi222 & ~n46899;
  assign n46903 = ~n46900 & n46902;
  assign n46904 = ~n46899 & n46901;
  assign n46905 = ~pi224 & ~pi879;
  assign n46906 = ~n30613 & n46905;
  assign n46907 = pi224 & ~pi279;
  assign n46908 = ~pi222 & ~n46907;
  assign n46909 = ~n46906 & n46908;
  assign n46910 = ~n64982 & ~n46909;
  assign n46911 = ~pi223 & ~n46910;
  assign n46912 = ~n46646 & n46911;
  assign n46913 = n46898 & ~n46912;
  assign n46914 = ~pi39 & ~n46913;
  assign n46915 = ~n46896 & n46914;
  assign n46916 = ~n46897 & ~n46911;
  assign n46917 = ~pi299 & ~n46916;
  assign n46918 = n38189 & ~n46878;
  assign n46919 = n46917 & ~n46918;
  assign n46920 = pi228 & n46881;
  assign n46921 = ~pi879 & n62380;
  assign n46922 = pi161 & ~pi228;
  assign n46923 = ~n34059 & ~n46922;
  assign n46924 = ~n46921 & ~n46923;
  assign n46925 = ~n46920 & ~n46924;
  assign n46926 = ~pi216 & ~n46925;
  assign n46927 = ~n46869 & ~n46926;
  assign n46928 = ~pi221 & ~n46927;
  assign n46929 = ~n64980 & ~n46928;
  assign n46930 = ~pi215 & ~n46929;
  assign n46931 = ~n46894 & ~n46930;
  assign n46932 = pi299 & ~n46931;
  assign n46933 = ~n46919 & ~n46932;
  assign n46934 = pi39 & ~n46933;
  assign n46935 = ~pi38 & ~n46934;
  assign n46936 = ~n46915 & n46935;
  assign n46937 = ~n46920 & ~n46922;
  assign n46938 = ~pi216 & ~n46937;
  assign n46939 = ~n46869 & ~n46938;
  assign n46940 = ~pi221 & ~n46939;
  assign n46941 = ~n64980 & ~n46940;
  assign n46942 = ~pi215 & ~n46941;
  assign n46943 = ~n46894 & ~n46942;
  assign n46944 = pi299 & ~n46943;
  assign n46945 = ~n46919 & ~n46944;
  assign n46946 = pi38 & n46945;
  assign n46947 = ~pi100 & ~n46946;
  assign n46948 = ~n46936 & n46947;
  assign n46949 = ~pi879 & n64892;
  assign n46950 = pi161 & ~n46949;
  assign n46951 = ~pi152 & ~pi166;
  assign n46952 = ~n64892 & ~n46951;
  assign n46953 = ~n30857 & n46951;
  assign n46954 = pi879 & ~n46953;
  assign n46955 = ~n46952 & n46954;
  assign n46956 = ~n46950 & ~n46955;
  assign n46957 = ~pi228 & ~n46956;
  assign n46958 = ~n46920 & ~n46957;
  assign n46959 = ~pi216 & ~n46958;
  assign n46960 = ~n46869 & ~n46959;
  assign n46961 = ~pi221 & ~n46960;
  assign n46962 = ~n64980 & ~n46961;
  assign n46963 = ~pi215 & ~n46962;
  assign n46964 = ~n46894 & ~n46963;
  assign n46965 = pi299 & ~n46964;
  assign n46966 = n2764 & ~n46919;
  assign n46967 = ~n46965 & n46966;
  assign n46968 = ~n2764 & n46945;
  assign n46969 = pi100 & ~n46968;
  assign n46970 = ~n46967 & n46969;
  assign n46971 = ~n46948 & ~n46970;
  assign n46972 = ~pi87 & ~n46971;
  assign n46973 = ~n62373 & n46945;
  assign n46974 = n62373 & n46933;
  assign n46975 = ~n46973 & ~n46974;
  assign n46976 = pi87 & n46975;
  assign n46977 = ~pi75 & ~n46976;
  assign n46978 = ~n46972 & n46977;
  assign n46979 = pi75 & n46945;
  assign n46980 = ~pi92 & ~n46979;
  assign n46981 = ~n46978 & n46980;
  assign n46982 = n6795 & ~n46975;
  assign n46983 = ~n6795 & n46945;
  assign n46984 = pi92 & ~n46983;
  assign n46985 = ~n46982 & n46984;
  assign n46986 = n6792 & ~n46985;
  assign n46987 = ~n46981 & n46986;
  assign n46988 = ~n6792 & n46945;
  assign n46989 = ~pi55 & ~n46988;
  assign n46990 = ~n46987 & n46989;
  assign n46991 = n64082 & n46931;
  assign n46992 = ~n64082 & n46943;
  assign n46993 = pi55 & ~n46992;
  assign n46994 = ~n46991 & n46993;
  assign n46995 = ~pi56 & ~n46994;
  assign n46996 = ~n46990 & n46995;
  assign n46997 = n64084 & ~n46931;
  assign n46998 = ~n64084 & ~n46943;
  assign n46999 = pi56 & ~n46998;
  assign n47000 = ~n64084 & n46943;
  assign n47001 = ~pi55 & n46991;
  assign n47002 = ~n47000 & ~n47001;
  assign n47003 = pi56 & ~n47002;
  assign n47004 = ~n46997 & n46999;
  assign n47005 = ~pi62 & ~n64983;
  assign n47006 = ~n46996 & n47005;
  assign n47007 = n44475 & n46931;
  assign n47008 = ~n44475 & n46943;
  assign n47009 = pi62 & ~n47008;
  assign n47010 = ~n47007 & n47009;
  assign n47011 = n3472 & ~n47010;
  assign n47012 = ~n47006 & n47011;
  assign n47013 = ~n3472 & n46943;
  assign n47014 = ~pi244 & ~n47013;
  assign n47015 = ~n47012 & n47014;
  assign n47016 = ~pi161 & ~n43706;
  assign n47017 = pi879 & ~n47016;
  assign n47018 = pi161 & n44316;
  assign n47019 = ~pi161 & ~n44327;
  assign n47020 = ~pi879 & ~n47019;
  assign n47021 = ~n47018 & n47020;
  assign n47022 = ~pi228 & ~n47021;
  assign n47023 = ~pi228 & ~n47017;
  assign n47024 = ~n47021 & n47023;
  assign n47025 = ~n47017 & n47022;
  assign n47026 = n46883 & ~n64984;
  assign n47027 = ~n46869 & ~n47026;
  assign n47028 = ~pi221 & ~n47027;
  assign n47029 = ~n64980 & ~n47028;
  assign n47030 = ~pi215 & ~n47029;
  assign n47031 = n46895 & ~n47030;
  assign n47032 = ~n46646 & n46910;
  assign n47033 = ~pi223 & ~n47032;
  assign n47034 = n46898 & ~n47033;
  assign n47035 = ~pi39 & ~n47034;
  assign n47036 = ~n47031 & n47035;
  assign n47037 = ~n44384 & ~n46920;
  assign n47038 = ~n46924 & n47037;
  assign n47039 = ~pi216 & ~n47038;
  assign n47040 = ~n46869 & ~n47039;
  assign n47041 = ~pi221 & ~n47040;
  assign n47042 = ~n64980 & ~n47041;
  assign n47043 = ~pi215 & ~n47042;
  assign n47044 = ~n46894 & ~n47043;
  assign n47045 = pi299 & ~n47044;
  assign n47046 = ~n46917 & ~n47045;
  assign n47047 = pi39 & ~n47046;
  assign n47048 = ~pi38 & ~n47047;
  assign n47049 = ~n47036 & n47048;
  assign n47050 = ~n44399 & n46943;
  assign n47051 = pi299 & ~n47050;
  assign n47052 = ~n46917 & ~n47051;
  assign n47053 = pi38 & n47052;
  assign n47054 = ~pi100 & ~n47053;
  assign n47055 = ~n47049 & n47054;
  assign n47056 = ~n46957 & n47037;
  assign n47057 = ~pi216 & ~n47056;
  assign n47058 = ~n46869 & ~n47057;
  assign n47059 = ~pi221 & ~n47058;
  assign n47060 = ~n64980 & ~n47059;
  assign n47061 = ~pi215 & ~n47060;
  assign n47062 = ~n46894 & ~n47061;
  assign n47063 = pi299 & ~n47062;
  assign n47064 = n2764 & ~n46917;
  assign n47065 = ~n47063 & n47064;
  assign n47066 = ~n2764 & n47052;
  assign n47067 = pi100 & ~n47066;
  assign n47068 = ~n47065 & n47067;
  assign n47069 = ~n47055 & ~n47068;
  assign n47070 = ~pi87 & ~n47069;
  assign n47071 = ~n62373 & n47052;
  assign n47072 = n62373 & n47046;
  assign n47073 = ~n47071 & ~n47072;
  assign n47074 = pi87 & n47073;
  assign n47075 = ~pi75 & ~n47074;
  assign n47076 = ~n47070 & n47075;
  assign n47077 = pi75 & n47052;
  assign n47078 = ~pi92 & ~n47077;
  assign n47079 = ~n47076 & n47078;
  assign n47080 = n6795 & ~n47073;
  assign n47081 = ~n6795 & n47052;
  assign n47082 = pi92 & ~n47081;
  assign n47083 = ~n47080 & n47082;
  assign n47084 = n6792 & ~n47083;
  assign n47085 = ~n47079 & n47084;
  assign n47086 = ~n6792 & n47052;
  assign n47087 = ~pi55 & ~n47086;
  assign n47088 = ~n47085 & n47087;
  assign n47089 = n64082 & n47044;
  assign n47090 = ~n64082 & n47050;
  assign n47091 = pi55 & ~n47090;
  assign n47092 = ~n47089 & n47091;
  assign n47093 = ~pi56 & ~n47092;
  assign n47094 = ~n47088 & n47093;
  assign n47095 = n64084 & ~n47044;
  assign n47096 = ~n64084 & ~n47050;
  assign n47097 = pi56 & ~n47096;
  assign n47098 = ~pi55 & n47089;
  assign n47099 = ~n64084 & n47050;
  assign n47100 = ~n47098 & ~n47099;
  assign n47101 = pi56 & ~n47100;
  assign n47102 = ~n47095 & n47097;
  assign n47103 = ~pi62 & ~n64985;
  assign n47104 = ~n47094 & n47103;
  assign n47105 = n44475 & n47044;
  assign n47106 = ~n44475 & n47050;
  assign n47107 = pi62 & ~n47106;
  assign n47108 = ~n47105 & n47107;
  assign n47109 = n3472 & ~n47108;
  assign n47110 = ~n47104 & n47109;
  assign n47111 = ~n3472 & n47050;
  assign n47112 = pi244 & ~n47111;
  assign n47113 = ~n47110 & n47112;
  assign n47114 = ~n47015 & ~n47113;
  assign n47115 = pi833 & ~pi930;
  assign n47116 = n2958 & n47115;
  assign n47117 = pi216 & pi278;
  assign n47118 = ~pi221 & ~n47117;
  assign n47119 = ~pi105 & pi152;
  assign n47120 = pi228 & ~n47119;
  assign n47121 = ~pi846 & n44321;
  assign n47122 = pi105 & ~n47121;
  assign n47123 = n47120 & ~n47122;
  assign n47124 = ~pi216 & ~n47123;
  assign n47125 = pi152 & ~n44316;
  assign n47126 = ~pi152 & n44327;
  assign n47127 = ~pi846 & ~n47126;
  assign n47128 = ~n47125 & n47127;
  assign n47129 = ~pi152 & pi846;
  assign n47130 = ~n43706 & n47129;
  assign n47131 = ~n47128 & ~n47130;
  assign n47132 = ~pi228 & ~n47131;
  assign n47133 = n47124 & ~n47132;
  assign n47134 = n47118 & ~n47133;
  assign n47135 = ~n47116 & ~n47134;
  assign n47136 = pi221 & ~n41020;
  assign n47137 = n2959 & ~n47136;
  assign n47138 = n47135 & n47137;
  assign n47139 = pi224 & pi278;
  assign n47140 = ~pi222 & ~n47139;
  assign n47141 = ~pi224 & ~n47121;
  assign n47142 = n47140 & ~n47141;
  assign n47143 = n2978 & n47115;
  assign n47144 = n2979 & ~n41470;
  assign n47145 = ~n47143 & n47144;
  assign n47146 = ~n47142 & ~n47143;
  assign n47147 = n47144 & n47146;
  assign n47148 = ~n47142 & n47145;
  assign n47149 = ~pi39 & ~n64986;
  assign n47150 = ~n47138 & n47149;
  assign n47151 = pi846 & ~n30613;
  assign n47152 = ~pi224 & n47151;
  assign n47153 = n47140 & ~n47152;
  assign n47154 = n41471 & ~n47143;
  assign n47155 = ~n47153 & n47154;
  assign n47156 = ~pi299 & ~n47155;
  assign n47157 = ~n44372 & n47156;
  assign n47158 = ~pi215 & ~n47136;
  assign n47159 = ~n47116 & n47158;
  assign n47160 = pi105 & n47151;
  assign n47161 = ~n47119 & ~n47160;
  assign n47162 = pi228 & ~n47161;
  assign n47163 = ~n44384 & ~n47162;
  assign n47164 = ~pi846 & n62380;
  assign n47165 = ~pi152 & ~n62380;
  assign n47166 = ~pi228 & ~n47165;
  assign n47167 = ~pi228 & ~n47164;
  assign n47168 = ~n47165 & n47167;
  assign n47169 = ~n47164 & n47166;
  assign n47170 = n47163 & ~n64987;
  assign n47171 = ~pi216 & ~n47170;
  assign n47172 = n47118 & ~n47171;
  assign n47173 = n47159 & ~n47172;
  assign n47174 = pi299 & ~n47173;
  assign n47175 = ~n47157 & ~n47174;
  assign n47176 = pi39 & ~n47175;
  assign n47177 = ~pi38 & ~n47176;
  assign n47178 = ~n47150 & n47177;
  assign n47179 = pi152 & ~pi228;
  assign n47180 = ~n47162 & ~n47179;
  assign n47181 = ~pi216 & ~n47180;
  assign n47182 = n47118 & ~n47181;
  assign n47183 = n47159 & ~n47182;
  assign n47184 = ~n44399 & ~n47183;
  assign n47185 = pi299 & n47184;
  assign n47186 = ~n47157 & ~n47185;
  assign n47187 = pi38 & n47186;
  assign n47188 = ~pi100 & ~n47187;
  assign n47189 = ~n47178 & n47188;
  assign n47190 = pi846 & ~n44421;
  assign n47191 = ~n44417 & ~n47190;
  assign n47192 = ~pi228 & ~n47191;
  assign n47193 = n47163 & ~n47192;
  assign n47194 = ~pi216 & ~n47193;
  assign n47195 = n47118 & ~n47194;
  assign n47196 = n47159 & ~n47195;
  assign n47197 = pi299 & ~n47196;
  assign n47198 = n2764 & ~n47157;
  assign n47199 = ~n47197 & n47198;
  assign n47200 = ~n2764 & n47186;
  assign n47201 = pi100 & ~n47200;
  assign n47202 = ~n47199 & n47201;
  assign n47203 = ~n47189 & ~n47202;
  assign n47204 = ~pi87 & ~n47203;
  assign n47205 = ~n62373 & n47186;
  assign n47206 = n62373 & n47175;
  assign n47207 = ~n47205 & ~n47206;
  assign n47208 = pi87 & n47207;
  assign n47209 = ~pi75 & ~n47208;
  assign n47210 = ~n47204 & n47209;
  assign n47211 = pi75 & n47186;
  assign n47212 = ~pi92 & ~n47211;
  assign n47213 = ~n47210 & n47212;
  assign n47214 = n6795 & ~n47207;
  assign n47215 = ~n6795 & n47186;
  assign n47216 = pi92 & ~n47215;
  assign n47217 = ~n47214 & n47216;
  assign n47218 = n6792 & ~n47217;
  assign n47219 = ~n47213 & n47218;
  assign n47220 = ~n6792 & n47186;
  assign n47221 = ~pi55 & ~n47220;
  assign n47222 = ~n47219 & n47221;
  assign n47223 = n64082 & n47173;
  assign n47224 = ~n64082 & ~n47184;
  assign n47225 = pi55 & ~n47224;
  assign n47226 = ~n47223 & n47225;
  assign n47227 = ~pi56 & ~n47226;
  assign n47228 = ~n47222 & n47227;
  assign n47229 = n64084 & ~n47173;
  assign n47230 = ~n64084 & n47184;
  assign n47231 = pi56 & ~n47230;
  assign n47232 = ~n64084 & ~n47184;
  assign n47233 = ~pi55 & n47223;
  assign n47234 = ~n47232 & ~n47233;
  assign n47235 = pi56 & ~n47234;
  assign n47236 = ~n47229 & n47231;
  assign n47237 = ~pi62 & ~n64988;
  assign n47238 = ~n47228 & n47237;
  assign n47239 = n44475 & n47173;
  assign n47240 = ~n44475 & ~n47184;
  assign n47241 = pi62 & ~n47240;
  assign n47242 = ~n47239 & n47241;
  assign n47243 = n3472 & ~n47242;
  assign n47244 = ~n47238 & n47243;
  assign n47245 = ~n3472 & ~n47184;
  assign n47246 = pi242 & ~n47245;
  assign n47247 = ~n47244 & n47246;
  assign n47248 = ~pi152 & ~n44316;
  assign n47249 = pi152 & n44327;
  assign n47250 = pi846 & ~n47249;
  assign n47251 = ~n47248 & n47250;
  assign n47252 = pi152 & ~pi846;
  assign n47253 = ~n43706 & n47252;
  assign n47254 = ~pi228 & ~n47253;
  assign n47255 = ~n47251 & n47254;
  assign n47256 = ~n44321 & n47120;
  assign n47257 = n47124 & ~n47256;
  assign n47258 = ~n47255 & n47257;
  assign n47259 = n47118 & ~n47258;
  assign n47260 = ~n47116 & ~n47259;
  assign n47261 = n47137 & n47260;
  assign n47262 = ~n44320 & n47152;
  assign n47263 = n47140 & ~n47262;
  assign n47264 = n47145 & ~n47263;
  assign n47265 = ~pi39 & ~n47264;
  assign n47266 = ~n47261 & n47265;
  assign n47267 = ~n47162 & ~n64987;
  assign n47268 = ~pi216 & ~n47267;
  assign n47269 = n47118 & ~n47268;
  assign n47270 = n47159 & ~n47269;
  assign n47271 = pi299 & ~n47270;
  assign n47272 = ~n47156 & ~n47271;
  assign n47273 = pi39 & ~n47272;
  assign n47274 = ~pi38 & ~n47273;
  assign n47275 = ~n47266 & n47274;
  assign n47276 = pi299 & ~n47183;
  assign n47277 = ~n47156 & ~n47276;
  assign n47278 = pi38 & n47277;
  assign n47279 = ~pi100 & ~n47278;
  assign n47280 = ~n47275 & n47279;
  assign n47281 = ~n47162 & ~n47192;
  assign n47282 = ~pi216 & ~n47281;
  assign n47283 = n47118 & ~n47282;
  assign n47284 = n47159 & ~n47283;
  assign n47285 = pi299 & ~n47284;
  assign n47286 = n2764 & ~n47156;
  assign n47287 = ~n47285 & n47286;
  assign n47288 = ~n2764 & n47277;
  assign n47289 = pi100 & ~n47288;
  assign n47290 = ~n47287 & n47289;
  assign n47291 = ~n47280 & ~n47290;
  assign n47292 = ~pi87 & ~n47291;
  assign n47293 = ~n62373 & n47277;
  assign n47294 = n62373 & n47272;
  assign n47295 = ~n47293 & ~n47294;
  assign n47296 = pi87 & n47295;
  assign n47297 = ~pi75 & ~n47296;
  assign n47298 = ~n47292 & n47297;
  assign n47299 = pi75 & n47277;
  assign n47300 = ~pi92 & ~n47299;
  assign n47301 = ~n47298 & n47300;
  assign n47302 = n6795 & ~n47295;
  assign n47303 = ~n6795 & n47277;
  assign n47304 = pi92 & ~n47303;
  assign n47305 = ~n47302 & n47304;
  assign n47306 = n6792 & ~n47305;
  assign n47307 = ~n47301 & n47306;
  assign n47308 = ~n6792 & n47277;
  assign n47309 = ~pi55 & ~n47308;
  assign n47310 = ~n47307 & n47309;
  assign n47311 = n64082 & n47270;
  assign n47312 = ~n64082 & n47183;
  assign n47313 = pi55 & ~n47312;
  assign n47314 = ~n47311 & n47313;
  assign n47315 = ~pi56 & ~n47314;
  assign n47316 = ~n47310 & n47315;
  assign n47317 = n64084 & ~n47270;
  assign n47318 = ~n64084 & ~n47183;
  assign n47319 = pi56 & ~n47318;
  assign n47320 = ~n64084 & n47183;
  assign n47321 = ~pi55 & n47311;
  assign n47322 = ~n47320 & ~n47321;
  assign n47323 = pi56 & ~n47322;
  assign n47324 = ~n47317 & n47319;
  assign n47325 = ~pi62 & ~n64989;
  assign n47326 = ~n47316 & n47325;
  assign n47327 = n44475 & n47270;
  assign n47328 = ~n44475 & n47183;
  assign n47329 = pi62 & ~n47328;
  assign n47330 = ~n47327 & n47329;
  assign n47331 = n3472 & ~n47330;
  assign n47332 = ~n47326 & n47331;
  assign n47333 = ~n3472 & n47183;
  assign n47334 = ~pi242 & ~n47333;
  assign n47335 = ~n47332 & n47334;
  assign n47336 = ~n47247 & ~n47335;
  assign n47337 = ~pi1134 & ~n47336;
  assign n47338 = n2979 & ~n47146;
  assign n47339 = ~pi39 & ~n47338;
  assign n47340 = n2959 & ~n47135;
  assign n47341 = n47339 & ~n47340;
  assign n47342 = n41471 & n47157;
  assign n47343 = ~pi299 & ~n47342;
  assign n47344 = ~n47116 & ~n47172;
  assign n47345 = ~pi215 & ~n47344;
  assign n47346 = pi299 & ~n47345;
  assign n47347 = ~n47343 & ~n47346;
  assign n47348 = pi39 & ~n47347;
  assign n47349 = ~pi38 & ~n47348;
  assign n47350 = ~n47341 & n47349;
  assign n47351 = ~n47116 & ~n47182;
  assign n47352 = ~pi215 & ~n47351;
  assign n47353 = ~n44399 & n47352;
  assign n47354 = pi299 & ~n47353;
  assign n47355 = ~n47343 & ~n47354;
  assign n47356 = pi38 & n47355;
  assign n47357 = ~pi100 & ~n47356;
  assign n47358 = ~n47350 & n47357;
  assign n47359 = ~n47116 & ~n47195;
  assign n47360 = ~pi215 & ~n47359;
  assign n47361 = pi299 & ~n47360;
  assign n47362 = n2764 & ~n47343;
  assign n47363 = ~n47361 & n47362;
  assign n47364 = ~n2764 & n47355;
  assign n47365 = pi100 & ~n47364;
  assign n47366 = ~n47363 & n47365;
  assign n47367 = ~n47358 & ~n47366;
  assign n47368 = ~pi87 & ~n47367;
  assign n47369 = ~n62373 & n47355;
  assign n47370 = n62373 & n47347;
  assign n47371 = ~n47369 & ~n47370;
  assign n47372 = pi87 & n47371;
  assign n47373 = ~pi75 & ~n47372;
  assign n47374 = ~n47368 & n47373;
  assign n47375 = pi75 & n47355;
  assign n47376 = ~pi92 & ~n47375;
  assign n47377 = ~n47374 & n47376;
  assign n47378 = n6795 & ~n47371;
  assign n47379 = ~n6795 & n47355;
  assign n47380 = pi92 & ~n47379;
  assign n47381 = ~n47378 & n47380;
  assign n47382 = n6792 & ~n47381;
  assign n47383 = ~n47377 & n47382;
  assign n47384 = ~n6792 & n47355;
  assign n47385 = ~pi55 & ~n47384;
  assign n47386 = ~n47383 & n47385;
  assign n47387 = n64082 & n47345;
  assign n47388 = ~n64082 & n47353;
  assign n47389 = pi55 & ~n47388;
  assign n47390 = ~n47387 & n47389;
  assign n47391 = ~pi56 & ~n47390;
  assign n47392 = ~n47386 & n47391;
  assign n47393 = n64084 & ~n47345;
  assign n47394 = ~n64084 & ~n47353;
  assign n47395 = pi56 & ~n47394;
  assign n47396 = ~pi55 & n47387;
  assign n47397 = ~n64084 & n47353;
  assign n47398 = ~n47396 & ~n47397;
  assign n47399 = pi56 & ~n47398;
  assign n47400 = ~n47393 & n47395;
  assign n47401 = ~pi62 & ~n64990;
  assign n47402 = ~n47392 & n47401;
  assign n47403 = n44475 & n47345;
  assign n47404 = ~n44475 & n47353;
  assign n47405 = pi62 & ~n47404;
  assign n47406 = ~n47403 & n47405;
  assign n47407 = n3472 & ~n47406;
  assign n47408 = ~n47402 & n47407;
  assign n47409 = ~n3472 & n47353;
  assign n47410 = pi242 & ~n47409;
  assign n47411 = ~n47408 & n47410;
  assign n47412 = n2959 & ~n47260;
  assign n47413 = n2979 & n47263;
  assign n47414 = n47339 & ~n47413;
  assign n47415 = ~n47412 & n47414;
  assign n47416 = ~pi223 & n47153;
  assign n47417 = n47343 & ~n47416;
  assign n47418 = ~n47116 & ~n47269;
  assign n47419 = ~pi215 & ~n47418;
  assign n47420 = pi299 & ~n47419;
  assign n47421 = ~n47417 & ~n47420;
  assign n47422 = pi39 & ~n47421;
  assign n47423 = ~pi38 & ~n47422;
  assign n47424 = ~n47415 & n47423;
  assign n47425 = pi299 & ~n47352;
  assign n47426 = ~n47417 & ~n47425;
  assign n47427 = pi38 & n47426;
  assign n47428 = ~pi100 & ~n47427;
  assign n47429 = ~n47424 & n47428;
  assign n47430 = ~n47116 & ~n47283;
  assign n47431 = ~pi215 & ~n47430;
  assign n47432 = pi299 & ~n47431;
  assign n47433 = n2764 & ~n47417;
  assign n47434 = ~n47432 & n47433;
  assign n47435 = ~n2764 & n47426;
  assign n47436 = pi100 & ~n47435;
  assign n47437 = ~n47434 & n47436;
  assign n47438 = ~n47429 & ~n47437;
  assign n47439 = ~pi87 & ~n47438;
  assign n47440 = ~n62373 & n47426;
  assign n47441 = n62373 & n47421;
  assign n47442 = ~n47440 & ~n47441;
  assign n47443 = pi87 & n47442;
  assign n47444 = ~pi75 & ~n47443;
  assign n47445 = ~n47439 & n47444;
  assign n47446 = pi75 & n47426;
  assign n47447 = ~pi92 & ~n47446;
  assign n47448 = ~n47445 & n47447;
  assign n47449 = n6795 & ~n47442;
  assign n47450 = ~n6795 & n47426;
  assign n47451 = pi92 & ~n47450;
  assign n47452 = ~n47449 & n47451;
  assign n47453 = n6792 & ~n47452;
  assign n47454 = ~n47448 & n47453;
  assign n47455 = ~n6792 & n47426;
  assign n47456 = ~pi55 & ~n47455;
  assign n47457 = ~n47454 & n47456;
  assign n47458 = n64082 & n47419;
  assign n47459 = ~n64082 & n47352;
  assign n47460 = pi55 & ~n47459;
  assign n47461 = ~n47458 & n47460;
  assign n47462 = ~pi56 & ~n47461;
  assign n47463 = ~n47457 & n47462;
  assign n47464 = n64084 & ~n47419;
  assign n47465 = ~n64084 & ~n47352;
  assign n47466 = pi56 & ~n47465;
  assign n47467 = ~n64084 & n47352;
  assign n47468 = ~pi55 & n47458;
  assign n47469 = ~n47467 & ~n47468;
  assign n47470 = pi56 & ~n47469;
  assign n47471 = ~n47464 & n47466;
  assign n47472 = ~pi62 & ~n64991;
  assign n47473 = ~n47463 & n47472;
  assign n47474 = n44475 & n47419;
  assign n47475 = ~n44475 & n47352;
  assign n47476 = pi62 & ~n47475;
  assign n47477 = ~n47474 & n47476;
  assign n47478 = n3472 & ~n47477;
  assign n47479 = ~n47473 & n47478;
  assign n47480 = ~n3472 & n47352;
  assign n47481 = ~pi242 & ~n47480;
  assign n47482 = ~n47479 & n47481;
  assign n47483 = pi1134 & ~n47482;
  assign n47484 = ~n47411 & n47483;
  assign po165 = ~n47337 & ~n47484;
  assign n47486 = ~pi39 & ~n41912;
  assign n47487 = pi39 & ~n42562;
  assign n47488 = n2766 & ~n47487;
  assign n47489 = ~n47486 & n47488;
  assign n47490 = ~n43148 & ~n47489;
  assign n47491 = ~pi87 & ~n47490;
  assign n47492 = n64706 & ~n47491;
  assign n47493 = ~n64706 & ~n41788;
  assign n47494 = n41783 & ~n47493;
  assign n47495 = n41782 & n41783;
  assign n47496 = ~n47493 & n47495;
  assign n47497 = n41782 & n47494;
  assign n47498 = ~n64706 & n41788;
  assign n47499 = n6796 & n35113;
  assign n47500 = ~n47490 & n47499;
  assign n47501 = ~n47498 & ~n47500;
  assign n47502 = n47495 & ~n47501;
  assign n47503 = ~n47492 & n64992;
  assign n47504 = ~pi72 & n64082;
  assign n47505 = n64082 & ~n39223;
  assign n47506 = ~n39190 & n47504;
  assign n47507 = ~n3036 & n64994;
  assign n47508 = pi286 & n47507;
  assign n47509 = pi288 & pi289;
  assign n47510 = n47508 & n47509;
  assign n47511 = pi285 & n64994;
  assign n47512 = ~n47510 & ~n47511;
  assign n47513 = pi285 & n47510;
  assign n47514 = n62455 & ~n47513;
  assign n47515 = n62455 & ~n47512;
  assign n47516 = ~n47513 & n47515;
  assign n47517 = ~n47512 & n47514;
  assign n47518 = n62455 & n47510;
  assign n47519 = ~pi286 & n3036;
  assign n47520 = ~pi288 & n47519;
  assign n47521 = ~pi289 & n47520;
  assign n47522 = pi285 & ~n47521;
  assign n47523 = ~n47518 & n47522;
  assign n47524 = ~n64995 & ~n47523;
  assign po442 = ~pi793 & ~n47524;
  assign n47526 = ~pi288 & ~n3317;
  assign n47527 = n3036 & ~n64994;
  assign n47528 = pi286 & ~n47527;
  assign n47529 = ~n64994 & n47519;
  assign n47530 = ~n47528 & ~n47529;
  assign n47531 = n47526 & ~n47530;
  assign n47532 = ~pi286 & ~n47507;
  assign n47533 = pi288 & ~n47508;
  assign n47534 = ~n47532 & n47533;
  assign n47535 = n62455 & ~n47534;
  assign n47536 = n62455 & ~n47531;
  assign n47537 = ~n47534 & n47536;
  assign n47538 = ~n47531 & n47535;
  assign n47539 = n3036 & n47526;
  assign n47540 = ~pi286 & n47539;
  assign n47541 = pi286 & ~n47539;
  assign n47542 = ~n62455 & ~n47541;
  assign n47543 = ~n62455 & ~n47540;
  assign n47544 = ~n47541 & n47543;
  assign n47545 = ~n47540 & n47542;
  assign n47546 = ~pi793 & ~n64997;
  assign po443 = ~n64996 & n47546;
  assign n47548 = pi288 & ~n3036;
  assign n47549 = ~n47539 & ~n47548;
  assign n47550 = ~n39223 & n64705;
  assign n47551 = n62455 & n64994;
  assign n47552 = ~n47549 & po637;
  assign n47553 = n47549 & ~po637;
  assign n47554 = ~pi793 & ~n47553;
  assign n47555 = ~pi793 & ~n47552;
  assign n47556 = ~n47553 & n47555;
  assign n47557 = ~n47552 & n47554;
  assign n47558 = pi289 & ~n47529;
  assign n47559 = pi285 & ~pi289;
  assign n47560 = n47529 & n47559;
  assign n47561 = ~pi288 & ~n47560;
  assign n47562 = ~pi288 & ~n47558;
  assign n47563 = ~n47560 & n47562;
  assign n47564 = ~n47558 & n47561;
  assign n47565 = ~pi289 & n47533;
  assign n47566 = ~n47510 & ~n47565;
  assign n47567 = ~n47510 & ~n65000;
  assign n47568 = ~n47565 & n47567;
  assign n47569 = ~n65000 & n47566;
  assign n47570 = n62455 & ~n65001;
  assign n47571 = n47520 & n47559;
  assign n47572 = pi289 & ~n47520;
  assign n47573 = ~n62455 & ~n47572;
  assign n47574 = ~n62455 & ~n47571;
  assign n47575 = ~n47572 & n47574;
  assign n47576 = ~n47571 & n47573;
  assign n47577 = ~pi793 & ~n65002;
  assign po446 = ~n47570 & n47577;
  assign n47579 = pi233 & pi237;
  assign n47580 = ~pi332 & ~n2904;
  assign n47581 = ~pi947 & ~n47580;
  assign n47582 = pi96 & pi210;
  assign n47583 = pi332 & n47582;
  assign n47584 = ~pi32 & pi70;
  assign n47585 = ~pi70 & ~pi841;
  assign n47586 = pi32 & n47585;
  assign n47587 = ~n47584 & ~n47586;
  assign n47588 = ~pi210 & ~n47587;
  assign n47589 = ~pi32 & ~pi96;
  assign n47590 = pi70 & n47589;
  assign n47591 = ~pi332 & ~n47590;
  assign n47592 = ~n47588 & n47591;
  assign n47593 = ~n47583 & ~n47592;
  assign n47594 = ~n2814 & n47593;
  assign n47595 = n2904 & ~n47594;
  assign n47596 = n47581 & ~n47595;
  assign n47597 = pi332 & pi468;
  assign n47598 = ~pi468 & ~n47592;
  assign n47599 = ~n47597 & ~n47598;
  assign n47600 = ~n2904 & n47599;
  assign n47601 = n2904 & ~n47593;
  assign n47602 = pi947 & ~n47601;
  assign n47603 = ~n47600 & n47602;
  assign n47604 = ~n47596 & ~n47603;
  assign n47605 = ~n64082 & n47604;
  assign n47606 = ~pi95 & n64731;
  assign n47607 = ~pi70 & ~n47606;
  assign n47608 = n47589 & ~n47607;
  assign n47609 = pi210 & n47608;
  assign n47610 = ~pi95 & n2726;
  assign n47611 = pi32 & ~n47585;
  assign n47612 = ~pi96 & ~n47611;
  assign n47613 = ~pi95 & n2730;
  assign n47614 = ~n47611 & n47613;
  assign n47615 = n47610 & n47612;
  assign n47616 = n6829 & n65003;
  assign n47617 = n62363 & n47616;
  assign n47618 = n47587 & ~n47617;
  assign n47619 = ~pi210 & ~n47618;
  assign n47620 = ~pi332 & ~n47619;
  assign n47621 = ~n47609 & n47620;
  assign n47622 = ~n47583 & ~n47621;
  assign n47623 = ~n2814 & n47622;
  assign n47624 = n2904 & ~n47623;
  assign n47625 = n47581 & ~n47624;
  assign n47626 = ~pi468 & ~n47621;
  assign n47627 = ~n47597 & ~n47626;
  assign n47628 = ~n2904 & n47627;
  assign n47629 = n2904 & ~n47622;
  assign n47630 = pi947 & ~n47629;
  assign n47631 = ~n47628 & n47630;
  assign n47632 = ~n47625 & ~n47631;
  assign n47633 = n64082 & n47632;
  assign n47634 = ~n47605 & ~n47633;
  assign n47635 = n3471 & ~n47634;
  assign n47636 = ~n3471 & n47604;
  assign n47637 = pi59 & ~n47636;
  assign n47638 = ~n47635 & n47637;
  assign n47639 = n2743 & n41093;
  assign n47640 = n47610 & n47639;
  assign n47641 = ~pi70 & ~n47640;
  assign n47642 = n47589 & ~n47641;
  assign n47643 = pi210 & n47642;
  assign n47644 = n65003 & n47639;
  assign n47645 = n47587 & ~n47644;
  assign n47646 = ~pi210 & ~n47645;
  assign n47647 = ~pi332 & ~n47646;
  assign n47648 = ~n47643 & n47647;
  assign n47649 = ~pi468 & ~n47648;
  assign n47650 = ~n47597 & ~n47649;
  assign n47651 = pi947 & ~n47650;
  assign n47652 = pi332 & ~pi947;
  assign n47653 = ~n2904 & ~n47652;
  assign n47654 = ~n47651 & n47653;
  assign n47655 = ~n47583 & ~n47648;
  assign n47656 = n2904 & ~n47655;
  assign n47657 = pi299 & ~n34208;
  assign n47658 = ~n47656 & n47657;
  assign n47659 = ~n47654 & n47658;
  assign n47660 = pi198 & n47642;
  assign n47661 = ~pi198 & ~n47645;
  assign n47662 = ~pi332 & ~n47661;
  assign n47663 = ~n47660 & n47662;
  assign n47664 = ~pi468 & ~n47663;
  assign n47665 = ~n2904 & ~n47597;
  assign n47666 = ~n47664 & n47665;
  assign n47667 = pi587 & ~n47666;
  assign n47668 = pi468 & n2904;
  assign n47669 = ~pi332 & ~n47668;
  assign n47670 = ~pi587 & ~n47669;
  assign n47671 = ~n47667 & ~n47670;
  assign n47672 = pi96 & pi198;
  assign n47673 = pi332 & n47672;
  assign n47674 = ~n47663 & ~n47673;
  assign n47675 = n2904 & ~n47674;
  assign n47676 = ~pi299 & ~n47675;
  assign n47677 = ~n47671 & n47676;
  assign n47678 = n64086 & ~n47677;
  assign n47679 = ~n2814 & n47655;
  assign n47680 = n2904 & ~n47679;
  assign n47681 = n47581 & ~n47680;
  assign n47682 = ~n2904 & n47650;
  assign n47683 = pi947 & ~n47656;
  assign n47684 = ~n47682 & n47683;
  assign n47685 = pi299 & ~n47684;
  assign n47686 = pi299 & ~n47681;
  assign n47687 = ~n47684 & n47686;
  assign n47688 = ~n47681 & n47685;
  assign n47689 = ~pi587 & ~n47580;
  assign n47690 = ~n2814 & n47674;
  assign n47691 = n2904 & ~n47690;
  assign n47692 = n47689 & ~n47691;
  assign n47693 = pi587 & ~n47675;
  assign n47694 = ~n47666 & n47693;
  assign n47695 = n47667 & ~n47675;
  assign n47696 = ~pi299 & ~n65005;
  assign n47697 = ~n47671 & ~n47675;
  assign n47698 = ~pi299 & ~n47697;
  assign n47699 = ~pi299 & ~n47692;
  assign n47700 = ~n65005 & n47699;
  assign n47701 = ~n47692 & n47696;
  assign n47702 = ~n65004 & ~n65006;
  assign n47703 = n64086 & ~n47702;
  assign n47704 = ~n47659 & n47678;
  assign n47705 = pi299 & ~n47632;
  assign n47706 = pi198 & n47608;
  assign n47707 = ~pi198 & ~n47618;
  assign n47708 = ~pi332 & ~n47707;
  assign n47709 = ~n47706 & n47708;
  assign n47710 = ~pi468 & ~n47709;
  assign n47711 = n47665 & ~n47710;
  assign n47712 = pi587 & ~n47711;
  assign n47713 = ~n47670 & ~n47712;
  assign n47714 = ~n47673 & ~n47709;
  assign n47715 = n2904 & ~n47714;
  assign n47716 = ~pi299 & ~n47715;
  assign n47717 = ~n2814 & n47714;
  assign n47718 = n2904 & ~n47717;
  assign n47719 = n47689 & ~n47718;
  assign n47720 = pi587 & ~n47715;
  assign n47721 = ~n47711 & n47720;
  assign n47722 = n47712 & ~n47715;
  assign n47723 = ~n47719 & ~n65008;
  assign n47724 = ~pi299 & ~n47723;
  assign n47725 = ~n47713 & n47716;
  assign n47726 = n43656 & ~n65009;
  assign n47727 = n43656 & ~n47705;
  assign n47728 = ~n65009 & n47727;
  assign n47729 = ~n47705 & n47726;
  assign n47730 = ~n65007 & ~n65010;
  assign n47731 = ~pi74 & ~n47730;
  assign n47732 = pi299 & ~n47604;
  assign n47733 = ~pi74 & n64081;
  assign n47734 = ~pi198 & ~n47587;
  assign n47735 = n47591 & ~n47734;
  assign n47736 = ~n47673 & ~n47735;
  assign n47737 = n2904 & ~n47736;
  assign n47738 = n34213 & ~n47735;
  assign n47739 = n47580 & ~n47738;
  assign n47740 = ~pi299 & ~n34212;
  assign n47741 = ~n47739 & n47740;
  assign n47742 = ~n47737 & n47740;
  assign n47743 = ~n47739 & n47742;
  assign n47744 = ~n47737 & n47741;
  assign n47745 = ~n47733 & ~n65011;
  assign n47746 = ~n47732 & n47745;
  assign n47747 = ~pi55 & ~n47746;
  assign n47748 = ~n47731 & n47747;
  assign n47749 = pi55 & n47634;
  assign n47750 = n3470 & ~n47749;
  assign n47751 = ~n47748 & n47750;
  assign n47752 = ~n3470 & n47604;
  assign n47753 = ~pi59 & ~n47752;
  assign n47754 = ~n47751 & n47753;
  assign n47755 = ~n47638 & ~n47754;
  assign n47756 = ~pi57 & ~n47755;
  assign n47757 = pi57 & ~n47604;
  assign n47758 = ~n47756 & ~n47757;
  assign n47759 = n47579 & ~n47758;
  assign n47760 = pi57 & pi332;
  assign n47761 = pi332 & ~n3470;
  assign n47762 = ~pi59 & ~n47761;
  assign n47763 = pi74 & pi332;
  assign n47764 = ~pi55 & ~n47763;
  assign n47765 = ~pi299 & pi587;
  assign n47766 = ~n35595 & ~n47765;
  assign n47767 = ~pi468 & ~n47766;
  assign n47768 = pi468 & ~n2904;
  assign n47769 = ~pi468 & ~n35595;
  assign n47770 = ~n47765 & n47769;
  assign n47771 = ~n47768 & ~n47770;
  assign n47772 = ~n47668 & ~n47767;
  assign n47773 = n35400 & n41093;
  assign n47774 = n65012 & n47773;
  assign n47775 = ~pi332 & ~n47774;
  assign n47776 = n64086 & ~n47775;
  assign n47777 = n62380 & n34256;
  assign n47778 = ~pi332 & ~n47777;
  assign n47779 = n43656 & ~n47778;
  assign n47780 = pi332 & ~n64081;
  assign n47781 = ~n47779 & ~n47780;
  assign n47782 = ~n47776 & n47781;
  assign n47783 = ~pi74 & ~n47782;
  assign n47784 = n47764 & ~n47783;
  assign n47785 = n64082 & n34209;
  assign n47786 = n64109 & n34209;
  assign n47787 = n62380 & n47785;
  assign n47788 = ~pi332 & ~n65013;
  assign n47789 = pi55 & n47788;
  assign n47790 = n3470 & ~n47789;
  assign n47791 = ~n47784 & n47790;
  assign n47792 = n47762 & ~n47791;
  assign n47793 = n3471 & ~n47788;
  assign n47794 = pi332 & ~n3471;
  assign n47795 = pi59 & ~n47794;
  assign n47796 = ~n47793 & n47795;
  assign n47797 = ~pi57 & ~n47796;
  assign n47798 = ~n47792 & n47797;
  assign n47799 = ~n47760 & ~n47798;
  assign n47800 = ~n47579 & ~n47799;
  assign n47801 = ~n47759 & ~n47800;
  assign n47802 = ~pi201 & ~n47801;
  assign n47803 = ~pi299 & n3475;
  assign n47804 = ~pi57 & n47803;
  assign n47805 = ~pi299 & n62455;
  assign n47806 = n34213 & n47672;
  assign n47807 = n65014 & ~n47806;
  assign n47808 = ~n34209 & ~n65014;
  assign n47809 = ~n47582 & ~n65014;
  assign n47810 = ~n47808 & ~n47809;
  assign n47811 = ~n47807 & ~n47809;
  assign n47812 = ~n47808 & n47811;
  assign n47813 = ~n47807 & ~n47808;
  assign n47814 = ~n47809 & n47813;
  assign n47815 = ~n47807 & n47810;
  assign n47816 = n47579 & n65015;
  assign n47817 = pi201 & ~n47816;
  assign po358 = ~n47802 & ~n47817;
  assign n47819 = ~pi233 & pi237;
  assign n47820 = ~n47758 & n47819;
  assign n47821 = ~n47799 & ~n47819;
  assign n47822 = ~n47820 & ~n47821;
  assign n47823 = ~pi202 & ~n47822;
  assign n47824 = n65015 & n47819;
  assign n47825 = pi202 & ~n47824;
  assign po359 = ~n47823 & ~n47825;
  assign n47827 = ~pi233 & ~pi237;
  assign n47828 = ~n47758 & n47827;
  assign n47829 = ~n47799 & ~n47827;
  assign n47830 = ~n47828 & ~n47829;
  assign n47831 = ~pi203 & ~n47830;
  assign n47832 = n65015 & n47827;
  assign n47833 = pi203 & ~n47832;
  assign po360 = ~n47831 & ~n47833;
  assign n47835 = ~pi332 & ~n2907;
  assign n47836 = ~pi907 & ~n47835;
  assign n47837 = n2907 & ~n47594;
  assign n47838 = n47836 & ~n47837;
  assign n47839 = ~n2907 & n47599;
  assign n47840 = n2907 & ~n47593;
  assign n47841 = pi907 & ~n47840;
  assign n47842 = ~n47839 & n47841;
  assign n47843 = ~n47838 & ~n47842;
  assign n47844 = ~n64082 & n47843;
  assign n47845 = ~n2907 & n47627;
  assign n47846 = n2907 & ~n47622;
  assign n47847 = pi907 & ~n47846;
  assign n47848 = ~n47845 & n47847;
  assign n47849 = pi332 & ~n7008;
  assign n47850 = pi680 & ~n47849;
  assign n47851 = ~n47623 & n47850;
  assign n47852 = n47836 & ~n47851;
  assign n47853 = ~n47848 & ~n47852;
  assign n47854 = n64082 & n47853;
  assign n47855 = ~n47844 & ~n47854;
  assign n47856 = n3471 & ~n47855;
  assign n47857 = ~n3471 & n47843;
  assign n47858 = pi59 & ~n47857;
  assign n47859 = ~n47856 & n47858;
  assign n47860 = pi299 & n47853;
  assign n47861 = n34078 & n47714;
  assign n47862 = n2907 & n47672;
  assign n47863 = pi332 & ~n47862;
  assign n47864 = ~pi299 & ~n47863;
  assign n47865 = ~n47861 & n47864;
  assign n47866 = ~n47860 & ~n47865;
  assign n47867 = n43656 & ~n47866;
  assign n47868 = n34078 & n47674;
  assign n47869 = n47864 & ~n47868;
  assign n47870 = pi907 & ~n47650;
  assign n47871 = pi332 & ~pi907;
  assign n47872 = ~n2907 & ~n47871;
  assign n47873 = ~n47870 & n47872;
  assign n47874 = n2907 & ~n47655;
  assign n47875 = ~n34056 & ~n47874;
  assign n47876 = ~n47873 & n47875;
  assign n47877 = ~n2907 & n47650;
  assign n47878 = pi907 & ~n47874;
  assign n47879 = ~n47877 & n47878;
  assign n47880 = n2907 & ~n47679;
  assign n47881 = n47836 & ~n47880;
  assign n47882 = pi299 & ~n47881;
  assign n47883 = ~n47879 & n47882;
  assign n47884 = pi299 & ~n47879;
  assign n47885 = ~n47881 & n47884;
  assign n47886 = pi299 & ~n47876;
  assign n47887 = ~n47869 & ~n65016;
  assign n47888 = n64086 & ~n47887;
  assign n47889 = ~n47867 & ~n47888;
  assign n47890 = ~pi74 & ~n47889;
  assign n47891 = pi299 & ~n47843;
  assign n47892 = ~pi468 & pi602;
  assign n47893 = pi468 & n2907;
  assign n47894 = ~n47892 & ~n47893;
  assign n47895 = n47736 & ~n47894;
  assign n47896 = ~n47863 & ~n47895;
  assign n47897 = ~pi299 & ~n47896;
  assign n47898 = ~n47733 & ~n47897;
  assign n47899 = ~n47891 & n47898;
  assign n47900 = ~pi55 & ~n47899;
  assign n47901 = ~n47890 & n47900;
  assign n47902 = pi55 & n47855;
  assign n47903 = n3470 & ~n47902;
  assign n47904 = ~n47901 & n47903;
  assign n47905 = ~n3470 & n47843;
  assign n47906 = ~pi59 & ~n47905;
  assign n47907 = ~n47904 & n47906;
  assign n47908 = ~n47859 & ~n47907;
  assign n47909 = ~pi57 & ~n47908;
  assign n47910 = pi57 & ~n47843;
  assign n47911 = ~n47909 & ~n47910;
  assign n47912 = n47579 & ~n47911;
  assign n47913 = ~pi299 & ~n47894;
  assign n47914 = ~n34127 & ~n47913;
  assign n47915 = n62380 & ~n47914;
  assign n47916 = ~pi332 & ~n47915;
  assign n47917 = n43656 & ~n47916;
  assign n47918 = pi299 & ~pi907;
  assign n47919 = ~pi299 & ~pi602;
  assign n47920 = ~pi468 & ~n47919;
  assign n47921 = ~pi468 & ~n47918;
  assign n47922 = ~n47919 & n47921;
  assign n47923 = ~n47918 & n47920;
  assign n47924 = ~n47893 & ~n65017;
  assign n47925 = n47773 & ~n47924;
  assign n47926 = ~pi332 & ~n47925;
  assign n47927 = n64086 & ~n47926;
  assign n47928 = ~n47917 & ~n47927;
  assign n47929 = ~pi74 & ~n47928;
  assign n47930 = n47764 & ~n47780;
  assign n47931 = ~n47929 & n47930;
  assign n47932 = n64082 & n34057;
  assign n47933 = n64109 & n34057;
  assign n47934 = n62380 & n47932;
  assign n47935 = ~pi332 & ~n65018;
  assign n47936 = pi55 & n47935;
  assign n47937 = n3470 & ~n47936;
  assign n47938 = ~n47931 & n47937;
  assign n47939 = n47762 & ~n47938;
  assign n47940 = n3471 & ~n47935;
  assign n47941 = n47795 & ~n47940;
  assign n47942 = ~pi57 & ~n47941;
  assign n47943 = ~n47939 & n47942;
  assign n47944 = ~n47760 & ~n47943;
  assign n47945 = ~n47579 & ~n47944;
  assign n47946 = ~n47912 & ~n47945;
  assign n47947 = ~pi204 & ~n47946;
  assign n47948 = n34078 & n47672;
  assign n47949 = n65014 & ~n47948;
  assign n47950 = ~n34057 & ~n65014;
  assign n47951 = ~n47809 & ~n47950;
  assign n47952 = ~n47949 & n47951;
  assign n47953 = n47579 & n47952;
  assign n47954 = pi204 & ~n47953;
  assign po361 = ~n47947 & ~n47954;
  assign n47956 = n47819 & ~n47911;
  assign n47957 = ~n47819 & ~n47944;
  assign n47958 = ~n47956 & ~n47957;
  assign n47959 = ~pi205 & ~n47958;
  assign n47960 = n47819 & n47952;
  assign n47961 = pi205 & ~n47960;
  assign po362 = ~n47959 & ~n47961;
  assign n47963 = pi233 & ~pi237;
  assign n47964 = ~n47911 & n47963;
  assign n47965 = ~n47944 & ~n47963;
  assign n47966 = ~n47964 & ~n47965;
  assign n47967 = ~pi206 & ~n47966;
  assign n47968 = n47952 & n47963;
  assign n47969 = pi206 & ~n47968;
  assign po363 = ~n47967 & ~n47969;
  assign n47971 = n47827 & ~n47911;
  assign n47972 = ~n47827 & ~n47944;
  assign n47973 = ~n47971 & ~n47972;
  assign n47974 = ~pi218 & ~n47973;
  assign n47975 = n47827 & n47952;
  assign n47976 = pi218 & ~n47975;
  assign po375 = ~n47974 & ~n47976;
  assign n47978 = ~n47758 & n47963;
  assign n47979 = ~n47799 & ~n47963;
  assign n47980 = ~n47978 & ~n47979;
  assign n47981 = ~pi220 & ~n47980;
  assign n47982 = n65015 & n47963;
  assign n47983 = pi220 & ~n47982;
  assign po377 = ~n47981 & ~n47983;
  assign n47985 = n33956 & n38182;
  assign n47986 = n64339 & n38225;
  assign n47987 = n30617 & n38181;
  assign n47988 = n9738 & n65019;
  assign n47989 = n62951 & n65019;
  assign n47990 = pi74 & n34066;
  assign n47991 = n47989 & n47990;
  assign n47992 = ~pi54 & n47988;
  assign n47993 = pi74 & n47992;
  assign n47994 = n45942 & n47988;
  assign n47995 = ~pi96 & ~pi1093;
  assign n47996 = n2852 & n47995;
  assign n47997 = n64082 & ~n47996;
  assign n47998 = ~pi96 & n64148;
  assign n47999 = pi479 & ~n47998;
  assign n48000 = n38261 & ~n47999;
  assign n48001 = n47997 & n48000;
  assign n48002 = n62370 & n48001;
  assign n48003 = ~n38975 & n48001;
  assign n48004 = n62370 & n48003;
  assign n48005 = ~n38975 & n48002;
  assign n48006 = ~n65020 & ~n65021;
  assign po232 = n62455 & ~n48006;
  assign n48008 = ~pi39 & pi137;
  assign n48009 = n62952 & n39239;
  assign n48010 = ~pi210 & n40653;
  assign n48011 = pi299 & n48010;
  assign n48012 = n31512 & n40653;
  assign n48013 = ~pi198 & n40668;
  assign n48014 = n65014 & n48013;
  assign n48015 = ~n65022 & ~n48014;
  assign n48016 = ~n48009 & ~n48015;
  assign n48017 = ~pi210 & ~n62455;
  assign n48018 = ~n62455 & n48010;
  assign n48019 = n40653 & n48017;
  assign n48020 = ~n48016 & ~n65023;
  assign n48021 = n33664 & ~n48020;
  assign n48022 = ~n48008 & ~n48021;
  assign n48023 = n34046 & n35420;
  assign n48024 = n34059 & n44475;
  assign n48025 = ~n41010 & ~n65024;
  assign n48026 = pi62 & ~n48025;
  assign n48027 = ~pi100 & n45154;
  assign n48028 = n62380 & ~n34149;
  assign n48029 = ~pi299 & ~n48028;
  assign n48030 = pi299 & ~n44422;
  assign n48031 = ~n48029 & ~n48030;
  assign n48032 = pi100 & n34059;
  assign n48033 = n48031 & n48032;
  assign n48034 = ~pi39 & ~n48033;
  assign n48035 = ~n48027 & n48034;
  assign n48036 = pi39 & ~n34062;
  assign n48037 = ~pi38 & ~n48036;
  assign n48038 = ~n48035 & n48037;
  assign n48039 = ~n41010 & ~n48038;
  assign n48040 = ~pi87 & ~n48039;
  assign n48041 = ~n35420 & ~n41010;
  assign n48042 = pi87 & ~n48041;
  assign n48043 = ~pi75 & ~n48042;
  assign n48044 = ~n48040 & n48043;
  assign n48045 = pi75 & ~n41010;
  assign n48046 = ~pi92 & ~n48045;
  assign n48047 = ~n48044 & n48046;
  assign n48048 = ~n64341 & ~n41010;
  assign n48049 = pi92 & ~n48048;
  assign n48050 = n6792 & ~n48049;
  assign n48051 = ~n48047 & n48050;
  assign n48052 = ~n6792 & ~n41010;
  assign n48053 = ~pi55 & ~n48052;
  assign n48054 = ~n48051 & n48053;
  assign n48055 = ~n64305 & ~n41010;
  assign n48056 = pi55 & ~n48055;
  assign n48057 = ~pi56 & ~n48056;
  assign n48058 = ~n48054 & n48057;
  assign n48059 = n30584 & n35420;
  assign n48060 = n64084 & n34059;
  assign n48061 = pi56 & ~n41010;
  assign n48062 = ~n65025 & n48061;
  assign n48063 = ~pi62 & ~n48062;
  assign n48064 = ~n48058 & n48063;
  assign n48065 = ~n48026 & ~n48064;
  assign n48066 = n3472 & ~n48065;
  assign n48067 = ~n3472 & n41010;
  assign n48068 = ~n48066 & ~n48067;
  assign n48069 = pi40 & ~pi287;
  assign n48070 = n40055 & n48069;
  assign n48071 = ~n40220 & n48070;
  assign n48072 = ~n64705 & ~n48071;
  assign n48073 = n33899 & n39975;
  assign n48074 = ~pi102 & ~n48073;
  assign n48075 = n62355 & n6803;
  assign n48076 = n64196 & n48075;
  assign n48077 = n62355 & n64196;
  assign n48078 = n6803 & n48077;
  assign n48079 = n40591 & n43199;
  assign n48080 = ~n48074 & n65026;
  assign n48081 = n6822 & n48080;
  assign n48082 = ~n48070 & ~n48081;
  assign n48083 = ~n2852 & n48082;
  assign n48084 = n2852 & ~n48081;
  assign n48085 = pi1093 & ~n48084;
  assign n48086 = ~n2852 & ~n48082;
  assign n48087 = n2852 & n48081;
  assign n48088 = ~n48086 & ~n48087;
  assign n48089 = pi1093 & ~n48088;
  assign n48090 = ~n48083 & n48085;
  assign n48091 = ~n2584 & n48082;
  assign n48092 = n2584 & ~n48081;
  assign n48093 = ~pi1093 & ~n48092;
  assign n48094 = ~n2584 & ~n48082;
  assign n48095 = n2584 & n48081;
  assign n48096 = ~n48091 & ~n48092;
  assign n48097 = ~n48094 & ~n48095;
  assign n48098 = ~pi1093 & n65028;
  assign n48099 = ~n48091 & n48093;
  assign n48100 = ~n65027 & ~n65029;
  assign n48101 = ~pi1091 & ~n48100;
  assign n48102 = ~n3008 & n48082;
  assign n48103 = ~n3007 & n48092;
  assign n48104 = pi1091 & ~n48103;
  assign n48105 = ~n48102 & n48104;
  assign n48106 = n64705 & ~n48105;
  assign n48107 = ~n3007 & n65028;
  assign n48108 = n3007 & ~n48082;
  assign n48109 = pi1091 & ~n48108;
  assign n48110 = ~n48107 & n48109;
  assign n48111 = ~pi1091 & ~n65027;
  assign n48112 = ~pi1091 & ~n65029;
  assign n48113 = ~n65027 & n48112;
  assign n48114 = ~n65029 & n48111;
  assign n48115 = ~n48110 & ~n65030;
  assign n48116 = n64705 & ~n48115;
  assign n48117 = ~n48101 & n48106;
  assign po624 = ~n48072 & ~n65031;
  assign n48119 = n39880 & n64701;
  assign n48120 = n2852 & n48119;
  assign n48121 = ~pi1093 & ~n48120;
  assign n48122 = pi1093 & ~n43205;
  assign n48123 = ~n6899 & n64082;
  assign n48124 = ~n48122 & n48123;
  assign n48125 = ~n48121 & n48124;
  assign n48126 = n3318 & ~n48125;
  assign n48127 = ~pi1093 & n2726;
  assign n48128 = ~pi1093 & n64339;
  assign n48129 = n35394 & n48127;
  assign n48130 = ~pi1093 & n2728;
  assign n48131 = n64082 & n48130;
  assign n48132 = n62952 & n65032;
  assign n48133 = n39897 & n65033;
  assign n48134 = n38941 & n48133;
  assign n48135 = n38944 & n48133;
  assign n48136 = n6873 & n48134;
  assign n48137 = ~n3318 & ~n65034;
  assign n48138 = n62455 & ~n48137;
  assign po246 = ~n48126 & n48138;
  assign n48140 = pi1092 & ~n2924;
  assign n48141 = ~n62455 & n48140;
  assign n48142 = ~pi330 & n48141;
  assign n48143 = n62455 & n48140;
  assign n48144 = ~pi340 & n64994;
  assign n48145 = ~pi330 & ~n64994;
  assign n48146 = ~n48144 & ~n48145;
  assign n48147 = pi330 & ~n64994;
  assign n48148 = pi340 & n64994;
  assign n48149 = n48143 & ~n48148;
  assign n48150 = ~n48147 & n48149;
  assign n48151 = n48143 & ~n48146;
  assign n48152 = ~n48142 & ~n65035;
  assign n48153 = ~pi331 & n48141;
  assign n48154 = ~pi341 & n64994;
  assign n48155 = ~pi331 & ~n64994;
  assign n48156 = ~n48154 & ~n48155;
  assign n48157 = pi331 & ~n64994;
  assign n48158 = pi341 & n64994;
  assign n48159 = n48143 & ~n48158;
  assign n48160 = ~n48157 & n48159;
  assign n48161 = n48143 & ~n48156;
  assign n48162 = ~n48153 & ~n65036;
  assign n48163 = pi340 & n48141;
  assign n48164 = ~pi331 & n64994;
  assign n48165 = ~pi340 & ~n64994;
  assign n48166 = n48143 & ~n48165;
  assign n48167 = n48143 & ~n48164;
  assign n48168 = ~n48165 & n48167;
  assign n48169 = ~n48164 & n48166;
  assign po497 = ~n48163 & ~n65037;
  assign n48171 = ~pi330 & po637;
  assign n48172 = ~pi341 & ~po637;
  assign n48173 = ~n48171 & ~n48172;
  assign po498 = n48140 & ~n48173;
  assign n48175 = n38226 & n39025;
  assign n48176 = n38262 & n41393;
  assign n48177 = pi96 & n2750;
  assign n48178 = pi96 & n2585;
  assign n48179 = n2750 & n48178;
  assign n48180 = n2585 & n48177;
  assign n48181 = ~n38262 & n65038;
  assign n48182 = n41048 & n48181;
  assign n48183 = ~n48176 & ~n48182;
  assign n48184 = ~pi95 & ~n48183;
  assign n48185 = ~n48175 & ~n48184;
  assign po254 = n64705 & ~n48185;
  assign n48187 = n39702 & n48031;
  assign n48188 = ~n46299 & ~n48187;
  assign n48189 = ~pi38 & ~n48188;
  assign n48190 = ~pi87 & ~n48189;
  assign n48191 = n34034 & ~n48190;
  assign n48192 = ~pi92 & ~n48191;
  assign n48193 = ~pi74 & n37887;
  assign n48194 = ~n48192 & n48193;
  assign n48195 = ~pi55 & ~n48194;
  assign n48196 = ~n30903 & ~n48195;
  assign n48197 = ~pi56 & ~n48196;
  assign n48198 = ~n34043 & ~n48197;
  assign n48199 = ~pi62 & ~n48198;
  assign n48200 = ~pi57 & n34049;
  assign po275 = ~n48199 & n48200;
  assign n48202 = ~pi58 & n2858;
  assign n48203 = n2663 & n39887;
  assign n48204 = ~n48202 & ~n48203;
  assign n48205 = n64196 & ~n48204;
  assign n48206 = n3007 & ~n48205;
  assign n48207 = ~n2582 & n48205;
  assign n48208 = n6921 & n48119;
  assign n48209 = pi829 & ~n48208;
  assign n48210 = ~n48207 & n48209;
  assign n48211 = ~n2824 & n48210;
  assign n48212 = ~n48206 & ~n48211;
  assign n48213 = pi1091 & ~n48212;
  assign n48214 = ~n2852 & n48205;
  assign n48215 = ~pi829 & ~n48214;
  assign n48216 = ~n48210 & ~n48215;
  assign n48217 = ~pi1093 & ~n48216;
  assign n48218 = ~n39846 & ~n48202;
  assign n48219 = n43203 & ~n48218;
  assign n48220 = ~n3032 & ~n30822;
  assign n48221 = ~n48219 & ~n48220;
  assign n48222 = ~n48214 & n48221;
  assign n48223 = n64705 & ~n48222;
  assign n48224 = ~n48217 & n48223;
  assign po205 = ~n48213 & n48224;
  assign n48226 = pi1093 & n64528;
  assign n48227 = ~pi96 & ~n48226;
  assign n48228 = n2806 & ~n33973;
  assign n48229 = pi96 & ~pi1093;
  assign n48230 = n2927 & ~n38975;
  assign n48231 = ~n48229 & ~n48230;
  assign n48232 = n2806 & ~n48231;
  assign n48233 = ~n48227 & n48228;
  assign n48234 = n62392 & n65039;
  assign n48235 = ~pi75 & ~n48234;
  assign n48236 = pi75 & ~n47989;
  assign n48237 = n40103 & ~n48236;
  assign po233 = ~n48235 & n48237;
  assign n48239 = ~pi340 & po637;
  assign n48240 = n62455 & n48144;
  assign n48241 = pi315 & ~n65040;
  assign n48242 = pi1080 & n65040;
  assign n48243 = ~n48241 & ~n48242;
  assign n48244 = pi316 & ~n65040;
  assign n48245 = pi1047 & n65040;
  assign n48246 = ~n48244 & ~n48245;
  assign n48247 = pi317 & ~n48171;
  assign n48248 = pi1078 & n48171;
  assign n48249 = ~n48247 & ~n48248;
  assign n48250 = ~pi341 & po637;
  assign n48251 = n62455 & n48154;
  assign n48252 = pi318 & ~n65041;
  assign n48253 = pi1074 & n65041;
  assign n48254 = ~n48252 & ~n48253;
  assign n48255 = pi319 & ~n65041;
  assign n48256 = pi1072 & n65041;
  assign n48257 = ~n48255 & ~n48256;
  assign n48258 = pi320 & ~n65040;
  assign n48259 = pi1048 & n65040;
  assign n48260 = ~n48258 & ~n48259;
  assign n48261 = pi321 & ~n65040;
  assign n48262 = pi1058 & n65040;
  assign n48263 = ~n48261 & ~n48262;
  assign n48264 = pi322 & ~n65040;
  assign n48265 = pi1051 & n65040;
  assign n48266 = ~n48264 & ~n48265;
  assign n48267 = pi323 & ~n65040;
  assign n48268 = pi1065 & n65040;
  assign n48269 = ~n48267 & ~n48268;
  assign n48270 = pi324 & ~n65041;
  assign n48271 = pi1086 & n65041;
  assign n48272 = ~n48270 & ~n48271;
  assign n48273 = pi325 & ~n65041;
  assign n48274 = pi1063 & n65041;
  assign n48275 = ~n48273 & ~n48274;
  assign n48276 = pi326 & ~n65041;
  assign n48277 = pi1057 & n65041;
  assign n48278 = ~n48276 & ~n48277;
  assign n48279 = pi327 & ~n65040;
  assign n48280 = pi1040 & n65040;
  assign n48281 = ~n48279 & ~n48280;
  assign n48282 = pi328 & ~n65041;
  assign n48283 = pi1058 & n65041;
  assign n48284 = ~n48282 & ~n48283;
  assign n48285 = pi329 & ~n65041;
  assign n48286 = pi1043 & n65041;
  assign n48287 = ~n48285 & ~n48286;
  assign n48288 = pi333 & ~n65041;
  assign n48289 = pi1040 & n65041;
  assign n48290 = ~n48288 & ~n48289;
  assign n48291 = pi334 & ~n65041;
  assign n48292 = pi1065 & n65041;
  assign n48293 = ~n48291 & ~n48292;
  assign n48294 = pi335 & ~n65041;
  assign n48295 = pi1069 & n65041;
  assign n48296 = ~n48294 & ~n48295;
  assign n48297 = pi338 & ~n48171;
  assign n48298 = pi1072 & n48171;
  assign n48299 = ~n48297 & ~n48298;
  assign n48300 = pi339 & ~n48171;
  assign n48301 = pi1086 & n48171;
  assign n48302 = ~n48300 & ~n48301;
  assign n48303 = pi344 & ~n65040;
  assign n48304 = pi1069 & n65040;
  assign n48305 = ~n48303 & ~n48304;
  assign n48306 = pi349 & ~n65040;
  assign n48307 = pi1043 & n65040;
  assign n48308 = ~n48306 & ~n48307;
  assign n48309 = pi352 & ~n65040;
  assign n48310 = pi1078 & n65040;
  assign n48311 = ~n48309 & ~n48310;
  assign n48312 = pi353 & ~n65040;
  assign n48313 = pi1063 & n65040;
  assign n48314 = ~n48312 & ~n48313;
  assign n48315 = pi365 & ~n48171;
  assign n48316 = pi1065 & n48171;
  assign n48317 = ~n48315 & ~n48316;
  assign n48318 = pi366 & ~n48171;
  assign n48319 = pi1069 & n48171;
  assign n48320 = ~n48318 & ~n48319;
  assign n48321 = pi369 & ~n48171;
  assign n48322 = pi1080 & n48171;
  assign n48323 = ~n48321 & ~n48322;
  assign n48324 = pi371 & ~n48171;
  assign n48325 = pi1051 & n48171;
  assign n48326 = ~n48324 & ~n48325;
  assign n48327 = pi372 & ~n48171;
  assign n48328 = pi1048 & n48171;
  assign n48329 = ~n48327 & ~n48328;
  assign n48330 = pi375 & ~n48171;
  assign n48331 = pi1047 & n48171;
  assign n48332 = ~n48330 & ~n48331;
  assign n48333 = pi377 & ~n48171;
  assign n48334 = pi1074 & n48171;
  assign n48335 = ~n48333 & ~n48334;
  assign n48336 = pi378 & ~n48171;
  assign n48337 = pi1063 & n48171;
  assign n48338 = ~n48336 & ~n48337;
  assign n48339 = pi394 & ~n65041;
  assign n48340 = pi1080 & n65041;
  assign n48341 = ~n48339 & ~n48340;
  assign n48342 = pi396 & ~n65041;
  assign n48343 = pi1051 & n65041;
  assign n48344 = ~n48342 & ~n48343;
  assign n48345 = pi397 & ~n65041;
  assign n48346 = pi1048 & n65041;
  assign n48347 = ~n48345 & ~n48346;
  assign n48348 = pi399 & ~n65041;
  assign n48349 = pi1047 & n65041;
  assign n48350 = ~n48348 & ~n48349;
  assign n48351 = pi402 & ~n65041;
  assign n48352 = pi1078 & n65041;
  assign n48353 = ~n48351 & ~n48352;
  assign n48354 = n62455 & n48164;
  assign n48355 = pi416 & ~n48354;
  assign n48356 = pi1069 & n48354;
  assign n48357 = ~n48355 & ~n48356;
  assign n48358 = pi419 & ~n48354;
  assign n48359 = pi1080 & n48354;
  assign n48360 = ~n48358 & ~n48359;
  assign n48361 = pi421 & ~n48354;
  assign n48362 = pi1051 & n48354;
  assign n48363 = ~n48361 & ~n48362;
  assign n48364 = pi422 & ~n48354;
  assign n48365 = pi1048 & n48354;
  assign n48366 = ~n48364 & ~n48365;
  assign n48367 = pi424 & ~n48354;
  assign n48368 = pi1047 & n48354;
  assign n48369 = ~n48367 & ~n48368;
  assign n48370 = pi427 & ~n48354;
  assign n48371 = pi1078 & n48354;
  assign n48372 = ~n48370 & ~n48371;
  assign n48373 = pi439 & ~n48171;
  assign n48374 = pi1057 & n48171;
  assign n48375 = ~n48373 & ~n48374;
  assign n48376 = pi440 & ~n48171;
  assign n48377 = pi1043 & n48171;
  assign n48378 = ~n48376 & ~n48377;
  assign n48379 = pi442 & ~n48171;
  assign n48380 = pi1058 & n48171;
  assign n48381 = ~n48379 & ~n48380;
  assign n48382 = pi444 & ~n48354;
  assign n48383 = pi1072 & n48354;
  assign n48384 = ~n48382 & ~n48383;
  assign n48385 = pi446 & ~n48354;
  assign n48386 = pi1086 & n48354;
  assign n48387 = ~n48385 & ~n48386;
  assign n48388 = pi447 & ~n48171;
  assign n48389 = pi1040 & n48171;
  assign n48390 = ~n48388 & ~n48389;
  assign n48391 = pi448 & ~n48354;
  assign n48392 = pi1074 & n48354;
  assign n48393 = ~n48391 & ~n48392;
  assign n48394 = pi449 & ~n48354;
  assign n48395 = pi1057 & n48354;
  assign n48396 = ~n48394 & ~n48395;
  assign n48397 = pi451 & ~n48354;
  assign n48398 = pi1063 & n48354;
  assign n48399 = ~n48397 & ~n48398;
  assign n48400 = pi453 & ~n48354;
  assign n48401 = pi1040 & n48354;
  assign n48402 = ~n48400 & ~n48401;
  assign n48403 = pi454 & ~n48354;
  assign n48404 = pi1043 & n48354;
  assign n48405 = ~n48403 & ~n48404;
  assign n48406 = pi458 & ~n65040;
  assign n48407 = pi1072 & n65040;
  assign n48408 = ~n48406 & ~n48407;
  assign n48409 = pi459 & ~n48354;
  assign n48410 = pi1058 & n48354;
  assign n48411 = ~n48409 & ~n48410;
  assign n48412 = pi460 & ~n65040;
  assign n48413 = pi1086 & n65040;
  assign n48414 = ~n48412 & ~n48413;
  assign n48415 = pi461 & ~n65040;
  assign n48416 = pi1057 & n65040;
  assign n48417 = ~n48415 & ~n48416;
  assign n48418 = pi462 & ~n65040;
  assign n48419 = pi1074 & n65040;
  assign n48420 = ~n48418 & ~n48419;
  assign n48421 = pi464 & ~n48354;
  assign n48422 = pi1065 & n48354;
  assign n48423 = ~n48421 & ~n48422;
  assign n48424 = ~pi97 & n62359;
  assign n48425 = ~pi108 & ~n48424;
  assign n48426 = n2664 & n2696;
  assign n48427 = ~n38903 & n48426;
  assign n48428 = ~n48425 & n48427;
  assign n48429 = n64582 & n48428;
  assign n48430 = n62362 & n38903;
  assign n48431 = ~pi51 & ~n48430;
  assign n48432 = n2664 & ~n48425;
  assign n48433 = n64582 & n48432;
  assign n48434 = ~pi314 & ~n48433;
  assign n48435 = pi314 & ~n2708;
  assign n48436 = n2696 & ~n38902;
  assign n48437 = ~n48435 & n48436;
  assign n48438 = ~n48434 & n48437;
  assign n48439 = n2696 & n38902;
  assign n48440 = n48433 & n48439;
  assign n48441 = ~pi51 & ~n48440;
  assign n48442 = ~n48438 & n48441;
  assign n48443 = ~n48429 & n48431;
  assign n48444 = n62367 & n62373;
  assign n48445 = ~n65042 & n48444;
  assign n48446 = ~pi87 & ~n48445;
  assign n48447 = n34034 & n40103;
  assign po266 = ~n48446 & n48447;
  assign n48449 = pi39 & ~pi979;
  assign n48450 = ~n2934 & n48449;
  assign n48451 = n2935 & n48450;
  assign n48452 = n2933 & n48451;
  assign n48453 = n64325 & n48452;
  assign n48454 = n10335 & n63888;
  assign n48455 = n62384 & n48454;
  assign n48456 = pi468 & ~n48455;
  assign n48457 = ~n48453 & ~n48456;
  assign n48458 = n62355 & n31435;
  assign n48459 = pi24 & n64196;
  assign n48460 = ~pi39 & n48459;
  assign n48461 = ~pi39 & n48458;
  assign n48462 = n48459 & n48461;
  assign n48463 = n48458 & n48460;
  assign n48464 = n30638 & n65043;
  assign n48465 = ~n48452 & ~n48464;
  assign po218 = n64325 & ~n48465;
  assign n48467 = po740 & n64866;
  assign po194 = ~n48218 & n48467;
  assign n48469 = n2602 & n30677;
  assign n48470 = n39874 & n48469;
  assign n48471 = ~pi64 & n6811;
  assign n48472 = n48470 & n48471;
  assign n48473 = ~pi81 & ~n48472;
  assign n48474 = ~pi199 & pi200;
  assign n48475 = ~pi299 & n48474;
  assign n48476 = pi211 & ~pi219;
  assign n48477 = pi299 & n48476;
  assign n48478 = ~n48475 & ~n48477;
  assign n48479 = pi314 & ~n48478;
  assign n48480 = n64196 & n48479;
  assign n48481 = ~n48473 & n48480;
  assign n48482 = n34955 & n48481;
  assign n48483 = pi314 & n2613;
  assign n48484 = n64701 & n48483;
  assign n48485 = n64663 & n48478;
  assign n48486 = n48484 & n48485;
  assign n48487 = n48470 & n48486;
  assign n48488 = ~n48482 & ~n48487;
  assign po229 = n64705 & ~n48488;
  assign n48490 = pi81 & ~pi102;
  assign n48491 = n48484 & n48490;
  assign n48492 = n2632 & n48491;
  assign n48493 = n64082 & n48492;
  assign n48494 = pi211 & pi299;
  assign n48495 = pi219 & pi299;
  assign n48496 = ~n48494 & ~n48495;
  assign n48497 = ~pi299 & n39538;
  assign n48498 = ~pi211 & pi299;
  assign n48499 = ~pi219 & n48498;
  assign n48500 = ~n48497 & ~n48499;
  assign n48501 = ~n39539 & n48496;
  assign n48502 = n62455 & ~n65044;
  assign po242 = n48493 & n48502;
  assign n48504 = ~n39166 & ~n43691;
  assign n48505 = ~pi314 & n43691;
  assign n48506 = po740 & ~n48505;
  assign n48507 = n64866 & ~n48506;
  assign n48508 = ~n48504 & n48507;
  assign n48509 = pi53 & n2682;
  assign n48510 = n62361 & n48509;
  assign n48511 = n64092 & n48510;
  assign n48512 = n48459 & n48511;
  assign n48513 = ~pi39 & ~n48512;
  assign n48514 = ~pi287 & ~pi979;
  assign n48515 = n2934 & n48514;
  assign n48516 = pi39 & ~n48515;
  assign n48517 = n64325 & ~n48516;
  assign n48518 = ~n40219 & n48517;
  assign n48519 = ~n48513 & n48517;
  assign n48520 = ~n40219 & n48519;
  assign n48521 = ~n48513 & n48518;
  assign n48522 = ~n41056 & ~n41325;
  assign n48523 = ~pi70 & ~n48522;
  assign n48524 = ~pi51 & ~n48523;
  assign n48525 = n2733 & ~n48524;
  assign n48526 = n33868 & ~n48525;
  assign n48527 = n33860 & ~n48526;
  assign n48528 = n33859 & ~n48527;
  assign n48529 = ~n33959 & ~n48528;
  assign n48530 = ~pi95 & ~n48529;
  assign n48531 = n41047 & ~n48530;
  assign n48532 = ~pi39 & ~n48531;
  assign n48533 = ~pi38 & ~n40219;
  assign n48534 = ~n48532 & n48533;
  assign n48535 = ~pi100 & n48534;
  assign n48536 = n40229 & ~n48535;
  assign n48537 = ~n34033 & ~n48536;
  assign n48538 = ~pi75 & ~n48537;
  assign n48539 = ~n30600 & ~n48538;
  assign n48540 = ~pi92 & ~n48539;
  assign n48541 = n37887 & ~n48540;
  assign n48542 = ~pi74 & ~n48541;
  assign n48543 = n33857 & ~n48542;
  assign n48544 = ~pi56 & ~n48543;
  assign n48545 = ~n34043 & ~n48544;
  assign n48546 = ~pi62 & ~n48545;
  assign po393 = n48200 & ~n48546;
  assign n48548 = ~n62455 & n48476;
  assign n48549 = pi71 & n48548;
  assign n48550 = pi71 & ~n48478;
  assign n48551 = pi84 & n31456;
  assign n48552 = n41810 & n48551;
  assign n48553 = n2588 & n48552;
  assign n48554 = n62352 & n43682;
  assign n48555 = n2665 & n48554;
  assign n48556 = n62356 & n43682;
  assign n48557 = n48478 & n65046;
  assign n48558 = n64337 & ~n48478;
  assign n48559 = n38940 & n48558;
  assign n48560 = ~n48557 & ~n48559;
  assign n48561 = n64082 & n64196;
  assign n48562 = ~n48560 & n48561;
  assign n48563 = n48553 & n48562;
  assign n48564 = ~n48550 & ~n48563;
  assign n48565 = n62455 & ~n48564;
  assign n48566 = ~n48549 & ~n48565;
  assign n48567 = ~pi199 & ~pi299;
  assign n48568 = n48493 & ~n48567;
  assign n48569 = pi219 & ~n48568;
  assign n48570 = pi199 & ~pi299;
  assign n48571 = n2805 & n48570;
  assign n48572 = n43880 & n48571;
  assign n48573 = n48492 & n48572;
  assign n48574 = ~pi219 & ~n48573;
  assign n48575 = n62455 & ~n48574;
  assign po224 = ~n48569 & n48575;
  assign n48577 = pi54 & n62380;
  assign n48578 = ~pi49 & ~pi76;
  assign n48579 = n6809 & n48578;
  assign n48580 = ~pi60 & ~pi85;
  assign n48581 = pi106 & n48580;
  assign n48582 = n2598 & n38884;
  assign n48583 = n48581 & n48582;
  assign n48584 = n48579 & n48583;
  assign n48585 = n6808 & n39981;
  assign n48586 = n48584 & n48585;
  assign n48587 = n43524 & n48586;
  assign n48588 = ~pi53 & ~n48587;
  assign n48589 = n32085 & ~n48588;
  assign n48590 = ~pi54 & n40591;
  assign n48591 = n48589 & n48590;
  assign n48592 = ~n48577 & ~n48591;
  assign n48593 = n9738 & n64498;
  assign n48594 = ~n48592 & n48593;
  assign n48595 = ~pi39 & ~n48594;
  assign po456 = ~n48516 & ~n48595;
  assign n48597 = pi38 & ~n65019;
  assign n48598 = pi332 & n38242;
  assign n48599 = ~pi64 & ~n48598;
  assign n48600 = ~pi39 & ~pi841;
  assign n48601 = n2614 & n48600;
  assign n48602 = ~pi39 & ~pi81;
  assign n48603 = ~pi841 & n48602;
  assign n48604 = n2626 & n48603;
  assign n48605 = n2613 & n48601;
  assign n48606 = n64701 & n65047;
  assign n48607 = ~n48599 & n65047;
  assign n48608 = n64701 & n48607;
  assign n48609 = ~n48599 & n48606;
  assign n48610 = ~pi81 & ~n33875;
  assign n48611 = n2626 & n48600;
  assign n48612 = n64701 & n48611;
  assign n48613 = ~n48599 & n48611;
  assign n48614 = n64701 & n48613;
  assign n48615 = ~n48599 & n48612;
  assign n48616 = n48610 & n65049;
  assign n48617 = ~n33875 & n65048;
  assign n48618 = ~pi38 & ~n65050;
  assign n48619 = n63888 & ~n48618;
  assign po196 = ~n48597 & n48619;
  assign n48621 = pi979 & n39838;
  assign po203 = n2933 & n48621;
  assign n48623 = n38228 & n43526;
  assign n48624 = n38228 & n48579;
  assign n48625 = n43526 & n48624;
  assign n48626 = n48579 & n48623;
  assign n48627 = pi61 & ~pi82;
  assign n48628 = ~pi83 & ~pi89;
  assign n48629 = n48627 & n48628;
  assign n48630 = n2687 & n39978;
  assign n48631 = n48629 & n48630;
  assign n48632 = n39983 & n48631;
  assign n48633 = n38890 & n48632;
  assign n48634 = n65051 & n48633;
  assign n48635 = n62356 & n48634;
  assign n48636 = ~pi841 & n48635;
  assign n48637 = n2665 & n30630;
  assign n48638 = pi24 & n48637;
  assign n48639 = ~n48636 & ~n48638;
  assign po204 = n64866 & ~n48639;
  assign n48641 = pi74 & ~n62384;
  assign n48642 = pi841 & n2694;
  assign n48643 = pi841 & n2771;
  assign n48644 = n2694 & n48643;
  assign n48645 = n2728 & n48644;
  assign n48646 = ~pi72 & pi841;
  assign n48647 = ~pi70 & pi841;
  assign n48648 = n2729 & n48647;
  assign n48649 = n2771 & n48646;
  assign n48650 = n2694 & n65053;
  assign n48651 = n2751 & n48650;
  assign n48652 = n32374 & n65053;
  assign n48653 = n62378 & n48642;
  assign n48654 = n43537 & n65052;
  assign n48655 = ~pi74 & ~n48654;
  assign n48656 = n40691 & ~n48655;
  assign po207 = ~n48641 & n48656;
  assign n48658 = pi54 & ~n47988;
  assign n48659 = n48458 & n48587;
  assign n48660 = n6829 & n64081;
  assign n48661 = n43538 & n48660;
  assign n48662 = n48659 & n48661;
  assign n48663 = ~pi54 & ~n48662;
  assign n48664 = n64498 & ~n48663;
  assign n48665 = pi54 & n47988;
  assign n48666 = ~pi54 & n6829;
  assign n48667 = n64081 & n48666;
  assign n48668 = n43538 & n48667;
  assign n48669 = n48659 & n48668;
  assign n48670 = ~n48665 & ~n48669;
  assign n48671 = n64498 & ~n48670;
  assign n48672 = ~n48658 & n48664;
  assign n48673 = pi55 & n40045;
  assign n48674 = ~n43668 & ~n48673;
  assign n48675 = n2727 & n64084;
  assign n48676 = n33953 & n48675;
  assign n48677 = pi56 & ~n48676;
  assign n48678 = n3472 & ~n48677;
  assign po214 = ~n48674 & n48678;
  assign n48680 = pi841 & n48635;
  assign n48681 = ~pi24 & n48458;
  assign n48682 = n31435 & n64761;
  assign n48683 = n30638 & n65055;
  assign n48684 = ~n48680 & ~n48683;
  assign po219 = n64866 & ~n48684;
  assign n48686 = pi57 & ~n40046;
  assign n48687 = n43669 & n48676;
  assign n48688 = ~pi57 & ~n48687;
  assign n48689 = ~pi59 & ~n48688;
  assign n48690 = ~pi59 & ~n48686;
  assign n48691 = ~n48688 & n48690;
  assign n48692 = ~n48686 & n48689;
  assign n48693 = pi841 & n2696;
  assign n48694 = n38243 & n48693;
  assign n48695 = ~pi24 & pi70;
  assign n48696 = n62364 & n48695;
  assign n48697 = ~n48694 & ~n48696;
  assign n48698 = n62381 & n64705;
  assign n48699 = pi70 & ~n2818;
  assign n48700 = pi841 & n2695;
  assign n48701 = n38243 & n48700;
  assign n48702 = ~pi70 & ~n48701;
  assign n48703 = n48698 & ~n48702;
  assign n48704 = ~n48699 & n48703;
  assign n48705 = ~n48697 & n48698;
  assign n48706 = ~pi1050 & n32114;
  assign n48707 = ~pi90 & ~n48706;
  assign n48708 = ~pi93 & n35400;
  assign n48709 = n2585 & n48698;
  assign n48710 = n35400 & n64705;
  assign n48711 = ~pi93 & n65058;
  assign n48712 = n64705 & n48708;
  assign n48713 = ~n48707 & n65059;
  assign n48714 = ~n48707 & n65058;
  assign n48715 = n34979 & n48714;
  assign n48716 = ~n30627 & n48713;
  assign po248 = ~n2675 & n65060;
  assign n48718 = pi93 & n35400;
  assign n48719 = n30624 & n48718;
  assign n48720 = ~pi92 & ~n48719;
  assign n48721 = ~pi1050 & n62380;
  assign n48722 = pi92 & ~n48721;
  assign n48723 = n40697 & ~n48722;
  assign n48724 = n40697 & ~n48720;
  assign n48725 = ~n48722 & n48724;
  assign n48726 = ~n48720 & n48723;
  assign n48727 = ~pi92 & n64197;
  assign n48728 = ~n38966 & ~n48727;
  assign n48729 = pi314 & pi1050;
  assign n48730 = n40697 & n48729;
  assign po256 = ~n48728 & n48730;
  assign n48732 = pi24 & n48659;
  assign n48733 = n41823 & n48589;
  assign n48734 = ~n48732 & ~n48733;
  assign n48735 = pi841 & ~n48734;
  assign n48736 = n40148 & n48511;
  assign n48737 = ~n48735 & ~n48736;
  assign po264 = n64866 & ~n48737;
  assign n48739 = pi72 & n39025;
  assign n48740 = n62768 & n48505;
  assign n48741 = ~n48739 & ~n48740;
  assign po269 = n43679 & ~n48741;
  assign n48743 = n38244 & n48637;
  assign n48744 = ~n38243 & ~n48637;
  assign n48745 = n2695 & ~n48744;
  assign n48746 = ~pi70 & ~n48745;
  assign n48747 = pi332 & n32075;
  assign n48748 = ~n48746 & n48747;
  assign n48749 = ~n48743 & ~n48748;
  assign n48750 = ~pi39 & ~n48749;
  assign n48751 = pi39 & n39239;
  assign n48752 = ~pi38 & ~n48751;
  assign n48753 = ~n48750 & n48752;
  assign po489 = n38727 & ~n48753;
  assign n48755 = ~pi93 & pi102;
  assign n48756 = pi102 & n2715;
  assign n48757 = n2586 & n48755;
  assign n48758 = n2613 & n65062;
  assign n48759 = n62382 & n48758;
  assign n48760 = pi102 & n2613;
  assign n48761 = n62382 & n48760;
  assign n48762 = n2716 & n48761;
  assign n48763 = n62354 & n48759;
  assign n48764 = n2633 & n65063;
  assign n48765 = ~pi40 & ~n48764;
  assign n48766 = n6802 & ~n48765;
  assign n48767 = ~pi1082 & ~n48766;
  assign n48768 = n2751 & n48764;
  assign n48769 = pi1082 & ~n48768;
  assign n48770 = n64705 & ~n48769;
  assign po198 = ~n48767 & n48770;
  assign n48772 = pi841 & n64705;
  assign n48773 = n38897 & n48772;
  assign n48774 = ~pi51 & n65053;
  assign n48775 = n38897 & n48774;
  assign n48776 = n64705 & n48775;
  assign n48777 = n40604 & n48776;
  assign n48778 = n64701 & n48773;
  assign n48779 = n6792 & n47988;
  assign n48780 = ~pi74 & n47992;
  assign n48781 = n62952 & n65019;
  assign n48782 = pi55 & ~n65065;
  assign n48783 = n2626 & n64082;
  assign n48784 = n64701 & n48783;
  assign n48785 = n2626 & n64701;
  assign n48786 = n6819 & n64082;
  assign n48787 = n48785 & n48786;
  assign n48788 = n6819 & n48784;
  assign n48789 = ~pi55 & ~n65066;
  assign n48790 = n3473 & ~n48789;
  assign po213 = ~n48782 & n48790;
  assign po216 = n2675 & n65059;
  assign n48793 = n2663 & n64866;
  assign n48794 = n2655 & n48793;
  assign n48795 = ~pi107 & pi841;
  assign n48796 = pi64 & ~n48795;
  assign n48797 = ~pi64 & ~pi107;
  assign n48798 = ~pi63 & ~pi81;
  assign n48799 = ~n48797 & n48798;
  assign n48800 = ~n48796 & n48799;
  assign n48801 = n2626 & n48800;
  assign n48802 = n48794 & n48801;
  assign n48803 = ~pi63 & pi107;
  assign n48804 = n2625 & n48803;
  assign n48805 = ~pi64 & ~n48804;
  assign n48806 = n2626 & ~n48805;
  assign n48807 = n48610 & n48806;
  assign n48808 = pi841 & ~n48807;
  assign n48809 = n62348 & n48803;
  assign n48810 = ~pi841 & ~n48809;
  assign n48811 = n48794 & ~n48810;
  assign n48812 = ~n48808 & n48811;
  assign n48813 = n2625 & n48802;
  assign n48814 = pi83 & ~pi103;
  assign n48815 = n43682 & n48814;
  assign n48816 = n64705 & n48814;
  assign n48817 = n43682 & n48816;
  assign n48818 = n64705 & n48815;
  assign n48819 = n48484 & n65068;
  assign n48820 = n62345 & n65068;
  assign n48821 = n48484 & n48820;
  assign n48822 = n62345 & n48819;
  assign n48823 = pi69 & n6807;
  assign n48824 = n35357 & n48823;
  assign n48825 = ~pi71 & ~n48824;
  assign n48826 = ~pi81 & ~pi314;
  assign n48827 = n2626 & n48826;
  assign n48828 = n30696 & n48827;
  assign n48829 = ~n48825 & n48828;
  assign n48830 = pi71 & pi314;
  assign n48831 = n2687 & n48830;
  assign n48832 = n64337 & n48831;
  assign n48833 = n2610 & n48832;
  assign n48834 = ~n48829 & ~n48833;
  assign po227 = n48794 & ~n48834;
  assign n48836 = ~pi314 & ~n41857;
  assign n48837 = pi314 & ~n41855;
  assign n48838 = n64866 & ~n48837;
  assign po235 = ~n48836 & n48838;
  assign n48840 = n62455 & n48784;
  assign n48841 = n64705 & n48785;
  assign n48842 = pi81 & ~pi314;
  assign n48843 = n2632 & n48842;
  assign n48844 = pi68 & ~pi81;
  assign n48845 = n2599 & n48844;
  assign n48846 = n39874 & n48845;
  assign n48847 = n48471 & n48846;
  assign n48848 = n30651 & n48847;
  assign n48849 = ~n48843 & ~n48848;
  assign po239 = n65070 & ~n48849;
  assign n48851 = pi69 & pi314;
  assign n48852 = n2607 & n48851;
  assign n48853 = pi66 & ~pi73;
  assign n48854 = n2606 & n48853;
  assign n48855 = n2600 & n48854;
  assign n48856 = n2603 & n48854;
  assign n48857 = n2596 & n48855;
  assign n48858 = ~n48852 & ~n65071;
  assign n48859 = n43683 & n48794;
  assign po240 = ~n48858 & n48859;
  assign n48861 = ~pi83 & ~n48552;
  assign n48862 = n30648 & n65046;
  assign n48863 = n65046 & ~n48861;
  assign n48864 = n30648 & n48863;
  assign n48865 = ~n48861 & n48862;
  assign n48866 = ~pi314 & ~n65072;
  assign n48867 = n48553 & n65046;
  assign n48868 = pi314 & ~n48867;
  assign n48869 = n64866 & ~n48868;
  assign po241 = ~n48866 & n48869;
  assign n48871 = n30688 & n43684;
  assign n48872 = ~pi314 & n43685;
  assign n48873 = n48469 & n48872;
  assign n48874 = ~n48871 & ~n48873;
  assign po243 = n48794 & ~n48874;
  assign n48876 = n64095 & n48554;
  assign n48877 = pi314 & n64866;
  assign n48878 = n2665 & n48877;
  assign po245 = n48876 & n48878;
  assign n48880 = ~pi109 & ~n48876;
  assign n48881 = n30749 & ~n48880;
  assign n48882 = ~pi314 & ~n48881;
  assign n48883 = pi109 & n2866;
  assign n48884 = n2671 & n48883;
  assign n48885 = pi314 & ~n48884;
  assign n48886 = n48793 & ~n48885;
  assign po261 = ~n48882 & n48886;
  assign po267 = n41937 & n48877;
  assign n48889 = n62373 & n64700;
  assign n48890 = ~n30856 & ~n48889;
  assign n48891 = ~pi75 & ~n48890;
  assign n48892 = n30884 & n40025;
  assign n48893 = ~n48891 & ~n48892;
  assign n48894 = ~pi87 & ~pi250;
  assign n48895 = n40103 & n48894;
  assign po407 = ~n48893 & n48895;
  assign n48897 = n43685 & n48794;
  assign n48898 = n64094 & n43685;
  assign n48899 = n48794 & n48898;
  assign n48900 = n64094 & n48897;
  assign po260 = n48073 & n65070;
  assign n48902 = n62455 & n34255;
  assign n48903 = ~n47808 & ~n48902;
  assign n48904 = ~pi202 & n48903;
  assign n48905 = ~n34078 & n65014;
  assign n48906 = ~n47950 & ~n48905;
  assign n48907 = ~pi205 & n48906;
  assign n48908 = ~pi233 & ~n48907;
  assign n48909 = ~pi233 & ~n48904;
  assign n48910 = ~n48907 & n48909;
  assign n48911 = ~n48904 & n48908;
  assign n48912 = ~pi201 & n48903;
  assign n48913 = ~pi204 & n48906;
  assign n48914 = pi233 & ~n48913;
  assign n48915 = pi233 & ~n48912;
  assign n48916 = ~n48913 & n48915;
  assign n48917 = ~n48912 & n48914;
  assign n48918 = ~n65074 & ~n65075;
  assign n48919 = pi237 & ~n48918;
  assign n48920 = ~pi203 & n48903;
  assign n48921 = ~pi218 & n48906;
  assign n48922 = ~pi233 & ~n48921;
  assign n48923 = ~pi233 & ~n48920;
  assign n48924 = ~n48921 & n48923;
  assign n48925 = ~n48920 & n48922;
  assign n48926 = ~pi220 & n48903;
  assign n48927 = ~pi206 & n48906;
  assign n48928 = pi233 & ~n48927;
  assign n48929 = pi233 & ~n48926;
  assign n48930 = ~n48927 & n48929;
  assign n48931 = ~n48926 & n48928;
  assign n48932 = ~n65076 & ~n65077;
  assign n48933 = ~pi237 & ~n48932;
  assign po746 = ~n48919 & ~n48933;
  assign n48935 = ~pi211 & ~n62455;
  assign n48936 = ~pi219 & n48935;
  assign n48937 = ~n62455 & n39421;
  assign n48938 = ~n48502 & ~n65078;
  assign po635 = pi71 & ~n48938;
  assign n48940 = ~pi270 & ~pi277;
  assign n48941 = ~pi282 & n48940;
  assign n48942 = pi266 & ~pi269;
  assign n48943 = pi278 & pi279;
  assign n48944 = ~pi280 & n48943;
  assign n48945 = n48942 & n48944;
  assign n48946 = ~pi281 & n48945;
  assign n48947 = n48941 & n48946;
  assign n48948 = pi264 & ~n48947;
  assign n48949 = ~pi264 & n48947;
  assign po953 = ~n48948 & ~n48949;
  assign n48951 = n5530 & n31067;
  assign n48952 = ~n30913 & ~n48951;
  assign n48953 = ~pi982 & ~n6899;
  assign n48954 = n3032 & n5530;
  assign n48955 = ~n48953 & ~n48954;
  assign po981 = n2582 & ~n48955;
  assign po997 = ~pi33 & n33321;
  assign n48958 = n2924 & n5530;
  assign n48959 = pi951 & ~n48958;
  assign po986 = pi1092 & ~n48959;
  assign n48961 = ~pi832 & pi1091;
  assign n48962 = pi1162 & n48961;
  assign po989 = n5534 & n48962;
  assign n48964 = pi281 & ~n48945;
  assign po987 = ~n48946 & ~n48964;
  assign n48966 = pi833 & ~n2923;
  assign n48967 = ~n62394 & ~n48966;
  assign po1107 = n2887 & ~n3032;
  assign n48969 = pi24 & ~pi954;
  assign n48970 = pi786 & pi954;
  assign n48971 = ~pi786 & pi954;
  assign n48972 = ~pi24 & ~pi954;
  assign n48973 = ~n48971 & ~n48972;
  assign n48974 = ~n48969 & ~n48970;
  assign n48975 = pi1093 & pi1139;
  assign n48976 = pi920 & ~pi1093;
  assign n48977 = ~pi920 & ~pi1093;
  assign n48978 = pi1093 & ~pi1139;
  assign n48979 = ~n48977 & ~n48978;
  assign n48980 = ~n48975 & ~n48976;
  assign n48981 = pi1093 & pi1140;
  assign n48982 = pi921 & ~pi1093;
  assign n48983 = ~n48981 & ~n48982;
  assign n48984 = ~pi927 & ~pi1093;
  assign n48985 = pi1093 & ~pi1145;
  assign n48986 = pi1093 & pi1145;
  assign n48987 = pi927 & ~pi1093;
  assign n48988 = ~n48986 & ~n48987;
  assign n48989 = ~n48984 & ~n48985;
  assign n48990 = pi1093 & ~pi1136;
  assign n48991 = ~pi928 & ~pi1093;
  assign po1084 = ~n48990 & ~n48991;
  assign n48993 = ~pi929 & ~pi1093;
  assign n48994 = pi1093 & ~pi1144;
  assign n48995 = pi1093 & pi1144;
  assign n48996 = pi929 & ~pi1093;
  assign n48997 = ~n48995 & ~n48996;
  assign n48998 = ~n48993 & ~n48994;
  assign n48999 = ~pi930 & ~pi1093;
  assign n49000 = pi1093 & ~pi1134;
  assign n49001 = pi1093 & pi1134;
  assign n49002 = pi930 & ~pi1093;
  assign n49003 = ~n49001 & ~n49002;
  assign n49004 = ~n48999 & ~n49000;
  assign n49005 = pi1093 & pi1142;
  assign n49006 = pi932 & ~pi1093;
  assign n49007 = ~n49005 & ~n49006;
  assign n49008 = pi1093 & pi1137;
  assign n49009 = pi933 & ~pi1093;
  assign n49010 = ~n49008 & ~n49009;
  assign n49011 = pi1093 & pi1141;
  assign n49012 = pi935 & ~pi1093;
  assign n49013 = ~n49011 & ~n49012;
  assign n49014 = pi1093 & pi1135;
  assign n49015 = pi938 & ~pi1093;
  assign n49016 = ~n49014 & ~n49015;
  assign n49017 = ~pi939 & ~pi1093;
  assign n49018 = pi1093 & ~pi1146;
  assign n49019 = pi1093 & pi1146;
  assign n49020 = pi939 & ~pi1093;
  assign n49021 = ~n49019 & ~n49020;
  assign n49022 = ~n49017 & ~n49018;
  assign n49023 = pi1093 & pi1138;
  assign n49024 = pi940 & ~pi1093;
  assign n49025 = ~n49023 & ~n49024;
  assign n49026 = pi1093 & pi1143;
  assign n49027 = pi944 & ~pi1093;
  assign n49028 = ~pi944 & ~pi1093;
  assign n49029 = pi1093 & ~pi1143;
  assign n49030 = ~n49028 & ~n49029;
  assign n49031 = ~n49026 & ~n49027;
  assign n49032 = pi957 & pi1092;
  assign n49033 = ~pi31 & ~n49032;
  assign po1135 = pi824 & pi1092;
  assign n49035 = ~pi567 & pi1092;
  assign n49036 = ~pi230 & ~n49035;
  assign n49037 = ~pi1093 & n49035;
  assign n49038 = pi603 & n7224;
  assign n49039 = n13344 & n49038;
  assign n49040 = ~n8334 & n49039;
  assign n49041 = ~n63011 & n11313;
  assign n49042 = pi603 & ~n8135;
  assign n49043 = n7224 & ~n63011;
  assign n49044 = ~n63012 & n49043;
  assign n49045 = n49042 & n49044;
  assign n49046 = ~n63011 & n49038;
  assign n49047 = n11313 & n49046;
  assign n49048 = n49038 & n49041;
  assign n49049 = ~n11306 & n65086;
  assign n49050 = ~pi789 & ~n49037;
  assign n49051 = ~n65086 & n49050;
  assign n49052 = ~pi619 & n65086;
  assign n49053 = ~n49037 & ~n49052;
  assign n49054 = ~pi1159 & ~n49053;
  assign n49055 = pi619 & n65086;
  assign n49056 = ~n49037 & ~n49055;
  assign n49057 = pi1159 & ~n49056;
  assign n49058 = pi789 & ~n49057;
  assign n49059 = pi789 & ~n49054;
  assign n49060 = ~n49057 & n49059;
  assign n49061 = ~n49054 & n49058;
  assign n49062 = ~n49051 & ~n65087;
  assign n49063 = ~n49037 & ~n49049;
  assign n49064 = n8595 & ~n49037;
  assign n49065 = ~n8595 & n65088;
  assign n49066 = n8595 & n49037;
  assign n49067 = ~n49065 & ~n49066;
  assign n49068 = n65088 & ~n49064;
  assign n49069 = n8334 & ~n49037;
  assign n49070 = ~n65089 & ~n49069;
  assign n49071 = ~n8334 & n65089;
  assign n49072 = ~n49069 & ~n49071;
  assign n49073 = ~n8334 & ~n65089;
  assign n49074 = n8334 & n49037;
  assign n49075 = ~n49073 & ~n49074;
  assign n49076 = ~n49037 & ~n49040;
  assign n49077 = ~pi647 & n65090;
  assign n49078 = pi1157 & ~n49077;
  assign n49079 = pi680 & n7952;
  assign n49080 = ~n62964 & n49079;
  assign n49081 = ~n49037 & ~n49080;
  assign n49082 = n10106 & ~n49081;
  assign n49083 = n10206 & n49082;
  assign n49084 = ~n8257 & n49082;
  assign n49085 = ~n8303 & n49084;
  assign n49086 = n10207 & ~n49081;
  assign n49087 = ~n62892 & n65091;
  assign n49088 = ~pi647 & n49087;
  assign n49089 = ~pi1157 & ~n49037;
  assign n49090 = ~n49088 & n49089;
  assign n49091 = pi630 & ~n49090;
  assign n49092 = ~n49078 & n49091;
  assign n49093 = pi647 & n65090;
  assign n49094 = ~pi1157 & ~n49093;
  assign n49095 = pi647 & n49087;
  assign n49096 = pi1157 & ~n49037;
  assign n49097 = ~n49095 & n49096;
  assign n49098 = ~pi630 & ~n49097;
  assign n49099 = ~n49094 & n49098;
  assign n49100 = ~n49092 & ~n49099;
  assign n49101 = pi787 & ~n49100;
  assign n49102 = pi628 & n65091;
  assign n49103 = pi629 & n49039;
  assign n49104 = ~n49102 & ~n49103;
  assign n49105 = pi1156 & ~n49104;
  assign n49106 = ~pi628 & n65091;
  assign n49107 = ~pi629 & n49039;
  assign n49108 = ~n49106 & ~n49107;
  assign n49109 = ~pi1156 & ~n49108;
  assign n49110 = ~n49039 & ~n65091;
  assign n49111 = ~pi792 & ~n49110;
  assign n49112 = ~n49037 & ~n49111;
  assign n49113 = ~n49109 & n49112;
  assign n49114 = pi788 & ~n8524;
  assign n49115 = ~n8257 & n49114;
  assign n49116 = n49082 & n49115;
  assign n49117 = ~n49037 & ~n49116;
  assign n49118 = ~n8418 & ~n49117;
  assign n49119 = n11305 & n65086;
  assign n49120 = n8257 & ~n49037;
  assign n49121 = ~n62884 & n65087;
  assign n49122 = ~n49119 & n49120;
  assign n49123 = n62894 & n49082;
  assign n49124 = ~n65092 & n49123;
  assign n49125 = ~n49065 & ~n49124;
  assign n49126 = n49082 & ~n65092;
  assign n49127 = ~n65088 & ~n49126;
  assign n49128 = n62894 & ~n49127;
  assign n49129 = n12979 & n65088;
  assign n49130 = pi641 & n49084;
  assign n49131 = ~n49037 & ~n49130;
  assign n49132 = n8416 & ~n49131;
  assign n49133 = ~pi641 & n49084;
  assign n49134 = ~n49037 & ~n49133;
  assign n49135 = n8417 & ~n49134;
  assign n49136 = ~n49132 & ~n49135;
  assign n49137 = ~n49129 & n49136;
  assign n49138 = pi788 & ~n49137;
  assign n49139 = ~n49128 & ~n49138;
  assign n49140 = ~n49118 & n49125;
  assign n49141 = ~n63030 & ~n65093;
  assign n49142 = n8499 & ~n65089;
  assign n49143 = ~n49037 & ~n49102;
  assign n49144 = pi1156 & ~n49143;
  assign n49145 = ~pi629 & ~n49144;
  assign n49146 = ~pi629 & ~n49142;
  assign n49147 = ~n49144 & n49146;
  assign n49148 = ~n49142 & n49145;
  assign n49149 = n8498 & ~n65089;
  assign n49150 = ~n49037 & ~n49106;
  assign n49151 = ~pi1156 & ~n49150;
  assign n49152 = pi629 & ~n49151;
  assign n49153 = pi629 & ~n49149;
  assign n49154 = ~n49151 & n49153;
  assign n49155 = ~n49149 & n49152;
  assign n49156 = pi792 & ~n65095;
  assign n49157 = pi792 & ~n65094;
  assign n49158 = ~n65095 & n49157;
  assign n49159 = ~n65094 & n49156;
  assign n49160 = ~n49141 & ~n65096;
  assign n49161 = ~n49105 & n49113;
  assign n49162 = pi647 & n49091;
  assign n49163 = n8645 & ~n49096;
  assign n49164 = pi787 & ~n49163;
  assign n49165 = ~n49162 & n49164;
  assign n49166 = ~n65097 & ~n49165;
  assign n49167 = ~pi647 & ~n65097;
  assign n49168 = n49094 & ~n49167;
  assign n49169 = n49098 & ~n49168;
  assign n49170 = pi647 & ~n65097;
  assign n49171 = n49078 & ~n49170;
  assign n49172 = n49091 & ~n49171;
  assign n49173 = ~n49169 & ~n49172;
  assign n49174 = pi787 & ~n49173;
  assign n49175 = ~pi787 & ~n65097;
  assign n49176 = ~n49174 & ~n49175;
  assign n49177 = ~n49101 & ~n49166;
  assign n49178 = ~n11547 & ~n65098;
  assign n49179 = ~n11539 & n49037;
  assign n49180 = n29310 & n49039;
  assign n49181 = ~n49179 & ~n49180;
  assign n49182 = ~pi644 & ~n49181;
  assign n49183 = n11556 & n49087;
  assign n49184 = n29299 & n49039;
  assign n49185 = ~n49037 & ~n49184;
  assign n49186 = n11542 & ~n49185;
  assign n49187 = ~n49183 & ~n49186;
  assign n49188 = ~n49182 & n49187;
  assign n49189 = pi790 & ~n49188;
  assign n49190 = pi230 & ~n49189;
  assign n49191 = ~n49178 & n49190;
  assign n49192 = ~pi790 & ~n65098;
  assign n49193 = ~pi644 & ~n65098;
  assign n49194 = ~n10298 & n49087;
  assign n49195 = ~n49037 & ~n49194;
  assign n49196 = pi644 & ~n49195;
  assign n49197 = ~pi715 & ~n49196;
  assign n49198 = ~n49193 & n49197;
  assign n49199 = ~n8376 & n49073;
  assign n49200 = n8685 & ~n65089;
  assign n49201 = ~pi644 & n65099;
  assign n49202 = pi715 & ~n49037;
  assign n49203 = ~n49201 & n49202;
  assign n49204 = ~n49198 & ~n49203;
  assign n49205 = ~pi1160 & ~n49204;
  assign n49206 = pi644 & n65098;
  assign n49207 = ~pi644 & n49195;
  assign n49208 = pi715 & ~n49207;
  assign n49209 = ~n49206 & n49208;
  assign n49210 = pi644 & n65099;
  assign n49211 = ~n49037 & ~n49210;
  assign n49212 = ~pi715 & ~n49211;
  assign n49213 = pi1160 & ~n49212;
  assign n49214 = ~n49209 & n49213;
  assign n49215 = pi790 & ~n49214;
  assign n49216 = ~pi1160 & ~n49203;
  assign n49217 = ~n49198 & n49216;
  assign n49218 = pi644 & ~n65098;
  assign n49219 = ~pi644 & ~n49195;
  assign n49220 = pi715 & ~n49219;
  assign n49221 = ~n49218 & n49220;
  assign n49222 = ~pi715 & ~n49037;
  assign n49223 = ~n49210 & n49222;
  assign n49224 = pi1160 & ~n49223;
  assign n49225 = ~n49221 & n49224;
  assign n49226 = ~n49217 & ~n49225;
  assign n49227 = pi790 & ~n49226;
  assign n49228 = ~n49205 & n49215;
  assign n49229 = ~n49192 & ~n65100;
  assign n49230 = pi230 & ~n49229;
  assign n49231 = ~pi230 & n49035;
  assign n49232 = ~n49230 & ~n49231;
  assign n49233 = ~n49036 & ~n49191;
  assign n49234 = pi243 & ~pi1091;
  assign n49235 = ~pi83 & ~pi85;
  assign n49236 = pi314 & ~n49235;
  assign n49237 = pi802 & n49236;
  assign n49238 = pi276 & n49237;
  assign n49239 = ~pi1091 & ~n49238;
  assign n49240 = pi271 & ~n49239;
  assign n49241 = ~pi1091 & ~n49240;
  assign n49242 = pi273 & ~n49241;
  assign n49243 = ~pi1091 & ~n49242;
  assign n49244 = ~pi200 & ~n49243;
  assign n49245 = pi199 & ~n49243;
  assign n49246 = ~pi81 & n49235;
  assign n49247 = pi314 & ~n49246;
  assign n49248 = pi802 & n49247;
  assign n49249 = pi276 & n49248;
  assign n49250 = ~pi1091 & n49249;
  assign n49251 = pi271 & n49250;
  assign n49252 = pi273 & n49251;
  assign n49253 = ~n49242 & ~n49252;
  assign n49254 = ~pi1091 & n49253;
  assign n49255 = ~pi199 & ~n49254;
  assign n49256 = ~n49245 & ~n49255;
  assign n49257 = n49250 & ~n49256;
  assign n49258 = ~pi299 & ~n49257;
  assign n49259 = ~n49245 & n49258;
  assign n49260 = ~n49244 & n49259;
  assign n49261 = pi299 & ~n49252;
  assign n49262 = ~n49260 & ~n49261;
  assign n49263 = ~n49234 & ~n49262;
  assign n49264 = pi299 & n49243;
  assign n49265 = ~n49252 & n49264;
  assign n49266 = ~pi200 & ~n49250;
  assign n49267 = ~n49256 & ~n49266;
  assign n49268 = ~pi299 & ~n49267;
  assign n49269 = ~n49255 & n49268;
  assign n49270 = ~n49260 & ~n49269;
  assign n49271 = ~n49265 & n49270;
  assign n49272 = ~pi243 & ~n49271;
  assign n49273 = ~n49245 & n49268;
  assign n49274 = ~n49261 & ~n49273;
  assign n49275 = ~n49244 & n49258;
  assign n49276 = ~n49255 & n49275;
  assign n49277 = pi243 & ~n49276;
  assign n49278 = n49274 & n49277;
  assign n49279 = ~n49272 & ~n49278;
  assign n49280 = ~pi1155 & ~n49279;
  assign n49281 = ~pi1091 & n49238;
  assign n49282 = pi271 & n49281;
  assign n49283 = pi273 & n49282;
  assign n49284 = pi299 & ~n49283;
  assign n49285 = ~n49276 & ~n49284;
  assign n49286 = ~n49273 & n49285;
  assign n49287 = ~n49264 & ~n49275;
  assign n49288 = pi243 & ~n49287;
  assign n49289 = ~n49286 & n49288;
  assign n49290 = pi1155 & ~n49289;
  assign n49291 = ~n49265 & ~n49276;
  assign n49292 = pi1155 & n49291;
  assign n49293 = ~n49290 & ~n49292;
  assign n49294 = ~n49261 & ~n49268;
  assign n49295 = ~pi243 & n49294;
  assign n49296 = ~n49265 & ~n49268;
  assign n49297 = n49262 & n49296;
  assign n49298 = ~n49260 & n49294;
  assign n49299 = ~pi243 & n65102;
  assign n49300 = ~n49260 & n49295;
  assign n49301 = ~n49293 & ~n65103;
  assign n49302 = ~n49280 & ~n49301;
  assign n49303 = ~n49263 & n49302;
  assign n49304 = pi1156 & ~n49303;
  assign n49305 = ~n49264 & ~n49269;
  assign n49306 = ~pi243 & ~n49305;
  assign n49307 = ~pi1155 & ~n49306;
  assign n49308 = ~n49258 & ~n49261;
  assign n49309 = ~pi1155 & n49308;
  assign n49310 = ~n49307 & ~n49309;
  assign n49311 = ~n49259 & ~n49261;
  assign n49312 = ~n49275 & n49311;
  assign n49313 = ~n49261 & ~n49275;
  assign n49314 = pi243 & n49313;
  assign n49315 = ~n49259 & n49314;
  assign n49316 = pi243 & n49312;
  assign n49317 = ~n49310 & ~n65104;
  assign n49318 = ~pi1156 & ~n49317;
  assign n49319 = ~pi243 & ~n49296;
  assign n49320 = pi1155 & ~n49319;
  assign n49321 = ~n49314 & n49320;
  assign n49322 = n49318 & ~n49321;
  assign n49323 = pi1157 & ~n49322;
  assign n49324 = ~n49304 & n49323;
  assign n49325 = pi243 & n49308;
  assign n49326 = ~pi243 & ~pi1091;
  assign n49327 = ~n49258 & ~n49284;
  assign n49328 = n49326 & ~n49327;
  assign n49329 = ~pi1155 & ~n49328;
  assign n49330 = ~n49309 & ~n49329;
  assign n49331 = ~n49325 & ~n49330;
  assign n49332 = ~pi1156 & ~n49331;
  assign n49333 = pi1155 & ~n49234;
  assign n49334 = n49245 & n49333;
  assign n49335 = ~n49321 & ~n49334;
  assign n49336 = n49332 & n49335;
  assign n49337 = ~n49255 & n49258;
  assign n49338 = ~n49265 & ~n49337;
  assign n49339 = pi243 & ~n49338;
  assign n49340 = ~pi243 & n49311;
  assign n49341 = ~n49339 & ~n49340;
  assign n49342 = ~pi1155 & n49313;
  assign n49343 = ~n49250 & n49342;
  assign n49344 = pi1156 & ~n49343;
  assign n49345 = pi1156 & n49341;
  assign n49346 = ~n49343 & n49345;
  assign n49347 = n49341 & n49344;
  assign n49348 = ~pi1157 & ~n65105;
  assign n49349 = ~n49336 & n49348;
  assign n49350 = pi211 & ~n49349;
  assign n49351 = ~n49324 & n49350;
  assign n49352 = pi1156 & ~n49302;
  assign n49353 = ~n49265 & ~n49275;
  assign n49354 = pi243 & ~n49353;
  assign n49355 = ~n49295 & ~n49354;
  assign n49356 = n49318 & n49355;
  assign n49357 = pi1157 & ~n49356;
  assign n49358 = ~n49352 & n49357;
  assign n49359 = ~pi1155 & n49353;
  assign n49360 = ~n49294 & n49359;
  assign n49361 = n65105 & ~n49360;
  assign n49362 = n49341 & n49355;
  assign n49363 = pi1155 & ~n49362;
  assign n49364 = n49332 & ~n49363;
  assign n49365 = ~pi1157 & ~n49364;
  assign n49366 = ~pi1157 & ~n49361;
  assign n49367 = ~n49364 & n49366;
  assign n49368 = ~n49361 & n49365;
  assign n49369 = ~pi211 & ~n65106;
  assign n49370 = ~n49358 & n49369;
  assign n49371 = ~pi219 & ~n49370;
  assign n49372 = ~n49351 & n49371;
  assign n49373 = pi253 & pi254;
  assign n49374 = pi267 & n49373;
  assign n49375 = ~pi263 & n49374;
  assign n49376 = ~n49260 & ~n49264;
  assign n49377 = ~pi243 & n49376;
  assign n49378 = ~n49268 & ~n49284;
  assign n49379 = n49377 & n49378;
  assign n49380 = n49290 & ~n49379;
  assign n49381 = pi243 & ~n49286;
  assign n49382 = ~n49377 & ~n49381;
  assign n49383 = ~n49263 & ~n49306;
  assign n49384 = ~n49382 & n49383;
  assign n49385 = ~pi1155 & ~n49384;
  assign n49386 = ~n49380 & ~n49385;
  assign n49387 = pi1156 & ~n49386;
  assign n49388 = ~pi211 & pi1157;
  assign n49389 = ~n49269 & ~n49284;
  assign n49390 = ~pi243 & ~n49389;
  assign n49391 = pi243 & ~n49259;
  assign n49392 = ~pi1155 & ~n49391;
  assign n49393 = ~n49390 & n49392;
  assign n49394 = ~pi243 & pi1155;
  assign n49395 = n49378 & n49394;
  assign n49396 = ~pi1156 & ~n49395;
  assign n49397 = ~n49288 & n49396;
  assign n49398 = ~n49393 & n49397;
  assign n49399 = n49388 & ~n49398;
  assign n49400 = ~n49387 & n49399;
  assign n49401 = pi243 & n49285;
  assign n49402 = n49320 & ~n49401;
  assign n49403 = ~n49307 & ~n49402;
  assign n49404 = ~n49382 & ~n49403;
  assign n49405 = pi1156 & ~n49404;
  assign n49406 = pi211 & pi1157;
  assign n49407 = ~n49275 & ~n49284;
  assign n49408 = pi243 & n49407;
  assign n49409 = ~n49319 & ~n49408;
  assign n49410 = pi1155 & ~n49409;
  assign n49411 = ~n49259 & n49407;
  assign n49412 = pi243 & n49411;
  assign n49413 = n49391 & n49407;
  assign n49414 = ~n49306 & ~n65107;
  assign n49415 = ~n49410 & n49414;
  assign n49416 = ~pi1156 & ~n49415;
  assign n49417 = n49406 & ~n49416;
  assign n49418 = ~n49405 & n49417;
  assign n49419 = ~n49284 & ~n49337;
  assign n49420 = pi1155 & n49419;
  assign n49421 = ~n49268 & n49419;
  assign n49422 = ~n49420 & ~n49421;
  assign n49423 = pi243 & ~n49422;
  assign n49424 = ~n49259 & ~n49264;
  assign n49425 = ~pi243 & ~n49424;
  assign n49426 = ~n49343 & n49425;
  assign n49427 = ~n49423 & ~n49426;
  assign n49428 = pi1156 & ~n49427;
  assign n49429 = ~n49337 & n49408;
  assign n49430 = ~n49264 & ~n49273;
  assign n49431 = ~pi243 & ~n49430;
  assign n49432 = pi1155 & ~n49431;
  assign n49433 = ~n49429 & n49432;
  assign n49434 = pi243 & n49327;
  assign n49435 = n49329 & ~n49434;
  assign n49436 = ~pi1156 & ~n49435;
  assign n49437 = ~n49433 & n49436;
  assign n49438 = ~pi1157 & ~n49437;
  assign n49439 = ~n49428 & n49438;
  assign n49440 = ~n49418 & ~n49439;
  assign n49441 = ~n49400 & n49440;
  assign n49442 = pi219 & ~n49441;
  assign n49443 = n49375 & ~n49442;
  assign n49444 = ~n49372 & n49443;
  assign n49445 = pi199 & pi200;
  assign n49446 = ~pi1155 & n39538;
  assign n49447 = ~n49445 & ~n65108;
  assign n49448 = ~pi299 & pi1091;
  assign n49449 = n49447 & n49448;
  assign n49450 = ~n49326 & ~n49449;
  assign n49451 = pi1156 & ~n49450;
  assign n49452 = ~pi299 & n49445;
  assign n49453 = pi1156 & ~n49452;
  assign n49454 = pi1091 & ~n48497;
  assign n49455 = n49453 & n49454;
  assign n49456 = ~n49451 & ~n49455;
  assign n49457 = pi199 & ~pi200;
  assign n49458 = ~pi299 & n49457;
  assign n49459 = pi1091 & ~n49458;
  assign n49460 = ~n49234 & ~n49459;
  assign n49461 = ~pi200 & ~pi299;
  assign n49462 = ~pi1155 & ~n49326;
  assign n49463 = ~n49234 & ~n49462;
  assign n49464 = n49461 & n49463;
  assign n49465 = ~n49460 & ~n49464;
  assign n49466 = ~pi1156 & ~n49465;
  assign n49467 = pi1157 & ~n49466;
  assign n49468 = n49456 & n49467;
  assign n49469 = ~n49454 & n49463;
  assign n49470 = ~pi1156 & ~n49469;
  assign n49471 = pi199 & pi1091;
  assign n49472 = ~pi299 & n49471;
  assign n49473 = n49333 & ~n49472;
  assign n49474 = pi1156 & ~n49473;
  assign n49475 = ~pi1155 & ~n49234;
  assign n49476 = ~n48474 & n49448;
  assign n49477 = n49475 & ~n49476;
  assign n49478 = n49474 & ~n49477;
  assign n49479 = ~n49470 & ~n49478;
  assign n49480 = ~pi1157 & ~n49479;
  assign n49481 = pi211 & ~n49480;
  assign n49482 = n49456 & ~n49466;
  assign n49483 = pi1157 & ~n49482;
  assign n49484 = ~pi1157 & ~n49478;
  assign n49485 = ~pi1157 & ~n49470;
  assign n49486 = ~n49478 & n49485;
  assign n49487 = ~n49470 & n49484;
  assign n49488 = ~n49483 & ~n65109;
  assign n49489 = pi211 & ~n49488;
  assign n49490 = ~n49468 & n49481;
  assign n49491 = n49450 & n49474;
  assign n49492 = ~pi1155 & n49460;
  assign n49493 = pi200 & pi1091;
  assign n49494 = pi200 & ~pi299;
  assign n49495 = pi1091 & n49494;
  assign n49496 = ~pi299 & n49493;
  assign n49497 = n49333 & ~n65111;
  assign n49498 = ~pi1156 & ~n49497;
  assign n49499 = ~n49492 & n49498;
  assign n49500 = ~n49491 & ~n49499;
  assign n49501 = pi1157 & ~n49500;
  assign n49502 = pi1091 & ~n48475;
  assign n49503 = n49475 & ~n49502;
  assign n49504 = ~n49473 & ~n49503;
  assign n49505 = pi200 & ~pi1156;
  assign n49506 = n49448 & n49505;
  assign n49507 = ~n49504 & ~n49506;
  assign n49508 = ~pi1157 & ~n49507;
  assign n49509 = ~pi211 & ~n49508;
  assign n49510 = ~n49501 & n49509;
  assign n49511 = ~n65110 & ~n49510;
  assign n49512 = ~pi219 & ~n49511;
  assign n49513 = n49406 & ~n49451;
  assign n49514 = ~n49466 & n49513;
  assign n49515 = pi219 & ~n49514;
  assign n49516 = pi299 & pi1091;
  assign n49517 = n49507 & ~n49516;
  assign n49518 = ~pi1157 & ~n49517;
  assign n49519 = ~pi299 & ~n49457;
  assign n49520 = pi1091 & n49519;
  assign n49521 = n49475 & ~n49520;
  assign n49522 = ~n49497 & ~n49521;
  assign n49523 = ~pi1156 & ~n49522;
  assign n49524 = n49388 & ~n49523;
  assign n49525 = n49456 & n49524;
  assign n49526 = ~n49518 & ~n49525;
  assign n49527 = pi219 & ~n49518;
  assign n49528 = ~n49514 & ~n49525;
  assign n49529 = n49527 & n49528;
  assign n49530 = n49515 & n49526;
  assign n49531 = ~n49512 & ~n65112;
  assign n49532 = ~n49375 & ~n49531;
  assign n49533 = n62455 & ~n49532;
  assign n49534 = ~n49444 & n49533;
  assign n49535 = pi272 & pi283;
  assign n49536 = pi275 & n49535;
  assign n49537 = pi268 & n49536;
  assign n49538 = pi243 & n49254;
  assign n49539 = n49234 & n49253;
  assign n49540 = ~pi243 & n49252;
  assign n49541 = pi211 & pi1156;
  assign n49542 = ~pi211 & pi1155;
  assign n49543 = ~n49541 & ~n49542;
  assign n49544 = pi1091 & n49543;
  assign n49545 = ~n49540 & ~n49544;
  assign n49546 = ~n65113 & n49545;
  assign n49547 = ~pi219 & ~n49546;
  assign n49548 = ~pi243 & n49243;
  assign n49549 = pi243 & n49283;
  assign n49550 = ~n49234 & n49388;
  assign n49551 = ~n49281 & n49550;
  assign n49552 = pi219 & ~n49551;
  assign n49553 = ~n49549 & n49552;
  assign n49554 = ~n49548 & n49553;
  assign n49555 = n49375 & ~n49554;
  assign n49556 = ~n49549 & ~n49551;
  assign n49557 = ~n49548 & n49556;
  assign n49558 = pi219 & ~n49557;
  assign n49559 = ~pi219 & ~n49544;
  assign n49560 = ~n49540 & n49559;
  assign n49561 = ~n65113 & n49560;
  assign n49562 = ~n49558 & ~n49561;
  assign n49563 = n49375 & ~n49562;
  assign n49564 = ~n49547 & n49555;
  assign n49565 = ~pi219 & ~n49543;
  assign n49566 = pi219 & n49388;
  assign n49567 = pi1157 & n39423;
  assign n49568 = ~n49565 & ~n65115;
  assign n49569 = pi1091 & ~n49568;
  assign n49570 = ~n49326 & ~n49569;
  assign n49571 = ~n49375 & ~n49570;
  assign n49572 = ~n62455 & ~n49571;
  assign n49573 = ~n65114 & n49572;
  assign n49574 = n49537 & ~n49573;
  assign n49575 = ~n49534 & n49574;
  assign n49576 = n62455 & n49531;
  assign n49577 = ~n62455 & n49570;
  assign n49578 = ~n49537 & ~n49577;
  assign n49579 = ~n49576 & n49578;
  assign n49580 = ~pi230 & ~n49579;
  assign n49581 = ~n49575 & n49580;
  assign n49582 = ~pi200 & pi1157;
  assign n49583 = pi199 & ~n49582;
  assign n49584 = ~n65108 & ~n49505;
  assign n49585 = ~n49583 & n49584;
  assign n49586 = n65014 & n49585;
  assign n49587 = ~n65014 & ~n49568;
  assign n49588 = pi230 & ~n49587;
  assign n49589 = pi230 & ~n49586;
  assign n49590 = ~n49587 & n49589;
  assign n49591 = ~n49586 & n49588;
  assign po400 = ~n49581 & ~n65116;
  assign n49593 = pi1154 & ~n39539;
  assign n49594 = pi200 & ~pi1155;
  assign n49595 = ~pi299 & ~n49445;
  assign n49596 = pi199 & pi1156;
  assign n49597 = ~pi200 & ~n49596;
  assign n49598 = ~n39538 & ~n49445;
  assign n49599 = ~pi299 & n49598;
  assign n49600 = ~pi1156 & ~n49494;
  assign n49601 = n49599 & ~n49600;
  assign n49602 = n49595 & ~n49597;
  assign n49603 = ~n49594 & n65117;
  assign n49604 = ~n49593 & ~n49603;
  assign n49605 = ~pi211 & ~n49604;
  assign n49606 = ~pi219 & ~n49605;
  assign n49607 = pi299 & pi1155;
  assign n49608 = ~pi199 & pi1155;
  assign n49609 = pi200 & ~n49608;
  assign n49610 = ~pi299 & ~n49609;
  assign n49611 = ~pi199 & pi1154;
  assign n49612 = n49597 & ~n49611;
  assign n49613 = pi1156 & n49457;
  assign n49614 = ~pi199 & ~n49594;
  assign n49615 = ~pi200 & ~pi1154;
  assign n49616 = n49614 & ~n49615;
  assign n49617 = ~n49613 & ~n49616;
  assign n49618 = ~pi299 & ~n49617;
  assign n49619 = ~pi299 & pi1155;
  assign n49620 = n49494 & n49608;
  assign n49621 = n48474 & n49619;
  assign n49622 = ~pi1154 & ~n65119;
  assign n49623 = n48567 & ~n49594;
  assign n49624 = ~n49622 & n49623;
  assign n49625 = ~pi1156 & ~n49624;
  assign n49626 = ~pi199 & ~pi1154;
  assign n49627 = ~pi200 & n49626;
  assign n49628 = n49610 & ~n65120;
  assign n49629 = ~n49625 & n49628;
  assign n49630 = n49610 & ~n49612;
  assign n49631 = ~n49607 & ~n65118;
  assign n49632 = pi211 & ~n49631;
  assign n49633 = n49606 & ~n49632;
  assign n49634 = pi1156 & n48498;
  assign n49635 = pi219 & ~n49634;
  assign n49636 = pi1154 & ~n49609;
  assign n49637 = pi1156 & ~n49636;
  assign n49638 = ~pi299 & ~n49637;
  assign n49639 = n39539 & ~n49609;
  assign n49640 = ~pi1154 & n49639;
  assign n49641 = ~n48498 & ~n49640;
  assign n49642 = ~n49638 & n49641;
  assign n49643 = pi1156 & ~n49642;
  assign n49644 = ~n49593 & ~n65119;
  assign n49645 = n49638 & ~n49644;
  assign n49646 = pi219 & ~n49645;
  assign n49647 = ~n49643 & n49646;
  assign n49648 = ~n65118 & n49635;
  assign n49649 = n62455 & ~n65121;
  assign n49650 = ~n49633 & n49649;
  assign n49651 = ~pi211 & pi1156;
  assign n49652 = pi219 & ~n49651;
  assign n49653 = ~pi211 & pi1154;
  assign n49654 = pi211 & pi1155;
  assign n49655 = ~pi219 & ~n49654;
  assign n49656 = ~n49653 & n49655;
  assign n49657 = ~n49652 & ~n49656;
  assign n49658 = ~n62455 & n49657;
  assign n49659 = pi230 & ~n49658;
  assign n49660 = ~n49650 & n49659;
  assign n49661 = ~pi1091 & ~n49419;
  assign n49662 = ~pi1155 & n49661;
  assign n49663 = ~n49338 & n49662;
  assign n49664 = pi1155 & ~n49262;
  assign n49665 = ~pi1154 & ~n49664;
  assign n49666 = ~n49663 & n49665;
  assign n49667 = ~pi1156 & ~n49666;
  assign n49668 = pi1155 & ~n49376;
  assign n49669 = ~pi1154 & ~n49668;
  assign n49670 = ~n49662 & n49669;
  assign n49671 = pi1155 & ~n49311;
  assign n49672 = pi1154 & ~n49671;
  assign n49673 = n49274 & n49672;
  assign n49674 = ~n49670 & ~n49673;
  assign n49675 = n49667 & n49674;
  assign n49676 = ~pi1155 & n49305;
  assign n49677 = ~n49261 & n49270;
  assign n49678 = ~n49676 & ~n49677;
  assign n49679 = ~pi1154 & ~n49678;
  assign n49680 = pi1156 & ~n49679;
  assign n49681 = n49305 & n49669;
  assign n49682 = ~n49266 & n49673;
  assign n49683 = ~n49681 & ~n49682;
  assign n49684 = n49680 & n49683;
  assign n49685 = ~pi211 & ~n49684;
  assign n49686 = ~pi211 & ~n49675;
  assign n49687 = ~n49684 & n49686;
  assign n49688 = ~n49675 & n49685;
  assign n49689 = ~n49265 & ~n49273;
  assign n49690 = n49672 & n49689;
  assign n49691 = n49667 & ~n49690;
  assign n49692 = n49296 & n49672;
  assign n49693 = n49680 & ~n49692;
  assign n49694 = pi211 & ~n49693;
  assign n49695 = pi211 & ~n49691;
  assign n49696 = ~n49693 & n49695;
  assign n49697 = ~n49691 & n49694;
  assign n49698 = ~pi219 & ~n65123;
  assign n49699 = ~pi219 & ~n65122;
  assign n49700 = ~n65123 & n49699;
  assign n49701 = ~n65122 & n49698;
  assign n49702 = pi1155 & n49260;
  assign n49703 = pi1154 & n49430;
  assign n49704 = ~n49702 & n49703;
  assign n49705 = ~n49670 & ~n49704;
  assign n49706 = ~pi1156 & ~n49705;
  assign n49707 = ~n49268 & n49704;
  assign n49708 = ~n49681 & ~n49707;
  assign n49709 = n49541 & ~n49708;
  assign n49710 = ~pi1154 & n49419;
  assign n49711 = ~n49378 & ~n49710;
  assign n49712 = n49651 & ~n49702;
  assign n49713 = ~n49711 & n49712;
  assign n49714 = pi219 & ~n49713;
  assign n49715 = ~n49709 & n49714;
  assign n49716 = ~n49706 & n49714;
  assign n49717 = ~n49709 & n49716;
  assign n49718 = ~n49706 & n49715;
  assign n49719 = ~pi263 & ~n65125;
  assign n49720 = ~n65124 & n49719;
  assign n49721 = pi1156 & n49312;
  assign n49722 = ~n49268 & n49338;
  assign n49723 = n49654 & n49722;
  assign n49724 = n49294 & ~n49337;
  assign n49725 = n49542 & n49724;
  assign n49726 = ~n49309 & ~n49725;
  assign n49727 = ~n49723 & n49726;
  assign n49728 = ~n49721 & n49727;
  assign n49729 = ~pi1154 & ~n49728;
  assign n49730 = ~n49292 & ~n49359;
  assign n49731 = ~n49269 & ~n49730;
  assign n49732 = ~pi1156 & ~n49731;
  assign n49733 = pi211 & n49342;
  assign n49734 = ~pi211 & n49359;
  assign n49735 = ~n49292 & ~n49734;
  assign n49736 = ~n49733 & n49735;
  assign n49737 = pi1154 & ~n49736;
  assign n49738 = ~n49732 & n49737;
  assign n49739 = ~n49729 & ~n49738;
  assign n49740 = pi1154 & ~n49292;
  assign n49741 = ~n49342 & n49740;
  assign n49742 = ~pi1154 & ~n49309;
  assign n49743 = pi1155 & n49722;
  assign n49744 = n49742 & ~n49743;
  assign n49745 = ~n49359 & n49740;
  assign n49746 = pi1154 & n49269;
  assign n49747 = ~pi1156 & ~n49746;
  assign n49748 = ~n49745 & n49747;
  assign n49749 = ~pi1156 & ~n49748;
  assign n49750 = ~n49744 & ~n49749;
  assign n49751 = ~n49721 & ~n49750;
  assign n49752 = ~n49741 & ~n49751;
  assign n49753 = pi211 & ~n49752;
  assign n49754 = pi1155 & n49724;
  assign n49755 = n49742 & ~n49754;
  assign n49756 = n49748 & ~n49755;
  assign n49757 = ~n49312 & n49755;
  assign n49758 = pi1156 & ~n49757;
  assign n49759 = ~n49745 & n49758;
  assign n49760 = ~pi211 & ~n49759;
  assign n49761 = ~n49756 & n49760;
  assign n49762 = ~pi219 & ~n49761;
  assign n49763 = ~n49753 & n49762;
  assign n49764 = ~pi219 & ~n49739;
  assign n49765 = ~n49287 & ~n49420;
  assign n49766 = pi1154 & n49273;
  assign n49767 = ~n49286 & ~n49766;
  assign n49768 = ~n49765 & ~n49767;
  assign n49769 = ~n49337 & n49768;
  assign n49770 = ~pi1156 & ~n49769;
  assign n49771 = n49541 & ~n49768;
  assign n49772 = ~n49275 & n49424;
  assign n49773 = ~pi1155 & ~n49772;
  assign n49774 = ~n49276 & n49430;
  assign n49775 = pi1155 & ~n49774;
  assign n49776 = ~pi1154 & ~n49775;
  assign n49777 = ~pi1154 & ~n49773;
  assign n49778 = ~n49775 & n49777;
  assign n49779 = ~n49773 & n49776;
  assign n49780 = pi1154 & ~n49765;
  assign n49781 = n49651 & ~n49780;
  assign n49782 = ~n65127 & n49781;
  assign n49783 = pi219 & ~n49782;
  assign n49784 = pi219 & ~n49771;
  assign n49785 = ~n49782 & n49784;
  assign n49786 = ~n49771 & n49783;
  assign n49787 = ~n49770 & n65128;
  assign n49788 = pi263 & ~n49787;
  assign n49789 = ~n65126 & n49788;
  assign n49790 = n49374 & ~n49789;
  assign n49791 = n49374 & ~n49720;
  assign n49792 = ~n49789 & n49791;
  assign n49793 = ~n49720 & n49790;
  assign n49794 = pi1155 & ~n49452;
  assign n49795 = n65111 & ~n49794;
  assign n49796 = pi1091 & ~n49599;
  assign n49797 = ~pi1154 & n49796;
  assign n49798 = ~n49795 & ~n49797;
  assign n49799 = ~pi211 & ~n49798;
  assign n49800 = ~pi299 & ~n48474;
  assign n49801 = pi1155 & ~n49800;
  assign n49802 = pi211 & pi1091;
  assign n49803 = n49461 & ~n49626;
  assign n49804 = n49802 & ~n49803;
  assign n49805 = ~n49801 & n49804;
  assign n49806 = pi1156 & ~n49805;
  assign n49807 = ~n49799 & n49806;
  assign n49808 = pi1091 & ~pi1154;
  assign n49809 = ~n49454 & ~n49808;
  assign n49810 = ~n49801 & ~n49809;
  assign n49811 = pi211 & n49810;
  assign n49812 = ~pi211 & pi1091;
  assign n49813 = ~n65119 & n49812;
  assign n49814 = n49644 & n49812;
  assign n49815 = ~n49593 & n49813;
  assign n49816 = ~pi1156 & ~n65130;
  assign n49817 = ~n49811 & n49816;
  assign n49818 = ~n49807 & ~n49817;
  assign n49819 = ~n49799 & ~n49805;
  assign n49820 = pi1156 & ~n49819;
  assign n49821 = ~n49811 & ~n65130;
  assign n49822 = ~pi1156 & ~n49821;
  assign n49823 = ~pi219 & ~n49822;
  assign n49824 = ~n49820 & n49823;
  assign n49825 = ~pi219 & ~n49818;
  assign n49826 = ~n49516 & n49798;
  assign n49827 = n49541 & ~n49826;
  assign n49828 = ~pi1156 & ~n65119;
  assign n49829 = ~n49809 & n49828;
  assign n49830 = pi200 & n49608;
  assign n49831 = ~pi1155 & ~n49519;
  assign n49832 = ~pi299 & ~n49598;
  assign n49833 = pi1155 & ~n49832;
  assign n49834 = ~n49831 & ~n49833;
  assign n49835 = n49519 & ~n49830;
  assign n49836 = ~pi1154 & ~n65132;
  assign n49837 = n49494 & ~n49608;
  assign n49838 = pi1154 & ~n49837;
  assign n49839 = pi1091 & n49651;
  assign n49840 = ~n49838 & n49839;
  assign n49841 = ~n49836 & n49840;
  assign n49842 = pi219 & ~n49841;
  assign n49843 = pi219 & ~n49829;
  assign n49844 = ~n49841 & n49843;
  assign n49845 = ~n49829 & n49842;
  assign n49846 = ~n49827 & n65133;
  assign n49847 = ~n65131 & ~n49846;
  assign n49848 = ~pi263 & ~n49847;
  assign n49849 = ~pi1155 & ~n39539;
  assign n49850 = n49836 & ~n49849;
  assign n49851 = pi1155 & ~n48570;
  assign n49852 = ~n49461 & ~n49851;
  assign n49853 = pi1154 & ~n49852;
  assign n49854 = pi1156 & ~n49853;
  assign n49855 = ~n49850 & n49854;
  assign n49856 = ~pi1156 & n49810;
  assign n49857 = pi211 & ~n49856;
  assign n49858 = ~n49855 & n49857;
  assign n49859 = n49606 & ~n49858;
  assign n49860 = pi263 & pi1091;
  assign n49861 = ~n65121 & n49860;
  assign n49862 = ~n49859 & n49861;
  assign n49863 = ~n49848 & ~n49862;
  assign n49864 = ~n49374 & ~n49863;
  assign n49865 = n62455 & ~n49864;
  assign n49866 = ~n65129 & n49865;
  assign n49867 = pi211 & n49243;
  assign n49868 = ~pi211 & ~n49808;
  assign n49869 = ~n49654 & ~n49868;
  assign n49870 = ~n49867 & n49869;
  assign n49871 = ~n49252 & ~n49870;
  assign n49872 = ~pi219 & ~n49871;
  assign n49873 = pi219 & ~n49243;
  assign n49874 = ~pi211 & ~n49281;
  assign n49875 = n49873 & ~n49874;
  assign n49876 = ~pi263 & ~n49875;
  assign n49877 = ~n49872 & n49876;
  assign n49878 = ~pi219 & ~n49252;
  assign n49879 = pi1154 & n49812;
  assign n49880 = ~n49654 & ~n49879;
  assign n49881 = ~n49867 & ~n49880;
  assign n49882 = n49878 & ~n49881;
  assign n49883 = ~pi211 & ~n49243;
  assign n49884 = pi211 & n49283;
  assign n49885 = pi219 & ~n49884;
  assign n49886 = ~n49883 & n49885;
  assign n49887 = pi263 & ~n49886;
  assign n49888 = ~n49882 & n49887;
  assign n49889 = ~n49877 & ~n49888;
  assign n49890 = pi1091 & n49652;
  assign n49891 = n49374 & ~n49890;
  assign n49892 = ~n49889 & n49891;
  assign n49893 = pi1091 & ~n49657;
  assign n49894 = pi263 & ~pi1091;
  assign n49895 = ~n49893 & ~n49894;
  assign n49896 = ~n49374 & n49895;
  assign n49897 = ~n62455 & ~n49896;
  assign n49898 = ~n49892 & n49897;
  assign n49899 = n49537 & ~n49898;
  assign n49900 = ~n49866 & n49899;
  assign n49901 = n62455 & n49863;
  assign n49902 = ~n62455 & ~n49895;
  assign n49903 = ~n49537 & ~n49902;
  assign n49904 = ~n49901 & n49903;
  assign n49905 = ~pi230 & ~n49904;
  assign n49906 = ~n49900 & n49905;
  assign po420 = ~n49660 & ~n49906;
  assign n49908 = ~pi1153 & n49338;
  assign n49909 = ~n49689 & ~n49908;
  assign n49910 = n49376 & ~n49909;
  assign n49911 = pi1154 & ~n49910;
  assign n49912 = ~pi1153 & ~n49661;
  assign n49913 = ~pi1154 & ~n49430;
  assign n49914 = ~n49912 & n49913;
  assign n49915 = ~pi1155 & ~n49914;
  assign n49916 = ~n49911 & n49915;
  assign n49917 = ~pi211 & ~n49252;
  assign n49918 = ~pi211 & n49261;
  assign n49919 = pi299 & n49917;
  assign n49920 = n49689 & ~n65134;
  assign n49921 = ~n49260 & n49305;
  assign n49922 = n49920 & n49921;
  assign n49923 = ~n49389 & ~n49922;
  assign n49924 = pi1153 & ~n49296;
  assign n49925 = pi1155 & ~n49924;
  assign n49926 = n49260 & ~n49710;
  assign n49927 = n49925 & ~n49926;
  assign n49928 = ~n49923 & n49927;
  assign n49929 = pi267 & ~n49928;
  assign n49930 = ~n49916 & n49929;
  assign n49931 = ~pi1153 & ~n49327;
  assign n49932 = ~n49275 & n49419;
  assign n49933 = ~n49931 & n49932;
  assign n49934 = ~pi1154 & ~n49411;
  assign n49935 = ~n49933 & n49934;
  assign n49936 = pi1153 & n49285;
  assign n49937 = pi1154 & pi1155;
  assign n49938 = ~n49286 & n49937;
  assign n49939 = ~n49936 & n49938;
  assign n49940 = ~n49935 & ~n49939;
  assign n49941 = pi211 & ~n49940;
  assign n49942 = pi1154 & n49774;
  assign n49943 = pi1153 & n49287;
  assign n49944 = n49542 & ~n49772;
  assign n49945 = ~n49943 & n49944;
  assign n49946 = ~n49942 & n49945;
  assign n49947 = pi1154 & ~n49268;
  assign n49948 = pi1154 & n49421;
  assign n49949 = n49419 & n49947;
  assign n49950 = ~pi1155 & ~n65135;
  assign n49951 = ~pi1155 & ~n49933;
  assign n49952 = ~n65135 & n49951;
  assign n49953 = ~n49933 & n49950;
  assign n49954 = ~pi267 & ~n65136;
  assign n49955 = ~pi267 & ~n49946;
  assign n49956 = ~n65136 & n49955;
  assign n49957 = ~n49946 & n49954;
  assign n49958 = ~n49941 & n65137;
  assign n49959 = ~n49930 & ~n49958;
  assign n49960 = ~n49946 & ~n65136;
  assign n49961 = ~n49941 & n49960;
  assign n49962 = ~pi267 & ~n49961;
  assign n49963 = ~n49916 & ~n49928;
  assign n49964 = pi267 & ~n49963;
  assign n49965 = pi219 & ~n49964;
  assign n49966 = ~n49962 & n49965;
  assign n49967 = pi219 & ~n49959;
  assign n49968 = n49262 & ~n49910;
  assign n49969 = n49775 & ~n49968;
  assign n49970 = pi1154 & ~n49969;
  assign n49971 = ~pi1153 & ~n49311;
  assign n49972 = ~pi1154 & ~n49971;
  assign n49973 = pi1155 & ~n49972;
  assign n49974 = n49313 & ~n49973;
  assign n49975 = ~n49970 & ~n49974;
  assign n49976 = ~pi1155 & ~n49722;
  assign n49977 = ~n49722 & n49951;
  assign n49978 = ~n49933 & n49976;
  assign n49979 = pi211 & ~n65139;
  assign n49980 = ~n49975 & n49979;
  assign n49981 = ~n49312 & ~n49943;
  assign n49982 = pi1155 & ~n49981;
  assign n49983 = pi1153 & ~pi1155;
  assign n49984 = ~n49724 & ~n49983;
  assign n49985 = pi1153 & ~n49338;
  assign n49986 = ~pi1155 & n49985;
  assign n49987 = ~n49984 & ~n49986;
  assign n49988 = ~pi1155 & ~n49985;
  assign n49989 = ~pi1153 & ~n49724;
  assign n49990 = n49988 & ~n49989;
  assign n49991 = pi1154 & ~n49754;
  assign n49992 = ~n49990 & n49991;
  assign n49993 = pi1154 & ~n49987;
  assign n49994 = ~pi1153 & ~n49308;
  assign n49995 = ~n49275 & ~n49994;
  assign n49996 = ~pi1155 & n49995;
  assign n49997 = n49988 & n49995;
  assign n49998 = ~n49985 & n49996;
  assign n49999 = ~pi1154 & ~n65141;
  assign n50000 = ~n65140 & ~n49999;
  assign n50001 = ~n49982 & ~n50000;
  assign n50002 = ~n49982 & n49991;
  assign n50003 = ~n49990 & n50002;
  assign n50004 = ~n49982 & n65140;
  assign n50005 = ~pi1154 & ~n49982;
  assign n50006 = ~n65141 & n50005;
  assign n50007 = ~pi211 & ~n50006;
  assign n50008 = ~n65142 & n50007;
  assign n50009 = ~pi211 & ~n65142;
  assign n50010 = ~n50006 & n50009;
  assign n50011 = ~pi211 & ~n50001;
  assign n50012 = ~pi267 & ~n65143;
  assign n50013 = ~n49980 & n50012;
  assign n50014 = n49677 & n49925;
  assign n50015 = ~pi1153 & n49353;
  assign n50016 = ~n49311 & ~n50015;
  assign n50017 = ~pi1155 & n49262;
  assign n50018 = ~n50016 & n50017;
  assign n50019 = pi1154 & ~n50018;
  assign n50020 = pi1154 & ~n50014;
  assign n50021 = ~n50018 & n50020;
  assign n50022 = ~n50014 & n50019;
  assign n50023 = ~pi1154 & ~n49908;
  assign n50024 = ~n49274 & n50023;
  assign n50025 = ~pi1155 & ~n50024;
  assign n50026 = ~n49296 & n50023;
  assign n50027 = ~n50025 & n50026;
  assign n50028 = ~n65144 & ~n50027;
  assign n50029 = pi211 & ~n50028;
  assign n50030 = pi1154 & n50016;
  assign n50031 = n50025 & ~n50030;
  assign n50032 = ~pi1153 & n49305;
  assign n50033 = ~n49294 & ~n50032;
  assign n50034 = pi1154 & n49260;
  assign n50035 = pi1155 & ~n50034;
  assign n50036 = ~n50033 & n50035;
  assign n50037 = ~pi211 & ~n50036;
  assign n50038 = ~n50031 & n50037;
  assign n50039 = pi267 & ~n50038;
  assign n50040 = ~n50029 & n50039;
  assign n50041 = ~pi219 & ~n50040;
  assign n50042 = ~n50013 & n50041;
  assign n50043 = ~n65138 & ~n50042;
  assign n50044 = n49373 & ~n50043;
  assign n50045 = ~pi1153 & ~n49454;
  assign n50046 = pi1091 & n49794;
  assign n50047 = ~n50045 & n50046;
  assign n50048 = pi1154 & ~n50047;
  assign n50049 = pi1091 & ~pi1155;
  assign n50050 = ~pi200 & ~pi1153;
  assign n50051 = ~pi199 & ~n50050;
  assign n50052 = ~pi299 & n50051;
  assign n50053 = n50049 & n50052;
  assign n50054 = n50048 & ~n50053;
  assign n50055 = ~pi1153 & n39538;
  assign n50056 = n49595 & ~n50055;
  assign n50057 = pi1155 & n50056;
  assign n50058 = pi1154 & ~n50057;
  assign n50059 = n49794 & n50058;
  assign n50060 = ~n50054 & ~n50059;
  assign n50061 = pi211 & ~n50060;
  assign n50062 = ~pi211 & ~pi1154;
  assign n50063 = ~n50054 & ~n50062;
  assign n50064 = pi1153 & ~n49494;
  assign n50065 = ~pi1153 & ~n49519;
  assign n50066 = ~n50064 & ~n50065;
  assign n50067 = n49808 & ~n49831;
  assign n50068 = ~n50066 & n50067;
  assign n50069 = ~n50063 & ~n50068;
  assign n50070 = pi1154 & ~n50054;
  assign n50071 = ~pi211 & ~n50068;
  assign n50072 = ~n50070 & n50071;
  assign n50073 = ~n50061 & ~n50072;
  assign n50074 = ~n50061 & ~n50069;
  assign n50075 = pi219 & ~n65145;
  assign n50076 = ~pi1153 & ~n39539;
  assign n50077 = ~pi200 & pi1155;
  assign n50078 = n48570 & ~n50077;
  assign n50079 = ~pi1154 & n49494;
  assign n50080 = ~n50078 & ~n50079;
  assign n50081 = ~n50076 & n50080;
  assign n50082 = pi1091 & n50081;
  assign n50083 = ~pi211 & ~n50082;
  assign n50084 = pi211 & pi1154;
  assign n50085 = ~pi299 & ~n50051;
  assign n50086 = n50049 & ~n50085;
  assign n50087 = n50084 & ~n50086;
  assign n50088 = ~n50047 & n50087;
  assign n50089 = ~n50083 & ~n50088;
  assign n50090 = ~pi219 & ~n50089;
  assign n50091 = pi1153 & ~n39539;
  assign n50092 = ~pi1155 & ~n50091;
  assign n50093 = pi1091 & ~pi1153;
  assign n50094 = n49458 & n50093;
  assign n50095 = pi1091 & pi1153;
  assign n50096 = n49461 & n50095;
  assign n50097 = ~n50094 & ~n50096;
  assign n50098 = ~n50092 & ~n50097;
  assign n50099 = pi211 & ~pi1154;
  assign n50100 = ~n50098 & n50099;
  assign n50101 = ~n50090 & ~n50100;
  assign n50102 = ~n50075 & n50101;
  assign n50103 = ~pi267 & ~n50102;
  assign n50104 = pi1153 & ~n65111;
  assign n50105 = pi1155 & ~n50104;
  assign n50106 = n49796 & n50105;
  assign n50107 = ~pi1153 & ~n49502;
  assign n50108 = pi1153 & ~n49472;
  assign n50109 = ~pi1155 & ~n50108;
  assign n50110 = ~n50107 & n50109;
  assign n50111 = ~n50106 & ~n50110;
  assign n50112 = pi1154 & ~n50111;
  assign n50113 = n49458 & ~n49831;
  assign n50114 = n48570 & n50077;
  assign n50115 = n49808 & ~n65146;
  assign n50116 = ~pi1153 & ~n49459;
  assign n50117 = n50105 & ~n50116;
  assign n50118 = pi1091 & n50092;
  assign n50119 = ~n50117 & ~n50118;
  assign n50120 = ~pi1154 & ~n50119;
  assign n50121 = ~n50091 & n50115;
  assign n50122 = ~pi219 & ~n65147;
  assign n50123 = ~pi219 & ~n50112;
  assign n50124 = ~n65147 & n50123;
  assign n50125 = ~n50112 & n50122;
  assign n50126 = pi1091 & ~n50052;
  assign n50127 = n50048 & n50126;
  assign n50128 = pi1155 & ~n50066;
  assign n50129 = pi1153 & n48497;
  assign n50130 = ~pi1154 & ~n50129;
  assign n50131 = pi1091 & n50130;
  assign n50132 = n49808 & ~n50129;
  assign n50133 = ~n50128 & n65149;
  assign n50134 = pi219 & ~n50133;
  assign n50135 = ~n50127 & n50134;
  assign n50136 = ~n65148 & ~n50135;
  assign n50137 = ~pi211 & ~n50136;
  assign n50138 = ~pi1155 & ~n50085;
  assign n50139 = ~n49833 & ~n50138;
  assign n50140 = ~n48495 & ~n50139;
  assign n50141 = pi1091 & n50058;
  assign n50142 = ~n50140 & n50141;
  assign n50143 = ~n49459 & ~n49831;
  assign n50144 = n65149 & ~n50143;
  assign n50145 = ~n65146 & n65149;
  assign n50146 = pi211 & ~n65150;
  assign n50147 = ~n50142 & n50146;
  assign n50148 = pi267 & ~n50147;
  assign n50149 = ~n50137 & n50148;
  assign n50150 = ~n50137 & ~n50147;
  assign n50151 = pi267 & ~n50150;
  assign n50152 = ~pi219 & ~n50083;
  assign n50153 = ~pi219 & ~n50088;
  assign n50154 = ~n50083 & n50153;
  assign n50155 = ~n50088 & n50152;
  assign n50156 = pi219 & ~n50072;
  assign n50157 = pi219 & ~n50061;
  assign n50158 = ~n50072 & n50157;
  assign n50159 = ~n50061 & n50156;
  assign n50160 = ~n65151 & ~n65152;
  assign n50161 = ~pi267 & ~n50100;
  assign n50162 = ~n50160 & n50161;
  assign n50163 = ~n50151 & ~n50162;
  assign n50164 = ~n50103 & ~n50149;
  assign n50165 = ~n49373 & ~n65153;
  assign n50166 = n62455 & ~n50165;
  assign n50167 = ~n50044 & n50166;
  assign n50168 = ~pi219 & n49252;
  assign n50169 = ~n49875 & ~n50168;
  assign n50170 = pi267 & n50169;
  assign n50171 = ~pi267 & ~n49254;
  assign n50172 = ~n49886 & n50171;
  assign n50173 = n49373 & ~n50172;
  assign n50174 = ~n50170 & n50173;
  assign n50175 = pi219 & ~n49542;
  assign n50176 = ~pi211 & pi1153;
  assign n50177 = ~pi219 & ~n50084;
  assign n50178 = ~n50176 & n50177;
  assign n50179 = ~n50175 & ~n50178;
  assign n50180 = pi1091 & ~n50179;
  assign n50181 = ~pi267 & ~pi1091;
  assign n50182 = ~n49373 & n50181;
  assign n50183 = ~n50180 & ~n50182;
  assign n50184 = ~n50174 & n50183;
  assign n50185 = ~n62455 & ~n50184;
  assign n50186 = n49537 & ~n50185;
  assign n50187 = ~n50167 & n50186;
  assign n50188 = n62455 & n65153;
  assign n50189 = ~n50180 & ~n50181;
  assign n50190 = ~n62455 & ~n50189;
  assign n50191 = ~n49537 & ~n50190;
  assign n50192 = ~n50188 & n50191;
  assign n50193 = ~pi230 & ~n50192;
  assign n50194 = ~n50187 & n50193;
  assign n50195 = ~pi199 & ~pi1153;
  assign n50196 = n49461 & ~n50195;
  assign n50197 = pi1155 & n50196;
  assign n50198 = ~n50085 & ~n50130;
  assign n50199 = ~pi1155 & n50129;
  assign n50200 = ~pi1154 & ~n50199;
  assign n50201 = ~n50085 & ~n50200;
  assign n50202 = ~n50197 & ~n50201;
  assign n50203 = ~n50197 & ~n50198;
  assign n50204 = pi219 & ~n50056;
  assign n50205 = pi211 & ~n50204;
  assign n50206 = ~n65154 & n50205;
  assign n50207 = ~pi219 & ~n50081;
  assign n50208 = pi200 & ~n49611;
  assign n50209 = ~pi1155 & ~n48567;
  assign n50210 = ~n50055 & ~n50209;
  assign n50211 = ~n50208 & n50210;
  assign n50212 = pi219 & ~n49607;
  assign n50213 = ~n50211 & n50212;
  assign n50214 = ~pi211 & ~n50213;
  assign n50215 = ~n50207 & n50214;
  assign n50216 = ~n50206 & ~n50215;
  assign n50217 = ~n65154 & ~n50204;
  assign n50218 = pi211 & ~n50217;
  assign n50219 = ~n49607 & ~n50211;
  assign n50220 = pi219 & ~n50219;
  assign n50221 = ~pi219 & n50081;
  assign n50222 = ~pi211 & ~n50221;
  assign n50223 = ~n50220 & n50222;
  assign n50224 = n62455 & ~n50223;
  assign n50225 = ~n50218 & n50224;
  assign n50226 = n62455 & ~n50216;
  assign n50227 = ~n62455 & n50179;
  assign n50228 = pi230 & ~n50227;
  assign n50229 = ~n65155 & n50228;
  assign po424 = ~n50194 & ~n50229;
  assign n50231 = pi1153 & ~pi1154;
  assign n50232 = ~n49800 & n50231;
  assign n50233 = ~pi1153 & ~n49461;
  assign n50234 = ~n49832 & ~n50233;
  assign n50235 = pi1154 & n50234;
  assign n50236 = ~n50232 & ~n50235;
  assign n50237 = n48476 & ~n50236;
  assign n50238 = ~pi199 & pi1153;
  assign n50239 = pi200 & n50238;
  assign n50240 = pi1153 & n48474;
  assign n50241 = ~pi299 & n65156;
  assign n50242 = ~pi1154 & ~n50241;
  assign n50243 = pi299 & n39423;
  assign n50244 = n49599 & ~n50195;
  assign n50245 = ~n48476 & n50244;
  assign n50246 = ~n50243 & ~n50245;
  assign n50247 = ~n50242 & ~n50246;
  assign n50248 = ~n50237 & ~n50247;
  assign n50249 = n62455 & ~n50248;
  assign n50250 = pi219 & ~n49653;
  assign n50251 = pi211 & pi1153;
  assign n50252 = ~pi219 & ~n50251;
  assign n50253 = ~n50250 & ~n50252;
  assign n50254 = ~n62455 & n50253;
  assign n50255 = ~pi1152 & ~n50254;
  assign n50256 = ~n50249 & n50255;
  assign n50257 = ~n48498 & ~n49461;
  assign n50258 = pi1154 & ~n50257;
  assign n50259 = pi200 & ~pi1153;
  assign n50260 = n48567 & ~n50259;
  assign n50261 = pi219 & ~n50260;
  assign n50262 = pi1153 & ~n49595;
  assign n50263 = ~n50233 & ~n50262;
  assign n50264 = n50084 & ~n50263;
  assign n50265 = pi1154 & n49494;
  assign n50266 = ~n50238 & n50265;
  assign n50267 = ~pi1154 & ~n50260;
  assign n50268 = ~n50266 & ~n50267;
  assign n50269 = ~n50264 & n50268;
  assign n50270 = pi219 & ~n50269;
  assign n50271 = ~n50258 & n50261;
  assign n50272 = ~pi200 & pi1154;
  assign n50273 = n48570 & ~n50272;
  assign n50274 = ~n48498 & n50233;
  assign n50275 = ~n50273 & ~n50274;
  assign n50276 = ~pi219 & ~n50275;
  assign n50277 = n62455 & ~n50276;
  assign n50278 = ~n65157 & n50277;
  assign n50279 = ~n62455 & ~n50250;
  assign n50280 = n48476 & ~n50251;
  assign n50281 = n50279 & ~n50280;
  assign n50282 = pi1152 & ~n50281;
  assign n50283 = ~n50278 & n50282;
  assign n50284 = ~n50256 & ~n50283;
  assign n50285 = pi230 & ~n50284;
  assign n50286 = ~n49265 & ~n49269;
  assign n50287 = ~pi1153 & ~n50286;
  assign n50288 = ~n49276 & n49920;
  assign n50289 = ~n50287 & n50288;
  assign n50290 = ~pi1153 & n50289;
  assign n50291 = ~n49311 & ~n50290;
  assign n50292 = ~pi1154 & ~n50291;
  assign n50293 = pi1153 & ~n65102;
  assign n50294 = n49920 & n49947;
  assign n50295 = ~n50293 & n50294;
  assign n50296 = pi254 & ~n50295;
  assign n50297 = ~n50292 & n50296;
  assign n50298 = ~n49338 & ~n49942;
  assign n50299 = pi211 & n49261;
  assign n50300 = ~n49275 & ~n50299;
  assign n50301 = ~pi1153 & ~n50300;
  assign n50302 = ~pi254 & ~n50301;
  assign n50303 = ~n50298 & n50302;
  assign n50304 = ~n50297 & ~n50303;
  assign n50305 = ~pi219 & ~n50304;
  assign n50306 = ~n49378 & ~n49922;
  assign n50307 = pi1153 & ~n49922;
  assign n50308 = pi1154 & ~n50307;
  assign n50309 = ~n50306 & n50308;
  assign n50310 = pi1153 & ~n49424;
  assign n50311 = ~pi1153 & ~n49430;
  assign n50312 = ~pi1154 & ~n50311;
  assign n50313 = ~n50310 & n50312;
  assign n50314 = pi254 & ~n50313;
  assign n50315 = ~n50309 & n50314;
  assign n50316 = n49421 & ~n49931;
  assign n50317 = ~pi1154 & ~n50316;
  assign n50318 = ~n49932 & n50317;
  assign n50319 = ~pi1153 & ~n49424;
  assign n50320 = n49774 & ~n50319;
  assign n50321 = n49653 & ~n50320;
  assign n50322 = ~n49244 & n50321;
  assign n50323 = ~n49407 & n50084;
  assign n50324 = ~n49936 & n50323;
  assign n50325 = ~pi254 & ~n50324;
  assign n50326 = ~n50322 & n50325;
  assign n50327 = ~n50318 & n50325;
  assign n50328 = ~n50322 & n50327;
  assign n50329 = ~n50318 & n50326;
  assign n50330 = ~n50315 & ~n65158;
  assign n50331 = pi219 & ~n50330;
  assign n50332 = pi253 & ~n50331;
  assign n50333 = ~n50305 & n50332;
  assign n50334 = pi219 & pi1091;
  assign n50335 = ~n49879 & ~n50334;
  assign n50336 = ~n50269 & ~n50335;
  assign n50337 = ~pi211 & n50076;
  assign n50338 = ~pi1154 & ~n50108;
  assign n50339 = ~n50045 & n50338;
  assign n50340 = ~n50045 & ~n50337;
  assign n50341 = n50338 & n50340;
  assign n50342 = ~n50337 & n50339;
  assign n50343 = pi1153 & ~n48570;
  assign n50344 = pi1091 & n50084;
  assign n50345 = ~n49461 & n50344;
  assign n50346 = ~n50343 & n50345;
  assign n50347 = ~n65159 & ~n50346;
  assign n50348 = ~pi219 & ~n50347;
  assign n50349 = ~n50336 & ~n50348;
  assign n50350 = pi254 & ~n50349;
  assign n50351 = ~pi254 & ~pi1091;
  assign n50352 = ~n65157 & ~n50276;
  assign n50353 = ~pi254 & ~n50352;
  assign n50354 = ~n50351 & ~n50353;
  assign n50355 = ~n50350 & n50354;
  assign n50356 = ~pi253 & ~n50355;
  assign n50357 = n62455 & ~n50356;
  assign n50358 = ~n50333 & n50357;
  assign n50359 = n49878 & ~n49883;
  assign n50360 = ~n50095 & n50359;
  assign n50361 = pi1091 & n50250;
  assign n50362 = ~pi254 & ~n50361;
  assign n50363 = ~n49886 & n50362;
  assign n50364 = ~n50360 & n50363;
  assign n50365 = n48476 & n50093;
  assign n50366 = pi254 & ~n50365;
  assign n50367 = ~n50361 & n50366;
  assign n50368 = n50169 & n50367;
  assign n50369 = pi253 & ~n50368;
  assign n50370 = pi253 & ~n50364;
  assign n50371 = ~n50368 & n50370;
  assign n50372 = ~n50364 & n50369;
  assign n50373 = pi1091 & ~n50253;
  assign n50374 = ~n62455 & ~n50351;
  assign n50375 = ~n50373 & n50374;
  assign n50376 = ~pi219 & n49812;
  assign n50377 = ~pi219 & ~n49254;
  assign n50378 = ~n49917 & n50377;
  assign n50379 = ~pi219 & ~n50378;
  assign n50380 = ~n62455 & n50379;
  assign n50381 = ~n49243 & n50380;
  assign n50382 = ~n62455 & n50376;
  assign n50383 = ~n50375 & ~n65161;
  assign n50384 = pi253 & ~n62455;
  assign n50385 = n50383 & ~n50384;
  assign n50386 = ~n65160 & ~n50385;
  assign n50387 = pi1152 & ~n50386;
  assign n50388 = ~n50358 & n50387;
  assign n50389 = ~pi211 & n49772;
  assign n50390 = ~n49262 & ~n50389;
  assign n50391 = ~n50032 & n50390;
  assign n50392 = ~pi219 & ~n49746;
  assign n50393 = ~n50391 & n50392;
  assign n50394 = ~pi1154 & ~n49934;
  assign n50395 = ~pi1154 & n49411;
  assign n50396 = ~n49921 & ~n50032;
  assign n50397 = ~n65162 & n50396;
  assign n50398 = ~n49389 & n49653;
  assign n50399 = pi219 & ~n50398;
  assign n50400 = ~n50397 & n50399;
  assign n50401 = ~n50393 & ~n50400;
  assign n50402 = pi254 & ~n50401;
  assign n50403 = n49286 & ~n50319;
  assign n50404 = n50084 & ~n50403;
  assign n50405 = pi219 & ~n50321;
  assign n50406 = pi219 & ~n50317;
  assign n50407 = ~n50321 & n50406;
  assign n50408 = ~n50317 & n50405;
  assign n50409 = ~n50404 & n65163;
  assign n50410 = n49722 & ~n49994;
  assign n50411 = pi1154 & n49312;
  assign n50412 = ~n50410 & ~n50411;
  assign n50413 = ~n49261 & ~n49766;
  assign n50414 = ~pi211 & ~n50413;
  assign n50415 = ~pi219 & ~n50414;
  assign n50416 = pi1154 & ~n49312;
  assign n50417 = ~n50410 & n50416;
  assign n50418 = ~pi1154 & ~n50410;
  assign n50419 = n50415 & ~n50418;
  assign n50420 = ~n50417 & n50419;
  assign n50421 = n50415 & ~n50417;
  assign n50422 = ~n50418 & n50421;
  assign n50423 = ~n50412 & n50415;
  assign n50424 = ~pi254 & ~n65164;
  assign n50425 = ~n50409 & n50424;
  assign n50426 = ~n50402 & ~n50425;
  assign n50427 = pi253 & ~n50426;
  assign n50428 = pi1153 & ~n49832;
  assign n50429 = pi1091 & n50428;
  assign n50430 = ~n50094 & ~n50429;
  assign n50431 = pi211 & ~n50338;
  assign n50432 = ~n50430 & n50431;
  assign n50433 = pi1091 & n50244;
  assign n50434 = pi1154 & ~n50433;
  assign n50435 = n48475 & n50095;
  assign n50436 = ~pi1154 & ~n50435;
  assign n50437 = ~pi211 & ~n50436;
  assign n50438 = ~n50434 & n50437;
  assign n50439 = ~n50432 & ~n50438;
  assign n50440 = ~pi219 & ~n50439;
  assign n50441 = pi211 & n50434;
  assign n50442 = pi1091 & n50065;
  assign n50443 = n49653 & ~n50442;
  assign n50444 = ~n50429 & n50443;
  assign n50445 = pi219 & ~n50436;
  assign n50446 = ~n50444 & n50445;
  assign n50447 = ~n50441 & n50446;
  assign n50448 = ~n50440 & ~n50447;
  assign n50449 = ~pi254 & ~n50448;
  assign n50450 = pi1091 & ~n48476;
  assign n50451 = ~n50241 & n50450;
  assign n50452 = ~pi1154 & ~n50451;
  assign n50453 = ~n39423 & ~n48476;
  assign n50454 = n49448 & ~n49598;
  assign n50455 = pi1153 & ~n50454;
  assign n50456 = ~n50116 & ~n50455;
  assign n50457 = ~n49796 & ~n50456;
  assign n50458 = n50453 & ~n50457;
  assign n50459 = n39423 & ~n50455;
  assign n50460 = n49520 & n50459;
  assign n50461 = pi1154 & ~n50460;
  assign n50462 = ~n50458 & n50461;
  assign n50463 = ~n50452 & ~n50462;
  assign n50464 = n49800 & n49808;
  assign n50465 = ~pi1154 & n49476;
  assign n50466 = ~n50456 & ~n65165;
  assign n50467 = n48476 & ~n50466;
  assign n50468 = pi254 & ~n50467;
  assign n50469 = ~n50463 & n50468;
  assign n50470 = ~n50449 & ~n50469;
  assign n50471 = ~pi253 & n50470;
  assign n50472 = n62455 & ~n50471;
  assign n50473 = ~n50427 & n50472;
  assign n50474 = ~n50375 & ~n50384;
  assign n50475 = n50364 & ~n50379;
  assign n50476 = ~n50359 & n50377;
  assign n50477 = n50368 & ~n50476;
  assign n50478 = pi253 & ~n50477;
  assign n50479 = pi253 & ~n50475;
  assign n50480 = ~n50477 & n50479;
  assign n50481 = ~n50475 & n50478;
  assign n50482 = ~n50474 & ~n65166;
  assign n50483 = ~pi1152 & ~n50482;
  assign n50484 = ~n50473 & n50483;
  assign n50485 = n49537 & ~n50484;
  assign n50486 = ~n50388 & n50485;
  assign n50487 = n62455 & ~n50470;
  assign n50488 = ~pi1152 & ~n50375;
  assign n50489 = ~n50487 & n50488;
  assign n50490 = n62455 & n50355;
  assign n50491 = pi1152 & n50383;
  assign n50492 = ~n50490 & n50491;
  assign n50493 = ~n49537 & ~n50492;
  assign n50494 = ~n50489 & n50493;
  assign n50495 = ~pi230 & ~n50494;
  assign n50496 = ~n50486 & n50495;
  assign po411 = ~n50285 & ~n50496;
  assign n50498 = ~pi230 & pi587;
  assign n50499 = pi230 & n7187;
  assign n50500 = ~n63011 & n50499;
  assign n50501 = ~n27509 & n50500;
  assign n50502 = n63013 & n50501;
  assign n50503 = n11558 & n50502;
  assign n50504 = n13393 & n50501;
  assign n50505 = ~n50498 & ~n65167;
  assign n50506 = ~pi230 & pi602;
  assign n50507 = pi230 & n7563;
  assign n50508 = ~n62892 & n50507;
  assign n50509 = pi790 & ~n11539;
  assign n50510 = pi790 & ~n11541;
  assign n50511 = ~n11539 & n50510;
  assign n50512 = ~n11541 & n50509;
  assign n50513 = ~n62964 & ~n10298;
  assign n50514 = ~n65168 & n50513;
  assign n50515 = n50508 & n50514;
  assign n50516 = n10206 & n50508;
  assign n50517 = n10106 & n50508;
  assign n50518 = n10206 & n50517;
  assign n50519 = n10106 & n50516;
  assign n50520 = n50514 & n65169;
  assign n50521 = n10207 & n50515;
  assign n50522 = ~n50506 & ~n65170;
  assign n50523 = ~pi219 & pi299;
  assign n50524 = ~n48494 & ~n50523;
  assign n50525 = ~n49519 & n50524;
  assign n50526 = n62455 & n50525;
  assign n50527 = pi219 & n48935;
  assign n50528 = ~n50526 & ~n50527;
  assign n50529 = ~pi1151 & pi1153;
  assign n50530 = ~n50528 & n50529;
  assign n50531 = ~n50064 & ~n50076;
  assign n50532 = n39421 & n50531;
  assign n50533 = pi199 & ~pi1153;
  assign n50534 = n49461 & ~n50533;
  assign n50535 = pi211 & ~n50534;
  assign n50536 = ~n50532 & ~n50535;
  assign n50537 = pi1151 & n62455;
  assign n50538 = ~pi1153 & ~n48567;
  assign n50539 = ~n49494 & ~n50538;
  assign n50540 = n39423 & ~n50539;
  assign n50541 = n50537 & ~n50540;
  assign n50542 = n50536 & n50541;
  assign n50543 = ~n50530 & ~n50542;
  assign n50544 = ~pi1152 & ~n50543;
  assign n50545 = n39423 & n50428;
  assign n50546 = n49599 & ~n50533;
  assign n50547 = ~pi1151 & ~n48477;
  assign n50548 = ~n50546 & n50547;
  assign n50549 = ~n50545 & n50548;
  assign n50550 = pi1152 & n62455;
  assign n50551 = pi1153 & ~n50257;
  assign n50552 = ~n48567 & ~n50523;
  assign n50553 = pi1151 & n50552;
  assign n50554 = ~n50551 & n50553;
  assign n50555 = n50550 & ~n50554;
  assign n50556 = ~n50549 & n50555;
  assign n50557 = pi219 & ~n50176;
  assign n50558 = ~pi219 & ~n62455;
  assign n50559 = pi1153 & n48935;
  assign n50560 = ~n62455 & n50176;
  assign n50561 = ~n50558 & ~n65171;
  assign n50562 = ~n62455 & ~n50557;
  assign n50563 = pi1152 & ~n39421;
  assign n50564 = pi1151 & ~n48476;
  assign n50565 = ~n50563 & ~n50564;
  assign n50566 = ~n65172 & ~n50565;
  assign n50567 = pi230 & ~n50566;
  assign n50568 = pi230 & ~n50556;
  assign n50569 = ~n50566 & n50568;
  assign n50570 = ~n50556 & n50567;
  assign n50571 = pi1153 & ~n50528;
  assign n50572 = ~pi1151 & ~n50571;
  assign n50573 = n62455 & ~n50540;
  assign n50574 = n50536 & n50573;
  assign n50575 = ~n48476 & ~n65172;
  assign n50576 = pi1151 & ~n50575;
  assign n50577 = pi1151 & ~n50574;
  assign n50578 = ~n50575 & n50577;
  assign n50579 = ~n50574 & n50576;
  assign n50580 = ~n50572 & ~n65174;
  assign n50581 = ~pi1152 & ~n50580;
  assign n50582 = n62455 & ~n50554;
  assign n50583 = ~n50549 & n50582;
  assign n50584 = ~pi1151 & n39421;
  assign n50585 = ~n50557 & ~n50584;
  assign n50586 = ~n65172 & ~n50584;
  assign n50587 = ~n62455 & n50585;
  assign n50588 = pi1152 & ~n65175;
  assign n50589 = pi1152 & ~n50583;
  assign n50590 = ~n65175 & n50589;
  assign n50591 = ~n50583 & n50588;
  assign n50592 = ~n50581 & ~n65176;
  assign n50593 = pi230 & ~n50592;
  assign n50594 = ~n50544 & n65173;
  assign n50595 = pi219 & ~n50319;
  assign n50596 = ~n50307 & n50595;
  assign n50597 = ~pi219 & ~n49971;
  assign n50598 = ~n50293 & n50597;
  assign n50599 = pi253 & ~n50598;
  assign n50600 = pi253 & ~n50596;
  assign n50601 = ~n50598 & n50600;
  assign n50602 = ~n50596 & n50599;
  assign n50603 = ~n49285 & ~n50389;
  assign n50604 = pi1153 & ~n50603;
  assign n50605 = ~n49419 & ~n50604;
  assign n50606 = pi219 & n50605;
  assign n50607 = pi1153 & n49291;
  assign n50608 = ~pi219 & ~n49908;
  assign n50609 = ~n50607 & n50608;
  assign n50610 = ~pi253 & ~n50609;
  assign n50611 = ~n50606 & n50610;
  assign n50612 = ~n65178 & ~n50611;
  assign n50613 = n62455 & ~n50612;
  assign n50614 = pi253 & ~n49283;
  assign n50615 = ~n50377 & n50614;
  assign n50616 = ~pi253 & ~n49878;
  assign n50617 = ~n49886 & n50616;
  assign n50618 = ~n50615 & ~n50617;
  assign n50619 = ~n50176 & n50334;
  assign n50620 = ~n62455 & ~n50619;
  assign n50621 = ~n49878 & ~n50619;
  assign n50622 = ~n49886 & n50621;
  assign n50623 = ~pi253 & ~n50622;
  assign n50624 = ~n49283 & ~n50619;
  assign n50625 = ~n50377 & n50624;
  assign n50626 = pi253 & ~n50625;
  assign n50627 = ~n62455 & ~n50626;
  assign n50628 = ~n50623 & n50627;
  assign n50629 = ~n62455 & ~n50623;
  assign n50630 = ~n50626 & n50629;
  assign n50631 = ~n50618 & n50620;
  assign n50632 = pi1151 & ~n65161;
  assign n50633 = pi1151 & ~n65179;
  assign n50634 = ~n65161 & n50633;
  assign n50635 = ~n65179 & n50632;
  assign n50636 = ~n50613 & n65180;
  assign n50637 = ~pi219 & ~n50289;
  assign n50638 = pi219 & n49273;
  assign n50639 = ~n50637 & ~n50638;
  assign n50640 = ~n50606 & n50639;
  assign n50641 = ~pi253 & ~n50640;
  assign n50642 = n50377 & ~n50390;
  assign n50643 = ~n49270 & ~n50287;
  assign n50644 = n50642 & ~n50643;
  assign n50645 = pi219 & n49376;
  assign n50646 = ~n49389 & n50307;
  assign n50647 = n50645 & ~n50646;
  assign n50648 = ~n50644 & ~n50647;
  assign n50649 = pi253 & ~n50648;
  assign n50650 = n62455 & ~n50649;
  assign n50651 = ~n50641 & n50650;
  assign n50652 = ~pi1151 & ~n50651;
  assign n50653 = ~n50636 & ~n50652;
  assign n50654 = ~n62455 & ~n49873;
  assign n50655 = ~n50476 & n50654;
  assign n50656 = ~n49243 & n50655;
  assign n50657 = ~n65179 & ~n50656;
  assign n50658 = ~n50653 & n50657;
  assign n50659 = pi1152 & ~n50658;
  assign n50660 = pi219 & ~n50605;
  assign n50661 = ~n50609 & n50642;
  assign n50662 = ~n50660 & ~n50661;
  assign n50663 = ~n49275 & ~n50662;
  assign n50664 = ~pi253 & ~n50663;
  assign n50665 = n49920 & n50377;
  assign n50666 = ~n49924 & n50665;
  assign n50667 = pi1153 & n50306;
  assign n50668 = pi219 & ~n50311;
  assign n50669 = ~n50667 & n50668;
  assign n50670 = ~n50666 & ~n50669;
  assign n50671 = pi253 & ~n50670;
  assign n50672 = n62455 & ~n50671;
  assign n50673 = ~n50664 & n50672;
  assign n50674 = n65180 & ~n50673;
  assign n50675 = ~n49259 & n50660;
  assign n50676 = ~pi219 & n49311;
  assign n50677 = n49995 & n50676;
  assign n50678 = ~pi253 & ~n50677;
  assign n50679 = ~n50675 & n50678;
  assign n50680 = ~pi219 & n50286;
  assign n50681 = ~n49912 & ~n50680;
  assign n50682 = n49923 & n50681;
  assign n50683 = pi253 & ~n50682;
  assign n50684 = n62455 & ~n50683;
  assign n50685 = ~n50679 & n50684;
  assign n50686 = ~pi1151 & ~n65179;
  assign n50687 = ~n50685 & n50686;
  assign n50688 = ~pi1152 & ~n50687;
  assign n50689 = ~n50674 & n50688;
  assign n50690 = ~n50659 & ~n50689;
  assign n50691 = n49537 & ~n50690;
  assign n50692 = pi1091 & ~n50536;
  assign n50693 = n39423 & ~n50104;
  assign n50694 = ~n50045 & n50693;
  assign n50695 = ~n50692 & ~n50694;
  assign n50696 = pi253 & ~n50695;
  assign n50697 = n65044 & ~n50551;
  assign n50698 = pi1091 & ~n50697;
  assign n50699 = ~pi253 & ~n50698;
  assign n50700 = n62455 & ~n50699;
  assign n50701 = ~n50696 & n50700;
  assign n50702 = ~pi253 & ~pi1091;
  assign n50703 = ~n62455 & ~n50702;
  assign n50704 = pi219 & n50093;
  assign n50705 = ~n49802 & ~n50704;
  assign n50706 = n50703 & n50705;
  assign n50707 = pi1151 & ~n50706;
  assign n50708 = ~n50701 & n50707;
  assign n50709 = ~n50619 & n50703;
  assign n50710 = pi219 & n50709;
  assign n50711 = n50095 & n50526;
  assign n50712 = pi253 & ~pi1091;
  assign n50713 = ~pi1151 & ~n50712;
  assign n50714 = ~n50711 & n50713;
  assign n50715 = ~n50710 & n50714;
  assign n50716 = ~n50708 & ~n50715;
  assign n50717 = ~pi1152 & ~n50716;
  assign n50718 = pi1091 & n50546;
  assign n50719 = pi211 & ~n49516;
  assign n50720 = ~n50718 & n50719;
  assign n50721 = n65111 & n50195;
  assign n50722 = n39423 & ~n50721;
  assign n50723 = ~n50429 & n50722;
  assign n50724 = ~pi253 & ~n50723;
  assign n50725 = ~pi253 & ~n50720;
  assign n50726 = ~n50723 & n50725;
  assign n50727 = ~n50720 & n50724;
  assign n50728 = ~n50107 & n50459;
  assign n50729 = n48476 & n49448;
  assign n50730 = ~n50546 & n50729;
  assign n50731 = pi253 & ~n50730;
  assign n50732 = ~n50728 & n50731;
  assign n50733 = ~n65181 & ~n50732;
  assign n50734 = ~pi57 & ~pi1151;
  assign n50735 = ~pi1151 & n62455;
  assign n50736 = n3475 & n50734;
  assign n50737 = n50453 & ~n50712;
  assign n50738 = ~n50718 & n50737;
  assign n50739 = n65182 & ~n50738;
  assign n50740 = ~n50733 & n50739;
  assign n50741 = ~pi1151 & n50376;
  assign n50742 = n50709 & ~n50741;
  assign n50743 = n50257 & ~n50712;
  assign n50744 = ~n50093 & ~n50743;
  assign n50745 = n50552 & ~n50744;
  assign n50746 = n50537 & ~n50702;
  assign n50747 = ~n50745 & n50746;
  assign n50748 = pi1152 & ~n50747;
  assign n50749 = n62455 & ~n50702;
  assign n50750 = ~n50745 & n50749;
  assign n50751 = ~n50709 & ~n50750;
  assign n50752 = pi1151 & ~n50751;
  assign n50753 = ~n50376 & n50709;
  assign n50754 = pi1152 & ~n50753;
  assign n50755 = ~n50752 & n50754;
  assign n50756 = ~n50742 & n50748;
  assign n50757 = ~n50740 & n65183;
  assign n50758 = ~n49537 & ~n50757;
  assign n50759 = ~n50717 & n50758;
  assign n50760 = ~pi230 & ~n50759;
  assign n50761 = ~n50691 & n50760;
  assign po410 = ~n65177 & ~n50761;
  assign n50763 = ~pi1137 & ~pi1138;
  assign n50764 = ~pi1134 & n50763;
  assign n50765 = ~pi680 & pi1135;
  assign n50766 = ~pi603 & ~pi1135;
  assign n50767 = pi1136 & ~n50766;
  assign n50768 = pi1136 & ~n50765;
  assign n50769 = ~n50766 & n50768;
  assign n50770 = ~n50765 & n50767;
  assign n50771 = ~pi778 & pi1135;
  assign n50772 = ~pi981 & ~pi1135;
  assign n50773 = ~pi1136 & ~n50772;
  assign n50774 = ~pi1136 & ~n50771;
  assign n50775 = ~n50772 & n50774;
  assign n50776 = ~n50771 & n50773;
  assign n50777 = ~n65184 & ~n65185;
  assign n50778 = n50764 & ~n50777;
  assign n50779 = pi1135 & n50763;
  assign n50780 = pi1136 & ~n50779;
  assign n50781 = ~pi759 & n50780;
  assign n50782 = pi1135 & ~pi1136;
  assign n50783 = pi1134 & n50763;
  assign n50784 = ~n50782 & n50783;
  assign n50785 = ~pi696 & pi1135;
  assign n50786 = ~pi837 & ~pi1136;
  assign n50787 = ~n50785 & ~n50786;
  assign n50788 = n50784 & n50787;
  assign n50789 = ~n50781 & n50788;
  assign n50790 = ~n50778 & ~n50789;
  assign n50791 = ~n5530 & ~n50790;
  assign n50792 = ~pi590 & pi592;
  assign n50793 = ~pi588 & ~n50792;
  assign n50794 = ~pi590 & pi591;
  assign n50795 = pi390 & n50794;
  assign n50796 = n50793 & ~n50795;
  assign n50797 = pi363 & ~pi591;
  assign n50798 = pi592 & ~n50797;
  assign n50799 = ~n50796 & ~n50798;
  assign n50800 = pi590 & ~pi591;
  assign n50801 = ~pi592 & n50800;
  assign n50802 = pi342 & n50801;
  assign n50803 = ~n50799 & ~n50802;
  assign n50804 = ~pi223 & ~pi224;
  assign n50805 = pi414 & n5481;
  assign n50806 = pi588 & ~n50805;
  assign n50807 = n50804 & ~n50806;
  assign n50808 = ~n50803 & n50807;
  assign n50809 = pi199 & ~pi1049;
  assign n50810 = ~pi199 & ~pi291;
  assign n50811 = ~n50804 & ~n50810;
  assign n50812 = ~n50804 & ~n50809;
  assign n50813 = ~n50810 & n50812;
  assign n50814 = ~n50809 & n50811;
  assign n50815 = ~n50808 & ~n65186;
  assign n50816 = n5530 & ~n50815;
  assign n50817 = ~n50791 & ~n50816;
  assign n50818 = ~pi661 & pi1135;
  assign n50819 = ~pi616 & ~pi1135;
  assign n50820 = pi1136 & ~n50819;
  assign n50821 = pi1136 & ~n50818;
  assign n50822 = ~n50819 & n50821;
  assign n50823 = ~n50818 & n50820;
  assign n50824 = ~pi781 & pi1135;
  assign n50825 = ~pi808 & ~pi1135;
  assign n50826 = ~pi1136 & ~n50825;
  assign n50827 = ~pi1136 & ~n50824;
  assign n50828 = ~n50825 & n50827;
  assign n50829 = ~n50824 & n50826;
  assign n50830 = ~n65187 & ~n65188;
  assign n50831 = n50764 & ~n50830;
  assign n50832 = ~pi758 & n50780;
  assign n50833 = ~pi736 & pi1135;
  assign n50834 = ~pi850 & ~pi1136;
  assign n50835 = ~n50833 & ~n50834;
  assign n50836 = n50784 & n50835;
  assign n50837 = ~n50832 & n50836;
  assign n50838 = ~n50831 & ~n50837;
  assign n50839 = ~n5530 & ~n50838;
  assign n50840 = pi397 & n50794;
  assign n50841 = n50793 & ~n50840;
  assign n50842 = pi372 & ~pi591;
  assign n50843 = pi592 & ~n50842;
  assign n50844 = ~n50841 & ~n50843;
  assign n50845 = pi320 & n50801;
  assign n50846 = ~n50844 & ~n50845;
  assign n50847 = pi422 & n5481;
  assign n50848 = pi588 & ~n50847;
  assign n50849 = n50804 & ~n50848;
  assign n50850 = ~n50846 & n50849;
  assign n50851 = pi199 & ~pi1048;
  assign n50852 = ~pi199 & ~pi290;
  assign n50853 = ~n50804 & ~n50852;
  assign n50854 = ~n50804 & ~n50851;
  assign n50855 = ~n50852 & n50854;
  assign n50856 = ~n50851 & n50853;
  assign n50857 = ~n50850 & ~n65189;
  assign n50858 = n5530 & ~n50857;
  assign n50859 = ~n50839 & ~n50858;
  assign n50860 = ~pi637 & pi1135;
  assign n50861 = ~pi617 & ~pi1135;
  assign n50862 = pi1136 & ~n50861;
  assign n50863 = pi1136 & ~n50860;
  assign n50864 = ~n50861 & n50863;
  assign n50865 = ~n50860 & n50862;
  assign n50866 = pi814 & ~pi1135;
  assign n50867 = ~pi788 & pi1135;
  assign n50868 = ~pi1136 & ~n50867;
  assign n50869 = ~pi1136 & ~n50866;
  assign n50870 = ~n50867 & n50869;
  assign n50871 = ~n50866 & n50868;
  assign n50872 = ~n65190 & ~n65191;
  assign n50873 = n50764 & ~n50872;
  assign n50874 = ~pi749 & n50780;
  assign n50875 = ~pi706 & pi1135;
  assign n50876 = ~pi866 & ~pi1136;
  assign n50877 = ~n50875 & ~n50876;
  assign n50878 = n50784 & n50877;
  assign n50879 = ~n50874 & n50878;
  assign n50880 = ~n50873 & ~n50879;
  assign n50881 = ~n5530 & ~n50880;
  assign n50882 = pi411 & n50794;
  assign n50883 = n50793 & ~n50882;
  assign n50884 = pi387 & ~pi591;
  assign n50885 = pi592 & ~n50884;
  assign n50886 = ~n50883 & ~n50885;
  assign n50887 = pi452 & n50801;
  assign n50888 = ~n50886 & ~n50887;
  assign n50889 = pi435 & n5481;
  assign n50890 = pi588 & ~n50889;
  assign n50891 = n50804 & ~n50890;
  assign n50892 = ~n50888 & n50891;
  assign n50893 = pi199 & ~pi1053;
  assign n50894 = ~pi199 & ~pi295;
  assign n50895 = ~n50804 & ~n50894;
  assign n50896 = ~n50804 & ~n50893;
  assign n50897 = ~n50894 & n50896;
  assign n50898 = ~n50893 & n50895;
  assign n50899 = ~n50892 & ~n65192;
  assign n50900 = n5530 & ~n50899;
  assign n50901 = ~n50881 & ~n50900;
  assign n50902 = pi199 & ~pi1070;
  assign n50903 = ~pi199 & ~pi256;
  assign n50904 = ~n50804 & ~n50903;
  assign n50905 = ~n50804 & ~n50902;
  assign n50906 = ~n50903 & n50905;
  assign n50907 = ~n50902 & n50904;
  assign n50908 = ~pi591 & pi592;
  assign n50909 = pi336 & n50908;
  assign n50910 = pi463 & pi591;
  assign n50911 = ~pi592 & n50910;
  assign n50912 = ~n50909 & ~n50911;
  assign n50913 = ~pi590 & ~n50912;
  assign n50914 = pi362 & n50801;
  assign n50915 = ~pi588 & ~n50914;
  assign n50916 = ~n50913 & n50915;
  assign n50917 = pi437 & n5481;
  assign n50918 = pi588 & ~n50917;
  assign n50919 = n50804 & ~n50918;
  assign n50920 = ~n50916 & n50919;
  assign n50921 = ~n65193 & ~n50920;
  assign n50922 = n5530 & ~n50921;
  assign n50923 = pi639 & pi1135;
  assign n50924 = pi622 & ~pi1135;
  assign n50925 = pi1136 & ~n50924;
  assign n50926 = pi1136 & ~n50923;
  assign n50927 = ~n50924 & n50926;
  assign n50928 = ~n50923 & n50925;
  assign n50929 = pi783 & pi1135;
  assign n50930 = pi804 & ~pi1135;
  assign n50931 = ~pi1136 & ~n50930;
  assign n50932 = ~pi1136 & ~n50929;
  assign n50933 = ~n50930 & n50932;
  assign n50934 = ~n50929 & n50931;
  assign n50935 = ~n65194 & ~n65195;
  assign n50936 = ~pi1134 & ~n50935;
  assign n50937 = ~n5530 & n50763;
  assign n50938 = ~pi735 & pi1135;
  assign n50939 = ~pi743 & ~pi1135;
  assign n50940 = pi1136 & ~n50939;
  assign n50941 = pi1136 & ~n50938;
  assign n50942 = ~n50939 & n50941;
  assign n50943 = ~n50938 & n50940;
  assign n50944 = ~pi1135 & ~pi1136;
  assign n50945 = pi859 & n50944;
  assign n50946 = pi1134 & ~n50945;
  assign n50947 = ~n65196 & n50946;
  assign n50948 = n50937 & ~n50947;
  assign n50949 = ~n50936 & n50948;
  assign n50950 = ~n50922 & ~n50949;
  assign n50951 = pi876 & n50944;
  assign n50952 = ~pi730 & pi1135;
  assign n50953 = ~pi748 & ~pi1135;
  assign n50954 = pi1136 & ~n50953;
  assign n50955 = pi1136 & ~n50952;
  assign n50956 = ~n50953 & n50955;
  assign n50957 = ~n50952 & n50954;
  assign n50958 = ~n50951 & ~n65197;
  assign n50959 = n50783 & ~n50958;
  assign n50960 = ~pi710 & pi1135;
  assign n50961 = pi1136 & ~n50960;
  assign n50962 = ~pi803 & ~pi1135;
  assign n50963 = pi789 & n50782;
  assign n50964 = ~n50962 & ~n50963;
  assign n50965 = pi803 & ~pi1136;
  assign n50966 = ~pi1135 & ~n50965;
  assign n50967 = pi710 & pi1136;
  assign n50968 = ~n50963 & ~n50967;
  assign n50969 = ~n50966 & n50968;
  assign n50970 = ~n50961 & ~n50962;
  assign n50971 = ~n50963 & n50970;
  assign n50972 = ~n50961 & n50964;
  assign n50973 = ~pi623 & n50780;
  assign n50974 = n50764 & ~n50973;
  assign n50975 = n50764 & ~n65198;
  assign n50976 = ~n50973 & n50975;
  assign n50977 = ~n65198 & n50974;
  assign n50978 = ~n50959 & ~n65199;
  assign n50979 = ~n5530 & ~n50978;
  assign n50980 = pi199 & ~pi1037;
  assign n50981 = ~pi199 & ~pi296;
  assign n50982 = ~n50804 & ~n50981;
  assign n50983 = ~n50804 & ~n50980;
  assign n50984 = ~n50981 & n50983;
  assign n50985 = ~n50980 & n50982;
  assign n50986 = pi412 & n50794;
  assign n50987 = n50793 & ~n50986;
  assign n50988 = pi388 & ~pi591;
  assign n50989 = pi592 & ~n50988;
  assign n50990 = ~n50987 & ~n50989;
  assign n50991 = pi455 & n50801;
  assign n50992 = ~n50990 & ~n50991;
  assign n50993 = pi436 & n5481;
  assign n50994 = pi588 & ~n50993;
  assign n50995 = n50804 & ~n50994;
  assign n50996 = ~n50992 & n50995;
  assign n50997 = ~n65200 & ~n50996;
  assign n50998 = n5530 & ~n50997;
  assign n50999 = ~n50979 & ~n50998;
  assign n51000 = ~pi643 & pi1135;
  assign n51001 = ~pi606 & ~pi1135;
  assign n51002 = pi1136 & ~n51001;
  assign n51003 = pi1136 & ~n51000;
  assign n51004 = ~n51001 & n51003;
  assign n51005 = ~n51000 & n51002;
  assign n51006 = pi812 & ~pi1135;
  assign n51007 = ~pi787 & pi1135;
  assign n51008 = ~pi1136 & ~n51007;
  assign n51009 = ~pi1136 & ~n51006;
  assign n51010 = ~n51007 & n51009;
  assign n51011 = ~n51006 & n51008;
  assign n51012 = ~n65201 & ~n65202;
  assign n51013 = n50764 & ~n51012;
  assign n51014 = ~pi746 & n50780;
  assign n51015 = ~pi729 & pi1135;
  assign n51016 = ~pi881 & ~pi1136;
  assign n51017 = ~n51015 & ~n51016;
  assign n51018 = n50784 & n51017;
  assign n51019 = ~n51014 & n51018;
  assign n51020 = ~n51013 & ~n51019;
  assign n51021 = ~n5530 & ~n51020;
  assign n51022 = pi410 & n50794;
  assign n51023 = n50793 & ~n51022;
  assign n51024 = pi386 & ~pi591;
  assign n51025 = pi592 & ~n51024;
  assign n51026 = ~n51023 & ~n51025;
  assign n51027 = pi361 & n50801;
  assign n51028 = ~n51026 & ~n51027;
  assign n51029 = pi434 & n5481;
  assign n51030 = pi588 & ~n51029;
  assign n51031 = n50804 & ~n51030;
  assign n51032 = ~n51028 & n51031;
  assign n51033 = pi199 & ~pi1059;
  assign n51034 = ~pi199 & ~pi293;
  assign n51035 = ~n50804 & ~n51034;
  assign n51036 = ~n50804 & ~n51033;
  assign n51037 = ~n51034 & n51036;
  assign n51038 = ~n51033 & n51035;
  assign n51039 = ~n51032 & ~n65203;
  assign n51040 = n5530 & ~n51039;
  assign n51041 = ~n51021 & ~n51040;
  assign n51042 = pi199 & ~pi1036;
  assign n51043 = ~pi199 & ~pi255;
  assign n51044 = ~n50804 & ~n51043;
  assign n51045 = ~n50804 & ~n51042;
  assign n51046 = ~n51043 & n51045;
  assign n51047 = ~n51042 & n51044;
  assign n51048 = pi389 & n50908;
  assign n51049 = pi413 & pi591;
  assign n51050 = ~pi592 & n51049;
  assign n51051 = ~n51048 & ~n51050;
  assign n51052 = ~pi590 & ~n51051;
  assign n51053 = pi450 & n50801;
  assign n51054 = ~pi588 & ~n51053;
  assign n51055 = ~n51052 & n51054;
  assign n51056 = pi438 & n5481;
  assign n51057 = pi588 & ~n51056;
  assign n51058 = n50804 & ~n51057;
  assign n51059 = ~n51055 & n51058;
  assign n51060 = ~n65204 & ~n51059;
  assign n51061 = n5530 & ~n51060;
  assign n51062 = ~pi665 & pi1136;
  assign n51063 = ~pi791 & ~pi1136;
  assign n51064 = pi1135 & ~n51063;
  assign n51065 = pi1135 & ~n51062;
  assign n51066 = ~n51063 & n51065;
  assign n51067 = ~n51062 & n51064;
  assign n51068 = ~pi621 & pi1136;
  assign n51069 = ~pi810 & ~pi1136;
  assign n51070 = ~pi1135 & ~n51069;
  assign n51071 = ~pi1135 & ~n51068;
  assign n51072 = ~n51069 & n51071;
  assign n51073 = ~n51068 & n51070;
  assign n51074 = ~n65205 & ~n65206;
  assign n51075 = n50764 & ~n51074;
  assign n51076 = ~pi739 & n50780;
  assign n51077 = ~pi874 & ~pi1136;
  assign n51078 = ~pi690 & pi1135;
  assign n51079 = ~n51077 & ~n51078;
  assign n51080 = n50784 & n51079;
  assign n51081 = ~n51076 & n51080;
  assign n51082 = ~n51075 & ~n51081;
  assign n51083 = ~n5530 & ~n51082;
  assign n51084 = ~n51061 & ~n51083;
  assign n51085 = pi590 & ~pi592;
  assign n51086 = pi357 & n51085;
  assign n51087 = pi382 & n50792;
  assign n51088 = ~n51086 & ~n51087;
  assign n51089 = ~pi591 & ~n51088;
  assign n51090 = pi406 & ~pi592;
  assign n51091 = n50794 & n51090;
  assign n51092 = ~n51089 & ~n51091;
  assign n51093 = ~pi588 & ~n51092;
  assign n51094 = pi588 & ~pi590;
  assign n51095 = ~pi591 & ~pi592;
  assign n51096 = pi430 & n51095;
  assign n51097 = pi430 & n51094;
  assign n51098 = n51095 & n51097;
  assign n51099 = n51094 & n51096;
  assign n51100 = ~n51093 & ~n65207;
  assign n51101 = n50804 & ~n51100;
  assign n51102 = pi200 & pi1067;
  assign n51103 = ~pi200 & pi1044;
  assign n51104 = ~pi199 & ~n51103;
  assign n51105 = ~pi199 & ~n51102;
  assign n51106 = ~n51103 & n51105;
  assign n51107 = ~n51102 & n51104;
  assign n51108 = pi199 & ~pi1076;
  assign n51109 = ~n50804 & ~n51108;
  assign n51110 = ~n65208 & n51109;
  assign n51111 = ~n51101 & ~n51110;
  assign n51112 = n5530 & ~n51111;
  assign n51113 = pi860 & n50944;
  assign n51114 = pi728 & pi1135;
  assign n51115 = pi744 & ~pi1135;
  assign n51116 = pi1136 & ~n51115;
  assign n51117 = pi1136 & ~n51114;
  assign n51118 = ~n51115 & n51117;
  assign n51119 = ~n51114 & n51116;
  assign n51120 = ~n51113 & ~n65209;
  assign n51121 = n50783 & ~n51120;
  assign n51122 = pi1136 & ~n50763;
  assign n51123 = ~pi1134 & ~n51122;
  assign n51124 = pi657 & pi1135;
  assign n51125 = ~pi652 & ~pi1135;
  assign n51126 = pi1136 & ~n51125;
  assign n51127 = pi1136 & ~n51124;
  assign n51128 = ~n51125 & n51127;
  assign n51129 = ~n51124 & n51126;
  assign n51130 = pi813 & n50763;
  assign n51131 = n50944 & n51130;
  assign n51132 = ~n65210 & ~n51131;
  assign n51133 = n51123 & ~n51132;
  assign n51134 = ~n51121 & ~n51133;
  assign n51135 = ~n5530 & ~n51134;
  assign n51136 = ~n51112 & ~n51135;
  assign n51137 = pi351 & n51085;
  assign n51138 = pi376 & n50792;
  assign n51139 = ~n51137 & ~n51138;
  assign n51140 = ~pi591 & ~n51139;
  assign n51141 = pi401 & ~pi592;
  assign n51142 = n50794 & n51141;
  assign n51143 = ~n51140 & ~n51142;
  assign n51144 = ~pi588 & ~n51143;
  assign n51145 = pi426 & n51095;
  assign n51146 = pi426 & n51094;
  assign n51147 = n51095 & n51146;
  assign n51148 = n51094 & n51145;
  assign n51149 = ~n51144 & ~n65211;
  assign n51150 = n50804 & ~n51149;
  assign n51151 = ~pi200 & pi1049;
  assign n51152 = pi200 & pi1036;
  assign n51153 = pi200 & ~pi1036;
  assign n51154 = ~pi200 & ~pi1049;
  assign n51155 = ~n51153 & ~n51154;
  assign n51156 = ~n51151 & ~n51152;
  assign n51157 = ~pi199 & ~n65212;
  assign n51158 = pi199 & ~pi1079;
  assign n51159 = ~n50804 & ~n51158;
  assign n51160 = ~n51157 & n51159;
  assign n51161 = ~n51150 & ~n51160;
  assign n51162 = n5530 & ~n51161;
  assign n51163 = pi798 & n50944;
  assign n51164 = pi655 & pi1135;
  assign n51165 = ~pi658 & ~pi1135;
  assign n51166 = pi1136 & ~n51165;
  assign n51167 = pi1136 & ~n51164;
  assign n51168 = ~n51165 & n51167;
  assign n51169 = ~n51164 & n51166;
  assign n51170 = ~n51163 & ~n65213;
  assign n51171 = n50764 & ~n51170;
  assign n51172 = pi752 & n50780;
  assign n51173 = ~pi703 & pi1135;
  assign n51174 = ~pi843 & ~pi1136;
  assign n51175 = ~n51173 & ~n51174;
  assign n51176 = n50784 & n51175;
  assign n51177 = ~n51172 & n51176;
  assign n51178 = ~n51171 & ~n51177;
  assign n51179 = ~n5530 & ~n51178;
  assign n51180 = ~n51162 & ~n51179;
  assign n51181 = pi352 & n51085;
  assign n51182 = pi317 & n50792;
  assign n51183 = ~n51181 & ~n51182;
  assign n51184 = ~pi591 & ~n51183;
  assign n51185 = pi402 & ~pi592;
  assign n51186 = n50794 & n51185;
  assign n51187 = ~n51184 & ~n51186;
  assign n51188 = ~pi588 & ~n51187;
  assign n51189 = pi427 & n51095;
  assign n51190 = pi427 & n51094;
  assign n51191 = n51095 & n51190;
  assign n51192 = n51094 & n51189;
  assign n51193 = ~n51188 & ~n65214;
  assign n51194 = n50804 & ~n51193;
  assign n51195 = ~pi200 & pi1084;
  assign n51196 = pi200 & pi1065;
  assign n51197 = pi200 & ~pi1065;
  assign n51198 = ~pi200 & ~pi1084;
  assign n51199 = ~n51197 & ~n51198;
  assign n51200 = ~n51195 & ~n51196;
  assign n51201 = ~pi199 & ~n65215;
  assign n51202 = pi199 & ~pi1078;
  assign n51203 = ~n50804 & ~n51202;
  assign n51204 = ~n51201 & n51203;
  assign n51205 = ~n51194 & ~n51204;
  assign n51206 = n5530 & ~n51205;
  assign n51207 = pi649 & pi1135;
  assign n51208 = ~pi656 & ~pi1135;
  assign n51209 = pi1136 & ~n51208;
  assign n51210 = pi1136 & ~n51207;
  assign n51211 = ~n51208 & n51210;
  assign n51212 = ~n51207 & n51209;
  assign n51213 = pi801 & n50944;
  assign n51214 = ~pi1134 & ~n51213;
  assign n51215 = ~n65216 & n51214;
  assign n51216 = pi770 & ~pi1135;
  assign n51217 = ~pi726 & pi1135;
  assign n51218 = pi1136 & ~n51217;
  assign n51219 = pi1136 & ~n51216;
  assign n51220 = ~n51217 & n51219;
  assign n51221 = ~n51216 & n51218;
  assign n51222 = pi844 & n50944;
  assign n51223 = pi1134 & ~n51222;
  assign n51224 = ~n65217 & n51223;
  assign n51225 = n50937 & ~n51224;
  assign n51226 = n50937 & ~n51215;
  assign n51227 = ~n51224 & n51226;
  assign n51228 = ~n51215 & n51225;
  assign n51229 = ~n51206 & ~n65218;
  assign n51230 = pi370 & n50908;
  assign n51231 = pi395 & pi591;
  assign n51232 = ~pi592 & n51231;
  assign n51233 = ~n51230 & ~n51232;
  assign n51234 = ~pi590 & ~n51233;
  assign n51235 = pi347 & n50801;
  assign n51236 = ~n51234 & ~n51235;
  assign n51237 = ~pi588 & n50804;
  assign n51238 = ~n51236 & n51237;
  assign n51239 = n5481 & n50804;
  assign n51240 = pi420 & pi588;
  assign n51241 = n51239 & n51240;
  assign n51242 = ~pi200 & ~pi304;
  assign n51243 = pi200 & ~pi1048;
  assign n51244 = ~n51242 & ~n51243;
  assign n51245 = pi200 & pi1048;
  assign n51246 = ~pi200 & pi304;
  assign n51247 = ~pi199 & ~n51246;
  assign n51248 = ~n51245 & n51247;
  assign n51249 = ~pi199 & ~n51244;
  assign n51250 = pi199 & ~pi1055;
  assign n51251 = ~n50804 & ~n51250;
  assign n51252 = ~n65219 & n51251;
  assign n51253 = n5530 & ~n51252;
  assign n51254 = n5530 & ~n51241;
  assign n51255 = ~n51252 & n51254;
  assign n51256 = ~n51241 & n51253;
  assign n51257 = ~n51238 & n65220;
  assign n51258 = pi753 & n50780;
  assign n51259 = pi702 & pi1135;
  assign n51260 = ~pi847 & ~pi1136;
  assign n51261 = ~n51259 & ~n51260;
  assign n51262 = n50784 & n51261;
  assign n51263 = ~n51258 & n51262;
  assign n51264 = pi1136 & n50763;
  assign n51265 = ~pi618 & ~pi1135;
  assign n51266 = ~pi627 & pi1135;
  assign n51267 = ~pi1134 & ~n51266;
  assign n51268 = ~pi1134 & ~n51265;
  assign n51269 = ~n51266 & n51268;
  assign n51270 = ~n51265 & n51267;
  assign n51271 = n51264 & n65221;
  assign n51272 = ~n5530 & ~n51271;
  assign n51273 = ~n51263 & n51272;
  assign n51274 = ~n51241 & ~n51252;
  assign n51275 = ~n51238 & n51274;
  assign n51276 = n5530 & ~n51275;
  assign n51277 = ~n51263 & ~n51271;
  assign n51278 = ~n5530 & ~n51277;
  assign n51279 = ~n51276 & ~n51278;
  assign n51280 = ~n51257 & ~n51273;
  assign n51281 = n50804 & n50908;
  assign n51282 = pi442 & n51281;
  assign n51283 = ~pi592 & n50804;
  assign n51284 = pi328 & pi591;
  assign n51285 = n51283 & n51284;
  assign n51286 = ~n51282 & ~n51285;
  assign n51287 = ~pi590 & ~n51286;
  assign n51288 = pi321 & n50804;
  assign n51289 = n50801 & n51288;
  assign n51290 = ~n51287 & ~n51289;
  assign n51291 = ~pi588 & ~n51290;
  assign n51292 = ~pi200 & ~pi305;
  assign n51293 = pi200 & ~pi1084;
  assign n51294 = ~n51292 & ~n51293;
  assign n51295 = pi200 & pi1084;
  assign n51296 = ~pi200 & pi305;
  assign n51297 = ~pi199 & ~n51296;
  assign n51298 = ~n51295 & n51297;
  assign n51299 = ~pi199 & ~n51294;
  assign n51300 = pi199 & ~pi1058;
  assign n51301 = ~n50804 & ~n51300;
  assign n51302 = ~n65223 & n51301;
  assign n51303 = n50804 & n51095;
  assign n51304 = pi459 & n51094;
  assign n51305 = n51303 & n51304;
  assign n51306 = n5530 & ~n51305;
  assign n51307 = ~n51302 & n51306;
  assign n51308 = ~n51291 & n51307;
  assign n51309 = pi754 & n50780;
  assign n51310 = pi709 & pi1135;
  assign n51311 = ~pi857 & ~pi1136;
  assign n51312 = ~n51310 & ~n51311;
  assign n51313 = n50763 & ~n50782;
  assign n51314 = pi1134 & ~n51311;
  assign n51315 = pi1134 & ~n51310;
  assign n51316 = ~n51311 & n51315;
  assign n51317 = ~n51310 & n51314;
  assign n51318 = n51313 & n65224;
  assign n51319 = n50784 & n51312;
  assign n51320 = ~n51309 & n65225;
  assign n51321 = ~pi609 & ~pi1135;
  assign n51322 = ~pi660 & pi1135;
  assign n51323 = ~pi1134 & ~n51322;
  assign n51324 = ~pi1134 & ~n51321;
  assign n51325 = ~n51322 & n51324;
  assign n51326 = ~n51321 & n51323;
  assign n51327 = n51264 & n65226;
  assign n51328 = ~n5530 & ~n51327;
  assign n51329 = ~n51320 & n51328;
  assign po865 = ~n51308 & ~n51329;
  assign n51331 = pi373 & n50908;
  assign n51332 = pi398 & pi591;
  assign n51333 = ~pi592 & n51332;
  assign n51334 = ~n51331 & ~n51333;
  assign n51335 = ~pi590 & ~n51334;
  assign n51336 = pi348 & n50801;
  assign n51337 = ~n51335 & ~n51336;
  assign n51338 = n51237 & ~n51337;
  assign n51339 = pi423 & pi588;
  assign n51340 = n51239 & n51339;
  assign n51341 = ~pi200 & ~pi306;
  assign n51342 = pi200 & ~pi1059;
  assign n51343 = ~n51341 & ~n51342;
  assign n51344 = pi200 & pi1059;
  assign n51345 = ~pi200 & pi306;
  assign n51346 = ~pi199 & ~n51345;
  assign n51347 = ~n51344 & n51346;
  assign n51348 = ~pi199 & ~n51343;
  assign n51349 = pi199 & ~pi1087;
  assign n51350 = ~n50804 & ~n51349;
  assign n51351 = ~n65227 & n51350;
  assign n51352 = n5530 & ~n51351;
  assign n51353 = n5530 & ~n51340;
  assign n51354 = ~n51351 & n51353;
  assign n51355 = ~n51340 & n51352;
  assign n51356 = ~n51338 & n65228;
  assign n51357 = pi755 & n50780;
  assign n51358 = pi725 & pi1135;
  assign n51359 = ~pi858 & ~pi1136;
  assign n51360 = ~n51358 & ~n51359;
  assign n51361 = n50784 & n51360;
  assign n51362 = ~n51357 & n51361;
  assign n51363 = ~pi630 & ~pi1135;
  assign n51364 = ~pi647 & pi1135;
  assign n51365 = ~pi1134 & ~n51364;
  assign n51366 = ~pi1134 & ~n51363;
  assign n51367 = ~n51364 & n51366;
  assign n51368 = ~n51363 & n51365;
  assign n51369 = n51264 & n65229;
  assign n51370 = ~n5530 & ~n51369;
  assign n51371 = ~n51362 & n51370;
  assign n51372 = ~n51340 & ~n51351;
  assign n51373 = ~n51338 & n51372;
  assign n51374 = n5530 & ~n51373;
  assign n51375 = ~n51362 & ~n51369;
  assign n51376 = ~n5530 & ~n51375;
  assign n51377 = ~n51374 & ~n51376;
  assign n51378 = ~n51356 & ~n51371;
  assign n51379 = ~pi644 & ~pi1135;
  assign n51380 = ~pi715 & pi1135;
  assign n51381 = ~pi1134 & ~n51380;
  assign n51382 = ~pi1134 & ~n51379;
  assign n51383 = ~n51380 & n51382;
  assign n51384 = ~n51379 & n51381;
  assign n51385 = n51264 & n65231;
  assign n51386 = pi751 & n50780;
  assign n51387 = pi701 & pi1135;
  assign n51388 = ~pi842 & ~pi1136;
  assign n51389 = ~n51387 & ~n51388;
  assign n51390 = pi1134 & ~n51388;
  assign n51391 = pi1134 & ~n51387;
  assign n51392 = ~n51388 & n51391;
  assign n51393 = ~n51387 & n51390;
  assign n51394 = n51313 & n65232;
  assign n51395 = n50784 & n51389;
  assign n51396 = ~n51386 & n65233;
  assign n51397 = ~n51385 & ~n51396;
  assign n51398 = ~n5530 & ~n51397;
  assign n51399 = pi374 & n50908;
  assign n51400 = pi400 & pi591;
  assign n51401 = ~pi592 & n51400;
  assign n51402 = ~n51399 & ~n51401;
  assign n51403 = ~pi590 & ~n51402;
  assign n51404 = pi350 & n50801;
  assign n51405 = ~n51403 & ~n51404;
  assign n51406 = ~pi588 & ~n51405;
  assign n51407 = pi425 & n51095;
  assign n51408 = pi425 & n51094;
  assign n51409 = n51095 & n51408;
  assign n51410 = n51094 & n51407;
  assign n51411 = n50804 & ~n65234;
  assign n51412 = ~n51406 & n51411;
  assign n51413 = pi1044 & n48474;
  assign n51414 = pi298 & n39538;
  assign n51415 = pi199 & pi1035;
  assign n51416 = ~n50804 & ~n51415;
  assign n51417 = ~n51414 & n51416;
  assign n51418 = ~n51413 & n51416;
  assign n51419 = ~n51414 & n51418;
  assign n51420 = ~n51413 & n51417;
  assign n51421 = n5530 & ~n65235;
  assign n51422 = ~n51412 & n51421;
  assign n51423 = ~n51398 & ~n51422;
  assign n51424 = pi371 & n50908;
  assign n51425 = pi396 & pi591;
  assign n51426 = ~pi592 & n51425;
  assign n51427 = ~n51424 & ~n51426;
  assign n51428 = ~pi590 & ~n51427;
  assign n51429 = pi322 & n50801;
  assign n51430 = ~n51428 & ~n51429;
  assign n51431 = n51237 & ~n51430;
  assign n51432 = pi421 & pi588;
  assign n51433 = n51239 & n51432;
  assign n51434 = ~pi200 & ~pi309;
  assign n51435 = pi200 & ~pi1072;
  assign n51436 = ~n51434 & ~n51435;
  assign n51437 = pi200 & pi1072;
  assign n51438 = ~pi200 & pi309;
  assign n51439 = ~pi199 & ~n51438;
  assign n51440 = ~n51437 & n51439;
  assign n51441 = ~pi199 & ~n51436;
  assign n51442 = pi199 & ~pi1051;
  assign n51443 = ~n50804 & ~n51442;
  assign n51444 = ~n65236 & n51443;
  assign n51445 = n5530 & ~n51444;
  assign n51446 = n5530 & ~n51433;
  assign n51447 = ~n51444 & n51446;
  assign n51448 = ~n51433 & n51445;
  assign n51449 = ~n51431 & n65237;
  assign n51450 = pi756 & n50780;
  assign n51451 = pi734 & pi1135;
  assign n51452 = ~pi854 & ~pi1136;
  assign n51453 = ~n51451 & ~n51452;
  assign n51454 = n50784 & n51453;
  assign n51455 = ~n51450 & n51454;
  assign n51456 = ~pi629 & ~pi1135;
  assign n51457 = ~pi628 & pi1135;
  assign n51458 = ~pi1134 & ~n51457;
  assign n51459 = ~pi1134 & ~n51456;
  assign n51460 = ~n51457 & n51459;
  assign n51461 = ~n51456 & n51458;
  assign n51462 = n51264 & n65238;
  assign n51463 = ~n5530 & ~n51462;
  assign n51464 = ~n51455 & n51463;
  assign n51465 = ~n51433 & ~n51444;
  assign n51466 = ~n51431 & n51465;
  assign n51467 = n5530 & ~n51466;
  assign n51468 = ~n51455 & ~n51462;
  assign n51469 = ~n5530 & ~n51468;
  assign n51470 = ~n51467 & ~n51469;
  assign n51471 = ~n51449 & ~n51464;
  assign n51472 = pi461 & n51085;
  assign n51473 = pi439 & n50792;
  assign n51474 = ~n51472 & ~n51473;
  assign n51475 = ~pi591 & ~n51474;
  assign n51476 = pi326 & ~pi592;
  assign n51477 = n50794 & n51476;
  assign n51478 = ~n51475 & ~n51477;
  assign n51479 = ~pi588 & ~n51478;
  assign n51480 = pi449 & n51095;
  assign n51481 = pi449 & n51094;
  assign n51482 = n51095 & n51481;
  assign n51483 = n51094 & n51480;
  assign n51484 = ~n51479 & ~n65240;
  assign n51485 = n50804 & ~n51484;
  assign n51486 = pi200 & pi1039;
  assign n51487 = ~pi200 & pi1053;
  assign n51488 = ~pi199 & ~n51487;
  assign n51489 = ~pi199 & ~n51486;
  assign n51490 = ~n51487 & n51489;
  assign n51491 = ~n51486 & n51488;
  assign n51492 = pi199 & ~pi1057;
  assign n51493 = ~n50804 & ~n51492;
  assign n51494 = ~n65241 & n51493;
  assign n51495 = ~n51485 & ~n51494;
  assign n51496 = n5530 & ~n51495;
  assign n51497 = pi867 & n50944;
  assign n51498 = pi697 & pi1135;
  assign n51499 = pi762 & ~pi1135;
  assign n51500 = pi1136 & ~n51499;
  assign n51501 = pi1136 & ~n51498;
  assign n51502 = ~n51499 & n51501;
  assign n51503 = ~n51498 & n51500;
  assign n51504 = ~n51497 & ~n65242;
  assign n51505 = n50783 & ~n51504;
  assign n51506 = pi693 & pi1135;
  assign n51507 = ~pi653 & ~pi1135;
  assign n51508 = pi1136 & ~n51507;
  assign n51509 = pi1136 & ~n51506;
  assign n51510 = ~n51507 & n51509;
  assign n51511 = ~n51506 & n51508;
  assign n51512 = pi816 & n50763;
  assign n51513 = n50944 & n51512;
  assign n51514 = ~n65243 & ~n51513;
  assign n51515 = n51123 & ~n51514;
  assign n51516 = ~n51505 & ~n51515;
  assign n51517 = ~n5530 & ~n51516;
  assign n51518 = ~n51496 & ~n51517;
  assign n51519 = pi440 & n51281;
  assign n51520 = pi329 & pi591;
  assign n51521 = n51283 & n51520;
  assign n51522 = ~n51519 & ~n51521;
  assign n51523 = ~pi590 & ~n51522;
  assign n51524 = pi349 & n50804;
  assign n51525 = n50801 & n51524;
  assign n51526 = ~n51523 & ~n51525;
  assign n51527 = ~pi588 & ~n51526;
  assign n51528 = ~pi200 & ~pi307;
  assign n51529 = pi200 & ~pi1053;
  assign n51530 = ~n51528 & ~n51529;
  assign n51531 = pi200 & pi1053;
  assign n51532 = ~pi200 & pi307;
  assign n51533 = ~pi199 & ~n51532;
  assign n51534 = ~n51531 & n51533;
  assign n51535 = ~pi199 & ~n51530;
  assign n51536 = pi199 & ~pi1043;
  assign n51537 = ~n50804 & ~n51536;
  assign n51538 = ~n65244 & n51537;
  assign n51539 = pi454 & n51094;
  assign n51540 = n51303 & n51539;
  assign n51541 = n5530 & ~n51540;
  assign n51542 = ~n51538 & n51541;
  assign n51543 = ~n51527 & n51542;
  assign n51544 = pi761 & n50780;
  assign n51545 = pi738 & pi1135;
  assign n51546 = ~pi845 & ~pi1136;
  assign n51547 = ~n51545 & ~n51546;
  assign n51548 = pi1134 & ~n51546;
  assign n51549 = pi1134 & ~n51545;
  assign n51550 = ~n51546 & n51549;
  assign n51551 = ~n51545 & n51548;
  assign n51552 = n51313 & n65245;
  assign n51553 = n50784 & n51547;
  assign n51554 = ~n51544 & n65246;
  assign n51555 = ~pi626 & ~pi1135;
  assign n51556 = ~pi641 & pi1135;
  assign n51557 = ~pi1134 & ~n51556;
  assign n51558 = ~pi1134 & ~n51555;
  assign n51559 = ~n51556 & n51558;
  assign n51560 = ~n51555 & n51557;
  assign n51561 = n51264 & n65247;
  assign n51562 = ~n5530 & ~n51561;
  assign n51563 = ~n51554 & n51562;
  assign po873 = ~n51543 & ~n51563;
  assign n51565 = ~pi591 & n4041;
  assign n51566 = pi377 & n50908;
  assign n51567 = pi318 & pi591;
  assign n51568 = ~pi592 & n51567;
  assign n51569 = ~n65248 & ~n51568;
  assign n51570 = ~pi590 & ~n51569;
  assign n51571 = pi462 & n50801;
  assign n51572 = ~n51570 & ~n51571;
  assign n51573 = n51237 & ~n51572;
  assign n51574 = ~pi200 & pi1048;
  assign n51575 = pi200 & pi1070;
  assign n51576 = pi200 & ~pi1070;
  assign n51577 = ~pi200 & ~pi1048;
  assign n51578 = ~n51576 & ~n51577;
  assign n51579 = ~n51574 & ~n51575;
  assign n51580 = ~pi199 & ~n65249;
  assign n51581 = pi199 & ~pi1074;
  assign n51582 = ~n50804 & ~n51581;
  assign n51583 = ~n51580 & n51582;
  assign n51584 = pi448 & pi588;
  assign n51585 = n51239 & n51584;
  assign n51586 = ~n51583 & ~n51585;
  assign n51587 = ~n51573 & n51586;
  assign n51588 = n5530 & ~n51587;
  assign n51589 = pi800 & n50944;
  assign n51590 = pi669 & pi1135;
  assign n51591 = ~pi645 & ~pi1135;
  assign n51592 = pi1136 & ~n51591;
  assign n51593 = pi1136 & ~n51590;
  assign n51594 = ~n51591 & n51593;
  assign n51595 = ~n51590 & n51592;
  assign n51596 = ~n51589 & ~n65250;
  assign n51597 = n50764 & ~n51596;
  assign n51598 = pi768 & n50780;
  assign n51599 = ~pi705 & pi1135;
  assign n51600 = ~pi839 & ~pi1136;
  assign n51601 = ~n51599 & ~n51600;
  assign n51602 = pi1134 & ~n51600;
  assign n51603 = pi1134 & ~n51599;
  assign n51604 = ~n51600 & n51603;
  assign n51605 = ~n51599 & n51602;
  assign n51606 = n51313 & n65251;
  assign n51607 = n50784 & n51601;
  assign n51608 = ~n51598 & n65252;
  assign n51609 = ~n51597 & ~n51608;
  assign n51610 = ~n5530 & ~n51609;
  assign n51611 = ~n51588 & ~n51610;
  assign n51612 = pi369 & n51281;
  assign n51613 = pi394 & pi591;
  assign n51614 = n51283 & n51613;
  assign n51615 = ~n51612 & ~n51614;
  assign n51616 = ~pi590 & ~n51615;
  assign n51617 = pi315 & n50804;
  assign n51618 = n50801 & n51617;
  assign n51619 = ~n51616 & ~n51618;
  assign n51620 = ~pi588 & ~n51619;
  assign n51621 = ~pi200 & ~pi303;
  assign n51622 = pi200 & ~pi1049;
  assign n51623 = ~n51621 & ~n51622;
  assign n51624 = pi200 & pi1049;
  assign n51625 = ~pi200 & pi303;
  assign n51626 = ~pi199 & ~n51625;
  assign n51627 = ~n51624 & n51626;
  assign n51628 = ~pi199 & ~n51623;
  assign n51629 = pi199 & ~pi1080;
  assign n51630 = ~n50804 & ~n51629;
  assign n51631 = ~n65253 & n51630;
  assign n51632 = pi419 & n51094;
  assign n51633 = n51303 & n51632;
  assign n51634 = n5530 & ~n51633;
  assign n51635 = ~n51631 & n51634;
  assign n51636 = ~n51620 & n51635;
  assign n51637 = pi767 & n50780;
  assign n51638 = pi698 & pi1135;
  assign n51639 = ~pi853 & ~pi1136;
  assign n51640 = ~n51638 & ~n51639;
  assign n51641 = pi1134 & ~n51639;
  assign n51642 = pi1134 & ~n51638;
  assign n51643 = ~n51639 & n51642;
  assign n51644 = ~n51638 & n51641;
  assign n51645 = n51313 & n65254;
  assign n51646 = n50784 & n51640;
  assign n51647 = ~n51637 & n65255;
  assign n51648 = ~pi608 & ~pi1135;
  assign n51649 = ~pi625 & pi1135;
  assign n51650 = ~pi1134 & ~n51649;
  assign n51651 = ~pi1134 & ~n51648;
  assign n51652 = ~n51649 & n51651;
  assign n51653 = ~n51648 & n51650;
  assign n51654 = n51264 & n65256;
  assign n51655 = ~n5530 & ~n51654;
  assign n51656 = ~n51647 & n51655;
  assign po875 = ~n51636 & ~n51656;
  assign n51658 = pi378 & n50908;
  assign n51659 = pi325 & pi591;
  assign n51660 = ~pi592 & n51659;
  assign n51661 = ~n51658 & ~n51660;
  assign n51662 = ~pi590 & ~n51661;
  assign n51663 = pi353 & n50801;
  assign n51664 = ~n51662 & ~n51663;
  assign n51665 = n51237 & ~n51664;
  assign n51666 = ~pi200 & pi1072;
  assign n51667 = pi200 & pi1062;
  assign n51668 = pi200 & ~pi1062;
  assign n51669 = ~pi200 & ~pi1072;
  assign n51670 = ~n51668 & ~n51669;
  assign n51671 = ~n51666 & ~n51667;
  assign n51672 = ~pi199 & ~n65257;
  assign n51673 = pi199 & ~pi1063;
  assign n51674 = ~n50804 & ~n51673;
  assign n51675 = ~n51672 & n51674;
  assign n51676 = pi451 & pi588;
  assign n51677 = n51239 & n51676;
  assign n51678 = ~n51675 & ~n51677;
  assign n51679 = ~n51665 & n51678;
  assign n51680 = n5530 & ~n51679;
  assign n51681 = pi807 & n50944;
  assign n51682 = pi650 & pi1135;
  assign n51683 = ~pi636 & ~pi1135;
  assign n51684 = pi1136 & ~n51683;
  assign n51685 = pi1136 & ~n51682;
  assign n51686 = ~n51683 & n51685;
  assign n51687 = ~n51682 & n51684;
  assign n51688 = ~n51681 & ~n65258;
  assign n51689 = n50764 & ~n51688;
  assign n51690 = pi774 & n50780;
  assign n51691 = ~pi687 & pi1135;
  assign n51692 = ~pi868 & ~pi1136;
  assign n51693 = ~n51691 & ~n51692;
  assign n51694 = pi1134 & ~n51692;
  assign n51695 = pi1134 & ~n51691;
  assign n51696 = ~n51692 & n51695;
  assign n51697 = ~n51691 & n51694;
  assign n51698 = n51313 & n65259;
  assign n51699 = n50784 & n51693;
  assign n51700 = ~n51690 & n65260;
  assign n51701 = ~n51689 & ~n51700;
  assign n51702 = ~n5530 & ~n51701;
  assign n51703 = ~n51680 & ~n51702;
  assign n51704 = pi356 & n51085;
  assign n51705 = pi381 & n50792;
  assign n51706 = ~n51704 & ~n51705;
  assign n51707 = ~pi591 & ~n51706;
  assign n51708 = pi405 & ~pi592;
  assign n51709 = n50794 & n51708;
  assign n51710 = ~n51707 & ~n51709;
  assign n51711 = ~pi588 & ~n51710;
  assign n51712 = pi445 & n51095;
  assign n51713 = pi445 & n51094;
  assign n51714 = n51095 & n51713;
  assign n51715 = n51094 & n51712;
  assign n51716 = ~n51711 & ~n65261;
  assign n51717 = n50804 & ~n51716;
  assign n51718 = pi200 & pi1040;
  assign n51719 = ~pi200 & pi1037;
  assign n51720 = ~pi199 & ~n51719;
  assign n51721 = ~pi199 & ~n51718;
  assign n51722 = ~n51719 & n51721;
  assign n51723 = ~n51718 & n51720;
  assign n51724 = pi199 & ~pi1081;
  assign n51725 = ~n50804 & ~n51724;
  assign n51726 = ~n65262 & n51725;
  assign n51727 = ~n51717 & ~n51726;
  assign n51728 = n5530 & ~n51727;
  assign n51729 = pi880 & n50944;
  assign n51730 = pi684 & pi1135;
  assign n51731 = pi750 & ~pi1135;
  assign n51732 = pi1136 & ~n51731;
  assign n51733 = pi1136 & ~n51730;
  assign n51734 = ~n51731 & n51733;
  assign n51735 = ~n51730 & n51732;
  assign n51736 = ~n51729 & ~n65263;
  assign n51737 = n50783 & ~n51736;
  assign n51738 = pi654 & pi1135;
  assign n51739 = ~pi651 & ~pi1135;
  assign n51740 = pi1136 & ~n51739;
  assign n51741 = pi1136 & ~n51738;
  assign n51742 = ~n51739 & n51741;
  assign n51743 = ~n51738 & n51740;
  assign n51744 = pi794 & n50763;
  assign n51745 = n50944 & n51744;
  assign n51746 = ~n65264 & ~n51745;
  assign n51747 = n51123 & ~n51746;
  assign n51748 = ~n51737 & ~n51747;
  assign n51749 = ~n5530 & ~n51748;
  assign n51750 = ~n51728 & ~n51749;
  assign n51751 = pi379 & n50908;
  assign n51752 = pi403 & pi591;
  assign n51753 = ~pi592 & n51752;
  assign n51754 = ~n51751 & ~n51753;
  assign n51755 = ~pi590 & ~n51754;
  assign n51756 = pi354 & n50801;
  assign n51757 = ~n51755 & ~n51756;
  assign n51758 = n51237 & ~n51757;
  assign n51759 = ~pi200 & pi1059;
  assign n51760 = pi200 & pi1069;
  assign n51761 = pi200 & ~pi1069;
  assign n51762 = ~pi200 & ~pi1059;
  assign n51763 = ~n51761 & ~n51762;
  assign n51764 = ~n51759 & ~n51760;
  assign n51765 = ~pi199 & ~n65265;
  assign n51766 = pi199 & ~pi1045;
  assign n51767 = ~n50804 & ~n51766;
  assign n51768 = ~n51765 & n51767;
  assign n51769 = pi428 & pi588;
  assign n51770 = n51239 & n51769;
  assign n51771 = ~n51768 & ~n51770;
  assign n51772 = ~n51758 & n51771;
  assign n51773 = n5530 & ~n51772;
  assign n51774 = ~pi851 & pi1134;
  assign n51775 = ~pi795 & ~pi1134;
  assign n51776 = ~pi1136 & ~n51775;
  assign n51777 = ~pi1136 & ~n51774;
  assign n51778 = ~n51775 & n51777;
  assign n51779 = ~n51774 & n51776;
  assign n51780 = pi776 & pi1134;
  assign n51781 = ~pi640 & ~pi1134;
  assign n51782 = pi1136 & ~n51781;
  assign n51783 = pi1136 & ~n51780;
  assign n51784 = ~n51781 & n51783;
  assign n51785 = ~n51780 & n51782;
  assign n51786 = ~n65266 & ~n65267;
  assign n51787 = ~pi1135 & ~n51786;
  assign n51788 = pi732 & ~pi1134;
  assign n51789 = pi694 & pi1134;
  assign n51790 = pi1135 & pi1136;
  assign n51791 = ~n51789 & n51790;
  assign n51792 = ~n51788 & n51790;
  assign n51793 = ~n51789 & n51792;
  assign n51794 = ~n51788 & n51791;
  assign n51795 = ~n51787 & ~n65268;
  assign n51796 = n50937 & ~n51795;
  assign n51797 = ~n51773 & ~n51796;
  assign n51798 = pi199 & ~pi1065;
  assign n51799 = ~pi199 & ~pi257;
  assign n51800 = ~n50804 & ~n51799;
  assign n51801 = ~n50804 & ~n51798;
  assign n51802 = ~n51799 & n51801;
  assign n51803 = ~n51798 & n51800;
  assign n51804 = pi365 & n50908;
  assign n51805 = pi334 & pi591;
  assign n51806 = ~pi592 & n51805;
  assign n51807 = ~n51804 & ~n51806;
  assign n51808 = ~pi590 & ~n51807;
  assign n51809 = pi323 & n50801;
  assign n51810 = ~pi588 & ~n51809;
  assign n51811 = ~n51808 & n51810;
  assign n51812 = pi464 & n5481;
  assign n51813 = pi588 & ~n51812;
  assign n51814 = n50804 & ~n51813;
  assign n51815 = ~n51811 & n51814;
  assign n51816 = ~n65269 & ~n51815;
  assign n51817 = n5530 & ~n51816;
  assign n51818 = ~pi634 & pi1136;
  assign n51819 = ~pi784 & ~pi1136;
  assign n51820 = pi1135 & ~n51819;
  assign n51821 = pi1135 & ~n51818;
  assign n51822 = ~n51819 & n51821;
  assign n51823 = ~n51818 & n51820;
  assign n51824 = ~pi633 & pi1136;
  assign n51825 = ~pi815 & ~pi1136;
  assign n51826 = ~pi1135 & ~n51825;
  assign n51827 = ~pi1135 & ~n51824;
  assign n51828 = ~n51825 & n51827;
  assign n51829 = ~n51824 & n51826;
  assign n51830 = ~n65270 & ~n65271;
  assign n51831 = n50764 & ~n51830;
  assign n51832 = ~pi766 & n50780;
  assign n51833 = ~pi855 & ~pi1136;
  assign n51834 = ~pi700 & pi1135;
  assign n51835 = ~n51833 & ~n51834;
  assign n51836 = n50784 & n51835;
  assign n51837 = ~n51832 & n51836;
  assign n51838 = ~n51831 & ~n51837;
  assign n51839 = ~n5530 & ~n51838;
  assign n51840 = ~n51817 & ~n51839;
  assign n51841 = pi404 & n50794;
  assign n51842 = n50793 & ~n51841;
  assign n51843 = pi380 & ~pi591;
  assign n51844 = pi592 & ~n51843;
  assign n51845 = ~n51842 & ~n51844;
  assign n51846 = pi355 & n50801;
  assign n51847 = ~n51845 & ~n51846;
  assign n51848 = pi429 & n5481;
  assign n51849 = pi588 & ~n51848;
  assign n51850 = n50804 & ~n51849;
  assign n51851 = ~n51847 & n51850;
  assign n51852 = pi199 & ~pi1084;
  assign n51853 = ~pi199 & ~pi292;
  assign n51854 = ~n50804 & ~n51853;
  assign n51855 = ~n50804 & ~n51852;
  assign n51856 = ~n51853 & n51855;
  assign n51857 = ~n51852 & n51854;
  assign n51858 = ~n51851 & ~n65272;
  assign n51859 = n5530 & ~n51858;
  assign n51860 = pi662 & pi1135;
  assign n51861 = pi614 & ~pi1135;
  assign n51862 = pi1136 & ~n51861;
  assign n51863 = pi1136 & ~n51860;
  assign n51864 = ~n51861 & n51863;
  assign n51865 = ~n51860 & n51862;
  assign n51866 = pi785 & pi1135;
  assign n51867 = pi811 & ~pi1135;
  assign n51868 = ~pi1136 & ~n51867;
  assign n51869 = ~pi1136 & ~n51866;
  assign n51870 = ~n51867 & n51869;
  assign n51871 = ~n51866 & n51868;
  assign n51872 = ~n65273 & ~n65274;
  assign n51873 = ~pi1134 & ~n51872;
  assign n51874 = ~pi727 & pi1135;
  assign n51875 = ~pi772 & ~pi1135;
  assign n51876 = pi1136 & ~n51875;
  assign n51877 = pi1136 & ~n51874;
  assign n51878 = ~n51875 & n51877;
  assign n51879 = ~n51874 & n51876;
  assign n51880 = pi872 & n50944;
  assign n51881 = pi1134 & ~n51880;
  assign n51882 = ~n65275 & n51881;
  assign n51883 = n50937 & ~n51882;
  assign n51884 = ~n51873 & n51883;
  assign n51885 = ~n51859 & ~n51884;
  assign n51886 = ~pi638 & pi1135;
  assign n51887 = ~pi607 & ~pi1135;
  assign n51888 = pi1136 & ~n51887;
  assign n51889 = pi1136 & ~n51886;
  assign n51890 = ~n51887 & n51889;
  assign n51891 = ~n51886 & n51888;
  assign n51892 = pi799 & ~pi1135;
  assign n51893 = ~pi790 & pi1135;
  assign n51894 = ~pi1136 & ~n51893;
  assign n51895 = ~pi1136 & ~n51892;
  assign n51896 = ~n51893 & n51895;
  assign n51897 = ~n51892 & n51894;
  assign n51898 = ~n65276 & ~n65277;
  assign n51899 = n50764 & ~n51898;
  assign n51900 = ~pi764 & n50780;
  assign n51901 = ~pi691 & pi1135;
  assign n51902 = ~pi873 & ~pi1136;
  assign n51903 = ~n51901 & ~n51902;
  assign n51904 = n50784 & n51903;
  assign n51905 = ~n51900 & n51904;
  assign n51906 = ~n51899 & ~n51905;
  assign n51907 = ~n5530 & ~n51906;
  assign n51908 = pi456 & n50794;
  assign n51909 = n50793 & ~n51908;
  assign n51910 = pi337 & ~pi591;
  assign n51911 = pi592 & ~n51910;
  assign n51912 = ~n51909 & ~n51911;
  assign n51913 = pi441 & n50801;
  assign n51914 = ~n51912 & ~n51913;
  assign n51915 = pi443 & n5481;
  assign n51916 = pi588 & ~n51915;
  assign n51917 = n50804 & ~n51916;
  assign n51918 = ~n51914 & n51917;
  assign n51919 = pi199 & ~pi1044;
  assign n51920 = ~pi199 & ~pi297;
  assign n51921 = ~n50804 & ~n51920;
  assign n51922 = ~n50804 & ~n51919;
  assign n51923 = ~n51920 & n51922;
  assign n51924 = ~n51919 & n51921;
  assign n51925 = ~n51918 & ~n65278;
  assign n51926 = n5530 & ~n51925;
  assign n51927 = ~n51907 & ~n51926;
  assign n51928 = pi319 & n50794;
  assign n51929 = n50793 & ~n51928;
  assign n51930 = pi338 & ~pi591;
  assign n51931 = pi592 & ~n51930;
  assign n51932 = ~n51929 & ~n51931;
  assign n51933 = pi458 & n50801;
  assign n51934 = ~n51932 & ~n51933;
  assign n51935 = pi444 & n5481;
  assign n51936 = pi588 & ~n51935;
  assign n51937 = n50804 & ~n51936;
  assign n51938 = ~n51934 & n51937;
  assign n51939 = pi199 & ~pi1072;
  assign n51940 = ~pi199 & ~pi294;
  assign n51941 = ~n50804 & ~n51940;
  assign n51942 = ~n50804 & ~n51939;
  assign n51943 = ~n51940 & n51942;
  assign n51944 = ~n51939 & n51941;
  assign n51945 = ~n51938 & ~n65279;
  assign n51946 = n5530 & ~n51945;
  assign n51947 = pi681 & pi1136;
  assign n51948 = pi792 & ~pi1136;
  assign n51949 = pi1135 & ~n51948;
  assign n51950 = pi1135 & ~n51947;
  assign n51951 = ~n51948 & n51950;
  assign n51952 = ~n51947 & n51949;
  assign n51953 = pi642 & pi1136;
  assign n51954 = ~pi809 & ~pi1136;
  assign n51955 = ~pi1135 & ~n51954;
  assign n51956 = ~pi1135 & ~n51953;
  assign n51957 = ~n51954 & n51956;
  assign n51958 = ~n51953 & n51955;
  assign n51959 = ~n65280 & ~n65281;
  assign n51960 = ~pi1134 & ~n51959;
  assign n51961 = ~pi699 & pi1135;
  assign n51962 = ~pi763 & ~pi1135;
  assign n51963 = pi1136 & ~n51962;
  assign n51964 = pi1136 & ~n51961;
  assign n51965 = ~n51962 & n51964;
  assign n51966 = ~n51961 & n51963;
  assign n51967 = pi871 & n50944;
  assign n51968 = pi1134 & ~n51967;
  assign n51969 = ~n65282 & n51968;
  assign n51970 = n50937 & ~n51969;
  assign n51971 = ~n51960 & n51970;
  assign n51972 = ~n51946 & ~n51971;
  assign n51973 = pi199 & ~pi1062;
  assign n51974 = ~pi199 & ~pi258;
  assign n51975 = ~n50804 & ~n51974;
  assign n51976 = ~n50804 & ~n51973;
  assign n51977 = ~n51974 & n51976;
  assign n51978 = ~n51973 & n51975;
  assign n51979 = pi364 & n50908;
  assign n51980 = pi391 & pi591;
  assign n51981 = ~pi592 & n51980;
  assign n51982 = ~n51979 & ~n51981;
  assign n51983 = ~pi590 & ~n51982;
  assign n51984 = pi343 & n50801;
  assign n51985 = ~pi588 & ~n51984;
  assign n51986 = ~n51983 & n51985;
  assign n51987 = pi415 & n5481;
  assign n51988 = pi588 & ~n51987;
  assign n51989 = n50804 & ~n51988;
  assign n51990 = ~n51986 & n51989;
  assign n51991 = ~n65283 & ~n51990;
  assign n51992 = n5530 & ~n51991;
  assign n51993 = ~pi612 & ~pi1135;
  assign n51994 = pi695 & pi1135;
  assign n51995 = ~pi1134 & ~n51994;
  assign n51996 = ~pi1134 & ~n51993;
  assign n51997 = ~n51994 & n51996;
  assign n51998 = ~n51993 & n51995;
  assign n51999 = n51264 & n65284;
  assign n52000 = pi745 & n50780;
  assign n52001 = pi723 & pi1135;
  assign n52002 = ~pi852 & ~pi1136;
  assign n52003 = ~n52001 & ~n52002;
  assign n52004 = n50784 & n52003;
  assign n52005 = ~n52000 & n52004;
  assign n52006 = ~n51999 & ~n52005;
  assign n52007 = ~n5530 & ~n52006;
  assign n52008 = ~n51992 & ~n52007;
  assign n52009 = pi199 & ~pi1040;
  assign n52010 = ~pi199 & ~pi261;
  assign n52011 = ~n50804 & ~n52010;
  assign n52012 = ~n50804 & ~n52009;
  assign n52013 = ~n52010 & n52012;
  assign n52014 = ~n52009 & n52011;
  assign n52015 = pi447 & n50908;
  assign n52016 = pi333 & pi591;
  assign n52017 = ~pi592 & n52016;
  assign n52018 = ~n52015 & ~n52017;
  assign n52019 = ~pi590 & ~n52018;
  assign n52020 = pi327 & n50801;
  assign n52021 = ~pi588 & ~n52020;
  assign n52022 = ~n52019 & n52021;
  assign n52023 = pi453 & n5481;
  assign n52024 = pi588 & ~n52023;
  assign n52025 = n50804 & ~n52024;
  assign n52026 = ~n52022 & n52025;
  assign n52027 = ~n65285 & ~n52026;
  assign n52028 = n5530 & ~n52027;
  assign n52029 = ~pi611 & ~pi1135;
  assign n52030 = pi646 & pi1135;
  assign n52031 = ~pi1134 & ~n52030;
  assign n52032 = ~pi1134 & ~n52029;
  assign n52033 = ~n52030 & n52032;
  assign n52034 = ~n52029 & n52031;
  assign n52035 = n51264 & n65286;
  assign n52036 = pi741 & n50780;
  assign n52037 = pi724 & pi1135;
  assign n52038 = ~pi865 & ~pi1136;
  assign n52039 = ~n52037 & ~n52038;
  assign n52040 = n50784 & n52039;
  assign n52041 = ~n52036 & n52040;
  assign n52042 = ~n52035 & ~n52041;
  assign n52043 = ~n5530 & ~n52042;
  assign n52044 = ~n52028 & ~n52043;
  assign n52045 = pi199 & ~pi1069;
  assign n52046 = ~pi199 & ~pi259;
  assign n52047 = ~n50804 & ~n52046;
  assign n52048 = ~n50804 & ~n52045;
  assign n52049 = ~n52046 & n52048;
  assign n52050 = ~n52045 & n52047;
  assign n52051 = pi366 & n50908;
  assign n52052 = pi335 & pi591;
  assign n52053 = ~pi592 & n52052;
  assign n52054 = ~n52051 & ~n52053;
  assign n52055 = ~pi590 & ~n52054;
  assign n52056 = pi344 & n50801;
  assign n52057 = ~pi588 & ~n52056;
  assign n52058 = ~n52055 & n52057;
  assign n52059 = pi416 & n5481;
  assign n52060 = pi588 & ~n52059;
  assign n52061 = n50804 & ~n52060;
  assign n52062 = ~n52058 & n52061;
  assign n52063 = ~n65287 & ~n52062;
  assign n52064 = n5530 & ~n52063;
  assign n52065 = ~pi620 & ~pi1135;
  assign n52066 = pi635 & pi1135;
  assign n52067 = ~pi1134 & ~n52066;
  assign n52068 = ~pi1134 & ~n52065;
  assign n52069 = ~n52066 & n52068;
  assign n52070 = ~n52065 & n52067;
  assign n52071 = n51264 & n65288;
  assign n52072 = pi742 & n50780;
  assign n52073 = pi704 & pi1135;
  assign n52074 = ~pi870 & ~pi1136;
  assign n52075 = ~n52073 & ~n52074;
  assign n52076 = n50784 & n52075;
  assign n52077 = ~n52072 & n52076;
  assign n52078 = ~n52071 & ~n52077;
  assign n52079 = ~n5530 & ~n52078;
  assign n52080 = ~n52064 & ~n52079;
  assign n52081 = pi199 & ~pi1067;
  assign n52082 = ~pi199 & ~pi260;
  assign n52083 = ~n50804 & ~n52082;
  assign n52084 = ~n50804 & ~n52081;
  assign n52085 = ~n52082 & n52084;
  assign n52086 = ~n52081 & n52083;
  assign n52087 = pi368 & n50908;
  assign n52088 = pi393 & pi591;
  assign n52089 = ~pi592 & n52088;
  assign n52090 = ~n52087 & ~n52089;
  assign n52091 = ~pi590 & ~n52090;
  assign n52092 = pi346 & n50801;
  assign n52093 = ~pi588 & ~n52092;
  assign n52094 = ~n52091 & n52093;
  assign n52095 = pi418 & n5481;
  assign n52096 = pi588 & ~n52095;
  assign n52097 = n50804 & ~n52096;
  assign n52098 = ~n52094 & n52097;
  assign n52099 = ~n65289 & ~n52098;
  assign n52100 = n5530 & ~n52099;
  assign n52101 = ~pi613 & ~pi1135;
  assign n52102 = pi632 & pi1135;
  assign n52103 = ~pi1134 & ~n52102;
  assign n52104 = ~pi1134 & ~n52101;
  assign n52105 = ~n52102 & n52104;
  assign n52106 = ~n52101 & n52103;
  assign n52107 = n51264 & n65290;
  assign n52108 = pi760 & n50780;
  assign n52109 = pi688 & pi1135;
  assign n52110 = ~pi856 & ~pi1136;
  assign n52111 = ~n52109 & ~n52110;
  assign n52112 = n50784 & n52111;
  assign n52113 = ~n52108 & n52112;
  assign n52114 = ~n52107 & ~n52113;
  assign n52115 = ~n5530 & ~n52114;
  assign n52116 = ~n52100 & ~n52115;
  assign n52117 = pi199 & ~pi1039;
  assign n52118 = ~pi199 & ~pi251;
  assign n52119 = ~n50804 & ~n52118;
  assign n52120 = ~n50804 & ~n52117;
  assign n52121 = ~n52118 & n52120;
  assign n52122 = ~n52117 & n52119;
  assign n52123 = pi367 & n50908;
  assign n52124 = pi392 & pi591;
  assign n52125 = ~pi592 & n52124;
  assign n52126 = ~n52123 & ~n52125;
  assign n52127 = ~pi590 & ~n52126;
  assign n52128 = pi345 & n50801;
  assign n52129 = ~pi588 & ~n52128;
  assign n52130 = ~n52127 & n52129;
  assign n52131 = pi417 & n5481;
  assign n52132 = pi588 & ~n52131;
  assign n52133 = n50804 & ~n52132;
  assign n52134 = ~n52130 & n52133;
  assign n52135 = ~n65291 & ~n52134;
  assign n52136 = n5530 & ~n52135;
  assign n52137 = ~pi610 & ~pi1135;
  assign n52138 = pi631 & pi1135;
  assign n52139 = ~pi1134 & ~n52138;
  assign n52140 = ~pi1134 & ~n52137;
  assign n52141 = ~n52138 & n52140;
  assign n52142 = ~n52137 & n52139;
  assign n52143 = n51264 & n65292;
  assign n52144 = pi757 & n50780;
  assign n52145 = pi686 & pi1135;
  assign n52146 = ~pi848 & ~pi1136;
  assign n52147 = ~n52145 & ~n52146;
  assign n52148 = n50784 & n52147;
  assign n52149 = ~n52144 & n52148;
  assign n52150 = ~n52143 & ~n52149;
  assign n52151 = ~n5530 & ~n52150;
  assign n52152 = ~n52136 & ~n52151;
  assign n52153 = pi897 & n39538;
  assign n52154 = ~pi476 & n48474;
  assign n52155 = ~n52153 & ~n52154;
  assign n52156 = ~n65241 & ~n52155;
  assign n52157 = pi251 & n52155;
  assign n52158 = ~n52156 & ~n52157;
  assign n52159 = ~n65212 & ~n52155;
  assign n52160 = ~pi255 & n52155;
  assign n52161 = n65212 & ~n52155;
  assign n52162 = pi255 & n52155;
  assign n52163 = ~n52161 & ~n52162;
  assign n52164 = ~n52159 & ~n52160;
  assign n52165 = ~n65249 & ~n52155;
  assign n52166 = ~pi256 & n52155;
  assign n52167 = n65249 & ~n52155;
  assign n52168 = pi256 & n52155;
  assign n52169 = ~n52167 & ~n52168;
  assign n52170 = ~n52165 & ~n52166;
  assign n52171 = ~n65215 & ~n52155;
  assign n52172 = ~pi257 & n52155;
  assign n52173 = n65215 & ~n52155;
  assign n52174 = pi257 & n52155;
  assign n52175 = ~n52173 & ~n52174;
  assign n52176 = ~n52171 & ~n52172;
  assign n52177 = ~n65257 & ~n52155;
  assign n52178 = ~pi258 & n52155;
  assign n52179 = n65257 & ~n52155;
  assign n52180 = pi258 & n52155;
  assign n52181 = ~n52179 & ~n52180;
  assign n52182 = ~n52177 & ~n52178;
  assign n52183 = ~n65265 & ~n52155;
  assign n52184 = ~pi259 & n52155;
  assign n52185 = n65265 & ~n52155;
  assign n52186 = pi259 & n52155;
  assign n52187 = ~n52185 & ~n52186;
  assign n52188 = ~n52183 & ~n52184;
  assign n52189 = ~n65208 & ~n52155;
  assign n52190 = pi260 & n52155;
  assign n52191 = ~n52189 & ~n52190;
  assign n52192 = ~n65262 & ~n52155;
  assign n52193 = pi261 & n52155;
  assign n52194 = ~n52192 & ~n52193;
  assign n52195 = ~pi290 & pi476;
  assign n52196 = ~pi476 & ~pi1048;
  assign n52197 = ~pi476 & pi1048;
  assign n52198 = pi290 & pi476;
  assign n52199 = ~n52197 & ~n52198;
  assign n52200 = ~n52195 & ~n52196;
  assign n52201 = ~pi291 & pi476;
  assign n52202 = ~pi476 & ~pi1049;
  assign n52203 = ~pi476 & pi1049;
  assign n52204 = pi291 & pi476;
  assign n52205 = ~n52203 & ~n52204;
  assign n52206 = ~n52201 & ~n52202;
  assign n52207 = ~pi292 & pi476;
  assign n52208 = ~pi476 & ~pi1084;
  assign n52209 = ~pi476 & pi1084;
  assign n52210 = pi292 & pi476;
  assign n52211 = ~n52209 & ~n52210;
  assign n52212 = ~n52207 & ~n52208;
  assign n52213 = ~pi293 & pi476;
  assign n52214 = ~pi476 & ~pi1059;
  assign n52215 = ~pi476 & pi1059;
  assign n52216 = pi293 & pi476;
  assign n52217 = ~n52215 & ~n52216;
  assign n52218 = ~n52213 & ~n52214;
  assign n52219 = ~pi294 & pi476;
  assign n52220 = ~pi476 & ~pi1072;
  assign n52221 = ~pi476 & pi1072;
  assign n52222 = pi294 & pi476;
  assign n52223 = ~n52221 & ~n52222;
  assign n52224 = ~n52219 & ~n52220;
  assign n52225 = ~pi295 & pi476;
  assign n52226 = ~pi476 & ~pi1053;
  assign n52227 = ~pi476 & pi1053;
  assign n52228 = pi295 & pi476;
  assign n52229 = ~n52227 & ~n52228;
  assign n52230 = ~n52225 & ~n52226;
  assign n52231 = ~pi296 & pi476;
  assign n52232 = ~pi476 & ~pi1037;
  assign n52233 = ~pi476 & pi1037;
  assign n52234 = pi296 & pi476;
  assign n52235 = ~n52233 & ~n52234;
  assign n52236 = ~n52231 & ~n52232;
  assign n52237 = ~pi297 & pi476;
  assign n52238 = ~pi476 & ~pi1044;
  assign n52239 = ~pi476 & pi1044;
  assign n52240 = pi297 & pi476;
  assign n52241 = ~n52239 & ~n52240;
  assign n52242 = ~n52237 & ~n52238;
  assign n52243 = pi375 & n51281;
  assign n52244 = pi399 & pi591;
  assign n52245 = n51283 & n52244;
  assign n52246 = ~n52243 & ~n52245;
  assign n52247 = ~pi590 & ~n52246;
  assign n52248 = pi316 & n50804;
  assign n52249 = n50801 & n52248;
  assign n52250 = ~n52247 & ~n52249;
  assign n52251 = ~pi588 & ~n52250;
  assign n52252 = ~pi200 & ~pi308;
  assign n52253 = pi200 & ~pi1037;
  assign n52254 = ~n52252 & ~n52253;
  assign n52255 = pi200 & pi1037;
  assign n52256 = ~pi200 & pi308;
  assign n52257 = ~pi199 & ~n52256;
  assign n52258 = ~n52255 & n52257;
  assign n52259 = ~pi199 & ~n52254;
  assign n52260 = pi199 & ~pi1047;
  assign n52261 = ~n50804 & ~n52260;
  assign n52262 = ~n65306 & n52261;
  assign n52263 = pi424 & n51094;
  assign n52264 = n51303 & n52263;
  assign n52265 = n5530 & ~n52264;
  assign n52266 = ~n52262 & n52265;
  assign n52267 = ~n52251 & n52266;
  assign n52268 = pi777 & n50780;
  assign n52269 = pi737 & pi1135;
  assign n52270 = ~pi838 & ~pi1136;
  assign n52271 = ~n52269 & ~n52270;
  assign n52272 = pi1134 & ~n52270;
  assign n52273 = pi1134 & ~n52269;
  assign n52274 = ~n52270 & n52273;
  assign n52275 = ~n52269 & n52272;
  assign n52276 = n51313 & n65307;
  assign n52277 = n50784 & n52271;
  assign n52278 = ~n52268 & n65308;
  assign n52279 = ~pi619 & ~pi1135;
  assign n52280 = ~pi648 & pi1135;
  assign n52281 = ~pi1134 & ~n52280;
  assign n52282 = ~pi1134 & ~n52279;
  assign n52283 = ~n52280 & n52282;
  assign n52284 = ~n52279 & n52281;
  assign n52285 = n51264 & n65309;
  assign n52286 = ~n5530 & ~n52285;
  assign n52287 = ~n52278 & n52286;
  assign po890 = ~n52267 & ~n52287;
  assign n52289 = ~n62455 & ~n49875;
  assign n52290 = ~n50378 & n52289;
  assign n52291 = pi219 & ~n50603;
  assign n52292 = ~n49273 & n52291;
  assign n52293 = ~n49276 & n50665;
  assign n52294 = ~n52292 & ~n52293;
  assign n52295 = ~n49378 & ~n50680;
  assign n52296 = ~n52294 & ~n52295;
  assign n52297 = n62455 & ~n52296;
  assign n52298 = ~n49283 & ~n50306;
  assign n52299 = n52297 & ~n52298;
  assign n52300 = ~n52290 & ~n52299;
  assign n52301 = ~pi1151 & ~n52300;
  assign n52302 = n62455 & ~n49922;
  assign n52303 = ~n49239 & n52302;
  assign n52304 = ~n50168 & n52289;
  assign n52305 = n62455 & ~n50676;
  assign n52306 = pi219 & n49424;
  assign n52307 = n52305 & ~n52306;
  assign n52308 = ~n52304 & ~n52307;
  assign n52309 = ~n52303 & n52308;
  assign n52310 = pi1151 & ~n52309;
  assign n52311 = pi268 & ~n52310;
  assign n52312 = ~n52301 & n52311;
  assign n52313 = ~n62455 & ~n49886;
  assign n52314 = ~n50359 & n52313;
  assign n52315 = pi219 & ~n49284;
  assign n52316 = ~n50642 & ~n52315;
  assign n52317 = ~n49275 & ~n52316;
  assign n52318 = ~n50389 & ~n52317;
  assign n52319 = n62455 & ~n52318;
  assign n52320 = ~n52314 & ~n52319;
  assign n52321 = ~pi1151 & ~n52320;
  assign n52322 = ~pi219 & n49291;
  assign n52323 = ~n52291 & ~n52322;
  assign n52324 = n62455 & ~n52323;
  assign n52325 = ~n50379 & n52313;
  assign n52326 = ~n50377 & n52289;
  assign n52327 = n52314 & ~n52326;
  assign n52328 = ~n52325 & ~n52327;
  assign n52329 = ~n52324 & n52328;
  assign n52330 = pi1151 & ~n52329;
  assign n52331 = ~pi268 & ~n52330;
  assign n52332 = ~n52321 & n52331;
  assign n52333 = ~n52312 & ~n52332;
  assign n52334 = pi1150 & ~n52333;
  assign n52335 = ~n50476 & n52289;
  assign n52336 = pi219 & ~n49923;
  assign n52337 = ~n50642 & ~n52336;
  assign n52338 = n49270 & ~n52337;
  assign n52339 = n62455 & ~n52338;
  assign n52340 = ~n52335 & ~n52339;
  assign n52341 = pi1151 & ~n52340;
  assign n52342 = n62455 & ~n50680;
  assign n52343 = ~n52336 & n52342;
  assign n52344 = ~n52326 & ~n52343;
  assign n52345 = ~pi1151 & ~n52344;
  assign n52346 = pi268 & ~n52345;
  assign n52347 = ~n52341 & n52346;
  assign n52348 = n62455 & ~n52294;
  assign n52349 = ~n52325 & ~n52348;
  assign n52350 = pi1151 & ~n52349;
  assign n52351 = ~n49878 & n52313;
  assign n52352 = ~pi219 & ~n49313;
  assign n52353 = ~n49259 & ~n52352;
  assign n52354 = n52324 & n52353;
  assign n52355 = ~n52351 & ~n52354;
  assign n52356 = ~pi1151 & ~n52355;
  assign n52357 = ~pi268 & ~n52356;
  assign n52358 = ~n52350 & n52357;
  assign n52359 = ~n52347 & ~n52358;
  assign n52360 = ~pi1150 & ~n52359;
  assign n52361 = pi1152 & ~n52360;
  assign n52362 = ~pi1150 & ~n52347;
  assign n52363 = ~n52358 & n52362;
  assign n52364 = pi1150 & ~n52332;
  assign n52365 = ~n52312 & n52364;
  assign n52366 = ~n52363 & ~n52365;
  assign n52367 = pi1152 & ~n52366;
  assign n52368 = ~n52334 & n52361;
  assign n52369 = n62455 & ~n50645;
  assign n52370 = ~n50642 & n52369;
  assign n52371 = ~n50655 & ~n52370;
  assign n52372 = pi1151 & ~n52371;
  assign n52373 = ~n50168 & n50654;
  assign n52374 = ~n52307 & ~n52373;
  assign n52375 = n49243 & ~n52374;
  assign n52376 = ~pi1151 & n52375;
  assign n52377 = pi268 & ~n52376;
  assign n52378 = ~n52372 & n52377;
  assign n52379 = pi219 & ~n62455;
  assign n52380 = ~n49283 & n52379;
  assign n52381 = ~n50380 & ~n52380;
  assign n52382 = ~n52297 & n52381;
  assign n52383 = pi1151 & n52382;
  assign n52384 = ~n49327 & n52305;
  assign n52385 = ~n49878 & ~n52380;
  assign n52386 = ~n52384 & n52385;
  assign n52387 = ~pi1151 & n52386;
  assign n52388 = ~pi268 & ~n52387;
  assign n52389 = ~n52383 & n52388;
  assign n52390 = ~n52378 & ~n52389;
  assign n52391 = ~pi1150 & ~n52390;
  assign n52392 = ~n50378 & n50654;
  assign n52393 = n52294 & n52302;
  assign n52394 = ~n52392 & ~n52393;
  assign n52395 = ~pi1151 & ~n52394;
  assign n52396 = pi1151 & ~n52374;
  assign n52397 = pi268 & ~n52396;
  assign n52398 = ~n52395 & n52397;
  assign n52399 = n62455 & ~n49337;
  assign n52400 = n52317 & n52399;
  assign n52401 = ~n52327 & ~n52400;
  assign n52402 = ~pi1151 & ~n52401;
  assign n52403 = ~n49243 & ~n52374;
  assign n52404 = ~n52386 & ~n52403;
  assign n52405 = pi1151 & ~n52404;
  assign n52406 = ~pi268 & ~n52405;
  assign n52407 = ~n52402 & n52406;
  assign n52408 = ~pi1151 & n52394;
  assign n52409 = pi1151 & n52374;
  assign n52410 = pi268 & ~n52409;
  assign n52411 = ~n52395 & ~n52396;
  assign n52412 = pi268 & ~n52411;
  assign n52413 = ~n52408 & n52410;
  assign n52414 = ~pi1151 & n52401;
  assign n52415 = pi1151 & n52404;
  assign n52416 = ~pi268 & ~n52415;
  assign n52417 = ~n52402 & ~n52405;
  assign n52418 = ~pi268 & ~n52417;
  assign n52419 = ~n52414 & n52416;
  assign n52420 = ~n65311 & ~n65312;
  assign n52421 = ~n52398 & ~n52407;
  assign n52422 = pi1150 & ~n65311;
  assign n52423 = ~n65312 & n52422;
  assign n52424 = pi1150 & n65313;
  assign n52425 = ~pi1152 & ~n65314;
  assign n52426 = ~n52391 & n52425;
  assign n52427 = ~pi1152 & ~n65313;
  assign n52428 = pi1152 & ~n52332;
  assign n52429 = ~n52312 & n52428;
  assign n52430 = ~n52427 & ~n52429;
  assign n52431 = pi1150 & ~n52430;
  assign n52432 = pi1152 & ~n52350;
  assign n52433 = pi1152 & ~n52356;
  assign n52434 = ~n52350 & n52433;
  assign n52435 = ~n52356 & n52432;
  assign n52436 = ~pi1152 & ~n52387;
  assign n52437 = ~n52383 & n52436;
  assign n52438 = ~n65315 & ~n52437;
  assign n52439 = ~pi268 & ~n52438;
  assign n52440 = pi1151 & n52340;
  assign n52441 = ~pi1151 & n52344;
  assign n52442 = pi1152 & ~n52441;
  assign n52443 = ~n52440 & n52442;
  assign n52444 = pi1151 & n52371;
  assign n52445 = ~pi1151 & ~n52375;
  assign n52446 = ~pi1152 & ~n52445;
  assign n52447 = ~n52444 & n52446;
  assign n52448 = pi268 & ~n52447;
  assign n52449 = ~n52443 & n52448;
  assign n52450 = ~pi1150 & ~n52449;
  assign n52451 = ~n52439 & n52450;
  assign n52452 = ~n52431 & ~n52451;
  assign n52453 = ~n65310 & ~n52426;
  assign n52454 = n49536 & ~n65316;
  assign n52455 = ~n65014 & n50453;
  assign n52456 = n62455 & n49832;
  assign n52457 = ~n65014 & ~n50453;
  assign n52458 = n65014 & ~n49445;
  assign n52459 = ~n39538 & n65317;
  assign n52460 = ~n52457 & ~n52459;
  assign n52461 = ~n52455 & ~n52456;
  assign n52462 = pi1151 & n65318;
  assign n52463 = pi1152 & n52462;
  assign n52464 = n62455 & ~n48478;
  assign n52465 = ~n48548 & ~n52464;
  assign n52466 = pi1151 & ~n52465;
  assign n52467 = ~pi1152 & ~n52466;
  assign n52468 = ~pi1151 & n50528;
  assign n52469 = ~pi1150 & ~n52468;
  assign n52470 = ~pi1150 & ~n52467;
  assign n52471 = ~n52468 & n52470;
  assign n52472 = ~n52467 & n52469;
  assign n52473 = ~n52463 & n65319;
  assign n52474 = ~pi199 & n65014;
  assign n52475 = ~pi219 & ~n65014;
  assign n52476 = ~n52474 & ~n52475;
  assign n52477 = pi1151 & ~n52476;
  assign n52478 = ~pi211 & ~n65014;
  assign n52479 = n62455 & n49461;
  assign n52480 = ~n52478 & ~n52479;
  assign n52481 = ~n52477 & n52480;
  assign n52482 = ~pi1152 & n52476;
  assign n52483 = pi1150 & ~n52482;
  assign n52484 = pi1150 & ~n52481;
  assign n52485 = ~n52482 & n52484;
  assign n52486 = pi1152 & ~n52480;
  assign n52487 = n52476 & ~n52486;
  assign n52488 = ~pi1151 & n52480;
  assign n52489 = pi1150 & ~n52488;
  assign n52490 = ~n52487 & n52489;
  assign n52491 = ~n52481 & n52483;
  assign n52492 = ~n52473 & ~n65320;
  assign n52493 = pi1091 & n52492;
  assign n52494 = ~pi268 & ~pi1091;
  assign n52495 = ~n49536 & ~n52494;
  assign n52496 = pi268 & pi1152;
  assign n52497 = n65320 & ~n52496;
  assign n52498 = ~n52473 & ~n52497;
  assign n52499 = pi1091 & ~n52498;
  assign n52500 = pi1152 & n52484;
  assign n52501 = pi1152 & n65320;
  assign n52502 = pi1091 & ~n65321;
  assign n52503 = pi268 & ~n52502;
  assign n52504 = ~n52499 & ~n52503;
  assign n52505 = ~n49536 & ~n52504;
  assign n52506 = ~n52493 & n52495;
  assign n52507 = ~pi230 & ~n65322;
  assign n52508 = ~n52454 & n52507;
  assign n52509 = pi230 & ~n65320;
  assign n52510 = ~n52473 & n52509;
  assign n52511 = ~n52454 & ~n65322;
  assign n52512 = ~pi230 & ~n52511;
  assign n52513 = pi230 & ~n52492;
  assign n52514 = ~n52512 & ~n52513;
  assign n52515 = ~n52508 & ~n52510;
  assign po1102 = pi230 & n2923;
  assign n52517 = ~pi212 & ~pi214;
  assign n52518 = ~pi211 & ~n52517;
  assign n52519 = pi219 & ~n52518;
  assign n52520 = ~n62455 & ~n52519;
  assign n52521 = pi1142 & ~n39346;
  assign n52522 = ~pi211 & pi1143;
  assign n52523 = n39342 & n52522;
  assign n52524 = pi211 & pi1143;
  assign n52525 = ~pi211 & pi1144;
  assign n52526 = ~n52524 & ~n52525;
  assign n52527 = ~pi212 & pi214;
  assign n52528 = pi212 & ~pi214;
  assign n52529 = ~n52527 & ~n52528;
  assign n52530 = ~n39342 & ~n52517;
  assign n52531 = ~n39342 & ~n52526;
  assign n52532 = ~n52517 & n52531;
  assign n52533 = ~n52526 & ~n65324;
  assign n52534 = ~n52523 & ~n65325;
  assign n52535 = ~pi219 & ~n52534;
  assign n52536 = ~n52521 & ~n52535;
  assign n52537 = n52520 & ~n52536;
  assign n52538 = pi199 & pi1142;
  assign n52539 = ~pi200 & ~n52538;
  assign n52540 = ~pi199 & pi1144;
  assign n52541 = n52539 & ~n52540;
  assign n52542 = ~pi199 & pi1143;
  assign n52543 = pi200 & ~n52542;
  assign n52544 = ~n52541 & ~n52543;
  assign n52545 = ~pi299 & ~n52544;
  assign n52546 = ~pi207 & ~n52545;
  assign n52547 = n52539 & ~n52542;
  assign n52548 = pi207 & ~pi299;
  assign n52549 = ~pi199 & pi1142;
  assign n52550 = pi200 & ~n52549;
  assign n52551 = n52548 & ~n52550;
  assign n52552 = ~n52547 & n52551;
  assign n52553 = ~n52546 & ~n52552;
  assign n52554 = pi208 & ~n52553;
  assign n52555 = pi207 & ~pi208;
  assign n52556 = n52544 & n52555;
  assign n52557 = ~n52554 & ~n52556;
  assign n52558 = ~pi299 & ~n52557;
  assign n52559 = pi211 & pi1142;
  assign n52560 = pi1142 & n64625;
  assign n52561 = n39342 & n52559;
  assign n52562 = ~n52523 & ~n65326;
  assign n52563 = ~n52523 & ~n52531;
  assign n52564 = ~n65326 & n52563;
  assign n52565 = ~n52531 & n52562;
  assign n52566 = ~pi219 & n65327;
  assign n52567 = ~pi211 & pi1142;
  assign n52568 = pi219 & ~n52567;
  assign n52569 = pi299 & ~n52517;
  assign n52570 = ~n52568 & n52569;
  assign n52571 = ~n52566 & n52570;
  assign n52572 = ~n52558 & ~n52571;
  assign n52573 = pi299 & ~n52526;
  assign n52574 = ~pi214 & ~n52558;
  assign n52575 = ~n52573 & n52574;
  assign n52576 = ~n52522 & ~n52559;
  assign n52577 = pi299 & ~n52576;
  assign n52578 = pi214 & ~n52577;
  assign n52579 = ~n52558 & n52578;
  assign n52580 = pi212 & ~n52579;
  assign n52581 = ~n52575 & n52580;
  assign n52582 = ~n52558 & ~n52573;
  assign n52583 = ~pi212 & ~n52582;
  assign n52584 = ~pi212 & ~n52574;
  assign n52585 = ~n52582 & n52584;
  assign n52586 = ~n52574 & n52583;
  assign n52587 = ~pi219 & ~n65328;
  assign n52588 = ~pi219 & ~n52581;
  assign n52589 = ~n65328 & n52588;
  assign n52590 = ~n52581 & n52587;
  assign n52591 = ~n52518 & n52558;
  assign n52592 = ~pi299 & n52557;
  assign n52593 = pi299 & ~pi1142;
  assign n52594 = n52518 & ~n52593;
  assign n52595 = ~n52592 & n52594;
  assign n52596 = pi219 & ~n52595;
  assign n52597 = pi219 & ~n52591;
  assign n52598 = ~n52595 & n52597;
  assign n52599 = ~n52591 & n52596;
  assign n52600 = n62455 & ~n65330;
  assign n52601 = ~n65329 & n52600;
  assign n52602 = n62455 & ~n52572;
  assign n52603 = ~n52537 & ~n65331;
  assign n52604 = pi213 & n52603;
  assign n52605 = ~n49542 & ~n50084;
  assign n52606 = pi214 & n52605;
  assign n52607 = ~n49651 & ~n49654;
  assign n52608 = ~pi214 & n52607;
  assign n52609 = pi212 & ~n52608;
  assign n52610 = pi212 & ~n52606;
  assign n52611 = ~n52608 & n52610;
  assign n52612 = ~pi214 & ~n52607;
  assign n52613 = pi214 & ~n52605;
  assign n52614 = ~n52612 & ~n52613;
  assign n52615 = pi212 & ~n52614;
  assign n52616 = ~n52606 & n52609;
  assign n52617 = ~n49388 & ~n49541;
  assign n52618 = pi214 & ~n52617;
  assign n52619 = ~pi212 & n52618;
  assign n52620 = n52527 & ~n52617;
  assign n52621 = ~pi219 & ~n65333;
  assign n52622 = ~pi212 & ~n52618;
  assign n52623 = pi212 & n52614;
  assign n52624 = ~n52622 & ~n52623;
  assign n52625 = ~n65332 & ~n65333;
  assign n52626 = ~pi219 & ~n65334;
  assign n52627 = ~n65332 & n52621;
  assign n52628 = ~pi211 & pi214;
  assign n52629 = pi1155 & n52628;
  assign n52630 = ~pi212 & ~n52629;
  assign n52631 = ~pi214 & ~n49653;
  assign n52632 = n39342 & ~n50176;
  assign n52633 = ~n52631 & ~n52632;
  assign n52634 = ~n52630 & n52633;
  assign n52635 = pi219 & ~n52634;
  assign n52636 = ~n62455 & ~n52635;
  assign n52637 = ~n65335 & n52636;
  assign n52638 = ~pi213 & ~n52637;
  assign n52639 = n49607 & n52527;
  assign n52640 = pi299 & pi1154;
  assign n52641 = ~pi214 & ~n52640;
  assign n52642 = pi299 & pi1153;
  assign n52643 = pi214 & ~n52642;
  assign n52644 = pi212 & ~n52643;
  assign n52645 = pi212 & ~n52641;
  assign n52646 = ~n52643 & n52645;
  assign n52647 = ~n52641 & n52644;
  assign n52648 = ~n52639 & ~n65336;
  assign n52649 = n39423 & ~n52648;
  assign n52650 = n50523 & n65334;
  assign n52651 = ~n52649 & ~n52650;
  assign n52652 = ~n52558 & n52651;
  assign n52653 = n62455 & ~n52652;
  assign n52654 = n52638 & ~n52653;
  assign n52655 = pi209 & ~n52654;
  assign n52656 = ~n52604 & n52655;
  assign n52657 = pi199 & n50077;
  assign n52658 = pi1155 & n49457;
  assign n52659 = ~pi299 & n65337;
  assign n52660 = ~pi1156 & ~n65146;
  assign n52661 = pi199 & ~pi1155;
  assign n52662 = ~pi200 & ~pi1155;
  assign n52663 = n49599 & ~n52662;
  assign n52664 = n49599 & ~n52661;
  assign n52665 = ~n52660 & n65338;
  assign n52666 = pi207 & n52665;
  assign n52667 = ~pi208 & ~n52666;
  assign n52668 = ~pi199 & ~pi1155;
  assign n52669 = ~pi1154 & ~n52668;
  assign n52670 = n50534 & n52669;
  assign n52671 = pi1154 & ~n50262;
  assign n52672 = n48567 & n50077;
  assign n52673 = n39538 & n49619;
  assign n52674 = pi1154 & n49598;
  assign n52675 = ~n50538 & n52674;
  assign n52676 = ~n65339 & ~n52675;
  assign n52677 = n52671 & ~n52676;
  assign n52678 = pi1155 & ~n50531;
  assign n52679 = ~pi1155 & n49458;
  assign n52680 = n48570 & n52662;
  assign n52681 = pi1153 & n65340;
  assign n52682 = ~n52678 & ~n52681;
  assign n52683 = ~pi1154 & ~n52682;
  assign n52684 = ~n49851 & ~n50546;
  assign n52685 = pi1154 & ~n52684;
  assign n52686 = ~n52683 & ~n52685;
  assign n52687 = ~pi299 & ~n52686;
  assign n52688 = ~n52670 & ~n52677;
  assign n52689 = pi207 & n65341;
  assign n52690 = pi1156 & n48567;
  assign n52691 = pi1156 & n49623;
  assign n52692 = ~n49594 & n52690;
  assign n52693 = ~n39538 & ~n49622;
  assign n52694 = n49610 & n52693;
  assign n52695 = ~n49622 & n49639;
  assign n52696 = ~n65342 & ~n65343;
  assign n52697 = ~pi207 & ~n52696;
  assign n52698 = pi208 & ~n52697;
  assign n52699 = pi207 & ~n65341;
  assign n52700 = ~pi207 & n52696;
  assign n52701 = ~n52699 & ~n52700;
  assign n52702 = pi208 & ~n52701;
  assign n52703 = ~n52689 & n52698;
  assign n52704 = ~n52667 & ~n65344;
  assign n52705 = ~pi1157 & ~n52704;
  assign n52706 = pi1156 & ~n52661;
  assign n52707 = n49595 & n52706;
  assign n52708 = ~pi1156 & ~n52661;
  assign n52709 = ~pi1156 & n49461;
  assign n52710 = ~n52661 & n52709;
  assign n52711 = n49461 & n52708;
  assign n52712 = ~n52707 & ~n65345;
  assign n52713 = pi207 & ~n52712;
  assign n52714 = ~pi208 & ~n52713;
  assign n52715 = ~n65344 & ~n52714;
  assign n52716 = pi1157 & ~n52715;
  assign n52717 = ~n52705 & ~n52716;
  assign n52718 = pi211 & ~n52717;
  assign n52719 = ~pi214 & ~n52717;
  assign n52720 = ~pi212 & ~n52719;
  assign n52721 = pi207 & n52686;
  assign n52722 = ~pi207 & ~n49607;
  assign n52723 = n52696 & n52722;
  assign n52724 = pi208 & ~n52723;
  assign n52725 = ~n52721 & n52724;
  assign n52726 = pi1155 & ~n49494;
  assign n52727 = ~n49607 & ~n50077;
  assign n52728 = ~n48567 & ~n65346;
  assign n52729 = pi1156 & ~n52728;
  assign n52730 = n49600 & ~n49831;
  assign n52731 = ~pi1156 & n49519;
  assign n52732 = ~pi1155 & ~n52731;
  assign n52733 = ~n49494 & ~n52732;
  assign n52734 = ~n52690 & ~n52733;
  assign n52735 = ~n52729 & ~n52730;
  assign n52736 = pi207 & n65347;
  assign n52737 = ~pi208 & pi1157;
  assign n52738 = ~pi208 & ~n52722;
  assign n52739 = pi1157 & n52738;
  assign n52740 = ~n52722 & n52737;
  assign n52741 = ~n52736 & n65348;
  assign n52742 = ~pi299 & n52660;
  assign n52743 = ~n49832 & ~n50209;
  assign n52744 = ~n52742 & n52743;
  assign n52745 = n52738 & n52744;
  assign n52746 = ~n52741 & ~n52745;
  assign n52747 = ~n52725 & n52746;
  assign n52748 = n52628 & n52747;
  assign n52749 = n52720 & ~n52748;
  assign n52750 = pi1154 & ~n65132;
  assign n52751 = n52696 & ~n52750;
  assign n52752 = ~pi207 & ~n52751;
  assign n52753 = ~pi299 & n52684;
  assign n52754 = pi1154 & ~n52753;
  assign n52755 = ~n52670 & ~n52754;
  assign n52756 = pi207 & ~n52755;
  assign n52757 = ~n52752 & ~n52756;
  assign n52758 = pi208 & ~n52757;
  assign n52759 = ~n49849 & ~n65346;
  assign n52760 = ~pi1156 & ~n52759;
  assign n52761 = pi1156 & ~n50078;
  assign n52762 = ~n52760 & ~n52761;
  assign n52763 = ~n52707 & n52759;
  assign n52764 = pi207 & n65349;
  assign n52765 = ~pi207 & ~pi299;
  assign n52766 = ~pi208 & ~n52765;
  assign n52767 = ~n52764 & n52766;
  assign n52768 = pi299 & ~pi1154;
  assign n52769 = pi1157 & ~n52768;
  assign n52770 = n52767 & n52769;
  assign n52771 = ~n52640 & ~n52666;
  assign n52772 = ~pi208 & ~n52771;
  assign n52773 = ~pi1157 & n52772;
  assign n52774 = ~n52770 & ~n52773;
  assign n52775 = ~n52758 & n52774;
  assign n52776 = ~pi211 & ~pi214;
  assign n52777 = n52775 & n52776;
  assign n52778 = pi1156 & ~n65337;
  assign n52779 = n49800 & n52778;
  assign n52780 = ~n52660 & ~n52779;
  assign n52781 = pi207 & n52780;
  assign n52782 = ~pi299 & ~n52781;
  assign n52783 = ~pi208 & ~n52782;
  assign n52784 = ~pi1157 & ~n52783;
  assign n52785 = pi1157 & ~n52767;
  assign n52786 = pi299 & ~pi1153;
  assign n52787 = ~n52785 & ~n52786;
  assign n52788 = ~pi1157 & n52783;
  assign n52789 = pi1157 & n52767;
  assign n52790 = ~n52784 & ~n52785;
  assign n52791 = ~n52788 & ~n52789;
  assign n52792 = ~n52786 & n65350;
  assign n52793 = ~n52784 & ~n52786;
  assign n52794 = ~n52785 & n52793;
  assign n52795 = ~n52784 & n52787;
  assign n52796 = pi1153 & ~n49519;
  assign n52797 = n52676 & ~n52796;
  assign n52798 = pi207 & ~n52797;
  assign n52799 = ~n49849 & ~n49851;
  assign n52800 = ~pi299 & ~n49614;
  assign n52801 = pi1156 & ~n65352;
  assign n52802 = pi299 & ~pi1155;
  assign n52803 = ~n49801 & ~n52802;
  assign n52804 = ~pi299 & ~n49830;
  assign n52805 = ~n52801 & n65353;
  assign n52806 = ~n52750 & ~n52801;
  assign n52807 = n65353 & n52806;
  assign n52808 = ~n52750 & n52805;
  assign n52809 = ~pi207 & ~n52786;
  assign n52810 = ~n65354 & n52809;
  assign n52811 = ~n52798 & ~n52810;
  assign n52812 = pi208 & ~n52811;
  assign n52813 = n52628 & ~n52812;
  assign n52814 = n52628 & ~n65351;
  assign n52815 = ~n52812 & n52814;
  assign n52816 = ~n65351 & n52813;
  assign n52817 = pi212 & ~n65355;
  assign n52818 = pi212 & ~n52777;
  assign n52819 = ~n65355 & n52818;
  assign n52820 = ~n52777 & n52817;
  assign n52821 = ~n52749 & ~n65356;
  assign n52822 = ~n52718 & ~n52821;
  assign n52823 = pi219 & ~n52822;
  assign n52824 = n52548 & n52797;
  assign n52825 = ~pi207 & n65354;
  assign n52826 = pi208 & ~n52825;
  assign n52827 = pi208 & ~n52824;
  assign n52828 = ~n52825 & n52827;
  assign n52829 = ~n52824 & n52826;
  assign n52830 = n52785 & ~n65357;
  assign n52831 = ~pi211 & ~n52830;
  assign n52832 = ~pi211 & ~n52705;
  assign n52833 = ~n52830 & n52832;
  assign n52834 = ~n52705 & n52831;
  assign n52835 = pi299 & pi1156;
  assign n52836 = pi207 & ~n52835;
  assign n52837 = ~n65343 & ~n52801;
  assign n52838 = ~pi207 & n52837;
  assign n52839 = ~pi207 & ~n52837;
  assign n52840 = pi207 & n52835;
  assign n52841 = ~n52839 & ~n52840;
  assign n52842 = ~n52836 & ~n52838;
  assign n52843 = ~n52689 & n65359;
  assign n52844 = pi208 & ~n52843;
  assign n52845 = ~n52660 & n52783;
  assign n52846 = ~n52713 & ~n52835;
  assign n52847 = n52737 & ~n52846;
  assign n52848 = ~n52845 & ~n52847;
  assign n52849 = ~n52844 & n52848;
  assign n52850 = pi211 & ~n52849;
  assign n52851 = pi214 & ~n52850;
  assign n52852 = ~n65358 & n52851;
  assign n52853 = n52720 & ~n52852;
  assign n52854 = n39343 & ~n52775;
  assign n52855 = ~n39343 & ~n52776;
  assign n52856 = ~n52747 & n52855;
  assign n52857 = n52776 & ~n52849;
  assign n52858 = ~n52856 & ~n52857;
  assign n52859 = ~n52854 & n52858;
  assign n52860 = pi212 & ~n52859;
  assign n52861 = ~pi219 & ~n52860;
  assign n52862 = ~n52853 & n52861;
  assign n52863 = n62455 & ~n52862;
  assign n52864 = ~n52853 & ~n52860;
  assign n52865 = ~pi219 & ~n52864;
  assign n52866 = n52527 & n52747;
  assign n52867 = ~n65351 & ~n52812;
  assign n52868 = pi214 & ~n52867;
  assign n52869 = ~pi214 & ~n52775;
  assign n52870 = pi212 & ~n52869;
  assign n52871 = ~n52868 & n52870;
  assign n52872 = ~n52866 & ~n52871;
  assign n52873 = ~pi211 & ~n52872;
  assign n52874 = ~n52518 & ~n52717;
  assign n52875 = pi219 & ~n52874;
  assign n52876 = ~n52873 & n52875;
  assign n52877 = ~n52865 & ~n52876;
  assign n52878 = n62455 & ~n52877;
  assign n52879 = ~n52823 & n52863;
  assign n52880 = n52638 & ~n65360;
  assign n52881 = pi299 & pi1143;
  assign n52882 = n52699 & ~n52881;
  assign n52883 = pi299 & ~pi1143;
  assign n52884 = n49833 & ~n52883;
  assign n52885 = ~pi1155 & n52881;
  assign n52886 = pi1154 & ~n65340;
  assign n52887 = ~n52885 & n52886;
  assign n52888 = ~n52884 & n52887;
  assign n52889 = n49622 & ~n52881;
  assign n52890 = ~pi1156 & ~n52889;
  assign n52891 = ~n52888 & n52890;
  assign n52892 = ~n65352 & ~n52883;
  assign n52893 = ~pi1154 & ~n52892;
  assign n52894 = pi1154 & ~n49610;
  assign n52895 = ~n52881 & n52894;
  assign n52896 = pi1156 & ~n52895;
  assign n52897 = ~n52893 & n52896;
  assign n52898 = ~n52891 & ~n52897;
  assign n52899 = ~pi207 & n52898;
  assign n52900 = pi208 & ~n52899;
  assign n52901 = pi208 & ~n52882;
  assign n52902 = ~n52899 & n52901;
  assign n52903 = ~n52882 & n52900;
  assign n52904 = n52788 & ~n52883;
  assign n52905 = pi207 & ~n52883;
  assign n52906 = ~n65349 & n52905;
  assign n52907 = ~n52881 & ~n52906;
  assign n52908 = n52737 & ~n52907;
  assign n52909 = ~pi211 & n39342;
  assign n52910 = pi211 & ~n65324;
  assign n52911 = pi211 & n52527;
  assign n52912 = pi212 & n52855;
  assign n52913 = ~n52911 & ~n52912;
  assign n52914 = ~n52909 & ~n52910;
  assign n52915 = ~n52908 & ~n65362;
  assign n52916 = ~n52904 & n52915;
  assign n52917 = ~n65361 & n52916;
  assign n52918 = pi299 & ~pi1144;
  assign n52919 = n49833 & ~n52918;
  assign n52920 = pi299 & pi1144;
  assign n52921 = ~pi1155 & n52920;
  assign n52922 = n52886 & ~n52921;
  assign n52923 = ~n52919 & n52922;
  assign n52924 = n49622 & ~n52920;
  assign n52925 = ~pi1156 & ~n52924;
  assign n52926 = ~n52923 & n52925;
  assign n52927 = ~n65352 & ~n52918;
  assign n52928 = ~pi1154 & ~n52927;
  assign n52929 = n52894 & ~n52920;
  assign n52930 = pi1156 & ~n52929;
  assign n52931 = ~n52928 & n52930;
  assign n52932 = ~n52926 & ~n52931;
  assign n52933 = ~pi207 & n52932;
  assign n52934 = n52699 & ~n52920;
  assign n52935 = pi208 & ~n52934;
  assign n52936 = pi208 & ~n52933;
  assign n52937 = ~n52934 & n52936;
  assign n52938 = ~n52933 & n52935;
  assign n52939 = n52788 & ~n52918;
  assign n52940 = pi207 & ~n52918;
  assign n52941 = ~n65349 & n52940;
  assign n52942 = ~n52920 & ~n52941;
  assign n52943 = n52737 & ~n52942;
  assign n52944 = n39424 & ~n52517;
  assign n52945 = ~pi211 & ~n65324;
  assign n52946 = ~n52943 & n65364;
  assign n52947 = ~n52939 & n52946;
  assign n52948 = ~n52939 & ~n52943;
  assign n52949 = ~n65363 & n52948;
  assign n52950 = ~pi211 & ~n52949;
  assign n52951 = ~n65324 & ~n52950;
  assign n52952 = ~pi211 & n52951;
  assign n52953 = ~n65363 & n52947;
  assign n52954 = ~n52904 & ~n52908;
  assign n52955 = ~n65361 & n52954;
  assign n52956 = ~n52909 & ~n52951;
  assign n52957 = n52955 & ~n52956;
  assign n52958 = ~n65365 & ~n52957;
  assign n52959 = n52909 & n52955;
  assign n52960 = pi211 & ~n52955;
  assign n52961 = ~n65324 & ~n52960;
  assign n52962 = ~n52950 & n52961;
  assign n52963 = n52951 & ~n52960;
  assign n52964 = ~n52959 & ~n65367;
  assign n52965 = ~n52917 & ~n65365;
  assign n52966 = ~pi219 & ~n65366;
  assign n52967 = ~pi219 & ~n52517;
  assign n52968 = ~n52518 & ~n52967;
  assign n52969 = ~n52717 & n52968;
  assign n52970 = ~n52593 & ~n52785;
  assign n52971 = ~n52593 & n65350;
  assign n52972 = ~n52593 & ~n52784;
  assign n52973 = ~n52785 & n52972;
  assign n52974 = ~n52784 & n52970;
  assign n52975 = pi299 & pi1142;
  assign n52976 = pi207 & ~n52975;
  assign n52977 = ~pi299 & n52686;
  assign n52978 = ~n52593 & ~n52977;
  assign n52979 = pi207 & ~n52978;
  assign n52980 = ~n65341 & n52976;
  assign n52981 = ~n52593 & ~n52806;
  assign n52982 = ~n65119 & ~n52975;
  assign n52983 = ~pi1154 & ~pi1156;
  assign n52984 = ~n52982 & n52983;
  assign n52985 = ~pi207 & ~n52984;
  assign n52986 = ~n52981 & n52985;
  assign n52987 = pi208 & ~n52986;
  assign n52988 = ~n65369 & n52987;
  assign n52989 = ~n39346 & ~n52968;
  assign n52990 = ~n52988 & n52989;
  assign n52991 = ~n65368 & n52989;
  assign n52992 = ~n52988 & n52991;
  assign n52993 = ~n65368 & n52990;
  assign n52994 = n62455 & ~n65370;
  assign n52995 = n62455 & ~n52969;
  assign n52996 = ~n65370 & n52995;
  assign n52997 = ~n52969 & n52994;
  assign n52998 = ~n52966 & n65371;
  assign n52999 = pi213 & ~n52537;
  assign n53000 = ~n52998 & n52999;
  assign n53001 = ~pi209 & ~n53000;
  assign n53002 = ~n52880 & n53001;
  assign n53003 = ~n52656 & ~n53002;
  assign n53004 = pi230 & ~n53003;
  assign n53005 = ~pi230 & ~pi233;
  assign n53006 = ~n53004 & ~n53005;
  assign n53007 = ~pi211 & pi1145;
  assign n53008 = pi211 & pi1144;
  assign n53009 = ~n53007 & ~n53008;
  assign n53010 = ~n39342 & n53009;
  assign n53011 = n39342 & n52526;
  assign n53012 = pi212 & ~n52526;
  assign n53013 = n65324 & ~n53012;
  assign n53014 = ~n52517 & ~n53011;
  assign n53015 = ~n52517 & ~n53010;
  assign n53016 = ~n53011 & n53015;
  assign n53017 = ~n53010 & ~n65372;
  assign n53018 = ~pi219 & ~n65373;
  assign n53019 = pi219 & ~n52522;
  assign n53020 = n52520 & ~n53019;
  assign n53021 = ~n53018 & n53020;
  assign n53022 = n50523 & n65373;
  assign n53023 = pi199 & pi1143;
  assign n53024 = ~pi200 & ~n53023;
  assign n53025 = ~n52540 & n53024;
  assign n53026 = pi208 & n52548;
  assign n53027 = ~n52543 & n53026;
  assign n53028 = ~n53025 & n53027;
  assign n53029 = ~pi199 & pi1145;
  assign n53030 = n53024 & ~n53029;
  assign n53031 = ~pi207 & ~pi208;
  assign n53032 = ~n38985 & ~n53031;
  assign n53033 = pi200 & ~n52540;
  assign n53034 = n53032 & ~n53033;
  assign n53035 = ~n53030 & n53034;
  assign n53036 = ~n53028 & ~n53035;
  assign n53037 = ~pi299 & ~n53036;
  assign n53038 = pi219 & ~n52517;
  assign n53039 = pi299 & n52522;
  assign n53040 = ~pi211 & n52881;
  assign n53041 = pi299 & n53038;
  assign n53042 = n52522 & n53041;
  assign n53043 = n53038 & n65374;
  assign n53044 = ~n53037 & ~n65375;
  assign n53045 = ~n53022 & ~n65375;
  assign n53046 = ~n53037 & n53045;
  assign n53047 = ~n53022 & n53044;
  assign n53048 = n62455 & ~n65376;
  assign n53049 = ~n53021 & ~n53048;
  assign n53050 = pi213 & n53049;
  assign n53051 = ~pi214 & n52617;
  assign n53052 = pi214 & n52607;
  assign n53053 = pi212 & ~n53052;
  assign n53054 = pi212 & ~n53051;
  assign n53055 = ~n53052 & n53054;
  assign n53056 = pi214 & ~n52607;
  assign n53057 = ~pi214 & ~n52617;
  assign n53058 = ~n53056 & ~n53057;
  assign n53059 = pi212 & ~n53058;
  assign n53060 = ~n53051 & n53053;
  assign n53061 = ~pi211 & pi1158;
  assign n53062 = ~n49406 & ~n53061;
  assign n53063 = n52527 & ~n53062;
  assign n53064 = ~pi219 & ~n53063;
  assign n53065 = ~pi219 & ~n65377;
  assign n53066 = ~n53063 & n53065;
  assign n53067 = ~n65377 & n53064;
  assign n53068 = ~pi212 & n52628;
  assign n53069 = pi1156 & n53068;
  assign n53070 = n49651 & n52527;
  assign n53071 = ~n62455 & n65379;
  assign n53072 = ~n50558 & ~n53071;
  assign n53073 = pi1155 & n52776;
  assign n53074 = ~pi214 & n49542;
  assign n53075 = pi214 & n49653;
  assign n53076 = pi1154 & n52628;
  assign n53077 = ~n65380 & ~n65381;
  assign n53078 = pi212 & ~n62455;
  assign n53079 = pi214 & ~n49653;
  assign n53080 = ~pi214 & ~n49542;
  assign n53081 = pi212 & ~n53080;
  assign n53082 = ~n53079 & n53081;
  assign n53083 = pi212 & ~n53077;
  assign n53084 = ~n62455 & n65382;
  assign n53085 = ~n53077 & n53078;
  assign n53086 = n53072 & ~n65383;
  assign n53087 = ~n65378 & ~n53086;
  assign n53088 = ~pi213 & ~n53087;
  assign n53089 = n50523 & ~n65378;
  assign n53090 = n52527 & n52835;
  assign n53091 = ~pi214 & ~n49607;
  assign n53092 = pi214 & ~n52640;
  assign n53093 = pi212 & ~n53092;
  assign n53094 = pi212 & ~n53091;
  assign n53095 = ~n53092 & n53094;
  assign n53096 = ~n53091 & n53093;
  assign n53097 = ~n53090 & ~n65384;
  assign n53098 = n39423 & ~n53097;
  assign n53099 = ~n53037 & ~n53098;
  assign n53100 = ~n53089 & n53099;
  assign n53101 = n62455 & ~n53100;
  assign n53102 = n53088 & ~n53101;
  assign n53103 = pi209 & ~n53102;
  assign n53104 = pi209 & ~n53050;
  assign n53105 = ~n53102 & n53104;
  assign n53106 = ~n53050 & n53103;
  assign n53107 = n49461 & n52555;
  assign n53108 = pi1158 & n48497;
  assign n53109 = ~pi199 & ~pi1158;
  assign n53110 = pi1156 & ~n53109;
  assign n53111 = ~pi1156 & ~n48497;
  assign n53112 = pi1158 & ~n53111;
  assign n53113 = ~n49596 & ~n53112;
  assign n53114 = ~n53108 & ~n53110;
  assign n53115 = n53107 & ~n65386;
  assign n53116 = pi207 & n52696;
  assign n53117 = ~pi207 & ~n52665;
  assign n53118 = pi208 & ~n53117;
  assign n53119 = ~n53116 & n53118;
  assign n53120 = ~n53115 & ~n53119;
  assign n53121 = ~pi1157 & ~n53120;
  assign n53122 = ~pi200 & ~pi1158;
  assign n53123 = ~pi199 & ~n53122;
  assign n53124 = ~n49613 & ~n53123;
  assign n53125 = ~pi1158 & ~n49599;
  assign n53126 = n49453 & ~n53125;
  assign n53127 = ~n53123 & ~n53126;
  assign n53128 = n52548 & ~n53127;
  assign n53129 = n52548 & ~n53124;
  assign n53130 = ~pi208 & n65387;
  assign n53131 = ~pi207 & n52712;
  assign n53132 = pi208 & ~n53131;
  assign n53133 = ~n53116 & n53132;
  assign n53134 = ~n53130 & ~n53133;
  assign n53135 = pi1157 & ~n53134;
  assign n53136 = ~n53121 & ~n53135;
  assign n53137 = ~n52518 & n53136;
  assign n53138 = pi207 & ~n52837;
  assign n53139 = ~pi207 & n52780;
  assign n53140 = pi208 & ~n53139;
  assign n53141 = ~n53138 & n53140;
  assign n53142 = ~pi208 & ~n52835;
  assign n53143 = ~pi200 & pi207;
  assign n53144 = ~n65386 & n53143;
  assign n53145 = n53142 & ~n53144;
  assign n53146 = ~pi1157 & ~n53145;
  assign n53147 = ~n53141 & n53146;
  assign n53148 = pi208 & pi1157;
  assign n53149 = ~n65345 & ~n52761;
  assign n53150 = ~pi207 & ~n53149;
  assign n53151 = ~n53138 & ~n53150;
  assign n53152 = n53148 & ~n53151;
  assign n53153 = ~n52835 & ~n65387;
  assign n53154 = n52737 & ~n53153;
  assign n53155 = ~n53152 & ~n53154;
  assign n53156 = ~n53147 & ~n53154;
  assign n53157 = ~n53152 & n53156;
  assign n53158 = ~n53147 & n53155;
  assign n53159 = n52527 & n65388;
  assign n53160 = ~pi207 & n52744;
  assign n53161 = ~n49607 & n52696;
  assign n53162 = pi207 & ~n53161;
  assign n53163 = ~n53160 & ~n53162;
  assign n53164 = pi208 & ~n53163;
  assign n53165 = ~pi208 & n49607;
  assign n53166 = ~n53115 & ~n53165;
  assign n53167 = ~n53164 & n53166;
  assign n53168 = ~pi1157 & ~n53167;
  assign n53169 = ~pi207 & ~n65347;
  assign n53170 = ~n53162 & ~n53169;
  assign n53171 = n53148 & ~n53170;
  assign n53172 = ~n49607 & ~n65387;
  assign n53173 = n52737 & ~n53172;
  assign n53174 = ~n53171 & ~n53173;
  assign n53175 = ~n53168 & n53174;
  assign n53176 = ~pi214 & ~n53175;
  assign n53177 = ~pi207 & ~n65349;
  assign n53178 = ~n52768 & n53177;
  assign n53179 = pi1157 & ~n53178;
  assign n53180 = pi1154 & ~n52779;
  assign n53181 = ~n65338 & ~n53180;
  assign n53182 = ~pi207 & ~n52742;
  assign n53183 = ~n53181 & n53182;
  assign n53184 = ~pi1157 & ~n53115;
  assign n53185 = ~n53183 & n53184;
  assign n53186 = ~n53179 & ~n53185;
  assign n53187 = pi207 & ~n52751;
  assign n53188 = pi208 & ~n53187;
  assign n53189 = ~n53186 & n53188;
  assign n53190 = n65387 & ~n53184;
  assign n53191 = ~pi208 & ~n52640;
  assign n53192 = ~n53190 & n53191;
  assign n53193 = pi214 & ~n53192;
  assign n53194 = ~n53189 & n53193;
  assign n53195 = pi212 & ~n53194;
  assign n53196 = ~n53176 & n53195;
  assign n53197 = ~n53159 & ~n53196;
  assign n53198 = ~pi211 & ~n53197;
  assign n53199 = ~n53137 & ~n53198;
  assign n53200 = pi219 & ~n53199;
  assign n53201 = ~pi214 & n53136;
  assign n53202 = ~pi212 & ~n53201;
  assign n53203 = ~pi299 & n53124;
  assign n53204 = n52766 & ~n53203;
  assign n53205 = pi207 & n65353;
  assign n53206 = pi207 & n52805;
  assign n53207 = ~n52801 & n53205;
  assign n53208 = n52806 & n53205;
  assign n53209 = ~n52750 & n65389;
  assign n53210 = ~pi207 & n65349;
  assign n53211 = pi208 & ~n53210;
  assign n53212 = ~n65390 & n53211;
  assign n53213 = ~n53204 & ~n53212;
  assign n53214 = pi1157 & ~n53213;
  assign n53215 = ~n53121 & ~n53214;
  assign n53216 = pi211 & n53215;
  assign n53217 = pi1158 & n65354;
  assign n53218 = ~pi1158 & n52696;
  assign n53219 = pi207 & ~n53218;
  assign n53220 = ~n53217 & n53219;
  assign n53221 = pi299 & ~pi1158;
  assign n53222 = n53177 & ~n53221;
  assign n53223 = ~n53220 & ~n53222;
  assign n53224 = n53148 & ~n53223;
  assign n53225 = ~pi299 & ~n52780;
  assign n53226 = ~pi207 & ~n53221;
  assign n53227 = ~n53225 & n53226;
  assign n53228 = pi208 & ~n53227;
  assign n53229 = ~n53220 & n53228;
  assign n53230 = pi207 & ~n39539;
  assign n53231 = ~pi299 & ~n53230;
  assign n53232 = pi1158 & ~n53231;
  assign n53233 = ~pi299 & n49613;
  assign n53234 = n49461 & n49596;
  assign n53235 = n49613 & n52548;
  assign n53236 = pi207 & n65391;
  assign n53237 = ~pi208 & ~n65392;
  assign n53238 = ~n53232 & n53237;
  assign n53239 = ~pi1157 & ~n53238;
  assign n53240 = ~n53229 & n53239;
  assign n53241 = pi1157 & ~n53108;
  assign n53242 = ~n65117 & n53241;
  assign n53243 = pi207 & ~n53242;
  assign n53244 = ~n53232 & ~n53243;
  assign n53245 = n52737 & ~n53244;
  assign n53246 = ~pi211 & ~n53245;
  assign n53247 = ~n53240 & n53246;
  assign n53248 = ~n53224 & n53246;
  assign n53249 = ~n53240 & n53248;
  assign n53250 = ~n53224 & n53247;
  assign n53251 = ~n53216 & ~n65393;
  assign n53252 = pi214 & ~n53251;
  assign n53253 = n53202 & ~n53252;
  assign n53254 = n39343 & ~n53175;
  assign n53255 = n52776 & ~n53215;
  assign n53256 = n52855 & ~n65388;
  assign n53257 = ~n53255 & ~n53256;
  assign n53258 = ~n53254 & ~n53256;
  assign n53259 = ~n53255 & n53258;
  assign n53260 = ~n53254 & n53257;
  assign n53261 = pi212 & ~n65394;
  assign n53262 = ~pi219 & ~n53261;
  assign n53263 = ~n53253 & n53262;
  assign n53264 = n62455 & ~n53263;
  assign n53265 = n62455 & ~n53200;
  assign n53266 = ~n53263 & n53265;
  assign n53267 = ~n53200 & n53264;
  assign n53268 = n53088 & ~n65395;
  assign n53269 = pi299 & ~pi1145;
  assign n53270 = ~n65132 & ~n53269;
  assign n53271 = pi1154 & ~n53270;
  assign n53272 = pi299 & pi1145;
  assign n53273 = n49622 & ~n53272;
  assign n53274 = ~pi1156 & ~n53273;
  assign n53275 = ~n53271 & n53274;
  assign n53276 = ~n65352 & ~n53269;
  assign n53277 = ~pi1154 & ~n53276;
  assign n53278 = n52894 & ~n53272;
  assign n53279 = pi1156 & ~n53278;
  assign n53280 = ~n53277 & n53279;
  assign n53281 = ~n53275 & ~n53280;
  assign n53282 = pi207 & ~n53281;
  assign n53283 = ~pi199 & n49582;
  assign n53284 = n53225 & ~n53283;
  assign n53285 = ~pi207 & ~n53269;
  assign n53286 = ~n53284 & n53285;
  assign n53287 = pi208 & ~n53286;
  assign n53288 = ~n53282 & n53287;
  assign n53289 = ~pi1157 & ~n65391;
  assign n53290 = ~pi1157 & ~n53108;
  assign n53291 = ~n65391 & n53290;
  assign n53292 = ~n53108 & n53289;
  assign n53293 = n53243 & ~n65396;
  assign n53294 = ~pi208 & ~n53272;
  assign n53295 = ~n53293 & n53294;
  assign n53296 = ~n53288 & ~n53295;
  assign n53297 = ~pi211 & ~n53296;
  assign n53298 = ~pi1157 & ~n53144;
  assign n53299 = ~pi208 & ~n53298;
  assign n53300 = n65387 & n53299;
  assign n53301 = n53130 & ~n53184;
  assign n53302 = ~pi208 & ~n65397;
  assign n53303 = ~n52920 & n53302;
  assign n53304 = pi207 & ~n52932;
  assign n53305 = ~pi207 & ~n52918;
  assign n53306 = ~n53284 & n53305;
  assign n53307 = pi208 & ~n53306;
  assign n53308 = ~n53304 & n53307;
  assign n53309 = ~n53303 & ~n53308;
  assign n53310 = pi211 & ~n53309;
  assign n53311 = ~n53297 & ~n53310;
  assign n53312 = ~pi214 & ~n53311;
  assign n53313 = ~n52881 & n53302;
  assign n53314 = pi207 & ~n52898;
  assign n53315 = ~pi207 & ~n52883;
  assign n53316 = ~n53284 & n53315;
  assign n53317 = pi208 & ~n53316;
  assign n53318 = ~n53314 & n53317;
  assign n53319 = ~n53313 & ~n53318;
  assign n53320 = pi211 & n53319;
  assign n53321 = ~pi211 & n53309;
  assign n53322 = pi214 & ~n53321;
  assign n53323 = pi214 & ~n53320;
  assign n53324 = ~n53321 & n53323;
  assign n53325 = ~n53320 & n53322;
  assign n53326 = pi212 & ~n65398;
  assign n53327 = ~n53312 & n53326;
  assign n53328 = pi214 & ~n53311;
  assign n53329 = n53202 & ~n53328;
  assign n53330 = ~pi219 & ~n53329;
  assign n53331 = ~pi219 & ~n53327;
  assign n53332 = ~n53329 & n53331;
  assign n53333 = ~n53327 & n53330;
  assign n53334 = n52518 & ~n53319;
  assign n53335 = ~n53137 & ~n53334;
  assign n53336 = pi219 & ~n53335;
  assign n53337 = n62455 & ~n53336;
  assign n53338 = ~n65399 & n53337;
  assign n53339 = pi213 & ~n53021;
  assign n53340 = ~n53338 & n53339;
  assign n53341 = ~pi209 & ~n53340;
  assign n53342 = ~n53268 & n53341;
  assign n53343 = ~n65385 & ~n53342;
  assign n53344 = pi230 & ~n53343;
  assign n53345 = ~pi230 & ~pi237;
  assign n53346 = ~n53344 & ~n53345;
  assign n53347 = n62455 & n49595;
  assign n53348 = ~pi1151 & n52465;
  assign n53349 = pi1150 & ~n53348;
  assign n53350 = ~n52462 & n53349;
  assign n53351 = ~pi1150 & pi1151;
  assign n53352 = ~n50528 & n53351;
  assign n53353 = ~pi1149 & ~n53352;
  assign n53354 = ~n53350 & n53353;
  assign n53355 = pi1149 & ~pi1150;
  assign n53356 = n52480 & n53355;
  assign n53357 = pi1151 & ~n52480;
  assign n53358 = pi1149 & n52476;
  assign n53359 = ~n53357 & n53358;
  assign n53360 = ~n53356 & ~n53359;
  assign n53361 = ~n53354 & n53360;
  assign n53362 = pi230 & ~n53361;
  assign n53363 = pi1149 & ~n53357;
  assign n53364 = n48938 & n53363;
  assign n53365 = pi1151 & ~n50528;
  assign n53366 = ~pi1149 & ~n53365;
  assign n53367 = ~pi1150 & ~n53366;
  assign n53368 = ~pi1151 & n48938;
  assign n53369 = pi1149 & ~n52480;
  assign n53370 = ~n53368 & n53369;
  assign n53371 = ~pi1149 & pi1151;
  assign n53372 = ~n50528 & n53371;
  assign n53373 = ~n53370 & ~n53372;
  assign n53374 = ~pi1150 & ~n53373;
  assign n53375 = ~n53364 & n53367;
  assign n53376 = ~pi1149 & n52462;
  assign n53377 = pi1150 & ~n53359;
  assign n53378 = ~n53376 & n53377;
  assign n53379 = pi1091 & ~n53378;
  assign n53380 = ~n53359 & ~n53376;
  assign n53381 = pi1150 & ~n53380;
  assign n53382 = ~pi1150 & ~n53372;
  assign n53383 = ~n53370 & n53382;
  assign n53384 = ~n53381 & ~n53383;
  assign n53385 = pi1091 & ~n53384;
  assign n53386 = ~n65400 & n53379;
  assign n53387 = ~n65014 & n50450;
  assign n53388 = n62455 & n49476;
  assign n53389 = ~n53387 & ~n53388;
  assign n53390 = ~pi1149 & pi1150;
  assign n53391 = ~pi1151 & n53390;
  assign n53392 = ~n53389 & n53391;
  assign n53393 = pi275 & ~n53392;
  assign n53394 = ~n65401 & n53393;
  assign n53395 = ~pi275 & pi1091;
  assign n53396 = n53361 & n53395;
  assign n53397 = ~n49535 & ~n53396;
  assign n53398 = ~n53394 & n53397;
  assign n53399 = ~pi1150 & ~n52394;
  assign n53400 = pi1150 & ~n52374;
  assign n53401 = ~pi1151 & ~n53400;
  assign n53402 = ~n53399 & n53401;
  assign n53403 = ~pi1150 & ~n52300;
  assign n53404 = pi1150 & ~n52309;
  assign n53405 = pi1151 & ~n53404;
  assign n53406 = ~n53403 & n53405;
  assign n53407 = ~n53402 & ~n53406;
  assign n53408 = ~n53403 & ~n53404;
  assign n53409 = pi1151 & ~n53408;
  assign n53410 = ~n53399 & ~n53400;
  assign n53411 = ~pi1151 & ~n53410;
  assign n53412 = pi275 & ~n53411;
  assign n53413 = ~n53409 & n53412;
  assign n53414 = pi275 & ~n53407;
  assign n53415 = pi1151 & ~n52320;
  assign n53416 = ~n52402 & ~n53415;
  assign n53417 = ~pi1150 & ~n53416;
  assign n53418 = ~pi1151 & ~n52404;
  assign n53419 = ~n52330 & ~n53418;
  assign n53420 = pi1150 & ~n53419;
  assign n53421 = ~pi275 & ~n53420;
  assign n53422 = ~n53417 & n53421;
  assign n53423 = pi1149 & ~n53422;
  assign n53424 = ~n65402 & n53423;
  assign n53425 = ~pi1150 & n52355;
  assign n53426 = pi1150 & n52349;
  assign n53427 = pi1151 & ~n53426;
  assign n53428 = ~n53425 & n53427;
  assign n53429 = pi1150 & ~n52382;
  assign n53430 = ~pi1150 & ~n52386;
  assign n53431 = ~pi1151 & ~n53430;
  assign n53432 = ~n53429 & n53431;
  assign n53433 = ~pi275 & ~n53432;
  assign n53434 = ~n53428 & n53433;
  assign n53435 = pi1150 & n52340;
  assign n53436 = ~pi1150 & n52344;
  assign n53437 = pi1151 & ~n53436;
  assign n53438 = ~n53435 & n53437;
  assign n53439 = pi1150 & n52371;
  assign n53440 = ~pi1150 & ~n52375;
  assign n53441 = ~pi1151 & ~n53440;
  assign n53442 = ~n53439 & n53441;
  assign n53443 = pi275 & ~n53442;
  assign n53444 = ~n53438 & n53443;
  assign n53445 = ~pi1149 & ~n53444;
  assign n53446 = ~n53434 & n53445;
  assign n53447 = n49535 & ~n53446;
  assign n53448 = ~n53424 & n53447;
  assign n53449 = ~n65401 & ~n53392;
  assign n53450 = pi275 & ~n53449;
  assign n53451 = pi1091 & n53361;
  assign n53452 = ~pi275 & ~n53451;
  assign n53453 = ~n49535 & ~n53452;
  assign n53454 = ~n53450 & n53453;
  assign n53455 = ~n53428 & ~n53432;
  assign n53456 = ~pi275 & ~n53455;
  assign n53457 = ~n53435 & ~n53436;
  assign n53458 = pi1151 & ~n53457;
  assign n53459 = ~n53439 & ~n53440;
  assign n53460 = ~pi1151 & ~n53459;
  assign n53461 = pi275 & ~n53460;
  assign n53462 = ~n53458 & n53461;
  assign n53463 = ~pi1149 & ~n53462;
  assign n53464 = ~n53456 & n53463;
  assign n53465 = pi1151 & ~n52300;
  assign n53466 = ~pi1150 & ~n52395;
  assign n53467 = ~n53465 & n53466;
  assign n53468 = ~pi1151 & ~n52374;
  assign n53469 = pi1150 & ~n53468;
  assign n53470 = ~n52310 & n53469;
  assign n53471 = pi275 & ~n53470;
  assign n53472 = ~n53467 & n53471;
  assign n53473 = ~pi1150 & ~n52320;
  assign n53474 = pi1150 & ~n52329;
  assign n53475 = pi1151 & ~n53474;
  assign n53476 = ~n53473 & n53475;
  assign n53477 = ~pi1150 & ~n52401;
  assign n53478 = pi1150 & ~n52404;
  assign n53479 = ~pi1151 & ~n53478;
  assign n53480 = ~n53477 & n53479;
  assign n53481 = ~pi275 & ~n53480;
  assign n53482 = ~n53476 & n53481;
  assign n53483 = pi1149 & ~n53482;
  assign n53484 = ~n53472 & n53483;
  assign n53485 = n49535 & ~n53484;
  assign n53486 = n49535 & ~n53464;
  assign n53487 = ~n53484 & n53486;
  assign n53488 = ~n53464 & n53485;
  assign n53489 = ~n53454 & ~n65403;
  assign n53490 = ~n53398 & ~n53448;
  assign n53491 = ~pi230 & n65404;
  assign n53492 = ~pi230 & ~n65404;
  assign n53493 = pi230 & n53361;
  assign n53494 = ~n53492 & ~n53493;
  assign n53495 = ~n53362 & ~n53491;
  assign n53496 = pi1150 & ~n52300;
  assign n53497 = ~pi1149 & ~n53399;
  assign n53498 = ~n53496 & n53497;
  assign n53499 = ~pi1150 & ~n52374;
  assign n53500 = pi1149 & ~n53499;
  assign n53501 = ~n53404 & n53500;
  assign n53502 = pi1150 & n52309;
  assign n53503 = ~pi1150 & n52374;
  assign n53504 = pi1149 & ~n53503;
  assign n53505 = ~n53502 & n53504;
  assign n53506 = pi1150 & n52300;
  assign n53507 = ~pi1150 & n52394;
  assign n53508 = ~pi1149 & ~n53507;
  assign n53509 = ~n53506 & n53508;
  assign n53510 = ~n53505 & ~n53509;
  assign n53511 = ~n53498 & ~n53501;
  assign n53512 = pi1148 & ~n65406;
  assign n53513 = ~pi1150 & n52371;
  assign n53514 = pi1149 & ~n53513;
  assign n53515 = ~n53435 & n53514;
  assign n53516 = pi1150 & n52344;
  assign n53517 = ~pi1149 & ~n53440;
  assign n53518 = ~n53516 & n53517;
  assign n53519 = ~n53515 & ~n53518;
  assign n53520 = ~pi1148 & ~n53519;
  assign n53521 = pi283 & ~n53520;
  assign n53522 = pi1148 & n65406;
  assign n53523 = ~pi1148 & ~n53518;
  assign n53524 = ~n53515 & n53523;
  assign n53525 = ~n53522 & ~n53524;
  assign n53526 = pi283 & ~n53525;
  assign n53527 = ~n53512 & n53521;
  assign n53528 = pi1091 & n65318;
  assign n53529 = pi1150 & ~n53528;
  assign n53530 = ~pi1150 & n53389;
  assign n53531 = ~pi1148 & pi1149;
  assign n53532 = ~n53530 & n53531;
  assign n53533 = ~n53529 & n53532;
  assign n53534 = ~pi1150 & n48938;
  assign n53535 = ~n52480 & ~n53534;
  assign n53536 = ~pi1149 & ~n53535;
  assign n53537 = pi1148 & ~n53536;
  assign n53538 = ~n52480 & ~n53355;
  assign n53539 = n52476 & ~n53538;
  assign n53540 = pi1148 & ~n53539;
  assign n53541 = ~n53536 & n53540;
  assign n53542 = ~n65317 & ~n52475;
  assign n53543 = ~n52475 & ~n52478;
  assign n53544 = ~n65317 & n53543;
  assign n53545 = ~n52478 & n53542;
  assign n53546 = pi1150 & ~n65409;
  assign n53547 = pi1149 & ~n53546;
  assign n53548 = n52476 & n53547;
  assign n53549 = n53537 & ~n53548;
  assign n53550 = n53537 & ~n53539;
  assign n53551 = pi1150 & ~n50528;
  assign n53552 = ~pi1149 & ~n53551;
  assign n53553 = ~pi1148 & ~n53552;
  assign n53554 = pi1091 & ~n53553;
  assign n53555 = ~n65408 & n53554;
  assign n53556 = ~n53533 & ~n53555;
  assign n53557 = pi1091 & n53552;
  assign n53558 = pi1149 & ~n53530;
  assign n53559 = ~n53529 & n53558;
  assign n53560 = ~pi1148 & ~n53559;
  assign n53561 = ~pi1148 & ~n53557;
  assign n53562 = ~n53559 & n53561;
  assign n53563 = ~n53557 & n53560;
  assign n53564 = ~n53536 & ~n53539;
  assign n53565 = pi1091 & ~n53564;
  assign n53566 = pi1148 & ~n53565;
  assign n53567 = ~pi283 & ~n53566;
  assign n53568 = ~n65410 & n53567;
  assign n53569 = ~pi283 & ~n65410;
  assign n53570 = ~n53566 & n53569;
  assign n53571 = ~pi283 & ~n53556;
  assign n53572 = pi272 & ~n65411;
  assign n53573 = ~n65407 & n53572;
  assign n53574 = ~pi1150 & ~n52382;
  assign n53575 = pi1149 & ~n53426;
  assign n53576 = ~n53574 & n53575;
  assign n53577 = pi1150 & n52355;
  assign n53578 = ~pi1149 & ~n53430;
  assign n53579 = ~n53577 & n53578;
  assign n53580 = ~n53576 & ~n53579;
  assign n53581 = ~pi1148 & ~n53580;
  assign n53582 = pi1150 & ~n52320;
  assign n53583 = ~pi1149 & ~n53477;
  assign n53584 = ~n53582 & n53583;
  assign n53585 = ~pi1150 & ~n52404;
  assign n53586 = pi1149 & ~n53585;
  assign n53587 = ~n53474 & n53586;
  assign n53588 = pi1148 & ~n53587;
  assign n53589 = ~n53584 & n53588;
  assign n53590 = pi283 & ~n53589;
  assign n53591 = ~n53584 & ~n53587;
  assign n53592 = pi1148 & ~n53591;
  assign n53593 = ~pi1148 & ~n53579;
  assign n53594 = ~n53576 & n53593;
  assign n53595 = ~n53592 & ~n53594;
  assign n53596 = pi283 & ~n53595;
  assign n53597 = ~n53581 & n53590;
  assign n53598 = pi1091 & n65408;
  assign n53599 = pi1150 & ~n65318;
  assign n53600 = ~pi1150 & ~n52465;
  assign n53601 = pi1149 & ~n53600;
  assign n53602 = pi1149 & n65318;
  assign n53603 = ~n53547 & ~n53602;
  assign n53604 = ~n53600 & ~n53603;
  assign n53605 = ~n53599 & n53601;
  assign n53606 = pi1091 & ~n65413;
  assign n53607 = pi1091 & n53553;
  assign n53608 = ~n65413 & n53607;
  assign n53609 = n53553 & n53606;
  assign n53610 = ~pi283 & ~n65414;
  assign n53611 = ~n53598 & n53610;
  assign n53612 = ~pi272 & ~n53611;
  assign n53613 = ~n65412 & n53612;
  assign n53614 = ~pi230 & ~n53613;
  assign n53615 = ~pi230 & ~n53573;
  assign n53616 = ~n53613 & n53615;
  assign n53617 = ~n53573 & n53614;
  assign n53618 = n53553 & ~n65413;
  assign n53619 = pi230 & ~n65408;
  assign n53620 = ~n53618 & n53619;
  assign po429 = ~n65415 & ~n53620;
  assign n53622 = pi1147 & n52320;
  assign n53623 = ~pi1147 & n52355;
  assign n53624 = pi1149 & ~n53623;
  assign n53625 = ~n53622 & n53624;
  assign n53626 = pi1147 & n52401;
  assign n53627 = ~pi1147 & ~n52386;
  assign n53628 = ~pi1149 & ~n53627;
  assign n53629 = ~n53626 & n53628;
  assign n53630 = ~pi1148 & ~n53629;
  assign n53631 = ~n53625 & n53630;
  assign n53632 = ~pi1147 & ~n52382;
  assign n53633 = pi1147 & n52404;
  assign n53634 = ~pi1149 & ~n53633;
  assign n53635 = ~n53632 & n53634;
  assign n53636 = ~pi1147 & n52349;
  assign n53637 = pi1147 & n52329;
  assign n53638 = pi1149 & ~n53637;
  assign n53639 = ~n53636 & n53638;
  assign n53640 = pi1148 & ~n53639;
  assign n53641 = ~n53635 & n53640;
  assign n53642 = ~pi283 & ~n53641;
  assign n53643 = ~pi283 & ~n53631;
  assign n53644 = ~n53641 & n53643;
  assign n53645 = ~n53631 & n53642;
  assign n53646 = pi1147 & n52300;
  assign n53647 = ~pi1147 & n52344;
  assign n53648 = ~pi1148 & ~n53647;
  assign n53649 = ~n53646 & n53648;
  assign n53650 = ~pi1147 & n52340;
  assign n53651 = pi1147 & n52309;
  assign n53652 = pi1148 & ~n53651;
  assign n53653 = ~n53650 & n53652;
  assign n53654 = pi1149 & ~n53653;
  assign n53655 = ~n53649 & n53654;
  assign n53656 = pi1147 & n52394;
  assign n53657 = ~pi1147 & ~n52375;
  assign n53658 = ~pi1148 & ~n53657;
  assign n53659 = ~n53656 & n53658;
  assign n53660 = ~pi1147 & n52371;
  assign n53661 = pi1147 & n52374;
  assign n53662 = pi1148 & ~n53661;
  assign n53663 = ~n53660 & n53662;
  assign n53664 = ~pi1149 & ~n53663;
  assign n53665 = ~n53659 & n53664;
  assign n53666 = pi283 & ~n53665;
  assign n53667 = ~n53655 & n53666;
  assign n53668 = ~pi230 & ~n53667;
  assign n53669 = ~n53649 & ~n53653;
  assign n53670 = pi283 & ~n53669;
  assign n53671 = ~pi1148 & ~n53623;
  assign n53672 = ~n53622 & n53671;
  assign n53673 = pi1148 & ~n53637;
  assign n53674 = ~n53636 & n53673;
  assign n53675 = ~n53672 & ~n53674;
  assign n53676 = ~pi283 & ~n53675;
  assign n53677 = pi1149 & ~n53676;
  assign n53678 = ~n53670 & n53677;
  assign n53679 = ~pi1148 & ~n53627;
  assign n53680 = ~n53626 & n53679;
  assign n53681 = pi1148 & ~n53633;
  assign n53682 = ~n53632 & n53681;
  assign n53683 = ~n53680 & ~n53682;
  assign n53684 = ~pi283 & ~n53683;
  assign n53685 = pi1147 & ~n52394;
  assign n53686 = ~pi1147 & n52375;
  assign n53687 = ~pi1148 & ~n53686;
  assign n53688 = ~n53685 & n53687;
  assign n53689 = ~pi1147 & ~n52371;
  assign n53690 = pi1147 & ~n52374;
  assign n53691 = pi1148 & ~n53690;
  assign n53692 = ~n53689 & n53691;
  assign n53693 = pi283 & ~n53692;
  assign n53694 = ~n53688 & n53693;
  assign n53695 = ~pi1149 & ~n53694;
  assign n53696 = ~n53684 & n53695;
  assign n53697 = ~n53635 & ~n53639;
  assign n53698 = pi1148 & ~n53697;
  assign n53699 = ~n53625 & ~n53629;
  assign n53700 = ~pi1148 & ~n53699;
  assign n53701 = ~pi283 & ~n53700;
  assign n53702 = ~n53698 & n53701;
  assign n53703 = pi1147 & ~n52300;
  assign n53704 = ~pi1147 & ~n52344;
  assign n53705 = ~pi1148 & ~n53704;
  assign n53706 = ~n53703 & n53705;
  assign n53707 = ~pi1147 & ~n52340;
  assign n53708 = pi1147 & ~n52309;
  assign n53709 = pi1148 & ~n53708;
  assign n53710 = ~n53707 & n53709;
  assign n53711 = pi1149 & ~n53710;
  assign n53712 = ~n53706 & n53711;
  assign n53713 = ~pi1149 & ~n53692;
  assign n53714 = ~n53688 & n53713;
  assign n53715 = pi283 & ~n53714;
  assign n53716 = ~n53712 & n53715;
  assign n53717 = ~n53702 & ~n53716;
  assign n53718 = ~n53678 & ~n53696;
  assign n53719 = ~pi230 & ~n65417;
  assign n53720 = ~pi230 & ~n65416;
  assign n53721 = ~n53667 & n53720;
  assign n53722 = ~n65416 & n53668;
  assign n53723 = pi1147 & ~n48938;
  assign n53724 = n53602 & ~n53723;
  assign n53725 = pi1147 & ~n52476;
  assign n53726 = ~pi1149 & n52465;
  assign n53727 = ~n53725 & n53726;
  assign n53728 = pi1148 & ~n53727;
  assign n53729 = pi1148 & ~n53724;
  assign n53730 = ~n53727 & n53729;
  assign n53731 = ~n53724 & n53728;
  assign n53732 = pi1149 & ~n50528;
  assign n53733 = ~n53723 & ~n53732;
  assign n53734 = ~pi1148 & ~n53733;
  assign n53735 = pi230 & ~n53734;
  assign n53736 = ~n65419 & n53735;
  assign po440 = ~n65418 & ~n53736;
  assign n53738 = ~pi230 & pi234;
  assign n53739 = ~n52835 & ~n53138;
  assign n53740 = ~pi208 & ~n53739;
  assign n53741 = ~pi1154 & ~n65339;
  assign n53742 = ~pi199 & n52662;
  assign n53743 = ~n65108 & n49595;
  assign n53744 = ~n53741 & n53743;
  assign n53745 = pi207 & n53744;
  assign n53746 = n65359 & ~n53745;
  assign n53747 = pi208 & ~n53746;
  assign n53748 = ~n53740 & ~n53747;
  assign n53749 = ~pi211 & ~n53748;
  assign n53750 = n52738 & ~n53161;
  assign n53751 = pi207 & ~n49607;
  assign n53752 = ~n53744 & n53751;
  assign n53753 = pi208 & ~n53752;
  assign n53754 = n52724 & ~n53752;
  assign n53755 = ~n52723 & n53753;
  assign n53756 = ~n53750 & ~n65420;
  assign n53757 = pi211 & ~n53756;
  assign n53758 = ~n53749 & ~n53757;
  assign n53759 = ~pi214 & n53758;
  assign n53760 = ~pi207 & n52640;
  assign n53761 = ~n53187 & ~n53760;
  assign n53762 = ~pi208 & ~n53761;
  assign n53763 = ~pi299 & ~n49447;
  assign n53764 = ~n53741 & ~n53763;
  assign n53765 = pi207 & n53764;
  assign n53766 = ~n52752 & ~n53765;
  assign n53767 = pi208 & ~n53766;
  assign n53768 = ~n53762 & ~n53767;
  assign n53769 = pi211 & ~n53768;
  assign n53770 = ~pi211 & ~n53756;
  assign n53771 = pi214 & ~n53770;
  assign n53772 = ~n53769 & n53771;
  assign n53773 = pi212 & ~n53772;
  assign n53774 = ~n53759 & n53773;
  assign n53775 = ~n38985 & n52696;
  assign n53776 = ~n53032 & ~n53745;
  assign n53777 = ~n53775 & ~n53776;
  assign n53778 = ~pi214 & ~n53777;
  assign n53779 = ~pi212 & ~n53778;
  assign n53780 = pi214 & n53758;
  assign n53781 = n53779 & ~n53780;
  assign n53782 = ~pi219 & ~n53781;
  assign n53783 = ~pi219 & ~n53774;
  assign n53784 = ~n53781 & n53783;
  assign n53785 = ~n53774 & n53782;
  assign n53786 = ~n52518 & n53777;
  assign n53787 = pi219 & ~n53786;
  assign n53788 = ~pi211 & ~n53768;
  assign n53789 = ~n52517 & n53788;
  assign n53790 = n53787 & ~n53789;
  assign n53791 = n37948 & ~n53790;
  assign n53792 = ~n65421 & n53791;
  assign n53793 = pi1153 & ~n52776;
  assign n53794 = ~n52628 & ~n52631;
  assign n53795 = ~n53793 & ~n53794;
  assign n53796 = pi212 & ~n53795;
  assign n53797 = ~n49653 & ~n50251;
  assign n53798 = n52527 & ~n53797;
  assign n53799 = ~pi219 & ~n53798;
  assign n53800 = ~n53796 & n53799;
  assign n53801 = n52520 & ~n53800;
  assign n53802 = pi1152 & ~n53801;
  assign n53803 = n52766 & ~n65390;
  assign n53804 = n52548 & ~n53764;
  assign n53805 = pi208 & ~n53804;
  assign n53806 = ~n52825 & n53805;
  assign n53807 = ~n53803 & ~n53806;
  assign n53808 = ~n52786 & ~n53807;
  assign n53809 = pi211 & n53808;
  assign n53810 = ~n53788 & ~n53809;
  assign n53811 = pi214 & n53810;
  assign n53812 = n53779 & ~n53811;
  assign n53813 = ~pi219 & ~n53812;
  assign n53814 = ~pi214 & ~n53810;
  assign n53815 = ~pi211 & ~pi1153;
  assign n53816 = pi299 & n53815;
  assign n53817 = ~pi211 & n52786;
  assign n53818 = pi214 & ~n65422;
  assign n53819 = ~pi211 & ~n53808;
  assign n53820 = pi214 & ~n53819;
  assign n53821 = ~n53807 & n53820;
  assign n53822 = ~n53807 & n53818;
  assign n53823 = ~n53814 & ~n65423;
  assign n53824 = pi212 & ~n53823;
  assign n53825 = n53813 & ~n53824;
  assign n53826 = n52518 & ~n53807;
  assign n53827 = n53787 & ~n53826;
  assign n53828 = n62455 & ~n53827;
  assign n53829 = ~n53825 & n53828;
  assign n53830 = n53802 & ~n53829;
  assign n53831 = ~n39342 & n53797;
  assign n53832 = n52967 & ~n53831;
  assign n53833 = ~n52632 & n53832;
  assign n53834 = ~n62455 & n53833;
  assign n53835 = ~pi1152 & ~n53834;
  assign n53836 = pi211 & ~n53777;
  assign n53837 = pi214 & ~n53836;
  assign n53838 = n53820 & ~n53836;
  assign n53839 = ~n53819 & n53837;
  assign n53840 = ~n53814 & ~n65424;
  assign n53841 = pi212 & ~n53840;
  assign n53842 = n53813 & ~n53841;
  assign n53843 = pi219 & ~n53777;
  assign n53844 = n62455 & ~n53843;
  assign n53845 = ~n53842 & n53844;
  assign n53846 = n53835 & ~n53845;
  assign n53847 = ~pi213 & ~n53846;
  assign n53848 = ~pi213 & ~n53830;
  assign n53849 = ~n53846 & n53848;
  assign n53850 = ~n53830 & n53847;
  assign n53851 = ~n53792 & ~n65425;
  assign n53852 = pi209 & ~n53851;
  assign n53853 = ~n50242 & ~n50266;
  assign n53854 = n49519 & ~n53853;
  assign n53855 = n52766 & ~n53854;
  assign n53856 = ~pi207 & n53854;
  assign n53857 = ~n49457 & n50085;
  assign n53858 = pi207 & n53857;
  assign n53859 = pi208 & ~n53858;
  assign n53860 = ~n53856 & n53859;
  assign n53861 = ~n53855 & ~n53860;
  assign n53862 = ~pi211 & ~n53861;
  assign n53863 = ~pi1153 & ~n48497;
  assign n53864 = n52671 & ~n53863;
  assign n53865 = ~n50244 & ~n53864;
  assign n53866 = ~n38985 & n53865;
  assign n53867 = n38985 & ~n50056;
  assign n53868 = ~n53031 & ~n53867;
  assign n53869 = ~n53866 & n53868;
  assign n53870 = pi211 & n53869;
  assign n53871 = ~pi211 & n53861;
  assign n53872 = pi211 & ~n53869;
  assign n53873 = ~n53871 & ~n53872;
  assign n53874 = ~n53862 & ~n53870;
  assign n53875 = ~n52517 & n65426;
  assign n53876 = pi219 & ~n53869;
  assign n53877 = ~n53038 & ~n53876;
  assign n53878 = ~n53875 & ~n53877;
  assign n53879 = n62455 & ~n53878;
  assign n53880 = ~pi214 & ~n53869;
  assign n53881 = ~pi212 & ~n53880;
  assign n53882 = pi207 & ~n53865;
  assign n53883 = ~n52640 & ~n53882;
  assign n53884 = ~pi208 & ~n53883;
  assign n53885 = pi207 & ~n53857;
  assign n53886 = ~n52768 & n53885;
  assign n53887 = ~n49593 & ~n53864;
  assign n53888 = ~n50244 & n53887;
  assign n53889 = ~pi207 & ~n53888;
  assign n53890 = ~n53886 & ~n53889;
  assign n53891 = pi208 & ~n53890;
  assign n53892 = ~n53884 & ~n53891;
  assign n53893 = ~pi211 & ~n53892;
  assign n53894 = ~pi207 & n52642;
  assign n53895 = pi1154 & ~n48570;
  assign n53896 = ~n50233 & n53895;
  assign n53897 = ~n50234 & ~n53896;
  assign n53898 = pi207 & ~n53897;
  assign n53899 = ~n53894 & ~n53898;
  assign n53900 = ~pi208 & ~n53899;
  assign n53901 = ~pi207 & ~n53897;
  assign n53902 = pi207 & ~n49452;
  assign n53903 = ~n50076 & n53902;
  assign n53904 = ~n53901 & ~n53903;
  assign n53905 = pi208 & ~n53904;
  assign n53906 = ~n53900 & ~n53905;
  assign n53907 = pi211 & ~n53906;
  assign n53908 = ~n53893 & ~n53907;
  assign n53909 = pi214 & n53908;
  assign n53910 = n53881 & ~n53909;
  assign n53911 = ~pi214 & n53908;
  assign n53912 = pi211 & ~n53861;
  assign n53913 = ~pi211 & ~n53906;
  assign n53914 = pi214 & ~n53913;
  assign n53915 = pi214 & ~n53912;
  assign n53916 = ~n53913 & n53915;
  assign n53917 = ~n53912 & n53914;
  assign n53918 = pi212 & ~n65427;
  assign n53919 = ~n53911 & n53918;
  assign n53920 = ~pi219 & ~n53919;
  assign n53921 = ~pi219 & ~n53910;
  assign n53922 = ~n53919 & n53921;
  assign n53923 = ~n53910 & n53920;
  assign n53924 = n53879 & ~n65428;
  assign n53925 = n53802 & ~n53924;
  assign n53926 = ~n50232 & ~n53896;
  assign n53927 = pi207 & ~n53926;
  assign n53928 = ~n53894 & ~n53927;
  assign n53929 = ~pi208 & ~n53928;
  assign n53930 = ~pi207 & ~n53926;
  assign n53931 = pi1153 & n53230;
  assign n53932 = ~n53930 & ~n53931;
  assign n53933 = pi208 & ~n53932;
  assign n53934 = ~n65362 & ~n53933;
  assign n53935 = ~n53929 & n53934;
  assign n53936 = ~n50076 & ~n50343;
  assign n53937 = pi1154 & ~n53936;
  assign n53938 = ~n50241 & ~n53937;
  assign n53939 = pi207 & ~n53938;
  assign n53940 = ~n53760 & ~n53939;
  assign n53941 = ~pi208 & ~n53940;
  assign n53942 = ~pi207 & n53938;
  assign n53943 = ~pi299 & ~pi1153;
  assign n53944 = ~n39539 & ~n53943;
  assign n53945 = ~n52768 & n53944;
  assign n53946 = pi207 & ~n53945;
  assign n53947 = pi208 & ~n53946;
  assign n53948 = ~n53942 & n53947;
  assign n53949 = ~n53941 & ~n53948;
  assign n53950 = n65364 & n53949;
  assign n53951 = ~n53929 & ~n53933;
  assign n53952 = n52909 & n53951;
  assign n53953 = ~pi211 & n53949;
  assign n53954 = pi211 & n53951;
  assign n53955 = ~n53953 & ~n53954;
  assign n53956 = ~n65324 & ~n53955;
  assign n53957 = ~n53952 & ~n53956;
  assign n53958 = ~n53935 & ~n53950;
  assign n53959 = ~pi219 & ~n65429;
  assign n53960 = pi1154 & ~n50260;
  assign n53961 = ~n50242 & ~n53960;
  assign n53962 = n53032 & n53961;
  assign n53963 = n50091 & n53026;
  assign n53964 = ~n53962 & ~n53963;
  assign n53965 = n39346 & ~n52517;
  assign n53966 = ~n64625 & n52967;
  assign n53967 = n53964 & ~n65430;
  assign n53968 = pi219 & n53964;
  assign n53969 = n62455 & ~n53968;
  assign n53970 = n65324 & ~n52628;
  assign n53971 = n53964 & n53970;
  assign n53972 = n53969 & ~n53971;
  assign n53973 = n62455 & ~n53967;
  assign n53974 = ~n53959 & n65431;
  assign n53975 = n53835 & ~n53974;
  assign n53976 = ~n53925 & ~n53975;
  assign n53977 = ~pi213 & ~n53976;
  assign n53978 = ~n52518 & n53869;
  assign n53979 = ~n52517 & n53893;
  assign n53980 = ~n53978 & ~n53979;
  assign n53981 = pi219 & ~n53980;
  assign n53982 = pi211 & ~n53892;
  assign n53983 = n52738 & ~n53854;
  assign n53984 = ~n53860 & ~n53983;
  assign n53985 = ~pi1154 & n39538;
  assign n53986 = n65120 & n52765;
  assign n53987 = ~n52802 & ~n53986;
  assign n53988 = ~n53984 & n53987;
  assign n53989 = ~pi211 & n53988;
  assign n53990 = n39342 & ~n53989;
  assign n53991 = ~n53982 & n53990;
  assign n53992 = pi211 & n53988;
  assign n53993 = ~n52835 & n53865;
  assign n53994 = ~pi207 & ~n53993;
  assign n53995 = pi299 & ~pi1156;
  assign n53996 = n53885 & ~n53995;
  assign n53997 = pi208 & ~n53996;
  assign n53998 = ~n53994 & n53997;
  assign n53999 = n53142 & ~n53882;
  assign n54000 = ~pi211 & ~n53999;
  assign n54001 = ~n53998 & n54000;
  assign n54002 = ~n65324 & ~n54001;
  assign n54003 = ~n53992 & n54002;
  assign n54004 = ~pi212 & n53880;
  assign n54005 = ~pi219 & ~n54004;
  assign n54006 = ~n54003 & n54005;
  assign n54007 = ~n53991 & n54006;
  assign n54008 = ~n53981 & ~n54007;
  assign n54009 = n50550 & ~n54008;
  assign n54010 = ~pi1152 & n62455;
  assign n54011 = n64625 & ~n53949;
  assign n54012 = ~pi211 & ~n52835;
  assign n54013 = n53964 & n54012;
  assign n54014 = ~n65324 & ~n54013;
  assign n54015 = ~pi211 & n54014;
  assign n54016 = ~n52909 & ~n54014;
  assign n54017 = ~pi299 & ~n65156;
  assign n54018 = ~pi1154 & ~n54017;
  assign n54019 = ~n52802 & n54018;
  assign n54020 = ~n50209 & n53937;
  assign n54021 = ~n54019 & ~n54020;
  assign n54022 = pi207 & n54021;
  assign n54023 = n52738 & ~n54022;
  assign n54024 = ~pi207 & n54021;
  assign n54025 = ~n52802 & n53944;
  assign n54026 = pi207 & ~n54025;
  assign n54027 = pi208 & ~n54026;
  assign n54028 = ~n54024 & n54027;
  assign n54029 = ~n54023 & ~n54028;
  assign n54030 = ~n54016 & ~n54029;
  assign n54031 = ~n54015 & ~n54030;
  assign n54032 = ~pi211 & n54029;
  assign n54033 = pi211 & n53949;
  assign n54034 = n39342 & ~n54033;
  assign n54035 = n39342 & ~n54032;
  assign n54036 = ~n54033 & n54035;
  assign n54037 = ~n54032 & n54034;
  assign n54038 = pi211 & n54029;
  assign n54039 = n54014 & ~n54038;
  assign n54040 = ~n65432 & ~n54039;
  assign n54041 = ~n54011 & n54031;
  assign n54042 = ~pi219 & ~n65433;
  assign n54043 = n52517 & ~n53964;
  assign n54044 = pi211 & n53964;
  assign n54045 = n53038 & ~n54044;
  assign n54046 = ~n53953 & n54045;
  assign n54047 = ~n54043 & ~n54046;
  assign n54048 = ~n54042 & n54047;
  assign n54049 = n54010 & ~n54048;
  assign n54050 = pi213 & ~n54049;
  assign n54051 = ~n54009 & n54050;
  assign n54052 = ~pi209 & ~n54051;
  assign n54053 = ~n53977 & n54052;
  assign n54054 = ~pi212 & n53056;
  assign n54055 = n52527 & ~n52607;
  assign n54056 = ~pi219 & ~n65434;
  assign n54057 = ~n65332 & n54056;
  assign n54058 = pi213 & ~n50250;
  assign n54059 = n52520 & n54058;
  assign n54060 = ~n54057 & n54059;
  assign n54061 = ~n54053 & ~n54060;
  assign n54062 = pi209 & ~n53792;
  assign n54063 = ~n65425 & n54062;
  assign n54064 = ~pi213 & n53976;
  assign n54065 = ~n54009 & ~n54049;
  assign n54066 = pi213 & ~n54065;
  assign n54067 = ~pi209 & ~n54066;
  assign n54068 = ~n54064 & n54067;
  assign n54069 = ~n54063 & ~n54068;
  assign n54070 = ~n54060 & ~n54069;
  assign n54071 = ~n53852 & n54061;
  assign n54072 = pi230 & ~n65435;
  assign n54073 = ~n53738 & ~n54072;
  assign n54074 = ~pi230 & ~pi235;
  assign n54075 = ~pi1156 & n65119;
  assign n54076 = ~n52801 & ~n54075;
  assign n54077 = pi207 & ~n54076;
  assign n54078 = ~n53139 & ~n54077;
  assign n54079 = pi208 & ~n54078;
  assign n54080 = ~n52845 & ~n54079;
  assign n54081 = ~pi1157 & ~n54080;
  assign n54082 = ~n53150 & ~n54077;
  assign n54083 = n53148 & ~n54082;
  assign n54084 = ~n52847 & ~n54083;
  assign n54085 = ~n54081 & n54084;
  assign n54086 = pi211 & ~n54085;
  assign n54087 = ~n65389 & n53211;
  assign n54088 = ~n52767 & ~n54087;
  assign n54089 = pi1157 & n54088;
  assign n54090 = n52785 & ~n54087;
  assign n54091 = n38985 & ~n65342;
  assign n54092 = ~n54075 & n54091;
  assign n54093 = ~n53117 & ~n54092;
  assign n54094 = ~n52667 & n54093;
  assign n54095 = ~pi1157 & ~n54094;
  assign n54096 = ~pi211 & ~n54095;
  assign n54097 = ~n65436 & n54096;
  assign n54098 = ~n65324 & ~n54097;
  assign n54099 = ~n54086 & n54098;
  assign n54100 = ~pi211 & ~n54085;
  assign n54101 = ~n49801 & ~n65342;
  assign n54102 = pi207 & ~n54101;
  assign n54103 = ~n53160 & ~n54102;
  assign n54104 = pi208 & ~n54103;
  assign n54105 = ~n52745 & ~n54104;
  assign n54106 = ~pi1157 & ~n54105;
  assign n54107 = ~n53169 & ~n54102;
  assign n54108 = n53148 & ~n54107;
  assign n54109 = ~n52741 & ~n54108;
  assign n54110 = ~n54106 & n54109;
  assign n54111 = pi211 & ~n54110;
  assign n54112 = n39342 & ~n54111;
  assign n54113 = n39342 & ~n54100;
  assign n54114 = ~n54111 & n54113;
  assign n54115 = ~n54100 & n54112;
  assign n54116 = ~n53131 & ~n54092;
  assign n54117 = ~n52714 & n54116;
  assign n54118 = pi1157 & ~n54117;
  assign n54119 = ~n54095 & ~n54118;
  assign n54120 = n52517 & ~n54119;
  assign n54121 = ~n65437 & ~n54120;
  assign n54122 = ~n54099 & ~n54120;
  assign n54123 = ~n65437 & n54122;
  assign n54124 = ~n54099 & n54121;
  assign n54125 = ~pi219 & ~n65438;
  assign n54126 = ~pi211 & n54110;
  assign n54127 = pi211 & ~n54119;
  assign n54128 = ~n65324 & ~n54127;
  assign n54129 = ~n54126 & n54128;
  assign n54130 = n65324 & n54119;
  assign n54131 = pi219 & ~n54130;
  assign n54132 = ~n54129 & n54131;
  assign n54133 = pi209 & ~n54132;
  assign n54134 = ~n54125 & n54133;
  assign n54135 = n38985 & ~n53961;
  assign n54136 = n65341 & ~n53031;
  assign n54137 = ~n38985 & ~n54136;
  assign n54138 = ~n54135 & ~n54137;
  assign n54139 = ~pi1157 & n54138;
  assign n54140 = n52766 & ~n52824;
  assign n54141 = n52765 & n52797;
  assign n54142 = ~n53937 & ~n54018;
  assign n54143 = pi207 & n54142;
  assign n54144 = pi208 & ~n54143;
  assign n54145 = pi208 & ~n54141;
  assign n54146 = ~n54143 & n54145;
  assign n54147 = ~n54141 & n54144;
  assign n54148 = ~n54140 & ~n65439;
  assign n54149 = pi1157 & ~n54148;
  assign n54150 = ~pi211 & ~n54149;
  assign n54151 = ~pi211 & ~n54139;
  assign n54152 = ~n54149 & n54151;
  assign n54153 = ~n54139 & n54150;
  assign n54154 = ~n52835 & ~n54138;
  assign n54155 = pi211 & n54154;
  assign n54156 = ~n65440 & ~n54155;
  assign n54157 = ~n65324 & ~n54156;
  assign n54158 = n52517 & ~n54138;
  assign n54159 = ~n52686 & n52738;
  assign n54160 = ~pi207 & n52686;
  assign n54161 = pi208 & ~n54022;
  assign n54162 = ~n54160 & n54161;
  assign n54163 = ~n54159 & ~n54162;
  assign n54164 = pi211 & ~n54163;
  assign n54165 = ~pi211 & ~n54154;
  assign n54166 = n39342 & ~n54165;
  assign n54167 = n39342 & ~n54164;
  assign n54168 = ~n54165 & n54167;
  assign n54169 = ~n54164 & n54166;
  assign n54170 = ~n54158 & ~n65441;
  assign n54171 = ~n54157 & n54170;
  assign n54172 = ~pi219 & ~n54171;
  assign n54173 = ~pi211 & n54163;
  assign n54174 = pi211 & ~n54138;
  assign n54175 = ~n65324 & ~n54174;
  assign n54176 = ~n54173 & n54175;
  assign n54177 = n65324 & n54138;
  assign n54178 = pi219 & ~n54177;
  assign n54179 = ~n54176 & n54178;
  assign n54180 = ~pi209 & ~n54179;
  assign n54181 = ~n54172 & n54180;
  assign n54182 = ~n54134 & ~n54181;
  assign n54183 = n62455 & ~n54182;
  assign n54184 = ~n65333 & n53065;
  assign n54185 = n52621 & ~n65377;
  assign n54186 = pi219 & n65324;
  assign n54187 = ~n62455 & ~n50175;
  assign n54188 = ~n50175 & ~n54186;
  assign n54189 = ~n62455 & n54188;
  assign n54190 = ~n54186 & n54187;
  assign n54191 = ~n65442 & n65443;
  assign n54192 = pi213 & ~n54191;
  assign n54193 = ~n54183 & n54192;
  assign n54194 = ~pi299 & ~pi1157;
  assign n54195 = ~n54081 & n54194;
  assign n54196 = n54080 & n54194;
  assign n54197 = ~n52786 & ~n65436;
  assign n54198 = pi1157 & ~n54088;
  assign n54199 = pi299 & ~pi1157;
  assign n54200 = ~n54081 & ~n54199;
  assign n54201 = ~n54198 & n54200;
  assign n54202 = ~n52786 & ~n54201;
  assign n54203 = ~n65444 & n54197;
  assign n54204 = ~pi211 & ~n65445;
  assign n54205 = n54128 & ~n54204;
  assign n54206 = n54131 & ~n54205;
  assign n54207 = pi211 & n65445;
  assign n54208 = ~n49622 & ~n65353;
  assign n54209 = ~n65342 & ~n54208;
  assign n54210 = pi207 & ~n54209;
  assign n54211 = ~n53183 & ~n54210;
  assign n54212 = pi208 & ~n54211;
  assign n54213 = ~n52772 & ~n54212;
  assign n54214 = ~pi1157 & ~n54213;
  assign n54215 = n52769 & ~n54088;
  assign n54216 = ~n54214 & ~n54215;
  assign n54217 = ~pi211 & ~n54216;
  assign n54218 = n39342 & ~n54217;
  assign n54219 = ~n54207 & n54218;
  assign n54220 = pi211 & n54216;
  assign n54221 = ~n54126 & ~n54220;
  assign n54222 = ~n65324 & ~n54221;
  assign n54223 = ~n54120 & ~n54222;
  assign n54224 = ~n54219 & n54223;
  assign n54225 = ~pi219 & ~n54224;
  assign n54226 = ~n54206 & ~n54225;
  assign n54227 = pi209 & ~n54226;
  assign n54228 = ~n52798 & ~n53894;
  assign n54229 = ~pi208 & ~n54228;
  assign n54230 = ~pi207 & ~n52797;
  assign n54231 = ~n53927 & ~n54230;
  assign n54232 = pi208 & ~n54231;
  assign n54233 = ~n54229 & ~n54232;
  assign n54234 = ~pi211 & n54233;
  assign n54235 = n54175 & ~n54234;
  assign n54236 = n54178 & ~n54235;
  assign n54237 = ~n52756 & ~n53760;
  assign n54238 = ~pi208 & ~n54237;
  assign n54239 = ~pi207 & ~n52755;
  assign n54240 = ~n53939 & ~n54239;
  assign n54241 = pi208 & ~n54240;
  assign n54242 = ~n65362 & ~n54241;
  assign n54243 = ~n54238 & n54242;
  assign n54244 = n65364 & n54163;
  assign n54245 = n64625 & n54233;
  assign n54246 = ~n54158 & ~n54245;
  assign n54247 = ~n54244 & n54246;
  assign n54248 = ~n54238 & ~n54241;
  assign n54249 = pi211 & n54248;
  assign n54250 = ~n54173 & ~n54249;
  assign n54251 = ~n65324 & ~n54250;
  assign n54252 = ~pi211 & ~n54248;
  assign n54253 = pi211 & ~n54233;
  assign n54254 = n39342 & ~n54253;
  assign n54255 = ~n54252 & n54254;
  assign n54256 = ~n54158 & ~n54255;
  assign n54257 = ~n54251 & n54256;
  assign n54258 = ~n54243 & n54247;
  assign n54259 = ~pi219 & ~n65446;
  assign n54260 = ~n54236 & ~n54259;
  assign n54261 = ~pi209 & ~n54260;
  assign n54262 = n62455 & ~n54261;
  assign n54263 = ~n54227 & n54262;
  assign n54264 = n39342 & ~n53797;
  assign n54265 = ~n65324 & ~n52605;
  assign n54266 = ~pi219 & ~n54265;
  assign n54267 = ~pi219 & ~n54264;
  assign n54268 = ~n54265 & n54267;
  assign n54269 = ~n54264 & n54266;
  assign n54270 = ~n65172 & ~n54186;
  assign n54271 = ~n54186 & ~n65447;
  assign n54272 = ~n65172 & n54271;
  assign n54273 = ~n65447 & n54270;
  assign n54274 = ~pi213 & ~n65448;
  assign n54275 = ~n54263 & n54274;
  assign n54276 = ~n54193 & ~n54275;
  assign n54277 = pi230 & ~n54276;
  assign po392 = ~n54074 & ~n54277;
  assign n54279 = ~pi230 & pi238;
  assign n54280 = n49599 & n50231;
  assign n54281 = n53887 & ~n54280;
  assign n54282 = pi207 & ~n54281;
  assign n54283 = ~n54239 & ~n54282;
  assign n54284 = pi208 & ~n54283;
  assign n54285 = ~n54238 & ~n54284;
  assign n54286 = pi211 & ~n54285;
  assign n54287 = ~n49595 & n54026;
  assign n54288 = ~pi1154 & ~n53943;
  assign n54289 = ~n49832 & n54288;
  assign n54290 = pi207 & ~n54289;
  assign n54291 = n53887 & n54290;
  assign n54292 = pi208 & ~n54291;
  assign n54293 = ~n54287 & n54292;
  assign n54294 = ~n54160 & n54293;
  assign n54295 = ~n54159 & ~n54294;
  assign n54296 = ~pi211 & ~n54295;
  assign n54297 = n52527 & ~n54296;
  assign n54298 = ~n54286 & n54297;
  assign n54299 = n52855 & ~n54285;
  assign n54300 = n52776 & ~n54295;
  assign n54301 = ~n50428 & ~n53864;
  assign n54302 = pi207 & ~n54301;
  assign n54303 = ~n54230 & ~n54302;
  assign n54304 = pi208 & ~n54303;
  assign n54305 = ~n54229 & ~n54304;
  assign n54306 = n39343 & ~n54305;
  assign n54307 = pi212 & ~n54306;
  assign n54308 = ~n54300 & n54307;
  assign n54309 = ~n54299 & n54308;
  assign n54310 = ~n54298 & ~n54309;
  assign n54311 = ~pi219 & ~n54310;
  assign n54312 = n38985 & ~n54280;
  assign n54313 = ~n53864 & n54312;
  assign n54314 = ~n54137 & ~n54313;
  assign n54315 = pi211 & n54314;
  assign n54316 = ~pi211 & ~n54305;
  assign n54317 = ~n54315 & ~n54316;
  assign n54318 = n53038 & n54317;
  assign n54319 = ~pi214 & ~n54314;
  assign n54320 = ~pi212 & n54319;
  assign n54321 = pi209 & n62455;
  assign n54322 = ~n54320 & n54321;
  assign n54323 = ~n54318 & n54322;
  assign n54324 = ~n54311 & n54323;
  assign n54325 = ~n48475 & ~n50343;
  assign n54326 = pi207 & ~n54325;
  assign n54327 = ~n53894 & ~n54326;
  assign n54328 = ~pi208 & ~n54327;
  assign n54329 = pi200 & pi207;
  assign n54330 = ~pi199 & ~n54329;
  assign n54331 = ~pi299 & ~n54330;
  assign n54332 = pi208 & ~n54331;
  assign n54333 = ~pi207 & n39538;
  assign n54334 = ~pi299 & ~n54333;
  assign n54335 = ~pi1153 & ~n54334;
  assign n54336 = n54332 & ~n54335;
  assign n54337 = ~n54328 & ~n54336;
  assign n54338 = pi211 & ~n54337;
  assign n54339 = ~pi207 & ~n50085;
  assign n54340 = ~n53230 & ~n54339;
  assign n54341 = pi208 & ~n54340;
  assign n54342 = ~n50085 & n52766;
  assign n54343 = ~n54341 & ~n54342;
  assign n54344 = ~pi211 & ~n52768;
  assign n54345 = ~n54343 & n54344;
  assign n54346 = ~n54338 & ~n54345;
  assign n54347 = n39342 & ~n54346;
  assign n54348 = ~n65324 & ~n54343;
  assign n54349 = pi299 & n52605;
  assign n54350 = n54348 & ~n54349;
  assign n54351 = ~n54347 & ~n54350;
  assign n54352 = ~pi219 & ~n54351;
  assign n54353 = ~n38985 & n50050;
  assign n54354 = ~pi299 & ~n53031;
  assign n54355 = pi200 & n38985;
  assign n54356 = pi208 & n54329;
  assign n54357 = ~pi199 & ~n65449;
  assign n54358 = ~n53032 & ~n53143;
  assign n54359 = n48567 & ~n54358;
  assign n54360 = n54354 & n54357;
  assign n54361 = ~n54353 & n65450;
  assign n54362 = ~pi211 & n52642;
  assign n54363 = ~n52517 & n54362;
  assign n54364 = ~n54361 & ~n54363;
  assign n54365 = ~n52967 & ~n54364;
  assign n54366 = ~n54352 & ~n54365;
  assign n54367 = n65182 & ~n54366;
  assign n54368 = n53857 & ~n53902;
  assign n54369 = pi208 & ~n54368;
  assign n54370 = n52766 & ~n53858;
  assign n54371 = ~n54369 & ~n54370;
  assign n54372 = ~pi211 & ~n54371;
  assign n54373 = ~n52802 & n54372;
  assign n54374 = pi211 & ~n54371;
  assign n54375 = ~n52768 & n54374;
  assign n54376 = ~n54373 & ~n54375;
  assign n54377 = ~n65324 & ~n54376;
  assign n54378 = n39538 & n53032;
  assign n54379 = ~pi299 & ~n54378;
  assign n54380 = n50251 & ~n54379;
  assign n54381 = n49598 & n52548;
  assign n54382 = pi208 & n49595;
  assign n54383 = ~n54333 & n54382;
  assign n54384 = ~n54381 & ~n54383;
  assign n54385 = ~n54380 & n54384;
  assign n54386 = ~n54345 & n54385;
  assign n54387 = n39342 & ~n54386;
  assign n54388 = n48497 & n53032;
  assign n54389 = pi1153 & n54388;
  assign n54390 = n54384 & ~n54389;
  assign n54391 = ~pi214 & n54384;
  assign n54392 = ~n54389 & n54391;
  assign n54393 = ~pi212 & ~n54392;
  assign n54394 = ~pi214 & n54393;
  assign n54395 = n52517 & ~n54390;
  assign n54396 = ~pi219 & ~n65451;
  assign n54397 = ~n54387 & n54396;
  assign n54398 = ~n54377 & n54397;
  assign n54399 = ~n48494 & ~n54379;
  assign n54400 = ~pi214 & ~n54388;
  assign n54401 = ~pi212 & n54400;
  assign n54402 = n54399 & ~n54401;
  assign n54403 = pi1153 & n54402;
  assign n54404 = pi219 & n54384;
  assign n54405 = ~n54403 & n54404;
  assign n54406 = n50537 & ~n54405;
  assign n54407 = ~n54398 & n54406;
  assign n54408 = pi1152 & ~n54407;
  assign n54409 = ~n54367 & n54408;
  assign n54410 = ~n38985 & n49461;
  assign n54411 = ~n53031 & n54410;
  assign n54412 = n49461 & n53032;
  assign n54413 = n49598 & n53026;
  assign n54414 = ~n49598 & n52548;
  assign n54415 = pi208 & ~n54414;
  assign n54416 = pi200 & n52765;
  assign n54417 = n54415 & ~n54416;
  assign n54418 = ~pi299 & n54417;
  assign n54419 = ~n53107 & ~n54418;
  assign n54420 = ~n65452 & ~n54413;
  assign n54421 = ~n50128 & ~n50196;
  assign n54422 = ~n52738 & ~n54415;
  assign n54423 = ~n54421 & ~n54422;
  assign n54424 = ~n54413 & ~n54423;
  assign n54425 = ~pi299 & ~n54424;
  assign n54426 = ~n50055 & ~n65453;
  assign n54427 = ~pi214 & ~n65454;
  assign n54428 = ~pi212 & ~n54427;
  assign n54429 = pi299 & ~n52605;
  assign n54430 = pi214 & ~n54429;
  assign n54431 = ~n65454 & n54430;
  assign n54432 = n54428 & ~n54431;
  assign n54433 = n52776 & n54424;
  assign n54434 = ~pi299 & ~n53143;
  assign n54435 = ~pi208 & ~n54434;
  assign n54436 = ~n54417 & ~n54435;
  assign n54437 = ~n50076 & ~n54436;
  assign n54438 = n39343 & ~n54437;
  assign n54439 = ~n52640 & n52855;
  assign n54440 = ~n65454 & n54439;
  assign n54441 = pi212 & ~n54440;
  assign n54442 = ~n54438 & n54441;
  assign n54443 = ~n54433 & n54442;
  assign n54444 = ~pi219 & ~n54443;
  assign n54445 = ~n54432 & n54444;
  assign n54446 = ~pi211 & ~n54436;
  assign n54447 = pi211 & ~n65453;
  assign n54448 = ~n54446 & ~n54447;
  assign n54449 = ~n50076 & ~n54448;
  assign n54450 = n52517 & ~n65454;
  assign n54451 = n54449 & ~n54450;
  assign n54452 = pi219 & ~n54451;
  assign n54453 = n50537 & ~n54452;
  assign n54454 = ~n54445 & n54453;
  assign n54455 = ~n52640 & ~n54389;
  assign n54456 = ~pi211 & ~n54455;
  assign n54457 = n39342 & ~n54380;
  assign n54458 = ~n54456 & n54457;
  assign n54459 = ~n65324 & ~n54429;
  assign n54460 = ~n54389 & n54459;
  assign n54461 = ~n54458 & ~n54460;
  assign n54462 = ~pi219 & ~n54461;
  assign n54463 = ~n52967 & ~n54403;
  assign n54464 = n65182 & ~n54463;
  assign n54465 = ~n54462 & n54464;
  assign n54466 = ~pi1152 & ~n54465;
  assign n54467 = ~n54454 & n54466;
  assign n54468 = ~pi209 & ~n54467;
  assign n54469 = ~n54409 & n54468;
  assign n54470 = pi219 & n53815;
  assign n54471 = ~pi1153 & n39423;
  assign n54472 = n52520 & ~n65455;
  assign n54473 = ~n65447 & n54472;
  assign n54474 = ~n54469 & ~n54473;
  assign n54475 = ~n54409 & ~n54467;
  assign n54476 = ~pi209 & ~n54475;
  assign n54477 = n62455 & ~n54320;
  assign n54478 = ~n54318 & n54477;
  assign n54479 = ~n54311 & n54478;
  assign n54480 = pi209 & ~n54479;
  assign n54481 = ~n54476 & ~n54480;
  assign n54482 = ~n54473 & ~n54481;
  assign n54483 = ~n54324 & n54474;
  assign n54484 = pi213 & ~n65456;
  assign n54485 = ~n62455 & n65430;
  assign n54486 = ~pi1153 & n39424;
  assign n54487 = ~n39342 & n53815;
  assign n54488 = ~n39425 & ~n50176;
  assign n54489 = ~n39342 & ~n53815;
  assign n54490 = ~n52909 & ~n54489;
  assign n54491 = ~n64625 & ~n65457;
  assign n54492 = n54485 & ~n65458;
  assign n54493 = n54485 & ~n65457;
  assign n54494 = ~n39346 & n52520;
  assign n54495 = pi1151 & ~n54494;
  assign n54496 = ~n65459 & n54495;
  assign n54497 = ~n54141 & n54292;
  assign n54498 = ~n54140 & ~n54497;
  assign n54499 = ~pi211 & ~n54498;
  assign n54500 = ~n54315 & ~n54499;
  assign n54501 = ~n52517 & n54500;
  assign n54502 = ~n54320 & ~n54501;
  assign n54503 = pi219 & ~n54502;
  assign n54504 = n62455 & ~n54503;
  assign n54505 = pi211 & ~n54498;
  assign n54506 = ~n54316 & ~n54505;
  assign n54507 = pi214 & n54506;
  assign n54508 = ~pi212 & ~n54319;
  assign n54509 = ~n54507 & n54508;
  assign n54510 = ~pi219 & ~n54509;
  assign n54511 = ~pi214 & ~n54506;
  assign n54512 = pi214 & ~n54498;
  assign n54513 = ~n54511 & ~n54512;
  assign n54514 = pi212 & ~n54513;
  assign n54515 = n54510 & ~n54514;
  assign n54516 = n54504 & ~n54515;
  assign n54517 = n54496 & ~n54516;
  assign n54518 = ~pi1151 & ~n65459;
  assign n54519 = pi214 & ~n54500;
  assign n54520 = ~n54511 & ~n54519;
  assign n54521 = pi212 & ~n54520;
  assign n54522 = n54510 & ~n54521;
  assign n54523 = pi219 & ~n54314;
  assign n54524 = n62455 & ~n54523;
  assign n54525 = ~n54522 & n54524;
  assign n54526 = n54518 & ~n54525;
  assign n54527 = pi1152 & ~n54526;
  assign n54528 = pi1152 & ~n54517;
  assign n54529 = ~n54526 & n54528;
  assign n54530 = ~n54517 & n54527;
  assign n54531 = pi1153 & n65364;
  assign n54532 = n50176 & ~n65324;
  assign n54533 = n39346 & ~n65461;
  assign n54534 = n52520 & ~n54533;
  assign n54535 = pi1151 & ~n54534;
  assign n54536 = pi214 & n54317;
  assign n54537 = ~n54319 & ~n54536;
  assign n54538 = ~pi212 & ~n54537;
  assign n54539 = ~pi211 & n54314;
  assign n54540 = ~n54505 & ~n54539;
  assign n54541 = pi214 & ~n54540;
  assign n54542 = ~pi214 & ~n54317;
  assign n54543 = pi212 & ~n54542;
  assign n54544 = pi212 & ~n54541;
  assign n54545 = ~n54542 & n54544;
  assign n54546 = ~n54541 & n54543;
  assign n54547 = ~n54538 & ~n65462;
  assign n54548 = ~pi219 & ~n54547;
  assign n54549 = n54504 & ~n54548;
  assign n54550 = n54535 & ~n54549;
  assign n54551 = n64656 & ~n52517;
  assign n54552 = n39424 & n52967;
  assign n54553 = n39421 & ~n65324;
  assign n54554 = ~pi219 & ~n65324;
  assign n54555 = n48935 & n54554;
  assign n54556 = n39346 & ~n65364;
  assign n54557 = n54485 & ~n54556;
  assign n54558 = n65364 & n54485;
  assign n54559 = ~n62455 & n65463;
  assign n54560 = pi1153 & n65464;
  assign n54561 = n50558 & n65461;
  assign n54562 = ~pi1151 & ~n65465;
  assign n54563 = n54317 & n54554;
  assign n54564 = ~n54314 & ~n54554;
  assign n54565 = n62455 & ~n54564;
  assign n54566 = ~n54563 & n54565;
  assign n54567 = n54562 & ~n54566;
  assign n54568 = ~pi1152 & ~n54567;
  assign n54569 = ~n54550 & n54568;
  assign n54570 = pi209 & ~n54569;
  assign n54571 = ~n54550 & ~n54567;
  assign n54572 = ~pi1152 & ~n54571;
  assign n54573 = ~n54517 & ~n54526;
  assign n54574 = pi1152 & ~n54573;
  assign n54575 = ~n54572 & ~n54574;
  assign n54576 = pi209 & ~n54575;
  assign n54577 = pi209 & ~n65460;
  assign n54578 = ~n54569 & n54577;
  assign n54579 = ~n65460 & n54570;
  assign n54580 = ~pi214 & n54449;
  assign n54581 = ~n48494 & ~n54389;
  assign n54582 = ~n65454 & n54581;
  assign n54583 = pi214 & ~n54582;
  assign n54584 = pi212 & ~n54583;
  assign n54585 = ~n54580 & n54584;
  assign n54586 = ~pi212 & ~n54451;
  assign n54587 = ~n54585 & ~n54586;
  assign n54588 = ~pi219 & ~n54587;
  assign n54589 = ~n48498 & ~n54389;
  assign n54590 = ~n65454 & n54589;
  assign n54591 = ~n54450 & ~n54590;
  assign n54592 = pi219 & ~n54591;
  assign n54593 = n62455 & ~n54592;
  assign n54594 = ~n54588 & n54593;
  assign n54595 = n54535 & ~n54594;
  assign n54596 = n54400 & n54403;
  assign n54597 = pi212 & ~n54400;
  assign n54598 = ~n54581 & n54597;
  assign n54599 = ~pi219 & ~n54598;
  assign n54600 = n52527 & n54362;
  assign n54601 = n52642 & n53068;
  assign n54602 = ~n54388 & ~n65467;
  assign n54603 = n54599 & n54602;
  assign n54604 = ~n54596 & n54603;
  assign n54605 = pi219 & ~n54388;
  assign n54606 = n62455 & ~n54605;
  assign n54607 = n54403 & n54606;
  assign n54608 = ~n54604 & n54607;
  assign n54609 = n54562 & ~n54608;
  assign n54610 = ~pi1152 & ~n54609;
  assign n54611 = ~n54595 & n54610;
  assign n54612 = ~n54372 & n54390;
  assign n54613 = ~pi212 & n54392;
  assign n54614 = pi214 & n54612;
  assign n54615 = ~n54392 & ~n54614;
  assign n54616 = ~pi212 & ~n54615;
  assign n54617 = ~n54612 & ~n54616;
  assign n54618 = ~n54612 & ~n54613;
  assign n54619 = pi219 & ~n65468;
  assign n54620 = n62455 & ~n54619;
  assign n54621 = pi1153 & ~n54379;
  assign n54622 = ~n54374 & ~n54621;
  assign n54623 = n54391 & n54622;
  assign n54624 = pi214 & n54371;
  assign n54625 = pi212 & ~n54624;
  assign n54626 = ~n54623 & n54625;
  assign n54627 = pi214 & n54384;
  assign n54628 = n54622 & n54627;
  assign n54629 = n54393 & ~n54628;
  assign n54630 = ~pi219 & ~n54629;
  assign n54631 = ~pi219 & ~n54626;
  assign n54632 = ~n54629 & n54631;
  assign n54633 = ~n54626 & n54630;
  assign n54634 = n54620 & ~n65469;
  assign n54635 = n54496 & ~n54634;
  assign n54636 = pi219 & ~n54361;
  assign n54637 = n62455 & ~n54636;
  assign n54638 = ~pi211 & n54337;
  assign n54639 = n54348 & ~n54638;
  assign n54640 = n65324 & n54361;
  assign n54641 = pi299 & n52909;
  assign n54642 = ~pi219 & ~n54641;
  assign n54643 = ~n54640 & n54642;
  assign n54644 = ~n54639 & n54643;
  assign n54645 = n54637 & ~n54644;
  assign n54646 = n54518 & ~n54645;
  assign n54647 = pi1152 & ~n54646;
  assign n54648 = ~n54635 & n54647;
  assign n54649 = ~n54635 & ~n54646;
  assign n54650 = pi1152 & ~n54649;
  assign n54651 = ~n54595 & ~n54609;
  assign n54652 = ~pi1152 & ~n54651;
  assign n54653 = ~n54650 & ~n54652;
  assign n54654 = ~n54611 & ~n54648;
  assign n54655 = ~pi209 & ~n65470;
  assign n54656 = ~pi213 & ~n54655;
  assign n54657 = ~n65466 & n54656;
  assign n54658 = ~n54484 & ~n54657;
  assign n54659 = pi230 & ~n54658;
  assign n54660 = ~n54279 & ~n54659;
  assign n54661 = ~pi230 & ~pi239;
  assign n54662 = n52555 & ~n52696;
  assign n54663 = ~pi214 & n54662;
  assign n54664 = ~pi212 & ~n54663;
  assign n54665 = ~pi219 & n54664;
  assign n54666 = ~pi208 & n53220;
  assign n54667 = pi299 & pi1158;
  assign n54668 = ~n52555 & n54667;
  assign n54669 = ~pi211 & ~n54668;
  assign n54670 = ~n54666 & n54669;
  assign n54671 = ~pi1157 & ~n54662;
  assign n54672 = pi208 & pi299;
  assign n54673 = pi1157 & ~n54672;
  assign n54674 = ~n53803 & n54673;
  assign n54675 = ~n54671 & ~n54674;
  assign n54676 = pi211 & ~n54675;
  assign n54677 = pi214 & ~n54676;
  assign n54678 = ~n54666 & ~n54668;
  assign n54679 = ~pi211 & ~n54678;
  assign n54680 = pi211 & ~n54671;
  assign n54681 = ~n54674 & n54680;
  assign n54682 = ~n54679 & ~n54681;
  assign n54683 = pi214 & ~n54682;
  assign n54684 = ~n54670 & n54677;
  assign n54685 = n54665 & ~n65471;
  assign n54686 = pi219 & n54664;
  assign n54687 = ~n53740 & n54012;
  assign n54688 = pi211 & ~n54662;
  assign n54689 = pi214 & ~n54688;
  assign n54690 = ~n54687 & n54689;
  assign n54691 = n54686 & ~n54690;
  assign n54692 = pi212 & ~n54662;
  assign n54693 = n62455 & ~n54692;
  assign n54694 = ~pi209 & n54693;
  assign n54695 = ~n54691 & n54694;
  assign n54696 = ~n54685 & n54695;
  assign n54697 = ~pi214 & n65397;
  assign n54698 = ~pi212 & ~n54697;
  assign n54699 = ~pi219 & n54698;
  assign n54700 = pi208 & ~n54667;
  assign n54701 = ~n52737 & ~n54700;
  assign n54702 = ~n53238 & n54701;
  assign n54703 = n53246 & ~n54702;
  assign n54704 = ~n53204 & n54673;
  assign n54705 = ~n53184 & ~n54704;
  assign n54706 = pi211 & ~n54705;
  assign n54707 = pi214 & ~n54706;
  assign n54708 = ~n54703 & n54707;
  assign n54709 = n54699 & ~n54708;
  assign n54710 = pi219 & n54698;
  assign n54711 = pi211 & ~n65397;
  assign n54712 = ~n65397 & n54012;
  assign n54713 = pi214 & ~n54712;
  assign n54714 = ~n54711 & n54713;
  assign n54715 = n54710 & ~n54714;
  assign n54716 = pi212 & ~n65397;
  assign n54717 = n62455 & ~n54716;
  assign n54718 = pi209 & n54717;
  assign n54719 = ~n54715 & n54718;
  assign n54720 = ~n54709 & n54718;
  assign n54721 = ~n54715 & n54720;
  assign n54722 = ~n54709 & n54719;
  assign n54723 = ~n53064 & ~n53072;
  assign n54724 = pi213 & ~n54723;
  assign n54725 = ~n65472 & n54724;
  assign n54726 = ~n54696 & n54725;
  assign n54727 = ~pi211 & ~n52640;
  assign n54728 = ~n65397 & n54727;
  assign n54729 = pi214 & ~n54711;
  assign n54730 = ~n54728 & n54729;
  assign n54731 = n54710 & ~n54730;
  assign n54732 = pi211 & ~n49607;
  assign n54733 = ~n65397 & n54732;
  assign n54734 = n54713 & ~n54733;
  assign n54735 = n54699 & ~n54734;
  assign n54736 = n54717 & ~n54735;
  assign n54737 = n54717 & ~n54731;
  assign n54738 = ~n54735 & n54737;
  assign n54739 = ~n54731 & n54736;
  assign n54740 = pi209 & ~n65473;
  assign n54741 = ~n52640 & ~n53762;
  assign n54742 = n54689 & ~n54741;
  assign n54743 = n54686 & ~n54742;
  assign n54744 = ~n53750 & n54732;
  assign n54745 = pi214 & ~n54744;
  assign n54746 = ~n54687 & n54745;
  assign n54747 = n54665 & ~n54746;
  assign n54748 = n54693 & ~n54747;
  assign n54749 = n54693 & ~n54743;
  assign n54750 = ~n54747 & n54749;
  assign n54751 = ~n54743 & n54748;
  assign n54752 = ~pi209 & ~n65474;
  assign n54753 = ~n54740 & ~n54752;
  assign n54754 = n52527 & ~n54056;
  assign n54755 = n50279 & n54754;
  assign n54756 = ~pi213 & ~n54755;
  assign n54757 = ~n54753 & n54756;
  assign n54758 = ~n54726 & ~n54757;
  assign n54759 = pi230 & ~n54758;
  assign po396 = ~n54661 & ~n54759;
  assign n54761 = ~pi211 & pi1146;
  assign n54762 = pi211 & pi1145;
  assign n54763 = ~n54761 & ~n54762;
  assign n54764 = pi214 & ~n54763;
  assign n54765 = pi211 & pi1146;
  assign n54766 = ~pi214 & n54765;
  assign n54767 = ~n54764 & ~n54766;
  assign n54768 = pi212 & ~n54767;
  assign n54769 = n52527 & n54765;
  assign n54770 = ~n54768 & ~n54769;
  assign n54771 = ~n53038 & n54770;
  assign n54772 = ~n62455 & n53007;
  assign n54773 = ~n50558 & ~n54772;
  assign n54774 = ~n54771 & ~n54773;
  assign n54775 = pi1147 & ~n65464;
  assign n54776 = ~n54774 & n54775;
  assign n54777 = n62455 & ~n52519;
  assign n54778 = ~pi211 & n53272;
  assign n54779 = pi219 & ~n54778;
  assign n54780 = n54777 & ~n54779;
  assign n54781 = pi219 & n65453;
  assign n54782 = n62455 & ~n54781;
  assign n54783 = ~n54780 & ~n54782;
  assign n54784 = pi299 & pi1146;
  assign n54785 = n65453 & ~n54784;
  assign n54786 = pi211 & ~n54785;
  assign n54787 = ~n54446 & ~n54786;
  assign n54788 = ~pi214 & n54787;
  assign n54789 = pi299 & ~n54763;
  assign n54790 = pi214 & ~n54789;
  assign n54791 = n65453 & n54790;
  assign n54792 = pi212 & ~n54791;
  assign n54793 = ~n54788 & n54792;
  assign n54794 = ~pi214 & n65453;
  assign n54795 = ~pi212 & ~n54794;
  assign n54796 = pi214 & n54787;
  assign n54797 = n54795 & ~n54796;
  assign n54798 = ~pi219 & ~n54797;
  assign n54799 = ~pi219 & ~n54793;
  assign n54800 = ~n54797 & n54799;
  assign n54801 = ~n54793 & n54798;
  assign n54802 = ~n54783 & ~n65475;
  assign n54803 = n54776 & ~n54802;
  assign n54804 = n65014 & n54378;
  assign n54805 = n62455 & n54388;
  assign n54806 = ~pi1147 & ~n54774;
  assign n54807 = pi219 & n54780;
  assign n54808 = pi299 & ~n54770;
  assign n54809 = n38010 & n54808;
  assign n54810 = ~n54807 & ~n54809;
  assign n54811 = n54806 & ~n54809;
  assign n54812 = ~n54807 & n54811;
  assign n54813 = n54806 & n54810;
  assign n54814 = ~n65476 & n65477;
  assign n54815 = ~pi1148 & ~n54814;
  assign n54816 = ~n54803 & n54815;
  assign n54817 = n48567 & n52555;
  assign n54818 = ~pi299 & ~n54817;
  assign n54819 = ~n48570 & n52766;
  assign n54820 = ~n54332 & ~n54819;
  assign n54821 = ~n54332 & n54818;
  assign n54822 = ~pi211 & ~n65478;
  assign n54823 = ~n52517 & n54822;
  assign n54824 = ~n52518 & n65450;
  assign n54825 = pi219 & ~n54824;
  assign n54826 = ~n54823 & n54825;
  assign n54827 = n62455 & ~n54826;
  assign n54828 = n48567 & n54827;
  assign n54829 = n52474 & ~n54826;
  assign n54830 = ~n54780 & ~n65479;
  assign n54831 = pi212 & ~n65478;
  assign n54832 = ~n65450 & n54767;
  assign n54833 = n54831 & ~n54832;
  assign n54834 = ~pi214 & ~n65450;
  assign n54835 = ~pi212 & ~n54834;
  assign n54836 = pi211 & n54784;
  assign n54837 = ~n65450 & ~n54836;
  assign n54838 = n54835 & ~n54837;
  assign n54839 = ~pi219 & ~n54838;
  assign n54840 = ~pi219 & ~n54833;
  assign n54841 = ~n54838 & n54840;
  assign n54842 = ~n54833 & n54839;
  assign n54843 = ~n54830 & ~n65480;
  assign n54844 = n54806 & ~n54843;
  assign n54845 = n49595 & ~n53031;
  assign n54846 = pi219 & ~n54845;
  assign n54847 = n62455 & ~n54846;
  assign n54848 = ~pi299 & ~n54845;
  assign n54849 = pi212 & ~n52776;
  assign n54850 = pi299 & n54849;
  assign n54851 = pi212 & ~n54850;
  assign n54852 = pi212 & ~n54848;
  assign n54853 = ~n54850 & n54852;
  assign n54854 = ~n54848 & n54851;
  assign n54855 = pi214 & pi299;
  assign n54856 = ~pi211 & n54855;
  assign n54857 = ~n54845 & ~n54856;
  assign n54858 = pi211 & ~n54845;
  assign n54859 = ~n54845 & ~n54855;
  assign n54860 = ~pi212 & ~n54859;
  assign n54861 = ~n54858 & n54860;
  assign n54862 = ~pi212 & ~n54857;
  assign n54863 = ~pi219 & ~n65482;
  assign n54864 = ~pi219 & ~n65481;
  assign n54865 = ~n65482 & n54864;
  assign n54866 = ~n65481 & n54863;
  assign n54867 = n54847 & ~n65483;
  assign n54868 = n54810 & ~n54867;
  assign n54869 = n54776 & n54810;
  assign n54870 = ~n54867 & n54869;
  assign n54871 = n54776 & n54868;
  assign n54872 = pi1148 & ~n65484;
  assign n54873 = ~n54844 & n54872;
  assign n54874 = pi1149 & ~n54873;
  assign n54875 = ~n54816 & n54874;
  assign n54876 = n54384 & ~n54789;
  assign n54877 = n39342 & ~n54876;
  assign n54878 = ~pi1146 & n48494;
  assign n54879 = ~n65324 & ~n54878;
  assign n54880 = ~n54877 & ~n54879;
  assign n54881 = n49519 & ~n54329;
  assign n54882 = pi208 & ~n54881;
  assign n54883 = ~pi199 & ~n54882;
  assign n54884 = ~n54384 & ~n54883;
  assign n54885 = ~pi299 & ~n54884;
  assign n54886 = ~pi219 & ~n54885;
  assign n54887 = ~n54880 & n54886;
  assign n54888 = n53007 & n53041;
  assign n54889 = n53038 & n54778;
  assign n54890 = ~n52967 & n54884;
  assign n54891 = ~n65485 & ~n54890;
  assign n54892 = pi219 & ~n54884;
  assign n54893 = ~n54885 & ~n54892;
  assign n54894 = ~n54879 & ~n54890;
  assign n54895 = ~n54877 & n54894;
  assign n54896 = n54893 & ~n54895;
  assign n54897 = ~n65485 & ~n54896;
  assign n54898 = ~n54887 & n54891;
  assign n54899 = n62455 & ~n65486;
  assign n54900 = n54776 & ~n54899;
  assign n54901 = ~pi1148 & ~n65477;
  assign n54902 = ~n54900 & n54901;
  assign n54903 = ~n53032 & ~n53230;
  assign n54904 = ~n38985 & n49800;
  assign n54905 = ~n54903 & ~n54904;
  assign n54906 = n54334 & n54905;
  assign n54907 = n62455 & n54906;
  assign n54908 = n65477 & ~n54907;
  assign n54909 = n62455 & ~n54384;
  assign n54910 = ~n54780 & ~n54909;
  assign n54911 = ~n48498 & ~n54836;
  assign n54912 = n54384 & n54911;
  assign n54913 = ~n65324 & ~n54912;
  assign n54914 = n52517 & ~n54384;
  assign n54915 = ~pi219 & ~n54914;
  assign n54916 = ~n54877 & n54915;
  assign n54917 = ~n54913 & n54915;
  assign n54918 = ~n54877 & n54917;
  assign n54919 = ~n54913 & n54916;
  assign n54920 = ~n54910 & ~n65487;
  assign n54921 = n54776 & ~n54920;
  assign n54922 = pi1148 & ~n54921;
  assign n54923 = pi1148 & ~n54908;
  assign n54924 = ~n54921 & n54923;
  assign n54925 = ~n54908 & n54922;
  assign n54926 = ~pi1149 & ~n65488;
  assign n54927 = ~pi1148 & ~n54900;
  assign n54928 = ~n54922 & ~n54927;
  assign n54929 = ~n65477 & ~n54928;
  assign n54930 = n54907 & n54922;
  assign n54931 = ~pi1149 & ~n54930;
  assign n54932 = ~n54929 & n54931;
  assign n54933 = ~pi1149 & ~n54902;
  assign n54934 = ~n65488 & n54933;
  assign n54935 = ~n54902 & n54926;
  assign n54936 = pi209 & ~n65489;
  assign n54937 = ~n54875 & n54936;
  assign n54938 = ~pi199 & pi1146;
  assign n54939 = pi200 & ~n54938;
  assign n54940 = ~pi299 & ~n54939;
  assign n54941 = pi199 & pi1145;
  assign n54942 = n49457 & ~n54941;
  assign n54943 = n54940 & ~n54942;
  assign n54944 = n52555 & n54943;
  assign n54945 = ~pi207 & n54943;
  assign n54946 = ~pi200 & ~n54941;
  assign n54947 = ~n54938 & n54946;
  assign n54948 = pi200 & ~n53029;
  assign n54949 = n52548 & ~n54948;
  assign n54950 = ~n54947 & n54949;
  assign n54951 = ~n54784 & ~n54950;
  assign n54952 = ~n54945 & n54951;
  assign n54953 = pi208 & ~n54952;
  assign n54954 = ~n54944 & ~n54953;
  assign n54955 = ~pi299 & n54954;
  assign n54956 = pi211 & ~n54955;
  assign n54957 = ~n53269 & n54956;
  assign n54958 = n54790 & n54954;
  assign n54959 = n39343 & ~n54955;
  assign n54960 = ~n54958 & ~n54959;
  assign n54961 = ~n54957 & ~n54960;
  assign n54962 = ~pi214 & n54911;
  assign n54963 = n54954 & n54962;
  assign n54964 = pi212 & ~n54963;
  assign n54965 = ~n54961 & n54964;
  assign n54966 = ~n53032 & ~n54950;
  assign n54967 = ~n38985 & ~n54943;
  assign n54968 = ~n54966 & ~n54967;
  assign n54969 = ~pi211 & ~n54955;
  assign n54970 = ~n54968 & ~n54969;
  assign n54971 = ~pi214 & ~n54968;
  assign n54972 = ~pi212 & ~n54971;
  assign n54973 = ~n54970 & n54972;
  assign n54974 = n54940 & ~n54946;
  assign n54975 = ~n38985 & ~n54974;
  assign n54976 = n54945 & n54946;
  assign n54977 = n54953 & ~n54976;
  assign n54978 = n52555 & n54974;
  assign n54979 = ~n54977 & ~n54978;
  assign n54980 = ~pi299 & ~n54979;
  assign n54981 = ~n54966 & ~n54975;
  assign n54982 = ~n54836 & ~n65490;
  assign n54983 = ~pi214 & ~n65490;
  assign n54984 = ~pi212 & ~n54983;
  assign n54985 = ~n54982 & n54984;
  assign n54986 = ~pi219 & ~n54985;
  assign n54987 = ~n54973 & n54986;
  assign n54988 = ~pi219 & ~n54973;
  assign n54989 = ~n54965 & ~n54985;
  assign n54990 = n54988 & n54989;
  assign n54991 = ~n54965 & n54987;
  assign n54992 = ~n52518 & n54968;
  assign n54993 = pi219 & ~n54992;
  assign n54994 = ~n53269 & n54969;
  assign n54995 = ~n52517 & n54994;
  assign n54996 = n54993 & ~n54995;
  assign n54997 = n62455 & ~n54996;
  assign n54998 = ~n65491 & n54997;
  assign n54999 = n54776 & ~n54998;
  assign n55000 = n54790 & ~n65490;
  assign n55001 = ~pi214 & n54982;
  assign n55002 = pi212 & ~n55001;
  assign n55003 = ~n55000 & n55002;
  assign n55004 = n54986 & ~n55003;
  assign n55005 = n52517 & n65490;
  assign n55006 = pi219 & ~n55005;
  assign n55007 = ~n52517 & n65490;
  assign n55008 = ~n52518 & ~n55007;
  assign n55009 = ~pi211 & ~n53272;
  assign n55010 = ~n65490 & n55009;
  assign n55011 = ~n55008 & ~n55010;
  assign n55012 = n55006 & ~n55011;
  assign n55013 = n62455 & ~n55012;
  assign n55014 = n62455 & ~n55004;
  assign n55015 = ~n55012 & n55014;
  assign n55016 = ~n55004 & n55013;
  assign n55017 = n54806 & ~n65492;
  assign n55018 = ~n54999 & ~n55017;
  assign n55019 = ~pi209 & n55018;
  assign n55020 = ~pi213 & ~n55019;
  assign n55021 = ~n54937 & n55020;
  assign n55022 = ~pi299 & n54979;
  assign n55023 = ~n52517 & n55022;
  assign n55024 = n39342 & n54970;
  assign n55025 = ~n55023 & ~n55024;
  assign n55026 = ~pi219 & ~n55025;
  assign n55027 = ~n52967 & ~n65490;
  assign n55028 = n62455 & ~n55027;
  assign n55029 = pi214 & n54970;
  assign n55030 = ~n55022 & ~n55029;
  assign n55031 = pi212 & ~n55030;
  assign n55032 = pi214 & ~n55022;
  assign n55033 = ~pi214 & n65490;
  assign n55034 = ~pi212 & ~n55033;
  assign n55035 = ~n55032 & n55034;
  assign n55036 = ~n55031 & ~n55035;
  assign n55037 = ~pi219 & ~n55036;
  assign n55038 = pi219 & ~n65490;
  assign n55039 = n62455 & ~n55038;
  assign n55040 = ~n55037 & n55039;
  assign n55041 = ~n55026 & n55028;
  assign n55042 = ~pi1147 & ~n54485;
  assign n55043 = ~n65493 & n55042;
  assign n55044 = ~n52517 & n54969;
  assign n55045 = n54993 & ~n55044;
  assign n55046 = n62455 & ~n55045;
  assign n55047 = ~pi219 & ~n54968;
  assign n55048 = ~n52569 & n55047;
  assign n55049 = n55046 & ~n55048;
  assign n55050 = ~n48935 & ~n50558;
  assign n55051 = ~n52517 & ~n55050;
  assign n55052 = pi1147 & ~n55051;
  assign n55053 = ~n55049 & n55052;
  assign n55054 = pi1149 & ~n55053;
  assign n55055 = ~n55043 & n55054;
  assign n55056 = n50558 & ~n65362;
  assign n55057 = ~pi1147 & ~n55056;
  assign n55058 = ~n54956 & ~n55032;
  assign n55059 = pi212 & ~n55058;
  assign n55060 = ~n54959 & n55047;
  assign n55061 = ~n55059 & n55060;
  assign n55062 = n65493 & ~n55061;
  assign n55063 = n55057 & ~n55062;
  assign n55064 = ~pi219 & ~n54849;
  assign n55065 = ~pi219 & ~n52911;
  assign n55066 = ~n54849 & n55065;
  assign n55067 = ~n52911 & n55064;
  assign n55068 = n52520 & ~n65494;
  assign n55069 = pi1147 & ~n55068;
  assign n55070 = n55046 & ~n55061;
  assign n55071 = n55069 & ~n55070;
  assign n55072 = ~pi1149 & ~n55071;
  assign n55073 = ~n55063 & n55072;
  assign n55074 = ~n55055 & ~n55073;
  assign n55075 = pi1148 & ~n55074;
  assign n55076 = pi212 & ~n52855;
  assign n55077 = ~n53068 & ~n55076;
  assign n55078 = ~n54955 & ~n55077;
  assign n55079 = ~n52855 & ~n54955;
  assign n55080 = ~n54968 & ~n55079;
  assign n55081 = pi214 & ~n54968;
  assign n55082 = ~n54956 & n55081;
  assign n55083 = ~n54969 & n54971;
  assign n55084 = pi212 & ~n55083;
  assign n55085 = ~n55082 & n55084;
  assign n55086 = pi212 & ~n55082;
  assign n55087 = ~n55083 & n55086;
  assign n55088 = pi212 & ~n55080;
  assign n55089 = n54988 & ~n65495;
  assign n55090 = n55047 & ~n55078;
  assign n55091 = n55070 & ~n65496;
  assign n55092 = ~n54494 & ~n55091;
  assign n55093 = pi1147 & ~n55092;
  assign n55094 = ~pi57 & ~pi1147;
  assign n55095 = n3475 & n55094;
  assign n55096 = ~pi1147 & n62455;
  assign n55097 = n65490 & n65497;
  assign n55098 = ~pi1149 & ~n55097;
  assign n55099 = ~n55093 & n55098;
  assign n55100 = n52520 & ~n54556;
  assign n55101 = n55046 & ~n65496;
  assign n55102 = ~n55100 & ~n55101;
  assign n55103 = pi1147 & ~n55102;
  assign n55104 = ~pi1147 & n65463;
  assign n55105 = ~n55097 & ~n55104;
  assign n55106 = n65014 & n65463;
  assign n55107 = n54979 & n55106;
  assign n55108 = ~n55105 & ~n55107;
  assign n55109 = pi1149 & ~n55108;
  assign n55110 = ~n55103 & n55109;
  assign n55111 = ~pi1148 & ~n55110;
  assign n55112 = ~n55099 & n55111;
  assign n55113 = ~n55075 & ~n55112;
  assign n55114 = ~pi209 & ~n55113;
  assign n55115 = pi211 & ~n54436;
  assign n55116 = ~pi211 & ~n65453;
  assign n55117 = pi214 & ~n55116;
  assign n55118 = pi214 & ~n55115;
  assign n55119 = ~n55116 & n55118;
  assign n55120 = ~n55115 & n55117;
  assign n55121 = n39342 & ~n65498;
  assign n55122 = pi214 & n54448;
  assign n55123 = n54795 & ~n55122;
  assign n55124 = ~pi219 & ~n55123;
  assign n55125 = pi212 & ~n65498;
  assign n55126 = ~n54448 & n55125;
  assign n55127 = n55124 & ~n55126;
  assign n55128 = ~n55121 & n55127;
  assign n55129 = pi212 & ~n54448;
  assign n55130 = pi219 & ~n55129;
  assign n55131 = ~n55123 & n55130;
  assign n55132 = n62455 & ~n55131;
  assign n55133 = ~n55128 & n55132;
  assign n55134 = ~n55100 & ~n55133;
  assign n55135 = pi1147 & n55134;
  assign n55136 = n52475 & n65364;
  assign n55137 = ~n65476 & ~n55136;
  assign n55138 = ~pi1147 & n55137;
  assign n55139 = pi1149 & ~n55138;
  assign n55140 = ~n55135 & n55139;
  assign n55141 = pi299 & n39343;
  assign n55142 = ~pi212 & ~n55141;
  assign n55143 = n54384 & n55142;
  assign n55144 = ~n48498 & n54384;
  assign n55145 = ~n54391 & ~n55144;
  assign n55146 = n54384 & ~n54856;
  assign n55147 = ~pi214 & n48494;
  assign n55148 = pi212 & ~n55147;
  assign n55149 = ~n65499 & n55148;
  assign n55150 = ~n55143 & ~n55149;
  assign n55151 = ~pi219 & ~n55150;
  assign n55152 = ~pi219 & n54885;
  assign n55153 = ~n55151 & ~n55152;
  assign n55154 = ~pi211 & ~n55153;
  assign n55155 = ~pi212 & n65499;
  assign n55156 = ~pi219 & ~n55155;
  assign n55157 = ~pi214 & n55144;
  assign n55158 = pi212 & ~n55157;
  assign n55159 = ~n48494 & n54627;
  assign n55160 = n55158 & ~n55159;
  assign n55161 = n55156 & ~n55160;
  assign n55162 = pi219 & ~n48498;
  assign n55163 = n54777 & ~n55162;
  assign n55164 = ~n54909 & ~n55163;
  assign n55165 = ~n55161 & ~n55164;
  assign n55166 = ~n54885 & n55165;
  assign n55167 = ~n55154 & n55166;
  assign n55168 = ~n54494 & ~n55167;
  assign n55169 = pi1147 & ~pi1149;
  assign n55170 = ~n55168 & n55169;
  assign n55171 = ~n55140 & ~n55170;
  assign n55172 = ~pi1148 & ~n55171;
  assign n55173 = n52569 & n54777;
  assign n55174 = ~n65494 & n55173;
  assign n55175 = ~n54909 & ~n55174;
  assign n55176 = ~n54909 & ~n55068;
  assign n55177 = ~n55174 & n55176;
  assign n55178 = ~n55068 & n55175;
  assign n55179 = pi1147 & n65500;
  assign n55180 = n55069 & n55175;
  assign n55181 = ~n54906 & ~n55141;
  assign n55182 = ~pi212 & ~n55181;
  assign n55183 = ~pi219 & ~n55182;
  assign n55184 = ~pi299 & ~n54905;
  assign n55185 = pi214 & ~n55184;
  assign n55186 = ~pi214 & n54906;
  assign n55187 = ~pi212 & ~n55186;
  assign n55188 = ~n55185 & n55187;
  assign n55189 = ~pi214 & ~n55184;
  assign n55190 = pi211 & ~n54334;
  assign n55191 = ~pi211 & ~n55184;
  assign n55192 = ~n54906 & ~n55191;
  assign n55193 = ~n55184 & ~n55190;
  assign n55194 = pi214 & ~n65502;
  assign n55195 = n55185 & ~n55190;
  assign n55196 = pi212 & ~n65503;
  assign n55197 = ~n55189 & n55196;
  assign n55198 = ~n55188 & ~n55197;
  assign n55199 = ~n48494 & ~n54906;
  assign n55200 = ~n55185 & n55199;
  assign n55201 = pi212 & ~n55200;
  assign n55202 = n55198 & n55201;
  assign n55203 = n55183 & ~n55202;
  assign n55204 = pi219 & ~n54906;
  assign n55205 = n62455 & ~n55204;
  assign n55206 = ~n55203 & n55205;
  assign n55207 = ~n55056 & ~n55206;
  assign n55208 = ~pi1147 & n55207;
  assign n55209 = n55057 & ~n55206;
  assign n55210 = ~n65501 & ~n65504;
  assign n55211 = ~pi1149 & ~n55210;
  assign n55212 = n62455 & n65450;
  assign n55213 = ~n54606 & ~n55212;
  assign n55214 = pi214 & n65478;
  assign n55215 = n54835 & ~n55214;
  assign n55216 = ~pi219 & ~n55215;
  assign n55217 = pi211 & n65450;
  assign n55218 = pi214 & ~n55217;
  assign n55219 = ~n54822 & n55218;
  assign n55220 = pi212 & ~n55219;
  assign n55221 = ~n65478 & n55220;
  assign n55222 = n55216 & ~n55221;
  assign n55223 = ~n55213 & ~n55222;
  assign n55224 = ~n54485 & ~n55223;
  assign n55225 = ~pi1147 & ~n55224;
  assign n55226 = n65317 & ~n53031;
  assign n55227 = n62455 & n54845;
  assign n55228 = ~n55173 & ~n65505;
  assign n55229 = ~n55051 & n55228;
  assign n55230 = pi1147 & ~n55229;
  assign n55231 = pi1149 & ~n55230;
  assign n55232 = ~n55225 & n55231;
  assign n55233 = pi1148 & ~n55232;
  assign n55234 = ~pi1147 & n55224;
  assign n55235 = pi1147 & n55229;
  assign n55236 = pi1149 & ~n55235;
  assign n55237 = ~n55234 & n55236;
  assign n55238 = ~pi1149 & ~n65501;
  assign n55239 = ~n65504 & n55238;
  assign n55240 = ~n55237 & ~n55239;
  assign n55241 = pi1148 & ~n55240;
  assign n55242 = ~n55211 & n55233;
  assign n55243 = ~n55172 & ~n65506;
  assign n55244 = pi209 & ~n55243;
  assign n55245 = pi213 & ~n55244;
  assign n55246 = ~n55114 & n55245;
  assign n55247 = pi213 & n55243;
  assign n55248 = ~n54902 & ~n65488;
  assign n55249 = ~pi1149 & ~n55248;
  assign n55250 = ~n54816 & ~n54873;
  assign n55251 = pi1149 & ~n55250;
  assign n55252 = ~n55249 & ~n55251;
  assign n55253 = ~n54875 & ~n65489;
  assign n55254 = ~pi213 & n65507;
  assign n55255 = pi209 & ~n55254;
  assign n55256 = ~n55247 & n55255;
  assign n55257 = pi213 & ~n55075;
  assign n55258 = ~n55112 & n55257;
  assign n55259 = ~pi213 & ~n55018;
  assign n55260 = ~pi209 & ~n55259;
  assign n55261 = ~n55258 & n55260;
  assign n55262 = ~n55256 & ~n55261;
  assign n55263 = pi213 & ~n55243;
  assign n55264 = ~pi213 & ~n65489;
  assign n55265 = ~pi213 & ~n65507;
  assign n55266 = ~n54875 & n55264;
  assign n55267 = pi209 & ~n65509;
  assign n55268 = ~n55263 & n55267;
  assign n55269 = ~n55093 & ~n55097;
  assign n55270 = ~pi1149 & ~n55269;
  assign n55271 = ~n55103 & ~n55108;
  assign n55272 = pi1149 & ~n55271;
  assign n55273 = ~pi1148 & ~n55272;
  assign n55274 = ~n55270 & n55273;
  assign n55275 = pi1148 & ~n55055;
  assign n55276 = ~n55073 & n55275;
  assign n55277 = pi213 & ~n55276;
  assign n55278 = pi213 & ~n55274;
  assign n55279 = ~n55276 & n55278;
  assign n55280 = ~n55274 & n55277;
  assign n55281 = ~pi213 & n55018;
  assign n55282 = ~pi209 & ~n55281;
  assign n55283 = ~n65510 & n55282;
  assign n55284 = ~n55268 & ~n55283;
  assign n55285 = ~n55021 & ~n55246;
  assign n55286 = pi230 & n65508;
  assign n55287 = ~pi230 & ~pi240;
  assign n55288 = pi230 & ~n65508;
  assign n55289 = ~pi230 & pi240;
  assign n55290 = ~n55288 & ~n55289;
  assign n55291 = ~n55286 & ~n55287;
  assign n55292 = ~pi1151 & ~n55068;
  assign n55293 = pi219 & ~n54389;
  assign n55294 = n62455 & ~n55293;
  assign n55295 = ~n55163 & ~n55294;
  assign n55296 = ~n54637 & n55295;
  assign n55297 = n39342 & n54343;
  assign n55298 = ~n54401 & ~n54581;
  assign n55299 = ~n39342 & ~n54361;
  assign n55300 = ~n55298 & n55299;
  assign n55301 = ~n55297 & ~n55300;
  assign n55302 = ~pi219 & ~n55301;
  assign n55303 = ~n55296 & ~n55302;
  assign n55304 = pi1152 & ~n55303;
  assign n55305 = ~pi212 & ~n54379;
  assign n55306 = ~n54400 & n55305;
  assign n55307 = ~n48498 & n55306;
  assign n55308 = ~pi219 & ~n55307;
  assign n55309 = pi214 & ~n54399;
  assign n55310 = ~pi211 & n54400;
  assign n55311 = pi212 & ~n54379;
  assign n55312 = ~n55310 & n55311;
  assign n55313 = ~n55309 & n55312;
  assign n55314 = n55308 & ~n55313;
  assign n55315 = ~n54389 & n54599;
  assign n55316 = ~pi299 & n55315;
  assign n55317 = ~n55314 & ~n55316;
  assign n55318 = n55294 & n55317;
  assign n55319 = ~pi1152 & ~n55318;
  assign n55320 = ~n55295 & ~n55315;
  assign n55321 = n55319 & ~n55320;
  assign n55322 = ~n55304 & ~n55321;
  assign n55323 = n55292 & ~n55322;
  assign n55324 = n54393 & ~n54624;
  assign n55325 = ~pi219 & ~n55324;
  assign n55326 = pi212 & ~n54371;
  assign n55327 = n55325 & ~n55326;
  assign n55328 = pi1152 & ~n55327;
  assign n55329 = n54620 & n55328;
  assign n55330 = pi1151 & ~n55051;
  assign n55331 = ~pi299 & ~n54437;
  assign n55332 = ~n54450 & ~n55331;
  assign n55333 = ~pi219 & ~n55332;
  assign n55334 = ~pi1152 & n54593;
  assign n55335 = ~n55333 & n55334;
  assign n55336 = n55330 & ~n55335;
  assign n55337 = ~n55329 & n55336;
  assign n55338 = pi1150 & ~n55337;
  assign n55339 = pi1150 & ~n55323;
  assign n55340 = ~n55337 & n55339;
  assign n55341 = ~n55323 & n55338;
  assign n55342 = ~n54371 & ~n55077;
  assign n55343 = ~pi219 & n54390;
  assign n55344 = ~n52855 & ~n54371;
  assign n55345 = pi212 & n54390;
  assign n55346 = ~n55344 & n55345;
  assign n55347 = ~n54616 & ~n55346;
  assign n55348 = ~pi219 & ~n55347;
  assign n55349 = ~n55342 & n55343;
  assign n55350 = pi1152 & ~n65513;
  assign n55351 = n54620 & n55350;
  assign n55352 = pi1151 & ~n55100;
  assign n55353 = ~pi214 & ~n54590;
  assign n55354 = n54584 & ~n55353;
  assign n55355 = ~pi212 & ~n54591;
  assign n55356 = ~n55354 & ~n55355;
  assign n55357 = ~pi219 & ~n55356;
  assign n55358 = n55334 & ~n55357;
  assign n55359 = n55352 & ~n55358;
  assign n55360 = ~n55351 & n55359;
  assign n55361 = ~pi1151 & ~n54494;
  assign n55362 = ~pi1152 & ~n55320;
  assign n55363 = pi1152 & ~n54361;
  assign n55364 = n54599 & n55363;
  assign n55365 = ~n55296 & ~n55364;
  assign n55366 = ~n55362 & n55365;
  assign n55367 = ~n54361 & n54599;
  assign n55368 = pi1152 & ~n55367;
  assign n55369 = pi1152 & ~n55296;
  assign n55370 = ~n55367 & n55369;
  assign n55371 = ~n55296 & n55368;
  assign n55372 = ~pi1152 & n55320;
  assign n55373 = n55361 & ~n55372;
  assign n55374 = ~n65514 & n55373;
  assign n55375 = n55361 & ~n65514;
  assign n55376 = ~n55372 & n55375;
  assign n55377 = n55361 & ~n55366;
  assign n55378 = ~pi1150 & ~n65515;
  assign n55379 = ~n55360 & n55378;
  assign n55380 = pi1149 & ~n55379;
  assign n55381 = pi1149 & ~n65512;
  assign n55382 = ~n55379 & n55381;
  assign n55383 = ~n65512 & n55380;
  assign n55384 = pi1151 & ~n54485;
  assign n55385 = ~pi214 & n54436;
  assign n55386 = pi212 & ~n55385;
  assign n55387 = ~n55122 & n55386;
  assign n55388 = ~n54428 & ~n55387;
  assign n55389 = ~n55331 & ~n55388;
  assign n55390 = ~pi219 & ~n55389;
  assign n55391 = ~n54781 & ~n55390;
  assign n55392 = ~pi1152 & ~n55391;
  assign n55393 = ~n54909 & ~n55294;
  assign n55394 = ~pi214 & n54371;
  assign n55395 = pi212 & ~n55394;
  assign n55396 = ~n54614 & n55395;
  assign n55397 = pi1152 & n55325;
  assign n55398 = ~n55396 & n55397;
  assign n55399 = ~n55393 & ~n55398;
  assign n55400 = n55325 & ~n55396;
  assign n55401 = pi1152 & ~n55400;
  assign n55402 = ~pi1152 & ~n54781;
  assign n55403 = ~n55390 & n55402;
  assign n55404 = ~n55401 & ~n55403;
  assign n55405 = ~n55393 & ~n55404;
  assign n55406 = ~n55392 & n55399;
  assign n55407 = n55384 & ~n65517;
  assign n55408 = ~pi1151 & ~n55056;
  assign n55409 = ~n54361 & ~n55317;
  assign n55410 = n54637 & ~n55409;
  assign n55411 = pi1152 & ~n55410;
  assign n55412 = ~n55319 & ~n55411;
  assign n55413 = n55408 & ~n55412;
  assign n55414 = pi1150 & ~n55413;
  assign n55415 = ~n55407 & n55414;
  assign n55416 = ~pi1152 & ~n54389;
  assign n55417 = n65182 & ~n55416;
  assign n55418 = pi1152 & n54361;
  assign n55419 = ~pi1152 & n54389;
  assign n55420 = ~n55418 & ~n55419;
  assign n55421 = n65182 & ~n55420;
  assign n55422 = ~n55363 & n55417;
  assign n55423 = n54372 & n54554;
  assign n55424 = ~n54371 & n65463;
  assign n55425 = n54390 & ~n65519;
  assign n55426 = pi1152 & ~n55425;
  assign n55427 = n50523 & n65364;
  assign n55428 = ~n65454 & ~n55427;
  assign n55429 = ~pi1152 & ~n55428;
  assign n55430 = n62455 & ~n55429;
  assign n55431 = pi1152 & n54390;
  assign n55432 = ~n65519 & n55431;
  assign n55433 = ~pi1152 & ~n55427;
  assign n55434 = ~n65454 & n55433;
  assign n55435 = ~n55432 & ~n55434;
  assign n55436 = n62455 & ~n55435;
  assign n55437 = ~n55426 & n55430;
  assign n55438 = ~n62455 & ~n65463;
  assign n55439 = pi1151 & ~n55438;
  assign n55440 = ~n65520 & n55439;
  assign n55441 = n62455 & ~n55426;
  assign n55442 = n55439 & ~n55441;
  assign n55443 = n65182 & n54389;
  assign n55444 = ~n55428 & n55439;
  assign n55445 = ~n55443 & ~n55444;
  assign n55446 = ~pi1152 & ~n55445;
  assign n55447 = pi1152 & n65182;
  assign n55448 = n54361 & n55447;
  assign n55449 = ~n55446 & ~n55448;
  assign n55450 = ~n55442 & n55449;
  assign n55451 = ~n65518 & ~n55440;
  assign n55452 = ~pi1150 & ~n65521;
  assign n55453 = ~pi1149 & ~n55452;
  assign n55454 = ~n55415 & n55453;
  assign n55455 = ~n55415 & ~n55452;
  assign n55456 = ~pi1149 & ~n55455;
  assign n55457 = ~n65512 & ~n55379;
  assign n55458 = pi1149 & ~n55457;
  assign n55459 = ~n55456 & ~n55458;
  assign n55460 = ~n65516 & ~n55454;
  assign n55461 = ~pi213 & ~n55454;
  assign n55462 = ~n65516 & n55461;
  assign n55463 = ~pi213 & ~n65522;
  assign n55464 = pi213 & n65470;
  assign n55465 = pi209 & ~n55464;
  assign n55466 = ~n65523 & n55465;
  assign n55467 = ~n65422 & ~n55184;
  assign n55468 = pi214 & n55467;
  assign n55469 = n55187 & ~n55468;
  assign n55470 = ~pi214 & n55467;
  assign n55471 = n55196 & ~n55470;
  assign n55472 = ~n55469 & ~n55471;
  assign n55473 = ~pi219 & ~n55472;
  assign n55474 = n55205 & ~n55473;
  assign n55475 = n54518 & ~n55474;
  assign n55476 = pi211 & ~n65478;
  assign n55477 = ~pi211 & ~n52786;
  assign n55478 = ~n65478 & n55477;
  assign n55479 = ~n55476 & ~n55478;
  assign n55480 = ~pi214 & n55479;
  assign n55481 = n54831 & ~n55480;
  assign n55482 = pi214 & n55479;
  assign n55483 = n54835 & ~n55482;
  assign n55484 = ~pi219 & ~n55483;
  assign n55485 = ~pi219 & ~n55481;
  assign n55486 = ~n55483 & n55485;
  assign n55487 = ~n55481 & n55484;
  assign n55488 = n54827 & ~n65524;
  assign n55489 = n54496 & ~n55488;
  assign n55490 = pi1152 & ~n55489;
  assign n55491 = ~n55475 & n55490;
  assign n55492 = ~n52855 & ~n65478;
  assign n55493 = ~n65450 & ~n55492;
  assign n55494 = ~n65450 & ~n55476;
  assign n55495 = pi214 & n55494;
  assign n55496 = ~n54822 & n54834;
  assign n55497 = pi212 & ~n55496;
  assign n55498 = ~n55495 & n55497;
  assign n55499 = pi212 & ~n55493;
  assign n55500 = ~n55479 & n65525;
  assign n55501 = ~n55217 & ~n55478;
  assign n55502 = n54835 & ~n55501;
  assign n55503 = ~pi219 & ~n55502;
  assign n55504 = ~n55500 & n55503;
  assign n55505 = n54827 & ~n55504;
  assign n55506 = n54535 & ~n55505;
  assign n55507 = ~n54554 & n54906;
  assign n55508 = ~n52786 & ~n55184;
  assign n55509 = ~pi211 & ~n55508;
  assign n55510 = n54554 & ~n55190;
  assign n55511 = n54554 & ~n65502;
  assign n55512 = ~n55184 & n55510;
  assign n55513 = ~n55509 & n65526;
  assign n55514 = ~n55507 & ~n55513;
  assign n55515 = n62455 & ~n55514;
  assign n55516 = n54562 & ~n55515;
  assign n55517 = ~pi1152 & ~n55516;
  assign n55518 = ~pi1152 & ~n55506;
  assign n55519 = ~n55516 & n55518;
  assign n55520 = ~n55506 & n55517;
  assign n55521 = pi1150 & ~n65527;
  assign n55522 = ~n55491 & n55521;
  assign n55523 = pi219 & ~n54402;
  assign n55524 = n62455 & ~n55523;
  assign n55525 = n55308 & ~n55312;
  assign n55526 = n55524 & ~n55525;
  assign n55527 = ~n54604 & n55524;
  assign n55528 = n54496 & ~n55527;
  assign n55529 = n54496 & ~n55526;
  assign n55530 = ~n55527 & n55529;
  assign n55531 = ~n55526 & n55528;
  assign n55532 = n39346 & n52569;
  assign n55533 = pi299 & n65430;
  assign n55534 = ~n65458 & n65529;
  assign n55535 = ~n65457 & n65529;
  assign n55536 = n54518 & ~n65530;
  assign n55537 = pi1152 & ~n55536;
  assign n55538 = ~n65528 & n55537;
  assign n55539 = pi1153 & n55427;
  assign n55540 = n54362 & n54554;
  assign n55541 = n50523 & n65461;
  assign n55542 = n54562 & ~n65531;
  assign n55543 = ~pi1152 & ~n55542;
  assign n55544 = n54535 & ~n55527;
  assign n55545 = n55543 & ~n55544;
  assign n55546 = ~pi1150 & ~n55545;
  assign n55547 = ~n55538 & n55546;
  assign n55548 = ~pi1149 & ~n55547;
  assign n55549 = ~n55522 & n55548;
  assign n55550 = ~n54794 & ~n65498;
  assign n55551 = ~pi219 & ~n55550;
  assign n55552 = ~n54451 & ~n54850;
  assign n55553 = ~pi219 & ~n54850;
  assign n55554 = ~n54451 & n55553;
  assign n55555 = ~n55550 & n55554;
  assign n55556 = n55551 & n55552;
  assign n55557 = n55132 & ~n65532;
  assign n55558 = n54496 & ~n55557;
  assign n55559 = ~n52569 & ~n54884;
  assign n55560 = ~n49599 & n65458;
  assign n55561 = ~n55559 & ~n55560;
  assign n55562 = ~pi219 & ~n55561;
  assign n55563 = n3475 & ~n54892;
  assign n55564 = ~pi57 & n55563;
  assign n55565 = n62455 & ~n54892;
  assign n55566 = ~n55562 & n65533;
  assign n55567 = n54518 & ~n55566;
  assign n55568 = pi1152 & ~n55567;
  assign n55569 = ~n55558 & n55568;
  assign n55570 = ~n54795 & ~n55125;
  assign n55571 = ~n52786 & n54446;
  assign n55572 = ~n54436 & n55477;
  assign n55573 = ~n54447 & ~n65534;
  assign n55574 = ~n55121 & n55573;
  assign n55575 = ~n55570 & ~n55574;
  assign n55576 = ~pi219 & ~n55575;
  assign n55577 = n55132 & ~n55576;
  assign n55578 = n54535 & ~n55577;
  assign n55579 = ~n54884 & ~n55427;
  assign n55580 = n62455 & ~n55579;
  assign n55581 = ~n65422 & n55580;
  assign n55582 = n54562 & ~n55581;
  assign n55583 = ~pi1152 & ~n55582;
  assign n55584 = ~n55578 & n55583;
  assign n55585 = ~pi1150 & ~n55584;
  assign n55586 = ~pi1150 & ~n55569;
  assign n55587 = ~n55584 & n55586;
  assign n55588 = ~n55569 & n55585;
  assign n55589 = n3475 & ~n54404;
  assign n55590 = ~pi57 & n55589;
  assign n55591 = n62455 & ~n54404;
  assign n55592 = ~pi299 & n54384;
  assign n55593 = ~n65324 & ~n65422;
  assign n55594 = ~n55592 & n55593;
  assign n55595 = n39342 & ~n55144;
  assign n55596 = n54915 & ~n55595;
  assign n55597 = n54915 & ~n55594;
  assign n55598 = ~n55595 & n55597;
  assign n55599 = ~n55594 & n55596;
  assign n55600 = n65536 & ~n65537;
  assign n55601 = n54518 & ~n55600;
  assign n55602 = ~pi219 & ~n54845;
  assign n55603 = ~n54850 & n55602;
  assign n55604 = ~pi1153 & n55603;
  assign n55605 = pi299 & n64625;
  assign n55606 = pi212 & n55141;
  assign n55607 = ~pi219 & ~n65538;
  assign n55608 = n55163 & ~n55607;
  assign n55609 = ~n54867 & ~n55608;
  assign n55610 = ~n55604 & ~n55609;
  assign n55611 = ~pi211 & n55603;
  assign n55612 = ~n55228 & ~n55611;
  assign n55613 = n54496 & ~n55612;
  assign n55614 = ~n55610 & n55613;
  assign n55615 = pi1152 & ~n55614;
  assign n55616 = pi1152 & ~n55601;
  assign n55617 = ~n55614 & n55616;
  assign n55618 = ~n55601 & n55615;
  assign n55619 = n54535 & ~n55610;
  assign n55620 = ~pi1151 & ~n54909;
  assign n55621 = ~pi1152 & ~n55620;
  assign n55622 = ~n55543 & ~n55621;
  assign n55623 = ~n55619 & ~n55622;
  assign n55624 = pi1150 & ~n55623;
  assign n55625 = pi1150 & ~n65539;
  assign n55626 = ~n55623 & n55625;
  assign n55627 = ~n65539 & n55624;
  assign n55628 = pi1149 & ~n65540;
  assign n55629 = ~n65535 & n55628;
  assign n55630 = ~n55522 & ~n55547;
  assign n55631 = ~pi1149 & ~n55630;
  assign n55632 = ~n55569 & ~n55584;
  assign n55633 = ~pi1150 & ~n55632;
  assign n55634 = ~n65539 & ~n55623;
  assign n55635 = pi1150 & ~n55634;
  assign n55636 = pi1149 & ~n55635;
  assign n55637 = ~n55633 & n55636;
  assign n55638 = ~n55631 & ~n55637;
  assign n55639 = ~n55549 & ~n55629;
  assign n55640 = pi213 & n65541;
  assign n55641 = ~n55206 & n55408;
  assign n55642 = ~n55223 & n55384;
  assign n55643 = pi1150 & ~n55642;
  assign n55644 = ~n55641 & n55643;
  assign n55645 = n53351 & ~n55137;
  assign n55646 = ~pi1149 & ~n55645;
  assign n55647 = ~n55644 & n55646;
  assign n55648 = ~n55133 & n55352;
  assign n55649 = ~n55167 & n55361;
  assign n55650 = ~pi1150 & ~n55649;
  assign n55651 = ~n55648 & n55650;
  assign n55652 = n55228 & n55330;
  assign n55653 = ~n55174 & n55292;
  assign n55654 = ~pi1151 & n65500;
  assign n55655 = ~n54909 & n55653;
  assign n55656 = pi1150 & ~n65542;
  assign n55657 = pi1150 & ~n55652;
  assign n55658 = ~n65542 & n55657;
  assign n55659 = ~n55652 & n55656;
  assign n55660 = pi1149 & ~n65543;
  assign n55661 = ~n55651 & n55660;
  assign n55662 = ~n55647 & ~n55661;
  assign n55663 = ~pi213 & n55662;
  assign n55664 = ~pi209 & ~n55663;
  assign n55665 = ~pi209 & ~n55640;
  assign n55666 = ~n55663 & n55665;
  assign n55667 = ~n55640 & n55664;
  assign n55668 = pi213 & ~n65541;
  assign n55669 = ~pi213 & ~n55662;
  assign n55670 = ~pi209 & ~n55669;
  assign n55671 = ~n55668 & n55670;
  assign n55672 = ~pi213 & n65522;
  assign n55673 = pi213 & ~n65470;
  assign n55674 = pi209 & ~n55673;
  assign n55675 = ~n55672 & n55674;
  assign n55676 = ~n55671 & ~n55675;
  assign n55677 = ~n55466 & ~n65544;
  assign n55678 = pi230 & n65545;
  assign n55679 = ~pi230 & ~pi241;
  assign n55680 = pi230 & ~n65545;
  assign n55681 = ~pi230 & pi241;
  assign n55682 = ~n55680 & ~n55681;
  assign n55683 = ~n55678 & ~n55679;
  assign n55684 = ~pi230 & ~pi242;
  assign n55685 = pi214 & ~n53009;
  assign n55686 = ~pi214 & ~n54763;
  assign n55687 = ~n55685 & ~n55686;
  assign n55688 = pi212 & ~n55687;
  assign n55689 = ~pi212 & n54764;
  assign n55690 = ~pi219 & ~n55689;
  assign n55691 = ~n55688 & n55690;
  assign n55692 = pi219 & ~n52525;
  assign n55693 = n52520 & ~n55692;
  assign n55694 = ~n55691 & n55693;
  assign n55695 = ~pi299 & ~n53033;
  assign n55696 = pi199 & pi1144;
  assign n55697 = ~pi200 & ~n55696;
  assign n55698 = ~n53029 & n55697;
  assign n55699 = n55695 & ~n55698;
  assign n55700 = pi207 & ~n55699;
  assign n55701 = ~n54938 & n55697;
  assign n55702 = ~pi299 & ~n54948;
  assign n55703 = ~n55701 & n55702;
  assign n55704 = ~pi207 & ~n55703;
  assign n55705 = pi208 & ~n55704;
  assign n55706 = pi208 & ~n55700;
  assign n55707 = ~n55704 & n55706;
  assign n55708 = ~n55700 & n55705;
  assign n55709 = n52555 & n55703;
  assign n55710 = ~n54784 & ~n55709;
  assign n55711 = ~n65547 & n55710;
  assign n55712 = ~pi211 & ~n55711;
  assign n55713 = ~n53272 & ~n55709;
  assign n55714 = ~n65547 & n55713;
  assign n55715 = pi211 & ~n55714;
  assign n55716 = ~n55712 & ~n55715;
  assign n55717 = ~pi214 & n55716;
  assign n55718 = ~pi211 & ~n55714;
  assign n55719 = ~n52920 & ~n55709;
  assign n55720 = ~n65547 & n55719;
  assign n55721 = pi211 & ~n55720;
  assign n55722 = pi214 & ~n55721;
  assign n55723 = pi214 & ~n55718;
  assign n55724 = ~n55721 & n55723;
  assign n55725 = ~n55718 & n55722;
  assign n55726 = pi212 & ~n65548;
  assign n55727 = pi212 & ~n55717;
  assign n55728 = ~n65548 & n55727;
  assign n55729 = ~n55717 & n55726;
  assign n55730 = n53032 & n55703;
  assign n55731 = ~pi299 & ~n55716;
  assign n55732 = ~n65547 & ~n55730;
  assign n55733 = ~pi214 & ~n65550;
  assign n55734 = ~pi212 & ~n55733;
  assign n55735 = pi214 & n55716;
  assign n55736 = n55734 & ~n55735;
  assign n55737 = ~pi219 & ~n55736;
  assign n55738 = ~n65549 & n55737;
  assign n55739 = ~n52518 & n65550;
  assign n55740 = pi219 & ~n55739;
  assign n55741 = n52518 & ~n55720;
  assign n55742 = n55740 & ~n55741;
  assign n55743 = n62455 & ~n55742;
  assign n55744 = ~n55738 & n55743;
  assign n55745 = ~n55694 & ~n55744;
  assign n55746 = pi213 & n55745;
  assign n55747 = pi211 & ~n55730;
  assign n55748 = n52518 & ~n52975;
  assign n55749 = ~n55709 & n55748;
  assign n55750 = ~n55747 & ~n55749;
  assign n55751 = pi219 & ~n55750;
  assign n55752 = n52517 & ~n55730;
  assign n55753 = pi299 & ~n65327;
  assign n55754 = n52967 & ~n55709;
  assign n55755 = n39342 & ~n52577;
  assign n55756 = ~n65324 & ~n52573;
  assign n55757 = ~n55755 & ~n55756;
  assign n55758 = ~pi219 & ~n55709;
  assign n55759 = ~n55757 & n55758;
  assign n55760 = ~n55753 & n55754;
  assign n55761 = ~n55752 & ~n65551;
  assign n55762 = ~n55751 & n55761;
  assign n55763 = ~n65547 & ~n55762;
  assign n55764 = n62455 & ~n55763;
  assign n55765 = ~pi213 & ~n52537;
  assign n55766 = ~n55764 & n55765;
  assign n55767 = ~n55746 & ~n55766;
  assign n55768 = pi209 & ~n55767;
  assign n55769 = ~pi213 & ~n52603;
  assign n55770 = ~n52517 & n52525;
  assign n55771 = pi219 & n52517;
  assign n55772 = ~n55692 & ~n55771;
  assign n55773 = pi219 & ~n55770;
  assign n55774 = ~n55691 & n65552;
  assign n55775 = pi299 & ~n55774;
  assign n55776 = n62455 & ~n55775;
  assign n55777 = pi299 & n65552;
  assign n55778 = ~n55691 & n55777;
  assign n55779 = ~n52558 & ~n55778;
  assign n55780 = n62455 & ~n55779;
  assign n55781 = ~n52592 & n55776;
  assign n55782 = ~n55694 & ~n65553;
  assign n55783 = pi213 & ~n55782;
  assign n55784 = ~pi209 & ~n55783;
  assign n55785 = ~pi209 & ~n55769;
  assign n55786 = ~n55783 & n55785;
  assign n55787 = ~n55769 & n55784;
  assign n55788 = ~n55768 & ~n65554;
  assign n55789 = pi230 & ~n55788;
  assign po399 = ~n55684 & ~n55789;
  assign n55791 = ~pi230 & ~pi244;
  assign n55792 = pi213 & ~n55018;
  assign n55793 = ~n52918 & n54956;
  assign n55794 = ~n54994 & ~n55793;
  assign n55795 = ~pi214 & n55794;
  assign n55796 = n52526 & n54855;
  assign n55797 = pi212 & ~n55796;
  assign n55798 = ~n55795 & n55797;
  assign n55799 = ~n55022 & n55798;
  assign n55800 = ~n55022 & ~n55794;
  assign n55801 = pi214 & ~n55800;
  assign n55802 = n54984 & ~n55801;
  assign n55803 = ~pi219 & ~n55802;
  assign n55804 = ~pi219 & ~n55799;
  assign n55805 = ~n55802 & n55804;
  assign n55806 = ~n55799 & n55803;
  assign n55807 = ~pi211 & ~n52881;
  assign n55808 = ~n65490 & n55807;
  assign n55809 = ~n55008 & ~n55808;
  assign n55810 = n55006 & ~n55809;
  assign n55811 = n65497 & ~n55810;
  assign n55812 = ~n65555 & n55811;
  assign n55813 = ~n54955 & n55798;
  assign n55814 = pi214 & n55794;
  assign n55815 = n54972 & ~n55814;
  assign n55816 = ~pi219 & ~n55815;
  assign n55817 = ~n55813 & n55816;
  assign n55818 = pi299 & n53019;
  assign n55819 = pi1147 & ~n55818;
  assign n55820 = n55046 & n55819;
  assign n55821 = ~n55817 & n55820;
  assign n55822 = ~pi213 & ~n53021;
  assign n55823 = ~n55821 & n55822;
  assign n55824 = ~n55812 & n55823;
  assign n55825 = ~n55792 & ~n55824;
  assign n55826 = ~n53021 & ~n55821;
  assign n55827 = ~n55812 & n55826;
  assign n55828 = ~pi213 & ~n55827;
  assign n55829 = pi213 & n55018;
  assign n55830 = pi209 & ~n55829;
  assign n55831 = ~n55828 & n55830;
  assign n55832 = pi209 & ~n55825;
  assign n55833 = ~n54776 & ~n54811;
  assign n55834 = n54806 & ~n54808;
  assign n55835 = n39342 & ~n54789;
  assign n55836 = ~n39342 & n54911;
  assign n55837 = n52967 & ~n55836;
  assign n55838 = n52967 & ~n55835;
  assign n55839 = ~n55836 & n55838;
  assign n55840 = ~n55835 & n55837;
  assign n55841 = ~n55834 & n65557;
  assign n55842 = ~n53037 & ~n65485;
  assign n55843 = ~n55841 & n55842;
  assign n55844 = n62455 & ~n55843;
  assign n55845 = ~n55833 & ~n55844;
  assign n55846 = pi213 & ~n55845;
  assign n55847 = ~pi213 & ~n53049;
  assign n55848 = ~pi209 & ~n55847;
  assign n55849 = ~n55846 & n55848;
  assign n55850 = ~n65556 & ~n55849;
  assign n55851 = pi230 & ~n55850;
  assign po401 = ~n55791 & ~n55851;
  assign n55853 = pi1146 & n54494;
  assign n55854 = pi1147 & ~n54485;
  assign n55855 = ~n55853 & n55854;
  assign n55856 = ~n55069 & ~n55855;
  assign n55857 = ~n52517 & n55712;
  assign n55858 = n52518 & ~n55711;
  assign n55859 = n55740 & ~n65558;
  assign n55860 = n62455 & ~n55859;
  assign n55861 = ~pi299 & n55714;
  assign n55862 = ~pi211 & ~n55861;
  assign n55863 = pi211 & ~n55711;
  assign n55864 = ~n55862 & ~n55863;
  assign n55865 = pi214 & ~n55864;
  assign n55866 = ~n48494 & ~n65550;
  assign n55867 = ~pi214 & ~n55866;
  assign n55868 = ~n55865 & ~n55867;
  assign n55869 = pi212 & ~n55868;
  assign n55870 = n55734 & ~n55866;
  assign n55871 = ~pi219 & ~n55870;
  assign n55872 = ~n55869 & n55871;
  assign n55873 = n55860 & ~n55872;
  assign n55874 = ~n55856 & ~n55873;
  assign n55875 = ~pi1147 & ~n55853;
  assign n55876 = pi214 & ~n54836;
  assign n55877 = ~n65550 & n55876;
  assign n55878 = pi212 & ~n55877;
  assign n55879 = ~n55733 & n55878;
  assign n55880 = ~pi212 & n65550;
  assign n55881 = ~pi219 & ~n55880;
  assign n55882 = ~n55879 & n55881;
  assign n55883 = n55860 & ~n55882;
  assign n55884 = n55875 & ~n55883;
  assign n55885 = ~pi1148 & ~n55884;
  assign n55886 = ~pi1148 & ~n55874;
  assign n55887 = ~n55884 & n55886;
  assign n55888 = ~n55874 & n55885;
  assign n55889 = ~pi214 & ~n55861;
  assign n55890 = ~n55865 & ~n55889;
  assign n55891 = pi212 & ~n55890;
  assign n55892 = n55734 & ~n55861;
  assign n55893 = ~pi219 & ~n55892;
  assign n55894 = ~n55891 & n55893;
  assign n55895 = n55860 & ~n55894;
  assign n55896 = n55855 & ~n55895;
  assign n55897 = ~n65464 & n55875;
  assign n55898 = ~n65550 & ~n55862;
  assign n55899 = ~pi214 & n55898;
  assign n55900 = n55878 & ~n55899;
  assign n55901 = n55734 & ~n55898;
  assign n55902 = ~pi219 & ~n55901;
  assign n55903 = ~n55900 & n55902;
  assign n55904 = n55860 & ~n55903;
  assign n55905 = n55897 & ~n55904;
  assign n55906 = pi1148 & ~n55905;
  assign n55907 = pi1148 & ~n55896;
  assign n55908 = ~n55905 & n55907;
  assign n55909 = ~n55896 & n55906;
  assign n55910 = ~n55896 & ~n55905;
  assign n55911 = pi1148 & ~n55910;
  assign n55912 = ~n55874 & ~n55884;
  assign n55913 = ~pi1148 & ~n55912;
  assign n55914 = ~n55911 & ~n55913;
  assign n55915 = ~n65559 & ~n65560;
  assign n55916 = pi213 & n65561;
  assign n55917 = ~pi213 & ~n55745;
  assign n55918 = ~pi209 & ~n55917;
  assign n55919 = ~n55916 & n55918;
  assign n55920 = pi199 & pi1146;
  assign n55921 = ~pi200 & ~n55920;
  assign n55922 = n54940 & ~n55921;
  assign n55923 = pi207 & n55922;
  assign n55924 = pi1146 & ~n49519;
  assign n55925 = ~n55923 & ~n55924;
  assign n55926 = pi208 & ~n55925;
  assign n55927 = n49457 & ~n55920;
  assign n55928 = n54940 & ~n55927;
  assign n55929 = pi208 & n55928;
  assign n55930 = ~pi207 & ~n55929;
  assign n55931 = n54410 & ~n55927;
  assign n55932 = ~n55930 & n55931;
  assign n55933 = n65452 & ~n55927;
  assign n55934 = ~n55926 & ~n65562;
  assign n55935 = ~pi208 & n54784;
  assign n55936 = ~n65562 & ~n55935;
  assign n55937 = n55934 & ~n55935;
  assign n55938 = ~n55926 & ~n55935;
  assign n55939 = ~n65562 & n55938;
  assign n55940 = ~n55926 & n55936;
  assign n55941 = ~pi299 & ~n65563;
  assign n55942 = ~pi299 & ~n55934;
  assign n55943 = ~pi214 & ~n65564;
  assign n55944 = ~pi212 & ~n55943;
  assign n55945 = ~n38985 & ~n65452;
  assign n55946 = n55922 & ~n55945;
  assign n55947 = pi211 & ~n55946;
  assign n55948 = ~pi299 & ~n55922;
  assign n55949 = ~n65563 & ~n55948;
  assign n55950 = ~pi299 & ~n55949;
  assign n55951 = ~pi211 & n55950;
  assign n55952 = ~n55947 & ~n55951;
  assign n55953 = ~n65564 & ~n55952;
  assign n55954 = n55944 & ~n55953;
  assign n55955 = ~pi219 & ~n55954;
  assign n55956 = n55876 & ~n65564;
  assign n55957 = ~pi214 & n55953;
  assign n55958 = pi212 & ~n55957;
  assign n55959 = ~n55956 & n55958;
  assign n55960 = n55955 & ~n55959;
  assign n55961 = ~n52518 & n65564;
  assign n55962 = pi219 & ~n55961;
  assign n55963 = n52518 & ~n65563;
  assign n55964 = n55962 & ~n55963;
  assign n55965 = n62455 & ~n55964;
  assign n55966 = ~n55960 & n55965;
  assign n55967 = n55897 & ~n55966;
  assign n55968 = ~pi1146 & ~n54357;
  assign n55969 = n49595 & ~n55927;
  assign n55970 = ~n38985 & ~n55969;
  assign n55971 = pi207 & ~n55927;
  assign n55972 = pi207 & n55928;
  assign n55973 = n54940 & n55971;
  assign n55974 = ~n53032 & ~n65565;
  assign n55975 = ~n55970 & ~n55974;
  assign n55976 = n49595 & ~n55921;
  assign n55977 = ~pi207 & n55976;
  assign n55978 = ~n54784 & ~n65565;
  assign n55979 = ~n54784 & ~n55977;
  assign n55980 = ~n65565 & n55979;
  assign n55981 = ~n55977 & n55978;
  assign n55982 = pi208 & ~n65567;
  assign n55983 = ~pi299 & n55982;
  assign n55984 = n52555 & n55969;
  assign n55985 = ~n55929 & ~n55984;
  assign n55986 = ~n55983 & n55985;
  assign n55987 = n54845 & ~n55968;
  assign n55988 = ~pi214 & ~n65566;
  assign n55989 = ~pi212 & ~n55988;
  assign n55990 = ~pi299 & ~n65566;
  assign n55991 = n55989 & ~n55990;
  assign n55992 = ~pi219 & ~n55991;
  assign n55993 = pi212 & ~n55990;
  assign n55994 = ~n54784 & ~n65566;
  assign n55995 = n39343 & n55994;
  assign n55996 = n55993 & ~n55995;
  assign n55997 = n55992 & ~n55996;
  assign n55998 = ~n52518 & n65566;
  assign n55999 = pi219 & ~n55998;
  assign n56000 = n52518 & ~n55994;
  assign n56001 = n55999 & ~n56000;
  assign n56002 = n62455 & ~n56001;
  assign n56003 = ~n55997 & n56002;
  assign n56004 = n55855 & ~n56003;
  assign n56005 = pi1148 & ~n56004;
  assign n56006 = ~n55967 & n56005;
  assign n56007 = ~n38985 & ~n55976;
  assign n56008 = ~n55974 & ~n56007;
  assign n56009 = ~n48494 & ~n56008;
  assign n56010 = pi214 & ~n56009;
  assign n56011 = ~pi214 & n56008;
  assign n56012 = ~pi212 & ~n56011;
  assign n56013 = ~n56010 & n56012;
  assign n56014 = ~pi214 & ~n56009;
  assign n56015 = n52555 & n55976;
  assign n56016 = ~n55982 & ~n56015;
  assign n56017 = ~n55935 & ~n56015;
  assign n56018 = ~n55935 & n56016;
  assign n56019 = ~n55982 & n56017;
  assign n56020 = ~pi299 & n65568;
  assign n56021 = ~pi299 & n56016;
  assign n56022 = pi214 & ~n65569;
  assign n56023 = ~pi211 & ~n55990;
  assign n56024 = ~n65566 & ~n56023;
  assign n56025 = n56022 & ~n56024;
  assign n56026 = pi212 & ~n56025;
  assign n56027 = ~n56014 & n56026;
  assign n56028 = ~n56013 & ~n56027;
  assign n56029 = ~pi219 & ~n56028;
  assign n56030 = ~pi1146 & ~n52855;
  assign n56031 = n54850 & ~n56030;
  assign n56032 = n56029 & ~n56031;
  assign n56033 = ~n52517 & n56008;
  assign n56034 = ~n52518 & ~n56033;
  assign n56035 = ~n65568 & ~n56034;
  assign n56036 = ~pi212 & n56011;
  assign n56037 = pi219 & ~n56036;
  assign n56038 = ~n56035 & n56037;
  assign n56039 = n62455 & ~n56038;
  assign n56040 = ~n56032 & n56039;
  assign n56041 = ~n55856 & ~n56040;
  assign n56042 = ~n65538 & ~n65564;
  assign n56043 = ~n55925 & ~n56042;
  assign n56044 = ~pi219 & ~n56043;
  assign n56045 = pi219 & ~n55946;
  assign n56046 = ~n53038 & ~n56045;
  assign n56047 = ~n52517 & ~n55947;
  assign n56048 = n55949 & n56047;
  assign n56049 = ~n56046 & ~n56048;
  assign n56050 = n62455 & ~n56049;
  assign n56051 = ~n56044 & n56050;
  assign n56052 = n55875 & ~n56051;
  assign n56053 = ~pi1148 & ~n56052;
  assign n56054 = ~n56041 & n56053;
  assign n56055 = ~n56006 & ~n56054;
  assign n56056 = pi213 & ~n56055;
  assign n56057 = ~pi214 & n55946;
  assign n56058 = ~n54789 & ~n65564;
  assign n56059 = pi214 & ~n55950;
  assign n56060 = ~n56058 & n56059;
  assign n56061 = ~n56057 & ~n56060;
  assign n56062 = ~pi212 & ~n56061;
  assign n56063 = pi299 & ~n55687;
  assign n56064 = ~n65564 & ~n56063;
  assign n56065 = pi212 & ~n56064;
  assign n56066 = ~n55948 & n56065;
  assign n56067 = ~pi219 & ~n56066;
  assign n56068 = ~n56062 & n56067;
  assign n56069 = ~n52918 & ~n55950;
  assign n56070 = ~pi211 & ~n56069;
  assign n56071 = n56047 & ~n56070;
  assign n56072 = ~n56046 & ~n56071;
  assign n56073 = n65497 & ~n56072;
  assign n56074 = ~n56068 & n56073;
  assign n56075 = ~n54789 & ~n65566;
  assign n56076 = n56022 & ~n56075;
  assign n56077 = ~n56011 & ~n56076;
  assign n56078 = ~pi212 & ~n56077;
  assign n56079 = ~n65566 & ~n56063;
  assign n56080 = pi212 & ~n56079;
  assign n56081 = ~n65569 & n56080;
  assign n56082 = ~pi219 & ~n56081;
  assign n56083 = ~n56078 & n56082;
  assign n56084 = ~pi57 & pi1147;
  assign n56085 = pi1147 & n62455;
  assign n56086 = n3475 & n56084;
  assign n56087 = ~n52920 & ~n65566;
  assign n56088 = ~n65569 & ~n56087;
  assign n56089 = ~pi211 & ~n56088;
  assign n56090 = ~n56034 & ~n56089;
  assign n56091 = n56037 & ~n56090;
  assign n56092 = n65570 & ~n56091;
  assign n56093 = ~n56083 & n65570;
  assign n56094 = ~n56091 & n56093;
  assign n56095 = ~n56083 & n56092;
  assign n56096 = ~pi1148 & ~n55694;
  assign n56097 = ~n65571 & n56096;
  assign n56098 = ~n56074 & n56097;
  assign n56099 = n55944 & ~n56058;
  assign n56100 = ~pi219 & ~n56065;
  assign n56101 = ~n56099 & n56100;
  assign n56102 = ~pi299 & n65563;
  assign n56103 = ~pi299 & n55934;
  assign n56104 = n52518 & ~n65572;
  assign n56105 = ~n52918 & n56104;
  assign n56106 = n55962 & ~n56105;
  assign n56107 = n65497 & ~n56106;
  assign n56108 = ~n56101 & n56107;
  assign n56109 = pi214 & n56075;
  assign n56110 = n55989 & ~n56109;
  assign n56111 = ~pi219 & ~n56080;
  assign n56112 = ~n56110 & n56111;
  assign n56113 = n52518 & ~n56087;
  assign n56114 = n55999 & ~n56113;
  assign n56115 = n65570 & ~n56114;
  assign n56116 = ~n56112 & n56115;
  assign n56117 = pi1148 & ~n55694;
  assign n56118 = ~n56116 & n56117;
  assign n56119 = ~n56108 & n56118;
  assign n56120 = ~pi213 & ~n56119;
  assign n56121 = ~n56098 & n56120;
  assign n56122 = pi209 & ~n56121;
  assign n56123 = ~n56056 & n56122;
  assign n56124 = pi213 & ~n65561;
  assign n56125 = ~pi213 & n55745;
  assign n56126 = ~pi209 & ~n56125;
  assign n56127 = ~n56124 & n56126;
  assign n56128 = pi213 & n56055;
  assign n56129 = ~n56098 & ~n56119;
  assign n56130 = ~pi213 & ~n56129;
  assign n56131 = pi209 & ~n56130;
  assign n56132 = ~n56128 & n56131;
  assign n56133 = ~n56127 & ~n56132;
  assign n56134 = ~n55919 & ~n56123;
  assign n56135 = pi230 & n65573;
  assign n56136 = ~pi230 & ~pi245;
  assign n56137 = pi230 & ~n65573;
  assign n56138 = ~pi230 & pi245;
  assign n56139 = ~n56137 & ~n56138;
  assign n56140 = ~n56135 & ~n56136;
  assign n56141 = ~pi209 & n56055;
  assign n56142 = pi219 & ~n54784;
  assign n56143 = n54777 & ~n56142;
  assign n56144 = ~n54782 & ~n56143;
  assign n56145 = ~n54796 & n55386;
  assign n56146 = ~pi212 & ~n65453;
  assign n56147 = ~pi219 & ~n56146;
  assign n56148 = ~n55306 & n56147;
  assign n56149 = ~n56145 & n56148;
  assign n56150 = ~n56144 & ~n56149;
  assign n56151 = n55855 & ~n56150;
  assign n56152 = ~n54786 & n55117;
  assign n56153 = ~pi214 & n54448;
  assign n56154 = pi212 & ~n56153;
  assign n56155 = ~n56152 & n56154;
  assign n56156 = n55124 & ~n56155;
  assign n56157 = ~n56144 & ~n56156;
  assign n56158 = n55897 & ~n56157;
  assign n56159 = ~n56151 & ~n56158;
  assign n56160 = pi1150 & ~n56159;
  assign n56161 = ~n55152 & ~n55161;
  assign n56162 = n55897 & ~n56161;
  assign n56163 = ~n54883 & n54909;
  assign n56164 = ~n56143 & ~n56163;
  assign n56165 = n65324 & n54878;
  assign n56166 = ~n54878 & ~n54885;
  assign n56167 = n65324 & ~n56166;
  assign n56168 = ~n55559 & ~n56167;
  assign n56169 = ~n55559 & ~n56165;
  assign n56170 = ~pi219 & ~n65575;
  assign n56171 = ~n56164 & ~n56170;
  assign n56172 = ~n56162 & n56171;
  assign n56173 = ~n55855 & ~n55897;
  assign n56174 = ~pi1150 & ~n56173;
  assign n56175 = ~n56172 & n56174;
  assign n56176 = pi1148 & ~n56175;
  assign n56177 = ~n56171 & ~n56173;
  assign n56178 = ~pi1150 & ~n56162;
  assign n56179 = ~n56177 & n56178;
  assign n56180 = pi1150 & ~n56158;
  assign n56181 = ~n56151 & n56180;
  assign n56182 = ~n56179 & ~n56181;
  assign n56183 = pi1148 & ~n56182;
  assign n56184 = ~n56160 & n56176;
  assign n56185 = ~pi219 & ~n54765;
  assign n56186 = ~n55607 & ~n56185;
  assign n56187 = n56143 & n56186;
  assign n56188 = n55875 & ~n56187;
  assign n56189 = ~n55856 & ~n56143;
  assign n56190 = ~n56188 & ~n56189;
  assign n56191 = pi1150 & n65476;
  assign n56192 = ~n56190 & ~n56191;
  assign n56193 = pi1150 & n54388;
  assign n56194 = pi299 & n52911;
  assign n56195 = ~pi219 & ~n56194;
  assign n56196 = ~n56031 & n56195;
  assign n56197 = ~n56193 & n56196;
  assign n56198 = ~n55856 & n56197;
  assign n56199 = ~pi1148 & ~n56198;
  assign n56200 = ~n56192 & n56199;
  assign n56201 = ~n65576 & ~n56200;
  assign n56202 = ~pi1149 & ~n56201;
  assign n56203 = n54765 & n54855;
  assign n56204 = ~n54906 & ~n56203;
  assign n56205 = n55203 & n56204;
  assign n56206 = n54777 & ~n55184;
  assign n56207 = ~n55205 & ~n56206;
  assign n56208 = ~pi1146 & n55204;
  assign n56209 = ~n56207 & ~n56208;
  assign n56210 = ~n56205 & n56209;
  assign n56211 = ~n55856 & ~n56210;
  assign n56212 = ~n55181 & ~n55305;
  assign n56213 = ~pi219 & ~n56212;
  assign n56214 = ~n56207 & ~n56213;
  assign n56215 = ~pi1146 & ~n54906;
  assign n56216 = n56214 & ~n56215;
  assign n56217 = n55875 & ~n56216;
  assign n56218 = ~pi1150 & ~n56217;
  assign n56219 = ~n56211 & n56218;
  assign n56220 = ~pi214 & n55494;
  assign n56221 = n55220 & ~n56220;
  assign n56222 = ~pi219 & ~n56221;
  assign n56223 = ~n54834 & ~n55494;
  assign n56224 = ~pi212 & n56223;
  assign n56225 = n56222 & ~n56224;
  assign n56226 = ~pi299 & n54332;
  assign n56227 = ~n54784 & ~n54817;
  assign n56228 = ~n56226 & n56227;
  assign n56229 = n56225 & n56228;
  assign n56230 = ~n65479 & ~n56143;
  assign n56231 = n56222 & ~n56223;
  assign n56232 = ~n56230 & ~n56231;
  assign n56233 = ~n56229 & n56232;
  assign n56234 = n54835 & ~n55219;
  assign n56235 = ~pi219 & ~n65525;
  assign n56236 = ~pi219 & ~n56234;
  assign n56237 = ~n65525 & n56236;
  assign n56238 = ~n56234 & n56235;
  assign n56239 = n54827 & ~n65577;
  assign n56240 = n56233 & n56239;
  assign n56241 = n55875 & ~n56240;
  assign n56242 = ~n55856 & ~n56233;
  assign n56243 = pi1150 & ~n56242;
  assign n56244 = ~n56241 & n56243;
  assign n56245 = ~pi1148 & ~n56244;
  assign n56246 = pi1150 & n56239;
  assign n56247 = n56233 & n56246;
  assign n56248 = ~pi1150 & ~n56215;
  assign n56249 = n56214 & n56248;
  assign n56250 = n55875 & ~n56249;
  assign n56251 = ~n56247 & n56250;
  assign n56252 = ~pi1150 & ~n56208;
  assign n56253 = ~n56207 & n56252;
  assign n56254 = ~n56205 & n56253;
  assign n56255 = pi1150 & n56233;
  assign n56256 = ~n55856 & ~n56255;
  assign n56257 = ~n56254 & n56256;
  assign n56258 = ~n56251 & ~n56257;
  assign n56259 = ~pi1148 & ~n56258;
  assign n56260 = ~n56219 & n56245;
  assign n56261 = ~n54909 & ~n56143;
  assign n56262 = ~n55144 & n55160;
  assign n56263 = ~n55150 & ~n56262;
  assign n56264 = ~n55897 & ~n56263;
  assign n56265 = n54384 & n55876;
  assign n56266 = n55158 & ~n56265;
  assign n56267 = n55156 & ~n56266;
  assign n56268 = ~n56264 & n56267;
  assign n56269 = ~n56261 & ~n56268;
  assign n56270 = ~n56173 & ~n56269;
  assign n56271 = ~pi1150 & ~n56270;
  assign n56272 = ~n54867 & ~n56187;
  assign n56273 = ~n65464 & ~n54867;
  assign n56274 = n56188 & n56273;
  assign n56275 = n55897 & n56272;
  assign n56276 = ~n54845 & ~n65529;
  assign n56277 = pi214 & n54858;
  assign n56278 = n54852 & ~n56277;
  assign n56279 = ~pi219 & ~n54860;
  assign n56280 = ~n56278 & n56279;
  assign n56281 = n54847 & ~n56280;
  assign n56282 = n62455 & ~n56276;
  assign n56283 = pi1146 & n55173;
  assign n56284 = ~n65580 & ~n56283;
  assign n56285 = n55855 & ~n56283;
  assign n56286 = ~n65580 & n56285;
  assign n56287 = n55855 & n56284;
  assign n56288 = pi1150 & ~n65581;
  assign n56289 = ~n65579 & n56288;
  assign n56290 = pi1148 & ~n56289;
  assign n56291 = ~n56271 & n56290;
  assign n56292 = pi1149 & ~n56291;
  assign n56293 = ~n65578 & n56292;
  assign n56294 = ~n56271 & ~n56289;
  assign n56295 = pi1148 & ~n56294;
  assign n56296 = ~pi1148 & ~n56257;
  assign n56297 = ~n56251 & n56296;
  assign n56298 = pi1149 & ~n56297;
  assign n56299 = ~n65578 & ~n56291;
  assign n56300 = pi1149 & ~n56299;
  assign n56301 = ~n56295 & n56298;
  assign n56302 = ~pi1149 & ~n56200;
  assign n56303 = ~n65576 & n56302;
  assign n56304 = ~n65582 & ~n56303;
  assign n56305 = ~n56202 & ~n56293;
  assign n56306 = pi209 & ~n65583;
  assign n56307 = ~pi213 & ~n56306;
  assign n56308 = ~n56141 & n56307;
  assign n56309 = ~pi212 & ~n56057;
  assign n56310 = ~n48494 & ~n55946;
  assign n56311 = pi214 & ~n56310;
  assign n56312 = n56309 & ~n56311;
  assign n56313 = pi214 & n55952;
  assign n56314 = pi212 & ~n56313;
  assign n56315 = ~pi214 & ~n56310;
  assign n56316 = n56314 & ~n56315;
  assign n56317 = ~n56312 & ~n56316;
  assign n56318 = ~pi219 & ~n56317;
  assign n56319 = n65497 & ~n56045;
  assign n56320 = ~n56318 & n56319;
  assign n56321 = ~pi1150 & ~n55056;
  assign n56322 = pi219 & ~n56008;
  assign n56323 = n65570 & ~n56322;
  assign n56324 = ~n56029 & n56323;
  assign n56325 = n56321 & ~n56324;
  assign n56326 = ~n56320 & n56325;
  assign n56327 = ~n56059 & n56309;
  assign n56328 = ~pi214 & ~n55950;
  assign n56329 = n56314 & ~n56328;
  assign n56330 = ~n56327 & ~n56329;
  assign n56331 = ~pi219 & ~n56330;
  assign n56332 = ~n56045 & ~n56331;
  assign n56333 = ~pi1147 & ~n56332;
  assign n56334 = n56012 & ~n56022;
  assign n56335 = ~pi214 & ~n65569;
  assign n56336 = n56026 & ~n56335;
  assign n56337 = ~n56334 & ~n56336;
  assign n56338 = ~pi219 & ~n56337;
  assign n56339 = ~n56322 & ~n56338;
  assign n56340 = pi1147 & ~n56339;
  assign n56341 = n62455 & ~n56340;
  assign n56342 = ~n56333 & n56341;
  assign n56343 = pi1150 & ~n54485;
  assign n56344 = ~n56342 & n56343;
  assign n56345 = ~n56326 & ~n56344;
  assign n56346 = pi1149 & ~n56345;
  assign n56347 = pi1150 & n65463;
  assign n56348 = ~pi1147 & n55949;
  assign n56349 = n65014 & ~n56348;
  assign n56350 = n56347 & ~n56349;
  assign n56351 = pi1147 & ~n56008;
  assign n56352 = n55946 & ~n56347;
  assign n56353 = ~pi1147 & ~n56352;
  assign n56354 = n62455 & ~n56353;
  assign n56355 = ~n56351 & n56354;
  assign n56356 = ~pi1149 & ~n56355;
  assign n56357 = ~n56350 & n56356;
  assign n56358 = ~pi1148 & ~n56357;
  assign n56359 = ~n56346 & n56358;
  assign n56360 = n55962 & ~n56104;
  assign n56361 = n65497 & ~n56360;
  assign n56362 = ~pi219 & n56042;
  assign n56363 = n55607 & ~n65564;
  assign n56364 = n56361 & ~n65584;
  assign n56365 = ~n52517 & n56023;
  assign n56366 = n55999 & ~n56365;
  assign n56367 = n3475 & ~n56366;
  assign n56368 = n56084 & n56367;
  assign n56369 = n65570 & ~n56366;
  assign n56370 = pi214 & ~n48494;
  assign n56371 = ~n65566 & n56370;
  assign n56372 = pi212 & ~n56371;
  assign n56373 = ~n55988 & n56372;
  assign n56374 = ~pi212 & n65566;
  assign n56375 = ~pi219 & ~n56374;
  assign n56376 = ~n56373 & n56375;
  assign n56377 = n65585 & ~n56376;
  assign n56378 = ~pi1150 & ~n54494;
  assign n56379 = ~n56377 & n56378;
  assign n56380 = ~n56364 & n56378;
  assign n56381 = ~n56377 & n56380;
  assign n56382 = ~n56364 & n56379;
  assign n56383 = pi214 & n56310;
  assign n56384 = ~n65564 & n56310;
  assign n56385 = pi214 & n56384;
  assign n56386 = ~n65564 & n56383;
  assign n56387 = n55958 & ~n65587;
  assign n56388 = n55955 & ~n56387;
  assign n56389 = n56361 & ~n56388;
  assign n56390 = ~pi214 & n56024;
  assign n56391 = n56372 & ~n56390;
  assign n56392 = n55989 & ~n56024;
  assign n56393 = ~pi219 & ~n56392;
  assign n56394 = ~pi219 & ~n56391;
  assign n56395 = ~n56392 & n56394;
  assign n56396 = ~n56391 & n56393;
  assign n56397 = n65585 & ~n65588;
  assign n56398 = pi1150 & ~n55100;
  assign n56399 = ~n56397 & n56398;
  assign n56400 = ~n56389 & n56399;
  assign n56401 = ~n65586 & ~n56400;
  assign n56402 = ~pi1149 & ~n56401;
  assign n56403 = n39342 & ~n55950;
  assign n56404 = ~n52517 & ~n56310;
  assign n56405 = ~pi219 & ~n56404;
  assign n56406 = ~n65564 & n56405;
  assign n56407 = ~n56059 & n56384;
  assign n56408 = pi212 & ~n56407;
  assign n56409 = n55944 & ~n65587;
  assign n56410 = ~pi219 & ~n56409;
  assign n56411 = ~n56408 & n56410;
  assign n56412 = ~n56403 & n56406;
  assign n56413 = n56361 & ~n65589;
  assign n56414 = n55992 & ~n55993;
  assign n56415 = ~n56366 & ~n56414;
  assign n56416 = n3475 & n56415;
  assign n56417 = n56367 & ~n56414;
  assign n56418 = ~n55611 & n56084;
  assign n56419 = ~n55611 & n65570;
  assign n56420 = n56415 & n56419;
  assign n56421 = n65590 & n56418;
  assign n56422 = ~n55068 & ~n65591;
  assign n56423 = ~n56413 & n56422;
  assign n56424 = ~pi1150 & ~n56423;
  assign n56425 = ~n3475 & ~n52968;
  assign n56426 = n56084 & ~n56425;
  assign n56427 = ~n65590 & n56426;
  assign n56428 = n62455 & n65572;
  assign n56429 = ~n47803 & n52968;
  assign n56430 = ~n56428 & ~n56429;
  assign n56431 = ~pi1147 & ~n56430;
  assign n56432 = pi57 & n52968;
  assign n56433 = pi1150 & ~n56432;
  assign n56434 = n3475 & ~n52967;
  assign n56435 = n55961 & n56434;
  assign n56436 = ~n52968 & ~n65572;
  assign n56437 = n55094 & ~n56425;
  assign n56438 = ~n56436 & n56437;
  assign n56439 = ~n56435 & n56438;
  assign n56440 = n56433 & ~n56439;
  assign n56441 = ~n56431 & n56433;
  assign n56442 = ~n56427 & n65592;
  assign n56443 = pi1149 & ~n56442;
  assign n56444 = ~n56424 & n56443;
  assign n56445 = pi1148 & ~n56444;
  assign n56446 = ~n56402 & n56445;
  assign n56447 = ~pi209 & ~n56446;
  assign n56448 = ~n56359 & n56447;
  assign n56449 = n53390 & ~n55137;
  assign n56450 = ~pi1150 & n55207;
  assign n56451 = ~n55206 & n56321;
  assign n56452 = pi1150 & n55224;
  assign n56453 = pi1149 & ~n56452;
  assign n56454 = ~n65593 & n56453;
  assign n56455 = ~n56449 & ~n56454;
  assign n56456 = ~pi1148 & ~n56455;
  assign n56457 = pi1150 & ~n55134;
  assign n56458 = ~pi1150 & ~n55168;
  assign n56459 = ~pi1149 & ~n56458;
  assign n56460 = ~n56457 & n56459;
  assign n56461 = ~pi1150 & ~n65500;
  assign n56462 = pi1150 & ~n55229;
  assign n56463 = pi1149 & ~n56462;
  assign n56464 = ~n56461 & n56463;
  assign n56465 = pi1148 & ~n56464;
  assign n56466 = ~pi1150 & n65500;
  assign n56467 = pi1150 & n55229;
  assign n56468 = pi1149 & ~n56467;
  assign n56469 = pi1149 & ~n56466;
  assign n56470 = ~n56467 & n56469;
  assign n56471 = ~n56466 & n56468;
  assign n56472 = pi1150 & n55134;
  assign n56473 = ~pi1150 & n55168;
  assign n56474 = ~pi1149 & ~n56473;
  assign n56475 = ~n56472 & n56474;
  assign n56476 = ~n65594 & ~n56475;
  assign n56477 = pi1148 & ~n56476;
  assign n56478 = ~n56460 & n56465;
  assign n56479 = ~n56456 & ~n65595;
  assign n56480 = pi209 & n56479;
  assign n56481 = pi213 & ~n56480;
  assign n56482 = ~n56448 & n56481;
  assign n56483 = ~pi213 & ~n56303;
  assign n56484 = ~pi213 & n65583;
  assign n56485 = ~n65582 & n56483;
  assign n56486 = pi213 & ~n56479;
  assign n56487 = pi209 & ~n56486;
  assign n56488 = pi209 & ~n65596;
  assign n56489 = ~n56486 & n56488;
  assign n56490 = ~n65596 & n56487;
  assign n56491 = ~n56359 & ~n56446;
  assign n56492 = ~n56346 & ~n56357;
  assign n56493 = ~pi1148 & ~n56492;
  assign n56494 = ~pi1149 & ~n65586;
  assign n56495 = ~n56400 & n56494;
  assign n56496 = ~n56432 & ~n56439;
  assign n56497 = ~n56427 & n56496;
  assign n56498 = pi1150 & ~n56497;
  assign n56499 = ~pi1150 & ~n55068;
  assign n56500 = ~n65591 & n56499;
  assign n56501 = ~n56413 & n56500;
  assign n56502 = pi1149 & ~n56501;
  assign n56503 = pi1149 & ~n56498;
  assign n56504 = ~n56501 & n56503;
  assign n56505 = ~n56498 & n56502;
  assign n56506 = pi1148 & ~n65598;
  assign n56507 = ~n56495 & n56506;
  assign n56508 = pi213 & ~n56507;
  assign n56509 = ~n56493 & n56508;
  assign n56510 = pi213 & ~n56491;
  assign n56511 = ~pi213 & ~n56055;
  assign n56512 = ~pi209 & ~n56511;
  assign n56513 = ~n65599 & n56512;
  assign n56514 = ~n65597 & ~n56513;
  assign n56515 = ~n56308 & ~n56482;
  assign n56516 = pi230 & ~n65600;
  assign n56517 = ~pi230 & ~pi246;
  assign n56518 = pi230 & n65600;
  assign n56519 = ~pi230 & pi246;
  assign n56520 = ~n56518 & ~n56519;
  assign n56521 = ~n56516 & ~n56517;
  assign n56522 = pi1147 & ~n55648;
  assign n56523 = ~pi1151 & ~n55100;
  assign n56524 = ~n55166 & n56523;
  assign n56525 = n56522 & ~n56524;
  assign n56526 = pi1151 & ~n65464;
  assign n56527 = n54782 & ~n55127;
  assign n56528 = ~n65464 & ~n56527;
  assign n56529 = pi1151 & n56528;
  assign n56530 = n56526 & ~n56527;
  assign n56531 = ~pi1151 & ~n65464;
  assign n56532 = ~n55580 & n56531;
  assign n56533 = ~pi1147 & ~n56532;
  assign n56534 = ~n65602 & n56533;
  assign n56535 = ~n56525 & ~n56534;
  assign n56536 = ~pi1150 & ~n56535;
  assign n56537 = n55352 & n55609;
  assign n56538 = pi1147 & ~n56537;
  assign n56539 = ~n55100 & ~n55165;
  assign n56540 = ~pi1151 & n56539;
  assign n56541 = n56538 & ~n56540;
  assign n56542 = n55156 & ~n56262;
  assign n56543 = n65536 & ~n56542;
  assign n56544 = n56531 & ~n56543;
  assign n56545 = ~n54867 & n56526;
  assign n56546 = ~pi1147 & ~n56545;
  assign n56547 = ~n56544 & n56546;
  assign n56548 = ~n56541 & ~n56547;
  assign n56549 = pi1150 & ~n56548;
  assign n56550 = ~pi1148 & ~n56549;
  assign n56551 = ~n56536 & n56550;
  assign n56552 = pi212 & ~n54436;
  assign n56553 = n56148 & ~n56552;
  assign n56554 = n55132 & ~n56553;
  assign n56555 = n55330 & ~n56554;
  assign n56556 = pi1147 & ~n56555;
  assign n56557 = n65324 & ~n65499;
  assign n56558 = n62455 & ~n56557;
  assign n56559 = ~n54885 & ~n56557;
  assign n56560 = n65533 & n56559;
  assign n56561 = ~n54885 & n65533;
  assign n56562 = ~n56557 & n56561;
  assign n56563 = n54893 & n56558;
  assign n56564 = ~pi1151 & ~n55051;
  assign n56565 = ~n65603 & n56564;
  assign n56566 = ~n55166 & n56565;
  assign n56567 = n56556 & ~n56566;
  assign n56568 = ~n55387 & n56148;
  assign n56569 = n54782 & ~n56568;
  assign n56570 = ~n54485 & ~n56569;
  assign n56571 = pi1151 & n56570;
  assign n56572 = n55384 & ~n56569;
  assign n56573 = ~pi1151 & ~n54485;
  assign n56574 = ~n65603 & n56573;
  assign n56575 = ~pi1147 & ~n56574;
  assign n56576 = ~n65604 & n56575;
  assign n56577 = ~n56567 & ~n56576;
  assign n56578 = ~pi1150 & ~n56577;
  assign n56579 = pi1147 & ~n55652;
  assign n56580 = ~n55051 & ~n55173;
  assign n56581 = n55620 & n56580;
  assign n56582 = n56579 & ~n56581;
  assign n56583 = ~n55151 & n65536;
  assign n56584 = ~n56543 & ~n56583;
  assign n56585 = n56573 & n56584;
  assign n56586 = n55384 & ~n65580;
  assign n56587 = ~pi1147 & ~n56586;
  assign n56588 = ~n56585 & n56587;
  assign n56589 = ~n56582 & ~n56588;
  assign n56590 = pi1150 & ~n56589;
  assign n56591 = pi1148 & ~n56590;
  assign n56592 = ~n56578 & n56591;
  assign n56593 = pi1149 & ~n56592;
  assign n56594 = ~n56551 & n56593;
  assign n56595 = ~pi1147 & ~n55641;
  assign n56596 = pi1151 & ~n55056;
  assign n56597 = ~n55213 & ~n56225;
  assign n56598 = n56596 & ~n56597;
  assign n56599 = n56595 & ~n56598;
  assign n56600 = n55183 & ~n55201;
  assign n56601 = ~n56207 & ~n56600;
  assign n56602 = ~n55068 & ~n56601;
  assign n56603 = ~pi1151 & n56602;
  assign n56604 = n54827 & ~n56231;
  assign n56605 = pi1151 & ~n55068;
  assign n56606 = ~n56604 & n56605;
  assign n56607 = pi1147 & ~n56606;
  assign n56608 = pi1147 & ~n56603;
  assign n56609 = ~n56606 & n56608;
  assign n56610 = ~n56603 & n56607;
  assign n56611 = ~n56599 & ~n65605;
  assign n56612 = pi1150 & ~n56611;
  assign n56613 = n52475 & ~n65362;
  assign n56614 = ~pi1151 & ~n56613;
  assign n56615 = ~pi1147 & ~n56614;
  assign n56616 = n54606 & ~n55314;
  assign n56617 = n56596 & ~n56616;
  assign n56618 = n56615 & ~n56617;
  assign n56619 = ~n55526 & n56605;
  assign n56620 = pi1147 & ~n55653;
  assign n56621 = ~n56619 & n56620;
  assign n56622 = ~n56618 & ~n56621;
  assign n56623 = ~pi1150 & ~n56622;
  assign n56624 = pi1148 & ~n56623;
  assign n56625 = ~n56612 & n56624;
  assign n56626 = ~n65577 & n56604;
  assign n56627 = n54495 & ~n56626;
  assign n56628 = ~n54494 & ~n56214;
  assign n56629 = ~pi1151 & n56628;
  assign n56630 = pi1147 & ~n56629;
  assign n56631 = ~n56627 & n56630;
  assign n56632 = ~pi1151 & ~n54907;
  assign n56633 = ~pi1147 & ~n56632;
  assign n56634 = pi1151 & ~n55212;
  assign n56635 = n56633 & ~n56634;
  assign n56636 = pi1150 & ~n56635;
  assign n56637 = ~n56631 & n56636;
  assign n56638 = ~n54388 & n55607;
  assign n56639 = n55524 & ~n56638;
  assign n56640 = n54495 & ~n56639;
  assign n56641 = n55361 & ~n55608;
  assign n56642 = pi1147 & ~n56641;
  assign n56643 = ~n56640 & n56642;
  assign n56644 = ~pi1147 & pi1151;
  assign n56645 = n65476 & n56644;
  assign n56646 = ~pi1150 & ~n56645;
  assign n56647 = ~n56643 & n56646;
  assign n56648 = ~n56637 & ~n56647;
  assign n56649 = ~pi1148 & ~n56648;
  assign n56650 = ~pi1149 & ~n56649;
  assign n56651 = ~n56625 & n56650;
  assign n56652 = ~pi1150 & ~n56534;
  assign n56653 = ~n56525 & n56652;
  assign n56654 = pi1150 & ~n56547;
  assign n56655 = pi1150 & ~n56541;
  assign n56656 = ~n56547 & n56655;
  assign n56657 = ~n56541 & n56654;
  assign n56658 = ~n56653 & ~n65606;
  assign n56659 = pi1149 & ~n56549;
  assign n56660 = ~n56536 & n56659;
  assign n56661 = pi1149 & ~n56658;
  assign n56662 = ~pi1149 & ~n56648;
  assign n56663 = ~n65607 & ~n56662;
  assign n56664 = ~pi1148 & ~n56663;
  assign n56665 = ~pi1149 & ~n65605;
  assign n56666 = ~n56599 & n56665;
  assign n56667 = pi1149 & ~n56582;
  assign n56668 = ~n56588 & n56667;
  assign n56669 = pi1150 & ~n56668;
  assign n56670 = ~n56666 & n56669;
  assign n56671 = pi1149 & ~n56576;
  assign n56672 = ~n56567 & n56671;
  assign n56673 = ~pi1149 & ~n56621;
  assign n56674 = ~pi1149 & ~n56618;
  assign n56675 = ~n56621 & n56674;
  assign n56676 = ~n56618 & n56673;
  assign n56677 = ~pi1150 & ~n65608;
  assign n56678 = ~n56672 & n56677;
  assign n56679 = pi1148 & ~n56678;
  assign n56680 = ~n56670 & n56679;
  assign n56681 = ~n56664 & ~n56680;
  assign n56682 = ~n56670 & ~n56678;
  assign n56683 = pi1148 & ~n56682;
  assign n56684 = ~pi1148 & ~n56662;
  assign n56685 = ~n65607 & n56684;
  assign n56686 = ~n56683 & ~n56685;
  assign n56687 = ~n56594 & ~n56651;
  assign n56688 = ~pi213 & n65609;
  assign n56689 = pi213 & n55662;
  assign n56690 = pi209 & ~n56689;
  assign n56691 = ~n56688 & n56690;
  assign n56692 = n55198 & n55205;
  assign n56693 = n55384 & ~n56692;
  assign n56694 = n56595 & ~n56693;
  assign n56695 = n55384 & n56584;
  assign n56696 = n55408 & ~n56583;
  assign n56697 = pi1147 & ~n56696;
  assign n56698 = ~n56695 & n56697;
  assign n56699 = pi1150 & ~n56698;
  assign n56700 = ~n56694 & n56699;
  assign n56701 = n56526 & ~n56543;
  assign n56702 = pi1147 & ~n55620;
  assign n56703 = ~n56701 & n56702;
  assign n56704 = n62455 & ~n55507;
  assign n56705 = ~n65526 & n56704;
  assign n56706 = ~n55438 & ~n56705;
  assign n56707 = n56633 & n56706;
  assign n56708 = ~pi1150 & ~n56707;
  assign n56709 = ~n56703 & n56708;
  assign n56710 = ~pi1149 & ~n56709;
  assign n56711 = ~n56700 & n56710;
  assign n56712 = n55361 & ~n56626;
  assign n56713 = ~n55100 & ~n56239;
  assign n56714 = pi1151 & n56713;
  assign n56715 = ~pi1147 & ~n56714;
  assign n56716 = ~n56712 & n56715;
  assign n56717 = ~n65505 & n56641;
  assign n56718 = n56538 & ~n56717;
  assign n56719 = ~pi1150 & ~n56718;
  assign n56720 = ~n56716 & n56719;
  assign n56721 = n55292 & ~n56604;
  assign n56722 = ~n54831 & n55216;
  assign n56723 = n54827 & ~n56722;
  assign n56724 = n55330 & ~n56723;
  assign n56725 = ~pi1147 & ~n56724;
  assign n56726 = ~n56721 & n56725;
  assign n56727 = ~n55068 & ~n55612;
  assign n56728 = ~pi1151 & n56727;
  assign n56729 = n56579 & ~n56728;
  assign n56730 = pi1150 & ~n56729;
  assign n56731 = ~n56726 & n56730;
  assign n56732 = pi1149 & ~n56731;
  assign n56733 = ~n56720 & n56732;
  assign n56734 = pi1148 & ~n56733;
  assign n56735 = ~n56711 & n56734;
  assign n56736 = ~pi219 & ~n55312;
  assign n56737 = ~n55312 & n55551;
  assign n56738 = ~n55550 & n56736;
  assign n56739 = n55132 & ~n65610;
  assign n56740 = ~n55128 & n56739;
  assign n56741 = n55361 & ~n56740;
  assign n56742 = n56522 & ~n56741;
  assign n56743 = n54402 & n54606;
  assign n56744 = ~n39342 & n56743;
  assign n56745 = ~n56639 & ~n56744;
  assign n56746 = n55352 & n56745;
  assign n56747 = ~pi1151 & ~n56639;
  assign n56748 = ~n54494 & n56747;
  assign n56749 = n55361 & ~n56639;
  assign n56750 = ~pi1147 & ~n65611;
  assign n56751 = ~pi1147 & ~n56746;
  assign n56752 = ~n65611 & n56751;
  assign n56753 = ~n56746 & n56750;
  assign n56754 = ~pi1150 & ~n65612;
  assign n56755 = ~n56742 & n56754;
  assign n56756 = ~n55068 & ~n56739;
  assign n56757 = ~pi1151 & n56756;
  assign n56758 = n56556 & ~n56757;
  assign n56759 = n55292 & ~n55526;
  assign n56760 = n55330 & ~n56743;
  assign n56761 = ~n55526 & n56760;
  assign n56762 = ~pi1147 & ~n56761;
  assign n56763 = ~pi1147 & ~n56759;
  assign n56764 = ~n56761 & n56763;
  assign n56765 = ~n56759 & n56762;
  assign n56766 = pi1150 & ~n65613;
  assign n56767 = ~n56758 & n56766;
  assign n56768 = pi1149 & ~n56767;
  assign n56769 = ~n56755 & n56768;
  assign n56770 = n55153 & n65533;
  assign n56771 = ~n55056 & ~n56770;
  assign n56772 = ~pi1151 & n56771;
  assign n56773 = n55408 & ~n56770;
  assign n56774 = n55384 & ~n65603;
  assign n56775 = pi1147 & ~n56774;
  assign n56776 = ~n65614 & n56775;
  assign n56777 = ~n65014 & n65430;
  assign n56778 = pi1151 & ~n56777;
  assign n56779 = n56615 & ~n56778;
  assign n56780 = pi1150 & ~n56779;
  assign n56781 = ~n56776 & n56780;
  assign n56782 = ~n65464 & ~n55580;
  assign n56783 = ~pi1151 & ~n56163;
  assign n56784 = pi1147 & ~n56783;
  assign n56785 = ~n56782 & n56784;
  assign n56786 = n55136 & n56644;
  assign n56787 = ~pi1150 & ~n56786;
  assign n56788 = ~n56785 & n56787;
  assign n56789 = ~pi1149 & ~n56788;
  assign n56790 = ~n56781 & n56789;
  assign n56791 = ~pi1148 & ~n56790;
  assign n56792 = ~n56769 & n56791;
  assign n56793 = pi213 & ~n56792;
  assign n56794 = ~n56700 & ~n56709;
  assign n56795 = ~pi1149 & ~n56794;
  assign n56796 = ~n56720 & ~n56731;
  assign n56797 = pi1149 & ~n56796;
  assign n56798 = pi1148 & ~n56797;
  assign n56799 = ~n56711 & ~n56733;
  assign n56800 = pi1148 & ~n56799;
  assign n56801 = ~n56795 & n56798;
  assign n56802 = ~n56755 & ~n56767;
  assign n56803 = pi1149 & ~n56802;
  assign n56804 = ~n56781 & ~n56788;
  assign n56805 = ~pi1149 & ~n56804;
  assign n56806 = ~pi1148 & ~n56805;
  assign n56807 = ~n56803 & n56806;
  assign n56808 = ~n65615 & ~n56807;
  assign n56809 = pi213 & ~n56808;
  assign n56810 = ~n56735 & n56793;
  assign n56811 = ~pi213 & ~n55243;
  assign n56812 = ~pi209 & ~n56811;
  assign n56813 = ~n65616 & n56812;
  assign n56814 = ~pi213 & ~n65609;
  assign n56815 = pi213 & ~n55662;
  assign n56816 = pi209 & ~n56815;
  assign n56817 = ~n56814 & n56816;
  assign n56818 = pi213 & ~n65615;
  assign n56819 = ~n56807 & n56818;
  assign n56820 = ~pi213 & n55243;
  assign n56821 = ~pi209 & ~n56820;
  assign n56822 = ~n56819 & n56821;
  assign n56823 = ~n56817 & ~n56822;
  assign n56824 = ~n56691 & ~n56813;
  assign n56825 = pi230 & n65617;
  assign n56826 = ~pi230 & ~pi247;
  assign n56827 = pi230 & ~n65617;
  assign n56828 = ~pi230 & pi247;
  assign n56829 = ~n56827 & ~n56828;
  assign n56830 = ~n56825 & ~n56826;
  assign n56831 = ~pi1151 & n55134;
  assign n56832 = ~n55133 & n56523;
  assign n56833 = pi1152 & ~n65619;
  assign n56834 = ~n56537 & n56833;
  assign n56835 = pi1151 & n56539;
  assign n56836 = ~pi1152 & ~n56524;
  assign n56837 = ~n56835 & n56836;
  assign n56838 = ~n56834 & ~n56837;
  assign n56839 = pi1150 & ~n56838;
  assign n56840 = pi1152 & ~n65611;
  assign n56841 = ~n56627 & n56840;
  assign n56842 = pi1151 & n56628;
  assign n56843 = ~pi1152 & ~n56641;
  assign n56844 = ~n56842 & n56843;
  assign n56845 = ~n56841 & ~n56844;
  assign n56846 = ~n56627 & ~n65611;
  assign n56847 = pi1152 & ~n56846;
  assign n56848 = ~n56641 & ~n56842;
  assign n56849 = ~pi1152 & ~n56848;
  assign n56850 = ~pi1150 & ~n56849;
  assign n56851 = ~n56847 & n56850;
  assign n56852 = ~pi1150 & ~n56845;
  assign n56853 = pi1148 & ~n65620;
  assign n56854 = ~n56839 & n56853;
  assign n56855 = pi1151 & ~pi1152;
  assign n56856 = n54907 & n56855;
  assign n56857 = ~pi1151 & ~n65476;
  assign n56858 = pi1152 & ~n56857;
  assign n56859 = pi1152 & ~n56634;
  assign n56860 = ~n56857 & n56859;
  assign n56861 = ~n56634 & n56858;
  assign n56862 = ~pi1150 & ~n65621;
  assign n56863 = ~pi1150 & ~n56856;
  assign n56864 = ~n65621 & n56863;
  assign n56865 = ~n56856 & n56862;
  assign n56866 = ~pi1151 & n56528;
  assign n56867 = ~n56527 & n56531;
  assign n56868 = pi1152 & ~n56545;
  assign n56869 = ~n65623 & n56868;
  assign n56870 = ~pi1152 & ~n56532;
  assign n56871 = ~n56701 & n56870;
  assign n56872 = pi1150 & ~n56871;
  assign n56873 = ~n56869 & n56872;
  assign n56874 = ~n65622 & ~n56873;
  assign n56875 = ~pi1148 & ~n56874;
  assign n56876 = ~pi1149 & ~n56875;
  assign n56877 = ~n56854 & n56876;
  assign n56878 = ~n55206 & n56596;
  assign n56879 = ~pi1152 & ~n56878;
  assign n56880 = ~n56614 & n56879;
  assign n56881 = n55408 & ~n56616;
  assign n56882 = pi1152 & ~n56881;
  assign n56883 = ~n56598 & n56882;
  assign n56884 = ~pi1150 & ~n56883;
  assign n56885 = ~n56880 & n56884;
  assign n56886 = ~pi1152 & ~n56574;
  assign n56887 = ~n56695 & n56886;
  assign n56888 = ~pi1151 & n56570;
  assign n56889 = ~n56569 & n56573;
  assign n56890 = pi1152 & ~n56586;
  assign n56891 = ~n65624 & n56890;
  assign n56892 = pi1150 & ~n56891;
  assign n56893 = pi1150 & ~n56887;
  assign n56894 = ~n56891 & n56893;
  assign n56895 = ~n56887 & n56892;
  assign n56896 = ~n56885 & ~n65625;
  assign n56897 = ~pi1148 & ~n56896;
  assign n56898 = pi1151 & n56602;
  assign n56899 = ~pi1152 & ~n55653;
  assign n56900 = ~n56898 & n56899;
  assign n56901 = pi1152 & ~n56759;
  assign n56902 = ~n56606 & n56901;
  assign n56903 = ~pi1150 & ~n56902;
  assign n56904 = ~pi1150 & ~n56900;
  assign n56905 = ~n56902 & n56904;
  assign n56906 = ~n56900 & n56903;
  assign n56907 = pi1152 & ~n55652;
  assign n56908 = ~n56554 & n56564;
  assign n56909 = n56907 & ~n56908;
  assign n56910 = pi1151 & ~n54909;
  assign n56911 = n56580 & n56910;
  assign n56912 = ~pi1152 & ~n56911;
  assign n56913 = ~n56566 & n56912;
  assign n56914 = pi1150 & ~n56913;
  assign n56915 = ~n56909 & n56914;
  assign n56916 = ~n65626 & ~n56915;
  assign n56917 = pi1148 & ~n56916;
  assign n56918 = pi1149 & ~n56917;
  assign n56919 = pi1148 & ~n56915;
  assign n56920 = pi1148 & ~n65626;
  assign n56921 = ~n56915 & n56920;
  assign n56922 = ~n65626 & n56919;
  assign n56923 = ~pi1148 & ~n65625;
  assign n56924 = ~n56885 & n56923;
  assign n56925 = ~n65627 & ~n56924;
  assign n56926 = pi1149 & ~n56925;
  assign n56927 = ~n56897 & n56918;
  assign n56928 = ~n56839 & ~n65620;
  assign n56929 = pi1148 & ~n56928;
  assign n56930 = ~pi1148 & ~n65622;
  assign n56931 = ~n56873 & n56930;
  assign n56932 = ~pi1149 & ~n56931;
  assign n56933 = ~n56929 & n56932;
  assign n56934 = pi1149 & ~n65627;
  assign n56935 = ~n56924 & n56934;
  assign n56936 = ~n56933 & ~n56935;
  assign n56937 = ~n56877 & ~n65628;
  assign n56938 = ~pi213 & n65629;
  assign n56939 = ~n55207 & n56855;
  assign n56940 = ~pi1151 & ~n55136;
  assign n56941 = ~n65476 & n56940;
  assign n56942 = pi1152 & ~n56941;
  assign n56943 = ~n55642 & n56942;
  assign n56944 = ~pi1150 & ~n56943;
  assign n56945 = ~n56939 & n56944;
  assign n56946 = ~n55652 & n56833;
  assign n56947 = ~n65619 & n56907;
  assign n56948 = pi1151 & n65500;
  assign n56949 = ~pi1152 & ~n56948;
  assign n56950 = ~n55649 & n56949;
  assign n56951 = pi1150 & ~n56950;
  assign n56952 = ~n65630 & n56951;
  assign n56953 = ~n56939 & ~n56943;
  assign n56954 = ~pi1150 & ~n56953;
  assign n56955 = ~n65630 & ~n56950;
  assign n56956 = pi1150 & ~n56955;
  assign n56957 = ~n56954 & ~n56956;
  assign n56958 = ~n56945 & ~n56952;
  assign n56959 = pi213 & ~n65631;
  assign n56960 = pi209 & ~n56959;
  assign n56961 = ~n56938 & n56960;
  assign n56962 = ~n56555 & n56833;
  assign n56963 = pi1151 & n56756;
  assign n56964 = ~pi1152 & ~n56741;
  assign n56965 = ~n56963 & n56964;
  assign n56966 = pi1150 & ~n56965;
  assign n56967 = pi1150 & ~n56962;
  assign n56968 = ~n56965 & n56967;
  assign n56969 = ~n56962 & n56966;
  assign n56970 = pi1151 & n56771;
  assign n56971 = n56596 & ~n56770;
  assign n56972 = ~pi1152 & ~n56783;
  assign n56973 = ~n65633 & n56972;
  assign n56974 = pi1152 & ~n56532;
  assign n56975 = ~n56774 & n56974;
  assign n56976 = ~pi1150 & ~n56975;
  assign n56977 = ~n56973 & n56976;
  assign n56978 = ~pi1149 & ~n56977;
  assign n56979 = ~n65632 & n56978;
  assign n56980 = pi1152 & ~n56544;
  assign n56981 = ~n56695 & n56980;
  assign n56982 = ~n56583 & n56596;
  assign n56983 = n55621 & ~n56982;
  assign n56984 = ~pi1150 & ~n56983;
  assign n56985 = ~n56981 & n56984;
  assign n56986 = n55609 & n56523;
  assign n56987 = n56907 & ~n56986;
  assign n56988 = pi1151 & n56727;
  assign n56989 = ~pi1152 & ~n56717;
  assign n56990 = ~n56988 & n56989;
  assign n56991 = pi1150 & ~n56990;
  assign n56992 = pi1150 & ~n56987;
  assign n56993 = ~n56990 & n56992;
  assign n56994 = ~n56987 & n56991;
  assign n56995 = pi1149 & ~n65634;
  assign n56996 = ~n56985 & n56995;
  assign n56997 = pi1148 & ~n56996;
  assign n56998 = ~n56979 & n56997;
  assign n56999 = ~n56632 & n56879;
  assign n57000 = ~pi1151 & ~n56706;
  assign n57001 = pi1152 & ~n57000;
  assign n57002 = ~n56693 & n57001;
  assign n57003 = ~pi1150 & ~n57002;
  assign n57004 = ~n56999 & n57003;
  assign n57005 = ~pi1152 & ~n56606;
  assign n57006 = ~n56712 & n57005;
  assign n57007 = ~pi1151 & n56713;
  assign n57008 = pi1152 & ~n56724;
  assign n57009 = ~n57007 & n57008;
  assign n57010 = pi1150 & ~n57009;
  assign n57011 = ~n57006 & n57010;
  assign n57012 = pi1149 & ~n57011;
  assign n57013 = ~n57004 & n57012;
  assign n57014 = n56523 & n56745;
  assign n57015 = pi1152 & ~n56761;
  assign n57016 = ~n57014 & n57015;
  assign n57017 = ~pi1152 & ~n65611;
  assign n57018 = ~pi1152 & ~n56619;
  assign n57019 = ~n65611 & n57018;
  assign n57020 = ~n56619 & n57017;
  assign n57021 = pi1150 & ~n65635;
  assign n57022 = ~n57016 & n57021;
  assign n57023 = pi1152 & ~n56778;
  assign n57024 = ~n56940 & n57023;
  assign n57025 = n56613 & n56855;
  assign n57026 = ~pi1150 & ~n57025;
  assign n57027 = ~n57024 & n57026;
  assign n57028 = ~pi1149 & ~n57027;
  assign n57029 = ~n57022 & n57028;
  assign n57030 = ~pi1148 & ~n57029;
  assign n57031 = ~n57013 & n57030;
  assign n57032 = pi213 & ~n57031;
  assign n57033 = pi213 & ~n56998;
  assign n57034 = ~n57031 & n57033;
  assign n57035 = ~n56998 & n57032;
  assign n57036 = ~pi213 & ~n56479;
  assign n57037 = ~pi209 & ~n57036;
  assign n57038 = ~n65636 & n57037;
  assign n57039 = ~pi213 & ~n65629;
  assign n57040 = pi213 & n65631;
  assign n57041 = pi209 & ~n57040;
  assign n57042 = ~n57039 & n57041;
  assign n57043 = ~n56962 & ~n56965;
  assign n57044 = pi1150 & ~n57043;
  assign n57045 = ~n56973 & ~n56975;
  assign n57046 = ~pi1150 & ~n57045;
  assign n57047 = ~pi1149 & ~n57046;
  assign n57048 = ~n57044 & n57047;
  assign n57049 = ~n56985 & ~n65634;
  assign n57050 = pi1149 & ~n57049;
  assign n57051 = pi1148 & ~n57050;
  assign n57052 = ~n57048 & n57051;
  assign n57053 = ~n57013 & ~n57029;
  assign n57054 = ~pi1148 & ~n57053;
  assign n57055 = pi213 & ~n57054;
  assign n57056 = ~n57052 & n57055;
  assign n57057 = ~pi213 & n56479;
  assign n57058 = ~pi209 & ~n57057;
  assign n57059 = ~n57056 & n57058;
  assign n57060 = ~n57042 & ~n57059;
  assign n57061 = ~n56961 & ~n57038;
  assign n57062 = pi230 & n65637;
  assign n57063 = ~pi230 & ~pi248;
  assign n57064 = pi230 & ~n65637;
  assign n57065 = ~pi230 & pi248;
  assign n57066 = ~n57064 & ~n57065;
  assign n57067 = ~n57062 & ~n57063;
  assign n57068 = pi209 & n53976;
  assign n57069 = pi57 & ~n53833;
  assign n57070 = pi299 & n53797;
  assign n57071 = ~n55592 & ~n57070;
  assign n57072 = ~pi214 & ~n57071;
  assign n57073 = ~n54362 & n54627;
  assign n57074 = pi212 & ~n57073;
  assign n57075 = ~n57072 & n57074;
  assign n57076 = pi214 & ~n57071;
  assign n57077 = ~pi212 & ~n54391;
  assign n57078 = ~n57076 & n57077;
  assign n57079 = ~pi219 & ~n57078;
  assign n57080 = ~pi219 & ~n57075;
  assign n57081 = ~n57078 & n57080;
  assign n57082 = ~n57075 & n57079;
  assign n57083 = n55589 & ~n65639;
  assign n57084 = ~n3475 & n53833;
  assign n57085 = ~pi57 & pi1151;
  assign n57086 = ~n57084 & n57085;
  assign n57087 = ~n57083 & n57086;
  assign n57088 = pi1151 & ~n57083;
  assign n57089 = ~pi57 & ~n57088;
  assign n57090 = ~n53834 & ~n57089;
  assign n57091 = ~n57069 & ~n57087;
  assign n57092 = ~n54885 & ~n57070;
  assign n57093 = ~n54391 & n57092;
  assign n57094 = ~pi212 & ~n57093;
  assign n57095 = ~pi214 & n57092;
  assign n57096 = ~n48498 & ~n54884;
  assign n57097 = n53818 & ~n57096;
  assign n57098 = pi212 & ~n57097;
  assign n57099 = ~n57095 & n57098;
  assign n57100 = ~n57094 & ~n57099;
  assign n57101 = ~pi219 & ~n57100;
  assign n57102 = n55563 & ~n57101;
  assign n57103 = n50734 & ~n57084;
  assign n57104 = ~n57102 & n57103;
  assign n57105 = ~n65640 & ~n57104;
  assign n57106 = ~pi1152 & ~n57105;
  assign n57107 = ~pi214 & ~n57070;
  assign n57108 = ~n53818 & ~n57107;
  assign n57109 = n55118 & ~n65534;
  assign n57110 = ~n54436 & ~n57070;
  assign n57111 = ~pi214 & ~n57110;
  assign n57112 = pi212 & ~n57111;
  assign n57113 = ~n57109 & n57112;
  assign n57114 = n56552 & ~n57108;
  assign n57115 = n55306 & ~n57070;
  assign n57116 = n56147 & ~n57115;
  assign n57117 = ~n65641 & n57116;
  assign n57118 = ~pi1151 & ~n57117;
  assign n57119 = n55132 & n57118;
  assign n57120 = pi299 & ~n53797;
  assign n57121 = ~n39342 & n57120;
  assign n57122 = ~n53796 & ~n57121;
  assign n57123 = n52569 & ~n57122;
  assign n57124 = n55602 & ~n57123;
  assign n57125 = ~n54847 & ~n55163;
  assign n57126 = pi1151 & ~n57125;
  assign n57127 = ~n57124 & n57126;
  assign n57128 = n53802 & ~n57127;
  assign n57129 = ~n57119 & n57128;
  assign n57130 = ~n57106 & ~n57129;
  assign n57131 = pi1150 & ~n57130;
  assign n57132 = n54834 & ~n57120;
  assign n57133 = pi212 & ~n57132;
  assign n57134 = ~n55482 & n57133;
  assign n57135 = ~pi212 & n65450;
  assign n57136 = ~pi219 & ~n57135;
  assign n57137 = ~n57115 & n57136;
  assign n57138 = ~n57134 & n57137;
  assign n57139 = n54827 & ~n57138;
  assign n57140 = pi1151 & ~n57139;
  assign n57141 = ~n56747 & ~n57140;
  assign n57142 = n53802 & ~n57141;
  assign n57143 = ~n55184 & ~n57070;
  assign n57144 = pi211 & n55508;
  assign n57145 = ~n52768 & n55191;
  assign n57146 = ~n65324 & ~n57145;
  assign n57147 = ~n57144 & n57146;
  assign n57148 = ~n65324 & ~n57144;
  assign n57149 = ~n57145 & n57148;
  assign n57150 = ~n65324 & ~n57143;
  assign n57151 = n39342 & n55509;
  assign n57152 = ~n65642 & ~n57151;
  assign n57153 = ~pi219 & ~n57152;
  assign n57154 = ~n65430 & ~n54906;
  assign n57155 = n50537 & ~n57154;
  assign n57156 = n53970 & ~n54906;
  assign n57157 = ~n65642 & ~n57156;
  assign n57158 = ~n57151 & ~n57156;
  assign n57159 = ~n65642 & n57158;
  assign n57160 = ~n57151 & n57157;
  assign n57161 = ~pi219 & ~n65643;
  assign n57162 = pi1151 & n55205;
  assign n57163 = ~n57161 & n57162;
  assign n57164 = ~n57153 & n57155;
  assign n57165 = n53835 & ~n65644;
  assign n57166 = ~n57142 & ~n57165;
  assign n57167 = ~n54362 & ~n57121;
  assign n57168 = n65182 & n53832;
  assign n57169 = ~n57167 & n57168;
  assign n57170 = ~pi1150 & ~n57169;
  assign n57171 = ~n57166 & n57170;
  assign n57172 = ~pi209 & ~n57171;
  assign n57173 = ~n57131 & n57172;
  assign n57174 = pi213 & ~n57173;
  assign n57175 = ~n57068 & n57174;
  assign n57176 = pi214 & ~n65426;
  assign n57177 = ~n53880 & ~n57176;
  assign n57178 = ~pi212 & ~n57177;
  assign n57179 = ~pi214 & n65426;
  assign n57180 = ~pi211 & n53869;
  assign n57181 = ~n53912 & ~n57180;
  assign n57182 = pi214 & ~n57181;
  assign n57183 = pi212 & ~n57182;
  assign n57184 = pi212 & ~n57179;
  assign n57185 = ~n57182 & n57184;
  assign n57186 = ~n57179 & n57183;
  assign n57187 = ~n57178 & ~n65645;
  assign n57188 = ~pi219 & ~n57187;
  assign n57189 = n53879 & ~n57188;
  assign n57190 = n56523 & ~n57189;
  assign n57191 = pi214 & n53861;
  assign n57192 = n53881 & ~n57191;
  assign n57193 = ~pi219 & ~n57192;
  assign n57194 = pi212 & ~n53861;
  assign n57195 = n57193 & ~n57194;
  assign n57196 = n53879 & ~n57195;
  assign n57197 = n55330 & ~n57196;
  assign n57198 = pi1152 & ~n57197;
  assign n57199 = ~n57190 & n57198;
  assign n57200 = n52766 & ~n54143;
  assign n57201 = ~pi207 & n54142;
  assign n57202 = pi207 & ~n52786;
  assign n57203 = ~n50091 & n57202;
  assign n57204 = pi208 & ~n57203;
  assign n57205 = ~n57201 & n57204;
  assign n57206 = ~n57200 & ~n57205;
  assign n57207 = ~pi211 & n57206;
  assign n57208 = ~n54044 & ~n57207;
  assign n57209 = ~n52517 & n57208;
  assign n57210 = pi219 & ~n54043;
  assign n57211 = ~n57209 & n57210;
  assign n57212 = n62455 & ~n57211;
  assign n57213 = ~n39343 & ~n53964;
  assign n57214 = pi211 & ~n57206;
  assign n57215 = pi214 & n57214;
  assign n57216 = ~n57213 & ~n57215;
  assign n57217 = ~pi212 & ~n57216;
  assign n57218 = ~pi219 & ~n57217;
  assign n57219 = ~pi211 & ~n53964;
  assign n57220 = ~pi214 & ~n57219;
  assign n57221 = ~n57214 & n57220;
  assign n57222 = pi212 & ~n57221;
  assign n57223 = pi214 & n57206;
  assign n57224 = n57222 & ~n57223;
  assign n57225 = n57218 & ~n57224;
  assign n57226 = n57212 & ~n57225;
  assign n57227 = n56605 & ~n57226;
  assign n57228 = pi212 & ~n57216;
  assign n57229 = ~pi212 & ~n53964;
  assign n57230 = ~pi219 & ~n57229;
  assign n57231 = ~n57228 & n57230;
  assign n57232 = n57212 & ~n57231;
  assign n57233 = n55361 & ~n57232;
  assign n57234 = ~pi1152 & ~n57233;
  assign n57235 = ~n57227 & n57234;
  assign n57236 = pi1150 & ~n57235;
  assign n57237 = ~n57199 & n57236;
  assign n57238 = ~n53964 & n54010;
  assign n57239 = ~n56855 & ~n57238;
  assign n57240 = pi214 & ~n57208;
  assign n57241 = n57222 & ~n57240;
  assign n57242 = n57218 & ~n57241;
  assign n57243 = n53969 & ~n57242;
  assign n57244 = n56596 & ~n57243;
  assign n57245 = ~n57239 & ~n57244;
  assign n57246 = ~pi214 & n53861;
  assign n57247 = pi212 & ~n57246;
  assign n57248 = ~n57176 & n57247;
  assign n57249 = n57193 & ~n57248;
  assign n57250 = n62455 & ~n53876;
  assign n57251 = ~n57249 & n57250;
  assign n57252 = n55384 & ~n57251;
  assign n57253 = ~n65426 & n54554;
  assign n57254 = ~n53869 & ~n54554;
  assign n57255 = n62455 & ~n57254;
  assign n57256 = ~n57253 & n57255;
  assign n57257 = n56531 & ~n57256;
  assign n57258 = pi1152 & ~n57257;
  assign n57259 = ~n57252 & n57258;
  assign n57260 = ~pi1150 & ~n57259;
  assign n57261 = ~n57245 & n57260;
  assign n57262 = ~n57245 & ~n57259;
  assign n57263 = ~pi1150 & ~n57262;
  assign n57264 = ~n57199 & ~n57235;
  assign n57265 = pi1150 & ~n57264;
  assign n57266 = ~n57263 & ~n57265;
  assign n57267 = ~n57237 & ~n57261;
  assign n57268 = pi209 & ~n65646;
  assign n57269 = ~pi209 & ~n65631;
  assign n57270 = ~pi213 & ~n57269;
  assign n57271 = ~n57268 & n57270;
  assign n57272 = pi209 & ~n53976;
  assign n57273 = pi1150 & ~n57129;
  assign n57274 = ~n57106 & n57273;
  assign n57275 = n53835 & ~n57169;
  assign n57276 = ~n65644 & n57275;
  assign n57277 = pi1151 & n54827;
  assign n57278 = n50537 & ~n54826;
  assign n57279 = ~n57138 & n65647;
  assign n57280 = ~pi1151 & n56639;
  assign n57281 = n53802 & ~n57169;
  assign n57282 = ~n57280 & n57281;
  assign n57283 = ~n57279 & n57282;
  assign n57284 = ~pi1150 & ~n57283;
  assign n57285 = ~n57276 & n57284;
  assign n57286 = ~pi209 & ~n57285;
  assign n57287 = ~n57274 & n57286;
  assign n57288 = pi213 & ~n57287;
  assign n57289 = ~n57272 & n57288;
  assign n57290 = pi209 & n65646;
  assign n57291 = ~pi209 & n65631;
  assign n57292 = ~pi213 & ~n57291;
  assign n57293 = ~n57290 & n57292;
  assign n57294 = ~n57289 & ~n57293;
  assign n57295 = ~pi213 & ~n65631;
  assign n57296 = ~n57274 & ~n57285;
  assign n57297 = pi213 & ~n57296;
  assign n57298 = ~pi209 & ~n57297;
  assign n57299 = ~n57295 & n57298;
  assign n57300 = ~pi213 & ~n57261;
  assign n57301 = ~pi213 & ~n65646;
  assign n57302 = ~n57237 & n57300;
  assign n57303 = pi213 & n53976;
  assign n57304 = pi209 & ~n57303;
  assign n57305 = ~n65649 & n57304;
  assign n57306 = ~n57299 & ~n57305;
  assign n57307 = ~n57175 & ~n57271;
  assign n57308 = pi230 & n65648;
  assign n57309 = ~pi230 & ~pi249;
  assign n57310 = pi230 & ~n65648;
  assign n57311 = ~pi230 & pi249;
  assign n57312 = ~n57310 & ~n57311;
  assign n57313 = ~n57308 & ~n57309;
  assign n57314 = ~pi273 & ~n49282;
  assign n57315 = ~n49242 & ~n57314;
  assign n57316 = pi219 & ~n57315;
  assign n57317 = ~pi273 & ~n49251;
  assign n57318 = n49253 & ~n57317;
  assign n57319 = pi1091 & pi1146;
  assign n57320 = ~pi211 & n57319;
  assign n57321 = ~pi219 & ~n57320;
  assign n57322 = ~n57318 & n57321;
  assign n57323 = ~n57316 & ~n57322;
  assign n57324 = pi299 & n57323;
  assign n57325 = ~pi200 & n57319;
  assign n57326 = ~pi199 & ~n57325;
  assign n57327 = ~n57318 & n57326;
  assign n57328 = pi199 & ~n57315;
  assign n57329 = ~pi299 & ~n57328;
  assign n57330 = ~n57327 & n57329;
  assign n57331 = ~n57324 & ~n57330;
  assign n57332 = ~n48477 & ~n49421;
  assign n57333 = pi1091 & ~n57332;
  assign n57334 = n57331 & ~n57333;
  assign n57335 = n62455 & ~n57334;
  assign n57336 = pi1091 & n50655;
  assign n57337 = ~n57335 & ~n57336;
  assign n57338 = pi1147 & ~n57337;
  assign n57339 = ~n62455 & n57323;
  assign n57340 = n65497 & ~n57331;
  assign n57341 = ~pi1148 & ~n57340;
  assign n57342 = pi1091 & n39423;
  assign n57343 = ~n57323 & ~n57342;
  assign n57344 = pi299 & ~n57343;
  assign n57345 = ~pi271 & ~n49281;
  assign n57346 = ~n49240 & ~n57345;
  assign n57347 = pi199 & ~n57346;
  assign n57348 = ~pi1091 & ~n49249;
  assign n57349 = pi271 & ~n57348;
  assign n57350 = ~pi271 & ~n49250;
  assign n57351 = ~n57349 & ~n57350;
  assign n57352 = ~n57319 & ~n57351;
  assign n57353 = ~pi199 & n57352;
  assign n57354 = ~n57347 & ~n57353;
  assign n57355 = pi200 & ~n57354;
  assign n57356 = n49472 & ~n57355;
  assign n57357 = ~n57330 & ~n57356;
  assign n57358 = ~n57344 & n57357;
  assign n57359 = n62455 & ~n57358;
  assign n57360 = n48935 & n50334;
  assign n57361 = pi1148 & ~n57360;
  assign n57362 = ~n57359 & n57361;
  assign n57363 = ~n57341 & ~n57362;
  assign n57364 = ~n57339 & ~n57363;
  assign n57365 = ~n57338 & n57364;
  assign n57366 = ~pi230 & ~n57365;
  assign n57367 = ~pi1146 & n39421;
  assign n57368 = pi1147 & n52475;
  assign n57369 = ~n52478 & ~n57368;
  assign n57370 = ~n57367 & ~n57369;
  assign n57371 = ~pi1146 & n39538;
  assign n57372 = ~pi199 & pi1147;
  assign n57373 = pi200 & ~n57372;
  assign n57374 = ~n57371 & ~n57373;
  assign n57375 = n65014 & n57374;
  assign n57376 = pi1148 & ~n57375;
  assign n57377 = ~n57370 & n57376;
  assign n57378 = ~pi211 & ~n54784;
  assign n57379 = n52475 & ~n57378;
  assign n57380 = n52474 & ~n57371;
  assign n57381 = ~n57379 & ~n57380;
  assign n57382 = pi1147 & ~n57381;
  assign n57383 = pi1146 & ~n65570;
  assign n57384 = ~n48938 & n57383;
  assign n57385 = ~pi1148 & ~n57384;
  assign n57386 = ~n57382 & n57385;
  assign n57387 = pi230 & ~n57386;
  assign n57388 = pi230 & ~n57377;
  assign n57389 = ~n57386 & n57388;
  assign n57390 = ~n57377 & n57387;
  assign n57391 = ~n57366 & ~n65651;
  assign n57392 = pi1147 & n49471;
  assign n57393 = pi1091 & pi1145;
  assign n57394 = n39538 & ~n57393;
  assign n57395 = ~n57351 & n57394;
  assign n57396 = ~n57347 & ~n57395;
  assign n57397 = ~n57392 & ~n57396;
  assign n57398 = ~pi199 & ~n57393;
  assign n57399 = ~n57351 & n57398;
  assign n57400 = ~n57347 & ~n57399;
  assign n57401 = ~pi200 & ~n57392;
  assign n57402 = ~n57400 & n57401;
  assign n57403 = ~n57355 & ~n57402;
  assign n57404 = ~n57355 & ~n57397;
  assign n57405 = n65014 & ~n65652;
  assign n57406 = pi219 & ~n57346;
  assign n57407 = ~n57320 & ~n57352;
  assign n57408 = pi1091 & n53007;
  assign n57409 = ~pi219 & ~n57408;
  assign n57410 = ~n57407 & n57409;
  assign n57411 = ~n57406 & ~n57410;
  assign n57412 = ~pi211 & pi1147;
  assign n57413 = n50334 & n57412;
  assign n57414 = ~n65014 & ~n57413;
  assign n57415 = ~n57411 & n57414;
  assign n57416 = ~n57405 & ~n57415;
  assign n57417 = ~pi230 & ~n57416;
  assign n57418 = ~n54778 & ~n54836;
  assign n57419 = ~pi219 & ~n57418;
  assign n57420 = pi1147 & n50525;
  assign n57421 = ~pi200 & ~n53029;
  assign n57422 = n54940 & ~n57421;
  assign n57423 = ~n57420 & ~n57422;
  assign n57424 = ~n57419 & ~n57420;
  assign n57425 = ~n57422 & n57424;
  assign n57426 = ~n57419 & n57423;
  assign n57427 = n62455 & ~n65653;
  assign n57428 = ~n53007 & n56185;
  assign n57429 = pi219 & ~n57412;
  assign n57430 = ~n62455 & ~n57429;
  assign n57431 = ~n57428 & ~n57429;
  assign n57432 = ~n62455 & n57431;
  assign n57433 = ~n57428 & n57430;
  assign n57434 = pi230 & ~n65654;
  assign n57435 = ~n57427 & n57434;
  assign po428 = ~n57417 & ~n57435;
  assign n57437 = pi264 & ~n49247;
  assign n57438 = ~pi796 & n49247;
  assign n57439 = ~pi1091 & ~n57438;
  assign n57440 = ~pi1091 & ~n57437;
  assign n57441 = ~n57438 & n57440;
  assign n57442 = ~n57437 & n57439;
  assign n57443 = pi1091 & pi1142;
  assign n57444 = ~n65655 & ~n57443;
  assign n57445 = pi200 & ~n57444;
  assign n57446 = pi1091 & pi1141;
  assign n57447 = ~n65655 & ~n57446;
  assign n57448 = ~pi200 & ~n57447;
  assign n57449 = ~pi199 & ~n57448;
  assign n57450 = ~pi199 & ~n57445;
  assign n57451 = ~n57448 & n57450;
  assign n57452 = ~n57445 & n57449;
  assign n57453 = pi264 & ~n49236;
  assign n57454 = ~pi796 & n49236;
  assign n57455 = ~pi1091 & ~n57454;
  assign n57456 = ~pi1091 & ~n57453;
  assign n57457 = ~n57454 & n57456;
  assign n57458 = ~n57453 & n57455;
  assign n57459 = pi1091 & pi1143;
  assign n57460 = ~pi200 & n57459;
  assign n57461 = pi199 & ~n57460;
  assign n57462 = ~n65657 & n57461;
  assign n57463 = n65014 & ~n57462;
  assign n57464 = ~n65656 & n57463;
  assign n57465 = pi211 & ~n57444;
  assign n57466 = ~pi211 & ~n57447;
  assign n57467 = ~pi219 & ~n57466;
  assign n57468 = ~pi219 & ~n57465;
  assign n57469 = ~n57466 & n57468;
  assign n57470 = ~n57465 & n57467;
  assign n57471 = pi219 & ~n49812;
  assign n57472 = ~n53019 & ~n57471;
  assign n57473 = ~n65657 & ~n57472;
  assign n57474 = ~n65014 & ~n57473;
  assign n57475 = ~n65658 & n57474;
  assign n57476 = ~n57464 & ~n57475;
  assign n57477 = ~pi230 & ~n57476;
  assign n57478 = ~pi199 & pi1141;
  assign n57479 = n53024 & ~n57478;
  assign n57480 = ~n52550 & ~n57479;
  assign n57481 = n65014 & ~n57480;
  assign n57482 = ~pi211 & pi1141;
  assign n57483 = ~pi219 & ~n57482;
  assign n57484 = ~pi219 & ~n52559;
  assign n57485 = ~n57482 & n57484;
  assign n57486 = ~n52559 & n57483;
  assign n57487 = ~n53019 & ~n65659;
  assign n57488 = ~n65014 & ~n57487;
  assign n57489 = pi230 & ~n57488;
  assign n57490 = pi230 & ~n57481;
  assign n57491 = ~n57488 & n57490;
  assign n57492 = ~n57481 & n57489;
  assign n57493 = ~n57477 & ~n65660;
  assign n57494 = pi265 & ~n49247;
  assign n57495 = ~pi819 & n49247;
  assign n57496 = ~pi1091 & ~n57495;
  assign n57497 = ~pi1091 & ~n57494;
  assign n57498 = ~n57495 & n57497;
  assign n57499 = ~n57494 & n57496;
  assign n57500 = ~n57459 & ~n65661;
  assign n57501 = pi200 & ~n57500;
  assign n57502 = ~n57443 & ~n65661;
  assign n57503 = ~pi200 & ~n57502;
  assign n57504 = ~pi199 & ~n57503;
  assign n57505 = ~pi199 & ~n57501;
  assign n57506 = ~n57503 & n57505;
  assign n57507 = ~n57501 & n57504;
  assign n57508 = pi265 & ~n49236;
  assign n57509 = ~pi819 & n49236;
  assign n57510 = ~pi1091 & ~n57509;
  assign n57511 = ~pi1091 & ~n57508;
  assign n57512 = ~n57509 & n57511;
  assign n57513 = ~n57508 & n57510;
  assign n57514 = pi1091 & pi1144;
  assign n57515 = ~pi200 & n57514;
  assign n57516 = pi199 & ~n57515;
  assign n57517 = ~n65663 & n57516;
  assign n57518 = n65014 & ~n57517;
  assign n57519 = ~n65662 & n57518;
  assign n57520 = pi211 & ~n57500;
  assign n57521 = ~pi211 & ~n57502;
  assign n57522 = ~pi219 & ~n57521;
  assign n57523 = ~pi219 & ~n57520;
  assign n57524 = ~n57521 & n57523;
  assign n57525 = ~n57520 & n57522;
  assign n57526 = ~n55692 & ~n57471;
  assign n57527 = ~n65663 & ~n57526;
  assign n57528 = ~n65014 & ~n57527;
  assign n57529 = ~n65664 & n57528;
  assign n57530 = ~n57519 & ~n57529;
  assign n57531 = ~pi230 & ~n57530;
  assign n57532 = ~n52549 & n55697;
  assign n57533 = ~n52543 & ~n57532;
  assign n57534 = n65014 & ~n57533;
  assign n57535 = ~pi219 & ~n52524;
  assign n57536 = ~n52567 & n57535;
  assign n57537 = ~n55692 & ~n57536;
  assign n57538 = ~n65014 & ~n57537;
  assign n57539 = pi230 & ~n57538;
  assign n57540 = pi230 & ~n57534;
  assign n57541 = ~n57538 & n57540;
  assign n57542 = ~n57534 & n57539;
  assign n57543 = ~n57531 & ~n65665;
  assign n57544 = ~pi211 & pi1136;
  assign n57545 = pi219 & ~n57544;
  assign n57546 = pi211 & ~pi1135;
  assign n57547 = ~n57545 & ~n57546;
  assign n57548 = ~n39421 & n57547;
  assign n57549 = pi299 & n57548;
  assign n57550 = pi199 & pi1136;
  assign n57551 = ~pi200 & ~n57550;
  assign n57552 = ~pi199 & pi1135;
  assign n57553 = pi200 & ~n57552;
  assign n57554 = ~pi299 & ~n57553;
  assign n57555 = ~pi299 & ~n57551;
  assign n57556 = ~n57553 & n57555;
  assign n57557 = ~n57551 & n57554;
  assign n57558 = ~n57549 & ~n65666;
  assign n57559 = n62455 & ~n57558;
  assign n57560 = ~n62455 & n57548;
  assign n57561 = pi230 & ~n57560;
  assign n57562 = ~n57559 & n57561;
  assign n57563 = ~pi948 & n49247;
  assign n57564 = ~pi266 & ~n49247;
  assign n57565 = ~pi1091 & ~n57564;
  assign n57566 = ~pi1091 & ~n57563;
  assign n57567 = ~n57564 & n57566;
  assign n57568 = ~n57563 & n57565;
  assign n57569 = ~pi199 & ~n65667;
  assign n57570 = pi1091 & pi1136;
  assign n57571 = ~pi948 & n49236;
  assign n57572 = ~pi266 & ~n49236;
  assign n57573 = ~pi1091 & ~n57572;
  assign n57574 = ~pi1091 & ~n57571;
  assign n57575 = ~n57572 & n57574;
  assign n57576 = ~n57571 & n57573;
  assign n57577 = pi199 & ~n65668;
  assign n57578 = ~n57570 & n57577;
  assign n57579 = ~n57569 & ~n57578;
  assign n57580 = ~pi200 & n57579;
  assign n57581 = pi1091 & pi1135;
  assign n57582 = n57569 & ~n57581;
  assign n57583 = pi200 & ~n57577;
  assign n57584 = ~n57582 & n57583;
  assign n57585 = ~n57580 & ~n57584;
  assign n57586 = n65014 & ~n57585;
  assign n57587 = ~n57471 & ~n57545;
  assign n57588 = ~n65668 & ~n57587;
  assign n57589 = ~n65014 & ~n57588;
  assign n57590 = ~pi219 & ~n65667;
  assign n57591 = pi1135 & n49802;
  assign n57592 = n57590 & ~n57591;
  assign n57593 = n57589 & ~n57592;
  assign n57594 = ~pi230 & ~n57593;
  assign n57595 = ~n57586 & n57594;
  assign n57596 = ~n57562 & ~n57595;
  assign n57597 = ~pi1134 & ~n57596;
  assign n57598 = ~n65014 & n57547;
  assign n57599 = n49457 & ~n57550;
  assign n57600 = ~n57553 & ~n57599;
  assign n57601 = n65014 & n57600;
  assign n57602 = pi230 & ~n57601;
  assign n57603 = pi230 & ~n57598;
  assign n57604 = ~n57601 & n57603;
  assign n57605 = ~n57598 & n57602;
  assign n57606 = ~pi199 & pi1091;
  assign n57607 = ~n57579 & ~n57606;
  assign n57608 = ~pi200 & ~n57607;
  assign n57609 = ~n57584 & ~n57608;
  assign n57610 = n65014 & ~n57609;
  assign n57611 = pi1091 & ~n57546;
  assign n57612 = n57590 & ~n57611;
  assign n57613 = n57589 & ~n57612;
  assign n57614 = ~pi230 & ~n57613;
  assign n57615 = ~n57610 & n57614;
  assign n57616 = ~n65669 & ~n57615;
  assign n57617 = pi1134 & ~n57616;
  assign po423 = ~n57597 & ~n57617;
  assign n57619 = pi211 & pi1137;
  assign n57620 = ~n57544 & ~n57619;
  assign n57621 = pi1091 & ~n57620;
  assign n57622 = n52475 & ~n57621;
  assign n57623 = ~pi200 & n57570;
  assign n57624 = pi1137 & n49493;
  assign n57625 = ~n57623 & ~n57624;
  assign n57626 = n52474 & n57625;
  assign n57627 = ~n57622 & ~n57626;
  assign n57628 = pi269 & ~n49247;
  assign n57629 = ~pi817 & n49247;
  assign n57630 = ~pi1091 & ~n57629;
  assign n57631 = ~pi1091 & ~n57628;
  assign n57632 = ~n57629 & n57631;
  assign n57633 = ~n57628 & n57630;
  assign n57634 = ~n57627 & ~n65670;
  assign n57635 = pi219 & ~n65014;
  assign n57636 = pi1138 & n49812;
  assign n57637 = n57635 & ~n57636;
  assign n57638 = ~pi200 & pi1091;
  assign n57639 = pi1138 & n57638;
  assign n57640 = pi199 & ~n57639;
  assign n57641 = n65014 & n57640;
  assign n57642 = ~n57637 & ~n57641;
  assign n57643 = pi269 & ~n49236;
  assign n57644 = ~pi817 & n49236;
  assign n57645 = ~pi1091 & ~n57644;
  assign n57646 = ~pi1091 & ~n57643;
  assign n57647 = ~n57644 & n57646;
  assign n57648 = ~n57643 & n57645;
  assign n57649 = ~n57642 & ~n65671;
  assign n57650 = ~n57634 & ~n57649;
  assign n57651 = ~pi230 & ~n57650;
  assign n57652 = ~pi199 & pi1137;
  assign n57653 = pi200 & ~n57652;
  assign n57654 = ~pi199 & pi1136;
  assign n57655 = pi199 & pi1138;
  assign n57656 = ~pi200 & ~n57655;
  assign n57657 = ~pi200 & ~n57654;
  assign n57658 = ~n57655 & n57657;
  assign n57659 = ~n57654 & n57656;
  assign n57660 = ~n57653 & ~n65672;
  assign n57661 = n65014 & ~n57660;
  assign n57662 = ~pi219 & ~n57620;
  assign n57663 = ~pi211 & pi1138;
  assign n57664 = pi219 & n57663;
  assign n57665 = ~n57662 & ~n57664;
  assign n57666 = ~n65014 & n57665;
  assign n57667 = ~n57661 & ~n57666;
  assign n57668 = pi230 & ~n57667;
  assign po426 = ~n57651 & ~n57668;
  assign n57670 = ~pi211 & pi1139;
  assign n57671 = pi211 & pi1140;
  assign n57672 = ~n57670 & ~n57671;
  assign n57673 = pi1091 & ~n57672;
  assign n57674 = n52475 & ~n57673;
  assign n57675 = pi1139 & n57638;
  assign n57676 = pi1091 & pi1140;
  assign n57677 = pi200 & n57676;
  assign n57678 = pi1140 & n49493;
  assign n57679 = ~n57675 & ~n65673;
  assign n57680 = n52474 & n57679;
  assign n57681 = ~n57674 & ~n57680;
  assign n57682 = pi270 & ~n49247;
  assign n57683 = ~pi805 & n49247;
  assign n57684 = ~pi1091 & ~n57683;
  assign n57685 = ~pi1091 & ~n57682;
  assign n57686 = ~n57683 & n57685;
  assign n57687 = ~n57682 & n57684;
  assign n57688 = ~n57681 & ~n65674;
  assign n57689 = n49812 & n57482;
  assign n57690 = pi1091 & n57482;
  assign n57691 = n57635 & ~n65675;
  assign n57692 = ~pi200 & n57446;
  assign n57693 = pi199 & ~n57692;
  assign n57694 = n65014 & n57693;
  assign n57695 = ~n57691 & ~n57694;
  assign n57696 = pi270 & ~n49236;
  assign n57697 = ~pi805 & n49236;
  assign n57698 = ~pi1091 & ~n57697;
  assign n57699 = ~pi1091 & ~n57696;
  assign n57700 = ~n57697 & n57699;
  assign n57701 = ~n57696 & n57698;
  assign n57702 = ~n57695 & ~n65676;
  assign n57703 = ~pi230 & ~n57702;
  assign n57704 = ~pi230 & ~n57688;
  assign n57705 = ~n57702 & n57704;
  assign n57706 = ~n57688 & n57703;
  assign n57707 = pi1140 & n48474;
  assign n57708 = pi199 & pi1141;
  assign n57709 = ~pi199 & pi1139;
  assign n57710 = ~n57708 & ~n57709;
  assign n57711 = ~pi200 & ~n57710;
  assign n57712 = ~pi199 & pi1140;
  assign n57713 = pi200 & ~n57712;
  assign n57714 = ~pi200 & ~n57709;
  assign n57715 = ~pi200 & ~n57708;
  assign n57716 = ~n57709 & n57715;
  assign n57717 = ~n57708 & n57714;
  assign n57718 = ~n57713 & ~n65678;
  assign n57719 = ~n57707 & ~n57711;
  assign n57720 = n65014 & ~n65679;
  assign n57721 = ~pi219 & ~n57672;
  assign n57722 = pi1141 & n39423;
  assign n57723 = pi219 & n57482;
  assign n57724 = pi219 & ~n57482;
  assign n57725 = ~pi219 & n57672;
  assign n57726 = ~n57724 & ~n57725;
  assign n57727 = ~n57721 & ~n65680;
  assign n57728 = ~n65014 & ~n65681;
  assign n57729 = pi230 & ~n57728;
  assign n57730 = pi230 & ~n57720;
  assign n57731 = ~n57728 & n57730;
  assign n57732 = ~n57720 & n57729;
  assign n57733 = ~n65677 & ~n65682;
  assign n57734 = pi274 & ~n49247;
  assign n57735 = ~pi659 & n49247;
  assign n57736 = ~pi1091 & ~n57735;
  assign n57737 = ~pi1091 & ~n57734;
  assign n57738 = ~n57735 & n57737;
  assign n57739 = ~n57734 & n57736;
  assign n57740 = ~n57459 & ~n65683;
  assign n57741 = ~pi211 & ~n57740;
  assign n57742 = ~n57514 & ~n65683;
  assign n57743 = pi211 & ~n57742;
  assign n57744 = ~pi219 & ~n57743;
  assign n57745 = ~pi219 & ~n57741;
  assign n57746 = ~n57743 & n57745;
  assign n57747 = ~n57741 & n57744;
  assign n57748 = pi274 & ~n49236;
  assign n57749 = ~pi659 & n49236;
  assign n57750 = ~pi1091 & ~n57749;
  assign n57751 = ~pi1091 & ~n57748;
  assign n57752 = ~n57749 & n57751;
  assign n57753 = ~n57748 & n57750;
  assign n57754 = pi219 & ~n57408;
  assign n57755 = ~n65685 & n57754;
  assign n57756 = ~n65014 & ~n57755;
  assign n57757 = ~n65684 & n57756;
  assign n57758 = ~pi200 & ~n57740;
  assign n57759 = pi200 & ~n57742;
  assign n57760 = ~pi199 & ~n57759;
  assign n57761 = ~pi199 & ~n57758;
  assign n57762 = ~n57759 & n57761;
  assign n57763 = ~n57758 & n57760;
  assign n57764 = ~pi200 & n57393;
  assign n57765 = pi199 & ~n57764;
  assign n57766 = ~n65685 & n57765;
  assign n57767 = n65014 & ~n57766;
  assign n57768 = ~n65686 & n57767;
  assign n57769 = ~pi230 & ~n57768;
  assign n57770 = ~pi230 & ~n57757;
  assign n57771 = ~n57768 & n57770;
  assign n57772 = ~n57757 & n57769;
  assign n57773 = ~pi219 & ~n52522;
  assign n57774 = ~n53008 & n57773;
  assign n57775 = ~n54773 & ~n57774;
  assign n57776 = ~n50523 & ~n54778;
  assign n57777 = ~n57774 & ~n57776;
  assign n57778 = ~n52542 & n54946;
  assign n57779 = n55695 & ~n57778;
  assign n57780 = ~n57777 & ~n57779;
  assign n57781 = n62455 & ~n57780;
  assign n57782 = pi230 & ~n57781;
  assign n57783 = ~n57775 & n57782;
  assign po431 = ~n65687 & ~n57783;
  assign n57785 = ~pi276 & ~n49237;
  assign n57786 = n49239 & ~n57785;
  assign n57787 = ~n57320 & n57635;
  assign n57788 = pi199 & ~n57325;
  assign n57789 = n65014 & n57788;
  assign n57790 = ~n57787 & ~n57789;
  assign n57791 = ~n57786 & ~n57790;
  assign n57792 = ~pi276 & ~n49248;
  assign n57793 = n57348 & ~n57792;
  assign n57794 = ~n52525 & ~n54762;
  assign n57795 = pi1091 & ~n57794;
  assign n57796 = n52475 & ~n57795;
  assign n57797 = pi1145 & n49493;
  assign n57798 = ~n57515 & ~n57797;
  assign n57799 = n52474 & n57798;
  assign n57800 = ~n57796 & ~n57799;
  assign n57801 = ~n57793 & ~n57800;
  assign n57802 = ~pi230 & ~n57801;
  assign n57803 = ~pi230 & ~n57791;
  assign n57804 = ~n57801 & n57803;
  assign n57805 = ~n57791 & n57802;
  assign n57806 = pi1146 & n39423;
  assign n57807 = pi219 & n54761;
  assign n57808 = ~pi219 & ~n57794;
  assign n57809 = ~n65689 & ~n57808;
  assign n57810 = ~n65014 & n57809;
  assign n57811 = ~n52540 & n55921;
  assign n57812 = ~n54948 & ~n57811;
  assign n57813 = n65014 & ~n57812;
  assign n57814 = pi230 & ~n57813;
  assign n57815 = pi230 & ~n57810;
  assign n57816 = ~n57813 & n57815;
  assign n57817 = ~n57810 & n57814;
  assign n57818 = ~n65688 & ~n65690;
  assign n57819 = pi277 & ~n49247;
  assign n57820 = ~pi820 & n49247;
  assign n57821 = ~pi1091 & ~n57820;
  assign n57822 = ~pi1091 & ~n57819;
  assign n57823 = ~n57820 & n57822;
  assign n57824 = ~n57819 & n57821;
  assign n57825 = ~n57446 & ~n65691;
  assign n57826 = pi200 & ~n57825;
  assign n57827 = ~n57676 & ~n65691;
  assign n57828 = ~pi200 & ~n57827;
  assign n57829 = ~pi199 & ~n57828;
  assign n57830 = ~pi199 & ~n57826;
  assign n57831 = ~n57828 & n57830;
  assign n57832 = ~n57826 & n57829;
  assign n57833 = pi277 & ~n49236;
  assign n57834 = ~pi820 & n49236;
  assign n57835 = ~pi1091 & ~n57834;
  assign n57836 = ~pi1091 & ~n57833;
  assign n57837 = ~n57834 & n57836;
  assign n57838 = ~n57833 & n57835;
  assign n57839 = ~pi200 & n57443;
  assign n57840 = pi199 & ~n57839;
  assign n57841 = ~n65693 & n57840;
  assign n57842 = n65014 & ~n57841;
  assign n57843 = ~n65692 & n57842;
  assign n57844 = pi211 & ~n57825;
  assign n57845 = ~pi211 & ~n57827;
  assign n57846 = ~pi219 & ~n57845;
  assign n57847 = ~pi219 & ~n57844;
  assign n57848 = ~n57845 & n57847;
  assign n57849 = ~n57844 & n57846;
  assign n57850 = ~n52568 & ~n57471;
  assign n57851 = ~n65693 & ~n57850;
  assign n57852 = ~n65014 & ~n57851;
  assign n57853 = ~n65694 & n57852;
  assign n57854 = ~n57843 & ~n57853;
  assign n57855 = ~pi230 & ~n57854;
  assign n57856 = n52539 & ~n57712;
  assign n57857 = pi200 & ~n57478;
  assign n57858 = ~n57856 & ~n57857;
  assign n57859 = n65014 & ~n57858;
  assign n57860 = ~pi211 & pi1140;
  assign n57861 = pi211 & pi1141;
  assign n57862 = ~pi219 & ~n57861;
  assign n57863 = ~pi219 & ~n57860;
  assign n57864 = ~n57861 & n57863;
  assign n57865 = ~n57860 & n57862;
  assign n57866 = ~n52568 & ~n65695;
  assign n57867 = ~n65014 & ~n57866;
  assign n57868 = pi230 & ~n57867;
  assign n57869 = pi230 & ~n57859;
  assign n57870 = ~n57867 & n57869;
  assign n57871 = ~n57859 & n57868;
  assign n57872 = ~n57855 & ~n65696;
  assign n57873 = ~pi976 & n49236;
  assign n57874 = ~pi278 & ~n49236;
  assign n57875 = ~pi1091 & ~n57874;
  assign n57876 = ~pi1091 & ~n57873;
  assign n57877 = ~n57874 & n57876;
  assign n57878 = ~n57873 & n57875;
  assign n57879 = pi199 & ~n65697;
  assign n57880 = pi1091 & ~pi1132;
  assign n57881 = pi278 & ~n49247;
  assign n57882 = pi976 & n49247;
  assign n57883 = ~pi1091 & ~n57882;
  assign n57884 = ~pi1091 & ~n57881;
  assign n57885 = ~n57882 & n57884;
  assign n57886 = ~n57881 & n57883;
  assign n57887 = ~n57880 & ~n65698;
  assign n57888 = ~pi199 & ~n57887;
  assign n57889 = ~n57879 & ~n57888;
  assign n57890 = ~pi200 & ~n57889;
  assign n57891 = pi1091 & ~pi1133;
  assign n57892 = ~n65698 & ~n57891;
  assign n57893 = ~pi199 & ~n57892;
  assign n57894 = ~n57879 & ~n57893;
  assign n57895 = pi200 & ~n57894;
  assign n57896 = ~pi299 & ~n57895;
  assign n57897 = ~n57890 & n57896;
  assign n57898 = pi219 & ~n65697;
  assign n57899 = pi211 & ~pi1133;
  assign n57900 = ~pi211 & ~pi1132;
  assign n57901 = ~pi211 & pi1132;
  assign n57902 = pi211 & pi1133;
  assign n57903 = ~n57901 & ~n57902;
  assign n57904 = ~n57899 & ~n57900;
  assign n57905 = pi1091 & n65699;
  assign n57906 = ~n65698 & ~n57905;
  assign n57907 = ~pi219 & ~n57906;
  assign n57908 = ~n57898 & ~n57907;
  assign n57909 = pi299 & n57908;
  assign n57910 = ~n57897 & ~n57909;
  assign n57911 = n62455 & ~n57910;
  assign n57912 = ~n62455 & n57908;
  assign n57913 = ~pi230 & ~n57912;
  assign n57914 = ~n57911 & n57913;
  assign n57915 = ~pi199 & pi1132;
  assign n57916 = ~pi200 & ~n57915;
  assign n57917 = ~pi199 & pi1133;
  assign n57918 = pi200 & ~n57917;
  assign n57919 = ~pi299 & ~n57918;
  assign n57920 = ~n57916 & n57919;
  assign n57921 = n50523 & ~n65699;
  assign n57922 = ~n57920 & ~n57921;
  assign n57923 = n62455 & ~n57922;
  assign n57924 = n50558 & ~n65699;
  assign n57925 = pi230 & ~n57924;
  assign n57926 = pi230 & ~n57923;
  assign n57927 = ~n57924 & n57926;
  assign n57928 = ~n57923 & n57925;
  assign n57929 = ~n57914 & ~n65700;
  assign n57930 = ~pi1134 & ~n57929;
  assign n57931 = ~pi219 & n65699;
  assign n57932 = ~n55050 & ~n57931;
  assign n57933 = n39538 & ~n57915;
  assign n57934 = n57919 & ~n57933;
  assign n57935 = ~n50243 & ~n57921;
  assign n57936 = ~n57934 & n57935;
  assign n57937 = n62455 & ~n57936;
  assign n57938 = pi230 & ~n57937;
  assign n57939 = ~n57932 & n57938;
  assign n57940 = ~n49471 & n57890;
  assign n57941 = n57896 & ~n57940;
  assign n57942 = n48495 & n49812;
  assign n57943 = ~n57909 & ~n57942;
  assign n57944 = ~n57941 & n57943;
  assign n57945 = n62455 & ~n57944;
  assign n57946 = ~n57360 & n57913;
  assign n57947 = ~n57945 & n57946;
  assign n57948 = ~n57939 & ~n57947;
  assign n57949 = pi1134 & ~n57948;
  assign po435 = ~n57930 & ~n57949;
  assign n57951 = ~pi958 & n49236;
  assign n57952 = ~pi279 & ~n49236;
  assign n57953 = ~pi1091 & ~n57952;
  assign n57954 = ~pi1091 & ~n57951;
  assign n57955 = ~n57952 & n57954;
  assign n57956 = ~n57951 & n57953;
  assign n57957 = pi1135 & n57638;
  assign n57958 = ~n65701 & ~n57957;
  assign n57959 = pi199 & ~n57958;
  assign n57960 = pi279 & ~n49247;
  assign n57961 = pi958 & n49247;
  assign n57962 = ~pi1091 & ~n57961;
  assign n57963 = ~pi1091 & ~n57960;
  assign n57964 = ~n57961 & n57963;
  assign n57965 = ~n57960 & n57962;
  assign n57966 = ~pi1133 & n57638;
  assign n57967 = ~pi199 & ~n57966;
  assign n57968 = ~n65702 & n57967;
  assign n57969 = ~n57959 & ~n57968;
  assign n57970 = n65014 & ~n57969;
  assign n57971 = ~n49493 & n57970;
  assign n57972 = ~n49802 & ~n57891;
  assign n57973 = ~n65702 & n57972;
  assign n57974 = ~pi219 & ~n57973;
  assign n57975 = pi1135 & n49812;
  assign n57976 = pi219 & ~n57975;
  assign n57977 = ~n65701 & n57976;
  assign n57978 = ~n65014 & ~n57977;
  assign n57979 = ~n57974 & n57978;
  assign n57980 = ~pi230 & ~n57979;
  assign n57981 = ~n57971 & n57980;
  assign n57982 = pi199 & pi1135;
  assign n57983 = ~n57917 & ~n57982;
  assign n57984 = n49461 & ~n57983;
  assign n57985 = pi1135 & n39423;
  assign n57986 = ~pi211 & ~pi1133;
  assign n57987 = ~pi219 & ~n57986;
  assign n57988 = ~pi211 & n57987;
  assign n57989 = ~n57985 & ~n57988;
  assign n57990 = pi299 & ~n57989;
  assign n57991 = ~n57984 & ~n57990;
  assign n57992 = n62455 & ~n57991;
  assign n57993 = ~n62455 & ~n57989;
  assign n57994 = pi230 & ~n57993;
  assign n57995 = ~n57992 & n57994;
  assign n57996 = ~n57981 & ~n57995;
  assign n57997 = ~pi1134 & ~n57996;
  assign n57998 = ~pi1133 & n39538;
  assign n57999 = ~pi200 & pi1135;
  assign n58000 = pi199 & ~n57999;
  assign n58001 = ~n57998 & ~n58000;
  assign n58002 = n65014 & n58001;
  assign n58003 = ~n57985 & ~n57987;
  assign n58004 = ~n65014 & ~n58003;
  assign n58005 = pi230 & ~n58004;
  assign n58006 = n65014 & ~n58001;
  assign n58007 = ~n65014 & n58003;
  assign n58008 = ~n58006 & ~n58007;
  assign n58009 = pi230 & ~n58008;
  assign n58010 = ~n58002 & n58005;
  assign n58011 = pi1091 & ~n57986;
  assign n58012 = n52475 & n58011;
  assign n58013 = ~n57970 & ~n58012;
  assign n58014 = n57980 & n58013;
  assign n58015 = ~n65703 & ~n58014;
  assign n58016 = pi1134 & ~n58015;
  assign po436 = ~n57997 & ~n58016;
  assign n58018 = pi914 & n49247;
  assign n58019 = ~pi280 & ~n49247;
  assign n58020 = ~pi1091 & ~n58019;
  assign n58021 = ~pi1091 & ~n58018;
  assign n58022 = ~n58019 & n58021;
  assign n58023 = ~n58018 & n58020;
  assign n58024 = pi200 & pi1136;
  assign n58025 = pi1091 & ~n57999;
  assign n58026 = ~n58024 & n58025;
  assign n58027 = ~pi199 & ~n58026;
  assign n58028 = ~n65704 & n58027;
  assign n58029 = pi280 & ~n49236;
  assign n58030 = ~pi914 & n49236;
  assign n58031 = ~pi1091 & ~n58030;
  assign n58032 = ~pi1091 & ~n58029;
  assign n58033 = ~n58030 & n58032;
  assign n58034 = ~n58029 & n58031;
  assign n58035 = pi1137 & n57638;
  assign n58036 = ~n65705 & ~n58035;
  assign n58037 = pi199 & ~n58036;
  assign n58038 = ~n58028 & ~n58037;
  assign n58039 = n65014 & ~n58038;
  assign n58040 = ~pi211 & pi1135;
  assign n58041 = pi211 & pi1136;
  assign n58042 = ~n58040 & ~n58041;
  assign n58043 = pi1091 & n58042;
  assign n58044 = ~n65704 & ~n58043;
  assign n58045 = ~pi219 & ~n58044;
  assign n58046 = ~pi211 & pi1137;
  assign n58047 = pi219 & ~n58046;
  assign n58048 = ~n57471 & ~n58047;
  assign n58049 = ~n65705 & ~n58048;
  assign n58050 = ~n65014 & ~n58049;
  assign n58051 = ~n58045 & n58050;
  assign n58052 = ~n58045 & ~n58049;
  assign n58053 = ~n65014 & ~n58052;
  assign n58054 = n65014 & ~n58037;
  assign n58055 = n65014 & ~n58028;
  assign n58056 = ~n58037 & n58055;
  assign n58057 = ~n58028 & n58054;
  assign n58058 = ~n58053 & ~n65706;
  assign n58059 = ~n58039 & ~n58051;
  assign n58060 = ~pi230 & ~n65707;
  assign n58061 = ~pi219 & n58042;
  assign n58062 = ~n58047 & ~n58061;
  assign n58063 = ~n65014 & n58062;
  assign n58064 = pi200 & ~n57654;
  assign n58065 = pi199 & pi1137;
  assign n58066 = ~pi200 & ~n57552;
  assign n58067 = ~n58065 & n58066;
  assign n58068 = ~n58064 & ~n58067;
  assign n58069 = n65014 & n58068;
  assign n58070 = pi230 & ~n58069;
  assign n58071 = pi230 & ~n58063;
  assign n58072 = ~n58069 & n58071;
  assign n58073 = ~n58063 & n58070;
  assign n58074 = ~pi230 & n65707;
  assign n58075 = n65014 & ~n58068;
  assign n58076 = ~n65014 & ~n58062;
  assign n58077 = pi230 & ~n58076;
  assign n58078 = ~n58075 & n58077;
  assign n58079 = ~n58074 & ~n58078;
  assign n58080 = ~n58060 & ~n65708;
  assign n58081 = pi211 & pi1138;
  assign n58082 = ~n58046 & ~n58081;
  assign n58083 = pi1091 & ~n58082;
  assign n58084 = n52475 & ~n58083;
  assign n58085 = pi1138 & n49493;
  assign n58086 = ~n58035 & ~n58085;
  assign n58087 = n52474 & n58086;
  assign n58088 = ~n58084 & ~n58087;
  assign n58089 = pi281 & ~n49247;
  assign n58090 = ~pi830 & n49247;
  assign n58091 = ~pi1091 & ~n58090;
  assign n58092 = ~pi1091 & ~n58089;
  assign n58093 = ~n58090 & n58092;
  assign n58094 = ~n58089 & n58091;
  assign n58095 = ~n58088 & ~n65710;
  assign n58096 = pi1139 & n49812;
  assign n58097 = n57635 & ~n58096;
  assign n58098 = pi199 & ~n57675;
  assign n58099 = n65014 & n58098;
  assign n58100 = ~n58097 & ~n58099;
  assign n58101 = pi281 & ~n49236;
  assign n58102 = ~pi830 & n49236;
  assign n58103 = ~pi1091 & ~n58102;
  assign n58104 = ~pi1091 & ~n58101;
  assign n58105 = ~n58102 & n58104;
  assign n58106 = ~n58101 & n58103;
  assign n58107 = ~n58100 & ~n65711;
  assign n58108 = ~n58095 & ~n58107;
  assign n58109 = ~pi230 & ~n58108;
  assign n58110 = ~pi199 & pi1138;
  assign n58111 = pi200 & ~n58110;
  assign n58112 = pi199 & pi1139;
  assign n58113 = ~pi200 & ~n57652;
  assign n58114 = ~n58112 & n58113;
  assign n58115 = ~n58111 & ~n58114;
  assign n58116 = n65014 & ~n58115;
  assign n58117 = pi219 & n57670;
  assign n58118 = ~pi219 & ~n58082;
  assign n58119 = ~n58117 & ~n58118;
  assign n58120 = ~n65014 & n58119;
  assign n58121 = ~n58116 & ~n58120;
  assign n58122 = pi230 & ~n58121;
  assign po438 = ~n58109 & ~n58122;
  assign n58124 = pi211 & pi1139;
  assign n58125 = ~n57663 & ~n58124;
  assign n58126 = pi1091 & ~n58125;
  assign n58127 = n52475 & ~n58126;
  assign n58128 = pi1139 & n49493;
  assign n58129 = ~n57639 & ~n58128;
  assign n58130 = n52474 & n58129;
  assign n58131 = ~n58127 & ~n58130;
  assign n58132 = pi282 & ~n49247;
  assign n58133 = ~pi836 & n49247;
  assign n58134 = ~pi1091 & ~n58133;
  assign n58135 = ~pi1091 & ~n58132;
  assign n58136 = ~n58133 & n58135;
  assign n58137 = ~n58132 & n58134;
  assign n58138 = ~n58131 & ~n65712;
  assign n58139 = pi1140 & n49812;
  assign n58140 = n57635 & ~n58139;
  assign n58141 = ~pi200 & n57676;
  assign n58142 = pi199 & ~n58141;
  assign n58143 = n65014 & n58142;
  assign n58144 = ~n58140 & ~n58143;
  assign n58145 = pi282 & ~n49236;
  assign n58146 = ~pi836 & n49236;
  assign n58147 = ~pi1091 & ~n58146;
  assign n58148 = ~pi1091 & ~n58145;
  assign n58149 = ~n58146 & n58148;
  assign n58150 = ~n58145 & n58147;
  assign n58151 = ~n58144 & ~n65713;
  assign n58152 = ~n58138 & ~n58151;
  assign n58153 = ~pi230 & ~n58152;
  assign n58154 = pi200 & ~n57709;
  assign n58155 = pi199 & pi1140;
  assign n58156 = ~pi200 & ~n58110;
  assign n58157 = ~n58155 & n58156;
  assign n58158 = ~n58154 & ~n58157;
  assign n58159 = n65014 & ~n58158;
  assign n58160 = pi219 & n57860;
  assign n58161 = ~pi219 & ~n58125;
  assign n58162 = ~n58160 & ~n58161;
  assign n58163 = ~n65014 & n58162;
  assign n58164 = ~n58159 & ~n58163;
  assign n58165 = pi230 & ~n58164;
  assign po439 = ~n58153 & ~n58165;
  assign n58167 = pi336 & ~n48171;
  assign n58168 = pi1070 & n48171;
  assign n58169 = ~n58167 & ~n58168;
  assign n58170 = pi337 & ~n48171;
  assign n58171 = pi1044 & n48171;
  assign n58172 = ~n58170 & ~n58171;
  assign n58173 = pi342 & ~n65040;
  assign n58174 = pi1049 & n65040;
  assign n58175 = ~n58173 & ~n58174;
  assign n58176 = pi343 & ~n65040;
  assign n58177 = pi1062 & n65040;
  assign n58178 = ~n58176 & ~n58177;
  assign n58179 = pi345 & ~n65040;
  assign n58180 = pi1039 & n65040;
  assign n58181 = ~n58179 & ~n58180;
  assign n58182 = pi346 & ~n65040;
  assign n58183 = pi1067 & n65040;
  assign n58184 = ~n58182 & ~n58183;
  assign n58185 = pi347 & ~n65040;
  assign n58186 = pi1055 & n65040;
  assign n58187 = ~n58185 & ~n58186;
  assign n58188 = pi348 & ~n65040;
  assign n58189 = pi1087 & n65040;
  assign n58190 = ~n58188 & ~n58189;
  assign n58191 = pi350 & ~n65040;
  assign n58192 = pi1035 & n65040;
  assign n58193 = ~n58191 & ~n58192;
  assign n58194 = pi351 & ~n65040;
  assign n58195 = pi1079 & n65040;
  assign n58196 = ~n58194 & ~n58195;
  assign n58197 = pi354 & ~n65040;
  assign n58198 = pi1045 & n65040;
  assign n58199 = ~n58197 & ~n58198;
  assign n58200 = pi355 & ~n65040;
  assign n58201 = pi1084 & n65040;
  assign n58202 = ~n58200 & ~n58201;
  assign n58203 = pi356 & ~n65040;
  assign n58204 = pi1081 & n65040;
  assign n58205 = ~n58203 & ~n58204;
  assign n58206 = pi357 & ~n65040;
  assign n58207 = pi1076 & n65040;
  assign n58208 = ~n58206 & ~n58207;
  assign n58209 = pi358 & ~n65040;
  assign n58210 = pi1071 & n65040;
  assign n58211 = ~n58209 & ~n58210;
  assign n58212 = pi359 & ~n65040;
  assign n58213 = pi1068 & n65040;
  assign n58214 = ~n58212 & ~n58213;
  assign n58215 = pi360 & ~n65040;
  assign n58216 = pi1042 & n65040;
  assign n58217 = ~n58215 & ~n58216;
  assign n58218 = pi361 & ~n65040;
  assign n58219 = pi1059 & n65040;
  assign n58220 = ~n58218 & ~n58219;
  assign n58221 = pi362 & ~n65040;
  assign n58222 = pi1070 & n65040;
  assign n58223 = ~n58221 & ~n58222;
  assign n58224 = pi363 & ~n48171;
  assign n58225 = pi1049 & n48171;
  assign n58226 = ~n58224 & ~n58225;
  assign n58227 = pi364 & ~n48171;
  assign n58228 = pi1062 & n48171;
  assign n58229 = ~n58227 & ~n58228;
  assign n58230 = pi367 & ~n48171;
  assign n58231 = pi1039 & n48171;
  assign n58232 = ~n58230 & ~n58231;
  assign n58233 = pi368 & ~n48171;
  assign n58234 = pi1067 & n48171;
  assign n58235 = ~n58233 & ~n58234;
  assign n58236 = pi370 & ~n48171;
  assign n58237 = pi1055 & n48171;
  assign n58238 = ~n58236 & ~n58237;
  assign n58239 = pi373 & ~n48171;
  assign n58240 = pi1087 & n48171;
  assign n58241 = ~n58239 & ~n58240;
  assign n58242 = pi374 & ~n48171;
  assign n58243 = pi1035 & n48171;
  assign n58244 = ~n58242 & ~n58243;
  assign n58245 = pi376 & ~n48171;
  assign n58246 = pi1079 & n48171;
  assign n58247 = ~n58245 & ~n58246;
  assign n58248 = pi379 & ~n48171;
  assign n58249 = pi1045 & n48171;
  assign n58250 = ~n58248 & ~n58249;
  assign n58251 = pi380 & ~n48171;
  assign n58252 = pi1084 & n48171;
  assign n58253 = ~n58251 & ~n58252;
  assign n58254 = pi381 & ~n48171;
  assign n58255 = pi1081 & n48171;
  assign n58256 = ~n58254 & ~n58255;
  assign n58257 = pi382 & ~n48171;
  assign n58258 = pi1076 & n48171;
  assign n58259 = ~n58257 & ~n58258;
  assign n58260 = pi383 & ~n48171;
  assign n58261 = pi1071 & n48171;
  assign n58262 = ~n58260 & ~n58261;
  assign n58263 = pi384 & ~n48171;
  assign n58264 = pi1068 & n48171;
  assign n58265 = ~n58263 & ~n58264;
  assign n58266 = pi385 & ~n48171;
  assign n58267 = pi1042 & n48171;
  assign n58268 = ~n58266 & ~n58267;
  assign n58269 = pi386 & ~n48171;
  assign n58270 = pi1059 & n48171;
  assign n58271 = ~n58269 & ~n58270;
  assign n58272 = pi387 & ~n48171;
  assign n58273 = pi1053 & n48171;
  assign n58274 = ~n58272 & ~n58273;
  assign n58275 = pi388 & ~n48171;
  assign n58276 = pi1037 & n48171;
  assign n58277 = ~n58275 & ~n58276;
  assign n58278 = pi389 & ~n48171;
  assign n58279 = pi1036 & n48171;
  assign n58280 = ~n58278 & ~n58279;
  assign n58281 = pi390 & ~n65041;
  assign n58282 = pi1049 & n65041;
  assign n58283 = ~n58281 & ~n58282;
  assign n58284 = pi391 & ~n65041;
  assign n58285 = pi1062 & n65041;
  assign n58286 = ~n58284 & ~n58285;
  assign n58287 = pi392 & ~n65041;
  assign n58288 = pi1039 & n65041;
  assign n58289 = ~n58287 & ~n58288;
  assign n58290 = pi393 & ~n65041;
  assign n58291 = pi1067 & n65041;
  assign n58292 = ~n58290 & ~n58291;
  assign n58293 = pi395 & ~n65041;
  assign n58294 = pi1055 & n65041;
  assign n58295 = ~n58293 & ~n58294;
  assign n58296 = pi398 & ~n65041;
  assign n58297 = pi1087 & n65041;
  assign n58298 = ~n58296 & ~n58297;
  assign n58299 = pi400 & ~n65041;
  assign n58300 = pi1035 & n65041;
  assign n58301 = ~n58299 & ~n58300;
  assign n58302 = pi401 & ~n65041;
  assign n58303 = pi1079 & n65041;
  assign n58304 = ~n58302 & ~n58303;
  assign n58305 = pi403 & ~n65041;
  assign n58306 = pi1045 & n65041;
  assign n58307 = ~n58305 & ~n58306;
  assign n58308 = pi404 & ~n65041;
  assign n58309 = pi1084 & n65041;
  assign n58310 = ~n58308 & ~n58309;
  assign n58311 = pi405 & ~n65041;
  assign n58312 = pi1081 & n65041;
  assign n58313 = ~n58311 & ~n58312;
  assign n58314 = pi406 & ~n65041;
  assign n58315 = pi1076 & n65041;
  assign n58316 = ~n58314 & ~n58315;
  assign n58317 = pi407 & ~n65041;
  assign n58318 = pi1071 & n65041;
  assign n58319 = ~n58317 & ~n58318;
  assign n58320 = pi408 & ~n65041;
  assign n58321 = pi1068 & n65041;
  assign n58322 = ~n58320 & ~n58321;
  assign n58323 = pi409 & ~n65041;
  assign n58324 = pi1042 & n65041;
  assign n58325 = ~n58323 & ~n58324;
  assign n58326 = pi410 & ~n65041;
  assign n58327 = pi1059 & n65041;
  assign n58328 = ~n58326 & ~n58327;
  assign n58329 = pi411 & ~n65041;
  assign n58330 = pi1053 & n65041;
  assign n58331 = ~n58329 & ~n58330;
  assign n58332 = pi412 & ~n65041;
  assign n58333 = pi1037 & n65041;
  assign n58334 = ~n58332 & ~n58333;
  assign n58335 = pi413 & ~n65041;
  assign n58336 = pi1036 & n65041;
  assign n58337 = ~n58335 & ~n58336;
  assign n58338 = pi414 & ~n48354;
  assign n58339 = pi1049 & n48354;
  assign n58340 = ~n58338 & ~n58339;
  assign n58341 = pi415 & ~n48354;
  assign n58342 = pi1062 & n48354;
  assign n58343 = ~n58341 & ~n58342;
  assign n58344 = pi417 & ~n48354;
  assign n58345 = pi1039 & n48354;
  assign n58346 = ~n58344 & ~n58345;
  assign n58347 = pi418 & ~n48354;
  assign n58348 = pi1067 & n48354;
  assign n58349 = ~n58347 & ~n58348;
  assign n58350 = pi420 & ~n48354;
  assign n58351 = pi1055 & n48354;
  assign n58352 = ~n58350 & ~n58351;
  assign n58353 = pi423 & ~n48354;
  assign n58354 = pi1087 & n48354;
  assign n58355 = ~n58353 & ~n58354;
  assign n58356 = pi425 & ~n48354;
  assign n58357 = pi1035 & n48354;
  assign n58358 = ~n58356 & ~n58357;
  assign n58359 = pi426 & ~n48354;
  assign n58360 = pi1079 & n48354;
  assign n58361 = ~n58359 & ~n58360;
  assign n58362 = pi428 & ~n48354;
  assign n58363 = pi1045 & n48354;
  assign n58364 = ~n58362 & ~n58363;
  assign n58365 = pi429 & ~n48354;
  assign n58366 = pi1084 & n48354;
  assign n58367 = ~n58365 & ~n58366;
  assign n58368 = pi430 & ~n48354;
  assign n58369 = pi1076 & n48354;
  assign n58370 = ~n58368 & ~n58369;
  assign n58371 = pi431 & ~n48354;
  assign n58372 = pi1071 & n48354;
  assign n58373 = ~n58371 & ~n58372;
  assign n58374 = pi432 & ~n48354;
  assign n58375 = pi1068 & n48354;
  assign n58376 = ~n58374 & ~n58375;
  assign n58377 = pi433 & ~n48354;
  assign n58378 = pi1042 & n48354;
  assign n58379 = ~n58377 & ~n58378;
  assign n58380 = pi434 & ~n48354;
  assign n58381 = pi1059 & n48354;
  assign n58382 = ~n58380 & ~n58381;
  assign n58383 = pi435 & ~n48354;
  assign n58384 = pi1053 & n48354;
  assign n58385 = ~n58383 & ~n58384;
  assign n58386 = pi436 & ~n48354;
  assign n58387 = pi1037 & n48354;
  assign n58388 = ~n58386 & ~n58387;
  assign n58389 = pi437 & ~n48354;
  assign n58390 = pi1070 & n48354;
  assign n58391 = ~n58389 & ~n58390;
  assign n58392 = pi438 & ~n48354;
  assign n58393 = pi1036 & n48354;
  assign n58394 = ~n58392 & ~n58393;
  assign n58395 = pi441 & ~n65040;
  assign n58396 = pi1044 & n65040;
  assign n58397 = ~n58395 & ~n58396;
  assign n58398 = pi443 & ~n48354;
  assign n58399 = pi1044 & n48354;
  assign n58400 = ~n58398 & ~n58399;
  assign n58401 = pi445 & ~n48354;
  assign n58402 = pi1081 & n48354;
  assign n58403 = ~n58401 & ~n58402;
  assign n58404 = pi450 & ~n65040;
  assign n58405 = pi1036 & n65040;
  assign n58406 = ~n58404 & ~n58405;
  assign n58407 = pi452 & ~n65040;
  assign n58408 = pi1053 & n65040;
  assign n58409 = ~n58407 & ~n58408;
  assign n58410 = pi455 & ~n65040;
  assign n58411 = pi1037 & n65040;
  assign n58412 = ~n58410 & ~n58411;
  assign n58413 = pi456 & ~n65041;
  assign n58414 = pi1044 & n65041;
  assign n58415 = ~n58413 & ~n58414;
  assign n58416 = pi463 & ~n65041;
  assign n58417 = pi1070 & n65041;
  assign n58418 = ~n58416 & ~n58417;
  assign n58419 = ~pi954 & ~n48508;
  assign n58420 = pi313 & pi954;
  assign po470 = ~n58419 & ~n58420;
  assign n58422 = pi228 & pi231;
  assign n58423 = ~pi228 & n48534;
  assign n58424 = ~n58422 & ~n58423;
  assign n58425 = ~pi100 & ~n58424;
  assign n58426 = ~n34060 & ~n58422;
  assign n58427 = pi100 & ~n58426;
  assign n58428 = ~pi87 & ~n58427;
  assign n58429 = ~n58425 & n58428;
  assign n58430 = pi87 & ~n58422;
  assign n58431 = ~n35420 & n58430;
  assign n58432 = ~pi75 & ~n58431;
  assign n58433 = ~n58429 & n58432;
  assign n58434 = ~n64304 & ~n58422;
  assign n58435 = pi75 & ~n58434;
  assign n58436 = ~pi92 & ~n58435;
  assign n58437 = ~n58433 & n58436;
  assign n58438 = pi92 & ~n58422;
  assign n58439 = ~n64341 & n58438;
  assign n58440 = ~n58437 & ~n58439;
  assign n58441 = ~pi54 & ~n58440;
  assign n58442 = pi54 & ~n58422;
  assign n58443 = ~pi74 & ~n58442;
  assign n58444 = ~n58441 & n58443;
  assign n58445 = ~n64306 & ~n58422;
  assign n58446 = ~n34066 & ~n58422;
  assign n58447 = pi74 & ~n58446;
  assign n58448 = ~n58434 & n58447;
  assign n58449 = pi74 & ~n58445;
  assign n58450 = ~pi55 & ~n65714;
  assign n58451 = ~n58444 & n58450;
  assign n58452 = pi55 & ~n58422;
  assign n58453 = ~pi56 & ~n58452;
  assign n58454 = ~n58451 & n58453;
  assign n58455 = ~n65025 & ~n58422;
  assign n58456 = pi56 & ~n58455;
  assign n58457 = ~pi62 & ~n58456;
  assign n58458 = ~n58454 & n58457;
  assign n58459 = pi62 & ~n58422;
  assign n58460 = ~n65024 & n58459;
  assign n58461 = ~n58458 & ~n58460;
  assign n58462 = n3472 & ~n58461;
  assign n58463 = ~n3472 & ~n58422;
  assign po383 = ~n58462 & ~n58463;
  assign n58465 = pi57 & ~pi59;
  assign n58466 = n40045 & n58465;
  assign n58467 = ~pi312 & n58466;
  assign n58468 = ~pi300 & pi301;
  assign n58469 = ~pi55 & n58468;
  assign n58470 = ~pi300 & n58467;
  assign n58471 = ~pi55 & pi301;
  assign n58472 = n58470 & n58471;
  assign n58473 = n58467 & n58469;
  assign n58474 = ~pi55 & ~pi311;
  assign n58475 = ~n65715 & ~n58474;
  assign n58476 = ~pi311 & n65715;
  assign n58477 = pi311 & ~n65715;
  assign n58478 = ~pi55 & ~n65715;
  assign n58479 = ~pi311 & ~n58478;
  assign n58480 = ~n58477 & ~n58479;
  assign n58481 = ~n58475 & ~n58476;
  assign n58482 = ~pi55 & ~n58470;
  assign n58483 = ~pi301 & n58482;
  assign n58484 = ~n65715 & ~n58483;
  assign n58485 = n6909 & n48675;
  assign n58486 = ~pi924 & n43669;
  assign n58487 = ~n43668 & ~n58486;
  assign n58488 = n58485 & ~n58487;
  assign n58489 = ~pi57 & ~n58488;
  assign n58490 = n3471 & n65065;
  assign n58491 = pi57 & ~n58490;
  assign n58492 = ~pi59 & ~n58491;
  assign n58493 = ~pi59 & ~n58489;
  assign n58494 = ~n58491 & n58493;
  assign n58495 = ~n58489 & n58492;
  assign n58496 = pi924 & n43669;
  assign n58497 = n58485 & n58496;
  assign n58498 = ~pi59 & ~n58497;
  assign n58499 = pi59 & ~n58490;
  assign n58500 = ~pi57 & ~n58499;
  assign n58501 = ~pi57 & ~n58498;
  assign n58502 = ~n58499 & n58501;
  assign n58503 = ~n58498 & n58500;
  assign n58504 = pi300 & ~n58467;
  assign n58505 = n58482 & ~n58504;
  assign n58506 = n62356 & n33908;
  assign n58507 = n2670 & n33909;
  assign n58508 = n62348 & n58506;
  assign n58509 = pi999 & n65719;
  assign n58510 = ~pi24 & n48637;
  assign n58511 = ~n58509 & ~n58510;
  assign po221 = n64866 & ~n58511;
  assign n58513 = pi312 & ~n58466;
  assign n58514 = ~n58467 & ~n58513;
  assign po469 = ~pi55 & ~n58514;
  assign n58516 = ~pi999 & n64866;
  assign po265 = n65719 & n58516;
  assign n58518 = pi481 & ~n47816;
  assign n58519 = pi248 & n47816;
  assign n58520 = ~n58518 & ~n58519;
  assign n58521 = pi482 & ~n47832;
  assign n58522 = pi249 & n47832;
  assign n58523 = ~n58521 & ~n58522;
  assign n58524 = pi483 & ~n47968;
  assign n58525 = pi242 & n47968;
  assign n58526 = ~n58524 & ~n58525;
  assign n58527 = pi484 & ~n47968;
  assign n58528 = pi249 & n47968;
  assign n58529 = ~n58527 & ~n58528;
  assign n58530 = pi485 & ~n47975;
  assign n58531 = pi234 & n47975;
  assign n58532 = ~n58530 & ~n58531;
  assign n58533 = pi486 & ~n47975;
  assign n58534 = pi244 & n47975;
  assign n58535 = ~n58533 & ~n58534;
  assign n58536 = pi487 & ~n47816;
  assign n58537 = pi246 & n47816;
  assign n58538 = ~n58536 & ~n58537;
  assign n58539 = pi488 & ~n47816;
  assign n58540 = ~pi239 & n47816;
  assign po645 = ~n58539 & ~n58540;
  assign n58542 = pi489 & ~n47975;
  assign n58543 = pi242 & n47975;
  assign n58544 = ~n58542 & ~n58543;
  assign n58545 = pi490 & ~n47968;
  assign n58546 = pi241 & n47968;
  assign n58547 = ~n58545 & ~n58546;
  assign n58548 = pi491 & ~n47968;
  assign n58549 = pi238 & n47968;
  assign n58550 = ~n58548 & ~n58549;
  assign n58551 = pi492 & ~n47968;
  assign n58552 = pi240 & n47968;
  assign n58553 = ~n58551 & ~n58552;
  assign n58554 = pi493 & ~n47968;
  assign n58555 = pi244 & n47968;
  assign n58556 = ~n58554 & ~n58555;
  assign n58557 = pi494 & ~n47968;
  assign n58558 = ~pi239 & n47968;
  assign po651 = ~n58557 & ~n58558;
  assign n58560 = pi495 & ~n47968;
  assign n58561 = pi235 & n47968;
  assign n58562 = ~n58560 & ~n58561;
  assign n58563 = pi496 & ~n47960;
  assign n58564 = pi249 & n47960;
  assign n58565 = ~n58563 & ~n58564;
  assign n58566 = pi497 & ~n47960;
  assign n58567 = ~pi239 & n47960;
  assign po654 = ~n58566 & ~n58567;
  assign n58569 = pi498 & ~n47832;
  assign n58570 = pi238 & n47832;
  assign n58571 = ~n58569 & ~n58570;
  assign n58572 = pi499 & ~n47960;
  assign n58573 = pi246 & n47960;
  assign n58574 = ~n58572 & ~n58573;
  assign n58575 = pi500 & ~n47960;
  assign n58576 = pi241 & n47960;
  assign n58577 = ~n58575 & ~n58576;
  assign n58578 = pi501 & ~n47960;
  assign n58579 = pi248 & n47960;
  assign n58580 = ~n58578 & ~n58579;
  assign n58581 = pi502 & ~n47960;
  assign n58582 = pi247 & n47960;
  assign n58583 = ~n58581 & ~n58582;
  assign n58584 = pi503 & ~n47960;
  assign n58585 = pi245 & n47960;
  assign n58586 = ~n58584 & ~n58585;
  assign n58587 = pi504 & ~n47953;
  assign n58588 = pi242 & n47953;
  assign n58589 = ~n58587 & ~n58588;
  assign n58590 = pi505 & ~n47960;
  assign n58591 = pi234 & n47952;
  assign n58592 = n47819 & n58591;
  assign n58593 = ~pi234 & n48906;
  assign n58594 = n47960 & n58593;
  assign n58595 = pi505 & ~n58594;
  assign n58596 = ~pi505 & n47819;
  assign n58597 = n58591 & n58596;
  assign n58598 = ~n58595 & ~n58597;
  assign n58599 = ~n58590 & ~n58592;
  assign n58600 = pi506 & ~n47953;
  assign n58601 = pi241 & n47953;
  assign n58602 = ~n58600 & ~n58601;
  assign n58603 = pi507 & ~n47953;
  assign n58604 = pi238 & n47953;
  assign n58605 = ~n58603 & ~n58604;
  assign n58606 = pi508 & ~n47953;
  assign n58607 = pi247 & n47953;
  assign n58608 = ~n58606 & ~n58607;
  assign n58609 = pi509 & ~n47953;
  assign n58610 = pi245 & n47953;
  assign n58611 = ~n58609 & ~n58610;
  assign n58612 = pi510 & ~n47816;
  assign n58613 = pi242 & n47816;
  assign n58614 = ~n58612 & ~n58613;
  assign n58615 = ~pi234 & n48903;
  assign n58616 = n47816 & ~n58615;
  assign n58617 = pi511 & ~n47816;
  assign n58618 = ~n58616 & ~n58617;
  assign n58619 = pi512 & ~n47816;
  assign n58620 = pi235 & n47816;
  assign n58621 = ~n58619 & ~n58620;
  assign n58622 = pi513 & ~n47816;
  assign n58623 = pi244 & n47816;
  assign n58624 = ~n58622 & ~n58623;
  assign n58625 = pi514 & ~n47816;
  assign n58626 = pi245 & n47816;
  assign n58627 = ~n58625 & ~n58626;
  assign n58628 = pi515 & ~n47816;
  assign n58629 = pi240 & n47816;
  assign n58630 = ~n58628 & ~n58629;
  assign n58631 = pi516 & ~n47816;
  assign n58632 = pi247 & n47816;
  assign n58633 = ~n58631 & ~n58632;
  assign n58634 = pi517 & ~n47816;
  assign n58635 = pi238 & n47816;
  assign n58636 = ~n58634 & ~n58635;
  assign n58637 = pi518 & ~n47824;
  assign n58638 = pi234 & n65015;
  assign n58639 = n47819 & n58638;
  assign n58640 = n47824 & n58615;
  assign n58641 = pi518 & ~n58640;
  assign n58642 = ~pi518 & n47819;
  assign n58643 = n58638 & n58642;
  assign n58644 = ~n58641 & ~n58643;
  assign n58645 = ~n58637 & ~n58639;
  assign n58646 = pi519 & ~n47824;
  assign n58647 = ~pi239 & n47824;
  assign po676 = ~n58646 & ~n58647;
  assign n58649 = pi520 & ~n47824;
  assign n58650 = pi246 & n47824;
  assign n58651 = ~n58649 & ~n58650;
  assign n58652 = pi521 & ~n47824;
  assign n58653 = pi248 & n47824;
  assign n58654 = ~n58652 & ~n58653;
  assign n58655 = pi522 & ~n47824;
  assign n58656 = pi238 & n47824;
  assign n58657 = ~n58655 & ~n58656;
  assign n58658 = pi523 & ~n47982;
  assign n58659 = n47963 & n58638;
  assign n58660 = n47982 & n58615;
  assign n58661 = pi523 & ~n58660;
  assign n58662 = ~pi523 & n47963;
  assign n58663 = n58638 & n58662;
  assign n58664 = ~n58661 & ~n58663;
  assign n58665 = ~n58658 & ~n58659;
  assign n58666 = pi524 & ~n47982;
  assign n58667 = ~pi239 & n47982;
  assign po681 = ~n58666 & ~n58667;
  assign n58669 = pi525 & ~n47982;
  assign n58670 = pi245 & n47982;
  assign n58671 = ~n58669 & ~n58670;
  assign n58672 = pi526 & ~n47982;
  assign n58673 = pi246 & n47982;
  assign n58674 = ~n58672 & ~n58673;
  assign n58675 = pi527 & ~n47982;
  assign n58676 = pi247 & n47982;
  assign n58677 = ~n58675 & ~n58676;
  assign n58678 = pi528 & ~n47982;
  assign n58679 = pi249 & n47982;
  assign n58680 = ~n58678 & ~n58679;
  assign n58681 = pi529 & ~n47982;
  assign n58682 = pi238 & n47982;
  assign n58683 = ~n58681 & ~n58682;
  assign n58684 = pi530 & ~n47982;
  assign n58685 = pi240 & n47982;
  assign n58686 = ~n58684 & ~n58685;
  assign n58687 = pi531 & ~n47832;
  assign n58688 = pi235 & n47832;
  assign n58689 = ~n58687 & ~n58688;
  assign n58690 = pi532 & ~n47832;
  assign n58691 = pi247 & n47832;
  assign n58692 = ~n58690 & ~n58691;
  assign n58693 = pi533 & ~n47953;
  assign n58694 = pi235 & n47953;
  assign n58695 = ~n58693 & ~n58694;
  assign n58696 = ~pi228 & ~pi1093;
  assign n58697 = pi123 & pi228;
  assign n58698 = ~pi123 & pi228;
  assign n58699 = ~pi228 & pi1093;
  assign n58700 = ~n58698 & ~n58699;
  assign n58701 = ~n58696 & ~n58697;
  assign n58702 = pi199 & ~n65723;
  assign n58703 = ~pi262 & ~pi1093;
  assign n58704 = ~n49005 & ~n58703;
  assign n58705 = ~pi228 & ~n58704;
  assign n58706 = pi123 & pi262;
  assign n58707 = ~pi123 & ~pi1142;
  assign n58708 = pi228 & ~n58707;
  assign n58709 = pi228 & ~n58706;
  assign n58710 = ~n58707 & n58709;
  assign n58711 = ~n58706 & n58708;
  assign n58712 = ~n58705 & ~n65724;
  assign n58713 = n54329 & ~n65723;
  assign n58714 = ~n58712 & ~n58713;
  assign n58715 = pi208 & ~n58714;
  assign n58716 = ~n58702 & ~n58715;
  assign n58717 = ~pi299 & ~n58716;
  assign n58718 = ~n52555 & ~n65529;
  assign n58719 = n58712 & ~n58718;
  assign n58720 = ~pi262 & n65723;
  assign n58721 = ~n54354 & ~n58720;
  assign n58722 = ~n65529 & n58721;
  assign n58723 = n62455 & ~n58722;
  assign n58724 = ~n58719 & n58723;
  assign n58725 = ~n65529 & ~n58720;
  assign n58726 = n52548 & ~n58702;
  assign n58727 = n58725 & ~n58726;
  assign n58728 = ~n58712 & ~n58727;
  assign n58729 = ~pi207 & n58720;
  assign n58730 = ~pi208 & ~n58729;
  assign n58731 = ~n65529 & ~n58730;
  assign n58732 = ~n58728 & ~n58731;
  assign n58733 = pi299 & ~n58725;
  assign n58734 = ~n54330 & ~n65723;
  assign n58735 = ~pi299 & ~n58734;
  assign n58736 = ~n58712 & n58735;
  assign n58737 = pi208 & ~n58736;
  assign n58738 = ~n58733 & n58737;
  assign n58739 = n62455 & ~n58738;
  assign n58740 = ~n58732 & n58739;
  assign n58741 = ~n58717 & n58724;
  assign n58742 = ~n65430 & ~n65723;
  assign n58743 = ~n62455 & ~n58712;
  assign n58744 = ~n58742 & n58743;
  assign n58745 = ~n65725 & ~n58744;
  assign n58746 = ~pi284 & n65723;
  assign n58747 = pi1143 & ~n65723;
  assign n58748 = ~n55137 & n58747;
  assign n58749 = ~n58746 & ~n58748;
  assign n58750 = pi266 & pi992;
  assign n58751 = ~pi280 & n58750;
  assign n58752 = ~pi269 & n58751;
  assign n58753 = ~pi281 & n58752;
  assign n58754 = n48941 & n58753;
  assign n58755 = ~pi264 & n58754;
  assign n58756 = ~pi265 & n58755;
  assign po959 = ~pi274 & n58756;
  assign n58758 = pi274 & ~n58756;
  assign po816 = ~po959 & ~n58758;
  assign n58760 = pi265 & ~n58755;
  assign po976 = ~n58756 & ~n58760;
  assign n58762 = ~pi282 & n58753;
  assign n58763 = ~pi270 & n58762;
  assign n58764 = pi277 & ~n58763;
  assign po977 = ~n58754 & ~n58764;
  assign n58766 = pi270 & ~n58762;
  assign po962 = ~n58763 & ~n58766;
  assign n58768 = pi282 & ~n58753;
  assign po992 = ~n58762 & ~n58768;
  assign n58770 = pi269 & ~n58751;
  assign po974 = ~n58752 & ~n58770;
  assign n58772 = pi280 & ~n58750;
  assign po1070 = ~n58751 & ~n58772;
  assign n58774 = pi311 & ~pi312;
  assign po1080 = n58468 & n58774;
  assign n58776 = ~pi266 & ~pi992;
  assign po1104 = ~n58750 & ~n58776;
  assign n58778 = ~pi313 & ~pi954;
  assign n58779 = pi949 & pi954;
  assign n58780 = ~pi949 & pi954;
  assign n58781 = pi313 & ~pi954;
  assign n58782 = ~n58780 & ~n58781;
  assign n58783 = ~n58778 & ~n58779;
  assign n58784 = n41471 & n65014;
  assign n58785 = n62455 & n47144;
  assign n58786 = ~pi222 & ~pi223;
  assign n58787 = pi937 & ~n58786;
  assign n58788 = pi273 & n28811;
  assign n58789 = ~n58787 & ~n58788;
  assign n58790 = n65727 & n58789;
  assign n58791 = n38199 & ~n65014;
  assign n58792 = ~n58790 & ~n58791;
  assign n58793 = pi237 & ~n58792;
  assign n58794 = n47158 & ~n65014;
  assign n58795 = ~n65727 & ~n58794;
  assign n58796 = ~pi1148 & n58795;
  assign n58797 = ~n7034 & n58790;
  assign n58798 = ~pi215 & n39839;
  assign n58799 = ~pi273 & n58798;
  assign n58800 = pi833 & n3056;
  assign n58801 = ~pi937 & n58800;
  assign n58802 = ~n58799 & ~n58801;
  assign n58803 = ~n65014 & ~n58802;
  assign n58804 = ~n58797 & ~n58803;
  assign n58805 = ~n58796 & n58804;
  assign n58806 = ~n58793 & n58804;
  assign n58807 = ~n58796 & n58806;
  assign n58808 = ~n58793 & n58805;
  assign n58809 = pi1147 & n58795;
  assign n58810 = ~n7118 & n58794;
  assign n58811 = pi934 & ~n41037;
  assign n58812 = pi271 & n39839;
  assign n58813 = ~n58811 & ~n58812;
  assign n58814 = n58810 & ~n58813;
  assign n58815 = pi222 & ~pi934;
  assign n58816 = ~pi271 & n28811;
  assign n58817 = ~n58815 & ~n58816;
  assign n58818 = n65727 & n58817;
  assign n58819 = ~n58791 & ~n58818;
  assign n58820 = ~n58814 & n58819;
  assign n58821 = ~n58809 & n58820;
  assign n58822 = ~pi233 & ~n58821;
  assign n58823 = n58794 & n58813;
  assign n58824 = n65727 & ~n58817;
  assign n58825 = n38189 & n65014;
  assign n58826 = n62455 & n38188;
  assign n58827 = pi1147 & ~n65729;
  assign n58828 = pi1147 & ~n58824;
  assign n58829 = ~n65729 & n58828;
  assign n58830 = ~n58824 & n58827;
  assign n58831 = ~n58823 & n65730;
  assign n58832 = ~n7034 & n65727;
  assign n58833 = ~n58810 & ~n58832;
  assign n58834 = ~pi1147 & ~n58833;
  assign n58835 = ~n58820 & n58834;
  assign n58836 = ~n58831 & ~n58835;
  assign n58837 = pi233 & ~n58836;
  assign n58838 = ~n58822 & ~n58837;
  assign n58839 = pi1157 & ~n47158;
  assign n58840 = pi926 & n58800;
  assign n58841 = ~pi243 & n58798;
  assign n58842 = ~n58840 & ~n58841;
  assign n58843 = ~n58839 & n58842;
  assign n58844 = ~n62455 & ~n58843;
  assign n58845 = ~n39840 & ~n39842;
  assign n58846 = ~pi243 & ~n58845;
  assign n58847 = ~n47137 & ~n47144;
  assign n58848 = ~pi1157 & n58847;
  assign n58849 = ~pi926 & ~n58847;
  assign n58850 = ~pi243 & pi1157;
  assign n58851 = pi299 & n41037;
  assign n58852 = ~pi299 & n58786;
  assign n58853 = ~pi222 & n2979;
  assign n58854 = ~n64521 & ~n65731;
  assign n58855 = ~n58850 & ~n58854;
  assign n58856 = ~n58849 & ~n58855;
  assign n58857 = ~n58848 & n58854;
  assign n58858 = ~n58850 & ~n58857;
  assign n58859 = ~n58849 & ~n58858;
  assign n58860 = ~n58848 & n58856;
  assign n58861 = ~n58846 & ~n65732;
  assign n58862 = pi299 & n38199;
  assign n58863 = ~n38188 & ~n64522;
  assign n58864 = pi926 & n58850;
  assign n58865 = ~n58863 & n58864;
  assign n58866 = n62455 & ~n58865;
  assign n58867 = ~n58861 & n58866;
  assign n58868 = pi926 & ~n58847;
  assign n58869 = pi1157 & n58847;
  assign n58870 = ~n58846 & ~n58869;
  assign n58871 = ~n58846 & ~n58868;
  assign n58872 = ~n58869 & n58871;
  assign n58873 = ~n58868 & n58870;
  assign n58874 = ~n58846 & n58855;
  assign n58875 = ~n58865 & ~n58874;
  assign n58876 = ~n65733 & n58875;
  assign n58877 = n62455 & ~n58876;
  assign n58878 = ~n62455 & ~n58841;
  assign n58879 = ~n58839 & ~n58840;
  assign n58880 = n58878 & n58879;
  assign n58881 = ~n58877 & ~n58880;
  assign n58882 = ~n58844 & ~n58867;
  assign n58883 = ~n62455 & ~n58798;
  assign n58884 = n62455 & n58845;
  assign n58885 = n62455 & ~n58845;
  assign n58886 = ~n62455 & n58798;
  assign n58887 = ~n58885 & ~n58886;
  assign n58888 = ~n58883 & ~n58884;
  assign n58889 = ~pi943 & n65735;
  assign n58890 = pi943 & n58833;
  assign n58891 = ~n58889 & ~n58890;
  assign n58892 = ~pi1151 & ~n58891;
  assign n58893 = ~n58791 & ~n65729;
  assign n58894 = pi943 & pi1151;
  assign n58895 = ~n58893 & n58894;
  assign n58896 = ~n58795 & n58889;
  assign n58897 = n62455 & ~n58854;
  assign n58898 = ~n62455 & n41037;
  assign n58899 = ~n62455 & ~n41037;
  assign n58900 = n62455 & n58854;
  assign n58901 = ~n58899 & ~n58900;
  assign n58902 = ~n58897 & ~n58898;
  assign n58903 = ~pi275 & n65736;
  assign n58904 = ~n58896 & ~n58903;
  assign n58905 = ~n58895 & ~n58903;
  assign n58906 = ~n58896 & n58905;
  assign n58907 = ~n58895 & n58904;
  assign po623 = ~n58892 & n65737;
  assign n58909 = pi1156 & ~n47158;
  assign n58910 = pi942 & n58800;
  assign n58911 = ~pi263 & n58798;
  assign n58912 = ~n58910 & ~n58911;
  assign n58913 = ~n58909 & n58912;
  assign n58914 = ~n62455 & ~n58913;
  assign n58915 = ~pi263 & ~n58845;
  assign n58916 = ~pi1156 & n58847;
  assign n58917 = ~pi942 & ~n58847;
  assign n58918 = ~pi263 & pi1156;
  assign n58919 = ~n58854 & ~n58918;
  assign n58920 = ~n58917 & ~n58919;
  assign n58921 = n58854 & ~n58916;
  assign n58922 = ~n58918 & ~n58921;
  assign n58923 = ~n58917 & ~n58922;
  assign n58924 = ~n58916 & n58920;
  assign n58925 = ~n58915 & ~n65738;
  assign n58926 = pi942 & n58918;
  assign n58927 = ~n58863 & n58926;
  assign n58928 = n62455 & ~n58927;
  assign n58929 = ~n58925 & n58928;
  assign n58930 = pi942 & ~n58847;
  assign n58931 = pi1156 & n58847;
  assign n58932 = ~n58915 & ~n58931;
  assign n58933 = ~n58915 & ~n58930;
  assign n58934 = ~n58931 & n58933;
  assign n58935 = ~n58930 & n58932;
  assign n58936 = ~n58915 & n58919;
  assign n58937 = ~n58927 & ~n58936;
  assign n58938 = ~n65739 & n58937;
  assign n58939 = n62455 & ~n58938;
  assign n58940 = ~n62455 & ~n58911;
  assign n58941 = ~n58909 & ~n58910;
  assign n58942 = n58940 & n58941;
  assign n58943 = ~n58939 & ~n58942;
  assign n58944 = ~n58914 & ~n58929;
  assign n58945 = pi1155 & ~n47158;
  assign n58946 = pi925 & n58800;
  assign n58947 = pi267 & n58798;
  assign n58948 = ~n58946 & ~n58947;
  assign n58949 = ~n58945 & n58948;
  assign n58950 = ~n62455 & ~n58949;
  assign n58951 = pi267 & ~n58845;
  assign n58952 = ~pi1155 & n58847;
  assign n58953 = ~pi925 & ~n58847;
  assign n58954 = pi267 & pi1155;
  assign n58955 = ~n58854 & ~n58954;
  assign n58956 = ~n58953 & ~n58955;
  assign n58957 = n58854 & ~n58952;
  assign n58958 = ~n58954 & ~n58957;
  assign n58959 = ~n58953 & ~n58958;
  assign n58960 = ~n58952 & n58956;
  assign n58961 = ~n58951 & ~n65741;
  assign n58962 = pi925 & n58954;
  assign n58963 = ~n58863 & n58962;
  assign n58964 = n62455 & ~n58963;
  assign n58965 = ~n58961 & n58964;
  assign n58966 = pi925 & ~n58847;
  assign n58967 = pi1155 & n58847;
  assign n58968 = ~n58951 & ~n58967;
  assign n58969 = ~n58951 & ~n58966;
  assign n58970 = ~n58967 & n58969;
  assign n58971 = ~n58966 & n58968;
  assign n58972 = ~n58951 & n58955;
  assign n58973 = ~n58963 & ~n58972;
  assign n58974 = ~n65742 & n58973;
  assign n58975 = n62455 & ~n58974;
  assign n58976 = ~n62455 & ~n58947;
  assign n58977 = ~n58945 & ~n58946;
  assign n58978 = n58976 & n58977;
  assign n58979 = ~n58975 & ~n58978;
  assign n58980 = ~n58950 & ~n58965;
  assign n58981 = pi1153 & ~n47158;
  assign n58982 = pi941 & n58800;
  assign n58983 = pi253 & n58798;
  assign n58984 = ~n58982 & ~n58983;
  assign n58985 = ~n58981 & n58984;
  assign n58986 = ~n62455 & ~n58985;
  assign n58987 = pi253 & ~n58845;
  assign n58988 = ~pi1153 & n58847;
  assign n58989 = ~pi941 & ~n58847;
  assign n58990 = pi253 & pi1153;
  assign n58991 = ~n58854 & ~n58990;
  assign n58992 = ~n58989 & ~n58991;
  assign n58993 = n58854 & ~n58988;
  assign n58994 = ~n58990 & ~n58993;
  assign n58995 = ~n58989 & ~n58994;
  assign n58996 = ~n58988 & n58992;
  assign n58997 = ~n58987 & ~n65744;
  assign n58998 = pi941 & n58990;
  assign n58999 = ~n58863 & n58998;
  assign n59000 = n62455 & ~n58999;
  assign n59001 = ~n58997 & n59000;
  assign n59002 = pi941 & ~n58847;
  assign n59003 = pi1153 & n58847;
  assign n59004 = ~n58987 & ~n59003;
  assign n59005 = ~n58987 & ~n59002;
  assign n59006 = ~n59003 & n59005;
  assign n59007 = ~n59002 & n59004;
  assign n59008 = ~n58987 & n58991;
  assign n59009 = ~n58999 & ~n59008;
  assign n59010 = ~n65745 & n59009;
  assign n59011 = n62455 & ~n59010;
  assign n59012 = ~n62455 & ~n58983;
  assign n59013 = ~n58981 & ~n58982;
  assign n59014 = n59012 & n59013;
  assign n59015 = ~n59011 & ~n59014;
  assign n59016 = ~n58986 & ~n59001;
  assign n59017 = pi1154 & ~n47158;
  assign n59018 = pi923 & n58800;
  assign n59019 = pi254 & n58798;
  assign n59020 = ~n59018 & ~n59019;
  assign n59021 = ~n59017 & n59020;
  assign n59022 = ~n62455 & ~n59021;
  assign n59023 = pi254 & ~n58845;
  assign n59024 = ~pi1154 & n58847;
  assign n59025 = ~pi923 & ~n58847;
  assign n59026 = pi254 & pi1154;
  assign n59027 = ~n58854 & ~n59026;
  assign n59028 = ~n59025 & ~n59027;
  assign n59029 = n58854 & ~n59024;
  assign n59030 = ~n59026 & ~n59029;
  assign n59031 = ~n59025 & ~n59030;
  assign n59032 = ~n59024 & n59028;
  assign n59033 = ~n59023 & ~n65747;
  assign n59034 = pi923 & n59026;
  assign n59035 = ~n58863 & n59034;
  assign n59036 = n62455 & ~n59035;
  assign n59037 = ~n59033 & n59036;
  assign n59038 = pi923 & ~n58847;
  assign n59039 = pi1154 & n58847;
  assign n59040 = ~n59023 & ~n59039;
  assign n59041 = ~n59023 & ~n59038;
  assign n59042 = ~n59039 & n59041;
  assign n59043 = ~n59038 & n59040;
  assign n59044 = ~n59023 & n59027;
  assign n59045 = ~n59035 & ~n59044;
  assign n59046 = ~n65748 & n59045;
  assign n59047 = n62455 & ~n59046;
  assign n59048 = ~n62455 & ~n59019;
  assign n59049 = ~n59017 & ~n59018;
  assign n59050 = n59048 & n59049;
  assign n59051 = ~n59047 & ~n59050;
  assign n59052 = ~n59022 & ~n59037;
  assign n59053 = ~pi922 & n65735;
  assign n59054 = pi922 & n58833;
  assign n59055 = ~n59053 & ~n59054;
  assign n59056 = ~pi1152 & ~n59055;
  assign n59057 = pi922 & pi1152;
  assign n59058 = ~n58893 & n59057;
  assign n59059 = ~n58795 & n59053;
  assign n59060 = ~pi268 & n65736;
  assign n59061 = ~n59059 & ~n59060;
  assign n59062 = ~n59058 & ~n59060;
  assign n59063 = ~n59059 & n59062;
  assign n59064 = ~n59058 & n59061;
  assign po630 = ~n59056 & n65750;
  assign n59066 = ~pi931 & n65735;
  assign n59067 = pi931 & n58833;
  assign n59068 = ~n59066 & ~n59067;
  assign n59069 = ~pi1150 & ~n59068;
  assign n59070 = pi931 & pi1150;
  assign n59071 = ~n58893 & n59070;
  assign n59072 = ~n58795 & n59066;
  assign n59073 = ~pi272 & n65736;
  assign n59074 = ~n59072 & ~n59073;
  assign n59075 = ~n59071 & ~n59073;
  assign n59076 = ~n59072 & n59075;
  assign n59077 = ~n59071 & n59074;
  assign po631 = ~n59069 & n65751;
  assign n59079 = ~pi936 & n65735;
  assign n59080 = pi936 & n58833;
  assign n59081 = ~n59079 & ~n59080;
  assign n59082 = ~pi1149 & ~n59081;
  assign n59083 = pi936 & pi1149;
  assign n59084 = ~n58893 & n59083;
  assign n59085 = ~n58795 & n59079;
  assign n59086 = ~pi283 & n65736;
  assign n59087 = ~n59085 & ~n59086;
  assign n59088 = ~n59084 & ~n59086;
  assign n59089 = ~n59085 & n59088;
  assign n59090 = ~n59084 & n59087;
  assign po632 = ~n59082 & n65752;
  assign n59092 = ~pi241 & ~pi506;
  assign n59093 = pi241 & pi506;
  assign n59094 = ~n59092 & ~n59093;
  assign n59095 = ~pi557 & ~n58593;
  assign n59096 = pi234 & n48906;
  assign n59097 = pi557 & ~n59096;
  assign n59098 = ~pi246 & ~pi536;
  assign n59099 = pi246 & pi536;
  assign n59100 = ~n59098 & ~n59099;
  assign n59101 = pi248 & ~pi537;
  assign n59102 = ~pi248 & pi537;
  assign n59103 = ~n59101 & ~n59102;
  assign n59104 = pi249 & ~pi538;
  assign n59105 = ~pi249 & pi538;
  assign n59106 = ~pi249 & ~pi538;
  assign n59107 = pi249 & pi538;
  assign n59108 = ~n59106 & ~n59107;
  assign n59109 = ~n59104 & ~n59105;
  assign n59110 = n59103 & ~n65753;
  assign n59111 = ~n59100 & n59110;
  assign n59112 = ~n59097 & n59111;
  assign n59113 = ~n59097 & ~n59100;
  assign n59114 = ~n59095 & ~n59100;
  assign n59115 = ~n59097 & n59114;
  assign n59116 = ~n59095 & n59113;
  assign n59117 = ~pi538 & n65754;
  assign n59118 = ~pi249 & ~n59117;
  assign n59119 = pi538 & n65754;
  assign n59120 = pi249 & ~n59119;
  assign n59121 = ~n59118 & ~n59120;
  assign n59122 = ~n65753 & n65754;
  assign n59123 = ~pi537 & n65755;
  assign n59124 = ~pi248 & ~n59123;
  assign n59125 = pi537 & n65755;
  assign n59126 = pi248 & ~n59125;
  assign n59127 = ~n59124 & ~n59126;
  assign n59128 = ~n59095 & n59112;
  assign n59129 = ~n59094 & n65756;
  assign n59130 = ~pi240 & ~pi535;
  assign n59131 = pi240 & pi535;
  assign n59132 = ~n59130 & ~n59131;
  assign n59133 = n59129 & ~n59132;
  assign n59134 = pi534 & n59133;
  assign n59135 = ~pi239 & ~n59134;
  assign n59136 = ~pi534 & n59133;
  assign n59137 = pi239 & ~n59136;
  assign n59138 = ~n59135 & ~n59137;
  assign n59139 = pi504 & n59138;
  assign n59140 = pi242 & ~n59139;
  assign n59141 = ~pi504 & n59138;
  assign n59142 = ~pi242 & ~n59141;
  assign n59143 = ~n59140 & ~n59142;
  assign n59144 = pi533 & n59143;
  assign n59145 = pi235 & ~n59144;
  assign n59146 = ~pi533 & n59143;
  assign n59147 = ~pi235 & ~n59146;
  assign n59148 = ~n59145 & ~n59147;
  assign n59149 = pi558 & n59148;
  assign n59150 = pi244 & ~n59149;
  assign n59151 = ~pi558 & n59148;
  assign n59152 = ~pi244 & ~n59151;
  assign n59153 = ~n59150 & ~n59152;
  assign n59154 = pi509 & n59153;
  assign n59155 = pi245 & ~n59154;
  assign n59156 = ~pi509 & n59153;
  assign n59157 = ~pi245 & ~n59156;
  assign n59158 = ~n59155 & ~n59157;
  assign n59159 = pi508 & n59158;
  assign n59160 = pi247 & ~n59159;
  assign n59161 = ~pi511 & ~n58615;
  assign n59162 = pi234 & n48903;
  assign n59163 = pi511 & ~n59162;
  assign n59164 = ~pi248 & ~pi481;
  assign n59165 = pi248 & pi481;
  assign n59166 = ~n59164 & ~n59165;
  assign n59167 = pi246 & ~pi487;
  assign n59168 = ~pi246 & pi487;
  assign n59169 = pi246 & pi487;
  assign n59170 = ~pi246 & ~pi487;
  assign n59171 = ~n59169 & ~n59170;
  assign n59172 = ~n59167 & ~n59168;
  assign n59173 = pi249 & ~pi579;
  assign n59174 = ~pi249 & pi579;
  assign n59175 = ~pi249 & ~pi579;
  assign n59176 = pi249 & pi579;
  assign n59177 = ~n59175 & ~n59176;
  assign n59178 = ~n59173 & ~n59174;
  assign n59179 = ~n65757 & ~n65758;
  assign n59180 = ~n59166 & n59179;
  assign n59181 = ~n59163 & n59180;
  assign n59182 = ~n59163 & ~n65757;
  assign n59183 = ~n59161 & ~n65757;
  assign n59184 = ~n59163 & n59183;
  assign n59185 = ~n59161 & n59182;
  assign n59186 = ~n65758 & n65759;
  assign n59187 = ~n59166 & n59186;
  assign n59188 = ~n59161 & n59181;
  assign n59189 = pi559 & n65760;
  assign n59190 = pi241 & ~n59189;
  assign n59191 = ~pi559 & n65760;
  assign n59192 = ~pi241 & ~n59191;
  assign n59193 = ~n59190 & ~n59192;
  assign n59194 = pi515 & n59193;
  assign n59195 = pi240 & ~n59194;
  assign n59196 = ~pi506 & n65756;
  assign n59197 = n59192 & ~n59196;
  assign n59198 = pi506 & n65756;
  assign n59199 = n59190 & ~n59198;
  assign n59200 = n59106 & n65754;
  assign n59201 = n65758 & ~n59200;
  assign n59202 = ~pi579 & ~n59186;
  assign n59203 = ~n59118 & n65759;
  assign n59204 = pi579 & ~n59203;
  assign n59205 = ~n59202 & ~n59204;
  assign n59206 = n65759 & ~n59201;
  assign n59207 = ~n65755 & ~n65761;
  assign n59208 = ~pi537 & ~n59207;
  assign n59209 = pi537 & n59186;
  assign n59210 = ~pi248 & ~n59209;
  assign n59211 = ~n59208 & n59210;
  assign n59212 = ~n59126 & ~n59211;
  assign n59213 = ~pi481 & ~n59212;
  assign n59214 = pi537 & ~n59207;
  assign n59215 = ~pi537 & n59186;
  assign n59216 = pi248 & ~n59215;
  assign n59217 = ~n59214 & n59216;
  assign n59218 = ~n59124 & ~n59217;
  assign n59219 = pi481 & ~n59218;
  assign n59220 = ~n59213 & ~n59219;
  assign n59221 = ~pi559 & n59220;
  assign n59222 = pi559 & n65756;
  assign n59223 = ~pi241 & ~n59222;
  assign n59224 = ~n59221 & n59223;
  assign n59225 = ~n59190 & ~n59224;
  assign n59226 = ~pi506 & ~n59225;
  assign n59227 = pi559 & n59220;
  assign n59228 = ~pi559 & n65756;
  assign n59229 = pi241 & ~n59228;
  assign n59230 = ~n59227 & n59229;
  assign n59231 = ~n59192 & ~n59230;
  assign n59232 = pi506 & ~n59231;
  assign n59233 = ~n59226 & ~n59232;
  assign n59234 = ~n59197 & ~n59199;
  assign n59235 = ~pi515 & n65762;
  assign n59236 = pi515 & n59129;
  assign n59237 = ~pi240 & ~n59236;
  assign n59238 = ~n59235 & n59237;
  assign n59239 = ~n59195 & ~n59238;
  assign n59240 = ~pi535 & ~n59239;
  assign n59241 = ~pi515 & n59193;
  assign n59242 = ~pi240 & ~n59241;
  assign n59243 = pi515 & n65762;
  assign n59244 = ~pi515 & n59129;
  assign n59245 = pi240 & ~n59244;
  assign n59246 = ~n59243 & n59245;
  assign n59247 = ~n59242 & ~n59246;
  assign n59248 = pi535 & ~n59247;
  assign n59249 = ~n59240 & ~n59248;
  assign n59250 = ~pi534 & n59249;
  assign n59251 = ~n59195 & ~n59242;
  assign n59252 = pi534 & n59251;
  assign n59253 = pi239 & ~n59252;
  assign n59254 = ~n59250 & n59253;
  assign n59255 = ~n59135 & ~n59254;
  assign n59256 = ~pi488 & ~n59255;
  assign n59257 = pi534 & n59249;
  assign n59258 = ~pi534 & n59251;
  assign n59259 = ~pi239 & ~n59258;
  assign n59260 = ~n59257 & n59259;
  assign n59261 = ~n59137 & ~n59260;
  assign n59262 = pi488 & ~n59261;
  assign n59263 = ~n59256 & ~n59262;
  assign n59264 = ~pi504 & n59263;
  assign n59265 = pi239 & ~pi488;
  assign n59266 = ~pi239 & pi488;
  assign n59267 = ~n59265 & ~n59266;
  assign n59268 = n59251 & ~n59267;
  assign n59269 = pi504 & n59268;
  assign n59270 = ~pi242 & ~n59269;
  assign n59271 = ~n59264 & n59270;
  assign n59272 = ~n59140 & ~n59271;
  assign n59273 = ~pi510 & ~n59272;
  assign n59274 = pi504 & n59263;
  assign n59275 = ~pi504 & n59268;
  assign n59276 = pi242 & ~n59275;
  assign n59277 = ~n59274 & n59276;
  assign n59278 = ~n59142 & ~n59277;
  assign n59279 = pi510 & ~n59278;
  assign n59280 = ~n59273 & ~n59279;
  assign n59281 = ~pi533 & n59280;
  assign n59282 = ~pi242 & ~pi510;
  assign n59283 = pi242 & pi510;
  assign n59284 = ~n59282 & ~n59283;
  assign n59285 = n59268 & ~n59284;
  assign n59286 = pi533 & n59285;
  assign n59287 = ~pi235 & ~n59286;
  assign n59288 = ~n59281 & n59287;
  assign n59289 = ~n59145 & ~n59288;
  assign n59290 = ~pi512 & ~n59289;
  assign n59291 = pi533 & n59280;
  assign n59292 = ~pi533 & n59285;
  assign n59293 = pi235 & ~n59292;
  assign n59294 = ~n59291 & n59293;
  assign n59295 = ~n59147 & ~n59294;
  assign n59296 = pi512 & ~n59295;
  assign n59297 = ~n59290 & ~n59296;
  assign n59298 = ~pi558 & n59297;
  assign n59299 = ~pi235 & ~pi512;
  assign n59300 = pi235 & pi512;
  assign n59301 = ~n59299 & ~n59300;
  assign n59302 = n59285 & ~n59301;
  assign n59303 = pi558 & n59302;
  assign n59304 = ~pi244 & ~n59303;
  assign n59305 = ~n59298 & n59304;
  assign n59306 = ~n59150 & ~n59305;
  assign n59307 = ~pi513 & ~n59306;
  assign n59308 = pi558 & n59297;
  assign n59309 = ~pi558 & n59302;
  assign n59310 = pi244 & ~n59309;
  assign n59311 = ~n59308 & n59310;
  assign n59312 = ~n59152 & ~n59311;
  assign n59313 = pi513 & ~n59312;
  assign n59314 = ~n59307 & ~n59313;
  assign n59315 = ~pi509 & n59314;
  assign n59316 = ~pi244 & ~pi513;
  assign n59317 = pi244 & pi513;
  assign n59318 = ~n59316 & ~n59317;
  assign n59319 = n59302 & ~n59318;
  assign n59320 = pi509 & n59319;
  assign n59321 = ~pi245 & ~n59320;
  assign n59322 = ~n59315 & n59321;
  assign n59323 = ~n59155 & ~n59322;
  assign n59324 = ~pi514 & ~n59323;
  assign n59325 = pi509 & n59314;
  assign n59326 = ~pi509 & n59319;
  assign n59327 = pi245 & ~n59326;
  assign n59328 = ~n59325 & n59327;
  assign n59329 = ~n59157 & ~n59328;
  assign n59330 = pi514 & ~n59329;
  assign n59331 = ~n59324 & ~n59330;
  assign n59332 = ~pi508 & n59331;
  assign n59333 = ~pi245 & ~pi514;
  assign n59334 = pi245 & pi514;
  assign n59335 = ~n59333 & ~n59334;
  assign n59336 = n59319 & ~n59335;
  assign n59337 = pi508 & n59336;
  assign n59338 = ~pi247 & ~n59337;
  assign n59339 = ~n59332 & n59338;
  assign n59340 = ~n59160 & ~n59339;
  assign n59341 = ~pi516 & ~n59340;
  assign n59342 = ~pi508 & n59158;
  assign n59343 = ~pi247 & ~n59342;
  assign n59344 = pi508 & n59331;
  assign n59345 = ~pi508 & n59336;
  assign n59346 = pi247 & ~n59345;
  assign n59347 = ~n59344 & n59346;
  assign n59348 = ~n59343 & ~n59347;
  assign n59349 = pi516 & ~n59348;
  assign n59350 = ~n59341 & ~n59349;
  assign n59351 = ~pi238 & n59350;
  assign n59352 = ~pi517 & ~n59351;
  assign n59353 = ~n59160 & ~n59343;
  assign n59354 = ~pi238 & n59353;
  assign n59355 = ~pi247 & ~pi516;
  assign n59356 = pi247 & pi516;
  assign n59357 = ~n59355 & ~n59356;
  assign n59358 = n59336 & ~n59357;
  assign n59359 = pi238 & n59358;
  assign n59360 = pi517 & ~n59359;
  assign n59361 = ~n59354 & n59360;
  assign n59362 = ~pi507 & ~n59361;
  assign n59363 = ~n59352 & n59362;
  assign n59364 = pi238 & n59350;
  assign n59365 = pi517 & ~n59364;
  assign n59366 = pi238 & n59353;
  assign n59367 = ~pi238 & n59358;
  assign n59368 = ~pi517 & ~n59367;
  assign n59369 = ~n59366 & n59368;
  assign n59370 = pi507 & ~n59369;
  assign n59371 = ~n59365 & n59370;
  assign n59372 = ~n59363 & ~n59371;
  assign n59373 = pi233 & ~n59372;
  assign n59374 = ~pi247 & ~pi561;
  assign n59375 = ~pi240 & ~pi542;
  assign n59376 = pi240 & pi542;
  assign n59377 = ~n59375 & ~n59376;
  assign n59378 = ~pi505 & ~n58593;
  assign n59379 = pi505 & ~n59096;
  assign n59380 = ~pi246 & pi499;
  assign n59381 = pi241 & ~pi500;
  assign n59382 = ~n59380 & ~n59381;
  assign n59383 = pi249 & ~pi496;
  assign n59384 = ~pi249 & pi496;
  assign n59385 = ~pi249 & ~pi496;
  assign n59386 = pi249 & pi496;
  assign n59387 = ~n59385 & ~n59386;
  assign n59388 = ~n59383 & ~n59384;
  assign n59389 = n59382 & ~n65763;
  assign n59390 = ~pi248 & ~pi501;
  assign n59391 = pi248 & pi501;
  assign n59392 = ~n59390 & ~n59391;
  assign n59393 = ~pi241 & pi500;
  assign n59394 = pi246 & ~pi499;
  assign n59395 = ~n59393 & ~n59394;
  assign n59396 = ~n59392 & n59395;
  assign n59397 = ~pi246 & ~pi499;
  assign n59398 = pi246 & pi499;
  assign n59399 = ~n59380 & ~n59394;
  assign n59400 = ~n59397 & ~n59398;
  assign n59401 = pi248 & ~pi501;
  assign n59402 = ~n59384 & ~n59401;
  assign n59403 = n65764 & n59402;
  assign n59404 = ~pi241 & ~pi500;
  assign n59405 = pi241 & pi500;
  assign n59406 = ~n59404 & ~n59405;
  assign n59407 = ~pi248 & pi501;
  assign n59408 = ~n59383 & ~n59407;
  assign n59409 = ~n59406 & n59408;
  assign n59410 = n59403 & n59409;
  assign n59411 = ~n59392 & n65764;
  assign n59412 = ~n65763 & ~n59406;
  assign n59413 = n59411 & n59412;
  assign n59414 = n59389 & n59396;
  assign n59415 = ~n59379 & n65765;
  assign n59416 = ~n65763 & n65764;
  assign n59417 = ~n65763 & ~n59392;
  assign n59418 = n65764 & n59417;
  assign n59419 = ~n59392 & n59416;
  assign n59420 = ~n59378 & n65766;
  assign n59421 = ~n59379 & n65766;
  assign n59422 = ~n59378 & n59421;
  assign n59423 = ~n59379 & n59420;
  assign n59424 = ~n59406 & n65767;
  assign n59425 = ~n59378 & n59415;
  assign n59426 = ~n59377 & n65768;
  assign n59427 = pi497 & n59426;
  assign n59428 = ~pi239 & ~n59427;
  assign n59429 = ~pi497 & n59426;
  assign n59430 = pi239 & ~n59429;
  assign n59431 = ~n59428 & ~n59430;
  assign n59432 = pi539 & n59431;
  assign n59433 = pi242 & ~n59432;
  assign n59434 = ~pi539 & n59431;
  assign n59435 = ~pi242 & ~n59434;
  assign n59436 = ~n59433 & ~n59435;
  assign n59437 = pi540 & n59436;
  assign n59438 = pi235 & ~n59437;
  assign n59439 = ~pi540 & n59436;
  assign n59440 = ~pi235 & ~n59439;
  assign n59441 = ~n59438 & ~n59440;
  assign n59442 = ~pi244 & ~pi541;
  assign n59443 = pi244 & pi541;
  assign n59444 = ~n59442 & ~n59443;
  assign n59445 = n59441 & ~n59444;
  assign n59446 = ~pi245 & ~pi503;
  assign n59447 = pi245 & pi503;
  assign n59448 = ~n59446 & ~n59447;
  assign n59449 = n59445 & ~n59448;
  assign n59450 = ~pi502 & n59449;
  assign n59451 = ~pi247 & ~n59450;
  assign n59452 = ~n59374 & ~n59451;
  assign n59453 = ~pi518 & ~n58615;
  assign n59454 = pi518 & ~n59162;
  assign n59455 = ~pi248 & pi521;
  assign n59456 = pi241 & ~pi574;
  assign n59457 = ~n59455 & ~n59456;
  assign n59458 = pi249 & ~pi578;
  assign n59459 = ~pi249 & pi578;
  assign n59460 = ~pi249 & ~pi578;
  assign n59461 = pi249 & pi578;
  assign n59462 = ~n59460 & ~n59461;
  assign n59463 = ~n59458 & ~n59459;
  assign n59464 = n59457 & ~n65769;
  assign n59465 = ~pi246 & ~pi520;
  assign n59466 = pi246 & pi520;
  assign n59467 = pi246 & ~pi520;
  assign n59468 = ~pi246 & pi520;
  assign n59469 = ~n59467 & ~n59468;
  assign n59470 = ~n59465 & ~n59466;
  assign n59471 = ~pi241 & pi574;
  assign n59472 = pi248 & ~pi521;
  assign n59473 = ~n59471 & ~n59472;
  assign n59474 = n65770 & n59473;
  assign n59475 = ~pi248 & ~pi521;
  assign n59476 = pi248 & pi521;
  assign n59477 = ~n59475 & ~n59476;
  assign n59478 = ~n59455 & ~n59472;
  assign n59479 = ~n65769 & ~n65771;
  assign n59480 = pi241 & pi574;
  assign n59481 = ~pi241 & ~pi574;
  assign n59482 = ~n59480 & ~n59481;
  assign n59483 = n65770 & ~n59482;
  assign n59484 = n59479 & n59483;
  assign n59485 = ~n59459 & ~n59467;
  assign n59486 = ~n65771 & n59485;
  assign n59487 = ~n59458 & ~n59468;
  assign n59488 = ~n59482 & n59487;
  assign n59489 = n59486 & n59488;
  assign n59490 = n65770 & ~n65771;
  assign n59491 = ~n65769 & ~n59482;
  assign n59492 = n59490 & n59491;
  assign n59493 = n59464 & n59474;
  assign n59494 = ~n59454 & n65772;
  assign n59495 = ~n59453 & n65772;
  assign n59496 = ~n59454 & n59495;
  assign n59497 = ~n59453 & n59494;
  assign n59498 = pi582 & n65773;
  assign n59499 = pi240 & ~n59498;
  assign n59500 = ~pi582 & n65773;
  assign n59501 = ~pi240 & ~n59500;
  assign n59502 = ~n59499 & ~n59501;
  assign n59503 = pi239 & ~pi519;
  assign n59504 = ~pi239 & pi519;
  assign n59505 = ~n59503 & ~n59504;
  assign n59506 = n59502 & ~n59505;
  assign n59507 = ~pi242 & ~pi586;
  assign n59508 = pi242 & pi586;
  assign n59509 = ~n59507 & ~n59508;
  assign n59510 = n59506 & ~n59509;
  assign n59511 = ~pi235 & ~pi581;
  assign n59512 = pi235 & pi581;
  assign n59513 = ~n59511 & ~n59512;
  assign n59514 = n59510 & ~n59513;
  assign n59515 = pi585 & n59514;
  assign n59516 = pi244 & ~n59515;
  assign n59517 = ~pi585 & n59514;
  assign n59518 = ~pi244 & ~n59517;
  assign n59519 = ~n59516 & ~n59518;
  assign n59520 = pi584 & n59519;
  assign n59521 = pi245 & ~n59520;
  assign n59522 = ~pi542 & n65768;
  assign n59523 = n59501 & ~n59522;
  assign n59524 = pi542 & n65768;
  assign n59525 = n59499 & ~n59524;
  assign n59526 = ~pi500 & n65768;
  assign n59527 = n59405 & n65767;
  assign n59528 = ~n65773 & ~n59527;
  assign n59529 = ~n59526 & n59528;
  assign n59530 = ~pi582 & ~n59529;
  assign n59531 = pi582 & n65768;
  assign n59532 = ~pi240 & ~n59531;
  assign n59533 = ~n59530 & n59532;
  assign n59534 = ~n59499 & ~n59533;
  assign n59535 = ~pi542 & ~n59534;
  assign n59536 = pi582 & ~n59529;
  assign n59537 = ~pi582 & n65768;
  assign n59538 = pi240 & ~n59537;
  assign n59539 = ~n59536 & n59538;
  assign n59540 = ~n59501 & ~n59539;
  assign n59541 = pi542 & ~n59540;
  assign n59542 = ~n59535 & ~n59541;
  assign n59543 = ~n59523 & ~n59525;
  assign n59544 = ~pi497 & n65774;
  assign n59545 = pi497 & n59502;
  assign n59546 = pi239 & ~n59545;
  assign n59547 = ~n59544 & n59546;
  assign n59548 = ~n59428 & ~n59547;
  assign n59549 = ~pi519 & ~n59548;
  assign n59550 = pi497 & n65774;
  assign n59551 = ~pi497 & n59502;
  assign n59552 = ~pi239 & ~n59551;
  assign n59553 = ~n59550 & n59552;
  assign n59554 = ~n59430 & ~n59553;
  assign n59555 = pi519 & ~n59554;
  assign n59556 = ~n59549 & ~n59555;
  assign n59557 = ~pi539 & n59556;
  assign n59558 = pi539 & n59506;
  assign n59559 = ~pi242 & ~n59558;
  assign n59560 = ~n59557 & n59559;
  assign n59561 = ~n59433 & ~n59560;
  assign n59562 = ~pi586 & ~n59561;
  assign n59563 = pi539 & n59556;
  assign n59564 = ~pi539 & n59506;
  assign n59565 = pi242 & ~n59564;
  assign n59566 = ~n59563 & n59565;
  assign n59567 = ~n59435 & ~n59566;
  assign n59568 = pi586 & ~n59567;
  assign n59569 = ~n59562 & ~n59568;
  assign n59570 = ~pi540 & n59569;
  assign n59571 = pi540 & n59510;
  assign n59572 = ~pi235 & ~n59571;
  assign n59573 = ~n59570 & n59572;
  assign n59574 = ~n59438 & ~n59573;
  assign n59575 = ~pi581 & ~n59574;
  assign n59576 = pi540 & n59569;
  assign n59577 = ~pi540 & n59510;
  assign n59578 = pi235 & ~n59577;
  assign n59579 = ~n59576 & n59578;
  assign n59580 = ~n59440 & ~n59579;
  assign n59581 = pi581 & ~n59580;
  assign n59582 = ~n59575 & ~n59581;
  assign n59583 = ~pi585 & n59582;
  assign n59584 = pi585 & n59441;
  assign n59585 = ~pi244 & ~n59584;
  assign n59586 = ~n59583 & n59585;
  assign n59587 = ~n59516 & ~n59586;
  assign n59588 = ~pi541 & ~n59587;
  assign n59589 = pi585 & n59582;
  assign n59590 = ~pi585 & n59441;
  assign n59591 = pi244 & ~n59590;
  assign n59592 = ~n59589 & n59591;
  assign n59593 = ~n59518 & ~n59592;
  assign n59594 = pi541 & ~n59593;
  assign n59595 = ~n59588 & ~n59594;
  assign n59596 = ~pi584 & n59595;
  assign n59597 = pi584 & n59445;
  assign n59598 = ~pi245 & ~n59597;
  assign n59599 = ~n59596 & n59598;
  assign n59600 = ~n59521 & ~n59599;
  assign n59601 = ~pi503 & ~n59600;
  assign n59602 = ~pi584 & n59519;
  assign n59603 = ~pi245 & ~n59602;
  assign n59604 = pi584 & n59595;
  assign n59605 = ~pi584 & n59445;
  assign n59606 = pi245 & ~n59605;
  assign n59607 = ~n59604 & n59606;
  assign n59608 = ~n59603 & ~n59607;
  assign n59609 = pi503 & ~n59608;
  assign n59610 = ~n59601 & ~n59609;
  assign n59611 = ~pi502 & ~n59610;
  assign n59612 = ~n59521 & ~n59603;
  assign n59613 = pi502 & ~n59612;
  assign n59614 = ~pi561 & ~n59613;
  assign n59615 = ~n59611 & n59614;
  assign n59616 = ~n59452 & ~n59615;
  assign n59617 = pi247 & pi561;
  assign n59618 = pi502 & n59449;
  assign n59619 = pi247 & ~n59618;
  assign n59620 = ~n59617 & ~n59619;
  assign n59621 = pi502 & ~n59610;
  assign n59622 = ~pi502 & ~n59612;
  assign n59623 = pi561 & ~n59622;
  assign n59624 = ~n59621 & n59623;
  assign n59625 = ~n59620 & ~n59624;
  assign n59626 = ~n59616 & ~n59625;
  assign n59627 = ~pi238 & n59626;
  assign n59628 = ~pi522 & ~n59627;
  assign n59629 = ~n59451 & ~n59619;
  assign n59630 = ~pi238 & n59629;
  assign n59631 = ~n59374 & ~n59617;
  assign n59632 = n59612 & ~n59631;
  assign n59633 = pi238 & n59632;
  assign n59634 = pi522 & ~n59633;
  assign n59635 = ~n59630 & n59634;
  assign n59636 = ~pi543 & ~n59635;
  assign n59637 = ~n59628 & n59636;
  assign n59638 = pi238 & n59626;
  assign n59639 = pi522 & ~n59638;
  assign n59640 = pi238 & n59629;
  assign n59641 = ~pi238 & n59632;
  assign n59642 = ~pi522 & ~n59641;
  assign n59643 = ~n59640 & n59642;
  assign n59644 = pi543 & ~n59643;
  assign n59645 = ~n59639 & n59644;
  assign n59646 = ~n59637 & ~n59645;
  assign n59647 = ~pi233 & ~n59646;
  assign n59648 = pi237 & ~n59647;
  assign n59649 = ~n59373 & n59648;
  assign n59650 = ~pi240 & ~pi492;
  assign n59651 = pi240 & pi492;
  assign n59652 = ~n59650 & ~n59651;
  assign n59653 = ~pi241 & ~pi490;
  assign n59654 = pi241 & pi490;
  assign n59655 = ~n59653 & ~n59654;
  assign n59656 = pi544 & ~n59096;
  assign n59657 = ~pi544 & ~n58593;
  assign n59658 = ~pi246 & ~pi546;
  assign n59659 = pi246 & pi546;
  assign n59660 = ~n59658 & ~n59659;
  assign n59661 = pi248 & ~pi548;
  assign n59662 = ~pi248 & pi548;
  assign n59663 = pi248 & pi548;
  assign n59664 = ~pi248 & ~pi548;
  assign n59665 = ~n59663 & ~n59664;
  assign n59666 = ~n59661 & ~n59662;
  assign n59667 = pi249 & ~pi484;
  assign n59668 = ~pi249 & pi484;
  assign n59669 = pi249 & pi484;
  assign n59670 = ~pi249 & ~pi484;
  assign n59671 = ~n59669 & ~n59670;
  assign n59672 = ~n59667 & ~n59668;
  assign n59673 = ~n65775 & ~n65776;
  assign n59674 = ~n59660 & ~n65775;
  assign n59675 = ~n65776 & n59674;
  assign n59676 = ~n59660 & n59673;
  assign n59677 = ~n59657 & n65777;
  assign n59678 = ~n59656 & n65777;
  assign n59679 = ~n59657 & n59678;
  assign n59680 = ~n59656 & n59677;
  assign n59681 = ~n59655 & n65778;
  assign n59682 = ~n59652 & n59681;
  assign n59683 = pi494 & n59682;
  assign n59684 = ~pi239 & ~n59683;
  assign n59685 = ~pi494 & n59682;
  assign n59686 = pi239 & ~n59685;
  assign n59687 = ~n59684 & ~n59686;
  assign n59688 = pi483 & n59687;
  assign n59689 = pi242 & ~n59688;
  assign n59690 = ~pi483 & n59687;
  assign n59691 = ~pi242 & ~n59690;
  assign n59692 = ~n59689 & ~n59691;
  assign n59693 = pi495 & n59692;
  assign n59694 = pi235 & ~n59693;
  assign n59695 = ~pi495 & n59692;
  assign n59696 = ~pi235 & ~n59695;
  assign n59697 = ~n59694 & ~n59696;
  assign n59698 = ~pi244 & ~pi493;
  assign n59699 = pi244 & pi493;
  assign n59700 = ~n59698 & ~n59699;
  assign n59701 = n59697 & ~n59700;
  assign n59702 = pi545 & n59701;
  assign n59703 = pi245 & ~n59702;
  assign n59704 = ~pi545 & n59701;
  assign n59705 = ~pi245 & ~n59704;
  assign n59706 = ~n59703 & ~n59705;
  assign n59707 = pi547 & n59706;
  assign n59708 = pi247 & ~n59707;
  assign n59709 = ~pi523 & ~n58615;
  assign n59710 = pi523 & ~n59162;
  assign n59711 = ~pi246 & ~pi526;
  assign n59712 = pi246 & pi526;
  assign n59713 = ~n59711 & ~n59712;
  assign n59714 = pi248 & ~pi576;
  assign n59715 = ~pi248 & pi576;
  assign n59716 = pi248 & pi576;
  assign n59717 = ~pi248 & ~pi576;
  assign n59718 = ~n59716 & ~n59717;
  assign n59719 = ~n59714 & ~n59715;
  assign n59720 = pi249 & ~pi528;
  assign n59721 = ~pi249 & pi528;
  assign n59722 = pi249 & pi528;
  assign n59723 = ~pi249 & ~pi528;
  assign n59724 = ~n59722 & ~n59723;
  assign n59725 = ~n59720 & ~n59721;
  assign n59726 = ~n65779 & ~n65780;
  assign n59727 = ~n59713 & ~n65779;
  assign n59728 = ~n65780 & n59727;
  assign n59729 = ~n59713 & n59726;
  assign n59730 = ~n59710 & n65781;
  assign n59731 = ~n59709 & n65781;
  assign n59732 = ~n59710 & n59731;
  assign n59733 = ~n59709 & n59730;
  assign n59734 = pi571 & n65782;
  assign n59735 = pi241 & ~n59734;
  assign n59736 = ~pi571 & n65782;
  assign n59737 = ~pi241 & ~n59736;
  assign n59738 = ~n59735 & ~n59737;
  assign n59739 = ~pi530 & n59738;
  assign n59740 = ~pi240 & ~n59739;
  assign n59741 = pi530 & n59738;
  assign n59742 = pi240 & ~n59741;
  assign n59743 = ~n59740 & ~n59742;
  assign n59744 = pi239 & ~pi524;
  assign n59745 = ~pi239 & pi524;
  assign n59746 = ~n59744 & ~n59745;
  assign n59747 = n59743 & ~n59746;
  assign n59748 = ~pi242 & ~pi573;
  assign n59749 = pi242 & pi573;
  assign n59750 = ~n59748 & ~n59749;
  assign n59751 = n59747 & ~n59750;
  assign n59752 = ~pi235 & ~pi575;
  assign n59753 = pi235 & pi575;
  assign n59754 = ~n59752 & ~n59753;
  assign n59755 = n59751 & ~n59754;
  assign n59756 = pi572 & n59755;
  assign n59757 = pi244 & ~n59756;
  assign n59758 = ~n59650 & ~n59740;
  assign n59759 = ~pi490 & n65778;
  assign n59760 = n59737 & ~n59759;
  assign n59761 = pi490 & n65778;
  assign n59762 = n59735 & ~n59761;
  assign n59763 = ~pi241 & ~n65778;
  assign n59764 = ~n59736 & n59763;
  assign n59765 = ~n59735 & ~n59764;
  assign n59766 = ~pi490 & ~n59765;
  assign n59767 = pi241 & ~n65778;
  assign n59768 = ~n59734 & n59767;
  assign n59769 = ~n59737 & ~n59768;
  assign n59770 = pi490 & ~n59769;
  assign n59771 = ~n59766 & ~n59770;
  assign n59772 = ~n59760 & ~n59762;
  assign n59773 = ~pi530 & ~n65783;
  assign n59774 = pi530 & ~n59681;
  assign n59775 = ~pi492 & ~n59774;
  assign n59776 = ~n59773 & n59775;
  assign n59777 = ~n59758 & ~n59776;
  assign n59778 = ~n59651 & ~n59742;
  assign n59779 = pi530 & ~n65783;
  assign n59780 = ~pi530 & ~n59681;
  assign n59781 = pi492 & ~n59780;
  assign n59782 = ~n59779 & n59781;
  assign n59783 = ~n59778 & ~n59782;
  assign n59784 = ~n59777 & ~n59783;
  assign n59785 = ~pi494 & n59784;
  assign n59786 = pi494 & n59743;
  assign n59787 = pi239 & ~n59786;
  assign n59788 = ~n59785 & n59787;
  assign n59789 = ~n59684 & ~n59788;
  assign n59790 = ~pi524 & ~n59789;
  assign n59791 = pi494 & n59784;
  assign n59792 = ~pi494 & n59743;
  assign n59793 = ~pi239 & ~n59792;
  assign n59794 = ~n59791 & n59793;
  assign n59795 = ~n59686 & ~n59794;
  assign n59796 = pi524 & ~n59795;
  assign n59797 = ~n59790 & ~n59796;
  assign n59798 = ~pi483 & n59797;
  assign n59799 = pi483 & n59747;
  assign n59800 = ~pi242 & ~n59799;
  assign n59801 = ~n59798 & n59800;
  assign n59802 = ~n59689 & ~n59801;
  assign n59803 = ~pi573 & ~n59802;
  assign n59804 = pi483 & n59797;
  assign n59805 = ~pi483 & n59747;
  assign n59806 = pi242 & ~n59805;
  assign n59807 = ~n59804 & n59806;
  assign n59808 = ~n59691 & ~n59807;
  assign n59809 = pi573 & ~n59808;
  assign n59810 = ~n59803 & ~n59809;
  assign n59811 = ~pi495 & n59810;
  assign n59812 = pi495 & n59751;
  assign n59813 = ~pi235 & ~n59812;
  assign n59814 = ~n59811 & n59813;
  assign n59815 = ~n59694 & ~n59814;
  assign n59816 = ~pi575 & ~n59815;
  assign n59817 = pi495 & n59810;
  assign n59818 = ~pi495 & n59751;
  assign n59819 = pi235 & ~n59818;
  assign n59820 = ~n59817 & n59819;
  assign n59821 = ~n59696 & ~n59820;
  assign n59822 = pi575 & ~n59821;
  assign n59823 = ~n59816 & ~n59822;
  assign n59824 = ~pi572 & n59823;
  assign n59825 = pi572 & n59697;
  assign n59826 = ~pi244 & ~n59825;
  assign n59827 = ~n59824 & n59826;
  assign n59828 = ~n59757 & ~n59827;
  assign n59829 = ~pi493 & ~n59828;
  assign n59830 = ~pi572 & n59755;
  assign n59831 = ~pi244 & ~n59830;
  assign n59832 = pi572 & n59823;
  assign n59833 = ~pi572 & n59697;
  assign n59834 = pi244 & ~n59833;
  assign n59835 = ~n59832 & n59834;
  assign n59836 = ~n59831 & ~n59835;
  assign n59837 = pi493 & ~n59836;
  assign n59838 = ~n59829 & ~n59837;
  assign n59839 = ~pi545 & n59838;
  assign n59840 = ~n59757 & ~n59831;
  assign n59841 = pi545 & n59840;
  assign n59842 = ~pi245 & ~n59841;
  assign n59843 = ~n59839 & n59842;
  assign n59844 = ~n59703 & ~n59843;
  assign n59845 = ~pi525 & ~n59844;
  assign n59846 = pi545 & n59838;
  assign n59847 = ~pi545 & n59840;
  assign n59848 = pi245 & ~n59847;
  assign n59849 = ~n59846 & n59848;
  assign n59850 = ~n59705 & ~n59849;
  assign n59851 = pi525 & ~n59850;
  assign n59852 = ~n59845 & ~n59851;
  assign n59853 = ~pi547 & n59852;
  assign n59854 = ~pi245 & ~pi525;
  assign n59855 = pi245 & pi525;
  assign n59856 = ~n59854 & ~n59855;
  assign n59857 = n59840 & ~n59856;
  assign n59858 = pi547 & n59857;
  assign n59859 = ~pi247 & ~n59858;
  assign n59860 = ~n59853 & n59859;
  assign n59861 = ~n59708 & ~n59860;
  assign n59862 = ~pi527 & ~n59861;
  assign n59863 = ~pi547 & n59706;
  assign n59864 = ~pi247 & ~n59863;
  assign n59865 = pi547 & n59852;
  assign n59866 = ~pi547 & n59857;
  assign n59867 = pi247 & ~n59866;
  assign n59868 = ~n59865 & n59867;
  assign n59869 = ~n59864 & ~n59868;
  assign n59870 = pi527 & ~n59869;
  assign n59871 = ~n59862 & ~n59870;
  assign n59872 = ~pi238 & n59871;
  assign n59873 = ~pi529 & ~n59872;
  assign n59874 = ~n59708 & ~n59864;
  assign n59875 = ~pi238 & n59874;
  assign n59876 = ~pi247 & ~pi527;
  assign n59877 = pi247 & pi527;
  assign n59878 = ~n59876 & ~n59877;
  assign n59879 = n59857 & ~n59878;
  assign n59880 = pi238 & n59879;
  assign n59881 = pi529 & ~n59880;
  assign n59882 = ~n59875 & n59881;
  assign n59883 = ~pi491 & ~n59882;
  assign n59884 = ~n59873 & n59883;
  assign n59885 = pi238 & n59871;
  assign n59886 = pi529 & ~n59885;
  assign n59887 = pi238 & n59874;
  assign n59888 = ~pi238 & n59879;
  assign n59889 = ~pi529 & ~n59888;
  assign n59890 = ~n59887 & n59889;
  assign n59891 = pi491 & ~n59890;
  assign n59892 = ~n59886 & n59891;
  assign n59893 = ~n59884 & ~n59892;
  assign n59894 = pi233 & ~n59893;
  assign n59895 = pi485 & ~n59096;
  assign n59896 = ~pi485 & ~n58593;
  assign n59897 = ~pi246 & pi563;
  assign n59898 = ~pi249 & pi555;
  assign n59899 = ~n59897 & ~n59898;
  assign n59900 = ~pi239 & ~pi550;
  assign n59901 = ~pi242 & pi489;
  assign n59902 = ~n59900 & ~n59901;
  assign n59903 = pi242 & ~pi489;
  assign n59904 = pi240 & ~pi551;
  assign n59905 = ~n59903 & ~n59904;
  assign n59906 = n59902 & n59905;
  assign n59907 = n59899 & n59906;
  assign n59908 = ~pi248 & pi554;
  assign n59909 = pi241 & ~pi553;
  assign n59910 = ~n59908 & ~n59909;
  assign n59911 = pi239 & pi550;
  assign n59912 = pi246 & ~pi563;
  assign n59913 = ~n59911 & ~n59912;
  assign n59914 = n59910 & n59913;
  assign n59915 = ~pi241 & pi553;
  assign n59916 = pi249 & ~pi555;
  assign n59917 = ~n59915 & ~n59916;
  assign n59918 = ~pi240 & pi551;
  assign n59919 = pi248 & ~pi554;
  assign n59920 = ~n59918 & ~n59919;
  assign n59921 = n59917 & n59920;
  assign n59922 = n59914 & n59921;
  assign n59923 = ~pi246 & ~pi563;
  assign n59924 = pi246 & pi563;
  assign n59925 = ~n59923 & ~n59924;
  assign n59926 = ~n59897 & ~n59912;
  assign n59927 = pi239 & ~pi550;
  assign n59928 = ~pi239 & pi550;
  assign n59929 = ~n59900 & ~n59911;
  assign n59930 = ~n59927 & ~n59928;
  assign n59931 = n59917 & n65785;
  assign n59932 = ~n65784 & n59931;
  assign n59933 = ~n59903 & ~n59918;
  assign n59934 = ~n59904 & ~n59909;
  assign n59935 = n59933 & n59934;
  assign n59936 = ~n59898 & ~n59908;
  assign n59937 = ~n59901 & ~n59919;
  assign n59938 = n59936 & n59937;
  assign n59939 = n59935 & n59938;
  assign n59940 = n59932 & n59939;
  assign n59941 = n59907 & n59922;
  assign n59942 = ~n59896 & n65786;
  assign n59943 = ~pi249 & ~pi555;
  assign n59944 = pi249 & pi555;
  assign n59945 = ~n59943 & ~n59944;
  assign n59946 = ~n59898 & ~n59916;
  assign n59947 = ~pi241 & ~pi553;
  assign n59948 = pi241 & pi553;
  assign n59949 = ~n59947 & ~n59948;
  assign n59950 = ~n59909 & ~n59915;
  assign n59951 = ~n65787 & ~n65788;
  assign n59952 = pi240 & pi551;
  assign n59953 = ~pi240 & ~pi551;
  assign n59954 = ~n59952 & ~n59953;
  assign n59955 = ~n59908 & ~n59919;
  assign n59956 = ~n65784 & n59955;
  assign n59957 = ~n59954 & n59956;
  assign n59958 = n59951 & ~n59954;
  assign n59959 = n59956 & n59958;
  assign n59960 = n59951 & n59957;
  assign n59961 = ~n59896 & n65789;
  assign n59962 = ~n59895 & n65789;
  assign n59963 = ~n59896 & n59962;
  assign n59964 = ~n59895 & n59961;
  assign n59965 = pi550 & n65790;
  assign n59966 = ~pi239 & ~n59965;
  assign n59967 = ~pi550 & n65790;
  assign n59968 = pi239 & ~n59967;
  assign n59969 = ~n59966 & ~n59968;
  assign n59970 = n65785 & n65790;
  assign n59971 = ~pi489 & n65791;
  assign n59972 = ~pi242 & ~n59971;
  assign n59973 = pi489 & n65791;
  assign n59974 = pi242 & ~n59973;
  assign n59975 = ~n59972 & ~n59974;
  assign n59976 = ~n59895 & n59942;
  assign n59977 = pi549 & n65792;
  assign n59978 = pi235 & ~n59977;
  assign n59979 = ~pi549 & n65792;
  assign n59980 = ~pi235 & ~n59979;
  assign n59981 = ~n59978 & ~n59980;
  assign n59982 = pi486 & n59981;
  assign n59983 = pi244 & ~n59982;
  assign n59984 = ~pi486 & n59981;
  assign n59985 = ~pi244 & ~n59984;
  assign n59986 = ~n59983 & ~n59985;
  assign n59987 = ~pi245 & ~pi580;
  assign n59988 = pi245 & pi580;
  assign n59989 = ~n59987 & ~n59988;
  assign n59990 = n59986 & ~n59989;
  assign n59991 = pi552 & n59990;
  assign n59992 = pi247 & ~n59991;
  assign n59993 = ~pi235 & ~pi531;
  assign n59994 = pi235 & pi531;
  assign n59995 = ~n59993 & ~n59994;
  assign n59996 = ~pi570 & ~n58615;
  assign n59997 = pi570 & ~n59162;
  assign n59998 = ~pi242 & ~pi556;
  assign n59999 = pi242 & pi556;
  assign n60000 = ~n59998 & ~n59999;
  assign n60001 = pi239 & pi569;
  assign n60002 = pi240 & ~pi560;
  assign n60003 = ~n60001 & ~n60002;
  assign n60004 = ~pi249 & pi482;
  assign n60005 = pi241 & ~pi562;
  assign n60006 = ~n60004 & ~n60005;
  assign n60007 = n60003 & n60006;
  assign n60008 = ~n60000 & n60007;
  assign n60009 = ~pi246 & pi564;
  assign n60010 = ~pi241 & pi562;
  assign n60011 = ~n60009 & ~n60010;
  assign n60012 = pi248 & ~pi565;
  assign n60013 = ~pi239 & ~pi569;
  assign n60014 = ~n60012 & ~n60013;
  assign n60015 = n60011 & n60014;
  assign n60016 = ~pi248 & pi565;
  assign n60017 = pi246 & ~pi564;
  assign n60018 = ~n60016 & ~n60017;
  assign n60019 = ~pi240 & pi560;
  assign n60020 = pi249 & ~pi482;
  assign n60021 = ~n60019 & ~n60020;
  assign n60022 = n60018 & n60021;
  assign n60023 = n60015 & n60022;
  assign n60024 = ~pi242 & pi556;
  assign n60025 = ~n60012 & ~n60024;
  assign n60026 = ~pi239 & pi569;
  assign n60027 = pi239 & ~pi569;
  assign n60028 = ~n60001 & ~n60013;
  assign n60029 = ~n60026 & ~n60027;
  assign n60030 = ~n60002 & ~n60010;
  assign n60031 = n65793 & n60030;
  assign n60032 = n60025 & n60031;
  assign n60033 = ~n60009 & ~n60020;
  assign n60034 = pi242 & ~pi556;
  assign n60035 = ~n60019 & ~n60034;
  assign n60036 = n60033 & n60035;
  assign n60037 = ~n60004 & ~n60017;
  assign n60038 = ~n60005 & ~n60016;
  assign n60039 = n60037 & n60038;
  assign n60040 = n60036 & n60039;
  assign n60041 = n60032 & n60040;
  assign n60042 = n60008 & n60023;
  assign n60043 = ~n59997 & n65794;
  assign n60044 = ~n60009 & ~n60012;
  assign n60045 = ~n60016 & ~n60020;
  assign n60046 = n60044 & n60045;
  assign n60047 = pi241 & pi562;
  assign n60048 = ~pi241 & ~pi562;
  assign n60049 = ~n60047 & ~n60048;
  assign n60050 = pi240 & pi560;
  assign n60051 = ~pi240 & ~pi560;
  assign n60052 = ~n60050 & ~n60051;
  assign n60053 = n60037 & ~n60052;
  assign n60054 = ~n60049 & n60053;
  assign n60055 = n60046 & n60054;
  assign n60056 = ~n59997 & n60055;
  assign n60057 = ~n60004 & ~n60009;
  assign n60058 = ~n60004 & n60033;
  assign n60059 = ~n60020 & n60057;
  assign n60060 = ~n60049 & n65795;
  assign n60061 = ~n59996 & n60060;
  assign n60062 = ~n59997 & n60060;
  assign n60063 = ~n59996 & n60062;
  assign n60064 = ~n59997 & n60061;
  assign n60065 = ~n60012 & ~n60016;
  assign n60066 = ~n60017 & ~n60052;
  assign n60067 = ~n60017 & n60065;
  assign n60068 = ~n60052 & n60067;
  assign n60069 = n60065 & n60066;
  assign n60070 = n65796 & n65797;
  assign n60071 = ~n59996 & n60056;
  assign n60072 = n65793 & n65798;
  assign n60073 = ~n60000 & n60072;
  assign n60074 = ~n59996 & n60043;
  assign n60075 = ~n59995 & n65799;
  assign n60076 = ~pi244 & ~pi566;
  assign n60077 = pi244 & pi566;
  assign n60078 = ~n60076 & ~n60077;
  assign n60079 = n60075 & ~n60078;
  assign n60080 = pi568 & n60079;
  assign n60081 = pi245 & ~n60080;
  assign n60082 = ~pi531 & n65799;
  assign n60083 = n59980 & ~n60082;
  assign n60084 = pi531 & n65799;
  assign n60085 = n59978 & ~n60084;
  assign n60086 = ~n59972 & ~n59998;
  assign n60087 = n59927 & n65790;
  assign n60088 = ~n65793 & ~n60087;
  assign n60089 = n65798 & ~n60088;
  assign n60090 = pi569 & ~n59968;
  assign n60091 = n65798 & n60090;
  assign n60092 = n60027 & n65798;
  assign n60093 = ~n65791 & ~n60092;
  assign n60094 = ~n60091 & n60093;
  assign n60095 = ~n65791 & ~n60089;
  assign n60096 = ~pi489 & n65800;
  assign n60097 = pi489 & ~n60072;
  assign n60098 = ~pi556 & ~n60097;
  assign n60099 = ~n60096 & n60098;
  assign n60100 = ~n60086 & ~n60099;
  assign n60101 = ~n59974 & ~n59999;
  assign n60102 = pi489 & n65800;
  assign n60103 = ~pi489 & ~n60072;
  assign n60104 = pi556 & ~n60103;
  assign n60105 = ~n60102 & n60104;
  assign n60106 = ~n60101 & ~n60105;
  assign n60107 = ~n60100 & ~n60106;
  assign n60108 = ~pi549 & n60107;
  assign n60109 = pi549 & n65799;
  assign n60110 = ~pi235 & ~n60109;
  assign n60111 = ~n60108 & n60110;
  assign n60112 = ~n59978 & ~n60111;
  assign n60113 = ~pi531 & ~n60112;
  assign n60114 = pi549 & n60107;
  assign n60115 = ~pi549 & n65799;
  assign n60116 = pi235 & ~n60115;
  assign n60117 = ~n60114 & n60116;
  assign n60118 = ~n59980 & ~n60117;
  assign n60119 = pi531 & ~n60118;
  assign n60120 = ~n60113 & ~n60119;
  assign n60121 = ~n60083 & ~n60085;
  assign n60122 = ~pi486 & n65801;
  assign n60123 = pi486 & n60075;
  assign n60124 = ~pi244 & ~n60123;
  assign n60125 = ~n60122 & n60124;
  assign n60126 = ~n59983 & ~n60125;
  assign n60127 = ~pi566 & ~n60126;
  assign n60128 = pi486 & n65801;
  assign n60129 = ~pi486 & n60075;
  assign n60130 = pi244 & ~n60129;
  assign n60131 = ~n60128 & n60130;
  assign n60132 = ~n59985 & ~n60131;
  assign n60133 = pi566 & ~n60132;
  assign n60134 = ~n60127 & ~n60133;
  assign n60135 = ~pi568 & n60134;
  assign n60136 = pi568 & n59986;
  assign n60137 = ~pi245 & ~n60136;
  assign n60138 = ~n60135 & n60137;
  assign n60139 = ~n60081 & ~n60138;
  assign n60140 = ~pi580 & ~n60139;
  assign n60141 = ~pi568 & n60079;
  assign n60142 = ~pi245 & ~n60141;
  assign n60143 = pi568 & n60134;
  assign n60144 = ~pi568 & n59986;
  assign n60145 = pi245 & ~n60144;
  assign n60146 = ~n60143 & n60145;
  assign n60147 = ~n60142 & ~n60146;
  assign n60148 = pi580 & ~n60147;
  assign n60149 = ~n60140 & ~n60148;
  assign n60150 = ~pi552 & n60149;
  assign n60151 = ~n60081 & ~n60142;
  assign n60152 = pi552 & n60151;
  assign n60153 = ~pi247 & ~n60152;
  assign n60154 = ~n60150 & n60153;
  assign n60155 = ~n59992 & ~n60154;
  assign n60156 = ~pi532 & ~n60155;
  assign n60157 = ~pi552 & n59990;
  assign n60158 = ~pi247 & ~n60157;
  assign n60159 = pi552 & n60149;
  assign n60160 = ~pi552 & n60151;
  assign n60161 = pi247 & ~n60160;
  assign n60162 = ~n60159 & n60161;
  assign n60163 = ~n60158 & ~n60162;
  assign n60164 = pi532 & ~n60163;
  assign n60165 = ~n60156 & ~n60164;
  assign n60166 = ~pi238 & n60165;
  assign n60167 = ~pi577 & ~n60166;
  assign n60168 = ~n59992 & ~n60158;
  assign n60169 = pi238 & n60168;
  assign n60170 = ~pi247 & ~pi532;
  assign n60171 = pi247 & pi532;
  assign n60172 = ~n60170 & ~n60171;
  assign n60173 = n60151 & ~n60172;
  assign n60174 = ~pi238 & n60173;
  assign n60175 = pi577 & ~n60174;
  assign n60176 = ~n60169 & n60175;
  assign n60177 = ~pi498 & ~n60176;
  assign n60178 = ~n60167 & n60177;
  assign n60179 = pi238 & n60165;
  assign n60180 = pi577 & ~n60179;
  assign n60181 = ~pi238 & n60168;
  assign n60182 = pi238 & n60173;
  assign n60183 = ~pi577 & ~n60182;
  assign n60184 = ~n60181 & n60183;
  assign n60185 = pi498 & ~n60184;
  assign n60186 = ~n60180 & n60185;
  assign n60187 = ~n60178 & ~n60186;
  assign n60188 = ~pi233 & ~n60187;
  assign n60189 = ~pi237 & ~n60188;
  assign n60190 = ~n59894 & n60189;
  assign po750 = ~n59649 & ~n60190;
  assign n60192 = pi534 & ~n47953;
  assign n60193 = ~pi239 & n47953;
  assign po691 = ~n60192 & ~n60193;
  assign n60195 = pi535 & ~n47953;
  assign n60196 = pi240 & n47953;
  assign n60197 = ~n60195 & ~n60196;
  assign n60198 = pi536 & ~n47953;
  assign n60199 = pi246 & n47953;
  assign n60200 = ~n60198 & ~n60199;
  assign n60201 = pi537 & ~n47953;
  assign n60202 = pi248 & n47953;
  assign n60203 = ~n60201 & ~n60202;
  assign n60204 = pi538 & ~n47953;
  assign n60205 = pi249 & n47953;
  assign n60206 = ~n60204 & ~n60205;
  assign n60207 = pi539 & ~n47960;
  assign n60208 = pi242 & n47960;
  assign n60209 = ~n60207 & ~n60208;
  assign n60210 = pi540 & ~n47960;
  assign n60211 = pi235 & n47960;
  assign n60212 = ~n60210 & ~n60211;
  assign n60213 = pi541 & ~n47960;
  assign n60214 = pi244 & n47960;
  assign n60215 = ~n60213 & ~n60214;
  assign n60216 = pi542 & ~n47960;
  assign n60217 = pi240 & n47960;
  assign n60218 = ~n60216 & ~n60217;
  assign n60219 = pi543 & ~n47960;
  assign n60220 = pi238 & n47960;
  assign n60221 = ~n60219 & ~n60220;
  assign n60222 = pi544 & ~n47968;
  assign n60223 = n47963 & n58591;
  assign n60224 = n47968 & n58593;
  assign n60225 = pi544 & ~n60224;
  assign n60226 = ~pi544 & n47963;
  assign n60227 = n58591 & n60226;
  assign n60228 = ~n60225 & ~n60227;
  assign n60229 = ~n60222 & ~n60223;
  assign n60230 = pi545 & ~n47968;
  assign n60231 = pi245 & n47968;
  assign n60232 = ~n60230 & ~n60231;
  assign n60233 = pi546 & ~n47968;
  assign n60234 = pi246 & n47968;
  assign n60235 = ~n60233 & ~n60234;
  assign n60236 = pi547 & ~n47968;
  assign n60237 = pi247 & n47968;
  assign n60238 = ~n60236 & ~n60237;
  assign n60239 = pi548 & ~n47968;
  assign n60240 = pi248 & n47968;
  assign n60241 = ~n60239 & ~n60240;
  assign n60242 = pi549 & ~n47975;
  assign n60243 = pi235 & n47975;
  assign n60244 = ~n60242 & ~n60243;
  assign n60245 = pi550 & ~n47975;
  assign n60246 = ~pi239 & n47975;
  assign po707 = ~n60245 & ~n60246;
  assign n60248 = pi551 & ~n47975;
  assign n60249 = pi240 & n47975;
  assign n60250 = ~n60248 & ~n60249;
  assign n60251 = pi552 & ~n47975;
  assign n60252 = pi247 & n47975;
  assign n60253 = ~n60251 & ~n60252;
  assign n60254 = pi553 & ~n47975;
  assign n60255 = pi241 & n47975;
  assign n60256 = ~n60254 & ~n60255;
  assign n60257 = pi554 & ~n47975;
  assign n60258 = pi248 & n47975;
  assign n60259 = ~n60257 & ~n60258;
  assign n60260 = pi555 & ~n47975;
  assign n60261 = pi249 & n47975;
  assign n60262 = ~n60260 & ~n60261;
  assign n60263 = pi556 & ~n47832;
  assign n60264 = pi242 & n47832;
  assign n60265 = ~n60263 & ~n60264;
  assign n60266 = pi557 & ~n47953;
  assign n60267 = n47579 & n58591;
  assign n60268 = n47953 & n58593;
  assign n60269 = pi557 & ~n60268;
  assign n60270 = ~pi557 & n47579;
  assign n60271 = n58591 & n60270;
  assign n60272 = ~n60269 & ~n60271;
  assign n60273 = ~n60266 & ~n60267;
  assign n60274 = pi558 & ~n47953;
  assign n60275 = pi244 & n47953;
  assign n60276 = ~n60274 & ~n60275;
  assign n60277 = pi559 & ~n47816;
  assign n60278 = pi241 & n47816;
  assign n60279 = ~n60277 & ~n60278;
  assign n60280 = pi560 & ~n47832;
  assign n60281 = pi240 & n47832;
  assign n60282 = ~n60280 & ~n60281;
  assign n60283 = pi561 & ~n47824;
  assign n60284 = pi247 & n47824;
  assign n60285 = ~n60283 & ~n60284;
  assign n60286 = pi562 & ~n47832;
  assign n60287 = pi241 & n47832;
  assign n60288 = ~n60286 & ~n60287;
  assign n60289 = pi563 & ~n47975;
  assign n60290 = pi246 & n47975;
  assign n60291 = ~n60289 & ~n60290;
  assign n60292 = pi564 & ~n47832;
  assign n60293 = pi246 & n47832;
  assign n60294 = ~n60292 & ~n60293;
  assign n60295 = pi565 & ~n47832;
  assign n60296 = pi248 & n47832;
  assign n60297 = ~n60295 & ~n60296;
  assign n60298 = pi566 & ~n47832;
  assign n60299 = pi244 & n47832;
  assign n60300 = ~n60298 & ~n60299;
  assign n60301 = pi568 & ~n47832;
  assign n60302 = pi245 & n47832;
  assign n60303 = ~n60301 & ~n60302;
  assign n60304 = pi569 & ~n47832;
  assign n60305 = ~pi239 & n47832;
  assign po726 = ~n60304 & ~n60305;
  assign n60307 = pi570 & ~n47832;
  assign n60308 = n47827 & n58638;
  assign n60309 = n47832 & n58615;
  assign n60310 = pi570 & ~n60309;
  assign n60311 = ~pi570 & n47827;
  assign n60312 = n58638 & n60311;
  assign n60313 = ~n60310 & ~n60312;
  assign n60314 = ~n60307 & ~n60308;
  assign n60315 = pi571 & ~n47982;
  assign n60316 = pi241 & n47982;
  assign n60317 = ~n60315 & ~n60316;
  assign n60318 = pi572 & ~n47982;
  assign n60319 = pi244 & n47982;
  assign n60320 = ~n60318 & ~n60319;
  assign n60321 = pi573 & ~n47982;
  assign n60322 = pi242 & n47982;
  assign n60323 = ~n60321 & ~n60322;
  assign n60324 = pi574 & ~n47824;
  assign n60325 = pi241 & n47824;
  assign n60326 = ~n60324 & ~n60325;
  assign n60327 = pi575 & ~n47982;
  assign n60328 = pi235 & n47982;
  assign n60329 = ~n60327 & ~n60328;
  assign n60330 = pi576 & ~n47982;
  assign n60331 = pi248 & n47982;
  assign n60332 = ~n60330 & ~n60331;
  assign n60333 = pi577 & ~n47975;
  assign n60334 = pi238 & n47975;
  assign n60335 = ~n60333 & ~n60334;
  assign n60336 = pi578 & ~n47824;
  assign n60337 = pi249 & n47824;
  assign n60338 = ~n60336 & ~n60337;
  assign n60339 = pi579 & ~n47816;
  assign n60340 = pi249 & n47816;
  assign n60341 = ~n60339 & ~n60340;
  assign n60342 = pi580 & ~n47975;
  assign n60343 = pi245 & n47975;
  assign n60344 = ~n60342 & ~n60343;
  assign n60345 = pi581 & ~n47824;
  assign n60346 = pi235 & n47824;
  assign n60347 = ~n60345 & ~n60346;
  assign n60348 = pi582 & ~n47824;
  assign n60349 = pi240 & n47824;
  assign n60350 = ~n60348 & ~n60349;
  assign n60351 = pi584 & ~n47824;
  assign n60352 = pi245 & n47824;
  assign n60353 = ~n60351 & ~n60352;
  assign n60354 = pi585 & ~n47824;
  assign n60355 = pi244 & n47824;
  assign n60356 = ~n60354 & ~n60355;
  assign n60357 = pi586 & ~n47824;
  assign n60358 = pi242 & n47824;
  assign n60359 = ~n60357 & ~n60358;
  assign n60360 = ~pi882 & n62455;
  assign n60361 = pi947 & n60360;
  assign n60362 = pi598 & ~n60361;
  assign n60363 = pi740 & pi780;
  assign n60364 = n2904 & n60363;
  assign n60365 = ~n60362 & ~n60364;
  assign n60366 = pi907 & n60360;
  assign n60367 = ~pi615 & ~n60366;
  assign n60368 = pi779 & pi797;
  assign n60369 = n2907 & n60368;
  assign n60370 = ~n60367 & ~n60369;
  assign n60371 = pi832 & ~pi973;
  assign n60372 = ~pi1054 & pi1066;
  assign n60373 = pi1088 & n60372;
  assign n60374 = n60371 & n60373;
  assign po954 = ~pi953 & n60374;
  assign n60376 = ~pi1116 & po954;
  assign n60377 = ~pi625 & ~po954;
  assign n60378 = ~pi962 & ~n60377;
  assign n60379 = ~pi962 & ~n60376;
  assign n60380 = ~n60377 & n60379;
  assign n60381 = ~n60376 & n60378;
  assign n60382 = ~pi1117 & po954;
  assign n60383 = ~pi627 & ~po954;
  assign n60384 = ~pi962 & ~n60383;
  assign n60385 = ~pi962 & ~n60382;
  assign n60386 = ~n60383 & n60385;
  assign n60387 = ~n60382 & n60384;
  assign n60388 = ~pi1119 & po954;
  assign n60389 = ~pi628 & ~po954;
  assign n60390 = ~pi962 & ~n60389;
  assign n60391 = ~pi962 & ~n60388;
  assign n60392 = ~n60389 & n60391;
  assign n60393 = ~n60388 & n60390;
  assign n60394 = ~pi980 & pi1038;
  assign n60395 = pi1060 & n60394;
  assign n60396 = pi832 & ~pi1061;
  assign n60397 = pi952 & n60396;
  assign n60398 = pi952 & ~pi1061;
  assign n60399 = n60395 & n60398;
  assign n60400 = pi832 & n60399;
  assign n60401 = n60395 & n60397;
  assign n60402 = ~pi1119 & po897;
  assign n60403 = ~pi629 & ~po897;
  assign n60404 = ~pi966 & ~n60403;
  assign n60405 = ~pi966 & ~n60402;
  assign n60406 = ~n60403 & n60405;
  assign n60407 = ~n60402 & n60404;
  assign n60408 = ~pi1120 & po897;
  assign n60409 = ~pi630 & ~po897;
  assign n60410 = ~pi966 & ~n60409;
  assign n60411 = ~pi966 & ~n60408;
  assign n60412 = ~n60409 & n60411;
  assign n60413 = ~n60408 & n60410;
  assign n60414 = pi631 & ~po954;
  assign n60415 = ~pi1113 & po954;
  assign n60416 = ~pi962 & ~n60415;
  assign n60417 = ~pi962 & ~n60414;
  assign n60418 = ~n60415 & n60417;
  assign n60419 = ~n60414 & n60416;
  assign n60420 = pi632 & ~po954;
  assign n60421 = ~pi1115 & po954;
  assign n60422 = ~pi962 & ~n60421;
  assign n60423 = ~pi962 & ~n60420;
  assign n60424 = ~n60421 & n60423;
  assign n60425 = ~n60420 & n60422;
  assign n60426 = ~pi1110 & po897;
  assign n60427 = ~pi633 & ~po897;
  assign n60428 = ~pi966 & ~n60427;
  assign n60429 = ~pi966 & ~n60426;
  assign n60430 = ~n60427 & n60429;
  assign n60431 = ~n60426 & n60428;
  assign n60432 = ~pi1110 & po954;
  assign n60433 = ~pi634 & ~po954;
  assign n60434 = ~pi962 & ~n60433;
  assign n60435 = ~pi962 & ~n60432;
  assign n60436 = ~n60433 & n60435;
  assign n60437 = ~n60432 & n60434;
  assign n60438 = pi635 & ~po954;
  assign n60439 = ~pi1112 & po954;
  assign n60440 = ~pi962 & ~n60439;
  assign n60441 = ~pi962 & ~n60438;
  assign n60442 = ~n60439 & n60441;
  assign n60443 = ~n60438 & n60440;
  assign n60444 = ~pi1127 & po897;
  assign n60445 = ~pi636 & ~po897;
  assign n60446 = ~pi966 & ~n60445;
  assign n60447 = ~pi966 & ~n60444;
  assign n60448 = ~n60445 & n60447;
  assign n60449 = ~n60444 & n60446;
  assign n60450 = ~pi1105 & po954;
  assign n60451 = ~pi637 & ~po954;
  assign n60452 = ~pi962 & ~n60451;
  assign n60453 = ~pi962 & ~n60450;
  assign n60454 = ~n60451 & n60453;
  assign n60455 = ~n60450 & n60452;
  assign n60456 = ~pi1107 & po954;
  assign n60457 = ~pi638 & ~po954;
  assign n60458 = ~pi962 & ~n60457;
  assign n60459 = ~pi962 & ~n60456;
  assign n60460 = ~n60457 & n60459;
  assign n60461 = ~n60456 & n60458;
  assign n60462 = ~pi1109 & po954;
  assign n60463 = ~pi639 & ~po954;
  assign n60464 = ~pi962 & ~n60463;
  assign n60465 = ~pi962 & ~n60462;
  assign n60466 = ~n60463 & n60465;
  assign n60467 = ~n60462 & n60464;
  assign n60468 = ~pi1128 & po897;
  assign n60469 = ~pi640 & ~po897;
  assign n60470 = ~pi966 & ~n60469;
  assign n60471 = ~pi966 & ~n60468;
  assign n60472 = ~n60469 & n60471;
  assign n60473 = ~n60468 & n60470;
  assign n60474 = ~pi1121 & po954;
  assign n60475 = ~pi641 & ~po954;
  assign n60476 = ~pi962 & ~n60475;
  assign n60477 = ~pi962 & ~n60474;
  assign n60478 = ~n60475 & n60477;
  assign n60479 = ~n60474 & n60476;
  assign n60480 = ~pi1104 & po954;
  assign n60481 = ~pi643 & ~po954;
  assign n60482 = ~pi962 & ~n60481;
  assign n60483 = ~pi962 & ~n60480;
  assign n60484 = ~n60481 & n60483;
  assign n60485 = ~n60480 & n60482;
  assign n60486 = ~pi1123 & po897;
  assign n60487 = ~pi644 & ~po897;
  assign n60488 = ~pi966 & ~n60487;
  assign n60489 = ~pi966 & ~n60486;
  assign n60490 = ~n60487 & n60489;
  assign n60491 = ~n60486 & n60488;
  assign n60492 = ~pi1125 & po897;
  assign n60493 = ~pi645 & ~po897;
  assign n60494 = ~pi966 & ~n60493;
  assign n60495 = ~pi966 & ~n60492;
  assign n60496 = ~n60493 & n60495;
  assign n60497 = ~n60492 & n60494;
  assign n60498 = pi646 & ~po954;
  assign n60499 = ~pi1114 & po954;
  assign n60500 = ~pi962 & ~n60499;
  assign n60501 = ~pi962 & ~n60498;
  assign n60502 = ~n60499 & n60501;
  assign n60503 = ~n60498 & n60500;
  assign n60504 = ~pi1120 & po954;
  assign n60505 = ~pi647 & ~po954;
  assign n60506 = ~pi962 & ~n60505;
  assign n60507 = ~pi962 & ~n60504;
  assign n60508 = ~n60505 & n60507;
  assign n60509 = ~n60504 & n60506;
  assign n60510 = ~pi1122 & po954;
  assign n60511 = ~pi648 & ~po954;
  assign n60512 = ~pi962 & ~n60511;
  assign n60513 = ~pi962 & ~n60510;
  assign n60514 = ~n60511 & n60513;
  assign n60515 = ~n60510 & n60512;
  assign n60516 = pi649 & ~po954;
  assign n60517 = ~pi1126 & po954;
  assign n60518 = ~pi962 & ~n60517;
  assign n60519 = ~pi962 & ~n60516;
  assign n60520 = ~n60517 & n60519;
  assign n60521 = ~n60516 & n60518;
  assign n60522 = pi650 & ~po954;
  assign n60523 = ~pi1127 & po954;
  assign n60524 = ~pi962 & ~n60523;
  assign n60525 = ~pi962 & ~n60522;
  assign n60526 = ~n60523 & n60525;
  assign n60527 = ~n60522 & n60524;
  assign n60528 = ~pi1130 & po897;
  assign n60529 = ~pi651 & ~po897;
  assign n60530 = ~pi966 & ~n60529;
  assign n60531 = ~pi966 & ~n60528;
  assign n60532 = ~n60529 & n60531;
  assign n60533 = ~n60528 & n60530;
  assign n60534 = ~pi1131 & po897;
  assign n60535 = ~pi652 & ~po897;
  assign n60536 = ~pi966 & ~n60535;
  assign n60537 = ~pi966 & ~n60534;
  assign n60538 = ~n60535 & n60537;
  assign n60539 = ~n60534 & n60536;
  assign n60540 = ~pi1129 & po897;
  assign n60541 = ~pi653 & ~po897;
  assign n60542 = ~pi966 & ~n60541;
  assign n60543 = ~pi966 & ~n60540;
  assign n60544 = ~n60541 & n60543;
  assign n60545 = ~n60540 & n60542;
  assign n60546 = pi654 & ~po954;
  assign n60547 = ~pi1130 & po954;
  assign n60548 = ~pi962 & ~n60547;
  assign n60549 = ~pi962 & ~n60546;
  assign n60550 = ~n60547 & n60549;
  assign n60551 = ~n60546 & n60548;
  assign n60552 = pi655 & ~po954;
  assign n60553 = ~pi1124 & po954;
  assign n60554 = ~pi962 & ~n60553;
  assign n60555 = ~pi962 & ~n60552;
  assign n60556 = ~n60553 & n60555;
  assign n60557 = ~n60552 & n60554;
  assign n60558 = ~pi1126 & po897;
  assign n60559 = ~pi656 & ~po897;
  assign n60560 = ~pi966 & ~n60559;
  assign n60561 = ~pi966 & ~n60558;
  assign n60562 = ~n60559 & n60561;
  assign n60563 = ~n60558 & n60560;
  assign n60564 = pi657 & ~po954;
  assign n60565 = ~pi1131 & po954;
  assign n60566 = ~pi962 & ~n60565;
  assign n60567 = ~pi962 & ~n60564;
  assign n60568 = ~n60565 & n60567;
  assign n60569 = ~n60564 & n60566;
  assign n60570 = ~pi1124 & po897;
  assign n60571 = ~pi658 & ~po897;
  assign n60572 = ~pi966 & ~n60571;
  assign n60573 = ~pi966 & ~n60570;
  assign n60574 = ~n60571 & n60573;
  assign n60575 = ~n60570 & n60572;
  assign n60576 = ~pi1118 & po954;
  assign n60577 = ~pi660 & ~po954;
  assign n60578 = ~pi962 & ~n60577;
  assign n60579 = ~pi962 & ~n60576;
  assign n60580 = ~n60577 & n60579;
  assign n60581 = ~n60576 & n60578;
  assign n60582 = ~pi1101 & po954;
  assign n60583 = ~pi661 & ~po954;
  assign n60584 = ~pi962 & ~n60583;
  assign n60585 = ~pi962 & ~n60582;
  assign n60586 = ~n60583 & n60585;
  assign n60587 = ~n60582 & n60584;
  assign n60588 = ~pi1102 & po954;
  assign n60589 = ~pi662 & ~po954;
  assign n60590 = ~pi962 & ~n60589;
  assign n60591 = ~pi962 & ~n60588;
  assign n60592 = ~n60589 & n60591;
  assign n60593 = ~n60588 & n60590;
  assign n60594 = ~pi1108 & po954;
  assign n60595 = ~pi665 & ~po954;
  assign n60596 = ~pi962 & ~n60595;
  assign n60597 = ~pi962 & ~n60594;
  assign n60598 = ~n60595 & n60597;
  assign n60599 = ~n60594 & n60596;
  assign n60600 = pi669 & ~po954;
  assign n60601 = ~pi1125 & po954;
  assign n60602 = ~pi962 & ~n60601;
  assign n60603 = ~pi962 & ~n60600;
  assign n60604 = ~n60601 & n60603;
  assign n60605 = ~n60600 & n60602;
  assign n60606 = ~pi1100 & po954;
  assign n60607 = ~pi680 & ~po954;
  assign n60608 = ~pi962 & ~n60607;
  assign n60609 = ~pi962 & ~n60606;
  assign n60610 = ~n60607 & n60609;
  assign n60611 = ~n60606 & n60608;
  assign n60612 = ~pi1103 & po954;
  assign n60613 = ~pi681 & ~po954;
  assign n60614 = ~pi962 & ~n60613;
  assign n60615 = ~pi962 & ~n60612;
  assign n60616 = ~n60613 & n60615;
  assign n60617 = ~n60612 & n60614;
  assign po980 = pi953 & n60374;
  assign n60619 = pi684 & ~po980;
  assign n60620 = ~pi1130 & po980;
  assign n60621 = ~pi962 & ~n60620;
  assign n60622 = ~pi962 & ~n60619;
  assign n60623 = ~n60620 & n60622;
  assign n60624 = ~n60619 & n60621;
  assign n60625 = pi686 & ~po980;
  assign n60626 = ~pi1113 & po980;
  assign n60627 = ~pi962 & ~n60626;
  assign n60628 = ~pi962 & ~n60625;
  assign n60629 = ~n60626 & n60628;
  assign n60630 = ~n60625 & n60627;
  assign n60631 = ~pi1127 & po980;
  assign n60632 = ~pi687 & ~po980;
  assign n60633 = ~pi962 & ~n60632;
  assign n60634 = ~pi962 & ~n60631;
  assign n60635 = ~n60632 & n60634;
  assign n60636 = ~n60631 & n60633;
  assign n60637 = pi688 & ~po980;
  assign n60638 = ~pi1115 & po980;
  assign n60639 = ~pi962 & ~n60638;
  assign n60640 = ~pi962 & ~n60637;
  assign n60641 = ~n60638 & n60640;
  assign n60642 = ~n60637 & n60639;
  assign n60643 = ~pi1108 & po980;
  assign n60644 = ~pi690 & ~po980;
  assign n60645 = ~pi962 & ~n60644;
  assign n60646 = ~pi962 & ~n60643;
  assign n60647 = ~n60644 & n60646;
  assign n60648 = ~n60643 & n60645;
  assign n60649 = ~pi1107 & po980;
  assign n60650 = ~pi691 & ~po980;
  assign n60651 = ~pi962 & ~n60650;
  assign n60652 = ~pi962 & ~n60649;
  assign n60653 = ~n60650 & n60652;
  assign n60654 = ~n60649 & n60651;
  assign n60655 = pi693 & ~po954;
  assign n60656 = ~pi1129 & po954;
  assign n60657 = ~pi962 & ~n60656;
  assign n60658 = ~pi962 & ~n60655;
  assign n60659 = ~n60656 & n60658;
  assign n60660 = ~n60655 & n60657;
  assign n60661 = pi694 & ~po980;
  assign n60662 = ~pi1128 & po980;
  assign n60663 = ~pi962 & ~n60662;
  assign n60664 = ~pi962 & ~n60661;
  assign n60665 = ~n60662 & n60664;
  assign n60666 = ~n60661 & n60663;
  assign n60667 = pi695 & ~po954;
  assign n60668 = ~pi1111 & po954;
  assign n60669 = ~pi962 & ~n60668;
  assign n60670 = ~pi962 & ~n60667;
  assign n60671 = ~n60668 & n60670;
  assign n60672 = ~n60667 & n60669;
  assign n60673 = ~pi1100 & po980;
  assign n60674 = ~pi696 & ~po980;
  assign n60675 = ~pi962 & ~n60674;
  assign n60676 = ~pi962 & ~n60673;
  assign n60677 = ~n60674 & n60676;
  assign n60678 = ~n60673 & n60675;
  assign n60679 = pi697 & ~po980;
  assign n60680 = ~pi1129 & po980;
  assign n60681 = ~pi962 & ~n60680;
  assign n60682 = ~pi962 & ~n60679;
  assign n60683 = ~n60680 & n60682;
  assign n60684 = ~n60679 & n60681;
  assign n60685 = pi698 & ~po980;
  assign n60686 = ~pi1116 & po980;
  assign n60687 = ~pi962 & ~n60686;
  assign n60688 = ~pi962 & ~n60685;
  assign n60689 = ~n60686 & n60688;
  assign n60690 = ~n60685 & n60687;
  assign n60691 = ~pi1103 & po980;
  assign n60692 = ~pi699 & ~po980;
  assign n60693 = ~pi962 & ~n60692;
  assign n60694 = ~pi962 & ~n60691;
  assign n60695 = ~n60692 & n60694;
  assign n60696 = ~n60691 & n60693;
  assign n60697 = ~pi1110 & po980;
  assign n60698 = ~pi700 & ~po980;
  assign n60699 = ~pi962 & ~n60698;
  assign n60700 = ~pi962 & ~n60697;
  assign n60701 = ~n60698 & n60700;
  assign n60702 = ~n60697 & n60699;
  assign n60703 = pi701 & ~po980;
  assign n60704 = ~pi1123 & po980;
  assign n60705 = ~pi962 & ~n60704;
  assign n60706 = ~pi962 & ~n60703;
  assign n60707 = ~n60704 & n60706;
  assign n60708 = ~n60703 & n60705;
  assign n60709 = pi702 & ~po980;
  assign n60710 = ~pi1117 & po980;
  assign n60711 = ~pi962 & ~n60710;
  assign n60712 = ~pi962 & ~n60709;
  assign n60713 = ~n60710 & n60712;
  assign n60714 = ~n60709 & n60711;
  assign n60715 = ~pi1124 & po980;
  assign n60716 = ~pi703 & ~po980;
  assign n60717 = ~pi962 & ~n60716;
  assign n60718 = ~pi962 & ~n60715;
  assign n60719 = ~n60716 & n60718;
  assign n60720 = ~n60715 & n60717;
  assign n60721 = pi704 & ~po980;
  assign n60722 = ~pi1112 & po980;
  assign n60723 = ~pi962 & ~n60722;
  assign n60724 = ~pi962 & ~n60721;
  assign n60725 = ~n60722 & n60724;
  assign n60726 = ~n60721 & n60723;
  assign n60727 = ~pi1125 & po980;
  assign n60728 = ~pi705 & ~po980;
  assign n60729 = ~pi962 & ~n60728;
  assign n60730 = ~pi962 & ~n60727;
  assign n60731 = ~n60728 & n60730;
  assign n60732 = ~n60727 & n60729;
  assign n60733 = ~pi1105 & po980;
  assign n60734 = ~pi706 & ~po980;
  assign n60735 = ~pi962 & ~n60734;
  assign n60736 = ~pi962 & ~n60733;
  assign n60737 = ~n60734 & n60736;
  assign n60738 = ~n60733 & n60735;
  assign n60739 = pi709 & ~po980;
  assign n60740 = ~pi1118 & po980;
  assign n60741 = ~pi962 & ~n60740;
  assign n60742 = ~pi962 & ~n60739;
  assign n60743 = ~n60740 & n60742;
  assign n60744 = ~n60739 & n60741;
  assign n60745 = ~pi1106 & po954;
  assign n60746 = ~pi710 & ~po954;
  assign n60747 = ~pi962 & ~n60746;
  assign n60748 = ~pi962 & ~n60745;
  assign n60749 = ~n60746 & n60748;
  assign n60750 = ~n60745 & n60747;
  assign n60751 = ~pi1123 & po954;
  assign n60752 = ~pi715 & ~po954;
  assign n60753 = ~pi962 & ~n60752;
  assign n60754 = ~pi962 & ~n60751;
  assign n60755 = ~n60752 & n60754;
  assign n60756 = ~n60751 & n60753;
  assign n60757 = pi723 & ~po980;
  assign n60758 = ~pi1111 & po980;
  assign n60759 = ~pi962 & ~n60758;
  assign n60760 = ~pi962 & ~n60757;
  assign n60761 = ~n60758 & n60760;
  assign n60762 = ~n60757 & n60759;
  assign n60763 = pi724 & ~po980;
  assign n60764 = ~pi1114 & po980;
  assign n60765 = ~pi962 & ~n60764;
  assign n60766 = ~pi962 & ~n60763;
  assign n60767 = ~n60764 & n60766;
  assign n60768 = ~n60763 & n60765;
  assign n60769 = pi725 & ~po980;
  assign n60770 = ~pi1120 & po980;
  assign n60771 = ~pi962 & ~n60770;
  assign n60772 = ~pi962 & ~n60769;
  assign n60773 = ~n60770 & n60772;
  assign n60774 = ~n60769 & n60771;
  assign n60775 = ~pi1126 & po980;
  assign n60776 = ~pi726 & ~po980;
  assign n60777 = ~pi962 & ~n60776;
  assign n60778 = ~pi962 & ~n60775;
  assign n60779 = ~n60776 & n60778;
  assign n60780 = ~n60775 & n60777;
  assign n60781 = ~pi1102 & po980;
  assign n60782 = ~pi727 & ~po980;
  assign n60783 = ~pi962 & ~n60782;
  assign n60784 = ~pi962 & ~n60781;
  assign n60785 = ~n60782 & n60784;
  assign n60786 = ~n60781 & n60783;
  assign n60787 = pi728 & ~po980;
  assign n60788 = ~pi1131 & po980;
  assign n60789 = ~pi962 & ~n60788;
  assign n60790 = ~pi962 & ~n60787;
  assign n60791 = ~n60788 & n60790;
  assign n60792 = ~n60787 & n60789;
  assign n60793 = ~pi1104 & po980;
  assign n60794 = ~pi729 & ~po980;
  assign n60795 = ~pi962 & ~n60794;
  assign n60796 = ~pi962 & ~n60793;
  assign n60797 = ~n60794 & n60796;
  assign n60798 = ~n60793 & n60795;
  assign n60799 = ~pi1106 & po980;
  assign n60800 = ~pi730 & ~po980;
  assign n60801 = ~pi962 & ~n60800;
  assign n60802 = ~pi962 & ~n60799;
  assign n60803 = ~n60800 & n60802;
  assign n60804 = ~n60799 & n60801;
  assign n60805 = pi732 & ~po954;
  assign n60806 = ~pi1128 & po954;
  assign n60807 = ~pi962 & ~n60806;
  assign n60808 = ~pi962 & ~n60805;
  assign n60809 = ~n60806 & n60808;
  assign n60810 = ~n60805 & n60807;
  assign n60811 = pi734 & ~po980;
  assign n60812 = ~pi1119 & po980;
  assign n60813 = ~pi962 & ~n60812;
  assign n60814 = ~pi962 & ~n60811;
  assign n60815 = ~n60812 & n60814;
  assign n60816 = ~n60811 & n60813;
  assign n60817 = ~pi1109 & po980;
  assign n60818 = ~pi735 & ~po980;
  assign n60819 = ~pi962 & ~n60818;
  assign n60820 = ~pi962 & ~n60817;
  assign n60821 = ~n60818 & n60820;
  assign n60822 = ~n60817 & n60819;
  assign n60823 = ~pi1101 & po980;
  assign n60824 = ~pi736 & ~po980;
  assign n60825 = ~pi962 & ~n60824;
  assign n60826 = ~pi962 & ~n60823;
  assign n60827 = ~n60824 & n60826;
  assign n60828 = ~n60823 & n60825;
  assign n60829 = pi737 & ~po980;
  assign n60830 = ~pi1122 & po980;
  assign n60831 = ~pi962 & ~n60830;
  assign n60832 = ~pi962 & ~n60829;
  assign n60833 = ~n60830 & n60832;
  assign n60834 = ~n60829 & n60831;
  assign n60835 = pi738 & ~po980;
  assign n60836 = ~pi1121 & po980;
  assign n60837 = ~pi962 & ~n60836;
  assign n60838 = ~pi962 & ~n60835;
  assign n60839 = ~n60836 & n60838;
  assign n60840 = ~n60835 & n60837;
  assign n60841 = ~pi952 & n60396;
  assign n60842 = ~pi952 & ~pi1061;
  assign n60843 = n60395 & n60842;
  assign n60844 = pi832 & n60843;
  assign n60845 = n60395 & n60841;
  assign n60846 = pi739 & ~po988;
  assign n60847 = pi1108 & po988;
  assign n60848 = ~pi966 & ~n60847;
  assign n60849 = ~pi966 & ~n60846;
  assign n60850 = ~n60847 & n60849;
  assign n60851 = ~n60846 & n60848;
  assign n60852 = pi1114 & po988;
  assign n60853 = ~pi741 & ~po988;
  assign n60854 = ~pi966 & ~n60853;
  assign n60855 = ~pi966 & ~n60852;
  assign n60856 = ~n60853 & n60855;
  assign n60857 = ~n60852 & n60854;
  assign n60858 = pi1112 & po988;
  assign n60859 = ~pi742 & ~po988;
  assign n60860 = ~pi966 & ~n60859;
  assign n60861 = ~pi966 & ~n60858;
  assign n60862 = ~n60859 & n60861;
  assign n60863 = ~n60858 & n60860;
  assign n60864 = pi743 & ~po988;
  assign n60865 = pi1109 & po988;
  assign n60866 = ~pi966 & ~n60865;
  assign n60867 = ~pi966 & ~n60864;
  assign n60868 = ~n60865 & n60867;
  assign n60869 = ~n60864 & n60866;
  assign n60870 = pi1131 & po988;
  assign n60871 = ~pi744 & ~po988;
  assign n60872 = ~pi966 & ~n60871;
  assign n60873 = ~pi966 & ~n60870;
  assign n60874 = ~n60871 & n60873;
  assign n60875 = ~n60870 & n60872;
  assign n60876 = pi1111 & po988;
  assign n60877 = ~pi745 & ~po988;
  assign n60878 = ~pi966 & ~n60877;
  assign n60879 = ~pi966 & ~n60876;
  assign n60880 = ~n60877 & n60879;
  assign n60881 = ~n60876 & n60878;
  assign n60882 = pi746 & ~po988;
  assign n60883 = pi1104 & po988;
  assign n60884 = ~pi966 & ~n60883;
  assign n60885 = ~pi966 & ~n60882;
  assign n60886 = ~n60883 & n60885;
  assign n60887 = ~n60882 & n60884;
  assign n60888 = pi748 & ~po988;
  assign n60889 = pi1106 & po988;
  assign n60890 = ~pi966 & ~n60889;
  assign n60891 = ~pi966 & ~n60888;
  assign n60892 = ~n60889 & n60891;
  assign n60893 = ~n60888 & n60890;
  assign n60894 = pi749 & ~po988;
  assign n60895 = pi1105 & po988;
  assign n60896 = ~pi966 & ~n60895;
  assign n60897 = ~pi966 & ~n60894;
  assign n60898 = ~n60895 & n60897;
  assign n60899 = ~n60894 & n60896;
  assign n60900 = pi1130 & po988;
  assign n60901 = ~pi750 & ~po988;
  assign n60902 = ~pi966 & ~n60901;
  assign n60903 = ~pi966 & ~n60900;
  assign n60904 = ~n60901 & n60903;
  assign n60905 = ~n60900 & n60902;
  assign n60906 = pi1123 & po988;
  assign n60907 = ~pi751 & ~po988;
  assign n60908 = ~pi966 & ~n60907;
  assign n60909 = ~pi966 & ~n60906;
  assign n60910 = ~n60907 & n60909;
  assign n60911 = ~n60906 & n60908;
  assign n60912 = pi1124 & po988;
  assign n60913 = ~pi752 & ~po988;
  assign n60914 = ~pi966 & ~n60913;
  assign n60915 = ~pi966 & ~n60912;
  assign n60916 = ~n60913 & n60915;
  assign n60917 = ~n60912 & n60914;
  assign n60918 = pi123 & n38189;
  assign n60919 = pi1131 & ~n60918;
  assign n60920 = pi1127 & ~n60918;
  assign n60921 = ~n60919 & ~n60920;
  assign n60922 = ~pi825 & n60918;
  assign n60923 = n60921 & ~n60922;
  assign n60924 = pi1131 & n60920;
  assign n60925 = ~n60923 & ~n60924;
  assign n60926 = pi1128 & ~pi1129;
  assign n60927 = ~pi1128 & pi1129;
  assign n60928 = ~pi1128 & ~pi1129;
  assign n60929 = pi1128 & pi1129;
  assign n60930 = ~n60928 & ~n60929;
  assign n60931 = ~n60926 & ~n60927;
  assign n60932 = ~pi1125 & ~pi1126;
  assign n60933 = pi1125 & pi1126;
  assign n60934 = pi1125 & ~pi1126;
  assign n60935 = ~pi1125 & pi1126;
  assign n60936 = ~n60934 & ~n60935;
  assign n60937 = ~n60932 & ~n60933;
  assign n60938 = ~pi1124 & ~pi1130;
  assign n60939 = pi1124 & pi1130;
  assign n60940 = pi1124 & ~pi1130;
  assign n60941 = ~pi1124 & pi1130;
  assign n60942 = ~n60940 & ~n60941;
  assign n60943 = ~n60938 & ~n60939;
  assign n60944 = ~n65896 & n65897;
  assign n60945 = n65896 & ~n65897;
  assign n60946 = ~n60944 & ~n60945;
  assign n60947 = ~n65895 & n60946;
  assign n60948 = n65895 & ~n60946;
  assign n60949 = n65895 & n65897;
  assign n60950 = ~n65895 & ~n65897;
  assign n60951 = ~n60949 & ~n60950;
  assign n60952 = n65896 & n60951;
  assign n60953 = ~n65896 & ~n60951;
  assign n60954 = ~n60952 & ~n60953;
  assign n60955 = n65895 & n65896;
  assign n60956 = ~n65895 & ~n65896;
  assign n60957 = ~n60955 & ~n60956;
  assign n60958 = n65897 & n60957;
  assign n60959 = ~n65897 & ~n60957;
  assign n60960 = ~n60958 & ~n60959;
  assign n60961 = ~n60947 & ~n60948;
  assign n60962 = ~n60925 & ~n65898;
  assign n60963 = pi825 & n60918;
  assign n60964 = n60921 & ~n60963;
  assign n60965 = ~n60924 & n65898;
  assign n60966 = ~n60964 & n60965;
  assign po982 = ~n60962 & ~n60966;
  assign n60968 = pi1123 & ~n60918;
  assign n60969 = pi1122 & ~n60918;
  assign n60970 = ~n60968 & ~n60969;
  assign n60971 = ~pi826 & n60918;
  assign n60972 = n60970 & ~n60971;
  assign n60973 = pi1123 & n60969;
  assign n60974 = ~n60972 & ~n60973;
  assign n60975 = pi1120 & ~pi1121;
  assign n60976 = ~pi1120 & pi1121;
  assign n60977 = ~pi1120 & ~pi1121;
  assign n60978 = pi1120 & pi1121;
  assign n60979 = ~n60977 & ~n60978;
  assign n60980 = ~n60975 & ~n60976;
  assign n60981 = ~pi1116 & ~pi1117;
  assign n60982 = pi1116 & pi1117;
  assign n60983 = pi1116 & ~pi1117;
  assign n60984 = ~pi1116 & pi1117;
  assign n60985 = ~n60983 & ~n60984;
  assign n60986 = ~n60981 & ~n60982;
  assign n60987 = ~pi1118 & ~pi1119;
  assign n60988 = pi1118 & pi1119;
  assign n60989 = pi1118 & ~pi1119;
  assign n60990 = ~pi1118 & pi1119;
  assign n60991 = ~n60989 & ~n60990;
  assign n60992 = ~n60987 & ~n60988;
  assign n60993 = ~n65900 & n65901;
  assign n60994 = n65900 & ~n65901;
  assign n60995 = ~n60993 & ~n60994;
  assign n60996 = ~n65899 & n60995;
  assign n60997 = n65899 & ~n60995;
  assign n60998 = n65899 & n65901;
  assign n60999 = ~n65899 & ~n65901;
  assign n61000 = ~n60998 & ~n60999;
  assign n61001 = n65900 & n61000;
  assign n61002 = ~n65900 & ~n61000;
  assign n61003 = ~n61001 & ~n61002;
  assign n61004 = n65899 & n65900;
  assign n61005 = ~n65899 & ~n65900;
  assign n61006 = ~n61004 & ~n61005;
  assign n61007 = n65901 & n61006;
  assign n61008 = ~n65901 & ~n61006;
  assign n61009 = ~n61007 & ~n61008;
  assign n61010 = ~n60996 & ~n60997;
  assign n61011 = ~n60974 & ~n65902;
  assign n61012 = pi826 & n60918;
  assign n61013 = n60970 & ~n61012;
  assign n61014 = ~n60973 & n65902;
  assign n61015 = ~n61013 & n61014;
  assign po983 = ~n61011 & ~n61015;
  assign n61017 = pi1100 & ~n60918;
  assign n61018 = pi1107 & ~n60918;
  assign n61019 = ~n61017 & ~n61018;
  assign n61020 = ~pi827 & n60918;
  assign n61021 = n61019 & ~n61020;
  assign n61022 = pi1100 & n61018;
  assign n61023 = ~n61021 & ~n61022;
  assign n61024 = pi1101 & ~pi1102;
  assign n61025 = ~pi1101 & pi1102;
  assign n61026 = ~pi1101 & ~pi1102;
  assign n61027 = pi1101 & pi1102;
  assign n61028 = ~n61026 & ~n61027;
  assign n61029 = ~n61024 & ~n61025;
  assign n61030 = ~pi1104 & ~pi1106;
  assign n61031 = pi1104 & pi1106;
  assign n61032 = pi1104 & ~pi1106;
  assign n61033 = ~pi1104 & pi1106;
  assign n61034 = ~n61032 & ~n61033;
  assign n61035 = ~n61030 & ~n61031;
  assign n61036 = ~pi1103 & ~pi1105;
  assign n61037 = pi1103 & pi1105;
  assign n61038 = pi1103 & ~pi1105;
  assign n61039 = ~pi1103 & pi1105;
  assign n61040 = ~n61038 & ~n61039;
  assign n61041 = ~n61036 & ~n61037;
  assign n61042 = ~n65904 & n65905;
  assign n61043 = n65904 & ~n65905;
  assign n61044 = ~n61042 & ~n61043;
  assign n61045 = ~n65903 & n61044;
  assign n61046 = n65903 & ~n61044;
  assign n61047 = n65903 & n65905;
  assign n61048 = ~n65903 & ~n65905;
  assign n61049 = ~n61047 & ~n61048;
  assign n61050 = n65904 & n61049;
  assign n61051 = ~n65904 & ~n61049;
  assign n61052 = ~n61050 & ~n61051;
  assign n61053 = n65903 & n65904;
  assign n61054 = ~n65903 & ~n65904;
  assign n61055 = ~n61053 & ~n61054;
  assign n61056 = n65905 & n61055;
  assign n61057 = ~n65905 & ~n61055;
  assign n61058 = ~n61056 & ~n61057;
  assign n61059 = ~n61045 & ~n61046;
  assign n61060 = ~n61023 & ~n65906;
  assign n61061 = pi827 & n60918;
  assign n61062 = n61019 & ~n61061;
  assign n61063 = ~n61022 & n65906;
  assign n61064 = ~n61062 & n61063;
  assign po984 = ~n61060 & ~n61064;
  assign n61066 = pi1115 & ~n60918;
  assign n61067 = pi1114 & ~n60918;
  assign n61068 = ~n61066 & ~n61067;
  assign n61069 = ~pi828 & n60918;
  assign n61070 = n61068 & ~n61069;
  assign n61071 = pi1115 & n61067;
  assign n61072 = ~n61070 & ~n61071;
  assign n61073 = pi1112 & ~pi1113;
  assign n61074 = ~pi1112 & pi1113;
  assign n61075 = ~pi1112 & ~pi1113;
  assign n61076 = pi1112 & pi1113;
  assign n61077 = ~n61075 & ~n61076;
  assign n61078 = ~n61073 & ~n61074;
  assign n61079 = ~pi1108 & ~pi1109;
  assign n61080 = pi1108 & pi1109;
  assign n61081 = pi1108 & ~pi1109;
  assign n61082 = ~pi1108 & pi1109;
  assign n61083 = ~n61081 & ~n61082;
  assign n61084 = ~n61079 & ~n61080;
  assign n61085 = ~pi1110 & ~pi1111;
  assign n61086 = pi1110 & pi1111;
  assign n61087 = pi1110 & ~pi1111;
  assign n61088 = ~pi1110 & pi1111;
  assign n61089 = ~n61087 & ~n61088;
  assign n61090 = ~n61085 & ~n61086;
  assign n61091 = ~n65908 & n65909;
  assign n61092 = n65908 & ~n65909;
  assign n61093 = ~n61091 & ~n61092;
  assign n61094 = ~n65907 & n61093;
  assign n61095 = n65907 & ~n61093;
  assign n61096 = n65907 & n65909;
  assign n61097 = ~n65907 & ~n65909;
  assign n61098 = ~n61096 & ~n61097;
  assign n61099 = n65908 & n61098;
  assign n61100 = ~n65908 & ~n61098;
  assign n61101 = ~n61099 & ~n61100;
  assign n61102 = n65907 & n65908;
  assign n61103 = ~n65907 & ~n65908;
  assign n61104 = ~n61102 & ~n61103;
  assign n61105 = n65909 & n61104;
  assign n61106 = ~n65909 & ~n61104;
  assign n61107 = ~n61105 & ~n61106;
  assign n61108 = ~n61094 & ~n61095;
  assign n61109 = ~n61072 & ~n65910;
  assign n61110 = pi828 & n60918;
  assign n61111 = n61068 & ~n61110;
  assign n61112 = ~n61071 & n65910;
  assign n61113 = ~n61111 & n61112;
  assign po985 = ~n61109 & ~n61113;
  assign n61115 = pi832 & ~pi1100;
  assign n61116 = n60399 & n61115;
  assign n61117 = ~pi1100 & po897;
  assign n61118 = ~pi603 & ~po897;
  assign n61119 = ~pi966 & ~n61118;
  assign n61120 = ~pi966 & ~n65911;
  assign n61121 = ~n61118 & n61120;
  assign n61122 = ~n65911 & n61119;
  assign n61123 = pi871 & pi966;
  assign n61124 = pi872 & pi966;
  assign n61125 = ~n61123 & ~n61124;
  assign n61126 = ~n65912 & n61125;
  assign n61127 = ~pi606 & ~po897;
  assign n61128 = ~pi1104 & po897;
  assign n61129 = pi606 & ~po897;
  assign n61130 = pi1104 & po897;
  assign n61131 = ~n61129 & ~n61130;
  assign n61132 = ~n61127 & ~n61128;
  assign n61133 = ~pi966 & n65913;
  assign n61134 = ~pi837 & pi966;
  assign n61135 = ~pi966 & ~n65913;
  assign n61136 = pi837 & pi966;
  assign n61137 = ~n61135 & ~n61136;
  assign n61138 = ~n61133 & ~n61134;
  assign n61139 = ~pi1102 & po897;
  assign n61140 = ~pi614 & ~po897;
  assign n61141 = ~pi966 & ~n61140;
  assign n61142 = ~pi966 & ~n61139;
  assign n61143 = ~n61140 & n61142;
  assign n61144 = ~n61139 & n61141;
  assign n61145 = ~n61123 & ~n65915;
  assign n61146 = ~pi1101 & po897;
  assign n61147 = ~pi616 & ~po897;
  assign n61148 = ~pi966 & ~n61147;
  assign n61149 = ~pi966 & ~n61146;
  assign n61150 = ~n61147 & n61149;
  assign n61151 = ~n61146 & n61148;
  assign n61152 = ~n61124 & ~n65916;
  assign n61153 = ~pi617 & ~po897;
  assign n61154 = ~pi1105 & po897;
  assign n61155 = pi617 & ~po897;
  assign n61156 = pi1105 & po897;
  assign n61157 = ~n61155 & ~n61156;
  assign n61158 = ~n61153 & ~n61154;
  assign n61159 = ~pi966 & n65917;
  assign n61160 = ~pi850 & pi966;
  assign n61161 = ~pi966 & ~n65917;
  assign n61162 = pi850 & pi966;
  assign n61163 = ~n61161 & ~n61162;
  assign n61164 = ~n61159 & ~n61160;
  assign n61165 = ~pi299 & pi983;
  assign n61166 = ~n40054 & ~n61165;
  assign n61167 = ~n60360 & n61166;
  assign n61168 = pi823 & n7008;
  assign n61169 = ~pi779 & n61168;
  assign n61170 = pi907 & n61165;
  assign n61171 = pi604 & ~n61170;
  assign n61172 = ~n61168 & n61171;
  assign n61173 = ~n61169 & ~n61172;
  assign n61174 = ~pi1107 & po897;
  assign n61175 = ~pi607 & ~po897;
  assign n61176 = ~pi966 & ~n61175;
  assign n61177 = ~pi966 & ~n61174;
  assign n61178 = ~n61175 & n61177;
  assign n61179 = ~n61174 & n61176;
  assign n61180 = ~pi1116 & po897;
  assign n61181 = ~pi608 & ~po897;
  assign n61182 = ~pi966 & ~n61181;
  assign n61183 = ~pi966 & ~n61180;
  assign n61184 = ~n61181 & n61183;
  assign n61185 = ~n61180 & n61182;
  assign n61186 = ~pi1118 & po897;
  assign n61187 = ~pi609 & ~po897;
  assign n61188 = ~pi966 & ~n61187;
  assign n61189 = ~pi966 & ~n61186;
  assign n61190 = ~n61187 & n61189;
  assign n61191 = ~n61186 & n61188;
  assign n61192 = ~pi1113 & po897;
  assign n61193 = ~pi610 & ~po897;
  assign n61194 = ~pi966 & ~n61193;
  assign n61195 = ~pi966 & ~n61192;
  assign n61196 = ~n61193 & n61195;
  assign n61197 = ~n61192 & n61194;
  assign n61198 = ~pi1114 & po897;
  assign n61199 = ~pi611 & ~po897;
  assign n61200 = ~pi966 & ~n61199;
  assign n61201 = ~pi966 & ~n61198;
  assign n61202 = ~n61199 & n61201;
  assign n61203 = ~n61198 & n61200;
  assign n61204 = ~pi1111 & po897;
  assign n61205 = ~pi612 & ~po897;
  assign n61206 = ~pi966 & ~n61205;
  assign n61207 = ~pi966 & ~n61204;
  assign n61208 = ~n61205 & n61207;
  assign n61209 = ~n61204 & n61206;
  assign n61210 = ~pi1115 & po897;
  assign n61211 = ~pi613 & ~po897;
  assign n61212 = ~pi966 & ~n61211;
  assign n61213 = ~pi966 & ~n61210;
  assign n61214 = ~n61211 & n61213;
  assign n61215 = ~n61210 & n61212;
  assign n61216 = ~pi1117 & po897;
  assign n61217 = ~pi618 & ~po897;
  assign n61218 = ~pi966 & ~n61217;
  assign n61219 = ~pi966 & ~n61216;
  assign n61220 = ~n61217 & n61219;
  assign n61221 = ~n61216 & n61218;
  assign n61222 = ~pi1122 & po897;
  assign n61223 = ~pi619 & ~po897;
  assign n61224 = ~pi966 & ~n61223;
  assign n61225 = ~pi966 & ~n61222;
  assign n61226 = ~n61223 & n61225;
  assign n61227 = ~n61222 & n61224;
  assign n61228 = ~pi1112 & po897;
  assign n61229 = ~pi620 & ~po897;
  assign n61230 = ~pi966 & ~n61229;
  assign n61231 = ~pi966 & ~n61228;
  assign n61232 = ~n61229 & n61231;
  assign n61233 = ~n61228 & n61230;
  assign n61234 = ~pi1108 & po897;
  assign n61235 = ~pi621 & ~po897;
  assign n61236 = ~pi966 & ~n61235;
  assign n61237 = ~pi966 & ~n61234;
  assign n61238 = ~n61235 & n61237;
  assign n61239 = ~n61234 & n61236;
  assign n61240 = ~pi1109 & po897;
  assign n61241 = ~pi622 & ~po897;
  assign n61242 = ~pi966 & ~n61241;
  assign n61243 = ~pi966 & ~n61240;
  assign n61244 = ~n61241 & n61243;
  assign n61245 = ~n61240 & n61242;
  assign n61246 = ~pi1106 & po897;
  assign n61247 = ~pi623 & ~po897;
  assign n61248 = ~pi966 & ~n61247;
  assign n61249 = ~pi966 & ~n61246;
  assign n61250 = ~n61247 & n61249;
  assign n61251 = ~n61246 & n61248;
  assign n61252 = pi831 & n7186;
  assign n61253 = ~pi780 & n61252;
  assign n61254 = pi947 & n61165;
  assign n61255 = pi624 & ~n61254;
  assign n61256 = ~n61252 & n61255;
  assign n61257 = ~n61253 & ~n61256;
  assign n61258 = ~pi1121 & po897;
  assign n61259 = ~pi626 & ~po897;
  assign n61260 = ~pi966 & ~n61259;
  assign n61261 = ~pi966 & ~n61258;
  assign n61262 = ~n61259 & n61261;
  assign n61263 = ~n61258 & n61260;
  assign n61264 = ~pi1103 & po897;
  assign n61265 = ~pi642 & ~po897;
  assign n61266 = ~pi966 & ~n61265;
  assign n61267 = ~pi966 & ~n61264;
  assign n61268 = ~n61265 & n61267;
  assign n61269 = ~n61264 & n61266;
  assign n61270 = pi1117 & po988;
  assign n61271 = ~pi753 & ~po988;
  assign n61272 = ~pi966 & ~n61271;
  assign n61273 = ~pi966 & ~n61270;
  assign n61274 = ~n61271 & n61273;
  assign n61275 = ~n61270 & n61272;
  assign n61276 = pi1118 & po988;
  assign n61277 = ~pi754 & ~po988;
  assign n61278 = ~pi966 & ~n61277;
  assign n61279 = ~pi966 & ~n61276;
  assign n61280 = ~n61277 & n61279;
  assign n61281 = ~n61276 & n61278;
  assign n61282 = pi1120 & po988;
  assign n61283 = ~pi755 & ~po988;
  assign n61284 = ~pi966 & ~n61283;
  assign n61285 = ~pi966 & ~n61282;
  assign n61286 = ~n61283 & n61285;
  assign n61287 = ~n61282 & n61284;
  assign n61288 = pi1119 & po988;
  assign n61289 = ~pi756 & ~po988;
  assign n61290 = ~pi966 & ~n61289;
  assign n61291 = ~pi966 & ~n61288;
  assign n61292 = ~n61289 & n61291;
  assign n61293 = ~n61288 & n61290;
  assign n61294 = pi1113 & po988;
  assign n61295 = ~pi757 & ~po988;
  assign n61296 = ~pi966 & ~n61295;
  assign n61297 = ~pi966 & ~n61294;
  assign n61298 = ~n61295 & n61297;
  assign n61299 = ~n61294 & n61296;
  assign n61300 = pi758 & ~po988;
  assign n61301 = pi1101 & po988;
  assign n61302 = ~pi966 & ~n61301;
  assign n61303 = ~pi966 & ~n61300;
  assign n61304 = ~n61301 & n61303;
  assign n61305 = ~n61300 & n61302;
  assign n61306 = pi759 & ~po988;
  assign n61307 = pi1100 & po988;
  assign n61308 = ~pi966 & ~n61307;
  assign n61309 = ~pi759 & ~po988;
  assign n61310 = n60843 & n61115;
  assign n61311 = ~n61309 & ~n61310;
  assign n61312 = ~pi966 & ~n61311;
  assign n61313 = ~n61306 & n61308;
  assign n61314 = pi1115 & po988;
  assign n61315 = ~pi760 & ~po988;
  assign n61316 = ~pi966 & ~n61315;
  assign n61317 = ~pi966 & ~n61314;
  assign n61318 = ~n61315 & n61317;
  assign n61319 = ~n61314 & n61316;
  assign n61320 = pi1121 & po988;
  assign n61321 = ~pi761 & ~po988;
  assign n61322 = ~pi966 & ~n61321;
  assign n61323 = ~pi966 & ~n61320;
  assign n61324 = ~n61321 & n61323;
  assign n61325 = ~n61320 & n61322;
  assign n61326 = pi1129 & po988;
  assign n61327 = ~pi762 & ~po988;
  assign n61328 = ~pi966 & ~n61327;
  assign n61329 = ~pi966 & ~n61326;
  assign n61330 = ~n61327 & n61329;
  assign n61331 = ~n61326 & n61328;
  assign n61332 = pi763 & ~po988;
  assign n61333 = pi1103 & po988;
  assign n61334 = ~pi966 & ~n61333;
  assign n61335 = ~pi966 & ~n61332;
  assign n61336 = ~n61333 & n61335;
  assign n61337 = ~n61332 & n61334;
  assign n61338 = pi764 & ~po988;
  assign n61339 = pi1107 & po988;
  assign n61340 = ~pi966 & ~n61339;
  assign n61341 = ~pi966 & ~n61338;
  assign n61342 = ~n61339 & n61341;
  assign n61343 = ~n61338 & n61340;
  assign n61344 = pi766 & ~po988;
  assign n61345 = pi1110 & po988;
  assign n61346 = ~pi966 & ~n61345;
  assign n61347 = ~pi966 & ~n61344;
  assign n61348 = ~n61345 & n61347;
  assign n61349 = ~n61344 & n61346;
  assign n61350 = pi1116 & po988;
  assign n61351 = ~pi767 & ~po988;
  assign n61352 = ~pi966 & ~n61351;
  assign n61353 = ~pi966 & ~n61350;
  assign n61354 = ~n61351 & n61353;
  assign n61355 = ~n61350 & n61352;
  assign n61356 = pi1125 & po988;
  assign n61357 = ~pi768 & ~po988;
  assign n61358 = ~pi966 & ~n61357;
  assign n61359 = ~pi966 & ~n61356;
  assign n61360 = ~n61357 & n61359;
  assign n61361 = ~n61356 & n61358;
  assign n61362 = pi1126 & po988;
  assign n61363 = ~pi770 & ~po988;
  assign n61364 = ~pi966 & ~n61363;
  assign n61365 = ~pi966 & ~n61362;
  assign n61366 = ~n61363 & n61365;
  assign n61367 = ~n61362 & n61364;
  assign n61368 = pi772 & ~po988;
  assign n61369 = pi1102 & po988;
  assign n61370 = ~pi966 & ~n61369;
  assign n61371 = ~pi966 & ~n61368;
  assign n61372 = ~n61369 & n61371;
  assign n61373 = ~n61368 & n61370;
  assign n61374 = pi1127 & po988;
  assign n61375 = ~pi774 & ~po988;
  assign n61376 = ~pi966 & ~n61375;
  assign n61377 = ~pi966 & ~n61374;
  assign n61378 = ~n61375 & n61377;
  assign n61379 = ~n61374 & n61376;
  assign n61380 = pi1128 & po988;
  assign n61381 = ~pi776 & ~po988;
  assign n61382 = ~pi966 & ~n61381;
  assign n61383 = ~pi966 & ~n61380;
  assign n61384 = ~n61381 & n61383;
  assign n61385 = ~n61380 & n61382;
  assign n61386 = pi1122 & po988;
  assign n61387 = ~pi777 & ~po988;
  assign n61388 = ~pi966 & ~n61387;
  assign n61389 = ~pi966 & ~n61386;
  assign n61390 = ~n61387 & n61389;
  assign n61391 = ~n61386 & n61388;
  assign n61392 = pi779 & ~n60366;
  assign n61393 = pi780 & ~n60361;
  assign n61394 = ~pi604 & ~pi979;
  assign n61395 = pi615 & pi979;
  assign n61396 = ~n61394 & ~n61395;
  assign n61397 = pi604 & ~pi979;
  assign n61398 = ~pi615 & pi979;
  assign n61399 = pi782 & ~n61398;
  assign n61400 = ~n61397 & n61399;
  assign n61401 = pi782 & ~n61396;
  assign n61402 = ~pi782 & ~pi907;
  assign n61403 = ~pi598 & pi979;
  assign n61404 = ~pi624 & ~pi979;
  assign n61405 = pi782 & ~n61404;
  assign n61406 = pi782 & ~n61403;
  assign n61407 = ~n61404 & n61406;
  assign n61408 = ~n61403 & n61405;
  assign n61409 = ~n61402 & ~n65955;
  assign n61410 = ~n65954 & ~n61402;
  assign n61411 = ~n65955 & n61410;
  assign n61412 = ~n65954 & n61409;
  assign n61413 = ~pi782 & pi947;
  assign n61414 = ~n65955 & ~n61413;
  assign n61415 = ~pi923 & ~pi1093;
  assign n61416 = pi1093 & ~pi1154;
  assign n61417 = pi1093 & pi1154;
  assign n61418 = pi923 & ~pi1093;
  assign n61419 = ~n61417 & ~n61418;
  assign n61420 = ~n61415 & ~n61416;
  assign n61421 = ~pi925 & ~pi1093;
  assign n61422 = pi1093 & ~pi1155;
  assign n61423 = pi1093 & pi1155;
  assign n61424 = pi925 & ~pi1093;
  assign n61425 = ~n61423 & ~n61424;
  assign n61426 = ~n61421 & ~n61422;
  assign n61427 = ~pi926 & ~pi1093;
  assign n61428 = pi1093 & ~pi1157;
  assign n61429 = pi1093 & pi1157;
  assign n61430 = pi926 & ~pi1093;
  assign n61431 = ~n61429 & ~n61430;
  assign n61432 = ~n61427 & ~n61428;
  assign n61433 = ~pi931 & ~pi1093;
  assign n61434 = pi1093 & ~pi1150;
  assign n61435 = pi1093 & pi1150;
  assign n61436 = pi931 & ~pi1093;
  assign n61437 = ~n61435 & ~n61436;
  assign n61438 = ~n61433 & ~n61434;
  assign n61439 = ~pi934 & ~pi1093;
  assign n61440 = pi1093 & ~pi1147;
  assign n61441 = pi1093 & pi1147;
  assign n61442 = pi934 & ~pi1093;
  assign n61443 = ~n61441 & ~n61442;
  assign n61444 = ~n61439 & ~n61440;
  assign n61445 = ~pi936 & ~pi1093;
  assign n61446 = pi1093 & ~pi1149;
  assign n61447 = pi1093 & pi1149;
  assign n61448 = pi936 & ~pi1093;
  assign n61449 = ~n61447 & ~n61448;
  assign n61450 = ~n61445 & ~n61446;
  assign n61451 = ~pi937 & ~pi1093;
  assign n61452 = pi1093 & ~pi1148;
  assign n61453 = pi1093 & pi1148;
  assign n61454 = pi937 & ~pi1093;
  assign n61455 = ~n61453 & ~n61454;
  assign n61456 = ~n61451 & ~n61452;
  assign n61457 = ~pi941 & ~pi1093;
  assign n61458 = pi1093 & ~pi1153;
  assign n61459 = pi1093 & pi1153;
  assign n61460 = pi941 & ~pi1093;
  assign n61461 = ~n61459 & ~n61460;
  assign n61462 = ~n61457 & ~n61458;
  assign n61463 = ~pi942 & ~pi1093;
  assign n61464 = pi1093 & ~pi1156;
  assign n61465 = pi1093 & pi1156;
  assign n61466 = pi942 & ~pi1093;
  assign n61467 = ~n61465 & ~n61466;
  assign n61468 = ~n61463 & ~n61464;
  assign n61469 = ~pi943 & ~pi1093;
  assign n61470 = pi1093 & ~pi1151;
  assign n61471 = pi1093 & pi1151;
  assign n61472 = pi943 & ~pi1093;
  assign n61473 = ~n61471 & ~n61472;
  assign n61474 = ~n61469 & ~n61470;
  assign n61475 = ~pi598 & pi615;
  assign n61476 = ~pi604 & ~pi624;
  assign n61477 = pi119 & pi1056;
  assign n61478 = ~pi228 & pi252;
  assign n61479 = ~pi119 & ~n61478;
  assign n61480 = ~pi468 & ~n61479;
  assign n61481 = ~n61477 & n61480;
  assign n61482 = pi119 & pi1077;
  assign n61483 = n61480 & ~n61482;
  assign n61484 = pi119 & pi1073;
  assign n61485 = n61480 & ~n61484;
  assign n61486 = pi119 & pi1041;
  assign n61487 = n61480 & ~n61486;
  assign n61488 = pi119 & pi232;
  assign po236 = ~pi468 & n61488;
  assign n61490 = pi124 & ~pi468;
  assign n61491 = ~pi478 & pi1044;
  assign n61492 = pi298 & pi478;
  assign n61493 = ~pi298 & pi478;
  assign n61494 = ~pi478 & ~pi1044;
  assign n61495 = ~n61493 & ~n61494;
  assign n61496 = ~n61491 & ~n61492;
  assign n61497 = ~pi478 & pi1049;
  assign n61498 = pi303 & pi478;
  assign n61499 = ~pi303 & pi478;
  assign n61500 = ~pi478 & ~pi1049;
  assign n61501 = ~n61499 & ~n61500;
  assign n61502 = ~n61497 & ~n61498;
  assign n61503 = ~pi478 & pi1048;
  assign n61504 = pi304 & pi478;
  assign n61505 = ~pi304 & pi478;
  assign n61506 = ~pi478 & ~pi1048;
  assign n61507 = ~n61505 & ~n61506;
  assign n61508 = ~n61503 & ~n61504;
  assign n61509 = ~pi478 & pi1084;
  assign n61510 = pi305 & pi478;
  assign n61511 = ~pi305 & pi478;
  assign n61512 = ~pi478 & ~pi1084;
  assign n61513 = ~n61511 & ~n61512;
  assign n61514 = ~n61509 & ~n61510;
  assign n61515 = ~pi478 & pi1059;
  assign n61516 = pi306 & pi478;
  assign n61517 = ~pi306 & pi478;
  assign n61518 = ~pi478 & ~pi1059;
  assign n61519 = ~n61517 & ~n61518;
  assign n61520 = ~n61515 & ~n61516;
  assign n61521 = ~pi478 & pi1053;
  assign n61522 = pi307 & pi478;
  assign n61523 = ~pi307 & pi478;
  assign n61524 = ~pi478 & ~pi1053;
  assign n61525 = ~n61523 & ~n61524;
  assign n61526 = ~n61521 & ~n61522;
  assign n61527 = ~pi478 & pi1037;
  assign n61528 = pi308 & pi478;
  assign n61529 = ~pi308 & pi478;
  assign n61530 = ~pi478 & ~pi1037;
  assign n61531 = ~n61529 & ~n61530;
  assign n61532 = ~n61527 & ~n61528;
  assign n61533 = ~pi478 & pi1072;
  assign n61534 = pi309 & pi478;
  assign n61535 = ~pi309 & pi478;
  assign n61536 = ~pi478 & ~pi1072;
  assign n61537 = ~n61535 & ~n61536;
  assign n61538 = ~n61533 & ~n61534;
  assign n61539 = ~pi599 & pi810;
  assign n61540 = pi596 & ~n61539;
  assign n61541 = pi804 & ~n61540;
  assign n61542 = pi815 & ~n61541;
  assign n61543 = pi595 & ~n61542;
  assign n61544 = ~pi804 & ~pi810;
  assign n61545 = ~pi595 & ~n61544;
  assign n61546 = pi594 & pi600;
  assign n61547 = pi597 & n61546;
  assign n61548 = pi601 & n61547;
  assign n61549 = ~n61545 & n61548;
  assign n61550 = ~pi595 & n61544;
  assign n61551 = pi595 & pi815;
  assign n61552 = ~n61541 & n61551;
  assign n61553 = ~n61550 & ~n61552;
  assign n61554 = n61548 & ~n61553;
  assign n61555 = ~n61543 & n61549;
  assign n61556 = ~pi601 & ~n61544;
  assign n61557 = pi600 & ~pi810;
  assign n61558 = pi804 & ~n61557;
  assign n61559 = ~pi815 & ~n61558;
  assign n61560 = ~pi815 & ~n61556;
  assign n61561 = ~n61558 & n61560;
  assign n61562 = ~n61556 & n61559;
  assign n61563 = ~n65975 & ~n65976;
  assign n61564 = pi605 & ~n61563;
  assign n61565 = pi990 & n61546;
  assign n61566 = ~pi815 & n61558;
  assign n61567 = n61565 & n61566;
  assign n61568 = ~n61564 & ~n61567;
  assign po614 = pi821 & ~n61568;
  assign n61570 = ~pi123 & n3112;
  assign n61571 = ~pi591 & n61570;
  assign n61572 = ~pi588 & ~n61570;
  assign n61573 = n48140 & ~n61572;
  assign n61574 = n48140 & ~n61571;
  assign n61575 = ~n61572 & n61574;
  assign n61576 = ~n61571 & n61573;
  assign n61577 = pi590 & ~n61570;
  assign n61578 = pi588 & n61570;
  assign n61579 = n48140 & ~n61578;
  assign n61580 = n48140 & ~n61577;
  assign n61581 = ~n61578 & n61580;
  assign n61582 = ~n61577 & n61579;
  assign n61583 = ~pi592 & n61570;
  assign n61584 = ~pi591 & ~n61570;
  assign n61585 = n48140 & ~n61584;
  assign n61586 = n48140 & ~n61583;
  assign n61587 = ~n61584 & n61586;
  assign n61588 = ~n61583 & n61585;
  assign n61589 = ~pi590 & n61570;
  assign n61590 = ~pi592 & ~n61570;
  assign n61591 = n48140 & ~n61590;
  assign n61592 = n48140 & ~n61589;
  assign n61593 = ~n61590 & n61592;
  assign n61594 = ~n61589 & n61591;
  assign n61595 = ~pi332 & ~pi806;
  assign n61596 = pi990 & n61595;
  assign n61597 = pi595 & n61547;
  assign n61598 = n61596 & n61597;
  assign n61599 = pi596 & n61598;
  assign n61600 = ~pi332 & pi599;
  assign n61601 = ~n61599 & ~n61600;
  assign n61602 = pi599 & n61599;
  assign po756 = ~n61601 & ~n61602;
  assign n61604 = pi605 & ~pi806;
  assign n61605 = n61548 & n61604;
  assign n61606 = ~pi595 & ~n61605;
  assign n61607 = pi595 & n61605;
  assign n61608 = ~pi332 & ~n61607;
  assign n61609 = ~pi332 & ~n61606;
  assign n61610 = ~n61607 & n61609;
  assign n61611 = ~n61606 & n61608;
  assign n61612 = ~pi332 & pi596;
  assign n61613 = ~n61598 & ~n61612;
  assign po753 = ~n61599 & ~n61613;
  assign n61615 = ~pi806 & n61565;
  assign n61616 = pi597 & n61615;
  assign n61617 = ~pi597 & ~n61615;
  assign n61618 = ~pi332 & ~n61617;
  assign n61619 = ~pi332 & ~n61616;
  assign n61620 = ~n61617 & n61619;
  assign n61621 = ~n61616 & n61618;
  assign n61622 = pi600 & n61596;
  assign n61623 = ~pi332 & pi594;
  assign n61624 = ~n61622 & ~n61623;
  assign po751 = ~n61615 & ~n61624;
  assign n61626 = ~pi332 & pi600;
  assign n61627 = ~n61596 & ~n61626;
  assign po757 = ~n61622 & ~n61627;
  assign n61629 = ~pi601 & pi806;
  assign n61630 = ~pi806 & ~pi989;
  assign n61631 = ~pi332 & ~n61630;
  assign n61632 = ~pi332 & ~n61629;
  assign n61633 = ~n61630 & n61632;
  assign n61634 = ~n61629 & n61631;
  assign n61635 = ~pi287 & pi457;
  assign po444 = ~pi332 & ~n61635;
  assign n61637 = ~pi605 & ~n61595;
  assign n61638 = ~pi332 & ~n61604;
  assign po762 = ~n61637 & n61638;
  assign n61640 = pi721 & pi813;
  assign n61641 = ~pi765 & ~pi798;
  assign n61642 = pi765 & pi798;
  assign n61643 = pi765 & ~pi798;
  assign n61644 = ~pi765 & pi798;
  assign n61645 = ~n61643 & ~n61644;
  assign n61646 = ~n61641 & ~n61642;
  assign n61647 = pi807 & n65984;
  assign n61648 = pi747 & n61647;
  assign n61649 = ~pi747 & ~pi807;
  assign n61650 = n65984 & n61649;
  assign n61651 = ~n61648 & ~n61650;
  assign n61652 = ~pi771 & ~pi800;
  assign n61653 = pi771 & pi800;
  assign n61654 = ~n61652 & ~n61653;
  assign n61655 = ~pi769 & ~pi794;
  assign n61656 = pi769 & pi794;
  assign n61657 = ~n61655 & ~n61656;
  assign n61658 = ~n61654 & ~n61657;
  assign n61659 = ~n61651 & ~n61657;
  assign n61660 = ~n61654 & n61659;
  assign n61661 = ~n61651 & n61658;
  assign n61662 = ~pi773 & ~pi801;
  assign n61663 = pi773 & pi801;
  assign n61664 = pi773 & ~pi801;
  assign n61665 = ~pi773 & pi801;
  assign n61666 = ~n61664 & ~n61665;
  assign n61667 = ~n61662 & ~n61663;
  assign n61668 = n65985 & n65986;
  assign n61669 = n61640 & n61668;
  assign n61670 = ~pi775 & ~pi816;
  assign n61671 = pi775 & pi816;
  assign n61672 = ~n61670 & ~n61671;
  assign n61673 = n61669 & ~n61672;
  assign n61674 = pi731 & ~pi945;
  assign n61675 = pi775 & n61674;
  assign n61676 = pi988 & n61675;
  assign n61677 = ~n61673 & ~n61676;
  assign n61678 = ~pi945 & pi988;
  assign n61679 = pi731 & n61678;
  assign n61680 = ~pi731 & ~pi795;
  assign n61681 = pi731 & pi795;
  assign n61682 = ~n61680 & ~n61681;
  assign n61683 = ~n61679 & n61682;
  assign n61684 = ~n61677 & ~n61683;
  assign n61685 = pi721 & ~pi775;
  assign n61686 = ~n61673 & n61685;
  assign n61687 = n61673 & ~n61682;
  assign n61688 = pi721 & ~n61679;
  assign n61689 = ~n61687 & n61688;
  assign n61690 = ~n61686 & ~n61689;
  assign n61691 = pi721 & ~n61684;
  assign n61692 = ~pi721 & ~pi813;
  assign n61693 = pi794 & pi801;
  assign n61694 = n61692 & n61693;
  assign n61695 = ~n61654 & n61694;
  assign n61696 = n61647 & ~n61654;
  assign n61697 = n61694 & n61696;
  assign n61698 = n61647 & n61695;
  assign n61699 = ~n61669 & ~n65988;
  assign n61700 = pi816 & ~n61699;
  assign n61701 = pi775 & ~n61700;
  assign n61702 = pi795 & ~n61701;
  assign n61703 = pi747 & pi773;
  assign n61704 = pi769 & pi775;
  assign n61705 = pi775 & n61703;
  assign n61706 = pi769 & n61705;
  assign n61707 = n61703 & n61704;
  assign n61708 = pi721 & n65989;
  assign n61709 = ~pi721 & ~n65989;
  assign n61710 = n61679 & ~n61709;
  assign n61711 = pi769 & n61703;
  assign n61712 = pi721 & n61711;
  assign n61713 = ~pi721 & ~n61711;
  assign n61714 = pi775 & ~n61713;
  assign n61715 = pi775 & ~n61712;
  assign n61716 = ~n61713 & n61715;
  assign n61717 = ~n61712 & n61714;
  assign n61718 = ~n61685 & ~n65990;
  assign n61719 = n61679 & ~n61718;
  assign n61720 = ~n61708 & n61710;
  assign n61721 = ~n61700 & n65990;
  assign n61722 = pi795 & ~n61721;
  assign n61723 = n65991 & ~n61722;
  assign n61724 = ~n61702 & n65991;
  assign n61725 = n65987 & ~n65992;
  assign n61726 = ~n61640 & ~n61692;
  assign n61727 = n61668 & ~n61726;
  assign n61728 = pi795 & ~n61672;
  assign n61729 = n61727 & n61728;
  assign n61730 = pi731 & n61729;
  assign n61731 = n61678 & n61703;
  assign n61732 = pi731 & n61731;
  assign n61733 = n61679 & n61703;
  assign n61734 = ~n61672 & ~n61726;
  assign n61735 = ~n61654 & n61734;
  assign n61736 = ~pi795 & pi801;
  assign n61737 = ~n61657 & n61736;
  assign n61738 = n61647 & n61737;
  assign n61739 = n61734 & n61737;
  assign n61740 = n61696 & n61739;
  assign n61741 = n61735 & n61738;
  assign n61742 = n61731 & ~n65994;
  assign n61743 = ~pi731 & ~n61742;
  assign n61744 = ~n65993 & ~n61743;
  assign n61745 = ~n61703 & ~n61729;
  assign n61746 = n61679 & ~n61745;
  assign n61747 = pi731 & ~n61729;
  assign n61748 = n61703 & ~n65994;
  assign n61749 = ~pi731 & ~n61748;
  assign n61750 = n61678 & ~n61749;
  assign n61751 = ~n61747 & ~n61750;
  assign n61752 = ~n61746 & ~n61751;
  assign n61753 = ~n61730 & n61744;
  assign n61754 = pi801 & n61650;
  assign n61755 = pi773 & n61678;
  assign n61756 = n65986 & ~n61755;
  assign n61757 = n61647 & n61756;
  assign n61758 = ~n61754 & ~n61757;
  assign n61759 = ~n61682 & n61734;
  assign n61760 = n61658 & n61759;
  assign n61761 = ~n61758 & n61760;
  assign n61762 = ~pi747 & ~n61755;
  assign n61763 = ~n61731 & ~n61762;
  assign po904 = ~n61761 & n61763;
  assign n61765 = n61671 & n61727;
  assign n61766 = pi794 & n65986;
  assign n61767 = ~n61654 & n61766;
  assign n61768 = n61734 & n61767;
  assign n61769 = n61735 & n61766;
  assign n61770 = ~n61651 & n65996;
  assign n61771 = ~pi775 & n61770;
  assign n61772 = ~n61765 & ~n61771;
  assign n61773 = pi795 & ~n61772;
  assign n61774 = ~pi769 & ~n61705;
  assign n61775 = n61679 & ~n65989;
  assign n61776 = pi769 & ~n61705;
  assign n61777 = ~pi769 & n61705;
  assign n61778 = ~n61776 & ~n61777;
  assign n61779 = n61679 & ~n61778;
  assign n61780 = ~n61774 & n61775;
  assign n61781 = ~n61773 & n65997;
  assign n61782 = ~n61682 & n61770;
  assign n61783 = pi769 & ~n61679;
  assign n61784 = ~n61782 & n61783;
  assign n61785 = ~n61781 & ~n61784;
  assign n61786 = ~pi765 & ~pi773;
  assign n61787 = ~n61653 & n61786;
  assign n61788 = ~n61656 & n61787;
  assign n61789 = ~n61648 & n61788;
  assign n61790 = ~pi765 & ~n61653;
  assign n61791 = ~n61656 & n61790;
  assign n61792 = ~n61648 & n61791;
  assign n61793 = n61662 & ~n61792;
  assign n61794 = ~n61663 & ~n61793;
  assign n61795 = n65985 & ~n61794;
  assign n61796 = n61668 & ~n61789;
  assign n61797 = ~pi721 & ~n65998;
  assign n61798 = n61670 & ~n61797;
  assign n61799 = ~n61671 & ~n61798;
  assign n61800 = n61680 & ~n61799;
  assign n61801 = ~n61672 & n61681;
  assign n61802 = ~n61800 & ~n61801;
  assign po963 = n61727 & ~n61802;
  assign n61804 = ~pi945 & pi987;
  assign n61805 = ~po963 & n61804;
  assign po978 = n61668 & n61759;
  assign n61807 = pi771 & pi945;
  assign n61808 = ~po978 & n61807;
  assign n61809 = ~n61805 & ~n61808;
  assign n61810 = ~pi801 & n65985;
  assign n61811 = po963 & n61810;
  assign n61812 = n61678 & ~n61811;
  assign n61813 = pi801 & n61759;
  assign n61814 = n65985 & n61813;
  assign n61815 = pi801 & ~n61759;
  assign n61816 = n61668 & ~n61815;
  assign n61817 = pi773 & ~n61816;
  assign n61818 = pi773 & ~n61814;
  assign n61819 = ~n61812 & ~n65999;
  assign po930 = ~n61755 & ~n61819;
  assign n61821 = pi765 & ~po978;
  assign n61822 = pi945 & ~n61821;
  assign n61823 = ~n61669 & ~n61692;
  assign n61824 = n61798 & ~n61823;
  assign n61825 = ~n61765 & ~n61824;
  assign n61826 = n61680 & ~n61825;
  assign n61827 = ~pi765 & ~n61730;
  assign n61828 = ~pi765 & ~n61765;
  assign n61829 = ~n61824 & n61828;
  assign n61830 = ~pi795 & ~n61829;
  assign n61831 = ~pi731 & ~n61830;
  assign n61832 = ~n61747 & ~n61831;
  assign n61833 = ~pi765 & ~n61832;
  assign n61834 = ~n61826 & n61827;
  assign n61835 = ~pi945 & ~n66000;
  assign po922 = ~n61822 & ~n61835;
  assign n61837 = pi765 & pi771;
  assign n61838 = n61703 & n61837;
  assign n61839 = ~n61729 & ~n61838;
  assign n61840 = n61675 & ~n61839;
  assign n61841 = pi775 & ~po978;
  assign n61842 = pi795 & pi800;
  assign n61843 = pi801 & ~pi816;
  assign n61844 = n61842 & n61843;
  assign n61845 = ~n61657 & n61844;
  assign n61846 = ~n61726 & n61845;
  assign n61847 = ~n61726 & n61844;
  assign n61848 = n61659 & n61847;
  assign n61849 = ~n61651 & n61846;
  assign n61850 = n61838 & ~n66001;
  assign n61851 = ~pi775 & ~n61850;
  assign n61852 = n61674 & ~n61851;
  assign n61853 = ~n61674 & po978;
  assign n61854 = pi775 & ~n61853;
  assign n61855 = n61674 & n61838;
  assign n61856 = ~n66001 & n61855;
  assign n61857 = ~n61854 & ~n61856;
  assign n61858 = ~n61841 & ~n61852;
  assign po932 = ~n61840 & ~n66002;
  assign n61860 = pi832 & pi956;
  assign n61861 = ~pi1046 & ~pi1083;
  assign n61862 = pi1085 & n61861;
  assign n61863 = n61860 & n61862;
  assign n61864 = ~pi968 & n61863;
  assign n61865 = pi778 & ~n61864;
  assign n61866 = pi1100 & n61864;
  assign n61867 = ~n61865 & ~n61866;
  assign n61868 = pi781 & ~n61864;
  assign n61869 = pi1101 & n61864;
  assign n61870 = ~n61868 & ~n61869;
  assign n61871 = pi783 & ~n61864;
  assign n61872 = pi1109 & n61864;
  assign n61873 = ~n61871 & ~n61872;
  assign n61874 = pi784 & ~n61864;
  assign n61875 = pi1110 & n61864;
  assign n61876 = ~n61874 & ~n61875;
  assign n61877 = pi785 & ~n61864;
  assign n61878 = pi1102 & n61864;
  assign n61879 = ~n61877 & ~n61878;
  assign n61880 = pi787 & ~n61864;
  assign n61881 = pi1104 & n61864;
  assign n61882 = ~n61880 & ~n61881;
  assign n61883 = pi788 & ~n61864;
  assign n61884 = pi1105 & n61864;
  assign n61885 = ~n61883 & ~n61884;
  assign n61886 = pi789 & ~n61864;
  assign n61887 = pi1106 & n61864;
  assign n61888 = ~n61886 & ~n61887;
  assign n61889 = pi790 & ~n61864;
  assign n61890 = pi1107 & n61864;
  assign n61891 = ~n61889 & ~n61890;
  assign n61892 = pi791 & ~n61864;
  assign n61893 = pi1108 & n61864;
  assign n61894 = ~n61892 & ~n61893;
  assign n61895 = pi792 & ~n61864;
  assign n61896 = pi1103 & n61864;
  assign n61897 = ~n61895 & ~n61896;
  assign n61898 = pi968 & n61863;
  assign n61899 = pi794 & ~n61898;
  assign n61900 = pi1130 & n61898;
  assign n61901 = ~n61899 & ~n61900;
  assign n61902 = pi795 & ~n61898;
  assign n61903 = pi1128 & n61898;
  assign n61904 = ~n61902 & ~n61903;
  assign n61905 = pi798 & ~n61898;
  assign n61906 = pi1124 & n61898;
  assign n61907 = ~n61905 & ~n61906;
  assign n61908 = pi799 & ~n61898;
  assign n61909 = ~pi1107 & n61898;
  assign po956 = ~n61908 & ~n61909;
  assign n61911 = pi800 & ~n61898;
  assign n61912 = pi1125 & n61898;
  assign n61913 = ~n61911 & ~n61912;
  assign n61914 = pi801 & ~n61898;
  assign n61915 = pi1126 & n61898;
  assign n61916 = ~n61914 & ~n61915;
  assign n61917 = pi803 & ~n61898;
  assign n61918 = ~pi1106 & n61898;
  assign po960 = ~n61917 & ~n61918;
  assign n61920 = pi804 & ~n61898;
  assign n61921 = pi1109 & n61898;
  assign n61922 = ~n61920 & ~n61921;
  assign n61923 = pi807 & ~n61898;
  assign n61924 = pi1127 & n61898;
  assign n61925 = ~n61923 & ~n61924;
  assign n61926 = pi808 & ~n61898;
  assign n61927 = pi1101 & n61898;
  assign n61928 = ~n61926 & ~n61927;
  assign n61929 = pi809 & ~n61898;
  assign n61930 = ~pi1103 & n61898;
  assign po966 = ~n61929 & ~n61930;
  assign n61932 = pi810 & ~n61898;
  assign n61933 = pi1108 & n61898;
  assign n61934 = ~n61932 & ~n61933;
  assign n61935 = pi811 & ~n61898;
  assign n61936 = pi1102 & n61898;
  assign n61937 = ~n61935 & ~n61936;
  assign n61938 = pi812 & ~n61898;
  assign n61939 = ~pi1104 & n61898;
  assign po969 = ~n61938 & ~n61939;
  assign n61941 = pi813 & ~n61898;
  assign n61942 = pi1131 & n61898;
  assign n61943 = ~n61941 & ~n61942;
  assign n61944 = pi814 & ~n61898;
  assign n61945 = ~pi1105 & n61898;
  assign po971 = ~n61944 & ~n61945;
  assign n61947 = pi815 & ~n61898;
  assign n61948 = pi1110 & n61898;
  assign n61949 = ~n61947 & ~n61948;
  assign n61950 = pi816 & ~n61898;
  assign n61951 = pi1129 & n61898;
  assign n61952 = ~n61950 & ~n61951;
  assign po979 = ~pi811 & ~pi893;
  assign n61954 = ~pi955 & pi1049;
  assign n61955 = pi837 & pi955;
  assign n61956 = ~pi837 & pi955;
  assign n61957 = ~pi955 & ~pi1049;
  assign n61958 = ~n61956 & ~n61957;
  assign n61959 = ~n61954 & ~n61955;
  assign n61960 = ~pi955 & pi1047;
  assign n61961 = pi838 & pi955;
  assign n61962 = ~pi838 & pi955;
  assign n61963 = ~pi955 & ~pi1047;
  assign n61964 = ~n61962 & ~n61963;
  assign n61965 = ~n61960 & ~n61961;
  assign n61966 = ~pi955 & pi1074;
  assign n61967 = pi839 & pi955;
  assign n61968 = ~pi839 & pi955;
  assign n61969 = ~pi955 & ~pi1074;
  assign n61970 = ~n61968 & ~n61969;
  assign n61971 = ~n61966 & ~n61967;
  assign n61972 = ~pi955 & pi1035;
  assign n61973 = pi842 & pi955;
  assign n61974 = ~pi842 & pi955;
  assign n61975 = ~pi955 & ~pi1035;
  assign n61976 = ~n61974 & ~n61975;
  assign n61977 = ~n61972 & ~n61973;
  assign n61978 = ~pi955 & pi1079;
  assign n61979 = pi843 & pi955;
  assign n61980 = ~pi843 & pi955;
  assign n61981 = ~pi955 & ~pi1079;
  assign n61982 = ~n61980 & ~n61981;
  assign n61983 = ~n61978 & ~n61979;
  assign n61984 = ~pi955 & pi1078;
  assign n61985 = pi844 & pi955;
  assign n61986 = ~pi844 & pi955;
  assign n61987 = ~pi955 & ~pi1078;
  assign n61988 = ~n61986 & ~n61987;
  assign n61989 = ~n61984 & ~n61985;
  assign n61990 = ~pi955 & pi1043;
  assign n61991 = pi845 & pi955;
  assign n61992 = ~pi845 & pi955;
  assign n61993 = ~pi955 & ~pi1043;
  assign n61994 = ~n61992 & ~n61993;
  assign n61995 = ~n61990 & ~n61991;
  assign n61996 = ~pi955 & pi1055;
  assign n61997 = pi847 & pi955;
  assign n61998 = ~pi847 & pi955;
  assign n61999 = ~pi955 & ~pi1055;
  assign n62000 = ~n61998 & ~n61999;
  assign n62001 = ~n61996 & ~n61997;
  assign n62002 = ~pi955 & pi1039;
  assign n62003 = pi848 & pi955;
  assign n62004 = ~pi848 & pi955;
  assign n62005 = ~pi955 & ~pi1039;
  assign n62006 = ~n62004 & ~n62005;
  assign n62007 = ~n62002 & ~n62003;
  assign n62008 = ~pi955 & pi1048;
  assign n62009 = pi850 & pi955;
  assign n62010 = ~pi850 & pi955;
  assign n62011 = ~pi955 & ~pi1048;
  assign n62012 = ~n62010 & ~n62011;
  assign n62013 = ~n62008 & ~n62009;
  assign n62014 = ~pi955 & pi1045;
  assign n62015 = pi851 & pi955;
  assign n62016 = ~pi851 & pi955;
  assign n62017 = ~pi955 & ~pi1045;
  assign n62018 = ~n62016 & ~n62017;
  assign n62019 = ~n62014 & ~n62015;
  assign n62020 = ~pi955 & pi1062;
  assign n62021 = pi852 & pi955;
  assign n62022 = ~pi852 & pi955;
  assign n62023 = ~pi955 & ~pi1062;
  assign n62024 = ~n62022 & ~n62023;
  assign n62025 = ~n62020 & ~n62021;
  assign n62026 = ~pi955 & pi1080;
  assign n62027 = pi853 & pi955;
  assign n62028 = ~pi853 & pi955;
  assign n62029 = ~pi955 & ~pi1080;
  assign n62030 = ~n62028 & ~n62029;
  assign n62031 = ~n62026 & ~n62027;
  assign n62032 = ~pi955 & pi1051;
  assign n62033 = pi854 & pi955;
  assign n62034 = ~pi854 & pi955;
  assign n62035 = ~pi955 & ~pi1051;
  assign n62036 = ~n62034 & ~n62035;
  assign n62037 = ~n62032 & ~n62033;
  assign n62038 = ~pi955 & pi1065;
  assign n62039 = pi855 & pi955;
  assign n62040 = ~pi855 & pi955;
  assign n62041 = ~pi955 & ~pi1065;
  assign n62042 = ~n62040 & ~n62041;
  assign n62043 = ~n62038 & ~n62039;
  assign n62044 = ~pi955 & pi1067;
  assign n62045 = pi856 & pi955;
  assign n62046 = ~pi856 & pi955;
  assign n62047 = ~pi955 & ~pi1067;
  assign n62048 = ~n62046 & ~n62047;
  assign n62049 = ~n62044 & ~n62045;
  assign n62050 = ~pi955 & pi1058;
  assign n62051 = pi857 & pi955;
  assign n62052 = ~pi857 & pi955;
  assign n62053 = ~pi955 & ~pi1058;
  assign n62054 = ~n62052 & ~n62053;
  assign n62055 = ~n62050 & ~n62051;
  assign n62056 = ~pi955 & pi1087;
  assign n62057 = pi858 & pi955;
  assign n62058 = ~pi858 & pi955;
  assign n62059 = ~pi955 & ~pi1087;
  assign n62060 = ~n62058 & ~n62059;
  assign n62061 = ~n62056 & ~n62057;
  assign n62062 = ~pi955 & pi1070;
  assign n62063 = pi859 & pi955;
  assign n62064 = ~pi859 & pi955;
  assign n62065 = ~pi955 & ~pi1070;
  assign n62066 = ~n62064 & ~n62065;
  assign n62067 = ~n62062 & ~n62063;
  assign n62068 = ~pi955 & pi1076;
  assign n62069 = pi860 & pi955;
  assign n62070 = ~pi860 & pi955;
  assign n62071 = ~pi955 & ~pi1076;
  assign n62072 = ~n62070 & ~n62071;
  assign n62073 = ~n62068 & ~n62069;
  assign n62074 = ~pi955 & pi1040;
  assign n62075 = pi865 & pi955;
  assign n62076 = ~pi865 & pi955;
  assign n62077 = ~pi955 & ~pi1040;
  assign n62078 = ~n62076 & ~n62077;
  assign n62079 = ~n62074 & ~n62075;
  assign n62080 = ~pi955 & pi1053;
  assign n62081 = pi866 & pi955;
  assign n62082 = ~pi866 & pi955;
  assign n62083 = ~pi955 & ~pi1053;
  assign n62084 = ~n62082 & ~n62083;
  assign n62085 = ~n62080 & ~n62081;
  assign n62086 = ~pi955 & pi1057;
  assign n62087 = pi867 & pi955;
  assign n62088 = ~pi867 & pi955;
  assign n62089 = ~pi955 & ~pi1057;
  assign n62090 = ~n62088 & ~n62089;
  assign n62091 = ~n62086 & ~n62087;
  assign n62092 = ~pi955 & pi1063;
  assign n62093 = pi868 & pi955;
  assign n62094 = ~pi868 & pi955;
  assign n62095 = ~pi955 & ~pi1063;
  assign n62096 = ~n62094 & ~n62095;
  assign n62097 = ~n62092 & ~n62093;
  assign n62098 = ~pi955 & pi1069;
  assign n62099 = pi870 & pi955;
  assign n62100 = ~pi870 & pi955;
  assign n62101 = ~pi955 & ~pi1069;
  assign n62102 = ~n62100 & ~n62101;
  assign n62103 = ~n62098 & ~n62099;
  assign n62104 = ~pi955 & pi1072;
  assign n62105 = pi871 & pi955;
  assign n62106 = ~pi871 & pi955;
  assign n62107 = ~pi955 & ~pi1072;
  assign n62108 = ~n62106 & ~n62107;
  assign n62109 = ~n62104 & ~n62105;
  assign n62110 = ~pi955 & pi1084;
  assign n62111 = pi872 & pi955;
  assign n62112 = ~pi872 & pi955;
  assign n62113 = ~pi955 & ~pi1084;
  assign n62114 = ~n62112 & ~n62113;
  assign n62115 = ~n62110 & ~n62111;
  assign n62116 = ~pi955 & pi1044;
  assign n62117 = pi873 & pi955;
  assign n62118 = ~pi873 & pi955;
  assign n62119 = ~pi955 & ~pi1044;
  assign n62120 = ~n62118 & ~n62119;
  assign n62121 = ~n62116 & ~n62117;
  assign n62122 = ~pi955 & pi1036;
  assign n62123 = pi874 & pi955;
  assign n62124 = ~pi874 & pi955;
  assign n62125 = ~pi955 & ~pi1036;
  assign n62126 = ~n62124 & ~n62125;
  assign n62127 = ~n62122 & ~n62123;
  assign n62128 = ~pi955 & pi1037;
  assign n62129 = pi876 & pi955;
  assign n62130 = ~pi876 & pi955;
  assign n62131 = ~pi955 & ~pi1037;
  assign n62132 = ~n62130 & ~n62131;
  assign n62133 = ~n62128 & ~n62129;
  assign n62134 = ~pi955 & pi1081;
  assign n62135 = pi880 & pi955;
  assign n62136 = ~pi880 & pi955;
  assign n62137 = ~pi955 & ~pi1081;
  assign n62138 = ~n62136 & ~n62137;
  assign n62139 = ~n62134 & ~n62135;
  assign n62140 = ~pi955 & pi1059;
  assign n62141 = pi881 & pi955;
  assign n62142 = ~pi881 & pi955;
  assign n62143 = ~pi955 & ~pi1059;
  assign n62144 = ~n62142 & ~n62143;
  assign n62145 = ~n62140 & ~n62141;
  assign n62146 = ~pi883 & n60918;
  assign n62147 = ~n61018 & ~n62146;
  assign n62148 = pi1124 & ~n60918;
  assign n62149 = ~pi884 & n60918;
  assign n62150 = ~n62148 & ~n62149;
  assign n62151 = pi1125 & ~n60918;
  assign n62152 = ~pi885 & n60918;
  assign n62153 = ~n62151 & ~n62152;
  assign n62154 = pi1109 & ~n60918;
  assign n62155 = ~pi886 & n60918;
  assign n62156 = ~n62154 & ~n62155;
  assign n62157 = ~pi887 & n60918;
  assign n62158 = ~n61017 & ~n62157;
  assign n62159 = pi1120 & ~n60918;
  assign n62160 = ~pi888 & n60918;
  assign n62161 = ~n62159 & ~n62160;
  assign n62162 = pi1103 & ~n60918;
  assign n62163 = ~pi889 & n60918;
  assign n62164 = ~n62162 & ~n62163;
  assign n62165 = pi1126 & ~n60918;
  assign n62166 = ~pi890 & n60918;
  assign n62167 = ~n62165 & ~n62166;
  assign n62168 = pi1116 & ~n60918;
  assign n62169 = ~pi891 & n60918;
  assign n62170 = ~n62168 & ~n62169;
  assign n62171 = pi1101 & ~n60918;
  assign n62172 = ~pi892 & n60918;
  assign n62173 = ~n62171 & ~n62172;
  assign n62174 = pi1119 & ~n60918;
  assign n62175 = ~pi894 & n60918;
  assign n62176 = ~n62174 & ~n62175;
  assign n62177 = pi1113 & ~n60918;
  assign n62178 = ~pi895 & n60918;
  assign n62179 = ~n62177 & ~n62178;
  assign n62180 = pi1118 & ~n60918;
  assign n62181 = ~pi896 & n60918;
  assign n62182 = ~n62180 & ~n62181;
  assign n62183 = pi1129 & ~n60918;
  assign n62184 = ~pi898 & n60918;
  assign n62185 = ~n62183 & ~n62184;
  assign n62186 = ~pi899 & n60918;
  assign n62187 = ~n61066 & ~n62186;
  assign n62188 = pi1110 & ~n60918;
  assign n62189 = ~pi900 & n60918;
  assign n62190 = ~n62188 & ~n62189;
  assign n62191 = pi1111 & ~n60918;
  assign n62192 = ~pi902 & n60918;
  assign n62193 = ~n62191 & ~n62192;
  assign n62194 = pi1121 & ~n60918;
  assign n62195 = ~pi903 & n60918;
  assign n62196 = ~n62194 & ~n62195;
  assign n62197 = ~pi904 & n60918;
  assign n62198 = ~n60920 & ~n62197;
  assign n62199 = ~pi905 & n60918;
  assign n62200 = ~n60919 & ~n62199;
  assign n62201 = pi1128 & ~n60918;
  assign n62202 = ~pi906 & n60918;
  assign n62203 = ~n62201 & ~n62202;
  assign n62204 = ~pi908 & n60918;
  assign n62205 = ~n60969 & ~n62204;
  assign n62206 = pi1105 & ~n60918;
  assign n62207 = ~pi909 & n60918;
  assign n62208 = ~n62206 & ~n62207;
  assign n62209 = pi1117 & ~n60918;
  assign n62210 = ~pi910 & n60918;
  assign n62211 = ~n62209 & ~n62210;
  assign n62212 = pi1130 & ~n60918;
  assign n62213 = ~pi911 & n60918;
  assign n62214 = ~n62212 & ~n62213;
  assign n62215 = ~pi912 & n60918;
  assign n62216 = ~n61067 & ~n62215;
  assign n62217 = pi1106 & ~n60918;
  assign n62218 = ~pi913 & n60918;
  assign n62219 = ~n62217 & ~n62218;
  assign n62220 = pi1108 & ~n60918;
  assign n62221 = ~pi915 & n60918;
  assign n62222 = ~n62220 & ~n62221;
  assign n62223 = ~pi916 & n60918;
  assign n62224 = ~n60968 & ~n62223;
  assign n62225 = pi1112 & ~n60918;
  assign n62226 = ~pi917 & n60918;
  assign n62227 = ~n62225 & ~n62226;
  assign n62228 = pi1104 & ~n60918;
  assign n62229 = ~pi918 & n60918;
  assign n62230 = ~n62228 & ~n62229;
  assign n62231 = pi1102 & ~n60918;
  assign n62232 = ~pi919 & n60918;
  assign n62233 = ~n62231 & ~n62232;
  assign n62234 = pi846 & n65723;
  assign n62235 = pi1134 & ~n65723;
  assign n62236 = ~n62234 & ~n62235;
  assign n62237 = pi861 & ~pi1093;
  assign n62238 = ~n49011 & ~n62237;
  assign n62239 = ~pi228 & ~n62238;
  assign n62240 = pi123 & ~pi861;
  assign n62241 = ~pi123 & ~pi1141;
  assign n62242 = pi228 & ~n62241;
  assign n62243 = pi228 & ~n62240;
  assign n62244 = ~n62241 & n62243;
  assign n62245 = ~n62240 & n62242;
  assign n62246 = ~n62239 & ~n66035;
  assign n62247 = pi862 & n65723;
  assign n62248 = pi1139 & ~n65723;
  assign n62249 = ~n62247 & ~n62248;
  assign n62250 = pi869 & ~pi1093;
  assign n62251 = ~n48981 & ~n62250;
  assign n62252 = ~pi228 & ~n62251;
  assign n62253 = pi123 & ~pi869;
  assign n62254 = ~pi123 & ~pi1140;
  assign n62255 = pi228 & ~n62254;
  assign n62256 = pi228 & ~n62253;
  assign n62257 = ~n62254 & n62256;
  assign n62258 = ~n62253 & n62255;
  assign n62259 = ~n62252 & ~n66036;
  assign n62260 = ~pi875 & ~pi1093;
  assign n62261 = ~n48990 & ~n62260;
  assign n62262 = ~pi228 & ~n62261;
  assign n62263 = pi123 & pi875;
  assign n62264 = ~pi123 & pi1136;
  assign n62265 = pi228 & ~n62264;
  assign n62266 = pi228 & ~n62263;
  assign n62267 = ~n62264 & n62266;
  assign n62268 = ~n62263 & n62265;
  assign po1031 = ~n62262 & ~n66037;
  assign n62270 = pi877 & ~pi1093;
  assign n62271 = ~n49023 & ~n62270;
  assign n62272 = ~pi228 & ~n62271;
  assign n62273 = pi123 & ~pi877;
  assign n62274 = ~pi123 & ~pi1138;
  assign n62275 = pi228 & ~n62274;
  assign n62276 = pi228 & ~n62273;
  assign n62277 = ~n62274 & n62276;
  assign n62278 = ~n62273 & n62275;
  assign n62279 = ~n62272 & ~n66038;
  assign n62280 = pi878 & ~pi1093;
  assign n62281 = ~n49008 & ~n62280;
  assign n62282 = ~pi228 & ~n62281;
  assign n62283 = pi123 & ~pi878;
  assign n62284 = ~pi123 & ~pi1137;
  assign n62285 = pi228 & ~n62284;
  assign n62286 = pi228 & ~n62283;
  assign n62287 = ~n62284 & n62286;
  assign n62288 = ~n62283 & n62285;
  assign n62289 = ~n62282 & ~n66039;
  assign n62290 = pi879 & ~pi1093;
  assign n62291 = ~n49014 & ~n62290;
  assign n62292 = ~pi228 & ~n62291;
  assign n62293 = pi123 & ~pi879;
  assign n62294 = ~pi123 & ~pi1135;
  assign n62295 = pi228 & ~n62294;
  assign n62296 = pi228 & ~n62293;
  assign n62297 = ~n62294 & n62296;
  assign n62298 = ~n62293 & n62295;
  assign n62299 = ~n62292 & ~n66040;
  assign n62300 = pi840 & ~n2923;
  assign n62301 = pi1196 & n2923;
  assign n62302 = ~n62300 & ~n62301;
  assign n62303 = pi849 & ~n2923;
  assign n62304 = pi1198 & n2923;
  assign n62305 = ~n62303 & ~n62304;
  assign n62306 = pi863 & ~n2923;
  assign n62307 = pi1199 & n2923;
  assign n62308 = ~n62306 & ~n62307;
  assign n62309 = pi864 & ~n2923;
  assign n62310 = pi1197 & n2923;
  assign n62311 = ~n62309 & ~n62310;
  assign po991 = pi946 & n2923;
  assign n62313 = ~pi922 & ~pi1093;
  assign n62314 = pi1093 & ~pi1152;
  assign n62315 = pi1093 & pi1152;
  assign n62316 = pi922 & ~pi1093;
  assign n62317 = ~n62315 & ~n62316;
  assign n62318 = ~n62313 & ~n62314;
  assign po1115 = ~pi782 & pi960;
  assign po1116 = ~pi230 & pi961;
  assign po1118 = ~pi782 & pi963;
  assign po1122 = ~pi230 & pi967;
  assign po1124 = ~pi230 & pi969;
  assign po1125 = ~pi782 & pi970;
  assign po1126 = ~pi230 & pi971;
  assign po1127 = ~pi782 & pi972;
  assign po1128 = ~pi230 & pi974;
  assign po1129 = ~pi782 & pi975;
  assign po1131 = ~pi230 & pi977;
  assign po1132 = ~pi782 & pi978;
  assign n62331 = n2441 | ~n2442;
  assign n62332 = n2447 | ~n2448;
  assign n62333 = n2456 | ~n2457;
  assign n62334 = n2467 | ~n2468;
  assign n62335 = n2474 | ~n2480 | n2489 | n2490;
  assign n62336 = n2495 | ~n2496;
  assign n62337 = n2504 | ~n2505;
  assign n62338 = n2510 | n2511;
  assign n62339 = n2516 | ~n2517;
  assign n62340 = n2528 | ~n2529;
  assign n62341 = n2534 | ~n2535;
  assign n62342 = n2549 | ~n2561 | ~n2570 | ~n2571;
  assign n62343 = n2576 | n2577;
  assign n62344 = n2604 | n2605;
  assign n62345 = n2608 | n2609;
  assign n62346 = n2618 | n2619;
  assign n62347 = n2622 | n2623;
  assign n62348 = n2628 | n2629;
  assign n62349 = n2635 | n2631 | n2634;
  assign n62350 = n2644 | n2645;
  assign n62351 = n2649 | n2646 | n2648;
  assign n62352 = n2651 | n2652;
  assign n62353 = n2653 | n2654;
  assign n62354 = n2656 | n2657;
  assign n62355 = n2666 | n2667;
  assign n62356 = n2668 | n2669;
  assign n62357 = n2672 | n2673;
  assign n62358 = n2679 | n2680;
  assign n62359 = n2691 | n2692;
  assign n62360 = n2700 | n2701 | n2703 | n2704;
  assign n62361 = n2705 | n2706;
  assign n62362 = n2713 | n2709 | n2712;
  assign n62363 = n2717 | n2718;
  assign n62364 = n2721 | n2722;
  assign n62365 = n2723 | n2724;
  assign n62366 = n2731 | n2732;
  assign n62367 = n2734 | n2735;
  assign n62368 = n2737 | n2738;
  assign n62369 = n2744 | n2745;
  assign n62370 = n2754 | n2749 | n2753;
  assign n62371 = n2756 | n2757;
  assign n62372 = n2759 | n2760;
  assign n62373 = n2767 | n2768;
  assign n62374 = n2769 | n2770;
  assign n62375 = n2774 | n2775;
  assign n62376 = n2776 | n2777;
  assign n62377 = n2782 | n2778 | n2781;
  assign n62378 = n2779 | n2780;
  assign n62379 = n2784 | n2785;
  assign n62380 = n2786 | n2790 | n2796 | n2797;
  assign n62381 = n2788 | n2789;
  assign n62382 = n2791 | n2792;
  assign n62383 = n2793 | n2794;
  assign n62384 = n2819 | n2820;
  assign n62385 = n2822 | n2823;
  assign n62386 = n2832 | n2833;
  assign n62387 = n2837 | n2834 | n2836;
  assign n62388 = n2840 | n2841;
  assign n62389 = n2862 | n2863;
  assign n62390 = n2875 | n2876;
  assign n62391 = n2885 | n2886;
  assign n62392 = n2888 | n2889;
  assign n62393 = n2917 | n2918;
  assign n62394 = n2925 | n2926;
  assign n62395 = n2932 | n2928 | n2931;
  assign n62396 = n2941 | n2942;
  assign n62397 = n2949 | n2943 | n2948;
  assign n62398 = n2944 | n2945;
  assign n62399 = n2946 | n2947;
  assign n62400 = n2956 | n2957;
  assign n62401 = n2962 | n2963;
  assign n62402 = n2976 | n2977;
  assign n62403 = n2981 | n2982;
  assign n62404 = n2983 | n2984;
  assign n62405 = n2988 | n2989;
  assign n62406 = n3001 | n3002;
  assign n62407 = n3012 | n3013;
  assign n62408 = n3016 | n3017;
  assign n62409 = n3038 | n3034 | n3037;
  assign n62410 = n3053 | ~n3054;
  assign n62411 = n3064 | n3060 | ~n3063;
  assign n62412 = n3068 | n3069;
  assign n62413 = n3071 | n3072;
  assign n62414 = n3080 | n3081;
  assign n62415 = n3083 | n3084;
  assign n62416 = n3089 | n3090;
  assign n62417 = n3094 | n3095;
  assign n62418 = n3101 | n3102;
  assign n62419 = n3108 | n3109;
  assign n62420 = n3114 | n3115;
  assign n62421 = n3116 | n3117;
  assign n62422 = n3133 | n3134;
  assign n62423 = n3145 | ~n3146;
  assign n62424 = n3151 | ~n3152;
  assign n62425 = n3166 | ~n3178 | n3184 | n3185;
  assign n62426 = n3193 | ~n3194;
  assign n62427 = n3210 | n3211;
  assign n62428 = n3213 | n3214;
  assign n62429 = ~n3230 | n3220 | ~n3229;
  assign n62430 = n3236 | ~n3237;
  assign n62431 = n3243 | ~n3244;
  assign n62432 = n3250 | ~n3251;
  assign n62433 = n3253 | n3254;
  assign n62434 = n3259 | n3255 | ~n3258;
  assign n62435 = n3265 | ~n3266;
  assign n62436 = n3274 | ~n3275;
  assign n62437 = n3284 | n3280 | ~n3283;
  assign n62438 = n3292 | n3293;
  assign n62439 = n3301 | n3302;
  assign n62440 = n3307 | n3308;
  assign n62441 = n3310 | n3311;
  assign n62442 = n3323 | n3324;
  assign n62443 = n3325 | n3326;
  assign n62444 = n3367 | n3368;
  assign n62445 = n3373 | n3374;
  assign n62446 = n3379 | n3376 | n3378;
  assign n62447 = n3386 | ~n3387;
  assign n62448 = n3398 | ~n3399;
  assign n62449 = n3403 | ~n3404;
  assign n62450 = n3410 | ~n3411;
  assign n62451 = n3419 | n3420;
  assign n62452 = n3447 | n3448;
  assign n62453 = n3455 | n3456;
  assign n62454 = n3461 | n3458 | n3460;
  assign n62455 = n3477 | n3474 | n3476;
  assign n62456 = n3486 | ~n3487;
  assign n62457 = n3501 | n3510 | ~n3516 | n3517;
  assign n62458 = n3522 | ~n3523;
  assign n62459 = n3538 | n3534 | ~n3537;
  assign n62460 = n3543 | n3544;
  assign n62461 = n3552 | ~n3553;
  assign n62462 = n3567 | n3568;
  assign n62463 = n3573 | ~n3574;
  assign n62464 = n3579 | ~n3580;
  assign n62465 = n3600 | n3593 | n3599;
  assign n62466 = n3603 | ~n3606 | n3612 | n3613;
  assign n62467 = n3621 | ~n3622;
  assign n62468 = n3627 | ~n3628;
  assign n62469 = n3633 | ~n3634;
  assign n62470 = n3659 | ~n3660;
  assign n62471 = n3663 | ~n3666 | n3678 | n3679;
  assign n62472 = n3684 | ~n3685;
  assign n62473 = n3688 | n3689;
  assign n62474 = n3761 | n3725 | n3760;
  assign n62475 = n3737 | n3738;
  assign n62476 = n3743 | n3744;
  assign n62477 = n3747 | n3748;
  assign n62478 = n3753 | n3754;
  assign n62479 = n3784 | ~n3785;
  assign n62480 = n3793 | ~n3794;
  assign n62481 = n3799 | ~n3800;
  assign n62482 = n3809 | n3810;
  assign n62483 = n3817 | n3818;
  assign n62484 = n3829 | ~n3830;
  assign n62485 = n3838 | ~n3839;
  assign n62486 = n3844 | ~n3845;
  assign n62487 = n3850 | ~n3851;
  assign n62488 = n3862 | ~n3863;
  assign n62489 = n3892 | n3893;
  assign n62490 = n3894 | n3895;
  assign n62491 = n3900 | ~n3901;
  assign n62492 = n3906 | ~n3907;
  assign n62493 = n3915 | ~n3916;
  assign n62494 = n3921 | ~n3922;
  assign n62495 = n3927 | ~n3928;
  assign n62496 = n3936 | n3937;
  assign n62497 = n3951 | ~n3952;
  assign n62498 = n3956 | n3953 | n3955;
  assign n62499 = n3962 | ~n3963;
  assign n62500 = n3971 | ~n3972;
  assign n62501 = n3977 | ~n3978;
  assign n62502 = n3995 | n3996;
  assign n62503 = n4014 | ~n4015;
  assign n62504 = n4022 | n4018 | ~n4021;
  assign n62505 = n4029 | n4025 | ~n4028;
  assign n62506 = ~n4059 | n4051 | ~n4058;
  assign n62507 = n4063 | ~n4064;
  assign n62508 = n4070 | ~n4071;
  assign n62509 = n4072 | n4073;
  assign n62510 = n4079 | ~n4080;
  assign n62511 = n4081 | n4082;
  assign n62512 = n4085 | ~n4086;
  assign n62513 = n4091 | ~n4092;
  assign n62514 = ~n4107 | n4103 | ~n4106;
  assign n62515 = n4127 | n4120 | n4126;
  assign n62516 = n4130 | n4131;
  assign n62517 = n4138 | ~n4139;
  assign n62518 = n4142 | ~n4145 | n4148 | ~n4149;
  assign n62519 = n4155 | ~n4156;
  assign n62520 = n4172 | ~n4173;
  assign n62521 = n4189 | ~n4190;
  assign n62522 = n4195 | ~n4196;
  assign n62523 = ~n4203 | n4199 | ~n4202;
  assign n62524 = n4216 | ~n4217;
  assign n62525 = n4228 | ~n4229;
  assign n62526 = n4237 | ~n4238;
  assign n62527 = n4248 | ~n4249;
  assign n62528 = n4252 | ~n4253;
  assign n62529 = ~n4270 | n4266 | n4269;
  assign n62530 = n4289 | n4276 | ~n4288;
  assign n62531 = n4284 | ~n4285;
  assign n62532 = n4296 | ~n4297;
  assign n62533 = n4305 | ~n4306;
  assign n62534 = n4314 | ~n4315;
  assign n62535 = n4335 | n4347 | ~n4359 | n4360;
  assign n62536 = n4366 | n4367;
  assign n62537 = n4378 | n4376 | n4377;
  assign n62538 = n4387 | n4385 | n4386;
  assign n62539 = n4389 | ~n4390;
  assign n62540 = n4392 | n4393;
  assign n62541 = n4394 | n4395;
  assign n62542 = n4396 | n4397;
  assign n62543 = n4398 | n4399;
  assign n62544 = n4412 | n4413;
  assign n62545 = n4414 | n4415;
  assign n62546 = n4421 | ~n4422;
  assign n62547 = n4430 | n4427 | n4429;
  assign n62548 = n4436 | n4433 | n4435;
  assign n62549 = n4471 | n4452 | n4470;
  assign n62550 = n4496 | n4497;
  assign n62551 = n4511 | n4512;
  assign n62552 = n4518 | n4519;
  assign n62553 = n4525 | n4522 | n4524;
  assign n62554 = n4539 | n4540;
  assign n62555 = n4556 | ~n4557;
  assign n62556 = n4565 | ~n4566;
  assign n62557 = n4586 | n4587;
  assign n62558 = n4620 | n4601 | n4619;
  assign n62559 = n4628 | n4629;
  assign n62560 = n4630 | n4631;
  assign n62561 = n4637 | n4638;
  assign n62562 = n4639 | n4640;
  assign n62563 = n4646 | n4643 | n4645;
  assign n62564 = n4678 | n4679;
  assign n62565 = ~n4690 | n4686 | ~n4689;
  assign n62566 = n4703 | ~n4704;
  assign n62567 = n4708 | ~n4709;
  assign n62568 = n4715 | ~n4716;
  assign n62569 = n4722 | n4723;
  assign n62570 = n4730 | n4731;
  assign n62571 = n4741 | n4734 | n4740;
  assign n62572 = n4746 | ~n4747;
  assign n62573 = n4760 | n4757 | n4759;
  assign n62574 = n4767 | n4768;
  assign n62575 = n4771 | n4772;
  assign n62576 = n4777 | n4778;
  assign n62577 = n4786 | n4783 | n4785;
  assign n62578 = n4810 | n4811;
  assign n62579 = n4812 | n4813;
  assign n62580 = n4821 | n4822;
  assign n62581 = n4832 | ~n4833;
  assign n62582 = n4839 | ~n4840;
  assign n62583 = ~n4862 | n4844 | n4861;
  assign n62584 = n4851 | n4852;
  assign n62585 = n4859 | n4860;
  assign n62586 = n4868 | ~n4869;
  assign n62587 = n4873 | n4874;
  assign n62588 = n4892 | n4893;
  assign n62589 = n4900 | n4901;
  assign n62590 = n4902 | ~n4903;
  assign n62591 = ~n4913 | n4909 | n4912;
  assign n62592 = n4917 | ~n4918;
  assign n62593 = n4924 | ~n4925;
  assign n62594 = n4929 | n4930;
  assign n62595 = n4935 | n4936;
  assign n62596 = n4939 | n4940;
  assign n62597 = n4949 | n4950;
  assign n62598 = n4962 | n4957 | ~n4961;
  assign n62599 = n4972 | ~n4973;
  assign n62600 = n4981 | n4982;
  assign n62601 = n5006 | n5007;
  assign n62602 = n5018 | n5019;
  assign n62603 = n5033 | n5034;
  assign n62604 = n5042 | n5039 | n5041;
  assign n62605 = n5046 | n5047;
  assign n62606 = n5063 | n5059 | ~n5062;
  assign n62607 = n5072 | n5073;
  assign n62608 = n5104 | n5105;
  assign n62609 = n5112 | n5113;
  assign n62610 = n5118 | n5115 | n5117;
  assign n62611 = n5124 | ~n5125;
  assign n62612 = n5129 | ~n5130;
  assign n62613 = n5134 | n5135;
  assign n62614 = n5140 | n5141;
  assign n62615 = n5144 | n5145;
  assign n62616 = n5168 | n5169;
  assign n62617 = n5174 | n5175;
  assign n62618 = n5178 | n5179;
  assign n62619 = n5186 | n5187;
  assign n62620 = n5189 | n5190;
  assign n62621 = n5193 | n5194;
  assign n62622 = n5197 | n5198;
  assign n62623 = n5203 | n5204;
  assign n62624 = n5219 | n5220;
  assign n62625 = n5257 | n5258;
  assign n62626 = n5263 | n5264;
  assign n62627 = ~n5271 | n5265 | n5270;
  assign n62628 = n5272 | n5273;
  assign n62629 = n5306 | n5307;
  assign n62630 = n5308 | n5309;
  assign n62631 = n5331 | ~n5332;
  assign n62632 = n5337 | n5338;
  assign n62633 = n5342 | n5343;
  assign n62634 = n5348 | n5349;
  assign n62635 = n5366 | n5367;
  assign n62636 = n5392 | n5393;
  assign n62637 = n5398 | n5399;
  assign n62638 = n5400 | n5401;
  assign n62639 = n5415 | n5416;
  assign n62640 = n5424 | n5425;
  assign n62641 = n5432 | ~n5433;
  assign n62642 = n5441 | n5442;
  assign n62643 = n5450 | ~n5451;
  assign n62644 = n5454 | ~n5455;
  assign n62645 = n5463 | n5464;
  assign n62646 = n5474 | n5475;
  assign n62647 = n5479 | n5480;
  assign n62648 = n5498 | n5499;
  assign n62649 = n5508 | n5509;
  assign n62650 = n5516 | n5517;
  assign n62651 = n5547 | n5548;
  assign n62652 = n5550 | n5551;
  assign n62653 = n5560 | n5561;
  assign n62654 = n5562 | n5563;
  assign n62655 = n5575 | n5576;
  assign n62656 = n5577 | n5578;
  assign n62657 = n5589 | n5590;
  assign n62658 = n5627 | n5628;
  assign n62659 = n5633 | n5634;
  assign n62660 = n5637 | n5638;
  assign n62661 = n5668 | n5669;
  assign n62662 = n5676 | n5677;
  assign n62663 = n5684 | ~n5685;
  assign n62664 = n5689 | n5690;
  assign n62665 = n5695 | n5696;
  assign n62666 = n5701 | n5698 | n5700;
  assign n62667 = n5720 | ~n5721;
  assign n62668 = n5725 | n5726;
  assign n62669 = n5731 | n5732;
  assign n62670 = n5735 | n5736;
  assign n62671 = n5751 | n5752;
  assign n62672 = n5755 | n5756;
  assign n62673 = n5770 | n5786 | n5788 | n5789;
  assign n62674 = n5777 | n5778;
  assign n62675 = n5783 | n5784;
  assign n62676 = n5810 | n5811;
  assign n62677 = n5816 | n5817;
  assign n62678 = n5822 | n5823;
  assign n62679 = n5828 | n5825 | n5827;
  assign n62680 = ~n5854 | n5844 | ~n5853;
  assign n62681 = n5857 | n5858;
  assign n62682 = n5865 | n5866;
  assign n62683 = n5870 | n5871;
  assign n62684 = n5903 | n5904;
  assign n62685 = n5907 | n5908;
  assign n62686 = n5927 | n5928;
  assign n62687 = n5945 | n5946;
  assign n62688 = n5956 | ~n5957;
  assign n62689 = n5965 | ~n5966;
  assign n62690 = n5979 | n6004 | n6006 | n6007;
  assign n62691 = n5982 | ~n5983;
  assign n62692 = n5993 | n5994;
  assign n62693 = n6001 | n6002;
  assign n62694 = n6037 | n6038;
  assign n62695 = n6043 | n6044;
  assign n62696 = n6045 | ~n6046;
  assign n62697 = n6056 | n6057;
  assign n62698 = n6062 | n6063;
  assign n62699 = n6068 | n6065 | n6067;
  assign n62700 = n6079 | ~n6080;
  assign n62701 = n6093 | n6094;
  assign n62702 = n6122 | n6123;
  assign n62703 = n6128 | n6129;
  assign n62704 = n6134 | n6131 | n6133;
  assign n62705 = n6141 | n6142;
  assign n62706 = n6156 | n6157;
  assign n62707 = n6185 | n6186;
  assign n62708 = n6191 | n6192;
  assign n62709 = n6195 | n6196;
  assign n62710 = n6213 | n6258 | n6260 | n6261;
  assign n62711 = n6228 | n6229;
  assign n62712 = n6236 | n6237;
  assign n62713 = n6244 | ~n6245;
  assign n62714 = n6249 | n6250;
  assign n62715 = n6255 | n6256;
  assign n62716 = n6271 | n6272;
  assign n62717 = n6285 | n6286;
  assign n62718 = n6305 | n6302 | n6304;
  assign n62719 = n6311 | ~n6312;
  assign n62720 = n6315 | n6316;
  assign n62721 = n6325 | n6326;
  assign n62722 = n6336 | n6337;
  assign n62723 = n6391 | n6392;
  assign n62724 = n6397 | n6398;
  assign n62725 = n6403 | n6400 | n6402;
  assign n62726 = n6408 | n6409;
  assign n62727 = n6414 | n6411 | n6413;
  assign n62728 = n6416 | n6417;
  assign n62729 = n6438 | n6439;
  assign n62730 = n6444 | n6445;
  assign n62731 = n6446 | ~n6447;
  assign n62732 = n6457 | n6458;
  assign n62733 = n6463 | n6464;
  assign n62734 = n6469 | n6466 | n6468;
  assign n62735 = n6480 | ~n6481;
  assign n62736 = n6491 | n6492;
  assign n62737 = n6520 | n6521;
  assign n62738 = n6526 | n6527;
  assign n62739 = n6532 | n6529 | n6531;
  assign n62740 = n6539 | n6540;
  assign n62741 = n6544 | n6545;
  assign n62742 = n6567 | n6568;
  assign n62743 = n6569 | n6570;
  assign n62744 = n6583 | n6580 | n6582;
  assign n62745 = n6603 | n6604;
  assign n62746 = n6609 | n6610;
  assign n62747 = n6613 | n6614;
  assign n62748 = n6618 | n6619;
  assign n62749 = n6648 | ~n6649;
  assign n62750 = n6656 | n6657;
  assign n62751 = n6661 | n6662;
  assign n62752 = n6663 | n6664;
  assign n62753 = n6668 | n6669;
  assign n62754 = n6674 | n6675;
  assign n62755 = n6680 | n6677 | n6679;
  assign n62756 = n6684 | n6685;
  assign n62757 = ~n6712 | n6694 | ~n6711;
  assign n62758 = n6701 | n6702;
  assign n62759 = n6709 | n6710;
  assign n62760 = ~n6722 | n6718 | n6721;
  assign n62761 = n6735 | ~n6736;
  assign n62762 = n6755 | n6771 | n6773 | n6774;
  assign n62763 = n6762 | n6763;
  assign n62764 = n6768 | n6769;
  assign n62765 = n6798 | n6799;
  assign n62766 = n6816 | n6817;
  assign n62767 = n6825 | n6826;
  assign n62768 = n6836 | n6827 | n6835;
  assign n62769 = n6834 | n6828 | n6833;
  assign n62770 = n6830 | n6831;
  assign n62771 = n6850 | n6851;
  assign n62772 = n6856 | n6857;
  assign n62773 = n6871 | n6872;
  assign n62774 = n6881 | n6882;
  assign n62775 = n6887 | n6888;
  assign n62776 = n6900 | n6901;
  assign n62777 = n6914 | n6915;
  assign n62778 = n6917 | n6918;
  assign n62779 = n6922 | n6923;
  assign n62780 = n6927 | n6928;
  assign n62781 = n6944 | ~n6945;
  assign n62782 = n6983 | n6984;
  assign n62783 = n6985 | n6986;
  assign n62784 = n7026 | ~n7027;
  assign n62785 = n7031 | ~n7032;
  assign n62786 = n7062 | ~n7063;
  assign n62787 = n7071 | n7072;
  assign n62788 = n7090 | n7091;
  assign n62789 = n7108 | ~n7109;
  assign n62790 = n7112 | n7113;
  assign n62791 = n7131 | n7132;
  assign n62792 = n7147 | ~n7148;
  assign n62793 = n7173 | ~n7174;
  assign n62794 = n7209 | n7206 | n7208;
  assign n62795 = n7210 | n7211;
  assign n62796 = n7231 | n7232;
  assign n62797 = n7243 | ~n7244;
  assign n62798 = n7255 | n7252 | n7254;
  assign n62799 = n7256 | n7257;
  assign n62800 = n7270 | ~n7271;
  assign n62801 = n7275 | ~n7276;
  assign n62802 = n7280 | ~n7281;
  assign n62803 = n7303 | ~n7304;
  assign n62804 = n7308 | ~n7309;
  assign n62805 = n7313 | n7314;
  assign n62806 = n7319 | n7317 | n7318;
  assign n62807 = n7335 | n7333 | n7334;
  assign n62808 = n7341 | n7342;
  assign n62809 = n7416 | n7417;
  assign n62810 = n7419 | n7420;
  assign n62811 = n7422 | n7423;
  assign n62812 = n7434 | n7435;
  assign n62813 = n7459 | n7460;
  assign n62814 = n7470 | ~n7471;
  assign n62815 = n7478 | ~n7479;
  assign n62816 = n7480 | n7481;
  assign n62817 = n7484 | n7485;
  assign n62818 = n7487 | n7488;
  assign n62819 = n7490 | n7491;
  assign n62820 = n7502 | ~n7503;
  assign n62821 = n7507 | ~n7508;
  assign n62822 = n7512 | ~n7513;
  assign n62823 = n7521 | ~n7522;
  assign n62824 = n7529 | n7530;
  assign n62825 = n7535 | n7536;
  assign n62826 = n7545 | n7546;
  assign n62827 = n7570 | n7566 | n7569;
  assign n62828 = n7567 | n7568;
  assign n62829 = n7573 | n7571 | n7572;
  assign n62830 = n7580 | n7581;
  assign n62831 = n7599 | n7588 | n7598;
  assign n62832 = n7595 | ~n7596;
  assign n62833 = n7607 | n7608;
  assign n62834 = n7617 | n7618;
  assign n62835 = n7621 | n7622;
  assign n62836 = n7628 | n7629;
  assign n62837 = n7646 | n7647;
  assign n62838 = n7661 | n7662;
  assign n62839 = n7671 | n7672;
  assign n62840 = n7673 | n7674;
  assign n62841 = n7721 | n7722;
  assign n62842 = n7730 | n7728 | n7729;
  assign n62843 = n7740 | ~n7741;
  assign n62844 = n7742 | n7743;
  assign n62845 = n7765 | n7766;
  assign n62846 = n7775 | ~n7776;
  assign n62847 = n7783 | ~n7784;
  assign n62848 = n7785 | n7786;
  assign n62849 = n7794 | n7795;
  assign n62850 = n7804 | ~n7805;
  assign n62851 = n7809 | ~n7810;
  assign n62852 = n7859 | n7860;
  assign n62853 = n7870 | n7871;
  assign n62854 = n7883 | n7884;
  assign n62855 = n7886 | n7887;
  assign n62856 = n7894 | n7891 | n7893;
  assign n62857 = n7899 | n7900;
  assign n62858 = n7911 | n7912;
  assign n62859 = n7914 | n7915;
  assign n62860 = n7918 | n7919;
  assign n62861 = n7924 | n7925;
  assign n62862 = n7953 | n7954;
  assign n62863 = n7960 | n7961;
  assign n62864 = n7969 | n7970;
  assign n62865 = n7977 | ~n7978;
  assign n62866 = n7984 | n7985;
  assign n62867 = n7992 | n7993;
  assign n62868 = n8000 | ~n8001;
  assign n62869 = n8005 | ~n8006;
  assign n62870 = n8026 | n8027;
  assign n62871 = n8046 | n8047;
  assign n62872 = n8049 | n8050;
  assign n62873 = n8054 | n8055;
  assign n62874 = n8062 | ~n8063;
  assign n62875 = n8070 | n8071;
  assign n62876 = n8080 | n8077 | n8079;
  assign n62877 = n8082 | n8083;
  assign n62878 = n8101 | n8102;
  assign n62879 = n8122 | ~n8123;
  assign n62880 = n8169 | n8166 | n8168;
  assign n62881 = n8174 | ~n8175;
  assign n62882 = n8215 | n8212 | n8214;
  assign n62883 = n8220 | ~n8221;
  assign n62884 = n8255 | ~n8256;
  assign n62885 = n8262 | ~n8263;
  assign n62886 = n8308 | ~n8309;
  assign n62887 = n8381 | ~n8382;
  assign n62888 = n8401 | n8402;
  assign n62889 = n8465 | ~n8466;
  assign n62890 = n8471 | ~n8472;
  assign n62891 = n8476 | ~n8477;
  assign n62892 = n8507 | n8504 | n8506;
  assign n62893 = n8591 | n8592;
  assign n62894 = n8596 | ~n8597;
  assign n62895 = n8640 | n8621 | n8639;
  assign n62896 = n8649 | ~n8650;
  assign n62897 = n8662 | n8663;
  assign n62898 = n8675 | ~n8676;
  assign n62899 = n8690 | n8691;
  assign n62900 = n8748 | n8749;
  assign n62901 = n8773 | n8774;
  assign n62902 = n8782 | n8783;
  assign n62903 = n8785 | n8786;
  assign n62904 = n8787 | n8788;
  assign n62905 = n8789 | n8790 | n8791 | n8792;
  assign n62906 = n8799 | n8800;
  assign n62907 = n8840 | n8841;
  assign n62908 = n8845 | ~n8846;
  assign n62909 = n8881 | ~n8882;
  assign n62910 = n8917 | ~n8918;
  assign n62911 = n8952 | ~n8953;
  assign n62912 = n8992 | ~n8993;
  assign n62913 = n9057 | ~n9058;
  assign n62914 = n9077 | n9078;
  assign n62915 = n9128 | ~n9129;
  assign n62916 = n9134 | ~n9135;
  assign n62917 = n9139 | ~n9140;
  assign n62918 = n9235 | n9236;
  assign n62919 = n9273 | n9274;
  assign n62920 = n9286 | n9287;
  assign n62921 = n9299 | ~n9300;
  assign n62922 = n9313 | n9314;
  assign n62923 = n9342 | n9343;
  assign n62924 = n9356 | ~n9357;
  assign n62925 = n9368 | ~n9369;
  assign n62926 = n9373 | ~n9374;
  assign n62927 = n9392 | ~n9393;
  assign n62928 = n9404 | ~n9405;
  assign n62929 = n9410 | n9411;
  assign n62930 = n9426 | ~n9427;
  assign n62931 = n9439 | n9440;
  assign n62932 = n9449 | ~n9450;
  assign n62933 = n9461 | ~n9462;
  assign n62934 = n9468 | n9469;
  assign n62935 = n9482 | ~n9483;
  assign n62936 = n9493 | ~n9494;
  assign n62937 = n9498 | ~n9499;
  assign n62938 = n9520 | n9521;
  assign n62939 = n9561 | n9562;
  assign n62940 = n9564 | n9565;
  assign n62941 = n9569 | ~n9570;
  assign n62942 = n9590 | n9591;
  assign n62943 = n9594 | n9592 | n9593;
  assign n62944 = n9612 | n9613;
  assign n62945 = n9653 | ~n9654;
  assign n62946 = n9664 | ~n9665;
  assign n62947 = n9669 | n9670;
  assign n62948 = n9684 | ~n9685;
  assign n62949 = n9712 | n9713;
  assign n62950 = n9718 | n9719;
  assign n62951 = n9736 | n9737;
  assign n62952 = n9741 | n9739 | n9740;
  assign n62953 = ~n9754 | n9752 | ~n9753;
  assign n62954 = n9772 | n9773;
  assign n62955 = n9780 | n9781;
  assign n62956 = n9837 | ~n9838;
  assign n62957 = n9873 | ~n9874;
  assign n62958 = n9908 | ~n9909;
  assign n62959 = n9948 | ~n9949;
  assign n62960 = n9975 | ~n9976;
  assign n62961 = n10016 | ~n10017;
  assign n62962 = n10036 | n10037;
  assign n62963 = n10094 | ~n10095;
  assign n62964 = n10103 | n10104;
  assign n62965 = n10110 | n10111;
  assign n62966 = n10112 | n10113;
  assign n62967 = ~n10160 | n10158 | n10159;
  assign n62968 = n10190 | n10191;
  assign n62969 = n10201 | ~n10202;
  assign n62970 = n10208 | n10209;
  assign n62971 = n10240 | ~n10241;
  assign n62972 = n10246 | ~n10247;
  assign n62973 = n10253 | ~n10254;
  assign n62974 = n10289 | ~n10290;
  assign n62975 = n10295 | ~n10296;
  assign n62976 = n10308 | ~n10309;
  assign n62977 = n10337 | n10338;
  assign n62978 = n10371 | n10372;
  assign n62979 = n10373 | ~n10374;
  assign n62980 = n10378 | n10375 | ~n10377;
  assign n62981 = n10386 | n10387;
  assign n62982 = n10406 | n10407;
  assign n62983 = n10432 | ~n10433;
  assign n62984 = n10468 | ~n10469;
  assign n62985 = n10504 | ~n10505;
  assign n62986 = n10539 | ~n10540;
  assign n62987 = n10579 | ~n10580;
  assign n62988 = n10644 | ~n10645;
  assign n62989 = n10664 | n10665;
  assign n62990 = n10715 | ~n10716;
  assign n62991 = n10721 | ~n10722;
  assign n62992 = n10726 | ~n10727;
  assign n62993 = n10822 | n10823;
  assign n62994 = n10860 | n10861;
  assign n62995 = n10873 | n10874;
  assign n62996 = n10886 | ~n10887;
  assign n62997 = n10900 | n10901;
  assign n62998 = n10944 | n10945;
  assign n62999 = n10962 | n10963;
  assign n63000 = n10978 | n10979;
  assign n63001 = n10995 | n10996;
  assign n63002 = n11010 | ~n11011;
  assign n63003 = n11044 | ~n11045;
  assign n63004 = n11071 | ~n11072;
  assign n63005 = n11105 | ~n11106;
  assign n63006 = n11140 | ~n11141;
  assign n63007 = n11180 | ~n11181;
  assign n63008 = n11245 | ~n11246;
  assign n63009 = n11265 | n11266;
  assign n63010 = n11291 | n11292;
  assign n63011 = n11299 | n11300;
  assign n63012 = n11311 | n11312;
  assign n63013 = n11315 | n11316;
  assign n63014 = n11330 | n11331;
  assign n63015 = n11332 | n11333;
  assign n63016 = n11334 | n11335;
  assign n63017 = n11342 | n11343;
  assign n63018 = n11373 | n11374;
  assign n63019 = n11381 | n11382;
  assign n63020 = n11418 | ~n11419;
  assign n63021 = ~n11433 | n11424 | n11432;
  assign n63022 = n11426 | n11427;
  assign n63023 = n11429 | n11430;
  assign n63024 = n11439 | n11440;
  assign n63025 = n11448 | n11449;
  assign n63026 = n11475 | n11476;
  assign n63027 = n11479 | n11480;
  assign n63028 = n11483 | n11484;
  assign n63029 = n11486 | n11487;
  assign n63030 = n11492 | n11489 | n11491;
  assign n63031 = n11494 | ~n11495;
  assign n63032 = n11510 | n11511;
  assign n63033 = n11519 | n11520;
  assign n63034 = n11534 | n11535;
  assign n63035 = n11545 | ~n11546;
  assign n63036 = n11554 | ~n11555;
  assign n63037 = n11559 | n11560;
  assign n63038 = n11596 | n11597;
  assign n63039 = n11629 | ~n11630;
  assign n63040 = n11635 | ~n11636;
  assign n63041 = n11640 | ~n11641;
  assign n63042 = n11663 | n11664;
  assign n63043 = n11674 | ~n11675;
  assign n63044 = n11680 | ~n11681;
  assign n63045 = n11706 | n11699 | ~n11705;
  assign n63046 = n11711 | ~n11712;
  assign n63047 = n11758 | ~n11759;
  assign n63048 = n11764 | ~n11765;
  assign n63049 = n11776 | ~n11777;
  assign n63050 = n11782 | ~n11783;
  assign n63051 = n11791 | ~n11792;
  assign n63052 = n11805 | ~n11806;
  assign n63053 = n11841 | n11842;
  assign n63054 = n11848 | n11849;
  assign n63055 = n11939 | n11940;
  assign n63056 = n11943 | n11944;
  assign n63057 = n11947 | n11948;
  assign n63058 = n11952 | n11953;
  assign n63059 = n11954 | n11955;
  assign n63060 = n12015 | ~n12016;
  assign n63061 = n12021 | ~n12022;
  assign n63062 = n12033 | ~n12034;
  assign n63063 = n12039 | ~n12040;
  assign n63064 = n12045 | n12046;
  assign n63065 = n12151 | n12152;
  assign n63066 = n12155 | n12156;
  assign n63067 = n12176 | n12169 | n12175;
  assign n63068 = n12193 | n12194;
  assign n63069 = n12247 | ~n12248;
  assign n63070 = n12253 | ~n12254;
  assign n63071 = n12258 | ~n12259;
  assign n63072 = n12281 | n12282;
  assign n63073 = n12292 | ~n12293;
  assign n63074 = n12298 | ~n12299;
  assign n63075 = n12324 | n12317 | ~n12323;
  assign n63076 = n12329 | ~n12330;
  assign n63077 = n12376 | ~n12377;
  assign n63078 = n12382 | ~n12383;
  assign n63079 = n12394 | ~n12395;
  assign n63080 = n12400 | ~n12401;
  assign n63081 = n12409 | ~n12410;
  assign n63082 = n12451 | n12452;
  assign n63083 = n12458 | n12459;
  assign n63084 = n12549 | n12550;
  assign n63085 = n12553 | n12554;
  assign n63086 = n12557 | n12558;
  assign n63087 = n12562 | n12563;
  assign n63088 = n12564 | n12565;
  assign n63089 = n12630 | ~n12631;
  assign n63090 = n12636 | ~n12637;
  assign n63091 = n12642 | n12643;
  assign n63092 = n12737 | n12738;
  assign n63093 = n12761 | n12754 | n12760;
  assign n63094 = n12778 | n12779;
  assign n63095 = n12824 | n12825;
  assign n63096 = n12833 | ~n12834;
  assign n63097 = n12872 | ~n12873;
  assign n63098 = n12887 | n12883 | ~n12886;
  assign n63099 = n12907 | ~n12908;
  assign n63100 = n12924 | ~n12925;
  assign n63101 = n12930 | ~n12931;
  assign n63102 = n12935 | ~n12936;
  assign n63103 = n12941 | ~n12942;
  assign n63104 = n12962 | n12963;
  assign n63105 = n13007 | n13008;
  assign n63106 = n13033 | n13034;
  assign n63107 = n13042 | n13043;
  assign n63108 = n13120 | n13121;
  assign n63109 = n13149 | ~n13150;
  assign n63110 = n13184 | ~n13185;
  assign n63111 = n13201 | n13202;
  assign n63112 = n13212 | n13213;
  assign n63113 = n13221 | n13222;
  assign n63114 = n13224 | n13225;
  assign n63115 = n13236 | n13237;
  assign n63116 = n13244 | n13245;
  assign n63117 = ~n13316 | n13310 | n13315;
  assign n63118 = n13339 | n13340;
  assign n63119 = n13345 | n13346;
  assign n63120 = n13349 | n13350;
  assign n63121 = n13355 | n13356;
  assign n63122 = n13383 | n13384;
  assign n63123 = n13385 | n13386;
  assign n63124 = n13394 | n13395;
  assign n63125 = n13414 | n13415;
  assign n63126 = n13425 | n13426;
  assign n63127 = n13435 | n13436;
  assign n63128 = n13470 | n13471;
  assign n63129 = n13477 | ~n13478;
  assign n63130 = n13483 | n13484;
  assign n63131 = n13524 | n13525;
  assign n63132 = n13602 | n13603;
  assign n63133 = n13606 | n13607;
  assign n63134 = n13627 | n13620 | n13626;
  assign n63135 = n13644 | n13645;
  assign n63136 = n13733 | ~n13734;
  assign n63137 = n13739 | ~n13740;
  assign n63138 = ~n13754 | n13750 | ~n13753;
  assign n63139 = n13789 | ~n13790;
  assign n63140 = n13795 | ~n13796;
  assign n63141 = n13800 | ~n13801;
  assign n63142 = ~n13822 | n13809 | ~n13821;
  assign n63143 = ~n13839 | n13826 | n13838;
  assign n63144 = n13844 | n13845;
  assign n63145 = n13858 | n13859;
  assign n63146 = n13861 | n13862;
  assign n63147 = n13881 | n13882;
  assign n63148 = n13899 | n13900;
  assign n63149 = n13915 | n13916;
  assign n63150 = n13968 | ~n13969;
  assign n63151 = n13990 | n13991;
  assign n63152 = n13994 | n13995;
  assign n63153 = n14007 | n14008;
  assign n63154 = n14015 | n14016;
  assign n63155 = n14018 | n14019;
  assign n63156 = n14021 | n14022;
  assign n63157 = n14025 | n14026;
  assign n63158 = n14030 | n14031;
  assign n63159 = n14034 | n14035;
  assign n63160 = n14038 | n14039;
  assign n63161 = n14082 | ~n14083;
  assign n63162 = n14088 | ~n14089;
  assign n63163 = n14094 | ~n14095;
  assign n63164 = n14100 | n14101;
  assign n63165 = n14141 | n14142;
  assign n63166 = n14216 | n14217;
  assign n63167 = n14220 | n14221;
  assign n63168 = n14241 | n14234 | n14240;
  assign n63169 = n14258 | n14259;
  assign n63170 = n14337 | ~n14338;
  assign n63171 = n14343 | ~n14344;
  assign n63172 = ~n14358 | n14354 | ~n14357;
  assign n63173 = n14393 | ~n14394;
  assign n63174 = n14399 | ~n14400;
  assign n63175 = n14404 | ~n14405;
  assign n63176 = ~n14426 | n14413 | ~n14425;
  assign n63177 = ~n14443 | n14430 | n14442;
  assign n63178 = n14448 | n14449;
  assign n63179 = n14462 | n14463;
  assign n63180 = n14465 | n14466;
  assign n63181 = n14490 | n14491;
  assign n63182 = n14494 | n14495;
  assign n63183 = n14570 | n14571;
  assign n63184 = n14574 | n14575;
  assign n63185 = n14587 | n14588;
  assign n63186 = n14597 | n14598;
  assign n63187 = n14600 | n14601;
  assign n63188 = n14603 | n14604;
  assign n63189 = n14606 | n14607;
  assign n63190 = n14610 | n14611;
  assign n63191 = n14614 | n14615;
  assign n63192 = n14618 | n14619;
  assign n63193 = n14622 | n14623;
  assign n63194 = n14666 | ~n14667;
  assign n63195 = n14672 | ~n14673;
  assign n63196 = n14678 | ~n14679;
  assign n63197 = n14684 | n14685;
  assign n63198 = n14725 | n14726;
  assign n63199 = n14800 | n14801;
  assign n63200 = n14804 | n14805;
  assign n63201 = n14825 | n14818 | n14824;
  assign n63202 = n14842 | n14843;
  assign n63203 = n14897 | ~n14898;
  assign n63204 = n14903 | ~n14904;
  assign n63205 = n14914 | ~n14915;
  assign n63206 = n14923 | n14924;
  assign n63207 = n14942 | ~n14943;
  assign n63208 = n14944 | n14945;
  assign n63209 = n14964 | ~n14965;
  assign n63210 = n15017 | ~n15018;
  assign n63211 = n15036 | n15037;
  assign n63212 = n15046 | n15047;
  assign n63213 = n15068 | n15069;
  assign n63214 = n15077 | n15078;
  assign n63215 = n15098 | ~n15099;
  assign n63216 = n15130 | n15131;
  assign n63217 = n15134 | n15135;
  assign n63218 = n15138 | n15139;
  assign n63219 = n15155 | n15156;
  assign n63220 = n15159 | n15160;
  assign n63221 = n15164 | n15165;
  assign n63222 = n15213 | ~n15214;
  assign n63223 = n15235 | ~n15236;
  assign n63224 = n15243 | n15239 | ~n15242;
  assign n63225 = n15271 | n15260 | n15270;
  assign n63226 = n15266 | n15267;
  assign n63227 = n15306 | n15307;
  assign n63228 = n15312 | ~n15313;
  assign n63229 = n15318 | n15319;
  assign n63230 = n15359 | n15360;
  assign n63231 = n15439 | n15440;
  assign n63232 = n15443 | n15444;
  assign n63233 = n15464 | n15457 | n15463;
  assign n63234 = n15481 | n15482;
  assign n63235 = n15534 | ~n15535;
  assign n63236 = n15540 | ~n15541;
  assign n63237 = n15545 | ~n15546;
  assign n63238 = n15567 | ~n15568;
  assign n63239 = n15569 | n15570;
  assign n63240 = n15580 | ~n15581;
  assign n63241 = n15586 | ~n15587;
  assign n63242 = n15606 | n15607;
  assign n63243 = n15655 | ~n15656;
  assign n63244 = n15661 | ~n15662;
  assign n63245 = ~n15676 | n15672 | ~n15675;
  assign n63246 = n15723 | n15724;
  assign n63247 = n15730 | n15731;
  assign n63248 = n15820 | n15821;
  assign n63249 = n15824 | n15825;
  assign n63250 = n15837 | n15838;
  assign n63251 = n15845 | n15846;
  assign n63252 = n15847 | n15848;
  assign n63253 = n15849 | n15850;
  assign n63254 = n15855 | n15856;
  assign n63255 = n15859 | n15860;
  assign n63256 = n15863 | n15864;
  assign n63257 = n15907 | ~n15908;
  assign n63258 = n15913 | ~n15914;
  assign n63259 = n15919 | ~n15920;
  assign n63260 = n15925 | n15926;
  assign n63261 = n15966 | n15967;
  assign n63262 = n16041 | n16042;
  assign n63263 = n16045 | n16046;
  assign n63264 = n16066 | n16059 | n16065;
  assign n63265 = n16083 | n16084;
  assign n63266 = n16112 | n16113;
  assign n63267 = n16168 | ~n16169;
  assign n63268 = n16209 | ~n16210;
  assign n63269 = n16215 | ~n16216;
  assign n63270 = n16220 | ~n16221;
  assign n63271 = n16226 | ~n16227;
  assign n63272 = n16246 | ~n16247;
  assign n63273 = n16254 | n16250 | ~n16253;
  assign n63274 = n16263 | n16264;
  assign n63275 = n16274 | n16275;
  assign n63276 = n16279 | n16280;
  assign n63277 = n16284 | n16285;
  assign n63278 = n16287 | n16288;
  assign n63279 = n16312 | n16313;
  assign n63280 = n16342 | n16343;
  assign n63281 = n16345 | n16346;
  assign n63282 = n16377 | ~n16378;
  assign n63283 = n16397 | ~n16398;
  assign n63284 = n16415 | n16407 | n16414;
  assign n63285 = n16417 | n16418;
  assign n63286 = n16431 | n16432;
  assign n63287 = n16459 | ~n16460;
  assign n63288 = n16476 | ~n16477;
  assign n63289 = n16481 | n16482;
  assign n63290 = n16498 | ~n16499;
  assign n63291 = n16537 | n16526 | n16536;
  assign n63292 = n16532 | n16533;
  assign n63293 = n16570 | n16571;
  assign n63294 = n16576 | ~n16577;
  assign n63295 = n16582 | n16583;
  assign n63296 = n16623 | n16624;
  assign n63297 = n16703 | n16704;
  assign n63298 = n16707 | n16708;
  assign n63299 = n16728 | n16721 | n16727;
  assign n63300 = n16745 | n16746;
  assign n63301 = n16798 | ~n16799;
  assign n63302 = n16804 | ~n16805;
  assign n63303 = n16809 | ~n16810;
  assign n63304 = n16831 | ~n16832;
  assign n63305 = n16833 | n16834;
  assign n63306 = n16844 | ~n16845;
  assign n63307 = n16850 | ~n16851;
  assign n63308 = n16920 | ~n16921;
  assign n63309 = n16926 | ~n16927;
  assign n63310 = ~n16941 | n16937 | ~n16940;
  assign n63311 = n16975 | n16976;
  assign n63312 = n17002 | n17003;
  assign n63313 = n17009 | n17010;
  assign n63314 = n17076 | ~n17077;
  assign n63315 = n17098 | n17099;
  assign n63316 = n17102 | n17103;
  assign n63317 = n17106 | n17107;
  assign n63318 = n17111 | n17112;
  assign n63319 = n17113 | n17114;
  assign n63320 = n17115 | n17116;
  assign n63321 = n17121 | n17122;
  assign n63322 = n17125 | n17126;
  assign n63323 = n17129 | n17130;
  assign n63324 = n17165 | n17166;
  assign n63325 = n17171 | ~n17172;
  assign n63326 = n17177 | n17178;
  assign n63327 = n17218 | n17219;
  assign n63328 = n17298 | n17299;
  assign n63329 = n17302 | n17303;
  assign n63330 = n17323 | n17316 | n17322;
  assign n63331 = n17340 | n17341;
  assign n63332 = n17393 | ~n17394;
  assign n63333 = n17399 | ~n17400;
  assign n63334 = n17404 | ~n17405;
  assign n63335 = n17426 | ~n17427;
  assign n63336 = n17428 | n17429;
  assign n63337 = n17439 | ~n17440;
  assign n63338 = n17445 | ~n17446;
  assign n63339 = n17515 | ~n17516;
  assign n63340 = n17521 | ~n17522;
  assign n63341 = ~n17536 | n17532 | ~n17535;
  assign n63342 = n17570 | n17571;
  assign n63343 = n17597 | n17598;
  assign n63344 = n17604 | n17605;
  assign n63345 = n17671 | ~n17672;
  assign n63346 = n17693 | n17694;
  assign n63347 = n17697 | n17698;
  assign n63348 = n17701 | n17702;
  assign n63349 = n17706 | n17707;
  assign n63350 = n17708 | n17709;
  assign n63351 = n17710 | n17711;
  assign n63352 = n17716 | n17717;
  assign n63353 = n17720 | n17721;
  assign n63354 = n17724 | n17725;
  assign n63355 = n17760 | n17761;
  assign n63356 = n17766 | ~n17767;
  assign n63357 = n17772 | n17773;
  assign n63358 = n17813 | n17814;
  assign n63359 = n17893 | n17894;
  assign n63360 = n17897 | n17898;
  assign n63361 = n17918 | n17911 | n17917;
  assign n63362 = n17935 | n17936;
  assign n63363 = n17988 | ~n17989;
  assign n63364 = n17994 | ~n17995;
  assign n63365 = n17999 | ~n18000;
  assign n63366 = n18021 | ~n18022;
  assign n63367 = n18023 | n18024;
  assign n63368 = n18034 | ~n18035;
  assign n63369 = n18040 | ~n18041;
  assign n63370 = n18060 | n18061;
  assign n63371 = n18109 | ~n18110;
  assign n63372 = n18115 | ~n18116;
  assign n63373 = ~n18130 | n18126 | ~n18129;
  assign n63374 = n18177 | n18178;
  assign n63375 = n18184 | n18185;
  assign n63376 = n18274 | n18275;
  assign n63377 = n18278 | n18279;
  assign n63378 = n18291 | n18292;
  assign n63379 = n18299 | n18300;
  assign n63380 = n18301 | n18302;
  assign n63381 = n18303 | n18304;
  assign n63382 = n18309 | n18310;
  assign n63383 = n18313 | n18314;
  assign n63384 = n18317 | n18318;
  assign n63385 = n18353 | n18354;
  assign n63386 = n18359 | ~n18360;
  assign n63387 = n18365 | n18366;
  assign n63388 = n18406 | n18407;
  assign n63389 = n18486 | n18487;
  assign n63390 = n18490 | n18491;
  assign n63391 = n18511 | n18504 | n18510;
  assign n63392 = n18528 | n18529;
  assign n63393 = n18581 | ~n18582;
  assign n63394 = n18587 | ~n18588;
  assign n63395 = n18592 | ~n18593;
  assign n63396 = n18614 | ~n18615;
  assign n63397 = n18616 | n18617;
  assign n63398 = n18627 | ~n18628;
  assign n63399 = n18633 | ~n18634;
  assign n63400 = n18653 | n18654;
  assign n63401 = n18702 | ~n18703;
  assign n63402 = n18708 | ~n18709;
  assign n63403 = ~n18723 | n18719 | ~n18722;
  assign n63404 = n18770 | n18771;
  assign n63405 = n18777 | n18778;
  assign n63406 = n18867 | n18868;
  assign n63407 = n18871 | n18872;
  assign n63408 = n18884 | n18885;
  assign n63409 = n18892 | n18893;
  assign n63410 = n18894 | n18895;
  assign n63411 = n18896 | n18897;
  assign n63412 = n18902 | n18903;
  assign n63413 = n18906 | n18907;
  assign n63414 = n18910 | n18911;
  assign n63415 = n18946 | n18947;
  assign n63416 = n18952 | ~n18953;
  assign n63417 = n18958 | n18959;
  assign n63418 = n18999 | n19000;
  assign n63419 = n19079 | n19080;
  assign n63420 = n19083 | n19084;
  assign n63421 = n19104 | n19097 | n19103;
  assign n63422 = n19121 | n19122;
  assign n63423 = n19174 | ~n19175;
  assign n63424 = n19180 | ~n19181;
  assign n63425 = n19185 | ~n19186;
  assign n63426 = n19207 | ~n19208;
  assign n63427 = n19209 | n19210;
  assign n63428 = n19220 | ~n19221;
  assign n63429 = n19226 | ~n19227;
  assign n63430 = n19246 | n19247;
  assign n63431 = n19295 | ~n19296;
  assign n63432 = n19301 | ~n19302;
  assign n63433 = ~n19316 | n19312 | ~n19315;
  assign n63434 = n19363 | n19364;
  assign n63435 = n19370 | n19371;
  assign n63436 = n19460 | n19461;
  assign n63437 = n19464 | n19465;
  assign n63438 = n19477 | n19478;
  assign n63439 = n19485 | n19486;
  assign n63440 = n19487 | n19488;
  assign n63441 = n19489 | n19490;
  assign n63442 = n19495 | n19496;
  assign n63443 = n19499 | n19500;
  assign n63444 = n19503 | n19504;
  assign n63445 = n19539 | n19540;
  assign n63446 = n19545 | ~n19546;
  assign n63447 = n19551 | n19552;
  assign n63448 = n19592 | n19593;
  assign n63449 = n19672 | n19673;
  assign n63450 = n19676 | n19677;
  assign n63451 = n19697 | n19690 | n19696;
  assign n63452 = n19714 | n19715;
  assign n63453 = n19767 | ~n19768;
  assign n63454 = n19773 | ~n19774;
  assign n63455 = n19778 | ~n19779;
  assign n63456 = n19800 | ~n19801;
  assign n63457 = n19802 | n19803;
  assign n63458 = n19813 | ~n19814;
  assign n63459 = n19819 | ~n19820;
  assign n63460 = n19889 | ~n19890;
  assign n63461 = n19895 | ~n19896;
  assign n63462 = ~n19910 | n19906 | ~n19909;
  assign n63463 = n19944 | n19945;
  assign n63464 = n19971 | n19972;
  assign n63465 = n19978 | n19979;
  assign n63466 = n20045 | ~n20046;
  assign n63467 = n20067 | n20068;
  assign n63468 = n20071 | n20072;
  assign n63469 = n20075 | n20076;
  assign n63470 = n20080 | n20081;
  assign n63471 = n20082 | n20083;
  assign n63472 = n20084 | n20085;
  assign n63473 = n20090 | n20091;
  assign n63474 = n20094 | n20095;
  assign n63475 = n20098 | n20099;
  assign n63476 = n20142 | ~n20143;
  assign n63477 = n20148 | ~n20149;
  assign n63478 = n20154 | ~n20155;
  assign n63479 = n20160 | n20161;
  assign n63480 = n20201 | n20202;
  assign n63481 = n20276 | n20277;
  assign n63482 = n20280 | n20281;
  assign n63483 = n20301 | n20294 | n20300;
  assign n63484 = n20318 | n20319;
  assign n63485 = n20402 | ~n20403;
  assign n63486 = n20424 | n20425;
  assign n63487 = n20443 | ~n20444;
  assign n63488 = n20449 | ~n20450;
  assign n63489 = n20454 | ~n20455;
  assign n63490 = n20460 | ~n20461;
  assign n63491 = n20469 | n20470;
  assign n63492 = n20483 | ~n20484;
  assign n63493 = n20485 | n20486;
  assign n63494 = n20500 | n20501;
  assign n63495 = n20526 | n20527;
  assign n63496 = n20558 | n20559;
  assign n63497 = n20579 | ~n20580;
  assign n63498 = n20599 | ~n20600;
  assign n63499 = n20617 | n20609 | n20616;
  assign n63500 = n20619 | n20620;
  assign n63501 = n20633 | n20634;
  assign n63502 = n20638 | n20639;
  assign n63503 = n20679 | ~n20680;
  assign n63504 = n20687 | n20688;
  assign n63505 = n20703 | ~n20704;
  assign n63506 = n20711 | n20707 | ~n20710;
  assign n63507 = n20749 | n20738 | n20748;
  assign n63508 = n20744 | n20745;
  assign n63509 = n20790 | ~n20791;
  assign n63510 = n20796 | ~n20797;
  assign n63511 = n20802 | ~n20803;
  assign n63512 = n20808 | n20809;
  assign n63513 = n20849 | n20850;
  assign n63514 = n20924 | n20925;
  assign n63515 = n20928 | n20929;
  assign n63516 = n20949 | n20942 | n20948;
  assign n63517 = n20966 | n20967;
  assign n63518 = n21021 | ~n21022;
  assign n63519 = n21027 | ~n21028;
  assign n63520 = n21032 | ~n21033;
  assign n63521 = n21038 | ~n21039;
  assign n63522 = n21047 | n21048;
  assign n63523 = n21063 | n21064;
  assign n63524 = n21087 | ~n21088;
  assign n63525 = n21140 | ~n21141;
  assign n63526 = n21159 | n21160;
  assign n63527 = n21164 | n21165;
  assign n63528 = n21190 | n21191;
  assign n63529 = n21222 | n21223;
  assign n63530 = n21243 | ~n21244;
  assign n63531 = n21263 | ~n21264;
  assign n63532 = n21281 | n21273 | n21280;
  assign n63533 = n21283 | n21284;
  assign n63534 = n21297 | n21298;
  assign n63535 = n21302 | n21303;
  assign n63536 = n21343 | ~n21344;
  assign n63537 = n21347 | n21348;
  assign n63538 = n21352 | n21353;
  assign n63539 = n21368 | ~n21369;
  assign n63540 = n21376 | n21372 | ~n21375;
  assign n63541 = n21384 | n21385;
  assign n63542 = n21391 | n21392;
  assign n63543 = n21395 | n21396;
  assign n63544 = n21437 | ~n21438;
  assign n63545 = n21443 | ~n21444;
  assign n63546 = n21449 | ~n21450;
  assign n63547 = n21455 | n21456;
  assign n63548 = n21496 | n21497;
  assign n63549 = n21571 | n21572;
  assign n63550 = n21575 | n21576;
  assign n63551 = n21596 | n21589 | n21595;
  assign n63552 = n21613 | n21614;
  assign n63553 = n21668 | ~n21669;
  assign n63554 = n21674 | ~n21675;
  assign n63555 = n21679 | ~n21680;
  assign n63556 = n21685 | ~n21686;
  assign n63557 = n21694 | n21695;
  assign n63558 = n21710 | n21711;
  assign n63559 = n21734 | ~n21735;
  assign n63560 = n21787 | ~n21788;
  assign n63561 = n21806 | n21807;
  assign n63562 = n21811 | n21812;
  assign n63563 = n21837 | n21838;
  assign n63564 = n21869 | n21870;
  assign n63565 = n21890 | ~n21891;
  assign n63566 = n21910 | ~n21911;
  assign n63567 = n21928 | n21920 | n21927;
  assign n63568 = n21930 | n21931;
  assign n63569 = n21944 | n21945;
  assign n63570 = n21949 | n21950;
  assign n63571 = n21990 | ~n21991;
  assign n63572 = n21994 | n21995;
  assign n63573 = n21999 | n22000;
  assign n63574 = n22015 | ~n22016;
  assign n63575 = n22023 | n22019 | ~n22022;
  assign n63576 = n22031 | n22032;
  assign n63577 = n22038 | n22039;
  assign n63578 = n22042 | n22043;
  assign n63579 = n22068 | n22069;
  assign n63580 = n22078 | ~n22079;
  assign n63581 = n22126 | ~n22127;
  assign n63582 = n22146 | ~n22147;
  assign n63583 = n22163 | ~n22164;
  assign n63584 = n22169 | ~n22170;
  assign n63585 = n22174 | ~n22175;
  assign n63586 = n22180 | ~n22181;
  assign n63587 = n22188 | n22189;
  assign n63588 = n22197 | ~n22198;
  assign n63589 = n22203 | ~n22204;
  assign n63590 = n22212 | n22213;
  assign n63591 = n22241 | n22242;
  assign n63592 = n22254 | n22255;
  assign n63593 = n22273 | n22274;
  assign n63594 = n22299 | n22300;
  assign n63595 = n22308 | n22309;
  assign n63596 = n22358 | n22359;
  assign n63597 = n22378 | n22379;
  assign n63598 = n22434 | ~n22435;
  assign n63599 = ~n22456 | n22439 | n22455;
  assign n63600 = n22486 | n22475 | n22485;
  assign n63601 = n22481 | n22482;
  assign n63602 = n22494 | n22495;
  assign n63603 = n22497 | n22498;
  assign n63604 = n22509 | n22510;
  assign n63605 = n22517 | n22518;
  assign n63606 = ~n22586 | n22580 | n22585;
  assign n63607 = n22609 | n22610;
  assign n63608 = n22613 | n22614;
  assign n63609 = n22617 | n22618;
  assign n63610 = n22623 | n22624;
  assign n63611 = n22649 | n22650;
  assign n63612 = n22657 | n22658;
  assign n63613 = n22694 | n22695;
  assign n63614 = n22725 | n22726;
  assign n63615 = n22731 | ~n22732;
  assign n63616 = n22737 | n22738;
  assign n63617 = n22778 | n22779;
  assign n63618 = n22858 | n22859;
  assign n63619 = n22862 | n22863;
  assign n63620 = n22883 | n22876 | n22882;
  assign n63621 = n22900 | n22901;
  assign n63622 = n22989 | ~n22990;
  assign n63623 = n22995 | ~n22996;
  assign n63624 = ~n23010 | n23006 | ~n23009;
  assign n63625 = n23045 | ~n23046;
  assign n63626 = n23051 | ~n23052;
  assign n63627 = n23056 | ~n23057;
  assign n63628 = ~n23078 | n23065 | ~n23077;
  assign n63629 = ~n23095 | n23082 | n23094;
  assign n63630 = n23100 | n23101;
  assign n63631 = n23114 | n23115;
  assign n63632 = n23117 | n23118;
  assign n63633 = n23137 | n23138;
  assign n63634 = n23155 | n23156;
  assign n63635 = n23170 | n23171;
  assign n63636 = n23223 | ~n23224;
  assign n63637 = n23245 | n23246;
  assign n63638 = n23249 | n23250;
  assign n63639 = n23262 | n23263;
  assign n63640 = n23270 | n23271;
  assign n63641 = n23273 | n23274;
  assign n63642 = n23276 | n23277;
  assign n63643 = n23280 | n23281;
  assign n63644 = n23284 | n23285;
  assign n63645 = n23288 | n23289;
  assign n63646 = n23292 | n23293;
  assign n63647 = n23328 | n23329;
  assign n63648 = n23334 | ~n23335;
  assign n63649 = n23340 | n23341;
  assign n63650 = n23381 | n23382;
  assign n63651 = n23461 | n23462;
  assign n63652 = n23465 | n23466;
  assign n63653 = n23486 | n23479 | n23485;
  assign n63654 = n23503 | n23504;
  assign n63655 = n23592 | ~n23593;
  assign n63656 = n23598 | ~n23599;
  assign n63657 = ~n23613 | n23609 | ~n23612;
  assign n63658 = n23648 | ~n23649;
  assign n63659 = n23654 | ~n23655;
  assign n63660 = n23659 | ~n23660;
  assign n63661 = ~n23681 | n23668 | ~n23680;
  assign n63662 = ~n23698 | n23685 | n23697;
  assign n63663 = n23703 | n23704;
  assign n63664 = n23717 | n23718;
  assign n63665 = n23720 | n23721;
  assign n63666 = n23740 | n23741;
  assign n63667 = n23758 | n23759;
  assign n63668 = n23773 | n23774;
  assign n63669 = n23826 | ~n23827;
  assign n63670 = n23848 | n23849;
  assign n63671 = n23852 | n23853;
  assign n63672 = n23865 | n23866;
  assign n63673 = n23873 | n23874;
  assign n63674 = n23876 | n23877;
  assign n63675 = n23879 | n23880;
  assign n63676 = n23883 | n23884;
  assign n63677 = n23887 | n23888;
  assign n63678 = n23891 | n23892;
  assign n63679 = n23895 | n23896;
  assign n63680 = n23931 | n23932;
  assign n63681 = n23937 | ~n23938;
  assign n63682 = n23943 | n23944;
  assign n63683 = n23984 | n23985;
  assign n63684 = n24064 | n24065;
  assign n63685 = n24068 | n24069;
  assign n63686 = n24089 | n24082 | n24088;
  assign n63687 = n24106 | n24107;
  assign n63688 = n24195 | ~n24196;
  assign n63689 = n24201 | ~n24202;
  assign n63690 = ~n24216 | n24212 | ~n24215;
  assign n63691 = n24251 | ~n24252;
  assign n63692 = n24257 | ~n24258;
  assign n63693 = n24262 | ~n24263;
  assign n63694 = ~n24284 | n24271 | ~n24283;
  assign n63695 = ~n24301 | n24288 | n24300;
  assign n63696 = n24306 | n24307;
  assign n63697 = n24320 | n24321;
  assign n63698 = n24323 | n24324;
  assign n63699 = n24343 | n24344;
  assign n63700 = n24361 | n24362;
  assign n63701 = n24376 | n24377;
  assign n63702 = n24429 | ~n24430;
  assign n63703 = n24451 | n24452;
  assign n63704 = n24455 | n24456;
  assign n63705 = n24468 | n24469;
  assign n63706 = n24476 | n24477;
  assign n63707 = n24479 | n24480;
  assign n63708 = n24482 | n24483;
  assign n63709 = n24486 | n24487;
  assign n63710 = n24490 | n24491;
  assign n63711 = n24494 | n24495;
  assign n63712 = n24498 | n24499;
  assign n63713 = n24534 | n24535;
  assign n63714 = n24540 | ~n24541;
  assign n63715 = n24546 | n24547;
  assign n63716 = n24587 | n24588;
  assign n63717 = n24667 | n24668;
  assign n63718 = n24671 | n24672;
  assign n63719 = n24692 | n24685 | n24691;
  assign n63720 = n24709 | n24710;
  assign n63721 = n24762 | ~n24763;
  assign n63722 = n24768 | ~n24769;
  assign n63723 = n24773 | ~n24774;
  assign n63724 = n24795 | ~n24796;
  assign n63725 = n24797 | n24798;
  assign n63726 = n24808 | ~n24809;
  assign n63727 = n24814 | ~n24815;
  assign n63728 = n24877 | ~n24878;
  assign n63729 = n24883 | ~n24884;
  assign n63730 = ~n24898 | n24894 | ~n24897;
  assign n63731 = n24949 | n24950;
  assign n63732 = n24952 | n24953;
  assign n63733 = n25043 | n25044;
  assign n63734 = n25047 | n25048;
  assign n63735 = n25060 | n25061;
  assign n63736 = n25068 | n25069;
  assign n63737 = n25070 | n25071;
  assign n63738 = n25072 | n25073;
  assign n63739 = n25078 | n25079;
  assign n63740 = n25082 | n25083;
  assign n63741 = n25086 | n25087;
  assign n63742 = n25154 | ~n25155;
  assign n63743 = n25188 | ~n25189;
  assign n63744 = n25194 | ~n25195;
  assign n63745 = n25199 | ~n25200;
  assign n63746 = n25205 | ~n25206;
  assign n63747 = n25225 | ~n25226;
  assign n63748 = n25233 | n25229 | ~n25232;
  assign n63749 = n25239 | ~n25240;
  assign n63750 = n25241 | n25242;
  assign n63751 = n25251 | ~n25252;
  assign n63752 = n25253 | n25254;
  assign n63753 = n25260 | n25261;
  assign n63754 = n25265 | n25266;
  assign n63755 = n25269 | n25270;
  assign n63756 = n25274 | n25275;
  assign n63757 = n25277 | n25278;
  assign n63758 = n25302 | n25303;
  assign n63759 = n25339 | n25340;
  assign n63760 = n25343 | n25344;
  assign n63761 = n25364 | ~n25365;
  assign n63762 = n25384 | ~n25385;
  assign n63763 = n25402 | n25394 | n25401;
  assign n63764 = n25404 | n25405;
  assign n63765 = n25418 | n25419;
  assign n63766 = n25446 | ~n25447;
  assign n63767 = n25463 | ~n25464;
  assign n63768 = n25468 | n25469;
  assign n63769 = n25485 | ~n25486;
  assign n63770 = n25517 | n25490 | n25516;
  assign n63771 = n25512 | n25513;
  assign n63772 = n25557 | ~n25558;
  assign n63773 = n25563 | ~n25564;
  assign n63774 = n25569 | ~n25570;
  assign n63775 = n25575 | n25576;
  assign n63776 = n25616 | n25617;
  assign n63777 = n25691 | n25692;
  assign n63778 = n25695 | n25696;
  assign n63779 = n25716 | n25709 | n25715;
  assign n63780 = n25733 | n25734;
  assign n63781 = n25772 | n25773;
  assign n63782 = n25797 | ~n25798;
  assign n63783 = n25803 | ~n25804;
  assign n63784 = n25808 | ~n25809;
  assign n63785 = n25814 | ~n25815;
  assign n63786 = n25822 | n25823;
  assign n63787 = n25831 | ~n25832;
  assign n63788 = n25837 | ~n25838;
  assign n63789 = n25845 | n25846;
  assign n63790 = n25872 | n25873;
  assign n63791 = n25879 | ~n25880;
  assign n63792 = n25930 | ~n25931;
  assign n63793 = n25933 | n25934;
  assign n63794 = n25950 | n25951;
  assign n63795 = n25959 | n25960;
  assign n63796 = n25974 | n25975;
  assign n63797 = n25981 | n25979 | n25980;
  assign n63798 = n26036 | n26037;
  assign n63799 = n26040 | n26041;
  assign n63800 = n26044 | n26045;
  assign n63801 = n26061 | n26062;
  assign n63802 = n26101 | ~n26102;
  assign n63803 = n26118 | ~n26119;
  assign n63804 = n26123 | n26124;
  assign n63805 = n26143 | ~n26144;
  assign n63806 = n26153 | ~n26154;
  assign n63807 = n26173 | n26174;
  assign n63808 = n26178 | ~n26179;
  assign n63809 = n26180 | n26181;
  assign po356 = n26184 | ~n26185;
  assign n63811 = n26207 | n26208;
  assign n63812 = n26219 | ~n26220;
  assign n63813 = n26236 | ~n26237;
  assign n63814 = n26242 | ~n26243;
  assign n63815 = n26247 | ~n26248;
  assign n63816 = n26292 | n26293;
  assign n63817 = n26299 | ~n26300;
  assign n63818 = n26338 | ~n26339;
  assign n63819 = ~n26353 | n26349 | ~n26352;
  assign n63820 = n26370 | n26371;
  assign n63821 = n26374 | n26375;
  assign n63822 = n26382 | n26383;
  assign n63823 = n26403 | n26404;
  assign n63824 = n26409 | n26410;
  assign n63825 = n26415 | ~n26416;
  assign n63826 = n26426 | n26427;
  assign n63827 = n26434 | n26435;
  assign n63828 = n26501 | n26502;
  assign n63829 = n26505 | n26506;
  assign n63830 = n26518 | n26519;
  assign n63831 = n26550 | ~n26551;
  assign po357 = n26555 | ~n26556;
  assign n63833 = n26574 | ~n26575;
  assign n63834 = n26580 | ~n26581;
  assign n63835 = n26585 | ~n26586;
  assign n63836 = n26591 | ~n26592;
  assign n63837 = n26597 | ~n26598;
  assign n63838 = n26603 | n26604;
  assign n63839 = n26662 | ~n26663;
  assign n63840 = n26682 | n26683;
  assign n63841 = n26689 | n26690;
  assign n63842 = n26710 | n26711;
  assign n63843 = n26753 | n26754;
  assign n63844 = n26764 | n26765;
  assign n63845 = n26802 | n26803;
  assign n63846 = n26804 | n26805;
  assign n63847 = n26813 | n26814;
  assign n63848 = n26818 | n26819;
  assign n63849 = n26837 | n26838;
  assign n63850 = n26852 | n26853;
  assign n63851 = n26869 | n26870;
  assign n63852 = n26873 | n26874;
  assign n63853 = n26894 | n26895;
  assign n63854 = n26898 | n26899;
  assign n63855 = n26910 | n26911;
  assign n63856 = n26927 | n26928;
  assign n63857 = n26934 | n26935;
  assign n63858 = n26939 | n26940;
  assign n63859 = n26974 | ~n26975;
  assign n63860 = n26989 | n26990;
  assign n63861 = n26993 | n26994;
  assign n63862 = n26996 | n26997;
  assign n63863 = n27001 | n27002;
  assign n63864 = n27006 | n27007;
  assign n63865 = n27026 | n27027;
  assign n63866 = n27062 | n27063;
  assign n63867 = n27068 | n27069;
  assign n63868 = n27072 | n27073;
  assign n63869 = n27088 | n27086 | n27087;
  assign n63870 = n27091 | ~n27092;
  assign n63871 = n27098 | n27099;
  assign n63872 = n27118 | n27119;
  assign n63873 = n27128 | n27129;
  assign n63874 = n27140 | n27141;
  assign n63875 = n27164 | ~n27165;
  assign n63876 = n27188 | n27189;
  assign n63877 = n27190 | ~n27191;
  assign po364 = n27196 | ~n27197;
  assign n63879 = n27221 | n27222;
  assign n63880 = n27228 | n27229;
  assign n63881 = n27257 | ~n27258;
  assign n63882 = n27281 | n27282;
  assign n63883 = n27283 | ~n27284;
  assign po365 = n27289 | ~n27290;
  assign n63885 = n27300 | n27301;
  assign n63886 = n27306 | n27307;
  assign n63887 = n27317 | ~n27318;
  assign n63888 = n27339 | n27340;
  assign n63889 = n27341 | n27342;
  assign n63890 = n27351 | n27352;
  assign n63891 = n27361 | ~n27362;
  assign n63892 = n27367 | ~n27368;
  assign n63893 = n27378 | ~n27379;
  assign n63894 = n27393 | n27394;
  assign n63895 = n27403 | n27404;
  assign n63896 = n27435 | n27436;
  assign n63897 = n27456 | n27457;
  assign n63898 = n27465 | n27466;
  assign n63899 = n27474 | n27475;
  assign n63900 = n27482 | n27483;
  assign n63901 = n27502 | n27503;
  assign n63902 = n27506 | n27507;
  assign n63903 = n27512 | n27513;
  assign n63904 = n27519 | n27520;
  assign n63905 = n27564 | n27565;
  assign n63906 = n27584 | n27585;
  assign n63907 = n27588 | n27589;
  assign n63908 = n27652 | n27653;
  assign n63909 = n27681 | n27682;
  assign n63910 = n27690 | ~n27691;
  assign n63911 = n27755 | ~n27756;
  assign n63912 = n27760 | ~n27761;
  assign n63913 = n27799 | n27800;
  assign n63914 = n27804 | n27805;
  assign n63915 = n27807 | n27808;
  assign n63916 = n27819 | n27820;
  assign n63917 = n27837 | n27838;
  assign n63918 = n27845 | n27846;
  assign n63919 = n27847 | n27848;
  assign n63920 = n27855 | n27856;
  assign n63921 = n27865 | n27866;
  assign n63922 = n27876 | n27877;
  assign n63923 = n27911 | ~n27912;
  assign n63924 = n27916 | ~n27917;
  assign n63925 = n27925 | n27926;
  assign n63926 = n27927 | n27928;
  assign n63927 = n27950 | n27951;
  assign n63928 = n27961 | n27962;
  assign n63929 = n27993 | n27994;
  assign n63930 = n28042 | n28043;
  assign n63931 = n28074 | n28075;
  assign n63932 = n28080 | ~n28081;
  assign n63933 = n28092 | n28093;
  assign n63934 = n28116 | n28117;
  assign n63935 = n28204 | n28205;
  assign n63936 = n28208 | n28209;
  assign n63937 = n28234 | n28235;
  assign n63938 = n28238 | n28239;
  assign n63939 = n28243 | n28244;
  assign n63940 = n28259 | ~n28260;
  assign n63941 = n28292 | n28293;
  assign n63942 = n28294 | n28295;
  assign n63943 = n28296 | n28297;
  assign n63944 = n28339 | ~n28340;
  assign n63945 = n28345 | n28346;
  assign n63946 = n28372 | n28373;
  assign n63947 = n28375 | n28376;
  assign n63948 = n28378 | n28379;
  assign n63949 = n28394 | n28395;
  assign n63950 = n28408 | n28409;
  assign n63951 = n28416 | n28417;
  assign n63952 = n28423 | n28424;
  assign n63953 = n28430 | n28431;
  assign n63954 = n28449 | ~n28450;
  assign n63955 = n28487 | ~n28488;
  assign n63956 = n28493 | ~n28494;
  assign n63957 = n28507 | n28508;
  assign n63958 = n28515 | n28516;
  assign n63959 = n28519 | n28520;
  assign n63960 = n28529 | n28530;
  assign n63961 = n28546 | n28547;
  assign n63962 = n28548 | n28549;
  assign n63963 = n28581 | n28582;
  assign n63964 = n28622 | ~n28623;
  assign n63965 = n28628 | ~n28629;
  assign n63966 = n28656 | n28657;
  assign n63967 = n28678 | ~n28679;
  assign n63968 = n28686 | ~n28687;
  assign n63969 = n28697 | n28698;
  assign n63970 = n28700 | n28701;
  assign n63971 = n28732 | n28733;
  assign n63972 = n28740 | n28741;
  assign n63973 = n28766 | n28767;
  assign n63974 = n28770 | n28771;
  assign n63975 = n28779 | n28780;
  assign n63976 = n28786 | n28787;
  assign n63977 = n28809 | n28810;
  assign n63978 = n28814 | ~n28815;
  assign n63979 = n28823 | n28824;
  assign n63980 = n28879 | n28885 | n28887 | n28888;
  assign n63981 = n28973 | n28974;
  assign n63982 = n28988 | n28989;
  assign n63983 = n28994 | n28995;
  assign n63984 = n29001 | n29002;
  assign n63985 = n29011 | n29012;
  assign n63986 = n29019 | n29020;
  assign n63987 = n29025 | n29026;
  assign n63988 = n29040 | n29041;
  assign n63989 = n29060 | n29061;
  assign po379 = n29084 | ~n29085;
  assign n63991 = n29108 | n29109;
  assign n63992 = n29160 | n29161;
  assign n63993 = n29206 | n29207;
  assign n63994 = n29223 | n29224;
  assign n63995 = n29238 | n29239;
  assign n63996 = n29252 | ~n29253;
  assign n63997 = n29290 | ~n29291;
  assign n63998 = n29296 | ~n29297;
  assign n63999 = n29301 | n29302;
  assign n64000 = n29311 | n29312;
  assign n64001 = n29324 | n29325;
  assign n64002 = n29332 | n29333;
  assign n64003 = n29336 | n29337;
  assign n64004 = n29338 | n29339;
  assign n64005 = n29355 | n29356;
  assign n64006 = n29381 | n29382;
  assign n64007 = n29388 | n29389;
  assign n64008 = n29391 | n29392;
  assign n64009 = n29407 | n29408;
  assign n64010 = n29427 | ~n29428;
  assign n64011 = n29433 | ~n29434;
  assign n64012 = n29442 | ~n29443;
  assign n64013 = n29460 | n29461;
  assign n64014 = n29466 | ~n29467;
  assign n64015 = n29493 | n29494;
  assign n64016 = n29508 | n29509;
  assign n64017 = n29512 | n29513;
  assign n64018 = n29540 | n29541;
  assign n64019 = n29547 | n29548;
  assign n64020 = n29564 | n29565;
  assign n64021 = n29578 | n29579;
  assign n64022 = n29584 | n29585;
  assign n64023 = n29592 | n29593;
  assign n64024 = n29596 | n29597;
  assign n64025 = n29616 | n29617;
  assign n64026 = n29634 | n29635;
  assign n64027 = n29642 | n29643;
  assign n64028 = n29652 | n29653;
  assign n64029 = n29670 | n29671;
  assign n64030 = n29672 | n29673;
  assign n64031 = n29677 | n29678;
  assign n64032 = n29683 | n29684;
  assign n64033 = n29764 | n29765;
  assign n64034 = n29768 | n29769;
  assign n64035 = n29782 | n29783;
  assign n64036 = ~n29824 | n29795 | ~n29823;
  assign n64037 = n29829 | ~n29830;
  assign n64038 = n29856 | n29857;
  assign n64039 = n29870 | n29871;
  assign n64040 = n29891 | n29892;
  assign n64041 = n29905 | n29906;
  assign n64042 = n29933 | n29934;
  assign n64043 = n29939 | n29940;
  assign n64044 = n29948 | n29949;
  assign n64045 = n29963 | n29964;
  assign n64046 = n29969 | n29970;
  assign n64047 = n29979 | ~n29980;
  assign n64048 = n30017 | ~n30018;
  assign n64049 = n30023 | ~n30024;
  assign n64050 = n30043 | n30044;
  assign n64051 = n30051 | n30052;
  assign n64052 = n30055 | n30056;
  assign n64053 = n30057 | n30058;
  assign n64054 = n30075 | n30076;
  assign n64055 = n30105 | n30106;
  assign n64056 = n30145 | ~n30146;
  assign n64057 = n30151 | ~n30152;
  assign n64058 = n30160 | ~n30161;
  assign n64059 = n30193 | ~n30194;
  assign n64060 = n30225 | n30226;
  assign n64061 = n30258 | n30259;
  assign n64062 = n30268 | n30265 | n30267;
  assign n64063 = n30287 | n30288;
  assign n64064 = n30301 | n30302;
  assign n64065 = n30315 | n30316;
  assign n64066 = n30322 | n30323;
  assign n64067 = n30332 | ~n30333;
  assign n64068 = n30346 | n30347;
  assign n64069 = n30349 | n30350;
  assign n64070 = n30363 | n30364;
  assign n64071 = n30368 | n30369;
  assign n64072 = n30371 | n30372;
  assign n64073 = n30378 | n30379;
  assign n64074 = n30387 | n30388;
  assign n64075 = n30393 | n30394;
  assign n64076 = n30496 | n30493 | n30495;
  assign n64077 = n30513 | n30514;
  assign n64078 = n30526 | n30527;
  assign n64079 = n30544 | n30545;
  assign n64080 = n30565 | n30566;
  assign n64081 = n30575 | n30573 | n30574;
  assign n64082 = n30581 | n30576 | n30577 | n30582 | n30583;
  assign n64083 = n30580 | n30578 | n30579;
  assign n64084 = n30585 | n30586;
  assign n64085 = n30587 | n30588;
  assign n64086 = n30593 | n30594;
  assign n64087 = n30596 | n30597;
  assign n64088 = n30601 | n30602;
  assign n64089 = n30615 | n30616;
  assign n64090 = n30622 | n30623;
  assign n64091 = n30632 | n30633;
  assign n64092 = n30636 | n30634 | n30635;
  assign n64093 = n30643 | n30644;
  assign n64094 = n30656 | n30657;
  assign n64095 = n30701 | n30702;
  assign n64096 = n30792 | n30793;
  assign n64097 = n30806 | ~n30807;
  assign n64098 = n30809 | n30810;
  assign n64099 = n30815 | n30816;
  assign n64100 = n30828 | ~n30829;
  assign n64101 = n30837 | ~n30838;
  assign n64102 = n30843 | n30840 | n30842;
  assign n64103 = n30845 | n30846;
  assign n64104 = n30847 | n30848;
  assign n64105 = n30865 | ~n30866;
  assign n64106 = n30879 | ~n30880;
  assign n64107 = n30882 | n30883;
  assign n64108 = n30888 | n30889;
  assign n64109 = n30902 | n30900 | n30901;
  assign n64110 = n30923 | n30924;
  assign n64111 = n30926 | ~n30927;
  assign n64112 = n30966 | n30967;
  assign n64113 = n30979 | n30980;
  assign n64114 = n30988 | n30989;
  assign n64115 = n30995 | n30996;
  assign n64116 = n31039 | n31040;
  assign n64117 = n31080 | n31081;
  assign n64118 = n31092 | n31088 | n31091;
  assign n64119 = n31093 | n31094;
  assign n64120 = n31127 | n31128;
  assign n64121 = n31136 | n31137;
  assign n64122 = n31140 | n31141;
  assign n64123 = n31146 | n31147;
  assign n64124 = n31157 | n31158;
  assign n64125 = n31166 | n31167;
  assign n64126 = n31170 | n31171;
  assign n64127 = n31226 | n31227;
  assign n64128 = n31229 | n31230;
  assign n64129 = n31236 | n31237;
  assign n64130 = n31239 | n31240;
  assign n64131 = n31249 | n31250;
  assign n64132 = n31252 | n31253;
  assign n64133 = n31298 | n31299;
  assign n64134 = n31306 | n31302 | n31305;
  assign n64135 = n31310 | n31311;
  assign n64136 = n31317 | n31318;
  assign n64137 = n31340 | n31341;
  assign n64138 = n31363 | n31364;
  assign n64139 = n31367 | n31368;
  assign n64140 = n31378 | n31379;
  assign n64141 = n31404 | n31405;
  assign n64142 = n31423 | ~n31424;
  assign n64143 = n31427 | n31428;
  assign n64144 = n31459 | n31460;
  assign n64145 = n31463 | n31464;
  assign n64146 = n31470 | n31471;
  assign n64147 = n31478 | n31475 | n31477;
  assign n64148 = n31515 | ~n31516;
  assign n64149 = n31605 | n31606;
  assign n64150 = n31634 | n31635;
  assign n64151 = n31659 | n31660;
  assign n64152 = n31685 | n31686;
  assign n64153 = n31728 | n31729;
  assign n64154 = n31752 | n31753;
  assign n64155 = n31759 | n31760;
  assign n64156 = n31771 | n31772;
  assign n64157 = n31780 | n31781;
  assign n64158 = n31791 | n31792;
  assign n64159 = n31799 | n31800;
  assign n64160 = n31818 | n31819;
  assign n64161 = n31861 | n31862;
  assign n64162 = n31870 | n31871;
  assign n64163 = n31874 | n31875;
  assign n64164 = n31878 | n31879;
  assign n64165 = n31880 | n31881;
  assign n64166 = n31924 | ~n31925;
  assign n64167 = n31932 | ~n31933;
  assign n64168 = n31950 | n31951;
  assign n64169 = n31957 | n31958;
  assign n64170 = n31972 | n31973;
  assign n64171 = n31974 | n31975;
  assign n64172 = n31991 | n31992;
  assign n64173 = n32000 | n32001;
  assign n64174 = n32002 | n32003;
  assign n64175 = n32011 | ~n32012;
  assign n64176 = n32021 | n32022;
  assign n64177 = n32025 | ~n32026;
  assign n64178 = n32063 | n32064;
  assign n64179 = n32084 | n32081 | n32083;
  assign n64180 = n32125 | n32126;
  assign n64181 = n32139 | n32140;
  assign n64182 = n32149 | n32150;
  assign n64183 = n32190 | n32191;
  assign n64184 = n32194 | n32195;
  assign n64185 = n32197 | n32198;
  assign n64186 = n32201 | n32202;
  assign n64187 = n32207 | n32208;
  assign n64188 = n32212 | n32213;
  assign n64189 = n32222 | n32223;
  assign n64190 = n32225 | n32226;
  assign n64191 = n32232 | n32233;
  assign n64192 = n32235 | n32236;
  assign n64193 = n32249 | ~n32250;
  assign n64194 = n32275 | n32276;
  assign n64195 = n32330 | n32327 | n32329;
  assign n64196 = n32376 | n32373 | n32375;
  assign n64197 = n32377 | n32378;
  assign n64198 = n32404 | n32405;
  assign n64199 = n32414 | n32415;
  assign n64200 = n32428 | n32429;
  assign n64201 = n32436 | n32437;
  assign n64202 = n32442 | n32439 | n32441;
  assign n64203 = n32452 | n32453;
  assign n64204 = n32462 | n32463;
  assign n64205 = n32468 | n32469;
  assign n64206 = n32474 | n32471 | n32473;
  assign n64207 = n32494 | n32495;
  assign n64208 = n32505 | n32506;
  assign n64209 = n32521 | n32522;
  assign n64210 = n32528 | n32529;
  assign n64211 = n32532 | n32533;
  assign n64212 = n32538 | n32539;
  assign n64213 = n32542 | n32543;
  assign n64214 = n32561 | n32562;
  assign n64215 = n32574 | n32575;
  assign n64216 = n32597 | ~n32598;
  assign n64217 = n32627 | ~n32628;
  assign n64218 = n32649 | n32650;
  assign n64219 = n32756 | n32757;
  assign n64220 = n32771 | n32772;
  assign n64221 = n32799 | n32800;
  assign n64222 = n32817 | n32818;
  assign n64223 = n32856 | n32857;
  assign n64224 = n32879 | n32880;
  assign n64225 = n32938 | n32939;
  assign n64226 = n32950 | n32951;
  assign n64227 = n32952 | n32953;
  assign n64228 = n32969 | n32970;
  assign n64229 = n33020 | n33021;
  assign n64230 = n33041 | n33042;
  assign n64231 = n33051 | n33052;
  assign n64232 = n33076 | n33077;
  assign n64233 = n33078 | n33079;
  assign n64234 = n33085 | n33086;
  assign n64235 = n33092 | n33093;
  assign n64236 = n33112 | n33113;
  assign n64237 = n33115 | n33116;
  assign n64238 = n33126 | n33127;
  assign n64239 = n33182 | n33183;
  assign n64240 = n33184 | n33185;
  assign n64241 = n33201 | n33202;
  assign n64242 = n33206 | n33207;
  assign n64243 = n33211 | n33208 | n33210;
  assign n64244 = n33212 | n33213;
  assign n64245 = n33216 | n33214 | n33215;
  assign n64246 = n33222 | n33223;
  assign n64247 = n33231 | n33232;
  assign n64248 = n33264 | n33265;
  assign n64249 = n33272 | n33273;
  assign n64250 = n33328 | ~n33329;
  assign n64251 = n33331 | n33332;
  assign n64252 = n33336 | n33337;
  assign n64253 = n33342 | n33343;
  assign n64254 = n33350 | n33351;
  assign n64255 = n33380 | n33381;
  assign n64256 = n33396 | n33392 | n33395;
  assign n64257 = n33409 | n33410;
  assign n64258 = n33417 | n33418;
  assign n64259 = n33425 | n33426;
  assign n64260 = n33466 | n33467;
  assign n64261 = n33470 | n33471;
  assign n64262 = n33481 | n33478 | n33480;
  assign n64263 = n33488 | n33485 | n33487;
  assign n64264 = n33495 | n33496;
  assign n64265 = n33502 | n33503;
  assign n64266 = n33508 | n33509;
  assign n64267 = n33517 | n33518;
  assign n64268 = n33523 | n33524;
  assign n64269 = n33533 | n33534;
  assign n64270 = n33550 | n33551;
  assign n64271 = n33562 | n33563;
  assign n64272 = n33570 | n33571;
  assign n64273 = n33572 | ~n33573;
  assign n64274 = n33595 | n33596;
  assign n64275 = n33614 | n33615;
  assign n64276 = n33631 | n33632;
  assign n64277 = n33642 | n33643;
  assign n64278 = n33651 | n33652;
  assign n64279 = n33654 | n33655;
  assign n64280 = n33701 | n33694 | n33700;
  assign n64281 = n33698 | n33699;
  assign n64282 = n33726 | n33727;
  assign n64283 = n33746 | n33747;
  assign n64284 = n33755 | n33756;
  assign n64285 = n33763 | n33764;
  assign n64286 = n33776 | n33777;
  assign n64287 = n33784 | n33785;
  assign n64288 = n33819 | n33820;
  assign n64289 = n33824 | n33825;
  assign n64290 = n33826 | n33827;
  assign n64291 = n33830 | n33831;
  assign n64292 = n33853 | n33854;
  assign n64293 = n33863 | n33864;
  assign n64294 = n33865 | n33866;
  assign n64295 = n33947 | n33948;
  assign n64296 = n33952 | n33950 | n33951;
  assign n64297 = n33970 | n33967 | n33969;
  assign n64298 = n33978 | n33979;
  assign n64299 = n34002 | n33999 | n34001;
  assign n64300 = n34020 | n34021;
  assign n64301 = n34026 | n34027;
  assign n64302 = n34029 | n34030;
  assign n64303 = n34041 | n34042;
  assign n64304 = n34064 | n34061 | n34063;
  assign n64305 = n34070 | n34065 | n34069;
  assign n64306 = n34067 | n34068;
  assign n64307 = n34073 | ~n34074;
  assign n64308 = n34105 | n34106;
  assign n64309 = n34147 | ~n34148;
  assign n64310 = n34234 | n34235;
  assign n64311 = n34250 | n34251;
  assign n64312 = n34268 | ~n34269;
  assign n64313 = n34405 | n34406;
  assign n64314 = n34414 | n34415;
  assign n64315 = n34944 | n34945;
  assign n64316 = n34946 | n34947;
  assign n64317 = n35007 | n35008;
  assign po281 = n35020 | ~n35021;
  assign n64319 = n35022 | n35023;
  assign n64320 = n35031 | n35032;
  assign n64321 = n35042 | n35043;
  assign n64322 = n35048 | n35049;
  assign n64323 = n35071 | ~n35072;
  assign n64324 = n35110 | n35111;
  assign n64325 = n35114 | n35115;
  assign n64326 = n35136 | n35137;
  assign n64327 = n35142 | n35143;
  assign n64328 = n35156 | n35157;
  assign n64329 = n35159 | n35160;
  assign n64330 = n35224 | n35225;
  assign n64331 = n35230 | n35231;
  assign n64332 = n35244 | n35245;
  assign n64333 = n35247 | n35248;
  assign n64334 = n35298 | n35299;
  assign n64335 = n35313 | n35314;
  assign n64336 = n35361 | n35362;
  assign n64337 = n35363 | n35364;
  assign n64338 = n35399 | n35395 | n35398;
  assign n64339 = n35396 | n35397;
  assign n64340 = n35401 | n35402;
  assign n64341 = n35423 | n35421 | n35422;
  assign n64342 = n35451 | n35452;
  assign n64343 = n35458 | ~n35459;
  assign n64344 = n35474 | n35475;
  assign n64345 = n35483 | ~n35484;
  assign n64346 = n35485 | n35486;
  assign n64347 = n35497 | n35498;
  assign n64348 = n35512 | n35513;
  assign n64349 = n35523 | n35524;
  assign n64350 = n35526 | n35527;
  assign n64351 = n35541 | n35542;
  assign n64352 = n35547 | n35548;
  assign n64353 = n35553 | n35550 | n35552;
  assign n64354 = n35557 | n35558;
  assign n64355 = n35561 | n35562;
  assign n64356 = n35598 | n35599;
  assign n64357 = n35608 | n35609;
  assign n64358 = n35613 | n35614;
  assign n64359 = n35620 | n35621;
  assign n64360 = n35624 | n35625;
  assign n64361 = n35626 | ~n35627;
  assign n64362 = n35645 | n35646;
  assign n64363 = n35682 | n35683;
  assign n64364 = n35685 | n35686;
  assign n64365 = n35702 | n35703;
  assign n64366 = n35711 | n35712;
  assign n64367 = n35735 | n35736;
  assign n64368 = n35768 | n35765 | n35767;
  assign n64369 = n35800 | n35801;
  assign n64370 = n35833 | n35834;
  assign n64371 = n35840 | n35841;
  assign n64372 = n35880 | n35881;
  assign n64373 = n35884 | n35885;
  assign n64374 = n35889 | n35890;
  assign n64375 = n35907 | n35908;
  assign n64376 = n35930 | n35931;
  assign n64377 = n35943 | n35941 | n35942;
  assign n64378 = n35952 | n35949 | n35951;
  assign n64379 = n35990 | n35991;
  assign n64380 = n35999 | n36000;
  assign n64381 = n36045 | n36046;
  assign n64382 = n36052 | n36053;
  assign n64383 = n36061 | n36058 | n36060;
  assign n64384 = n36087 | n36088;
  assign n64385 = n36102 | n36103;
  assign n64386 = n36128 | n36129;
  assign n64387 = n36135 | n36136;
  assign n64388 = n36140 | n36141;
  assign n64389 = n36183 | n36184;
  assign n64390 = n36215 | n36216;
  assign n64391 = n36225 | n36226;
  assign n64392 = n36238 | n36239;
  assign n64393 = n36242 | n36243;
  assign n64394 = n36245 | n36246;
  assign n64395 = n36250 | n36251;
  assign n64396 = n36272 | n36273;
  assign n64397 = n36283 | n36284;
  assign n64398 = n36320 | n36321;
  assign n64399 = n36350 | n36351;
  assign n64400 = n36361 | n36362;
  assign n64401 = n36366 | n36367 | n36368 | n36369;
  assign n64402 = n36378 | n36379;
  assign n64403 = n36404 | n36405;
  assign n64404 = n36416 | n36417;
  assign n64405 = n36430 | n36431;
  assign n64406 = n36436 | n36437;
  assign n64407 = n36448 | n36449;
  assign n64408 = n36455 | n36456;
  assign n64409 = n36493 | n36494;
  assign n64410 = n36497 | n36498;
  assign n64411 = n36502 | n36503;
  assign n64412 = n36520 | n36521;
  assign n64413 = n36543 | n36544;
  assign n64414 = n36556 | n36554 | n36555;
  assign n64415 = n36565 | n36562 | n36564;
  assign n64416 = n36596 | n36597;
  assign n64417 = n36619 | n36620;
  assign n64418 = n36632 | n36630 | n36631;
  assign n64419 = n36641 | n36638 | n36640;
  assign n64420 = n36691 | n36692;
  assign n64421 = n36697 | n36698;
  assign n64422 = n36736 | n36737;
  assign n64423 = n36740 | n36741;
  assign n64424 = n36745 | n36746;
  assign n64425 = n36764 | n36765;
  assign n64426 = n36779 | n36780;
  assign n64427 = n36801 | n36802;
  assign n64428 = n36808 | n36809;
  assign n64429 = n36813 | n36814;
  assign n64430 = n36859 | n36860;
  assign n64431 = n36884 | n36881 | n36883;
  assign n64432 = n36889 | n36890;
  assign n64433 = n36914 | n36915;
  assign n64434 = n36932 | n36930 | n36931;
  assign n64435 = n36935 | n36936;
  assign n64436 = n36940 | n36941;
  assign n64437 = n36964 | n36965;
  assign n64438 = n36971 | n36972;
  assign n64439 = n37010 | n37011;
  assign n64440 = n37014 | n37015;
  assign n64441 = n37019 | n37020;
  assign n64442 = n37067 | n37068;
  assign n64443 = n37112 | n37113;
  assign n64444 = n37146 | n37147;
  assign n64445 = n37152 | n37153;
  assign n64446 = n37164 | n37165;
  assign n64447 = n37168 | n37169;
  assign n64448 = n37176 | n37177;
  assign n64449 = n37182 | n37183;
  assign n64450 = n37184 | n37185;
  assign n64451 = n37189 | n37190;
  assign n64452 = n37254 | n37255;
  assign n64453 = n37264 | n37265;
  assign n64454 = n37280 | n37281;
  assign n64455 = n37289 | n37290;
  assign n64456 = n37321 | n37322;
  assign n64457 = n37331 | n37332;
  assign n64458 = n37344 | n37345;
  assign n64459 = n37348 | n37349;
  assign n64460 = n37351 | n37352;
  assign n64461 = n37356 | n37357;
  assign n64462 = n37378 | n37379;
  assign n64463 = n37389 | n37390;
  assign n64464 = n37398 | n37399;
  assign n64465 = n37430 | n37431;
  assign n64466 = n37440 | n37441;
  assign n64467 = n37453 | n37454;
  assign n64468 = n37457 | n37458;
  assign n64469 = n37460 | n37461;
  assign n64470 = n37465 | n37466;
  assign n64471 = n37487 | n37488;
  assign n64472 = n37498 | n37499;
  assign n64473 = n37512 | n37513;
  assign n64474 = n37560 | n37561;
  assign n64475 = n37588 | n37589;
  assign n64476 = n37620 | n37621;
  assign n64477 = n37630 | n37631;
  assign n64478 = n37643 | n37644;
  assign n64479 = n37647 | n37648;
  assign n64480 = n37650 | n37651;
  assign n64481 = n37655 | n37656;
  assign n64482 = n37677 | n37678;
  assign n64483 = n37688 | n37689;
  assign n64484 = n37697 | n37698;
  assign n64485 = n37704 | n37705;
  assign n64486 = n37713 | n37714;
  assign n64487 = n37727 | n37728;
  assign n64488 = n37760 | n37761;
  assign n64489 = n37767 | n37768;
  assign n64490 = n37772 | n37773;
  assign n64491 = n37782 | n37783;
  assign n64492 = n37793 | n37794;
  assign n64493 = n37818 | n37819;
  assign n64494 = n37856 | n37857;
  assign n64495 = n37860 | n37861;
  assign n64496 = n37865 | n37866;
  assign n64497 = n37882 | n37883;
  assign n64498 = n37886 | n37884 | n37885;
  assign n64499 = n37888 | n37889;
  assign n64500 = n37897 | n37898;
  assign n64501 = n37901 | n37902;
  assign n64502 = n37914 | n37915;
  assign n64503 = n37927 | n37928;
  assign n64504 = n37940 | n37941;
  assign n64505 = n37953 | n37954;
  assign n64506 = n37963 | n37964;
  assign n64507 = n37974 | n37975;
  assign n64508 = n37981 | n37982;
  assign n64509 = n37989 | n37990;
  assign n64510 = n38002 | n38003;
  assign n64511 = n38015 | n38016;
  assign n64512 = n38025 | n38026;
  assign n64513 = n38041 | n38042;
  assign n64514 = n38126 | n38127;
  assign n64515 = n38157 | n38158;
  assign n64516 = n38162 | n38163;
  assign n64517 = n38172 | n38173;
  assign n64518 = n38183 | n38184;
  assign n64519 = n38185 | n38186;
  assign n64520 = n38190 | n38191;
  assign n64521 = n38194 | n58851;
  assign n64522 = n58862 | n38195 | n38196;
  assign n64523 = n38201 | n38198 | n38200;
  assign n64524 = n38215 | n38216;
  assign n64525 = n38223 | n38224;
  assign n64526 = n38240 | n38241;
  assign n64527 = n38248 | n38249;
  assign n64528 = n38257 | n38258;
  assign n64529 = n38274 | n38275;
  assign n64530 = n38276 | n38277;
  assign n64531 = n38286 | n38287;
  assign n64532 = n38296 | n38293 | n38295;
  assign n64533 = n38307 | n38308;
  assign n64534 = n38311 | n38312;
  assign n64535 = n38314 | n38315;
  assign n64536 = n38357 | n38358;
  assign n64537 = n38396 | n38397;
  assign n64538 = n38402 | n38403;
  assign n64539 = n38408 | n38405 | n38407;
  assign n64540 = n38415 | n38416;
  assign n64541 = n38428 | n38429;
  assign n64542 = n38439 | n38440;
  assign n64543 = n38442 | n38443;
  assign n64544 = n38456 | n38457;
  assign n64545 = n38458 | n38459;
  assign n64546 = n38473 | n38474;
  assign n64547 = n38482 | n38483;
  assign n64548 = n38487 | n38488;
  assign n64549 = n38497 | n38493 | n38496;
  assign n64550 = n38504 | n38505;
  assign n64551 = n38515 | n38516;
  assign n64552 = n38533 | n38534;
  assign n64553 = n38561 | n38562;
  assign n64554 = n38567 | n38568;
  assign n64555 = n38573 | n38570 | n38572;
  assign n64556 = n38594 | n38595;
  assign n64557 = n38605 | n38606;
  assign n64558 = n38611 | n38612;
  assign n64559 = n38618 | n38619;
  assign n64560 = n38660 | n38661;
  assign n64561 = n38666 | n38667;
  assign n64562 = n38670 | n38671;
  assign n64563 = n38687 | n38688;
  assign n64564 = n38702 | n38703;
  assign n64565 = n38708 | n38709;
  assign n64566 = n38714 | n38711 | n38713;
  assign n64567 = n38721 | n38722;
  assign n64568 = n38770 | n38751 | n38769;
  assign n64569 = n38757 | n38758;
  assign n64570 = n38765 | n38766;
  assign n64571 = n38772 | n38773;
  assign n64572 = n38790 | n38791;
  assign n64573 = n38796 | n38797;
  assign n64574 = n38809 | n38810;
  assign n64575 = n38821 | n38822;
  assign n64576 = n38829 | n38830;
  assign n64577 = n38837 | n38838;
  assign n64578 = n38845 | n38846;
  assign n64579 = n38861 | n38862;
  assign n64580 = n38869 | n38870;
  assign n64581 = n38875 | n38876;
  assign n64582 = n38907 | n38908;
  assign n64583 = n38921 | n38922;
  assign po231 = n38937 | n38938;
  assign n64585 = n38945 | n38946;
  assign n64586 = n38954 | n38955;
  assign n64587 = n38964 | n38965;
  assign n64588 = n39017 | n39018;
  assign n64589 = n39023 | n39024;
  assign n64590 = n39048 | n39049;
  assign n64591 = n39054 | n39051 | n39053;
  assign n64592 = n39058 | n39056 | n39057;
  assign n64593 = n39062 | n39063;
  assign n64594 = n39065 | n39066;
  assign n64595 = n39071 | n39067 | n39070;
  assign n64596 = n39074 | n39075;
  assign n64597 = n39081 | n39082;
  assign n64598 = n39101 | n39102;
  assign n64599 = n39104 | n39105;
  assign n64600 = n39123 | n39124;
  assign n64601 = n39129 | n39130;
  assign n64602 = n39131 | n39132;
  assign n64603 = n39152 | n39153;
  assign n64604 = n39154 | n39155;
  assign n64605 = n39178 | n39179;
  assign n64606 = n39194 | n39195;
  assign n64607 = n39206 | n39207;
  assign n64608 = n39221 | n39222;
  assign n64609 = n39224 | n39225;
  assign n64610 = n39229 | n39230;
  assign n64611 = n39246 | n39247;
  assign n64612 = n39249 | n39250;
  assign n64613 = n39251 | n39252;
  assign n64614 = n39266 | n39267;
  assign n64615 = n39268 | n39269;
  assign n64616 = n39271 | n39272;
  assign n64617 = n39275 | ~n39276;
  assign n64618 = n39280 | n39281;
  assign n64619 = n39295 | n39296;
  assign n64620 = n39303 | n39304;
  assign n64621 = n39310 | n39311;
  assign n64622 = n39313 | n39314;
  assign n64623 = n39337 | ~n39338;
  assign n64624 = n39340 | n39341;
  assign n64625 = n39344 | n39345;
  assign n64626 = n39367 | n39368;
  assign n64627 = n39374 | n39375;
  assign n64628 = n39397 | n39398;
  assign n64629 = n39404 | n39405;
  assign n64630 = n39413 | n39414;
  assign n64631 = ~n39429 | n39426 | n39428;
  assign n64632 = n39440 | n39441;
  assign n64633 = n39443 | n39444;
  assign n64634 = n39449 | ~n39450;
  assign n64635 = n39485 | n39486;
  assign n64636 = n39489 | n39490;
  assign n64637 = n39493 | n39494;
  assign n64638 = n39507 | n39508;
  assign n64639 = n39513 | n39514;
  assign n64640 = n39516 | n39517;
  assign n64641 = n39529 | n39530;
  assign n64642 = n39625 | n39626;
  assign n64643 = n39644 | n39645;
  assign n64644 = n39651 | n39652;
  assign n64645 = n39668 | n39669;
  assign n64646 = n39671 | n39672;
  assign n64647 = n39680 | n39681;
  assign n64648 = n39683 | n39684;
  assign n64649 = n39690 | n39691;
  assign n64650 = n39703 | n39704;
  assign n64651 = n39717 | n39718;
  assign n64652 = n39729 | n39730;
  assign n64653 = n39734 | n39735;
  assign n64654 = n39746 | n39747;
  assign n64655 = n39750 | n39751;
  assign n64656 = n39752 | n39753;
  assign n64657 = n39767 | n39768;
  assign n64658 = n39782 | n39780 | n39781;
  assign n64659 = n39804 | n39805;
  assign n64660 = n39816 | n39817;
  assign n64661 = n39831 | n39832;
  assign n64662 = n39858 | n39854 | n39857;
  assign n64663 = n39871 | n39872;
  assign n64664 = n39891 | n39892;
  assign n64665 = n39900 | n39901;
  assign n64666 = n39910 | n39911;
  assign n64667 = n39928 | n39929;
  assign n64668 = n39934 | n39935;
  assign n64669 = n39957 | n39958;
  assign n64670 = n39964 | ~n39965;
  assign n64671 = n39973 | n39974;
  assign n64672 = n39988 | n39989;
  assign n64673 = n39990 | n39991;
  assign n64674 = n40005 | n40006;
  assign n64675 = n40009 | n40010;
  assign n64676 = n40016 | n40017;
  assign n64677 = n40034 | n40035;
  assign n64678 = n40075 | n40076;
  assign n64679 = n40081 | n40082;
  assign n64680 = n40085 | n40086;
  assign n64681 = n40110 | n40111;
  assign n64682 = n40114 | n40115;
  assign n64683 = n40130 | n40131;
  assign n64684 = n40133 | n40134;
  assign n64685 = n40147 | n40138 | n40146;
  assign n64686 = n40169 | n40170;
  assign po223 = n40173 | n40174;
  assign n64688 = n40182 | n40183;
  assign n64689 = n40268 | n40269;
  assign n64690 = n40285 | n40286;
  assign n64691 = n40308 | n40309;
  assign n64692 = n40356 | n40357;
  assign n64693 = n40374 | n40375;
  assign n64694 = n40382 | n40383;
  assign n64695 = n40403 | n40404;
  assign n64696 = n40479 | n40480;
  assign n64697 = n40514 | n40515;
  assign n64698 = n40519 | n40520;
  assign n64699 = n40556 | n40553 | n40555;
  assign n64700 = n40592 | n40593;
  assign n64701 = n40607 | n40605 | n40606;
  assign n64702 = n40661 | n40662;
  assign n64703 = n40676 | n40677;
  assign n64704 = n40686 | n40687;
  assign n64705 = n40696 | n40690 | n40692 | n40700 | n40698 | n40699;
  assign n64706 = n40695 | n40693 | n40694;
  assign n64707 = n40704 | n40705;
  assign n64708 = n40723 | n40724;
  assign n64709 = n40753 | n40754;
  assign n64710 = n40767 | n40768;
  assign n64711 = n40777 | n40778;
  assign po234 = n40787 | n40788;
  assign n64713 = n40839 | n40840;
  assign n64714 = n40843 | n40844;
  assign n64715 = n40852 | n40853;
  assign n64716 = n40864 | n40865;
  assign n64717 = n40873 | n40874;
  assign n64718 = n40889 | n40890;
  assign n64719 = n40899 | n40900;
  assign n64720 = n40912 | n40913;
  assign n64721 = n40926 | n40927;
  assign n64722 = n40956 | n40957;
  assign n64723 = n40984 | n40985;
  assign n64724 = n40986 | n40987;
  assign n64725 = n41025 | n41026;
  assign n64726 = n41051 | n41052;
  assign n64727 = n41106 | n41107;
  assign n64728 = n41111 | n41112;
  assign n64729 = n41117 | n41118;
  assign n64730 = n41127 | n41128;
  assign n64731 = n41129 | n41130;
  assign n64732 = n41165 | n41166;
  assign n64733 = n41169 | ~n41170;
  assign n64734 = n41212 | n41213;
  assign n64735 = n41217 | n41218;
  assign n64736 = n41222 | n41223;
  assign n64737 = n41243 | n41244;
  assign n64738 = n41260 | n41261;
  assign n64739 = n41285 | ~n41286;
  assign n64740 = n41305 | n41306;
  assign n64741 = n41421 | n41422;
  assign n64742 = n41427 | n41428;
  assign n64743 = n41448 | n41449;
  assign n64744 = n41458 | n41459;
  assign n64745 = n41461 | n41462;
  assign n64746 = n41499 | n41500;
  assign n64747 = n41505 | n41506;
  assign n64748 = n41510 | n41511;
  assign n64749 = n41537 | n41538;
  assign n64750 = n41543 | n41544;
  assign n64751 = n41572 | n41573;
  assign n64752 = n41579 | n41580;
  assign n64753 = n41607 | n41598 | n41606;
  assign n64754 = n41723 | ~n41724;
  assign n64755 = n41737 | n41738;
  assign n64756 = n41752 | n41753;
  assign n64757 = n41771 | n41772;
  assign n64758 = n41792 | n41793;
  assign n64759 = n41803 | n41804;
  assign n64760 = n41819 | n41820;
  assign n64761 = n41824 | n41825;
  assign n64762 = n41827 | n41828;
  assign n64763 = n41833 | n41834;
  assign n64764 = n41840 | n41841;
  assign n64765 = n41863 | n41864;
  assign n64766 = n41881 | n41882;
  assign n64767 = n41892 | n41893;
  assign n64768 = n41935 | n41936;
  assign n64769 = n41941 | n41939 | n41940;
  assign n64770 = n41965 | n41966;
  assign n64771 = n41970 | n41971;
  assign n64772 = n41983 | n41984;
  assign n64773 = n42006 | n42007;
  assign n64774 = n42034 | n42035;
  assign n64775 = n42044 | n42045;
  assign n64776 = n42098 | n42099;
  assign n64777 = n42113 | n42114;
  assign n64778 = n42120 | n42121;
  assign n64779 = n42163 | n42164;
  assign n64780 = n42195 | n42196;
  assign n64781 = n42208 | n42209;
  assign n64782 = n42216 | n42220 | n42222 | n42223;
  assign n64783 = n42227 | n42228;
  assign n64784 = n42248 | n42249;
  assign n64785 = n42307 | n42308;
  assign n64786 = n42333 | n42334;
  assign n64787 = n42343 | n42344;
  assign n64788 = n42370 | n42371;
  assign n64789 = n42399 | n42400;
  assign n64790 = n42408 | n42409;
  assign n64791 = n42412 | n42413;
  assign n64792 = n42422 | ~n42423;
  assign n64793 = n42431 | ~n42432;
  assign n64794 = n42467 | n42468;
  assign n64795 = n42472 | n42473;
  assign n64796 = n42488 | n42483 | n42487;
  assign n64797 = n42515 | n42512 | n42514;
  assign n64798 = n42518 | n42519;
  assign n64799 = n42525 | n42526;
  assign n64800 = n42575 | n42576;
  assign n64801 = n42588 | n42589;
  assign n64802 = n42623 | n42624;
  assign n64803 = n42676 | n42677;
  assign n64804 = n42690 | n42691;
  assign n64805 = n42714 | ~n42715;
  assign n64806 = n42724 | n42725;
  assign n64807 = n42733 | n42734;
  assign n64808 = n42741 | n42742;
  assign n64809 = n42759 | n42760;
  assign n64810 = n42769 | n42770;
  assign n64811 = n42786 | n42787;
  assign n64812 = n42788 | n42789;
  assign n64813 = n42806 | n42807;
  assign n64814 = n42843 | n42844;
  assign n64815 = n42851 | n42852;
  assign n64816 = n42892 | n42893;
  assign n64817 = n42904 | n42905;
  assign n64818 = n42919 | n42920;
  assign n64819 = n42941 | n42938 | n42940;
  assign n64820 = n42953 | n42948 | n42952;
  assign n64821 = n42957 | n42958;
  assign n64822 = n42971 | n42972;
  assign n64823 = n42993 | n42994;
  assign n64824 = n43005 | n43006;
  assign n64825 = n43057 | n43058;
  assign n64826 = n43062 | n43063;
  assign n64827 = n43068 | n43069;
  assign n64828 = n43075 | n43076;
  assign n64829 = n43086 | n43087;
  assign n64830 = n43104 | n43105;
  assign n64831 = n43108 | n43109;
  assign n64832 = n43140 | n43141;
  assign n64833 = n43154 | n43155;
  assign n64834 = n43166 | ~n43167;
  assign n64835 = n43187 | n43188;
  assign n64836 = n43192 | ~n43193;
  assign n64837 = n43197 | n43198;
  assign n64838 = n43200 | n43201;
  assign n64839 = n43230 | n43220 | n43229;
  assign n64840 = n43255 | n43256;
  assign n64841 = n43267 | n43268;
  assign n64842 = n43295 | n43296;
  assign n64843 = n43299 | n43300;
  assign n64844 = n43311 | n43306 | n43310;
  assign n64845 = n43315 | n43316;
  assign n64846 = n43324 | n43325;
  assign n64847 = n43352 | n43353;
  assign n64848 = n43369 | n43370;
  assign n64849 = n43405 | n43406;
  assign n64850 = n43409 | n43410;
  assign n64851 = n43432 | n43433;
  assign n64852 = n43450 | n43451;
  assign n64853 = n43454 | n43455;
  assign n64854 = n43472 | n43473;
  assign n64855 = n43494 | n43495;
  assign n64856 = n43514 | n43515;
  assign n64857 = n43531 | n43532;
  assign n64858 = n43555 | ~n43556;
  assign po252 = n43560 | n43561;
  assign n64860 = n43578 | n43579;
  assign n64861 = n43612 | n43613;
  assign n64862 = n43618 | n43619;
  assign n64863 = n43620 | n43621;
  assign n64864 = n43636 | n43637;
  assign n64865 = n43674 | n43675;
  assign n64866 = n43680 | n43681;
  assign n64867 = n43711 | n43712;
  assign n64868 = n43716 | n43717;
  assign n64869 = n43722 | n43723;
  assign n64870 = n43752 | n43753;
  assign n64871 = n43769 | n43770;
  assign n64872 = n43806 | n43807;
  assign n64873 = n43814 | ~n43815;
  assign n64874 = n43870 | n43871;
  assign n64875 = n43873 | n43874;
  assign n64876 = n43917 | n43914 | n43916;
  assign n64877 = n43946 | n43947;
  assign n64878 = n43990 | n43991;
  assign n64879 = n44003 | n44004;
  assign n64880 = n44070 | n44058 | n44069;
  assign n64881 = n44073 | n44074;
  assign n64882 = n44082 | n44083;
  assign n64883 = n44130 | n44131;
  assign n64884 = n44169 | n44170;
  assign n64885 = n44194 | n44195;
  assign n64886 = n44203 | n44204;
  assign n64887 = n44242 | n44243;
  assign n64888 = n44288 | n44289;
  assign n64889 = n44307 | n44308;
  assign n64890 = n44335 | n44336;
  assign n64891 = n44357 | n44358;
  assign n64892 = n44415 | n44416;
  assign n64893 = n44471 | n44472;
  assign n64894 = n44560 | n44561;
  assign n64895 = n44580 | n44581;
  assign n64896 = n44599 | n44600;
  assign n64897 = n44625 | n44626;
  assign n64898 = n44637 | n44638;
  assign n64899 = n44668 | n44669;
  assign n64900 = n44713 | n44714;
  assign n64901 = n44730 | n44731;
  assign n64902 = n44738 | n44739;
  assign n64903 = n44809 | n44810;
  assign po158 = n44825 | n44826;
  assign n64905 = n44833 | n44834;
  assign n64906 = n44852 | n44853;
  assign n64907 = n44887 | n44888;
  assign n64908 = n44917 | n44918;
  assign n64909 = n44962 | n44963;
  assign n64910 = n44979 | n44980;
  assign n64911 = n44987 | n44988;
  assign n64912 = n45058 | n45059;
  assign po159 = n45074 | n45075;
  assign n64914 = n45081 | n45082;
  assign n64915 = n45097 | n45098;
  assign n64916 = n45116 | n45117;
  assign n64917 = n45123 | n45124;
  assign n64918 = n45188 | n45189;
  assign n64919 = n45232 | n45233;
  assign n64920 = n45316 | n45317;
  assign n64921 = n45336 | n45337;
  assign n64922 = n45355 | n45356;
  assign n64923 = n45391 | n45392;
  assign n64924 = n45421 | n45422;
  assign n64925 = n45466 | n45467;
  assign n64926 = n45483 | n45484;
  assign n64927 = n45491 | n45492;
  assign n64928 = n45562 | n45563;
  assign po161 = n45578 | n45579;
  assign n64930 = n45586 | n45587;
  assign n64931 = n45605 | n45606;
  assign n64932 = n45641 | n45642;
  assign n64933 = n45671 | n45672;
  assign n64934 = n45716 | n45717;
  assign n64935 = n45733 | n45734;
  assign n64936 = n45741 | n45742;
  assign n64937 = n45812 | n45813;
  assign po162 = n45828 | n45829;
  assign n64939 = n45887 | n45888;
  assign n64940 = n45908 | n45909;
  assign n64941 = n45933 | n45934;
  assign n64942 = n45943 | n45944;
  assign n64943 = n45964 | n45965;
  assign n64944 = n45969 | n45970;
  assign n64945 = n45978 | n45979;
  assign n64946 = n45984 | n45985;
  assign n64947 = n45987 | n45988;
  assign n64948 = n46030 | n46031;
  assign n64949 = n46089 | n46090;
  assign n64950 = n46096 | n46097;
  assign n64951 = n46120 | n46121;
  assign n64952 = n46136 | n46137;
  assign n64953 = n46145 | n46146;
  assign n64954 = n46157 | n46158;
  assign n64955 = n46175 | n46176;
  assign n64956 = n46263 | n46264;
  assign n64957 = n46285 | n46286;
  assign n64958 = n46290 | n46291;
  assign n64959 = n46307 | n46308;
  assign n64960 = n46318 | n46319;
  assign n64961 = n46330 | n46331;
  assign n64962 = n46336 | n46337;
  assign n64963 = n46354 | n46355;
  assign n64964 = n46373 | n46374;
  assign n64965 = n46409 | n46410;
  assign n64966 = n46439 | n46440;
  assign n64967 = n46443 | n46444;
  assign n64968 = n46489 | n46490;
  assign n64969 = n46514 | n46515;
  assign n64970 = n46516 | n46517;
  assign n64971 = n46589 | n46590;
  assign po156 = n46605 | n46606;
  assign n64973 = n46611 | n46612;
  assign n64974 = n46632 | n46633;
  assign n64975 = n46652 | n46653;
  assign n64976 = n46675 | n46676;
  assign n64977 = n46755 | n46756;
  assign n64978 = n46776 | n46777;
  assign n64979 = n46849 | n46850;
  assign n64980 = n46867 | n46868;
  assign n64981 = n46888 | n46889;
  assign n64982 = n46903 | n46904;
  assign n64983 = n47003 | n47004;
  assign n64984 = n47024 | n47025;
  assign n64985 = n47101 | n47102;
  assign n64986 = n47147 | n47148;
  assign n64987 = n47168 | n47169;
  assign n64988 = n47235 | n47236;
  assign n64989 = n47323 | n47324;
  assign n64990 = n47399 | n47400;
  assign n64991 = n47470 | n47471;
  assign n64992 = n47496 | n47497;
  assign po471 = n47502 | n47503;
  assign n64994 = n47505 | n47506;
  assign n64995 = n47516 | n47517;
  assign n64996 = n47537 | n47538;
  assign n64997 = n47544 | n47545;
  assign po637 = n47550 | n47551;
  assign po445 = n47556 | n47557;
  assign n65000 = n47563 | n47564;
  assign n65001 = n47568 | n47569;
  assign n65002 = n47575 | n47576;
  assign n65003 = n47614 | n47615;
  assign n65004 = n47687 | n47688;
  assign n65005 = n47694 | n47695;
  assign n65006 = n47701 | n47698 | n47700;
  assign n65007 = n47703 | n47704;
  assign n65008 = n47721 | n47722;
  assign n65009 = n47724 | n47725;
  assign n65010 = n47728 | n47729;
  assign n65011 = n47743 | n47744;
  assign n65012 = n47771 | ~n47772;
  assign n65013 = n47786 | n47787;
  assign n65014 = n47804 | n47805;
  assign n65015 = n47815 | n47812 | n47814;
  assign n65016 = n47886 | n47883 | n47885;
  assign n65017 = n47922 | n47923;
  assign n65018 = n47933 | n47934;
  assign n65019 = n47987 | n47985 | n47986;
  assign n65020 = n47994 | n47991 | n47993;
  assign n65021 = n48004 | n48005;
  assign n65022 = n48011 | n48012;
  assign n65023 = n48018 | n48019;
  assign n65024 = n48023 | n48024;
  assign n65025 = n48059 | n48060;
  assign n65026 = n48079 | n48076 | n48078;
  assign n65027 = n48089 | n48090;
  assign n65028 = n48096 | ~n48097;
  assign n65029 = n48098 | n48099;
  assign n65030 = n48113 | n48114;
  assign n65031 = n48116 | n48117;
  assign n65032 = n48128 | n48129;
  assign n65033 = n48131 | n48132;
  assign n65034 = n48135 | n48136;
  assign n65035 = n48150 | n48151;
  assign n65036 = n48160 | n48161;
  assign n65037 = n48168 | n48169;
  assign n65038 = n48179 | n48180;
  assign n65039 = n48232 | n48233;
  assign n65040 = n48239 | n48240;
  assign n65041 = n48250 | n48251;
  assign n65042 = n48442 | n48443;
  assign n65043 = n48462 | n48463;
  assign n65044 = n48500 | ~n48501;
  assign po211 = n48520 | n48521;
  assign n65046 = n48555 | n48556;
  assign n65047 = n48604 | n48605;
  assign n65048 = n48608 | n48609;
  assign n65049 = n48614 | n48615;
  assign n65050 = n48616 | n48617;
  assign n65051 = n48625 | n48626;
  assign n65052 = n48645 | n48651 | n48652 | n48653;
  assign n65053 = n48648 | n48649;
  assign po212 = n48671 | n48672;
  assign n65055 = n48681 | n48682;
  assign po220 = n48691 | n48692;
  assign po247 = n48704 | n48705;
  assign n65058 = n48709 | n48710;
  assign n65059 = n48711 | n48712;
  assign n65060 = n48715 | n48716;
  assign po251 = n48725 | n48726;
  assign n65062 = n48756 | n48757;
  assign n65063 = n48762 | n48763;
  assign po206 = n48777 | n48778;
  assign n65065 = n48781 | n48779 | n48780;
  assign n65066 = n48787 | n48788;
  assign po222 = n48812 | n48813;
  assign n65068 = n48817 | n48818;
  assign po225 = n48821 | n48822;
  assign n65070 = n48840 | n48841;
  assign n65071 = n48856 | n48857;
  assign n65072 = n48864 | n48865;
  assign po209 = n48899 | n48900;
  assign n65074 = n48910 | n48911;
  assign n65075 = n48916 | n48917;
  assign n65076 = n48924 | n48925;
  assign n65077 = n48930 | n48931;
  assign n65078 = n48936 | n48937;
  assign n65079 = n48973 | ~n48974;
  assign po1076 = n48979 | ~n48980;
  assign n65081 = n48988 | ~n48989;
  assign n65082 = n48997 | ~n48998;
  assign n65083 = n49003 | ~n49004;
  assign n65084 = n49021 | ~n49022;
  assign po1100 = n49030 | ~n49031;
  assign n65086 = n49048 | n49045 | n49047;
  assign n65087 = n49060 | n49061;
  assign n65088 = n49062 | ~n49063;
  assign n65089 = n49067 | ~n49068;
  assign n65090 = n49070 | n49072 | ~n49075 | ~n49076;
  assign n65091 = n49086 | n49083 | n49085;
  assign n65092 = n49121 | n49122;
  assign n65093 = n49139 | n49140;
  assign n65094 = n49147 | n49148;
  assign n65095 = n49154 | n49155;
  assign n65096 = n49158 | n49159;
  assign n65097 = n49160 | n49161;
  assign n65098 = n49176 | n49177;
  assign n65099 = n49199 | n49200;
  assign n65100 = n49227 | n49228;
  assign n65101 = n49232 | ~n49233;
  assign n65102 = n49297 | n49298;
  assign n65103 = n49299 | n49300;
  assign n65104 = n49315 | n49316;
  assign n65105 = n49346 | n49347;
  assign n65106 = n49367 | n49368;
  assign n65107 = n49412 | n49413;
  assign n65108 = n49446 | n53742;
  assign n65109 = n49486 | n49487;
  assign n65110 = n49489 | n49490;
  assign n65111 = n49495 | n49496;
  assign n65112 = n49529 | n49530;
  assign n65113 = n49538 | n49539;
  assign n65114 = n49563 | n49564;
  assign n65115 = n49566 | n49567;
  assign n65116 = n49590 | n49591;
  assign n65117 = n49601 | n49602;
  assign n65118 = n49630 | n49618 | n49629;
  assign n65119 = n49620 | n49621;
  assign n65120 = n49627 | n53985;
  assign n65121 = n49647 | n49648;
  assign n65122 = n49687 | n49688;
  assign n65123 = n49696 | n49697;
  assign n65124 = n49700 | n49701;
  assign n65125 = n49717 | n49718;
  assign n65126 = n49763 | n49764;
  assign n65127 = n49778 | n49779;
  assign n65128 = n49785 | n49786;
  assign n65129 = n49792 | n49793;
  assign n65130 = n49814 | n49815;
  assign n65131 = n49824 | n49825;
  assign n65132 = n49834 | n49835;
  assign n65133 = n49844 | n49845;
  assign n65134 = n49918 | n49919;
  assign n65135 = n49948 | n49949;
  assign n65136 = n49952 | n49953;
  assign n65137 = n49956 | n49957;
  assign n65138 = n49966 | n49967;
  assign n65139 = n49977 | n49978;
  assign n65140 = n49992 | n49993;
  assign n65141 = n49997 | n49998;
  assign n65142 = n50003 | n50004;
  assign n65143 = n50011 | n50008 | n50010;
  assign n65144 = n50021 | n50022;
  assign n65145 = n50073 | n50074;
  assign n65146 = n52659 | n50113 | n50114;
  assign n65147 = n50120 | n50121;
  assign n65148 = n50124 | n50125;
  assign n65149 = n50131 | n50132;
  assign n65150 = n50144 | n50145;
  assign n65151 = n50154 | n50155;
  assign n65152 = n50158 | n50159;
  assign n65153 = n50163 | ~n50164;
  assign n65154 = n50202 | n50203;
  assign n65155 = n50225 | n50226;
  assign n65156 = n50239 | n50240;
  assign n65157 = n50270 | n50271;
  assign n65158 = n50328 | n50329;
  assign n65159 = n50341 | n50342;
  assign n65160 = n50371 | n50372;
  assign n65161 = n50381 | n50382;
  assign n65162 = n50394 | n50395;
  assign n65163 = n50407 | n50408;
  assign n65164 = n50423 | n50420 | n50422;
  assign n65165 = n50464 | n50465;
  assign n65166 = n50480 | n50481;
  assign n65167 = n50503 | n50504;
  assign n65168 = n50511 | n50512;
  assign n65169 = n50518 | n50519;
  assign n65170 = n50520 | n50521;
  assign n65171 = n50559 | n50560;
  assign n65172 = n50561 | ~n50562;
  assign n65173 = n50569 | n50570;
  assign n65174 = n50578 | n50579;
  assign n65175 = n50586 | n50587;
  assign n65176 = n50590 | n50591;
  assign n65177 = n50593 | n50594;
  assign n65178 = n50601 | n50602;
  assign n65179 = n50631 | n50628 | n50630;
  assign n65180 = n50634 | n50635;
  assign n65181 = n50726 | n50727;
  assign n65182 = n50735 | n50736;
  assign n65183 = n50755 | n50756;
  assign n65184 = n50769 | n50770;
  assign n65185 = n50775 | n50776;
  assign n65186 = n50813 | n50814;
  assign n65187 = n50822 | n50823;
  assign n65188 = n50828 | n50829;
  assign n65189 = n50855 | n50856;
  assign n65190 = n50864 | n50865;
  assign n65191 = n50870 | n50871;
  assign n65192 = n50897 | n50898;
  assign n65193 = n50906 | n50907;
  assign n65194 = n50927 | n50928;
  assign n65195 = n50933 | n50934;
  assign n65196 = n50942 | n50943;
  assign n65197 = n50956 | n50957;
  assign n65198 = n50972 | n50969 | n50971;
  assign n65199 = n50976 | n50977;
  assign n65200 = n50984 | n50985;
  assign n65201 = n51004 | n51005;
  assign n65202 = n51010 | n51011;
  assign n65203 = n51037 | n51038;
  assign n65204 = n51046 | n51047;
  assign n65205 = n51066 | n51067;
  assign n65206 = n51072 | n51073;
  assign n65207 = n51098 | n51099;
  assign n65208 = n51106 | n51107;
  assign n65209 = n51118 | n51119;
  assign n65210 = n51128 | n51129;
  assign n65211 = n51147 | n51148;
  assign n65212 = n51155 | ~n51156;
  assign n65213 = n51168 | n51169;
  assign n65214 = n51191 | n51192;
  assign n65215 = n51199 | ~n51200;
  assign n65216 = n51211 | n51212;
  assign n65217 = n51220 | n51221;
  assign n65218 = n51227 | n51228;
  assign n65219 = n51248 | n51249;
  assign n65220 = n51255 | n51256;
  assign n65221 = n51269 | n51270;
  assign n65222 = n51279 | ~n51280;
  assign n65223 = n51298 | n51299;
  assign n65224 = n51316 | n51317;
  assign n65225 = n51318 | n51319;
  assign n65226 = n51325 | n51326;
  assign n65227 = n51347 | n51348;
  assign n65228 = n51354 | n51355;
  assign n65229 = n51367 | n51368;
  assign n65230 = n51377 | ~n51378;
  assign n65231 = n51383 | n51384;
  assign n65232 = n51392 | n51393;
  assign n65233 = n51394 | n51395;
  assign n65234 = n51409 | n51410;
  assign n65235 = n51419 | n51420;
  assign n65236 = n51440 | n51441;
  assign n65237 = n51447 | n51448;
  assign n65238 = n51460 | n51461;
  assign n65239 = n51470 | ~n51471;
  assign n65240 = n51482 | n51483;
  assign n65241 = n51490 | n51491;
  assign n65242 = n51502 | n51503;
  assign n65243 = n51510 | n51511;
  assign n65244 = n51534 | n51535;
  assign n65245 = n51550 | n51551;
  assign n65246 = n51552 | n51553;
  assign n65247 = n51559 | n51560;
  assign n65248 = n51565 | n51566;
  assign n65249 = n51578 | ~n51579;
  assign n65250 = n51594 | n51595;
  assign n65251 = n51604 | n51605;
  assign n65252 = n51606 | n51607;
  assign n65253 = n51627 | n51628;
  assign n65254 = n51643 | n51644;
  assign n65255 = n51645 | n51646;
  assign n65256 = n51652 | n51653;
  assign n65257 = n51670 | ~n51671;
  assign n65258 = n51686 | n51687;
  assign n65259 = n51696 | n51697;
  assign n65260 = n51698 | n51699;
  assign n65261 = n51714 | n51715;
  assign n65262 = n51722 | n51723;
  assign n65263 = n51734 | n51735;
  assign n65264 = n51742 | n51743;
  assign n65265 = n51763 | ~n51764;
  assign n65266 = n51778 | n51779;
  assign n65267 = n51784 | n51785;
  assign n65268 = n51793 | n51794;
  assign n65269 = n51802 | n51803;
  assign n65270 = n51822 | n51823;
  assign n65271 = n51828 | n51829;
  assign n65272 = n51856 | n51857;
  assign n65273 = n51864 | n51865;
  assign n65274 = n51870 | n51871;
  assign n65275 = n51878 | n51879;
  assign n65276 = n51890 | n51891;
  assign n65277 = n51896 | n51897;
  assign n65278 = n51923 | n51924;
  assign n65279 = n51943 | n51944;
  assign n65280 = n51951 | n51952;
  assign n65281 = n51957 | n51958;
  assign n65282 = n51965 | n51966;
  assign n65283 = n51977 | n51978;
  assign n65284 = n51997 | n51998;
  assign n65285 = n52013 | n52014;
  assign n65286 = n52033 | n52034;
  assign n65287 = n52049 | n52050;
  assign n65288 = n52069 | n52070;
  assign n65289 = n52085 | n52086;
  assign n65290 = n52105 | n52106;
  assign n65291 = n52121 | n52122;
  assign n65292 = n52141 | n52142;
  assign n65293 = n52163 | ~n52164;
  assign n65294 = n52169 | ~n52170;
  assign n65295 = n52175 | ~n52176;
  assign n65296 = n52181 | ~n52182;
  assign n65297 = n52187 | ~n52188;
  assign n65298 = n52199 | ~n52200;
  assign n65299 = n52205 | ~n52206;
  assign n65300 = n52211 | ~n52212;
  assign n65301 = n52217 | ~n52218;
  assign n65302 = n52223 | ~n52224;
  assign n65303 = n52229 | ~n52230;
  assign n65304 = n52235 | ~n52236;
  assign n65305 = n52241 | ~n52242;
  assign n65306 = n52258 | n52259;
  assign n65307 = n52274 | n52275;
  assign n65308 = n52276 | n52277;
  assign n65309 = n52283 | n52284;
  assign n65310 = n52367 | n52368;
  assign n65311 = n52412 | n52413;
  assign n65312 = n52418 | n52419;
  assign n65313 = n52420 | ~n52421;
  assign n65314 = n52423 | n52424;
  assign n65315 = n52434 | n52435;
  assign n65316 = n52452 | n52453;
  assign n65317 = n52458 | n53347;
  assign n65318 = n52460 | ~n52461;
  assign n65319 = n52471 | n52472;
  assign n65320 = n52491 | n52485 | n52490;
  assign n65321 = n52500 | n52501;
  assign n65322 = n52505 | n52506;
  assign n65323 = n52514 | ~n52515;
  assign n65324 = n52529 | ~n52530;
  assign n65325 = n52532 | n52533;
  assign n65326 = n52560 | n52561;
  assign n65327 = n52564 | n52565;
  assign n65328 = n52585 | n52586;
  assign n65329 = n52589 | n52590;
  assign n65330 = n52598 | n52599;
  assign n65331 = n52601 | n52602;
  assign n65332 = n52616 | n52611 | n52615;
  assign n65333 = n52619 | n52620;
  assign n65334 = n52624 | ~n52625;
  assign n65335 = n52626 | n52627;
  assign n65336 = n52646 | n52647;
  assign n65337 = n52657 | n52658;
  assign n65338 = n52663 | n52664;
  assign n65339 = n52672 | n52673;
  assign n65340 = n52679 | n52680;
  assign n65341 = n52687 | ~n52688;
  assign n65342 = n52691 | n52692;
  assign n65343 = n52694 | n52695;
  assign n65344 = n52702 | n52703;
  assign n65345 = n52710 | n52711;
  assign n65346 = n52726 | ~n52727;
  assign n65347 = n52734 | n52735;
  assign n65348 = n52739 | n52740;
  assign n65349 = n52762 | n52763;
  assign n65350 = n52790 | ~n52791;
  assign n65351 = n52795 | n52792 | n52794;
  assign n65352 = n52799 | n52800;
  assign n65353 = n52803 | n52804;
  assign n65354 = n52807 | n52808;
  assign n65355 = n52815 | n52816;
  assign n65356 = n52819 | n52820;
  assign n65357 = n52828 | n52829;
  assign n65358 = n52833 | n52834;
  assign n65359 = n52841 | ~n52842;
  assign n65360 = n52878 | n52879;
  assign n65361 = n52902 | n52903;
  assign n65362 = n52913 | n52914;
  assign n65363 = n52937 | n52938;
  assign n65364 = n52944 | n52945;
  assign n65365 = n52952 | n52953;
  assign n65366 = n52965 | n52958 | n52964;
  assign n65367 = n52962 | n52963;
  assign n65368 = n52974 | n52971 | n52973;
  assign n65369 = n52979 | n52980;
  assign n65370 = n52992 | n52993;
  assign n65371 = n52996 | n52997;
  assign n65372 = n53013 | ~n53014;
  assign n65373 = n53016 | n53017;
  assign n65374 = n53039 | n53040;
  assign n65375 = n53042 | n53043;
  assign n65376 = n53046 | n53047;
  assign n65377 = n53060 | n53055 | n53059;
  assign n65378 = n53066 | n53067;
  assign n65379 = n53069 | n53070;
  assign n65380 = n53073 | n53074;
  assign n65381 = n53075 | n53076;
  assign n65382 = n53082 | n53083;
  assign n65383 = n53084 | n53085;
  assign n65384 = n53095 | n53096;
  assign n65385 = n53105 | n53106;
  assign n65386 = n53113 | n53114;
  assign n65387 = n53128 | n53129;
  assign n65388 = n53157 | n53158;
  assign n65389 = n53206 | n53207;
  assign n65390 = n53208 | n53209;
  assign n65391 = n53233 | n53234;
  assign n65392 = n53235 | n53236;
  assign n65393 = n53249 | n53250;
  assign n65394 = n53259 | n53260;
  assign n65395 = n53266 | n53267;
  assign n65396 = n53291 | n53292;
  assign n65397 = n53300 | n53301;
  assign n65398 = n53324 | n53325;
  assign n65399 = n53332 | n53333;
  assign n65400 = n53374 | n53375;
  assign n65401 = n53385 | n53386;
  assign n65402 = n53413 | n53414;
  assign n65403 = n53487 | n53488;
  assign n65404 = n53489 | ~n53490;
  assign n65405 = n53494 | ~n53495;
  assign n65406 = n53510 | ~n53511;
  assign n65407 = n53526 | n53527;
  assign n65408 = n53550 | n53541 | n53549;
  assign n65409 = n53544 | n53545;
  assign n65410 = n53562 | n53563;
  assign n65411 = n53571 | n53568 | n53570;
  assign n65412 = n53596 | n53597;
  assign n65413 = n53604 | n53605;
  assign n65414 = n53608 | n53609;
  assign n65415 = n53616 | n53617;
  assign n65416 = n53644 | n53645;
  assign n65417 = n53717 | n53718;
  assign n65418 = n53722 | n53719 | n53721;
  assign n65419 = n53730 | n53731;
  assign n65420 = n53754 | n53755;
  assign n65421 = n53784 | n53785;
  assign n65422 = n53816 | n53817;
  assign n65423 = n53821 | n53822;
  assign n65424 = n53838 | n53839;
  assign n65425 = n53849 | n53850;
  assign n65426 = n53873 | ~n53874;
  assign n65427 = n53916 | n53917;
  assign n65428 = n53922 | n53923;
  assign n65429 = n53957 | n53958;
  assign n65430 = n53965 | n53966;
  assign n65431 = n53972 | n53973;
  assign n65432 = n54036 | n54037;
  assign n65433 = n54040 | n54041;
  assign n65434 = n54054 | n54055;
  assign n65435 = n54070 | n54071;
  assign n65436 = n54089 | n54090;
  assign n65437 = n54114 | n54115;
  assign n65438 = n54123 | n54124;
  assign n65439 = n54146 | n54147;
  assign n65440 = n54152 | n54153;
  assign n65441 = n54168 | n54169;
  assign n65442 = n54184 | n54185;
  assign n65443 = n54189 | n54190;
  assign n65444 = n54195 | n54196;
  assign n65445 = n54202 | n54203;
  assign n65446 = n54257 | n54258;
  assign n65447 = n54268 | n54269;
  assign n65448 = n54272 | n54273;
  assign n65449 = n54355 | n54356;
  assign n65450 = n54359 | n54360;
  assign n65451 = n54394 | n54395;
  assign n65452 = n54411 | n54412;
  assign n65453 = n54419 | n54420;
  assign n65454 = n54425 | n54426;
  assign n65455 = n54470 | n54471;
  assign n65456 = n54482 | n54483;
  assign n65457 = n54486 | n54487;
  assign n65458 = ~n54491 | n54488 | n54490;
  assign n65459 = n54492 | n54493;
  assign n65460 = n54529 | n54530;
  assign n65461 = n54531 | n54532;
  assign n65462 = n54545 | n54546;
  assign n65463 = n54553 | n54551 | n54552;
  assign n65464 = n54555 | n54557 | n54558 | n54559;
  assign n65465 = n54560 | n54561;
  assign n65466 = n54579 | n54576 | n54578;
  assign n65467 = n54600 | n54601;
  assign n65468 = n54617 | n54618;
  assign n65469 = n54632 | n54633;
  assign n65470 = n54653 | ~n54654;
  assign n65471 = n54683 | n54684;
  assign n65472 = n54721 | n54722;
  assign n65473 = n54738 | n54739;
  assign n65474 = n54750 | n54751;
  assign n65475 = n54800 | n54801;
  assign n65476 = n54804 | n54805;
  assign n65477 = n54812 | n54813;
  assign n65478 = n54820 | n54821;
  assign n65479 = n54828 | n54829;
  assign n65480 = n54841 | n54842;
  assign n65481 = n54853 | n54854;
  assign n65482 = n54861 | n54862;
  assign n65483 = n54865 | n54866;
  assign n65484 = n54870 | n54871;
  assign n65485 = n54888 | n54889;
  assign n65486 = n54897 | n54898;
  assign n65487 = n54918 | n54919;
  assign n65488 = n54924 | n54925;
  assign n65489 = n54935 | n54932 | n54934;
  assign n65490 = n54980 | n54981;
  assign n65491 = n54990 | n54991;
  assign n65492 = n55015 | n55016;
  assign n65493 = n55040 | n55041;
  assign n65494 = n55066 | n55067;
  assign n65495 = n55088 | n55085 | n55087;
  assign n65496 = n55089 | n55090;
  assign n65497 = n55095 | n55096;
  assign n65498 = n55119 | n55120;
  assign n65499 = n55145 | ~n55146;
  assign n65500 = n55177 | n55178;
  assign n65501 = n55179 | n55180;
  assign n65502 = n55192 | ~n55193;
  assign n65503 = n55194 | n55195;
  assign n65504 = n55208 | n55209;
  assign n65505 = n55226 | n55227;
  assign n65506 = n55241 | n55242;
  assign n65507 = n55252 | ~n55253;
  assign n65508 = ~n55285 | n55262 | ~n55284;
  assign n65509 = n55265 | n55266;
  assign n65510 = n55279 | n55280;
  assign n65511 = n55290 | ~n55291;
  assign n65512 = n55340 | n55341;
  assign n65513 = n55348 | n55349;
  assign n65514 = n55370 | n55371;
  assign n65515 = n55377 | n55374 | n55376;
  assign n65516 = n55382 | n55383;
  assign n65517 = n55405 | n55406;
  assign n65518 = n55421 | n55422;
  assign n65519 = n55423 | n55424;
  assign n65520 = n55436 | n55437;
  assign n65521 = n55450 | n55451;
  assign n65522 = n55459 | ~n55460;
  assign n65523 = n55462 | n55463;
  assign n65524 = n55486 | n55487;
  assign n65525 = n55498 | n55499;
  assign n65526 = n55511 | n55512;
  assign n65527 = n55519 | n55520;
  assign n65528 = n55530 | n55531;
  assign n65529 = n55532 | n55533;
  assign n65530 = n55534 | n55535;
  assign n65531 = n55541 | n55539 | n55540;
  assign n65532 = n55555 | n55556;
  assign n65533 = n55564 | n55565;
  assign n65534 = n55571 | n55572;
  assign n65535 = n55587 | n55588;
  assign n65536 = n55590 | n55591;
  assign n65537 = n55598 | n55599;
  assign n65538 = n55605 | n55606;
  assign n65539 = n55617 | n55618;
  assign n65540 = n55626 | n55627;
  assign n65541 = n55638 | ~n55639;
  assign n65542 = n55654 | n55655;
  assign n65543 = n55658 | n55659;
  assign n65544 = n55666 | n55667;
  assign n65545 = n55676 | ~n55677;
  assign n65546 = n55682 | ~n55683;
  assign n65547 = n55707 | n55708;
  assign n65548 = n55724 | n55725;
  assign n65549 = n55728 | n55729;
  assign n65550 = n55731 | ~n55732;
  assign n65551 = n55759 | n55760;
  assign n65552 = n55772 | ~n55773;
  assign n65553 = n55780 | n55781;
  assign n65554 = n55786 | n55787;
  assign n65555 = n55805 | n55806;
  assign n65556 = n55831 | n55832;
  assign n65557 = n55839 | n55840;
  assign n65558 = n55857 | n55858;
  assign n65559 = n55887 | n55888;
  assign n65560 = n55908 | n55909;
  assign n65561 = n55914 | ~n55915;
  assign n65562 = n55932 | n55933;
  assign n65563 = n55940 | n55937 | n55939;
  assign n65564 = n55941 | n55942;
  assign n65565 = n55972 | n55973;
  assign n65566 = n55987 | n55975 | ~n55986;
  assign n65567 = n55980 | n55981;
  assign n65568 = n56018 | n56019;
  assign n65569 = n56020 | n56021;
  assign n65570 = n56085 | n56086;
  assign n65571 = n56094 | n56095;
  assign n65572 = n56102 | n56103;
  assign n65573 = n56133 | ~n56134;
  assign n65574 = n56139 | ~n56140;
  assign n65575 = n56168 | n56169;
  assign n65576 = n56183 | n56184;
  assign n65577 = n56237 | n56238;
  assign n65578 = n56259 | n56260;
  assign n65579 = n56274 | n56275;
  assign n65580 = n56281 | n56282;
  assign n65581 = n56286 | n56287;
  assign n65582 = n56300 | n56301;
  assign n65583 = n56304 | ~n56305;
  assign n65584 = n56362 | n56363;
  assign n65585 = n56368 | n56369;
  assign n65586 = n56381 | n56382;
  assign n65587 = n56385 | n56386;
  assign n65588 = n56395 | n56396;
  assign n65589 = n56411 | n56412;
  assign n65590 = n56416 | n56417;
  assign n65591 = n56420 | n56421;
  assign n65592 = n56440 | n56441;
  assign n65593 = n56450 | n56451;
  assign n65594 = n56470 | n56471;
  assign n65595 = n56477 | n56478;
  assign n65596 = n56484 | n56485;
  assign n65597 = n56489 | n56490;
  assign n65598 = n56504 | n56505;
  assign n65599 = n56509 | n56510;
  assign n65600 = n56514 | ~n56515;
  assign n65601 = n56520 | ~n56521;
  assign n65602 = n56529 | n56530;
  assign n65603 = n56563 | n56560 | n56562;
  assign n65604 = n56571 | n56572;
  assign n65605 = n56609 | n56610;
  assign n65606 = n56656 | n56657;
  assign n65607 = n56660 | n56661;
  assign n65608 = n56675 | n56676;
  assign n65609 = ~n56687 | n56681 | ~n56686;
  assign n65610 = n56737 | n56738;
  assign n65611 = n56748 | n56749;
  assign n65612 = n56752 | n56753;
  assign n65613 = n56764 | n56765;
  assign n65614 = n56772 | n56773;
  assign n65615 = n56800 | n56801;
  assign n65616 = n56809 | n56810;
  assign n65617 = n56823 | ~n56824;
  assign n65618 = n56829 | ~n56830;
  assign n65619 = n56831 | n56832;
  assign n65620 = n56851 | n56852;
  assign n65621 = n56860 | n56861;
  assign n65622 = n56864 | n56865;
  assign n65623 = n56866 | n56867;
  assign n65624 = n56888 | n56889;
  assign n65625 = n56894 | n56895;
  assign n65626 = n56905 | n56906;
  assign n65627 = n56921 | n56922;
  assign n65628 = n56926 | n56927;
  assign n65629 = n56936 | ~n56937;
  assign n65630 = n56946 | n56947;
  assign n65631 = n56957 | ~n56958;
  assign n65632 = n56968 | n56969;
  assign n65633 = n56970 | n56971;
  assign n65634 = n56993 | n56994;
  assign n65635 = n57019 | n57020;
  assign n65636 = n57034 | n57035;
  assign n65637 = n57060 | ~n57061;
  assign n65638 = n57066 | ~n57067;
  assign n65639 = n57081 | n57082;
  assign n65640 = n57090 | ~n57091;
  assign n65641 = n57113 | n57114;
  assign n65642 = n57150 | n57147 | n57149;
  assign n65643 = n57159 | n57160;
  assign n65644 = n57163 | n57164;
  assign n65645 = n57185 | n57186;
  assign n65646 = n57266 | ~n57267;
  assign n65647 = n57277 | n57278;
  assign n65648 = ~n57307 | n57294 | ~n57306;
  assign n65649 = n57301 | n57302;
  assign n65650 = n57312 | ~n57313;
  assign n65651 = n57389 | n57390;
  assign n65652 = n57403 | n57404;
  assign n65653 = n57425 | n57426;
  assign n65654 = n57432 | n57433;
  assign n65655 = n57441 | n57442;
  assign n65656 = n57451 | n57452;
  assign n65657 = n57457 | n57458;
  assign n65658 = n57469 | n57470;
  assign n65659 = n57485 | n57486;
  assign n65660 = n57491 | n57492;
  assign n65661 = n57498 | n57499;
  assign n65662 = n57506 | n57507;
  assign n65663 = n57512 | n57513;
  assign n65664 = n57524 | n57525;
  assign n65665 = n57541 | n57542;
  assign n65666 = n57556 | n57557;
  assign n65667 = n57567 | n57568;
  assign n65668 = n57575 | n57576;
  assign n65669 = n57604 | n57605;
  assign n65670 = n57632 | n57633;
  assign n65671 = n57647 | n57648;
  assign n65672 = n57658 | n57659;
  assign n65673 = n57677 | n57678;
  assign n65674 = n57686 | n57687;
  assign n65675 = n57689 | n57690;
  assign n65676 = n57700 | n57701;
  assign n65677 = n57705 | n57706;
  assign n65678 = n57716 | n57717;
  assign n65679 = n57718 | ~n57719;
  assign n65680 = n57722 | n57723;
  assign n65681 = n57726 | ~n57727;
  assign n65682 = n57731 | n57732;
  assign n65683 = n57738 | n57739;
  assign n65684 = n57746 | n57747;
  assign n65685 = n57752 | n57753;
  assign n65686 = n57762 | n57763;
  assign n65687 = n57771 | n57772;
  assign n65688 = n57804 | n57805;
  assign n65689 = n57806 | n57807;
  assign n65690 = n57816 | n57817;
  assign n65691 = n57823 | n57824;
  assign n65692 = n57831 | n57832;
  assign n65693 = n57837 | n57838;
  assign n65694 = n57848 | n57849;
  assign n65695 = n57864 | n57865;
  assign n65696 = n57870 | n57871;
  assign n65697 = n57877 | n57878;
  assign n65698 = n57885 | n57886;
  assign n65699 = n57903 | ~n57904;
  assign n65700 = n57927 | n57928;
  assign n65701 = n57955 | n57956;
  assign n65702 = n57964 | n57965;
  assign n65703 = n58009 | n58010;
  assign n65704 = n58022 | n58023;
  assign n65705 = n58033 | n58034;
  assign n65706 = n58056 | n58057;
  assign n65707 = n58058 | ~n58059;
  assign n65708 = n58072 | n58073;
  assign n65709 = n58079 | ~n58080;
  assign n65710 = n58093 | n58094;
  assign n65711 = n58105 | n58106;
  assign n65712 = n58136 | n58137;
  assign n65713 = n58149 | n58150;
  assign n65714 = n58448 | n58449;
  assign n65715 = n58472 | n58473;
  assign po468 = n58480 | n58481;
  assign po215 = n58494 | n58495;
  assign po217 = n58502 | n58503;
  assign n65719 = n58507 | n58508;
  assign n65720 = n58598 | n58599;
  assign n65721 = n58644 | n58645;
  assign n65722 = n58664 | n58665;
  assign n65723 = n58700 | ~n58701;
  assign n65724 = n58710 | n58711;
  assign n65725 = n58740 | n58741;
  assign po1105 = n58782 | ~n58783;
  assign n65727 = n58784 | n58785;
  assign po459 = n58807 | n58808;
  assign n65729 = n58825 | n58826;
  assign n65730 = n58829 | n58830;
  assign n65731 = n58852 | n58853;
  assign n65732 = n58859 | n58860;
  assign n65733 = n58872 | n58873;
  assign po622 = n58881 | ~n58882;
  assign n65735 = n58887 | ~n58888;
  assign n65736 = n58901 | ~n58902;
  assign n65737 = n58906 | n58907;
  assign n65738 = n58923 | n58924;
  assign n65739 = n58934 | n58935;
  assign po626 = n58943 | ~n58944;
  assign n65741 = n58959 | n58960;
  assign n65742 = n58970 | n58971;
  assign po627 = n58979 | ~n58980;
  assign n65744 = n58995 | n58996;
  assign n65745 = n59006 | n59007;
  assign po628 = n59015 | ~n59016;
  assign n65747 = n59031 | n59032;
  assign n65748 = n59042 | n59043;
  assign po629 = n59051 | ~n59052;
  assign n65750 = n59063 | n59064;
  assign n65751 = n59076 | n59077;
  assign n65752 = n59089 | n59090;
  assign n65753 = n59108 | ~n59109;
  assign n65754 = n59115 | n59116;
  assign n65755 = n59121 | n59122;
  assign n65756 = n59127 | n59128;
  assign n65757 = n59171 | ~n59172;
  assign n65758 = n59177 | ~n59178;
  assign n65759 = n59184 | n59185;
  assign n65760 = n59187 | n59188;
  assign n65761 = n59205 | n59206;
  assign n65762 = n59233 | n59234;
  assign n65763 = n59387 | ~n59388;
  assign n65764 = n59399 | ~n59400;
  assign n65765 = n59414 | n59410 | n59413;
  assign n65766 = n59418 | n59419;
  assign n65767 = n59422 | n59423;
  assign n65768 = n59424 | n59425;
  assign n65769 = n59462 | ~n59463;
  assign n65770 = n59469 | ~n59470;
  assign n65771 = n59477 | ~n59478;
  assign n65772 = n59484 | n59489 | n59492 | n59493;
  assign n65773 = n59496 | n59497;
  assign n65774 = n59542 | n59543;
  assign n65775 = n59665 | ~n59666;
  assign n65776 = n59671 | ~n59672;
  assign n65777 = n59675 | n59676;
  assign n65778 = n59679 | n59680;
  assign n65779 = n59718 | ~n59719;
  assign n65780 = n59724 | ~n59725;
  assign n65781 = n59728 | n59729;
  assign n65782 = n59732 | n59733;
  assign n65783 = n59771 | n59772;
  assign n65784 = n59925 | ~n59926;
  assign n65785 = n59929 | ~n59930;
  assign n65786 = n59940 | n59941;
  assign n65787 = n59945 | ~n59946;
  assign n65788 = n59949 | ~n59950;
  assign n65789 = n59959 | n59960;
  assign n65790 = n59963 | n59964;
  assign n65791 = n59969 | n59970;
  assign n65792 = n59975 | n59976;
  assign n65793 = n60028 | ~n60029;
  assign n65794 = n60041 | n60042;
  assign n65795 = n60058 | n60059;
  assign n65796 = n60063 | n60064;
  assign n65797 = n60068 | n60069;
  assign n65798 = n60070 | n60071;
  assign n65799 = n60073 | n60074;
  assign n65800 = n60094 | n60095;
  assign n65801 = n60120 | n60121;
  assign n65802 = n60228 | n60229;
  assign n65803 = n60272 | n60273;
  assign n65804 = n60313 | n60314;
  assign po782 = n60380 | n60381;
  assign po784 = n60386 | n60387;
  assign po785 = n60392 | n60393;
  assign po897 = n60400 | n60401;
  assign po786 = n60406 | n60407;
  assign po787 = n60412 | n60413;
  assign po788 = n60418 | n60419;
  assign po789 = n60424 | n60425;
  assign po790 = n60430 | n60431;
  assign po791 = n60436 | n60437;
  assign po792 = n60442 | n60443;
  assign po793 = n60448 | n60449;
  assign po794 = n60454 | n60455;
  assign po795 = n60460 | n60461;
  assign po796 = n60466 | n60467;
  assign po797 = n60472 | n60473;
  assign po798 = n60478 | n60479;
  assign po800 = n60484 | n60485;
  assign po801 = n60490 | n60491;
  assign po802 = n60496 | n60497;
  assign po803 = n60502 | n60503;
  assign po804 = n60508 | n60509;
  assign po805 = n60514 | n60515;
  assign po806 = n60520 | n60521;
  assign po807 = n60526 | n60527;
  assign po808 = n60532 | n60533;
  assign po809 = n60538 | n60539;
  assign po810 = n60544 | n60545;
  assign po811 = n60550 | n60551;
  assign po812 = n60556 | n60557;
  assign po813 = n60562 | n60563;
  assign po814 = n60568 | n60569;
  assign po815 = n60574 | n60575;
  assign po817 = n60580 | n60581;
  assign po818 = n60586 | n60587;
  assign po819 = n60592 | n60593;
  assign po822 = n60598 | n60599;
  assign po826 = n60604 | n60605;
  assign po837 = n60610 | n60611;
  assign po838 = n60616 | n60617;
  assign po841 = n60623 | n60624;
  assign po843 = n60629 | n60630;
  assign po844 = n60635 | n60636;
  assign po845 = n60641 | n60642;
  assign po847 = n60647 | n60648;
  assign po848 = n60653 | n60654;
  assign po850 = n60659 | n60660;
  assign po851 = n60665 | n60666;
  assign po852 = n60671 | n60672;
  assign po853 = n60677 | n60678;
  assign po854 = n60683 | n60684;
  assign po855 = n60689 | n60690;
  assign po856 = n60695 | n60696;
  assign po857 = n60701 | n60702;
  assign po858 = n60707 | n60708;
  assign po859 = n60713 | n60714;
  assign po860 = n60719 | n60720;
  assign po861 = n60725 | n60726;
  assign po862 = n60731 | n60732;
  assign po863 = n60737 | n60738;
  assign po866 = n60743 | n60744;
  assign po867 = n60749 | n60750;
  assign po872 = n60755 | n60756;
  assign po880 = n60761 | n60762;
  assign po881 = n60767 | n60768;
  assign po882 = n60773 | n60774;
  assign po883 = n60779 | n60780;
  assign po884 = n60785 | n60786;
  assign po885 = n60791 | n60792;
  assign po886 = n60797 | n60798;
  assign po887 = n60803 | n60804;
  assign po889 = n60809 | n60810;
  assign po891 = n60815 | n60816;
  assign po892 = n60821 | n60822;
  assign po893 = n60827 | n60828;
  assign po894 = n60833 | n60834;
  assign po895 = n60839 | n60840;
  assign po988 = n60844 | n60845;
  assign n65883 = n60850 | n60851;
  assign n65884 = n60856 | n60857;
  assign n65885 = n60862 | n60863;
  assign n65886 = n60868 | n60869;
  assign n65887 = n60874 | n60875;
  assign n65888 = n60880 | n60881;
  assign n65889 = n60886 | n60887;
  assign n65890 = n60892 | n60893;
  assign n65891 = n60898 | n60899;
  assign n65892 = n60904 | n60905;
  assign n65893 = n60910 | n60911;
  assign n65894 = n60916 | n60917;
  assign n65895 = n60930 | ~n60931;
  assign n65896 = n60936 | ~n60937;
  assign n65897 = n60942 | ~n60943;
  assign n65898 = n60961 | n60954 | n60960;
  assign n65899 = n60979 | ~n60980;
  assign n65900 = n60985 | ~n60986;
  assign n65901 = n60991 | ~n60992;
  assign n65902 = n61010 | n61003 | n61009;
  assign n65903 = n61028 | ~n61029;
  assign n65904 = n61034 | ~n61035;
  assign n65905 = n61040 | ~n61041;
  assign n65906 = n61059 | n61052 | n61058;
  assign n65907 = n61077 | ~n61078;
  assign n65908 = n61083 | ~n61084;
  assign n65909 = n61089 | ~n61090;
  assign n65910 = n61108 | n61101 | n61107;
  assign n65911 = n61116 | n61117;
  assign n65912 = n61121 | n61122;
  assign n65913 = n61131 | ~n61132;
  assign n65914 = n61137 | ~n61138;
  assign n65915 = n61143 | n61144;
  assign n65916 = n61150 | n61151;
  assign n65917 = n61157 | ~n61158;
  assign n65918 = n61163 | ~n61164;
  assign po764 = n61178 | n61179;
  assign po765 = n61184 | n61185;
  assign po766 = n61190 | n61191;
  assign po767 = n61196 | n61197;
  assign po768 = n61202 | n61203;
  assign po769 = n61208 | n61209;
  assign po770 = n61214 | n61215;
  assign po775 = n61220 | n61221;
  assign po776 = n61226 | n61227;
  assign po777 = n61232 | n61233;
  assign po778 = n61238 | n61239;
  assign po779 = n61244 | n61245;
  assign po780 = n61250 | n61251;
  assign po783 = n61262 | n61263;
  assign po799 = n61268 | n61269;
  assign n65934 = n61274 | n61275;
  assign n65935 = n61280 | n61281;
  assign n65936 = n61286 | n61287;
  assign n65937 = n61292 | n61293;
  assign n65938 = n61298 | n61299;
  assign n65939 = n61304 | n61305;
  assign n65940 = n61312 | n61313;
  assign n65941 = n61318 | n61319;
  assign n65942 = n61324 | n61325;
  assign n65943 = n61330 | n61331;
  assign n65944 = n61336 | n61337;
  assign n65945 = n61342 | n61343;
  assign n65946 = n61348 | n61349;
  assign n65947 = n61354 | n61355;
  assign n65948 = n61360 | n61361;
  assign n65949 = n61366 | n61367;
  assign n65950 = n61372 | n61373;
  assign n65951 = n61378 | n61379;
  assign n65952 = n61384 | n61385;
  assign n65953 = n61390 | n61391;
  assign n65954 = n61400 | n61401;
  assign n65955 = n61407 | n61408;
  assign po1063 = n61411 | n61412;
  assign n65957 = n61419 | ~n61420;
  assign n65958 = n61425 | ~n61426;
  assign n65959 = n61431 | ~n61432;
  assign n65960 = n61437 | ~n61438;
  assign n65961 = n61443 | ~n61444;
  assign n65962 = n61449 | ~n61450;
  assign n65963 = n61455 | ~n61456;
  assign n65964 = n61461 | ~n61462;
  assign n65965 = n61467 | ~n61468;
  assign n65966 = n61473 | ~n61474;
  assign po455 = n61495 | ~n61496;
  assign po460 = n61501 | ~n61502;
  assign po461 = n61507 | ~n61508;
  assign po462 = n61513 | ~n61514;
  assign po463 = n61519 | ~n61520;
  assign po464 = n61525 | ~n61526;
  assign po465 = n61531 | ~n61532;
  assign po466 = n61537 | ~n61538;
  assign n65975 = n61554 | n61555;
  assign n65976 = n61561 | n61562;
  assign po745 = n61575 | n61576;
  assign n65978 = n61581 | n61582;
  assign po748 = n61587 | n61588;
  assign po749 = n61593 | n61594;
  assign po752 = n61610 | n61611;
  assign po754 = n61620 | n61621;
  assign po758 = n61633 | n61634;
  assign n65984 = n61645 | ~n61646;
  assign n65985 = n61660 | n61661;
  assign n65986 = n61666 | ~n61667;
  assign n65987 = n61690 | ~n61691;
  assign n65988 = n61697 | n61698;
  assign n65989 = n61706 | n61707;
  assign n65990 = n61716 | n61717;
  assign n65991 = n61719 | n61720;
  assign n65992 = n61723 | n61724;
  assign n65993 = n61732 | n61733;
  assign n65994 = n61740 | n61741;
  assign po888 = n61752 | n61753;
  assign n65996 = n61768 | n61769;
  assign n65997 = n61779 | n61780;
  assign n65998 = n61795 | n61796;
  assign n65999 = n61817 | n61818;
  assign n66000 = n61833 | n61834;
  assign n66001 = n61848 | n61849;
  assign n66002 = n61857 | n61858;
  assign po993 = n61958 | ~n61959;
  assign po994 = n61964 | ~n61965;
  assign po995 = n61970 | ~n61971;
  assign po998 = n61976 | ~n61977;
  assign po999 = n61982 | ~n61983;
  assign po1000 = n61988 | ~n61989;
  assign po1001 = n61994 | ~n61995;
  assign po1003 = n62000 | ~n62001;
  assign po1004 = n62006 | ~n62007;
  assign po1006 = n62012 | ~n62013;
  assign po1007 = n62018 | ~n62019;
  assign po1008 = n62024 | ~n62025;
  assign po1009 = n62030 | ~n62031;
  assign po1010 = n62036 | ~n62037;
  assign po1011 = n62042 | ~n62043;
  assign po1012 = n62048 | ~n62049;
  assign po1013 = n62054 | ~n62055;
  assign po1014 = n62060 | ~n62061;
  assign po1015 = n62066 | ~n62067;
  assign po1016 = n62072 | ~n62073;
  assign po1021 = n62078 | ~n62079;
  assign po1022 = n62084 | ~n62085;
  assign po1023 = n62090 | ~n62091;
  assign po1024 = n62096 | ~n62097;
  assign po1026 = n62102 | ~n62103;
  assign po1027 = n62108 | ~n62109;
  assign po1028 = n62114 | ~n62115;
  assign po1029 = n62120 | ~n62121;
  assign po1030 = n62126 | ~n62127;
  assign po1032 = n62132 | ~n62133;
  assign po1036 = n62138 | ~n62139;
  assign po1037 = n62144 | ~n62145;
  assign n66035 = n62244 | n62245;
  assign n66036 = n62257 | n62258;
  assign n66037 = n62267 | n62268;
  assign n66038 = n62277 | n62278;
  assign n66039 = n62287 | n62288;
  assign n66040 = n62297 | n62298;
  assign n66041 = n62317 | ~n62318;
  assign po0 = pi668;
  assign po1 = pi672;
  assign po2 = pi664;
  assign po3 = pi667;
  assign po4 = pi676;
  assign po5 = pi673;
  assign po6 = pi675;
  assign po7 = pi666;
  assign po8 = pi679;
  assign po9 = pi674;
  assign po10 = pi663;
  assign po11 = pi670;
  assign po12 = pi677;
  assign po13 = pi682;
  assign po14 = pi671;
  assign po15 = pi678;
  assign po16 = pi718;
  assign po17 = pi707;
  assign po18 = pi708;
  assign po19 = pi713;
  assign po20 = pi711;
  assign po21 = pi716;
  assign po22 = pi733;
  assign po23 = pi712;
  assign po24 = pi689;
  assign po25 = pi717;
  assign po26 = pi692;
  assign po27 = pi719;
  assign po28 = pi722;
  assign po29 = pi714;
  assign po30 = pi720;
  assign po31 = pi685;
  assign po32 = pi837;
  assign po33 = pi850;
  assign po34 = pi872;
  assign po35 = pi871;
  assign po36 = pi881;
  assign po37 = pi866;
  assign po38 = pi876;
  assign po39 = pi873;
  assign po40 = pi874;
  assign po41 = pi859;
  assign po42 = pi855;
  assign po43 = pi852;
  assign po44 = pi870;
  assign po45 = pi848;
  assign po46 = pi865;
  assign po47 = pi856;
  assign po48 = pi853;
  assign po49 = pi847;
  assign po50 = pi857;
  assign po51 = pi854;
  assign po52 = pi858;
  assign po53 = pi845;
  assign po54 = pi838;
  assign po55 = pi842;
  assign po56 = pi843;
  assign po57 = pi839;
  assign po58 = pi844;
  assign po59 = pi868;
  assign po60 = pi851;
  assign po61 = pi867;
  assign po62 = pi880;
  assign po63 = pi860;
  assign po64 = pi1030;
  assign po65 = pi1034;
  assign po66 = pi1015;
  assign po67 = pi1020;
  assign po68 = pi1025;
  assign po69 = pi1005;
  assign po70 = pi996;
  assign po71 = pi1012;
  assign po72 = pi993;
  assign po73 = pi1016;
  assign po74 = pi1021;
  assign po75 = pi1010;
  assign po76 = pi1027;
  assign po77 = pi1018;
  assign po78 = pi1017;
  assign po79 = pi1024;
  assign po80 = pi1009;
  assign po81 = pi1032;
  assign po82 = pi1003;
  assign po83 = pi997;
  assign po84 = pi1013;
  assign po85 = pi1011;
  assign po86 = pi1008;
  assign po87 = pi1019;
  assign po88 = pi1031;
  assign po89 = pi1022;
  assign po90 = pi1000;
  assign po91 = pi1023;
  assign po92 = pi1002;
  assign po93 = pi1026;
  assign po94 = pi1006;
  assign po95 = pi998;
  assign po96 = pi31;
  assign po97 = pi80;
  assign po98 = pi893;
  assign po99 = pi467;
  assign po100 = pi78;
  assign po101 = pi112;
  assign po102 = pi13;
  assign po103 = pi25;
  assign po104 = pi226;
  assign po105 = pi127;
  assign po106 = pi822;
  assign po107 = pi808;
  assign po108 = pi227;
  assign po109 = pi477;
  assign po110 = pi834;
  assign po111 = pi229;
  assign po112 = pi12;
  assign po113 = pi11;
  assign po114 = pi10;
  assign po115 = pi9;
  assign po116 = pi8;
  assign po117 = pi7;
  assign po118 = pi6;
  assign po119 = pi5;
  assign po120 = pi4;
  assign po121 = pi3;
  assign po122 = pi0;
  assign po123 = pi2;
  assign po124 = pi1;
  assign po125 = pi310;
  assign po126 = pi302;
  assign po127 = pi475;
  assign po128 = pi474;
  assign po129 = pi466;
  assign po130 = pi473;
  assign po131 = pi471;
  assign po132 = pi472;
  assign po133 = pi470;
  assign po134 = pi469;
  assign po135 = pi465;
  assign po136 = pi1028;
  assign po137 = pi1033;
  assign po138 = pi995;
  assign po139 = pi994;
  assign po140 = pi28;
  assign po141 = pi27;
  assign po142 = pi26;
  assign po143 = pi29;
  assign po144 = pi15;
  assign po145 = pi14;
  assign po146 = pi21;
  assign po147 = pi20;
  assign po148 = pi19;
  assign po149 = pi18;
  assign po150 = pi17;
  assign po151 = pi16;
  assign po152 = pi1096;
  assign po153 = ~n41712;
  assign po154 = ~n46152;
  assign po157 = ~n44573;
  assign po160 = ~n45329;
  assign po163 = ~n46862;
  assign po164 = ~n47114;
  assign po168 = pi228;
  assign po169 = pi22;
  assign po170 = ~pi1090;
  assign po179 = pi1089;
  assign po180 = pi23;
  assign po181 = po167;
  assign po183 = ~n48068;
  assign po184 = ~n61481;
  assign po185 = ~n61483;
  assign po186 = ~n61485;
  assign po187 = ~n61487;
  assign po188 = pi37;
  assign po189 = ~n5537;
  assign po200 = ~n39419;
  assign po201 = ~n39631;
  assign po202 = ~n40418;
  assign po237 = ~n32930;
  assign po257 = ~n40495;
  assign po259 = ~n40589;
  assign po263 = pi117;
  assign po270 = ~n61490;
  assign po276 = ~n33320;
  assign po277 = ~n35428;
  assign po278 = ~n31346;
  assign po279 = ~n42275;
  assign po280 = ~n33855;
  assign po282 = ~n42797;
  assign po283 = ~n64836;
  assign po285 = pi131;
  assign po289 = ~n43523;
  assign po290 = ~n43950;
  assign po291 = ~n44084;
  assign po292 = ~n44207;
  assign po293 = ~n44300;
  assign po294 = ~n48022;
  assign po303 = ~n35568;
  assign po305 = ~n35814;
  assign po309 = ~n36179;
  assign po310 = ~n36288;
  assign po318 = ~n36852;
  assign po323 = ~n37228;
  assign po325 = ~n37394;
  assign po326 = ~n37503;
  assign po327 = ~n37584;
  assign po328 = ~n37693;
  assign po329 = ~n37798;
  assign po352 = ~n35261;
  assign po353 = ~n35345;
  assign po355 = ~n28298;
  assign po366 = ~n27522;
  assign po368 = ~n37922;
  assign po369 = ~n37947;
  assign po370 = ~n37984;
  assign po371 = ~n38009;
  assign po372 = ~n38419;
  assign po374 = ~n27541;
  assign po376 = ~n38044;
  assign po380 = ~n64037;
  assign po384 = ~n39920;
  assign po385 = ~n38984;
  assign po386 = pi232;
  assign po388 = pi236;
  assign po390 = ~n53006;
  assign po391 = ~n54073;
  assign po394 = ~n53346;
  assign po395 = ~n54660;
  assign po397 = ~n65511;
  assign po398 = ~n65546;
  assign po402 = ~n65574;
  assign po403 = ~n65601;
  assign po404 = ~n65618;
  assign po405 = ~n65638;
  assign po406 = ~n65650;
  assign po408 = ~n52158;
  assign po412 = ~n65293;
  assign po413 = ~n65294;
  assign po414 = ~n65295;
  assign po415 = ~n65296;
  assign po416 = ~n65297;
  assign po417 = ~n52191;
  assign po418 = ~n52194;
  assign po419 = ~n58745;
  assign po421 = ~n57493;
  assign po422 = ~n57543;
  assign po425 = ~n65323;
  assign po427 = ~n57733;
  assign po430 = ~n57391;
  assign po432 = ~n65405;
  assign po433 = ~n57818;
  assign po434 = ~n57872;
  assign po437 = ~n65709;
  assign po441 = ~n58749;
  assign po447 = ~n65298;
  assign po448 = ~n65299;
  assign po449 = ~n65300;
  assign po450 = ~n65301;
  assign po451 = ~n65302;
  assign po452 = ~n65303;
  assign po453 = ~n65304;
  assign po454 = ~n65305;
  assign po457 = ~n58505;
  assign po458 = ~n58484;
  assign po467 = ~n58838;
  assign po472 = ~n48243;
  assign po473 = ~n48246;
  assign po474 = ~n48249;
  assign po475 = ~n48254;
  assign po476 = ~n48257;
  assign po477 = ~n48260;
  assign po478 = ~n48263;
  assign po479 = ~n48266;
  assign po480 = ~n48269;
  assign po481 = ~n48272;
  assign po482 = ~n48275;
  assign po483 = ~n48278;
  assign po484 = ~n48281;
  assign po485 = ~n48284;
  assign po486 = ~n48287;
  assign po487 = ~n48152;
  assign po488 = ~n48162;
  assign po490 = ~n48290;
  assign po491 = ~n48293;
  assign po492 = ~n48296;
  assign po493 = ~n58169;
  assign po494 = ~n58172;
  assign po495 = ~n48299;
  assign po496 = ~n48302;
  assign po499 = ~n58175;
  assign po500 = ~n58178;
  assign po501 = ~n48305;
  assign po502 = ~n58181;
  assign po503 = ~n58184;
  assign po504 = ~n58187;
  assign po505 = ~n58190;
  assign po506 = ~n48308;
  assign po507 = ~n58193;
  assign po508 = ~n58196;
  assign po509 = ~n48311;
  assign po510 = ~n48314;
  assign po511 = ~n58199;
  assign po512 = ~n58202;
  assign po513 = ~n58205;
  assign po514 = ~n58208;
  assign po515 = ~n58211;
  assign po516 = ~n58214;
  assign po517 = ~n58217;
  assign po518 = ~n58220;
  assign po519 = ~n58223;
  assign po520 = ~n58226;
  assign po521 = ~n58229;
  assign po522 = ~n48317;
  assign po523 = ~n48320;
  assign po524 = ~n58232;
  assign po525 = ~n58235;
  assign po526 = ~n48323;
  assign po527 = ~n58238;
  assign po528 = ~n48326;
  assign po529 = ~n48329;
  assign po530 = ~n58241;
  assign po531 = ~n58244;
  assign po532 = ~n48332;
  assign po533 = ~n58247;
  assign po534 = ~n48335;
  assign po535 = ~n48338;
  assign po536 = ~n58250;
  assign po537 = ~n58253;
  assign po538 = ~n58256;
  assign po539 = ~n58259;
  assign po540 = ~n58262;
  assign po541 = ~n58265;
  assign po542 = ~n58268;
  assign po543 = ~n58271;
  assign po544 = ~n58274;
  assign po545 = ~n58277;
  assign po546 = ~n58280;
  assign po547 = ~n58283;
  assign po548 = ~n58286;
  assign po549 = ~n58289;
  assign po550 = ~n58292;
  assign po551 = ~n48341;
  assign po552 = ~n58295;
  assign po553 = ~n48344;
  assign po554 = ~n48347;
  assign po555 = ~n58298;
  assign po556 = ~n48350;
  assign po557 = ~n58301;
  assign po558 = ~n58304;
  assign po559 = ~n48353;
  assign po560 = ~n58307;
  assign po561 = ~n58310;
  assign po562 = ~n58313;
  assign po563 = ~n58316;
  assign po564 = ~n58319;
  assign po565 = ~n58322;
  assign po566 = ~n58325;
  assign po567 = ~n58328;
  assign po568 = ~n58331;
  assign po569 = ~n58334;
  assign po570 = ~n58337;
  assign po571 = ~n58340;
  assign po572 = ~n58343;
  assign po573 = ~n48357;
  assign po574 = ~n58346;
  assign po575 = ~n58349;
  assign po576 = ~n48360;
  assign po577 = ~n58352;
  assign po578 = ~n48363;
  assign po579 = ~n48366;
  assign po580 = ~n58355;
  assign po581 = ~n48369;
  assign po582 = ~n58358;
  assign po583 = ~n58361;
  assign po584 = ~n48372;
  assign po585 = ~n58364;
  assign po586 = ~n58367;
  assign po587 = ~n58370;
  assign po588 = ~n58373;
  assign po589 = ~n58376;
  assign po590 = ~n58379;
  assign po591 = ~n58382;
  assign po592 = ~n58385;
  assign po593 = ~n58388;
  assign po594 = ~n58391;
  assign po595 = ~n58394;
  assign po596 = ~n48375;
  assign po597 = ~n48378;
  assign po598 = ~n58397;
  assign po599 = ~n48381;
  assign po600 = ~n58400;
  assign po601 = ~n48384;
  assign po602 = ~n58403;
  assign po603 = ~n48387;
  assign po604 = ~n48390;
  assign po605 = ~n48393;
  assign po606 = ~n48396;
  assign po607 = ~n58406;
  assign po608 = ~n48399;
  assign po609 = ~n58409;
  assign po610 = ~n48402;
  assign po611 = ~n48405;
  assign po612 = ~n58412;
  assign po613 = ~n58415;
  assign po615 = ~n48408;
  assign po616 = ~n48411;
  assign po617 = ~n48414;
  assign po618 = ~n48417;
  assign po619 = ~n48420;
  assign po620 = ~n58418;
  assign po621 = ~n48423;
  assign po625 = ~n48457;
  assign po633 = ~n48566;
  assign po634 = ~n48508;
  assign po636 = pi583;
  assign po638 = ~n58520;
  assign po639 = ~n58523;
  assign po640 = ~n58526;
  assign po641 = ~n58529;
  assign po642 = ~n58532;
  assign po643 = ~n58535;
  assign po644 = ~n58538;
  assign po646 = ~n58544;
  assign po647 = ~n58547;
  assign po648 = ~n58550;
  assign po649 = ~n58553;
  assign po650 = ~n58556;
  assign po652 = ~n58562;
  assign po653 = ~n58565;
  assign po655 = ~n58571;
  assign po656 = ~n58574;
  assign po657 = ~n58577;
  assign po658 = ~n58580;
  assign po659 = ~n58583;
  assign po660 = ~n58586;
  assign po661 = ~n58589;
  assign po662 = ~n65720;
  assign po663 = ~n58602;
  assign po664 = ~n58605;
  assign po665 = ~n58608;
  assign po666 = ~n58611;
  assign po667 = ~n58614;
  assign po668 = ~n58618;
  assign po669 = ~n58621;
  assign po670 = ~n58624;
  assign po671 = ~n58627;
  assign po672 = ~n58630;
  assign po673 = ~n58633;
  assign po674 = ~n58636;
  assign po675 = ~n65721;
  assign po677 = ~n58651;
  assign po678 = ~n58654;
  assign po679 = ~n58657;
  assign po680 = ~n65722;
  assign po682 = ~n58671;
  assign po683 = ~n58674;
  assign po684 = ~n58677;
  assign po685 = ~n58680;
  assign po686 = ~n58683;
  assign po687 = ~n58686;
  assign po688 = ~n58689;
  assign po689 = ~n58692;
  assign po690 = ~n58695;
  assign po692 = ~n60197;
  assign po693 = ~n60200;
  assign po694 = ~n60203;
  assign po695 = ~n60206;
  assign po696 = ~n60209;
  assign po697 = ~n60212;
  assign po698 = ~n60215;
  assign po699 = ~n60218;
  assign po700 = ~n60221;
  assign po701 = ~n65802;
  assign po702 = ~n60232;
  assign po703 = ~n60235;
  assign po704 = ~n60238;
  assign po705 = ~n60241;
  assign po706 = ~n60244;
  assign po708 = ~n60250;
  assign po709 = ~n60253;
  assign po710 = ~n60256;
  assign po711 = ~n60259;
  assign po712 = ~n60262;
  assign po713 = ~n60265;
  assign po714 = ~n65803;
  assign po715 = ~n60276;
  assign po716 = ~n60279;
  assign po717 = ~n60282;
  assign po718 = ~n60285;
  assign po719 = ~n60288;
  assign po720 = ~n60291;
  assign po721 = ~n60294;
  assign po722 = ~n60297;
  assign po723 = ~n60300;
  assign po724 = ~n65101;
  assign po725 = ~n60303;
  assign po727 = ~n65804;
  assign po728 = ~n60317;
  assign po729 = ~n60320;
  assign po730 = ~n60323;
  assign po731 = ~n60326;
  assign po732 = ~n60329;
  assign po733 = ~n60332;
  assign po734 = ~n60335;
  assign po735 = ~n60338;
  assign po736 = ~n60341;
  assign po737 = ~n60344;
  assign po738 = ~n60347;
  assign po739 = ~n60350;
  assign po741 = ~n60353;
  assign po742 = ~n60356;
  assign po743 = ~n60359;
  assign po744 = ~n50505;
  assign po747 = ~n65978;
  assign po755 = ~n60365;
  assign po759 = ~n50522;
  assign po760 = ~n61126;
  assign po761 = ~n61173;
  assign po763 = ~n65914;
  assign po771 = ~n61145;
  assign po772 = ~n60370;
  assign po773 = ~n61152;
  assign po774 = ~n65918;
  assign po781 = ~n61257;
  assign po820 = ~n51840;
  assign po821 = ~n51885;
  assign po823 = ~n51927;
  assign po824 = ~n51972;
  assign po825 = ~n50817;
  assign po827 = ~n52008;
  assign po828 = ~n52044;
  assign po829 = ~n50859;
  assign po830 = ~n50901;
  assign po831 = ~n50950;
  assign po832 = ~n50999;
  assign po833 = ~n51041;
  assign po834 = ~n52080;
  assign po835 = ~n52116;
  assign po836 = ~n51084;
  assign po839 = ~n52152;
  assign po840 = ~n38261;
  assign po842 = ~n51136;
  assign po846 = ~n51180;
  assign po849 = ~n51229;
  assign po864 = ~n65222;
  assign po868 = ~n65230;
  assign po869 = ~n51423;
  assign po870 = ~n65239;
  assign po871 = ~n51518;
  assign po874 = ~n51611;
  assign po876 = ~n51703;
  assign po877 = ~n51750;
  assign po878 = ~n61725;
  assign po879 = ~n51797;
  assign po896 = ~n65883;
  assign po898 = ~n65884;
  assign po899 = ~n65885;
  assign po900 = ~n65886;
  assign po901 = ~n65887;
  assign po902 = ~n65888;
  assign po903 = ~n65889;
  assign po905 = ~n65890;
  assign po906 = ~n65891;
  assign po907 = ~n65892;
  assign po908 = ~n65893;
  assign po909 = ~n65894;
  assign po910 = ~n65934;
  assign po911 = ~n65935;
  assign po912 = ~n65936;
  assign po913 = ~n65937;
  assign po914 = ~n65938;
  assign po915 = ~n65939;
  assign po916 = ~n65940;
  assign po917 = ~n65941;
  assign po918 = ~n65942;
  assign po919 = ~n65943;
  assign po920 = ~n65944;
  assign po921 = ~n65945;
  assign po923 = ~n65946;
  assign po924 = ~n65947;
  assign po925 = ~n65948;
  assign po926 = ~n61785;
  assign po927 = ~n65949;
  assign po928 = ~n61809;
  assign po929 = ~n65950;
  assign po931 = ~n65951;
  assign po933 = ~n65952;
  assign po934 = ~n65953;
  assign po935 = ~n61867;
  assign po936 = ~n61392;
  assign po937 = ~n61393;
  assign po938 = ~n61870;
  assign po939 = ~n61167;
  assign po940 = ~n61873;
  assign po941 = ~n61876;
  assign po942 = ~n61879;
  assign po943 = ~n65079;
  assign po944 = ~n61882;
  assign po945 = ~n61885;
  assign po946 = ~n61888;
  assign po947 = ~n61891;
  assign po948 = ~n61894;
  assign po949 = ~n61897;
  assign po950 = ~n40220;
  assign po951 = ~n61901;
  assign po952 = ~n61904;
  assign po955 = ~n61907;
  assign po957 = ~n61913;
  assign po958 = ~n61916;
  assign po961 = ~n61922;
  assign po964 = ~n61925;
  assign po965 = ~n61928;
  assign po967 = ~n61934;
  assign po968 = ~n61937;
  assign po970 = ~n61943;
  assign po972 = ~n61949;
  assign po973 = ~n61952;
  assign po975 = ~n48952;
  assign po990 = ~n48967;
  assign po996 = ~n62302;
  assign po1002 = ~n62236;
  assign po1005 = ~n62305;
  assign po1017 = ~n62246;
  assign po1018 = ~n62249;
  assign po1019 = ~n62308;
  assign po1020 = ~n62311;
  assign po1025 = ~n62259;
  assign po1033 = ~n62279;
  assign po1034 = ~n62289;
  assign po1035 = ~n62299;
  assign po1038 = ~n62455;
  assign po1039 = ~n62147;
  assign po1040 = ~n62150;
  assign po1041 = ~n62153;
  assign po1042 = ~n62156;
  assign po1043 = ~n62158;
  assign po1044 = ~n62161;
  assign po1045 = ~n62164;
  assign po1046 = ~n62167;
  assign po1047 = ~n62170;
  assign po1048 = ~n62173;
  assign po1049 = ~n30695;
  assign po1050 = ~n62176;
  assign po1051 = ~n62179;
  assign po1052 = ~n62182;
  assign po1053 = pi67;
  assign po1054 = ~n62185;
  assign po1055 = ~n62187;
  assign po1056 = ~n62190;
  assign po1057 = ~n2843;
  assign po1058 = ~n62193;
  assign po1059 = ~n62196;
  assign po1060 = ~n62198;
  assign po1061 = ~n62200;
  assign po1062 = ~n62203;
  assign po1064 = ~n62205;
  assign po1065 = ~n62208;
  assign po1066 = ~n62211;
  assign po1067 = ~n62214;
  assign po1068 = ~n62216;
  assign po1069 = ~n62219;
  assign po1071 = ~n62222;
  assign po1072 = ~n62224;
  assign po1073 = ~n62227;
  assign po1074 = ~n62230;
  assign po1075 = ~n62233;
  assign po1077 = ~n48983;
  assign po1078 = ~n66041;
  assign po1079 = ~n65957;
  assign po1081 = ~n65958;
  assign po1082 = ~n65959;
  assign po1083 = ~n65081;
  assign po1085 = ~n65082;
  assign po1086 = ~n65083;
  assign po1087 = ~n65960;
  assign po1088 = ~n49007;
  assign po1089 = ~n49010;
  assign po1090 = ~n65961;
  assign po1091 = ~n49013;
  assign po1092 = ~n65962;
  assign po1093 = ~n65963;
  assign po1094 = ~n49016;
  assign po1095 = ~n65084;
  assign po1096 = ~n49025;
  assign po1097 = ~n65964;
  assign po1098 = ~n65965;
  assign po1099 = ~n65966;
  assign po1101 = ~n2908;
  assign po1103 = ~n61414;
  assign po1108 = pi1134;
  assign po1109 = pi964;
  assign po1110 = ~pi954;
  assign po1111 = pi965;
  assign po1112 = ~n49033;
  assign po1113 = pi991;
  assign po1114 = pi985;
  assign po1117 = pi1014;
  assign po1119 = pi1029;
  assign po1120 = pi1004;
  assign po1121 = pi1007;
  assign po1123 = pi1135;
  assign po1130 = ~pi278;
  assign po1133 = ~n61475;
  assign po1134 = pi1064;
  assign po1136 = pi299;
  assign po1137 = ~n61476;
  assign po1138 = pi1075;
  assign po1139 = pi1052;
  assign po1140 = pi771;
  assign po1141 = pi765;
  assign po1142 = pi605;
  assign po1143 = pi601;
  assign po1144 = pi278;
  assign po1145 = pi279;
  assign po1146 = ~pi915;
  assign po1147 = ~pi825;
  assign po1148 = ~pi826;
  assign po1149 = ~pi913;
  assign po1150 = ~pi894;
  assign po1151 = ~pi905;
  assign po1152 = pi1095;
  assign po1153 = ~pi890;
  assign po1154 = pi1094;
  assign po1155 = ~pi906;
  assign po1156 = ~pi896;
  assign po1157 = ~pi909;
  assign po1158 = ~pi911;
  assign po1159 = ~pi908;
  assign po1160 = ~pi891;
  assign po1161 = ~pi902;
  assign po1162 = ~pi903;
  assign po1163 = ~pi883;
  assign po1164 = ~pi888;
  assign po1165 = ~pi919;
  assign po1166 = ~pi886;
  assign po1167 = ~pi912;
  assign po1168 = ~pi895;
  assign po1169 = ~pi916;
  assign po1170 = ~pi889;
  assign po1171 = ~pi900;
  assign po1172 = ~pi885;
  assign po1173 = ~pi904;
  assign po1174 = ~pi899;
  assign po1175 = ~pi918;
  assign po1176 = ~pi898;
  assign po1177 = ~pi917;
  assign po1178 = ~pi827;
  assign po1179 = ~pi887;
  assign po1180 = ~pi884;
  assign po1181 = ~pi910;
  assign po1182 = ~pi828;
  assign po1183 = ~pi892;
  assign po1184 = pi1187;
  assign po1185 = pi1172;
  assign po1186 = pi1170;
  assign po1187 = pi1138;
  assign po1188 = pi1177;
  assign po1189 = pi1178;
  assign po1190 = pi863;
  assign po1191 = pi1203;
  assign po1192 = pi1185;
  assign po1193 = pi1171;
  assign po1194 = pi1192;
  assign po1195 = pi1137;
  assign po1196 = pi1186;
  assign po1197 = pi1165;
  assign po1198 = pi1164;
  assign po1199 = pi1098;
  assign po1200 = pi1183;
  assign po1201 = pi230;
  assign po1202 = pi1169;
  assign po1203 = pi1136;
  assign po1204 = pi1181;
  assign po1205 = pi849;
  assign po1206 = pi1193;
  assign po1207 = pi1182;
  assign po1208 = pi1168;
  assign po1209 = pi1175;
  assign po1210 = pi1191;
  assign po1211 = pi1099;
  assign po1212 = pi1174;
  assign po1213 = pi1179;
  assign po1214 = pi1202;
  assign po1215 = pi1176;
  assign po1216 = pi1173;
  assign po1217 = pi1201;
  assign po1218 = pi1167;
  assign po1219 = pi840;
  assign po1220 = pi1189;
  assign po1221 = pi1195;
  assign po1222 = pi864;
  assign po1223 = pi1190;
  assign po1224 = pi1188;
  assign po1225 = pi1180;
  assign po1226 = pi1194;
  assign po1227 = pi1097;
  assign po1228 = pi1166;
  assign po1229 = pi1200;
  assign po1230 = pi1184;
endmodule
