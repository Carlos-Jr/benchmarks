module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n493, n495, n496,
    n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n659,
    n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687,
    n688, n689, n690, n692, n693, n694, n695,
    n696, n697;
  assign n23 = pi08 & pi10;
  assign n24 = ~pi09 & pi11;
  assign n25 = ~pi13 & n24;
  assign n26 = n23 & n25;
  assign n27 = pi10 & ~pi11;
  assign n28 = ~pi08 & pi09;
  assign n29 = pi13 & n28;
  assign n30 = ~n27 & n29;
  assign n31 = pi08 & pi09;
  assign n32 = n27 & n31;
  assign n33 = ~n26 & ~n32;
  assign n34 = ~n30 & n33;
  assign n35 = ~pi04 & ~n34;
  assign n36 = ~pi08 & ~pi09;
  assign n37 = ~n31 & ~n36;
  assign n38 = ~pi10 & pi11;
  assign n39 = ~n37 & n38;
  assign n40 = pi13 & n39;
  assign n41 = ~pi09 & ~pi11;
  assign n42 = ~pi08 & pi10;
  assign n43 = n41 & n42;
  assign n44 = ~n40 & ~n43;
  assign n45 = pi00 & pi04;
  assign n46 = ~n44 & n45;
  assign n47 = ~pi00 & ~pi04;
  assign n48 = pi08 & ~pi09;
  assign n49 = pi10 & pi13;
  assign n50 = ~pi10 & ~pi11;
  assign n51 = ~pi13 & n50;
  assign n52 = ~n49 & ~n51;
  assign n53 = n48 & ~n52;
  assign n54 = ~n47 & n53;
  assign n55 = pi00 & ~pi04;
  assign n56 = ~pi00 & pi04;
  assign n57 = n27 & n56;
  assign n58 = ~n55 & ~n57;
  assign n59 = n29 & ~n58;
  assign n60 = pi09 & pi11;
  assign n61 = ~pi10 & ~pi13;
  assign n62 = ~n60 & n61;
  assign n63 = ~pi08 & n62;
  assign n64 = ~pi00 & n63;
  assign n65 = ~n59 & ~n64;
  assign n66 = ~n54 & n65;
  assign n67 = ~n35 & n66;
  assign n68 = ~n46 & n67;
  assign n69 = pi00 & pi11;
  assign n70 = ~n31 & n69;
  assign n71 = pi11 & n29;
  assign n72 = ~pi10 & n71;
  assign n73 = n45 & n72;
  assign n74 = ~pi00 & n68;
  assign n75 = n71 & ~n74;
  assign n76 = pi13 & n27;
  assign n77 = pi00 & ~n68;
  assign n78 = n31 & n77;
  assign n79 = n36 & n68;
  assign n80 = n45 & n48;
  assign n81 = ~n79 & ~n80;
  assign n82 = ~n78 & n81;
  assign n83 = n76 & ~n82;
  assign n84 = ~n75 & ~n83;
  assign n85 = ~pi09 & n27;
  assign n86 = pi13 & n85;
  assign n87 = pi08 & n86;
  assign n88 = n84 & n87;
  assign n89 = ~n73 & ~n88;
  assign n90 = pi08 & n41;
  assign n91 = ~n89 & n90;
  assign n92 = ~n70 & ~n91;
  assign n93 = pi10 & ~n92;
  assign n94 = ~pi10 & n31;
  assign n95 = n27 & n28;
  assign n96 = ~n94 & ~n95;
  assign n97 = ~n50 & ~n96;
  assign n98 = ~n93 & ~n97;
  assign n99 = n68 & ~n98;
  assign n100 = ~pi00 & ~pi08;
  assign n101 = n85 & n100;
  assign n102 = ~pi08 & ~pi10;
  assign n103 = pi09 & n102;
  assign n104 = pi11 & n103;
  assign n105 = n89 & n104;
  assign n106 = ~n101 & ~n105;
  assign n107 = ~n84 & ~n106;
  assign n108 = pi08 & ~pi10;
  assign n109 = pi04 & n108;
  assign n110 = pi00 & ~pi08;
  assign n111 = n84 & n110;
  assign n112 = ~n109 & ~n111;
  assign n113 = n41 & ~n112;
  assign n114 = pi09 & ~n68;
  assign n115 = ~pi00 & ~n114;
  assign n116 = ~pi11 & ~n115;
  assign n117 = pi00 & ~pi09;
  assign n118 = n68 & n117;
  assign n119 = ~n116 & ~n118;
  assign n120 = n102 & ~n119;
  assign n121 = ~pi09 & n108;
  assign n122 = ~n45 & ~n47;
  assign n123 = n121 & n122;
  assign n124 = ~pi00 & pi11;
  assign n125 = pi09 & n23;
  assign n126 = n124 & n125;
  assign n127 = pi08 & n85;
  assign n128 = n89 & n127;
  assign n129 = ~pi10 & ~n36;
  assign n130 = n124 & ~n129;
  assign n131 = ~n128 & ~n130;
  assign n132 = ~n68 & ~n131;
  assign n133 = ~n89 & n104;
  assign n134 = ~n32 & ~n133;
  assign n135 = n84 & ~n134;
  assign n136 = ~n123 & ~n126;
  assign n137 = ~n120 & n136;
  assign n138 = ~n113 & n137;
  assign n139 = ~n107 & n138;
  assign n140 = ~n132 & ~n135;
  assign n141 = n139 & n140;
  assign n142 = ~n99 & n141;
  assign n143 = pi13 & ~n142;
  assign n144 = pi12 & n143;
  assign n145 = ~pi12 & ~n143;
  assign n146 = ~n144 & ~n145;
  assign n147 = pi13 & ~n146;
  assign n148 = pi13 & n31;
  assign n149 = n50 & n148;
  assign n150 = n25 & n42;
  assign n151 = ~n149 & ~n150;
  assign n152 = n23 & n77;
  assign n153 = ~pi11 & ~n42;
  assign n154 = n45 & ~n153;
  assign n155 = ~pi08 & n27;
  assign n156 = n47 & n155;
  assign n157 = ~pi08 & pi11;
  assign n158 = pi04 & n157;
  assign n159 = ~n154 & ~n158;
  assign n160 = ~n156 & n159;
  assign n161 = ~n152 & n160;
  assign n162 = pi09 & ~n161;
  assign n163 = pi08 & n50;
  assign n164 = ~n42 & ~n163;
  assign n165 = n68 & ~n164;
  assign n166 = pi11 & n108;
  assign n167 = n56 & n166;
  assign n168 = pi08 & n27;
  assign n169 = ~pi04 & n168;
  assign n170 = pi11 & n55;
  assign n171 = ~n167 & ~n170;
  assign n172 = ~n169 & n171;
  assign n173 = ~n165 & n172;
  assign n174 = ~pi09 & ~n173;
  assign n175 = pi04 & n102;
  assign n176 = ~n31 & ~n129;
  assign n177 = ~n27 & n176;
  assign n178 = ~pi09 & n177;
  assign n179 = ~n175 & ~n178;
  assign n180 = ~n68 & ~n179;
  assign n181 = n69 & ~n129;
  assign n182 = ~n180 & ~n181;
  assign n183 = ~n174 & n182;
  assign n184 = ~n162 & n183;
  assign n185 = ~pi13 & ~n184;
  assign n186 = n151 & ~n185;
  assign po0 = n147 | ~n186;
  assign n188 = ~pi12 & n143;
  assign n189 = ~pi08 & pi13;
  assign n190 = ~pi09 & pi10;
  assign n191 = n69 & n190;
  assign n192 = pi01 & ~pi05;
  assign n193 = ~pi01 & pi05;
  assign n194 = n27 & n193;
  assign n195 = ~n192 & ~n194;
  assign n196 = ~n56 & ~n195;
  assign n197 = ~pi01 & ~pi05;
  assign n198 = n56 & n197;
  assign n199 = ~n196 & ~n198;
  assign n200 = pi09 & ~n199;
  assign n201 = ~n191 & ~n200;
  assign n202 = n189 & ~n201;
  assign n203 = pi01 & pi05;
  assign n204 = n44 & ~n86;
  assign n205 = n57 & n189;
  assign n206 = n204 & ~n205;
  assign n207 = n203 & ~n206;
  assign n208 = ~pi05 & ~n34;
  assign n209 = n53 & ~n197;
  assign n210 = ~pi01 & n63;
  assign n211 = ~n209 & ~n210;
  assign n212 = ~n208 & n211;
  assign n213 = ~n202 & n212;
  assign n214 = ~n207 & n213;
  assign n215 = ~n68 & ~n89;
  assign n216 = n72 & n203;
  assign n217 = ~pi01 & n214;
  assign n218 = n71 & ~n217;
  assign n219 = n36 & n214;
  assign n220 = pi09 & ~n214;
  assign n221 = pi05 & ~pi09;
  assign n222 = ~n220 & ~n221;
  assign n223 = pi01 & pi08;
  assign n224 = ~n222 & n223;
  assign n225 = ~n219 & ~n224;
  assign n226 = n76 & ~n225;
  assign n227 = ~n218 & ~n226;
  assign n228 = n87 & n227;
  assign n229 = ~n216 & ~n228;
  assign n230 = n215 & ~n229;
  assign n231 = ~n215 & n229;
  assign n232 = ~n230 & ~n231;
  assign n233 = ~n214 & ~n232;
  assign n234 = n214 & n232;
  assign n235 = ~n233 & ~n234;
  assign n236 = n23 & ~n235;
  assign n237 = pi05 & n108;
  assign n238 = pi00 & ~n84;
  assign n239 = n227 & n238;
  assign n240 = ~n227 & ~n238;
  assign n241 = ~n239 & ~n240;
  assign n242 = pi01 & ~pi08;
  assign n243 = n241 & n242;
  assign n244 = ~n237 & ~n243;
  assign n245 = ~n236 & n244;
  assign n246 = n41 & ~n245;
  assign n247 = ~n84 & ~n89;
  assign n248 = ~n229 & n247;
  assign n249 = n229 & ~n247;
  assign n250 = ~n248 & ~n249;
  assign n251 = ~n227 & ~n250;
  assign n252 = n227 & n250;
  assign n253 = ~n251 & ~n252;
  assign n254 = n104 & ~n253;
  assign n255 = n84 & n227;
  assign n256 = ~n84 & ~n227;
  assign n257 = ~n255 & ~n256;
  assign n258 = n125 & ~n257;
  assign n259 = n103 & ~n214;
  assign n260 = ~n258 & ~n259;
  assign n261 = ~pi11 & ~n260;
  assign n262 = pi11 & n176;
  assign n263 = n77 & ~n214;
  assign n264 = ~n77 & n214;
  assign n265 = ~n263 & ~n264;
  assign n266 = n262 & n265;
  assign n267 = n43 & ~n241;
  assign n268 = ~n266 & ~n267;
  assign n269 = ~pi01 & ~n268;
  assign n270 = n177 & ~n265;
  assign n271 = ~pi05 & ~n45;
  assign n272 = n121 & n271;
  assign n273 = n69 & n125;
  assign n274 = ~n31 & n50;
  assign n275 = ~n272 & ~n274;
  assign n276 = ~n273 & n275;
  assign n277 = ~n270 & n276;
  assign n278 = pi01 & ~n277;
  assign n279 = n68 & n214;
  assign n280 = n97 & n279;
  assign n281 = ~pi11 & n103;
  assign n282 = ~n97 & ~n281;
  assign n283 = ~n68 & ~n282;
  assign n284 = ~n214 & n283;
  assign n285 = ~pi00 & ~pi01;
  assign n286 = n125 & n285;
  assign n287 = n45 & n197;
  assign n288 = n121 & n287;
  assign n289 = ~n286 & ~n288;
  assign n290 = pi11 & ~n289;
  assign n291 = ~n45 & n193;
  assign n292 = n45 & n203;
  assign n293 = ~n291 & ~n292;
  assign n294 = n121 & ~n293;
  assign n295 = ~n290 & ~n294;
  assign n296 = ~n284 & n295;
  assign n297 = ~n280 & n296;
  assign n298 = ~n278 & n297;
  assign n299 = ~n261 & n298;
  assign n300 = ~n269 & n299;
  assign n301 = ~n254 & n300;
  assign n302 = ~n246 & n301;
  assign n303 = pi13 & ~n302;
  assign n304 = ~n188 & n303;
  assign n305 = n188 & ~n303;
  assign n306 = ~n304 & ~n305;
  assign n307 = pi13 & ~n306;
  assign n308 = ~n164 & n214;
  assign n309 = ~pi05 & n168;
  assign n310 = n166 & n193;
  assign n311 = pi11 & n192;
  assign n312 = ~n309 & ~n311;
  assign n313 = ~n310 & n312;
  assign n314 = ~n308 & n313;
  assign n315 = ~pi09 & ~n314;
  assign n316 = pi11 & ~n129;
  assign n317 = n125 & ~n214;
  assign n318 = ~n316 & ~n317;
  assign n319 = pi01 & ~n318;
  assign n320 = pi05 & n102;
  assign n321 = ~n178 & ~n320;
  assign n322 = ~n214 & ~n321;
  assign n323 = n155 & n197;
  assign n324 = ~n153 & n203;
  assign n325 = pi05 & n157;
  assign n326 = ~n323 & ~n325;
  assign n327 = ~n324 & n326;
  assign n328 = pi09 & ~n327;
  assign n329 = ~n322 & ~n328;
  assign n330 = ~n315 & n329;
  assign n331 = ~n319 & n330;
  assign n332 = ~pi13 & ~n331;
  assign n333 = n151 & ~n332;
  assign po1 = n307 | ~n333;
  assign n335 = n188 & n303;
  assign n336 = n56 & ~n192;
  assign n337 = ~n193 & ~n336;
  assign n338 = ~pi06 & ~n337;
  assign n339 = pi06 & n27;
  assign n340 = n337 & n339;
  assign n341 = ~n338 & ~n340;
  assign n342 = ~pi02 & pi09;
  assign n343 = ~n341 & n342;
  assign n344 = ~n337 & n339;
  assign n345 = ~pi06 & pi09;
  assign n346 = n337 & n345;
  assign n347 = ~n344 & ~n346;
  assign n348 = pi02 & ~n347;
  assign n349 = pi01 & pi11;
  assign n350 = n190 & n349;
  assign n351 = ~n343 & ~n350;
  assign n352 = ~n348 & n351;
  assign n353 = n189 & ~n352;
  assign n354 = pi02 & pi06;
  assign n355 = ~n204 & n354;
  assign n356 = ~pi06 & ~n34;
  assign n357 = ~pi02 & n63;
  assign n358 = ~pi02 & ~pi06;
  assign n359 = n53 & ~n358;
  assign n360 = ~n357 & ~n359;
  assign n361 = ~n356 & n360;
  assign n362 = ~n355 & n361;
  assign n363 = ~n353 & n362;
  assign n364 = n72 & n354;
  assign n365 = ~pi02 & n363;
  assign n366 = n71 & ~n365;
  assign n367 = n36 & n363;
  assign n368 = pi09 & ~n363;
  assign n369 = pi06 & ~pi09;
  assign n370 = ~n368 & ~n369;
  assign n371 = pi02 & pi08;
  assign n372 = ~n370 & n371;
  assign n373 = ~n367 & ~n372;
  assign n374 = n76 & ~n373;
  assign n375 = ~n366 & ~n374;
  assign n376 = n87 & n375;
  assign n377 = ~n364 & ~n376;
  assign n378 = n363 & n377;
  assign n379 = ~n363 & ~n377;
  assign n380 = ~n378 & ~n379;
  assign n381 = ~n231 & ~n234;
  assign n382 = ~n380 & n381;
  assign n383 = n380 & ~n381;
  assign n384 = ~n382 & ~n383;
  assign n385 = n23 & ~n384;
  assign n386 = pi06 & n108;
  assign n387 = ~pi01 & ~n238;
  assign n388 = ~n227 & ~n387;
  assign n389 = pi01 & n238;
  assign n390 = ~n388 & ~n389;
  assign n391 = ~n375 & n390;
  assign n392 = n375 & ~n390;
  assign n393 = ~n391 & ~n392;
  assign n394 = pi02 & ~pi08;
  assign n395 = n393 & n394;
  assign n396 = ~n386 & ~n395;
  assign n397 = ~n385 & n396;
  assign n398 = n41 & ~n397;
  assign n399 = ~n227 & ~n249;
  assign n400 = ~n248 & ~n399;
  assign n401 = ~n375 & n400;
  assign n402 = n375 & ~n400;
  assign n403 = ~n401 & ~n402;
  assign n404 = ~n377 & n403;
  assign n405 = n377 & ~n403;
  assign n406 = ~n404 & ~n405;
  assign n407 = n104 & ~n406;
  assign n408 = ~pi01 & ~n77;
  assign n409 = ~n214 & ~n408;
  assign n410 = pi01 & n77;
  assign n411 = ~n409 & ~n410;
  assign n412 = n262 & ~n363;
  assign n413 = n411 & n412;
  assign n414 = n43 & ~n393;
  assign n415 = ~n413 & ~n414;
  assign n416 = ~pi02 & ~n415;
  assign n417 = n255 & n375;
  assign n418 = ~n255 & ~n375;
  assign n419 = ~n417 & ~n418;
  assign n420 = ~pi11 & ~n419;
  assign n421 = ~pi02 & n285;
  assign n422 = pi11 & n421;
  assign n423 = pi02 & pi11;
  assign n424 = ~n285 & n423;
  assign n425 = ~n422 & ~n424;
  assign n426 = ~n420 & n425;
  assign n427 = n125 & ~n426;
  assign n428 = n177 & ~n363;
  assign n429 = ~n411 & n428;
  assign n430 = ~n274 & ~n429;
  assign n431 = pi02 & ~n430;
  assign n432 = pi02 & n177;
  assign n433 = n411 & n432;
  assign n434 = ~pi02 & n262;
  assign n435 = ~n411 & n434;
  assign n436 = ~n433 & ~n435;
  assign n437 = n363 & ~n436;
  assign n438 = ~n279 & ~n282;
  assign n439 = ~n281 & ~n438;
  assign n440 = ~n363 & ~n439;
  assign n441 = n45 & ~n197;
  assign n442 = ~n203 & ~n441;
  assign n443 = pi11 & n358;
  assign n444 = ~n354 & ~n443;
  assign n445 = ~n442 & ~n444;
  assign n446 = ~n354 & ~n358;
  assign n447 = n442 & n446;
  assign n448 = ~n445 & ~n447;
  assign n449 = n121 & ~n448;
  assign n450 = n279 & n363;
  assign n451 = n97 & n450;
  assign n452 = ~n449 & ~n451;
  assign n453 = ~n440 & n452;
  assign n454 = ~n431 & n453;
  assign n455 = ~n437 & n454;
  assign n456 = ~n427 & n455;
  assign n457 = ~n416 & n456;
  assign n458 = ~n407 & n457;
  assign n459 = ~n398 & n458;
  assign n460 = pi13 & ~n459;
  assign n461 = ~n335 & n460;
  assign n462 = n335 & ~n460;
  assign n463 = ~n461 & ~n462;
  assign n464 = pi13 & ~n463;
  assign n465 = ~n164 & n363;
  assign n466 = ~pi06 & n168;
  assign n467 = ~n465 & ~n466;
  assign n468 = ~pi09 & ~n467;
  assign n469 = pi06 & n102;
  assign n470 = pi02 & n125;
  assign n471 = ~n469 & ~n470;
  assign n472 = ~n178 & n471;
  assign n473 = ~n363 & ~n472;
  assign n474 = ~n153 & n354;
  assign n475 = n155 & n358;
  assign n476 = ~n474 & ~n475;
  assign n477 = pi09 & ~n476;
  assign n478 = pi09 & n157;
  assign n479 = ~pi02 & ~pi09;
  assign n480 = n166 & n479;
  assign n481 = ~n478 & ~n480;
  assign n482 = pi06 & ~n481;
  assign n483 = ~pi06 & ~pi09;
  assign n484 = n129 & ~n483;
  assign n485 = n423 & ~n484;
  assign n486 = ~n477 & ~n485;
  assign n487 = ~n482 & n486;
  assign n488 = ~n473 & n487;
  assign n489 = ~n468 & n488;
  assign n490 = ~pi13 & ~n489;
  assign n491 = n151 & ~n490;
  assign po2 = n464 | ~n491;
  assign n493 = n335 & n460;
  assign po5 = pi03 & pi07;
  assign n495 = n72 & po5;
  assign n496 = pi02 & ~pi06;
  assign n497 = ~pi02 & pi06;
  assign n498 = n337 & ~n497;
  assign n499 = ~n496 & ~n498;
  assign n500 = n76 & n499;
  assign n501 = ~n85 & ~n500;
  assign n502 = po5 & ~n501;
  assign n503 = pi07 & pi09;
  assign n504 = n76 & n503;
  assign n505 = ~n499 & n504;
  assign n506 = ~n62 & ~n505;
  assign n507 = ~pi03 & ~n506;
  assign n508 = n190 & n423;
  assign n509 = ~pi03 & ~pi07;
  assign n510 = pi09 & n509;
  assign n511 = n499 & n510;
  assign n512 = ~n508 & ~n511;
  assign n513 = pi13 & ~n512;
  assign n514 = ~n502 & ~n507;
  assign n515 = ~n513 & n514;
  assign n516 = ~pi08 & ~n515;
  assign n517 = pi03 & n29;
  assign n518 = ~n499 & n517;
  assign n519 = n34 & ~n518;
  assign n520 = ~pi07 & ~n519;
  assign n521 = ~n39 & ~n85;
  assign n522 = pi13 & po5;
  assign n523 = ~n521 & n522;
  assign n524 = n53 & ~n509;
  assign n525 = ~n523 & ~n524;
  assign n526 = ~n520 & n525;
  assign n527 = ~n516 & n526;
  assign n528 = ~pi03 & n527;
  assign n529 = n71 & ~n528;
  assign n530 = pi03 & ~n527;
  assign n531 = n31 & n530;
  assign n532 = n36 & n527;
  assign n533 = n48 & po5;
  assign n534 = ~n532 & ~n533;
  assign n535 = ~n531 & n534;
  assign n536 = n76 & ~n535;
  assign n537 = ~n529 & ~n536;
  assign n538 = n87 & n537;
  assign n539 = ~n495 & ~n538;
  assign n540 = n377 & n400;
  assign n541 = ~n375 & ~n540;
  assign n542 = ~n377 & ~n400;
  assign n543 = ~n541 & ~n542;
  assign n544 = ~n537 & n543;
  assign n545 = n537 & ~n543;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~n539 & n546;
  assign n548 = n539 & ~n546;
  assign n549 = ~n547 & ~n548;
  assign n550 = n103 & ~n549;
  assign n551 = ~pi03 & n125;
  assign n552 = n421 & n551;
  assign n553 = ~n358 & ~n447;
  assign n554 = n121 & n509;
  assign n555 = n553 & n554;
  assign n556 = ~n552 & ~n555;
  assign n557 = ~n550 & n556;
  assign n558 = pi11 & ~n557;
  assign n559 = ~pi02 & n390;
  assign n560 = ~n375 & ~n559;
  assign n561 = pi02 & ~n390;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~n537 & ~n562;
  assign n564 = n537 & n562;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~pi03 & ~pi08;
  assign n567 = n565 & n566;
  assign n568 = ~n527 & n539;
  assign n569 = n527 & ~n539;
  assign n570 = ~n568 & ~n569;
  assign n571 = ~n377 & n381;
  assign n572 = ~n363 & ~n383;
  assign n573 = ~n571 & ~n572;
  assign n574 = n570 & ~n573;
  assign n575 = ~n570 & n573;
  assign n576 = ~n574 & ~n575;
  assign n577 = pi08 & ~n576;
  assign n578 = ~n567 & ~n577;
  assign n579 = n85 & ~n578;
  assign n580 = pi03 & n36;
  assign n581 = ~n565 & n580;
  assign n582 = pi07 & n121;
  assign n583 = n417 & n537;
  assign n584 = ~n417 & ~n537;
  assign n585 = ~n583 & ~n584;
  assign n586 = n125 & ~n585;
  assign n587 = ~n582 & ~n586;
  assign n588 = ~n581 & n587;
  assign n589 = ~pi11 & ~n588;
  assign n590 = ~pi02 & n411;
  assign n591 = ~n363 & ~n590;
  assign n592 = pi02 & ~n411;
  assign n593 = ~n591 & ~n592;
  assign n594 = ~n527 & n593;
  assign n595 = n527 & ~n593;
  assign n596 = ~n594 & ~n595;
  assign n597 = n177 & n596;
  assign n598 = ~n274 & ~n597;
  assign n599 = pi03 & ~n598;
  assign n600 = n262 & ~n596;
  assign n601 = ~n553 & n582;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~pi03 & ~n602;
  assign n604 = ~n282 & ~n450;
  assign n605 = ~n281 & ~n604;
  assign n606 = ~n527 & ~n605;
  assign n607 = n450 & n527;
  assign n608 = n97 & n607;
  assign n609 = po5 & n553;
  assign n610 = ~n509 & n553;
  assign n611 = ~po5 & ~n610;
  assign n612 = pi03 & n611;
  assign n613 = ~n609 & ~n612;
  assign n614 = n121 & ~n613;
  assign n615 = pi03 & pi11;
  assign n616 = n125 & n615;
  assign n617 = ~n421 & n616;
  assign n618 = ~n614 & ~n617;
  assign n619 = ~n608 & n618;
  assign n620 = ~n606 & n619;
  assign n621 = ~n599 & n620;
  assign n622 = ~n603 & n621;
  assign n623 = ~n589 & n622;
  assign n624 = ~n579 & n623;
  assign n625 = ~n558 & n624;
  assign n626 = pi13 & ~n625;
  assign n627 = ~n493 & n626;
  assign n628 = n493 & ~n626;
  assign n629 = ~n627 & ~n628;
  assign n630 = pi13 & ~n629;
  assign n631 = n23 & n530;
  assign n632 = n155 & n509;
  assign n633 = ~n153 & po5;
  assign n634 = ~n632 & ~n633;
  assign n635 = ~n631 & n634;
  assign n636 = pi09 & ~n635;
  assign n637 = ~n164 & n527;
  assign n638 = ~pi07 & n168;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~pi09 & ~n639;
  assign n641 = pi07 & n102;
  assign n642 = ~n178 & ~n641;
  assign n643 = ~n527 & ~n642;
  assign n644 = ~pi07 & ~pi09;
  assign n645 = n129 & ~n644;
  assign n646 = n615 & ~n645;
  assign n647 = ~pi03 & ~pi09;
  assign n648 = n166 & n647;
  assign n649 = ~n478 & ~n648;
  assign n650 = pi07 & ~n649;
  assign n651 = ~n646 & ~n650;
  assign n652 = ~n643 & n651;
  assign n653 = ~n640 & n652;
  assign n654 = ~n636 & n653;
  assign n655 = ~pi13 & ~n654;
  assign n656 = n151 & ~n655;
  assign po3 = n630 | ~n656;
  assign po4 = po5 | n509;
  assign n659 = n493 & n626;
  assign n660 = ~pi03 & n562;
  assign n661 = ~n537 & ~n660;
  assign n662 = pi03 & ~n562;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~pi08 & ~n663;
  assign n665 = ~n527 & ~n573;
  assign n666 = ~n539 & ~n575;
  assign n667 = ~n665 & ~n666;
  assign n668 = pi08 & ~n667;
  assign n669 = ~n664 & ~n668;
  assign n670 = n190 & ~n669;
  assign n671 = n31 & n583;
  assign n672 = ~n94 & ~n671;
  assign n673 = ~n670 & n672;
  assign n674 = ~pi11 & ~n673;
  assign n675 = ~n96 & n607;
  assign n676 = ~n539 & ~n543;
  assign n677 = ~n537 & ~n548;
  assign n678 = ~n676 & ~n677;
  assign n679 = n103 & ~n678;
  assign n680 = ~n528 & ~n593;
  assign n681 = ~n530 & ~n680;
  assign n682 = n176 & ~n681;
  assign n683 = n121 & ~n611;
  assign n684 = ~n552 & ~n683;
  assign n685 = ~n682 & n684;
  assign n686 = ~n679 & n685;
  assign n687 = pi11 & ~n686;
  assign n688 = ~n675 & ~n687;
  assign n689 = ~n674 & n688;
  assign n690 = ~n659 & n689;
  assign po6 = pi13 & ~n690;
  assign n692 = n285 & ~n446;
  assign n693 = n337 & n692;
  assign n694 = ~n122 & n203;
  assign n695 = ~n287 & ~n694;
  assign n696 = ~n446 & ~n695;
  assign n697 = ~n693 & ~n696;
  assign po7 = po4 & ~n697;
endmodule
