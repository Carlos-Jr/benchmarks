module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7;
  wire n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n754, n755,
    n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798,
    n800, n801, n802, n803, n806, n807, n808,
    n809, n810, n811;
  assign n137 = pi118  & ~pi119 ;
  assign n138 = ~pi120  & ~n137;
  assign n139 = ~pi121  & ~n138;
  assign n140 = ~pi122  & ~n139;
  assign n141 = ~pi123  & ~n140;
  assign n142 = ~pi124  & ~n141;
  assign n143 = ~pi125  & ~n142;
  assign n144 = ~pi126  & ~n143;
  assign n145 = pi117  & n144;
  assign n146 = pi119  & ~pi120 ;
  assign n147 = ~pi121  & ~n146;
  assign n148 = ~pi122  & ~n147;
  assign n149 = ~pi123  & ~n148;
  assign n150 = ~pi124  & ~n149;
  assign n151 = ~pi125  & ~n150;
  assign n152 = ~pi117  & ~pi126 ;
  assign n153 = ~n151 & n152;
  assign n154 = ~pi127  & ~n153;
  assign n155 = ~n145 & n154;
  assign n156 = ~pi115  & ~n155;
  assign n157 = ~pi127  & ~n144;
  assign n158 = ~pi116  & ~n157;
  assign n159 = pi116  & ~n155;
  assign n160 = ~n158 & ~n159;
  assign n161 = pi115  & ~n160;
  assign n162 = ~n156 & ~n161;
  assign n163 = ~pi113  & ~n162;
  assign n164 = ~pi114  & ~n160;
  assign n165 = pi114  & ~n162;
  assign n166 = ~n164 & ~n165;
  assign n167 = pi113  & ~n166;
  assign n168 = ~n163 & ~n167;
  assign n169 = ~pi111  & ~n168;
  assign n170 = ~pi112  & ~n166;
  assign n171 = pi112  & ~n168;
  assign n172 = ~n170 & ~n171;
  assign n173 = pi111  & ~n172;
  assign n174 = ~n169 & ~n173;
  assign n175 = ~pi109  & ~n174;
  assign n176 = ~pi110  & ~n172;
  assign n177 = pi110  & ~n174;
  assign n178 = ~n176 & ~n177;
  assign n179 = pi109  & ~n178;
  assign n180 = ~n175 & ~n179;
  assign n181 = ~pi107  & ~n180;
  assign n182 = ~pi108  & ~n178;
  assign n183 = pi108  & ~n180;
  assign n184 = ~n182 & ~n183;
  assign n185 = pi107  & ~n184;
  assign n186 = ~n181 & ~n185;
  assign n187 = ~pi105  & ~n186;
  assign n188 = ~pi106  & ~n184;
  assign n189 = pi106  & ~n186;
  assign n190 = ~n188 & ~n189;
  assign n191 = pi105  & ~n190;
  assign n192 = ~n187 & ~n191;
  assign n193 = ~pi103  & ~n192;
  assign n194 = ~pi104  & ~n190;
  assign n195 = pi104  & ~n192;
  assign n196 = ~n194 & ~n195;
  assign n197 = pi103  & ~n196;
  assign n198 = ~n193 & ~n197;
  assign n199 = ~pi101  & ~n198;
  assign n200 = ~pi102  & ~n196;
  assign n201 = pi102  & ~n198;
  assign n202 = ~n200 & ~n201;
  assign n203 = pi101  & ~n202;
  assign n204 = ~n199 & ~n203;
  assign n205 = ~pi99  & ~n204;
  assign n206 = ~pi100  & ~n202;
  assign n207 = pi100  & ~n204;
  assign n208 = ~n206 & ~n207;
  assign n209 = pi99  & ~n208;
  assign n210 = ~n205 & ~n209;
  assign n211 = ~pi97  & ~n210;
  assign n212 = ~pi98  & ~n208;
  assign n213 = pi98  & ~n210;
  assign n214 = ~n212 & ~n213;
  assign n215 = pi97  & ~n214;
  assign n216 = ~n211 & ~n215;
  assign n217 = ~pi95  & ~n216;
  assign n218 = ~pi96  & ~n214;
  assign n219 = pi96  & ~n216;
  assign n220 = ~n218 & ~n219;
  assign n221 = pi95  & ~n220;
  assign n222 = ~n217 & ~n221;
  assign n223 = ~pi93  & ~n222;
  assign n224 = ~pi94  & ~n220;
  assign n225 = pi94  & ~n222;
  assign n226 = ~n224 & ~n225;
  assign n227 = pi93  & ~n226;
  assign n228 = ~n223 & ~n227;
  assign n229 = ~pi91  & ~n228;
  assign n230 = ~pi92  & ~n226;
  assign n231 = pi92  & ~n228;
  assign n232 = ~n230 & ~n231;
  assign n233 = pi91  & ~n232;
  assign n234 = ~n229 & ~n233;
  assign n235 = ~pi89  & ~n234;
  assign n236 = ~pi90  & ~n232;
  assign n237 = pi90  & ~n234;
  assign n238 = ~n236 & ~n237;
  assign n239 = pi89  & ~n238;
  assign n240 = ~n235 & ~n239;
  assign n241 = ~pi87  & ~n240;
  assign n242 = ~pi88  & ~n238;
  assign n243 = pi88  & ~n240;
  assign n244 = ~n242 & ~n243;
  assign n245 = pi87  & ~n244;
  assign n246 = ~n241 & ~n245;
  assign n247 = ~pi85  & ~n246;
  assign n248 = ~pi86  & ~n244;
  assign n249 = pi86  & ~n246;
  assign n250 = ~n248 & ~n249;
  assign n251 = pi85  & ~n250;
  assign n252 = ~n247 & ~n251;
  assign n253 = ~pi83  & ~n252;
  assign n254 = ~pi84  & ~n250;
  assign n255 = pi84  & ~n252;
  assign n256 = ~n254 & ~n255;
  assign n257 = pi83  & ~n256;
  assign n258 = ~n253 & ~n257;
  assign n259 = ~pi81  & ~n258;
  assign n260 = ~pi82  & ~n256;
  assign n261 = pi82  & ~n258;
  assign n262 = ~n260 & ~n261;
  assign n263 = pi81  & ~n262;
  assign n264 = ~n259 & ~n263;
  assign n265 = ~pi79  & ~n264;
  assign n266 = ~pi80  & ~n262;
  assign n267 = pi80  & ~n264;
  assign n268 = ~n266 & ~n267;
  assign n269 = pi79  & ~n268;
  assign n270 = ~n265 & ~n269;
  assign n271 = ~pi77  & ~n270;
  assign n272 = ~pi78  & ~n268;
  assign n273 = pi78  & ~n270;
  assign n274 = ~n272 & ~n273;
  assign n275 = pi77  & ~n274;
  assign n276 = ~n271 & ~n275;
  assign n277 = ~pi75  & ~n276;
  assign n278 = ~pi76  & ~n274;
  assign n279 = pi76  & ~n276;
  assign n280 = ~n278 & ~n279;
  assign n281 = pi75  & ~n280;
  assign n282 = ~n277 & ~n281;
  assign n283 = ~pi73  & ~n282;
  assign n284 = ~pi74  & ~n280;
  assign n285 = pi74  & ~n282;
  assign n286 = ~n284 & ~n285;
  assign n287 = pi73  & ~n286;
  assign n288 = ~n283 & ~n287;
  assign n289 = ~pi71  & ~n288;
  assign n290 = ~pi72  & ~n286;
  assign n291 = pi72  & ~n288;
  assign n292 = ~n290 & ~n291;
  assign n293 = pi71  & ~n292;
  assign n294 = ~n289 & ~n293;
  assign n295 = ~pi69  & ~n294;
  assign n296 = ~pi70  & ~n292;
  assign n297 = pi70  & ~n294;
  assign n298 = ~n296 & ~n297;
  assign n299 = pi69  & ~n298;
  assign n300 = ~n295 & ~n299;
  assign n301 = ~pi67  & ~n300;
  assign n302 = ~pi68  & ~n298;
  assign n303 = pi68  & ~n300;
  assign n304 = ~n302 & ~n303;
  assign n305 = pi67  & ~n304;
  assign n306 = ~n301 & ~n305;
  assign n307 = ~pi65  & ~n306;
  assign n308 = ~pi66  & ~n304;
  assign n309 = pi66  & ~n306;
  assign n310 = ~n308 & ~n309;
  assign n311 = pi65  & ~n310;
  assign n312 = ~n307 & ~n311;
  assign n313 = ~pi63  & ~n312;
  assign n314 = ~pi64  & ~n310;
  assign n315 = pi64  & ~n312;
  assign n316 = ~n314 & ~n315;
  assign n317 = pi63  & ~n316;
  assign n318 = ~n313 & ~n317;
  assign n319 = ~pi61  & ~n318;
  assign n320 = ~pi62  & ~n316;
  assign n321 = pi62  & ~n318;
  assign n322 = ~n320 & ~n321;
  assign n323 = pi61  & ~n322;
  assign n324 = ~n319 & ~n323;
  assign n325 = ~pi59  & ~n324;
  assign n326 = ~pi60  & ~n322;
  assign n327 = pi60  & ~n324;
  assign n328 = ~n326 & ~n327;
  assign n329 = pi59  & ~n328;
  assign n330 = ~n325 & ~n329;
  assign n331 = ~pi57  & ~n330;
  assign n332 = ~pi58  & ~n328;
  assign n333 = pi58  & ~n330;
  assign n334 = ~n332 & ~n333;
  assign n335 = pi57  & ~n334;
  assign n336 = ~n331 & ~n335;
  assign n337 = ~pi55  & ~n336;
  assign n338 = ~pi56  & ~n334;
  assign n339 = pi56  & ~n336;
  assign n340 = ~n338 & ~n339;
  assign n341 = pi55  & ~n340;
  assign n342 = ~n337 & ~n341;
  assign n343 = ~pi53  & ~n342;
  assign n344 = ~pi54  & ~n340;
  assign n345 = pi54  & ~n342;
  assign n346 = ~n344 & ~n345;
  assign n347 = pi53  & ~n346;
  assign n348 = ~n343 & ~n347;
  assign n349 = ~pi51  & ~n348;
  assign n350 = ~pi52  & ~n346;
  assign n351 = pi52  & ~n348;
  assign n352 = ~n350 & ~n351;
  assign n353 = pi51  & ~n352;
  assign n354 = ~n349 & ~n353;
  assign n355 = ~pi49  & ~n354;
  assign n356 = ~pi50  & ~n352;
  assign n357 = pi50  & ~n354;
  assign n358 = ~n356 & ~n357;
  assign n359 = pi49  & ~n358;
  assign n360 = ~n355 & ~n359;
  assign n361 = ~pi47  & ~n360;
  assign n362 = ~pi48  & ~n358;
  assign n363 = pi48  & ~n360;
  assign n364 = ~n362 & ~n363;
  assign n365 = pi47  & ~n364;
  assign n366 = ~n361 & ~n365;
  assign n367 = ~pi45  & ~n366;
  assign n368 = ~pi46  & ~n364;
  assign n369 = pi46  & ~n366;
  assign n370 = ~n368 & ~n369;
  assign n371 = pi45  & ~n370;
  assign n372 = ~n367 & ~n371;
  assign n373 = ~pi43  & ~n372;
  assign n374 = ~pi44  & ~n370;
  assign n375 = pi44  & ~n372;
  assign n376 = ~n374 & ~n375;
  assign n377 = pi43  & ~n376;
  assign n378 = ~n373 & ~n377;
  assign n379 = ~pi41  & ~n378;
  assign n380 = ~pi42  & ~n376;
  assign n381 = pi42  & ~n378;
  assign n382 = ~n380 & ~n381;
  assign n383 = pi41  & ~n382;
  assign n384 = ~n379 & ~n383;
  assign n385 = ~pi39  & ~n384;
  assign n386 = ~pi40  & ~n382;
  assign n387 = pi40  & ~n384;
  assign n388 = ~n386 & ~n387;
  assign n389 = pi39  & ~n388;
  assign n390 = ~n385 & ~n389;
  assign n391 = ~pi37  & ~n390;
  assign n392 = ~pi38  & ~n388;
  assign n393 = pi38  & ~n390;
  assign n394 = ~n392 & ~n393;
  assign n395 = pi37  & ~n394;
  assign n396 = ~n391 & ~n395;
  assign n397 = ~pi35  & ~n396;
  assign n398 = ~pi36  & ~n394;
  assign n399 = pi36  & ~n396;
  assign n400 = ~n398 & ~n399;
  assign n401 = pi35  & ~n400;
  assign n402 = ~n397 & ~n401;
  assign n403 = ~pi33  & ~n402;
  assign n404 = ~pi34  & ~n400;
  assign n405 = pi34  & ~n402;
  assign n406 = ~n404 & ~n405;
  assign n407 = pi33  & ~n406;
  assign n408 = ~n403 & ~n407;
  assign n409 = ~pi31  & ~n408;
  assign n410 = ~pi32  & ~n406;
  assign n411 = pi32  & ~n408;
  assign n412 = ~n410 & ~n411;
  assign n413 = pi31  & ~n412;
  assign n414 = ~n409 & ~n413;
  assign n415 = ~pi29  & ~n414;
  assign n416 = ~pi30  & ~n412;
  assign n417 = pi30  & ~n414;
  assign n418 = ~n416 & ~n417;
  assign n419 = pi29  & ~n418;
  assign n420 = ~n415 & ~n419;
  assign n421 = ~pi27  & ~n420;
  assign n422 = ~pi28  & ~n418;
  assign n423 = pi28  & ~n420;
  assign n424 = ~n422 & ~n423;
  assign n425 = pi27  & ~n424;
  assign n426 = ~n421 & ~n425;
  assign n427 = ~pi25  & ~n426;
  assign n428 = ~pi26  & ~n424;
  assign n429 = pi26  & ~n426;
  assign n430 = ~n428 & ~n429;
  assign n431 = pi25  & ~n430;
  assign n432 = ~n427 & ~n431;
  assign n433 = ~pi23  & ~n432;
  assign n434 = ~pi24  & ~n430;
  assign n435 = pi24  & ~n432;
  assign n436 = ~n434 & ~n435;
  assign n437 = pi23  & ~n436;
  assign n438 = ~n433 & ~n437;
  assign n439 = ~pi21  & ~n438;
  assign n440 = ~pi22  & ~n436;
  assign n441 = pi22  & ~n438;
  assign n442 = ~n440 & ~n441;
  assign n443 = pi21  & ~n442;
  assign n444 = pi1  & ~pi2 ;
  assign n445 = ~pi3  & ~n444;
  assign n446 = ~pi4  & ~n445;
  assign n447 = ~pi5  & ~n446;
  assign n448 = ~pi6  & ~n447;
  assign n449 = ~pi7  & ~n448;
  assign n450 = ~pi8  & ~n449;
  assign n451 = ~pi9  & ~n450;
  assign n452 = ~pi10  & ~n451;
  assign n453 = ~pi11  & ~n452;
  assign n454 = ~pi12  & ~n453;
  assign n455 = ~pi13  & ~n454;
  assign n456 = ~pi14  & ~n455;
  assign n457 = ~pi15  & ~n456;
  assign n458 = ~pi16  & ~n457;
  assign n459 = ~pi17  & ~n458;
  assign n460 = ~pi18  & ~n459;
  assign n461 = ~pi19  & ~n460;
  assign n462 = ~pi20  & ~n461;
  assign n463 = ~n439 & ~n462;
  assign n464 = ~n443 & n463;
  assign n465 = n442 & n462;
  assign po0  = ~n464 & ~n465;
  assign n467 = ~pi126  & ~pi127 ;
  assign n468 = ~pi124  & ~pi125 ;
  assign n469 = ~pi122  & ~pi123 ;
  assign n470 = ~pi120  & ~pi121 ;
  assign n471 = ~pi118  & ~pi119 ;
  assign n472 = ~pi116  & ~pi117 ;
  assign n473 = ~pi24  & ~pi25 ;
  assign n474 = ~pi22  & ~pi23 ;
  assign n475 = ~pi20  & ~pi21 ;
  assign n476 = ~pi18  & ~pi19 ;
  assign n477 = ~pi16  & ~pi17 ;
  assign n478 = ~pi14  & ~pi15 ;
  assign n479 = ~pi12  & ~pi13 ;
  assign n480 = ~pi10  & ~pi11 ;
  assign n481 = ~pi8  & ~pi9 ;
  assign n482 = ~pi6  & ~pi7 ;
  assign n483 = ~pi4  & ~pi5 ;
  assign n484 = ~pi2  & ~pi3 ;
  assign n485 = n483 & ~n484;
  assign n486 = n482 & ~n485;
  assign n487 = n481 & ~n486;
  assign n488 = n480 & ~n487;
  assign n489 = n479 & ~n488;
  assign n490 = n478 & ~n489;
  assign n491 = n477 & ~n490;
  assign n492 = n476 & ~n491;
  assign n493 = n475 & ~n492;
  assign n494 = n474 & ~n493;
  assign n495 = n473 & ~n494;
  assign n496 = ~pi26  & ~pi27 ;
  assign n497 = ~pi30  & ~pi31 ;
  assign n498 = ~pi32  & ~pi33 ;
  assign n499 = ~pi34  & ~pi35 ;
  assign n500 = ~pi36  & ~pi37 ;
  assign n501 = ~pi38  & ~pi39 ;
  assign n502 = ~pi40  & ~pi41 ;
  assign n503 = ~pi42  & ~pi43 ;
  assign n504 = ~pi44  & ~pi45 ;
  assign n505 = ~pi46  & ~pi47 ;
  assign n506 = ~pi48  & ~pi49 ;
  assign n507 = ~pi50  & ~pi51 ;
  assign n508 = ~pi52  & ~pi53 ;
  assign n509 = ~pi54  & ~pi55 ;
  assign n510 = ~pi56  & ~pi57 ;
  assign n511 = ~pi58  & ~pi59 ;
  assign n512 = ~pi60  & ~pi61 ;
  assign n513 = ~pi62  & ~pi63 ;
  assign n514 = ~pi64  & ~pi65 ;
  assign n515 = ~pi66  & ~pi67 ;
  assign n516 = ~pi68  & ~pi69 ;
  assign n517 = ~pi70  & ~pi71 ;
  assign n518 = ~pi72  & ~pi73 ;
  assign n519 = ~pi74  & ~pi75 ;
  assign n520 = ~pi76  & ~pi77 ;
  assign n521 = ~pi78  & ~pi79 ;
  assign n522 = ~pi80  & ~pi81 ;
  assign n523 = ~pi82  & ~pi83 ;
  assign n524 = ~pi84  & ~pi85 ;
  assign n525 = ~pi86  & ~pi87 ;
  assign n526 = ~pi88  & ~pi89 ;
  assign n527 = ~pi90  & ~pi91 ;
  assign n528 = ~pi92  & ~pi93 ;
  assign n529 = ~pi94  & ~pi95 ;
  assign n530 = ~pi96  & ~pi97 ;
  assign n531 = ~pi98  & ~pi99 ;
  assign n532 = ~pi102  & ~pi103 ;
  assign n533 = ~pi112  & ~pi113 ;
  assign n534 = ~pi110  & ~pi111 ;
  assign n535 = ~pi106  & ~pi107 ;
  assign n536 = ~pi108  & ~pi109 ;
  assign n537 = ~n535 & n536;
  assign n538 = n534 & ~n537;
  assign n539 = n533 & ~n538;
  assign n540 = n532 & ~n539;
  assign n541 = ~pi104  & ~pi105 ;
  assign n542 = n538 & ~n541;
  assign n543 = n534 & ~n536;
  assign n544 = n541 & n543;
  assign n545 = n533 & ~n544;
  assign n546 = ~n542 & n545;
  assign n547 = ~n532 & ~n546;
  assign n548 = ~n540 & ~n547;
  assign n549 = ~pi100  & ~pi101 ;
  assign n550 = n548 & ~n549;
  assign n551 = n546 & n549;
  assign n552 = ~n550 & ~n551;
  assign n553 = ~n531 & ~n552;
  assign n554 = n531 & n548;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~n530 & ~n555;
  assign n557 = n530 & ~n552;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~n529 & ~n558;
  assign n560 = n529 & ~n555;
  assign n561 = ~n559 & ~n560;
  assign n562 = ~n528 & ~n561;
  assign n563 = n528 & ~n558;
  assign n564 = ~n562 & ~n563;
  assign n565 = ~n527 & ~n564;
  assign n566 = n527 & ~n561;
  assign n567 = ~n565 & ~n566;
  assign n568 = ~n526 & ~n567;
  assign n569 = n526 & ~n564;
  assign n570 = ~n568 & ~n569;
  assign n571 = ~n525 & ~n570;
  assign n572 = n525 & ~n567;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~n524 & ~n573;
  assign n575 = n524 & ~n570;
  assign n576 = ~n574 & ~n575;
  assign n577 = ~n523 & ~n576;
  assign n578 = n523 & ~n573;
  assign n579 = ~n577 & ~n578;
  assign n580 = ~n522 & ~n579;
  assign n581 = n522 & ~n576;
  assign n582 = ~n580 & ~n581;
  assign n583 = ~n521 & ~n582;
  assign n584 = n521 & ~n579;
  assign n585 = ~n583 & ~n584;
  assign n586 = ~n520 & ~n585;
  assign n587 = n520 & ~n582;
  assign n588 = ~n586 & ~n587;
  assign n589 = ~n519 & ~n588;
  assign n590 = n519 & ~n585;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n518 & ~n591;
  assign n593 = n518 & ~n588;
  assign n594 = ~n592 & ~n593;
  assign n595 = ~n517 & ~n594;
  assign n596 = n517 & ~n591;
  assign n597 = ~n595 & ~n596;
  assign n598 = ~n516 & ~n597;
  assign n599 = n516 & ~n594;
  assign n600 = ~n598 & ~n599;
  assign n601 = ~n515 & ~n600;
  assign n602 = n515 & ~n597;
  assign n603 = ~n601 & ~n602;
  assign n604 = ~n514 & ~n603;
  assign n605 = n514 & ~n600;
  assign n606 = ~n604 & ~n605;
  assign n607 = ~n513 & ~n606;
  assign n608 = n513 & ~n603;
  assign n609 = ~n607 & ~n608;
  assign n610 = ~n512 & ~n609;
  assign n611 = n512 & ~n606;
  assign n612 = ~n610 & ~n611;
  assign n613 = ~n511 & ~n612;
  assign n614 = n511 & ~n609;
  assign n615 = ~n613 & ~n614;
  assign n616 = ~n510 & ~n615;
  assign n617 = n510 & ~n612;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~n509 & ~n618;
  assign n620 = n509 & ~n615;
  assign n621 = ~n619 & ~n620;
  assign n622 = ~n508 & ~n621;
  assign n623 = n508 & ~n618;
  assign n624 = ~n622 & ~n623;
  assign n625 = ~n507 & ~n624;
  assign n626 = n507 & ~n621;
  assign n627 = ~n625 & ~n626;
  assign n628 = ~n506 & ~n627;
  assign n629 = n506 & ~n624;
  assign n630 = ~n628 & ~n629;
  assign n631 = ~n505 & ~n630;
  assign n632 = n505 & ~n627;
  assign n633 = ~n631 & ~n632;
  assign n634 = ~n504 & ~n633;
  assign n635 = n504 & ~n630;
  assign n636 = ~n634 & ~n635;
  assign n637 = ~n503 & ~n636;
  assign n638 = n503 & ~n633;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~n502 & ~n639;
  assign n641 = n502 & ~n636;
  assign n642 = ~n640 & ~n641;
  assign n643 = ~n501 & ~n642;
  assign n644 = n501 & ~n639;
  assign n645 = ~n643 & ~n644;
  assign n646 = ~n500 & ~n645;
  assign n647 = n500 & ~n642;
  assign n648 = ~n646 & ~n647;
  assign n649 = ~n499 & ~n648;
  assign n650 = n499 & ~n645;
  assign n651 = ~n649 & ~n650;
  assign n652 = ~n498 & ~n651;
  assign n653 = n498 & ~n648;
  assign n654 = ~n652 & ~n653;
  assign n655 = ~n497 & ~n654;
  assign n656 = n497 & ~n651;
  assign n657 = ~n655 & ~n656;
  assign n658 = n496 & ~n657;
  assign n659 = ~pi114  & ~pi115 ;
  assign n660 = ~pi28  & ~pi29 ;
  assign n661 = ~n657 & ~n660;
  assign n662 = ~n654 & n660;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~n496 & ~n663;
  assign n665 = ~n495 & n659;
  assign n666 = ~n658 & n665;
  assign n667 = ~n664 & n666;
  assign n668 = n495 & n659;
  assign n669 = n663 & n668;
  assign n670 = n472 & ~n669;
  assign n671 = ~n667 & n670;
  assign n672 = n471 & ~n671;
  assign n673 = n470 & ~n672;
  assign n674 = n469 & ~n673;
  assign n675 = n468 & ~n674;
  assign po1  = ~n467 | n675;
  assign n677 = n467 & n468;
  assign n678 = n469 & n470;
  assign n679 = n471 & n472;
  assign n680 = n533 & n659;
  assign n681 = n524 & n525;
  assign n682 = n535 & n541;
  assign n683 = n526 & n527;
  assign n684 = n532 & n549;
  assign n685 = n530 & n531;
  assign n686 = n528 & n529;
  assign n687 = n685 & ~n686;
  assign n688 = n684 & ~n687;
  assign n689 = ~n683 & n688;
  assign n690 = n683 & n684;
  assign n691 = ~n685 & n690;
  assign n692 = n682 & ~n691;
  assign n693 = ~n689 & n692;
  assign n694 = ~n681 & n693;
  assign n695 = n534 & n536;
  assign n696 = n681 & n682;
  assign n697 = ~n688 & n696;
  assign n698 = n695 & ~n697;
  assign n699 = ~n694 & n698;
  assign n700 = n680 & ~n699;
  assign n701 = n679 & ~n700;
  assign n702 = n678 & ~n701;
  assign n703 = n522 & n523;
  assign n704 = n702 & ~n703;
  assign n705 = ~n693 & n695;
  assign n706 = n680 & ~n705;
  assign n707 = n679 & ~n706;
  assign n708 = n678 & n703;
  assign n709 = ~n707 & n708;
  assign n710 = n520 & n521;
  assign n711 = n518 & n519;
  assign n712 = n516 & n517;
  assign n713 = n514 & n515;
  assign n714 = n512 & n513;
  assign n715 = n510 & n511;
  assign n716 = n508 & n509;
  assign n717 = n506 & n507;
  assign n718 = n504 & n505;
  assign n719 = n502 & n503;
  assign n720 = n500 & n501;
  assign n721 = n498 & n499;
  assign n722 = n497 & n660;
  assign n723 = n473 & n496;
  assign n724 = n474 & n475;
  assign n725 = n476 & n477;
  assign n726 = n478 & n479;
  assign n727 = n480 & n481;
  assign n728 = n482 & n483;
  assign n729 = n727 & ~n728;
  assign n730 = n726 & ~n729;
  assign n731 = n725 & ~n730;
  assign n732 = n724 & ~n731;
  assign n733 = n723 & ~n732;
  assign n734 = n722 & ~n733;
  assign n735 = n721 & ~n734;
  assign n736 = n720 & ~n735;
  assign n737 = n719 & ~n736;
  assign n738 = n718 & ~n737;
  assign n739 = n717 & ~n738;
  assign n740 = n716 & ~n739;
  assign n741 = n715 & ~n740;
  assign n742 = n714 & ~n741;
  assign n743 = n713 & ~n742;
  assign n744 = n712 & ~n743;
  assign n745 = n711 & ~n744;
  assign n746 = n710 & ~n745;
  assign n747 = n677 & ~n709;
  assign n748 = ~n704 & n747;
  assign n749 = ~n746 & n748;
  assign n750 = n677 & n710;
  assign n751 = ~n702 & n750;
  assign n752 = ~n745 & n751;
  assign po2  = ~n749 & ~n752;
  assign n754 = n677 & n678;
  assign n755 = n681 & n703;
  assign n756 = n710 & n711;
  assign n757 = n712 & n713;
  assign n758 = n714 & n715;
  assign n759 = n716 & n717;
  assign n760 = n718 & n719;
  assign n761 = n720 & n721;
  assign n762 = n722 & n723;
  assign n763 = n724 & n725;
  assign n764 = n726 & n727;
  assign n765 = n763 & ~n764;
  assign n766 = n762 & ~n765;
  assign n767 = n761 & ~n766;
  assign n768 = n760 & ~n767;
  assign n769 = n759 & ~n768;
  assign n770 = n758 & ~n769;
  assign n771 = n757 & ~n770;
  assign n772 = n756 & ~n771;
  assign n773 = n755 & ~n772;
  assign n774 = n679 & n680;
  assign n775 = n682 & n695;
  assign n776 = n683 & n686;
  assign n777 = n684 & n685;
  assign n778 = ~n776 & n777;
  assign n779 = n775 & ~n778;
  assign n780 = n774 & ~n779;
  assign n781 = ~n773 & n780;
  assign n782 = n775 & ~n777;
  assign n783 = n774 & ~n782;
  assign n784 = n773 & n783;
  assign n785 = n754 & ~n781;
  assign po3  = n784 | ~n785;
  assign n787 = n754 & n774;
  assign n788 = n775 & n777;
  assign n789 = n755 & n776;
  assign n790 = n758 & n759;
  assign n791 = n762 & n763;
  assign n792 = n760 & n761;
  assign n793 = ~n791 & n792;
  assign n794 = n790 & ~n793;
  assign n795 = n756 & n757;
  assign n796 = ~n794 & n795;
  assign n797 = n789 & ~n796;
  assign n798 = n788 & ~n797;
  assign po4  = ~n787 | n798;
  assign n800 = n787 & n788;
  assign n801 = n789 & n795;
  assign n802 = n790 & n792;
  assign n803 = n801 & ~n802;
  assign po5  = ~n800 | n803;
  assign po6  = ~n800 | ~n801;
  assign n806 = ~pi0  & ~pi1 ;
  assign n807 = n484 & n806;
  assign n808 = n728 & n807;
  assign n809 = n764 & n808;
  assign n810 = n791 & n809;
  assign n811 = n802 & n810;
  assign po7 = po6  | ~n811;
endmodule
