module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330,
    n332, n333, n334;
  assign n92 = ~pi9  & ~pi10 ;
  assign n93 = pi9  & pi10 ;
  assign n94 = ~n92 & ~n93;
  assign n95 = pi11  & ~n92;
  assign n96 = ~pi11  & n92;
  assign n97 = ~n95 & ~n96;
  assign n98 = ~pi12  & ~n95;
  assign n99 = pi12  & n95;
  assign n100 = ~n98 & ~n99;
  assign n101 = ~pi13  & n98;
  assign n102 = pi13  & ~n98;
  assign n103 = ~n101 & ~n102;
  assign n104 = pi14  & ~n101;
  assign n105 = ~pi14  & n101;
  assign n106 = ~n104 & ~n105;
  assign n107 = pi15  & n104;
  assign n108 = ~pi16  & ~n107;
  assign n109 = pi16  & n107;
  assign n110 = ~n108 & ~n109;
  assign n111 = pi17  & ~n108;
  assign n112 = ~pi17  & n108;
  assign n113 = ~n111 & ~n112;
  assign n114 = ~pi18  & ~n111;
  assign n115 = pi18  & n111;
  assign n116 = ~n114 & ~n115;
  assign n117 = pi19  & ~n114;
  assign n118 = ~pi19  & n114;
  assign n119 = ~n117 & ~n118;
  assign n120 = pi20  & n117;
  assign n121 = ~pi21  & ~n120;
  assign n122 = pi21  & n120;
  assign n123 = ~n121 & ~n122;
  assign n124 = ~pi22  & n121;
  assign n125 = pi22  & ~n121;
  assign n126 = ~n124 & ~n125;
  assign n127 = pi23  & ~n124;
  assign n128 = ~pi23  & n124;
  assign n129 = ~n127 & ~n128;
  assign n130 = pi24  & n127;
  assign n131 = pi25  & n130;
  assign n132 = ~pi26  & ~n131;
  assign n133 = pi26  & n131;
  assign n134 = ~n132 & ~n133;
  assign n135 = pi27  & ~n132;
  assign n136 = ~pi27  & n132;
  assign n137 = ~n135 & ~n136;
  assign n138 = pi28  & n135;
  assign n139 = ~pi28  & ~n135;
  assign n140 = ~n138 & ~n139;
  assign n141 = ~pi9  & pi29 ;
  assign n142 = n140 & n141;
  assign n143 = n137 & n142;
  assign n144 = ~n134 & n143;
  assign n145 = ~pi25  & ~n130;
  assign n146 = ~n131 & ~n145;
  assign n147 = n144 & n146;
  assign n148 = ~pi24  & ~n127;
  assign n149 = ~n130 & ~n148;
  assign n150 = n147 & n149;
  assign n151 = n129 & n150;
  assign n152 = ~n126 & n151;
  assign n153 = ~n123 & n152;
  assign n154 = ~pi20  & ~n117;
  assign n155 = ~n120 & ~n154;
  assign n156 = n153 & n155;
  assign n157 = n119 & n156;
  assign n158 = ~n116 & n157;
  assign n159 = n113 & n158;
  assign n160 = ~n110 & n159;
  assign n161 = ~pi15  & ~n104;
  assign n162 = ~n107 & ~n161;
  assign n163 = n160 & n162;
  assign n164 = n106 & n163;
  assign n165 = ~n103 & n164;
  assign n166 = ~n100 & n165;
  assign n167 = n97 & n166;
  assign n168 = ~n94 & n167;
  assign n169 = pi8  & n168;
  assign n170 = pi7  & n169;
  assign n171 = pi6  & n170;
  assign n172 = pi5  & n171;
  assign n173 = pi4  & n172;
  assign n174 = pi3  & n173;
  assign n175 = pi2  & n174;
  assign n176 = pi1  & n175;
  assign n177 = pi0  & n176;
  assign n178 = pi29  & n138;
  assign n179 = ~n177 & ~n178;
  assign n180 = ~pi1  & ~pi2 ;
  assign n181 = ~pi3  & n180;
  assign n182 = ~pi4  & n181;
  assign n183 = ~pi5  & n182;
  assign n184 = ~pi6  & n183;
  assign n185 = ~pi7  & n184;
  assign n186 = ~pi8  & n185;
  assign n187 = n94 & n186;
  assign n188 = ~n97 & n187;
  assign n189 = n100 & n188;
  assign n190 = n103 & n189;
  assign n191 = ~n106 & n190;
  assign n192 = ~n162 & n191;
  assign n193 = n110 & n192;
  assign n194 = ~n113 & n193;
  assign n195 = n116 & n194;
  assign n196 = ~n119 & n195;
  assign n197 = ~n155 & n196;
  assign n198 = n123 & n197;
  assign n199 = n126 & n198;
  assign n200 = ~n129 & n199;
  assign n201 = ~n149 & n200;
  assign n202 = ~n146 & n201;
  assign n203 = n134 & n202;
  assign n204 = ~n137 & n203;
  assign n205 = ~n140 & n204;
  assign n206 = pi9  & n205;
  assign n207 = n178 & ~n206;
  assign po0  = n179 | n207;
  assign n209 = ~pi39  & ~pi40 ;
  assign n210 = pi41  & ~n209;
  assign n211 = ~pi42  & ~n210;
  assign n212 = ~pi43  & n211;
  assign n213 = pi44  & ~n212;
  assign n214 = pi45  & n213;
  assign n215 = ~pi46  & ~n214;
  assign n216 = pi47  & ~n215;
  assign n217 = ~pi48  & ~n216;
  assign n218 = pi49  & ~n217;
  assign n219 = pi50  & n218;
  assign n220 = ~pi51  & ~n219;
  assign n221 = ~pi52  & n220;
  assign n222 = pi53  & ~n221;
  assign n223 = pi54  & n222;
  assign n224 = pi55  & n223;
  assign n225 = ~pi56  & ~n224;
  assign n226 = pi57  & ~n225;
  assign n227 = pi58  & n226;
  assign n228 = pi59  & n227;
  assign n229 = pi0  & ~n228;
  assign n230 = ~pi0  & ~pi30 ;
  assign n231 = n228 & ~n230;
  assign n232 = pi39  & pi40 ;
  assign n233 = ~n209 & ~n232;
  assign n234 = ~pi41  & n209;
  assign n235 = ~n210 & ~n234;
  assign n236 = pi42  & n210;
  assign n237 = ~n211 & ~n236;
  assign n238 = pi43  & ~n211;
  assign n239 = ~n212 & ~n238;
  assign n240 = ~pi44  & n212;
  assign n241 = ~n213 & ~n240;
  assign n242 = pi46  & n214;
  assign n243 = ~n215 & ~n242;
  assign n244 = ~pi47  & n215;
  assign n245 = ~n216 & ~n244;
  assign n246 = pi48  & n216;
  assign n247 = ~n217 & ~n246;
  assign n248 = ~pi49  & n217;
  assign n249 = ~n218 & ~n248;
  assign n250 = pi51  & n219;
  assign n251 = ~n220 & ~n250;
  assign n252 = pi52  & ~n220;
  assign n253 = ~n221 & ~n252;
  assign n254 = ~pi53  & n221;
  assign n255 = ~n222 & ~n254;
  assign n256 = pi56  & n224;
  assign n257 = ~n225 & ~n256;
  assign n258 = ~pi57  & n225;
  assign n259 = ~n226 & ~n258;
  assign n260 = pi30  & ~pi39 ;
  assign n261 = pi59  & n260;
  assign n262 = ~pi58  & ~n226;
  assign n263 = ~n227 & ~n262;
  assign n264 = n261 & n263;
  assign n265 = n259 & n264;
  assign n266 = ~n257 & n265;
  assign n267 = ~pi55  & ~n223;
  assign n268 = ~n224 & ~n267;
  assign n269 = n266 & n268;
  assign n270 = ~pi54  & ~n222;
  assign n271 = ~n223 & ~n270;
  assign n272 = n269 & n271;
  assign n273 = n255 & n272;
  assign n274 = ~n253 & n273;
  assign n275 = ~n251 & n274;
  assign n276 = ~pi50  & ~n218;
  assign n277 = ~n219 & ~n276;
  assign n278 = n275 & n277;
  assign n279 = n249 & n278;
  assign n280 = ~n247 & n279;
  assign n281 = n245 & n280;
  assign n282 = ~n243 & n281;
  assign n283 = ~pi45  & ~n213;
  assign n284 = ~n214 & ~n283;
  assign n285 = n282 & n284;
  assign n286 = n241 & n285;
  assign n287 = ~n239 & n286;
  assign n288 = ~n237 & n287;
  assign n289 = n235 & n288;
  assign n290 = ~n233 & n289;
  assign n291 = pi38  & n290;
  assign n292 = pi37  & n291;
  assign n293 = pi36  & n292;
  assign n294 = pi35  & n293;
  assign n295 = pi34  & n294;
  assign n296 = pi33  & n295;
  assign n297 = pi32  & n296;
  assign n298 = pi31  & n297;
  assign n299 = ~pi31  & ~pi32 ;
  assign n300 = ~pi33  & n299;
  assign n301 = ~pi34  & n300;
  assign n302 = ~pi35  & n301;
  assign n303 = ~pi36  & n302;
  assign n304 = ~pi37  & n303;
  assign n305 = ~pi38  & n304;
  assign n306 = n233 & n305;
  assign n307 = ~n235 & n306;
  assign n308 = n237 & n307;
  assign n309 = n239 & n308;
  assign n310 = ~n241 & n309;
  assign n311 = ~n284 & n310;
  assign n312 = n243 & n311;
  assign n313 = ~n245 & n312;
  assign n314 = n247 & n313;
  assign n315 = ~n249 & n314;
  assign n316 = ~n277 & n315;
  assign n317 = n251 & n316;
  assign n318 = n253 & n317;
  assign n319 = ~n255 & n318;
  assign n320 = ~n271 & n319;
  assign n321 = ~n268 & n320;
  assign n322 = n257 & n321;
  assign n323 = ~n259 & n322;
  assign n324 = ~n263 & n323;
  assign n325 = pi39  & n324;
  assign n326 = n228 & ~n325;
  assign n327 = ~n298 & ~n326;
  assign n328 = ~n231 & n327;
  assign n329 = ~n179 & ~n328;
  assign n330 = ~n229 & n329;
  assign po1  = ~n207 & ~n330;
  assign n332 = pi0  & n228;
  assign n333 = pi30  & n332;
  assign n334 = ~n326 & ~n333;
  assign po2  = ~po0  & ~n334;
  assign po3  = 1'b0;
  assign po4  = 1'b0;
  assign po5  = 1'b0;
  assign po6  = 1'b0;
  assign po7  = 1'b0;
  assign po8  = 1'b0;
  assign po9  = 1'b0;
  assign po10  = 1'b0;
  assign po11  = 1'b0;
  assign po12  = 1'b0;
  assign po13  = 1'b0;
  assign po14  = 1'b0;
  assign po15  = 1'b0;
  assign po16  = 1'b0;
  assign po17  = 1'b0;
  assign po18  = 1'b0;
  assign po19  = 1'b0;
  assign po20  = 1'b0;
  assign po21  = 1'b0;
  assign po22  = 1'b0;
  assign po23  = 1'b0;
  assign po24  = 1'b0;
  assign po25  = 1'b0;
  assign po26  = 1'b0;
  assign po27  = 1'b0;
  assign po28  = 1'b0;
  assign po29  = 1'b0;
endmodule
