module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442,
    n444, n445, n446, n447, n448, n449, n450,
    n452, n453, n454, n455, n456, n457, n458,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n471, n472, n473, n474,
    n475, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n487, n488, n489, n490,
    n491, n492, n493, n495, n496, n497, n498,
    n499, n501, n502, n503, n504, n505, n506,
    n507, n508, n510, n511, n512, n513, n514,
    n515, n516, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n542, n543, n544,
    n545, n546, n547, n548, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n561, n562, n563, n564, n565, n566, n568,
    n569, n570, n571, n572, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590,
    n591, n593, n594, n595, n596, n597, n598,
    n599, n601, n602, n603, n604, n605, n606,
    n607, n609, n610, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n673,
    n674, n675, n676, n677, n678, n679, n681,
    n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760,
    n762, n763, n764, n765, n766, n767, n769,
    n770, n771, n772, n773, n774, n776, n777,
    n778, n779, n780, n781, n783, n784, n785,
    n786, n787, n788, n790, n791, n792, n793,
    n794, n795, n797, n798, n799, n800, n801,
    n802, n804, n805, n806, n807, n808, n809,
    n811, n812, n813, n814, n815, n816, n818,
    n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n843, n844, n845, n846, n847,
    n848, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862,
    n863, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n915,
    n916, n917, n918, n919, n920, n921, n923,
    n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952,
    n953, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967,
    n968, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1017,
    n1018, n1019, n1021, n1022, n1023, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1035, n1036, n1037, n1040,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1079,
    n1080, n1081, n1082, n1083, n1084, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1107, n1108, n1109, n1111, n1112,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1123, n1124, n1125, n1127,
    n1128, n1129, n1131, n1132, n1133, n1135,
    n1136, n1137, n1138, n1139, n1141, n1142,
    n1143, n1145, n1146, n1147, n1149, n1150,
    n1151, n1153, n1154, n1155, n1157, n1158,
    n1159, n1161, n1162, n1163, n1165, n1166,
    n1167, n1169, n1170, n1171, n1173, n1174,
    n1175, n1177, n1178, n1179, n1181, n1182,
    n1183, n1185, n1186, n1187, n1188, n1189,
    n1191, n1192, n1193, n1195, n1196, n1197,
    n1199, n1200, n1201, n1203, n1204, n1205,
    n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224,
    n1226, n1227, n1228, n1230, n1231, n1232,
    n1233, n1235, n1236, n1237, n1239, n1240,
    n1241, n1243, n1244, n1245, n1246, n1247,
    n1249, n1250, n1251, n1253, n1254, n1255,
    n1257, n1258, n1259, n1261, n1262, n1263,
    n1265, n1266, n1267, n1269, n1270, n1271,
    n1272, n1273, n1274, n1276, n1277, n1278,
    n1279, n1280, n1281, n1283, n1284, n1285,
    n1287, n1288, n1289, n1291, n1292, n1293,
    n1295, n1296, n1297, n1299, n1300, n1301,
    n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1321,
    n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1384, n1385,
    n1386, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404,
    n1406, n1407, n1408, n1409, n1410, n1411,
    n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1424,
    n1425, n1426, n1428, n1429, n1431, n1432,
    n1433, n1434, n1436, n1437, n1438, n1440,
    n1441, n1442, n1443, n1445, n1446, n1447,
    n1449, n1450, n1451, n1452, n1455, n1456,
    n1457, n1458, n1461, n1462, n1464, n1469,
    n1470, n1472;
  assign n291 = ~pi7 & ~pi13;
  assign n292 = ~pi14 & n291;
  assign n293 = ~pi4 & ~pi19;
  assign n294 = ~pi18 & n293;
  assign n295 = ~pi16 & n294;
  assign n296 = ~pi9 & ~pi11;
  assign n297 = ~pi6 & ~pi12;
  assign n298 = ~pi5 & n297;
  assign n299 = ~pi17 & ~pi21;
  assign n300 = ~pi8 & n299;
  assign n301 = ~pi22 & n296;
  assign n302 = n292 & n301;
  assign n303 = n298 & n300;
  assign n304 = n302 & n303;
  assign n305 = n295 & n304;
  assign n306 = pi54 & ~n305;
  assign n307 = ~pi0 & ~n306;
  assign n308 = ~pi5 & ~pi22;
  assign n309 = ~pi56 & ~n308;
  assign n310 = ~pi8 & ~pi21;
  assign n311 = n291 & n310;
  assign n312 = ~pi7 & n310;
  assign n313 = pi8 & pi21;
  assign n314 = ~pi13 & ~n313;
  assign n315 = ~n312 & ~n314;
  assign n316 = ~pi14 & ~n315;
  assign n317 = ~n311 & ~n316;
  assign n318 = pi7 & ~n310;
  assign n319 = ~n311 & ~n318;
  assign n320 = ~pi14 & ~n319;
  assign n321 = ~pi10 & ~n320;
  assign n322 = ~n317 & n321;
  assign n323 = ~pi14 & n310;
  assign n324 = pi10 & n291;
  assign n325 = n323 & n324;
  assign n326 = ~n322 & ~n325;
  assign n327 = ~pi17 & n297;
  assign n328 = n308 & n327;
  assign n329 = n295 & n328;
  assign n330 = ~n326 & n329;
  assign n331 = ~n309 & ~n330;
  assign n332 = n296 & ~n331;
  assign n333 = ~pi56 & ~n296;
  assign n334 = n308 & n333;
  assign n335 = ~n332 & ~n334;
  assign n336 = pi54 & ~n335;
  assign n337 = ~n307 & ~n336;
  assign n338 = ~pi3 & ~pi129;
  assign po15 = n337 | ~n338;
  assign n340 = ~pi17 & pi54;
  assign n341 = ~pi5 & ~pi6;
  assign n342 = n291 & n341;
  assign n343 = ~pi10 & ~pi22;
  assign n344 = n342 & n343;
  assign n345 = n295 & n344;
  assign n346 = ~pi11 & ~pi12;
  assign n347 = n323 & n346;
  assign n348 = n345 & n347;
  assign n349 = n340 & ~n348;
  assign n350 = ~pi1 & ~n349;
  assign n351 = ~pi14 & pi54;
  assign n352 = n343 & n351;
  assign n353 = ~pi5 & ~pi7;
  assign n354 = n297 & n353;
  assign n355 = pi13 & n354;
  assign n356 = pi6 & pi12;
  assign n357 = ~pi7 & ~n356;
  assign n358 = ~n298 & ~n357;
  assign n359 = ~n297 & ~n353;
  assign n360 = ~pi13 & ~n354;
  assign n361 = ~n359 & n360;
  assign n362 = ~n358 & n361;
  assign n363 = ~pi9 & ~n355;
  assign n364 = ~n362 & n363;
  assign n365 = ~pi8 & ~pi11;
  assign n366 = n299 & n365;
  assign n367 = n291 & n298;
  assign n368 = pi9 & ~n367;
  assign n369 = n352 & n366;
  assign n370 = n295 & n369;
  assign n371 = ~n368 & n370;
  assign n372 = ~n364 & n371;
  assign n373 = ~n350 & ~n372;
  assign po16 = ~n338 | n373;
  assign n375 = ~pi47 & ~pi48;
  assign n376 = ~pi45 & n375;
  assign n377 = ~pi41 & ~pi43;
  assign n378 = ~pi42 & ~pi44;
  assign n379 = ~pi38 & ~pi50;
  assign n380 = ~pi40 & ~pi46;
  assign n381 = n379 & n380;
  assign n382 = n378 & n381;
  assign n383 = n377 & n382;
  assign n384 = n376 & n383;
  assign n385 = pi82 & ~n384;
  assign n386 = pi122 & pi127;
  assign n387 = ~pi82 & n386;
  assign n388 = ~pi15 & ~pi20;
  assign n389 = ~pi24 & ~pi49;
  assign n390 = n388 & n389;
  assign n391 = pi82 & ~n390;
  assign n392 = ~n387 & ~n391;
  assign n393 = ~n385 & n392;
  assign n394 = pi2 & ~n393;
  assign n395 = ~pi40 & n378;
  assign n396 = ~pi41 & ~pi46;
  assign n397 = n379 & n396;
  assign n398 = ~pi45 & n390;
  assign n399 = ~pi43 & ~pi47;
  assign n400 = ~pi48 & n399;
  assign n401 = ~pi2 & n400;
  assign n402 = n398 & n401;
  assign n403 = n397 & n402;
  assign n404 = n395 & n403;
  assign n405 = pi82 & ~n404;
  assign n406 = ~pi65 & ~n386;
  assign n407 = ~n405 & n406;
  assign n408 = ~n394 & ~n407;
  assign po17 = ~pi129 & ~n408;
  assign n410 = pi0 & ~pi113;
  assign n411 = ~pi123 & n410;
  assign n412 = ~pi9 & ~pi14;
  assign n413 = ~pi12 & n366;
  assign n414 = n412 & n413;
  assign n415 = n345 & n414;
  assign n416 = ~pi61 & ~pi118;
  assign n417 = ~n415 & n416;
  assign n418 = ~n411 & ~n417;
  assign po18 = ~pi129 & ~n418;
  assign n420 = pi4 & ~pi54;
  assign n421 = ~pi16 & pi54;
  assign n422 = n294 & n421;
  assign n423 = n300 & n422;
  assign n424 = ~pi11 & n423;
  assign n425 = pi10 & ~pi22;
  assign n426 = n412 & n425;
  assign n427 = n367 & n426;
  assign n428 = n424 & n427;
  assign n429 = ~n420 & ~n428;
  assign po19 = n338 & ~n429;
  assign n431 = pi5 & ~pi54;
  assign n432 = n343 & n412;
  assign n433 = ~pi13 & n432;
  assign n434 = ~pi59 & n366;
  assign n435 = n433 & n434;
  assign n436 = n354 & n421;
  assign n437 = ~pi25 & pi28;
  assign n438 = ~pi29 & n437;
  assign n439 = n294 & n438;
  assign n440 = n436 & n439;
  assign n441 = n435 & n440;
  assign n442 = ~n431 & ~n441;
  assign po20 = n338 & ~n442;
  assign n444 = pi6 & ~pi54;
  assign n445 = ~pi28 & ~pi29;
  assign n446 = pi25 & n445;
  assign n447 = n294 & n446;
  assign n448 = n436 & n447;
  assign n449 = n435 & n448;
  assign n450 = ~n444 & ~n449;
  assign po21 = n338 & ~n450;
  assign n452 = pi7 & ~pi54;
  assign n453 = ~pi11 & n354;
  assign n454 = pi8 & n299;
  assign n455 = n422 & n454;
  assign n456 = n433 & n453;
  assign n457 = n455 & n456;
  assign n458 = ~n452 & ~n457;
  assign po22 = n338 & ~n458;
  assign n460 = pi8 & ~pi54;
  assign n461 = n342 & n432;
  assign n462 = ~pi12 & n461;
  assign n463 = n293 & n421;
  assign n464 = ~pi17 & ~pi18;
  assign n465 = n365 & n464;
  assign n466 = pi21 & n463;
  assign n467 = n465 & n466;
  assign n468 = n462 & n467;
  assign n469 = ~n460 & ~n468;
  assign po23 = n338 & ~n469;
  assign n471 = pi9 & ~pi54;
  assign n472 = pi11 & n354;
  assign n473 = n433 & n472;
  assign n474 = n423 & n473;
  assign n475 = ~n471 & ~n474;
  assign po24 = n338 & ~n475;
  assign n477 = pi10 & ~pi54;
  assign n478 = ~pi9 & ~pi18;
  assign n479 = n300 & n478;
  assign n480 = n343 & n479;
  assign n481 = ~pi13 & pi14;
  assign n482 = n463 & n481;
  assign n483 = n453 & n482;
  assign n484 = n480 & n483;
  assign n485 = ~n477 & ~n484;
  assign po25 = n338 & ~n485;
  assign n487 = pi11 & ~pi54;
  assign n488 = ~pi10 & ~pi11;
  assign n489 = pi22 & n488;
  assign n490 = n412 & n489;
  assign n491 = n367 & n490;
  assign n492 = n423 & n491;
  assign n493 = ~n487 & ~n492;
  assign po26 = n338 & ~n493;
  assign n495 = pi12 & ~pi54;
  assign n496 = pi18 & n463;
  assign n497 = n413 & n496;
  assign n498 = n461 & n497;
  assign n499 = ~n495 & ~n498;
  assign po27 = n338 & ~n499;
  assign n501 = pi13 & ~pi54;
  assign n502 = ~pi25 & ~pi28;
  assign n503 = pi29 & n502;
  assign n504 = n432 & n503;
  assign n505 = n367 & n504;
  assign n506 = n422 & n434;
  assign n507 = n505 & n506;
  assign n508 = ~n501 & ~n507;
  assign po28 = n338 & ~n508;
  assign n510 = pi14 & ~pi54;
  assign n511 = pi13 & ~pi16;
  assign n512 = n293 & n511;
  assign n513 = n352 & n512;
  assign n514 = n453 & n513;
  assign n515 = n479 & n514;
  assign n516 = ~n510 & ~n515;
  assign po29 = n338 & ~n516;
  assign n518 = pi15 & n387;
  assign n519 = ~pi45 & n389;
  assign n520 = n395 & n397;
  assign n521 = n400 & n519;
  assign n522 = n520 & n521;
  assign n523 = pi15 & ~n522;
  assign n524 = ~pi2 & ~pi20;
  assign n525 = ~pi15 & n389;
  assign n526 = ~n524 & n525;
  assign n527 = n376 & n526;
  assign n528 = n383 & n527;
  assign n529 = ~n523 & ~n528;
  assign n530 = pi82 & ~n529;
  assign n531 = ~pi47 & n377;
  assign n532 = ~pi48 & n519;
  assign n533 = ~pi15 & n531;
  assign n534 = n382 & n533;
  assign n535 = n532 & n534;
  assign n536 = pi82 & ~n535;
  assign n537 = ~pi70 & ~n386;
  assign n538 = ~n536 & n537;
  assign n539 = ~n518 & ~n530;
  assign n540 = ~n538 & n539;
  assign po30 = ~pi129 & ~n540;
  assign n542 = pi16 & ~pi54;
  assign n543 = ~pi5 & pi6;
  assign n544 = ~pi12 & n543;
  assign n545 = n291 & n544;
  assign n546 = n432 & n545;
  assign n547 = n424 & n546;
  assign n548 = ~n542 & ~n547;
  assign po31 = n338 & ~n548;
  assign n550 = pi17 & ~pi54;
  assign n551 = ~pi11 & n310;
  assign n552 = ~pi25 & pi59;
  assign n553 = n340 & n552;
  assign n554 = n445 & n553;
  assign n555 = n354 & n551;
  assign n556 = n554 & n555;
  assign n557 = n295 & n433;
  assign n558 = n556 & n557;
  assign n559 = ~n550 & ~n558;
  assign po32 = n338 & ~n559;
  assign n561 = pi18 & ~pi54;
  assign n562 = pi16 & pi54;
  assign n563 = n294 & n562;
  assign n564 = n366 & n563;
  assign n565 = n462 & n564;
  assign n566 = ~n561 & ~n565;
  assign po33 = n338 & ~n566;
  assign n568 = pi19 & ~pi54;
  assign n569 = pi17 & n551;
  assign n570 = n422 & n569;
  assign n571 = n462 & n570;
  assign n572 = ~n568 & ~n571;
  assign po34 = n338 & ~n572;
  assign n574 = pi20 & n387;
  assign n575 = ~pi43 & n396;
  assign n576 = n376 & n575;
  assign n577 = ~pi38 & n395;
  assign n578 = ~pi50 & n577;
  assign n579 = n576 & n578;
  assign n580 = n389 & n579;
  assign n581 = n388 & n580;
  assign n582 = pi2 & n581;
  assign n583 = ~pi15 & n580;
  assign n584 = pi20 & ~n583;
  assign n585 = ~n582 & ~n584;
  assign n586 = pi82 & ~n585;
  assign n587 = pi82 & ~n581;
  assign n588 = ~pi71 & ~n386;
  assign n589 = ~n587 & n588;
  assign n590 = ~n574 & ~n589;
  assign n591 = ~n586 & n590;
  assign po35 = ~pi129 & ~n591;
  assign n593 = pi21 & ~pi54;
  assign n594 = ~pi4 & pi19;
  assign n595 = ~pi21 & n594;
  assign n596 = n421 & n595;
  assign n597 = n465 & n596;
  assign n598 = n462 & n597;
  assign n599 = ~n593 & ~n598;
  assign po36 = n338 & ~n599;
  assign n601 = pi22 & ~pi54;
  assign n602 = pi5 & ~pi6;
  assign n603 = n346 & n602;
  assign n604 = n292 & n603;
  assign n605 = n463 & n604;
  assign n606 = n480 & n605;
  assign n607 = ~n601 & ~n606;
  assign po37 = n338 & ~n607;
  assign n609 = ~pi23 & pi55;
  assign n610 = pi61 & ~pi129;
  assign po38 = ~n609 & n610;
  assign n612 = pi24 & pi82;
  assign n613 = n579 & n612;
  assign n614 = ~pi2 & ~pi49;
  assign n615 = n388 & n614;
  assign n616 = pi82 & ~n615;
  assign n617 = n386 & ~n616;
  assign n618 = ~n385 & ~n617;
  assign n619 = ~pi24 & ~n618;
  assign n620 = n384 & n615;
  assign n621 = pi82 & ~n620;
  assign n622 = pi63 & ~n386;
  assign n623 = ~n621 & n622;
  assign n624 = ~pi129 & ~n613;
  assign n625 = ~n619 & n624;
  assign po39 = ~n623 & n625;
  assign n627 = pi85 & ~pi116;
  assign n628 = pi25 & n627;
  assign n629 = ~pi96 & ~pi110;
  assign n630 = ~pi85 & ~n629;
  assign n631 = pi100 & ~n627;
  assign n632 = ~n630 & n631;
  assign n633 = ~n628 & ~n632;
  assign n634 = ~pi26 & ~n633;
  assign n635 = pi25 & ~pi116;
  assign n636 = pi26 & n635;
  assign n637 = ~pi95 & ~pi100;
  assign n638 = ~pi97 & n637;
  assign n639 = ~pi110 & ~n638;
  assign n640 = pi25 & ~n639;
  assign n641 = pi26 & pi116;
  assign n642 = ~n640 & ~n641;
  assign n643 = ~pi51 & ~pi52;
  assign n644 = ~pi39 & n643;
  assign n645 = ~n642 & ~n644;
  assign n646 = ~n636 & ~n645;
  assign n647 = ~pi85 & ~n646;
  assign n648 = ~n634 & ~n647;
  assign n649 = ~pi27 & ~n648;
  assign n650 = ~pi39 & ~pi52;
  assign n651 = ~pi51 & n650;
  assign n652 = pi116 & n651;
  assign n653 = ~n635 & ~n652;
  assign n654 = pi27 & ~n653;
  assign n655 = n640 & n644;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~pi26 & ~pi85;
  assign n658 = ~n656 & n657;
  assign n659 = ~n649 & ~n658;
  assign n660 = ~pi53 & ~n659;
  assign n661 = ~pi26 & n635;
  assign n662 = pi53 & ~pi85;
  assign n663 = ~pi27 & n662;
  assign n664 = n661 & n663;
  assign n665 = ~n660 & ~n664;
  assign n666 = ~pi58 & ~n665;
  assign n667 = ~pi27 & ~pi85;
  assign n668 = ~pi53 & pi58;
  assign n669 = n667 & n668;
  assign n670 = n661 & n669;
  assign n671 = ~n666 & ~n670;
  assign po40 = n338 & ~n671;
  assign n673 = ~pi27 & ~pi53;
  assign n674 = ~pi58 & n673;
  assign n675 = ~pi85 & ~n652;
  assign n676 = pi26 & n675;
  assign n677 = n632 & ~n641;
  assign n678 = ~n676 & ~n677;
  assign n679 = n338 & n674;
  assign po41 = ~n678 & n679;
  assign n681 = ~pi53 & ~pi58;
  assign n682 = ~pi26 & n338;
  assign n683 = pi27 & n675;
  assign n684 = pi27 & pi116;
  assign n685 = pi85 & pi116;
  assign n686 = pi95 & ~n627;
  assign n687 = n629 & n686;
  assign n688 = ~n685 & ~n687;
  assign n689 = ~pi100 & ~n684;
  assign n690 = ~n688 & n689;
  assign n691 = ~n683 & ~n690;
  assign n692 = n681 & n682;
  assign po42 = ~n691 & n692;
  assign n694 = ~pi26 & ~pi27;
  assign n695 = ~pi28 & ~pi116;
  assign n696 = pi100 & pi116;
  assign n697 = n694 & ~n695;
  assign n698 = ~n696 & n697;
  assign n699 = pi85 & ~n698;
  assign n700 = ~pi26 & ~n644;
  assign n701 = n684 & n700;
  assign n702 = ~pi27 & n651;
  assign n703 = ~n700 & ~n702;
  assign n704 = ~n639 & ~n703;
  assign n705 = pi26 & ~pi27;
  assign n706 = ~pi26 & pi27;
  assign n707 = ~n705 & ~n706;
  assign n708 = ~pi116 & ~n707;
  assign n709 = ~n704 & ~n708;
  assign n710 = pi28 & ~n709;
  assign n711 = ~pi26 & pi95;
  assign n712 = ~pi100 & n711;
  assign n713 = n629 & n712;
  assign n714 = pi26 & n652;
  assign n715 = ~n713 & ~n714;
  assign n716 = ~pi27 & ~n715;
  assign n717 = ~pi85 & ~n701;
  assign n718 = ~n716 & n717;
  assign n719 = ~n710 & n718;
  assign n720 = ~pi53 & ~n699;
  assign n721 = ~n719 & n720;
  assign n722 = ~pi27 & pi28;
  assign n723 = ~pi116 & n722;
  assign n724 = ~pi26 & n662;
  assign n725 = n723 & n724;
  assign n726 = ~n721 & ~n725;
  assign n727 = ~pi58 & ~n726;
  assign n728 = n657 & n668;
  assign n729 = n723 & n728;
  assign n730 = ~n727 & ~n729;
  assign po43 = n338 & ~n730;
  assign n732 = pi97 & pi116;
  assign n733 = pi29 & ~pi116;
  assign n734 = pi58 & ~n732;
  assign n735 = ~n733 & n734;
  assign n736 = pi29 & pi110;
  assign n737 = ~pi29 & ~pi97;
  assign n738 = pi97 & ~n629;
  assign n739 = n637 & ~n737;
  assign n740 = ~n738 & n739;
  assign n741 = ~pi58 & ~n736;
  assign n742 = ~n740 & n741;
  assign n743 = ~pi53 & ~n735;
  assign n744 = ~n742 & n743;
  assign n745 = pi53 & ~pi58;
  assign n746 = n733 & n745;
  assign n747 = ~n744 & ~n746;
  assign n748 = ~pi27 & ~n747;
  assign n749 = pi27 & n681;
  assign n750 = n733 & n749;
  assign n751 = ~n748 & ~n750;
  assign n752 = ~pi85 & ~n751;
  assign n753 = pi85 & n733;
  assign n754 = n674 & n753;
  assign n755 = ~n752 & ~n754;
  assign n756 = ~pi26 & ~n755;
  assign n757 = ~pi85 & n681;
  assign n758 = n705 & n757;
  assign n759 = n733 & n758;
  assign n760 = ~n756 & ~n759;
  assign po44 = n338 & ~n760;
  assign n762 = ~pi88 & pi106;
  assign n763 = pi30 & ~pi109;
  assign n764 = pi60 & pi109;
  assign n765 = ~pi106 & ~n763;
  assign n766 = ~n764 & n765;
  assign n767 = ~pi129 & ~n762;
  assign po45 = ~n766 & n767;
  assign n769 = ~pi89 & pi106;
  assign n770 = pi31 & ~pi109;
  assign n771 = pi30 & pi109;
  assign n772 = ~pi106 & ~n770;
  assign n773 = ~n771 & n772;
  assign n774 = ~pi129 & ~n769;
  assign po46 = ~n773 & n774;
  assign n776 = ~pi99 & pi106;
  assign n777 = pi32 & ~pi109;
  assign n778 = pi31 & pi109;
  assign n779 = ~pi106 & ~n777;
  assign n780 = ~n778 & n779;
  assign n781 = ~pi129 & ~n776;
  assign po47 = ~n780 & n781;
  assign n783 = ~pi90 & pi106;
  assign n784 = pi33 & ~pi109;
  assign n785 = pi32 & pi109;
  assign n786 = ~pi106 & ~n784;
  assign n787 = ~n785 & n786;
  assign n788 = ~pi129 & ~n783;
  assign po48 = ~n787 & n788;
  assign n790 = ~pi91 & pi106;
  assign n791 = pi34 & ~pi109;
  assign n792 = pi33 & pi109;
  assign n793 = ~pi106 & ~n791;
  assign n794 = ~n792 & n793;
  assign n795 = ~pi129 & ~n790;
  assign po49 = ~n794 & n795;
  assign n797 = ~pi92 & pi106;
  assign n798 = pi35 & ~pi109;
  assign n799 = pi34 & pi109;
  assign n800 = ~pi106 & ~n798;
  assign n801 = ~n799 & n800;
  assign n802 = ~pi129 & ~n797;
  assign po50 = ~n801 & n802;
  assign n804 = ~pi98 & pi106;
  assign n805 = pi36 & ~pi109;
  assign n806 = pi35 & pi109;
  assign n807 = ~pi106 & ~n805;
  assign n808 = ~n806 & n807;
  assign n809 = ~pi129 & ~n804;
  assign po51 = ~n808 & n809;
  assign n811 = ~pi93 & pi106;
  assign n812 = pi37 & ~pi109;
  assign n813 = pi36 & pi109;
  assign n814 = ~pi106 & ~n812;
  assign n815 = ~n813 & n814;
  assign n816 = ~pi129 & ~n811;
  assign po52 = ~n815 & n816;
  assign n818 = ~pi40 & ~pi42;
  assign n819 = ~pi44 & pi82;
  assign n820 = n818 & n819;
  assign n821 = pi38 & n820;
  assign n822 = ~pi2 & n388;
  assign n823 = n532 & n822;
  assign n824 = n396 & n399;
  assign n825 = n823 & n824;
  assign n826 = ~pi50 & n395;
  assign n827 = n825 & n826;
  assign n828 = pi82 & ~n827;
  assign n829 = pi74 & ~n386;
  assign n830 = ~n828 & n829;
  assign n831 = pi82 & ~n395;
  assign n832 = n519 & n822;
  assign n833 = n375 & n575;
  assign n834 = ~pi50 & n833;
  assign n835 = n832 & n834;
  assign n836 = pi82 & ~n835;
  assign n837 = n386 & ~n836;
  assign n838 = ~n831 & ~n837;
  assign n839 = ~pi38 & ~n838;
  assign n840 = ~pi129 & ~n821;
  assign n841 = ~n830 & n840;
  assign po53 = ~n839 & n841;
  assign n843 = pi109 & n643;
  assign n844 = pi39 & ~n843;
  assign n845 = ~pi51 & pi109;
  assign n846 = n650 & n845;
  assign n847 = ~pi106 & ~n846;
  assign n848 = ~n844 & n847;
  assign po54 = ~pi129 & ~n848;
  assign n850 = ~pi42 & n819;
  assign n851 = pi40 & n850;
  assign n852 = n379 & n825;
  assign n853 = n378 & n852;
  assign n854 = pi82 & ~n853;
  assign n855 = pi73 & ~n386;
  assign n856 = ~n854 & n855;
  assign n857 = pi82 & ~n378;
  assign n858 = pi82 & ~n403;
  assign n859 = n386 & ~n858;
  assign n860 = ~n857 & ~n859;
  assign n861 = ~pi40 & ~n860;
  assign n862 = ~pi129 & ~n851;
  assign n863 = ~n856 & n862;
  assign po55 = ~n861 & n863;
  assign n865 = pi82 & ~n382;
  assign n866 = pi82 & ~n402;
  assign n867 = n386 & ~n866;
  assign n868 = ~n865 & ~n867;
  assign n869 = ~pi41 & ~n868;
  assign n870 = pi41 & n381;
  assign n871 = n850 & n870;
  assign n872 = ~pi46 & n399;
  assign n873 = n578 & n872;
  assign n874 = n823 & n873;
  assign n875 = pi82 & ~n874;
  assign n876 = pi76 & ~n386;
  assign n877 = ~n875 & n876;
  assign n878 = ~pi129 & ~n871;
  assign n879 = ~n869 & n878;
  assign po56 = ~n877 & n879;
  assign n881 = pi44 & pi82;
  assign n882 = n531 & n823;
  assign n883 = n381 & n882;
  assign n884 = pi82 & ~n883;
  assign n885 = n386 & ~n884;
  assign n886 = ~n881 & ~n885;
  assign n887 = ~pi42 & ~n886;
  assign n888 = pi42 & n819;
  assign n889 = ~pi40 & ~pi44;
  assign n890 = n852 & n889;
  assign n891 = pi82 & ~n890;
  assign n892 = pi72 & ~n386;
  assign n893 = ~n891 & n892;
  assign n894 = ~pi129 & ~n888;
  assign n895 = ~n893 & n894;
  assign po57 = ~n887 & n895;
  assign n897 = n397 & n818;
  assign n898 = pi43 & n819;
  assign n899 = n897 & n898;
  assign n900 = pi82 & ~n520;
  assign n901 = ~pi2 & n375;
  assign n902 = n398 & n901;
  assign n903 = pi82 & ~n902;
  assign n904 = n386 & ~n903;
  assign n905 = ~n900 & ~n904;
  assign n906 = ~pi43 & ~n905;
  assign n907 = ~pi47 & n520;
  assign n908 = n823 & n907;
  assign n909 = pi82 & ~n908;
  assign n910 = pi77 & ~n386;
  assign n911 = ~n909 & n910;
  assign n912 = ~pi129 & ~n899;
  assign n913 = ~n911 & n912;
  assign po58 = ~n906 & n913;
  assign n915 = ~pi42 & n883;
  assign n916 = pi82 & ~n915;
  assign n917 = ~pi67 & ~n386;
  assign n918 = pi44 & n386;
  assign n919 = ~n917 & ~n918;
  assign n920 = ~n916 & n919;
  assign n921 = ~pi129 & ~n881;
  assign po59 = ~n920 & n921;
  assign n923 = pi45 & pi82;
  assign n924 = n577 & n923;
  assign n925 = n834 & n924;
  assign n926 = ~pi2 & n390;
  assign n927 = pi82 & ~n926;
  assign n928 = n386 & ~n927;
  assign n929 = n578 & n833;
  assign n930 = pi82 & ~n929;
  assign n931 = ~n928 & ~n930;
  assign n932 = ~pi45 & ~n931;
  assign n933 = n390 & n901;
  assign n934 = n383 & n933;
  assign n935 = pi82 & ~n934;
  assign n936 = pi68 & ~n386;
  assign n937 = ~n935 & n936;
  assign n938 = ~pi129 & ~n925;
  assign n939 = ~n937 & n938;
  assign po60 = ~n932 & n939;
  assign n941 = pi82 & ~n578;
  assign n942 = pi82 & ~n882;
  assign n943 = n386 & ~n942;
  assign n944 = ~n941 & ~n943;
  assign n945 = ~pi46 & ~n944;
  assign n946 = pi46 & pi82;
  assign n947 = n578 & n946;
  assign n948 = n578 & n882;
  assign n949 = pi82 & ~n948;
  assign n950 = pi75 & ~n386;
  assign n951 = ~n949 & n950;
  assign n952 = ~pi129 & ~n947;
  assign n953 = ~n951 & n952;
  assign po61 = ~n945 & n953;
  assign n955 = pi47 & n379;
  assign n956 = n575 & n955;
  assign n957 = n820 & n956;
  assign n958 = pi82 & ~n383;
  assign n959 = pi82 & ~n823;
  assign n960 = n386 & ~n959;
  assign n961 = ~n958 & ~n960;
  assign n962 = ~pi47 & ~n961;
  assign n963 = n383 & n823;
  assign n964 = pi82 & ~n963;
  assign n965 = pi64 & ~n386;
  assign n966 = ~n964 & n965;
  assign n967 = ~pi129 & ~n957;
  assign n968 = ~n966 & n967;
  assign po62 = ~n962 & n968;
  assign n970 = pi48 & n399;
  assign n971 = n819 & n970;
  assign n972 = n897 & n971;
  assign n973 = pi82 & ~n832;
  assign n974 = n386 & ~n973;
  assign n975 = n578 & n824;
  assign n976 = pi82 & ~n975;
  assign n977 = ~n974 & ~n976;
  assign n978 = ~pi48 & ~n977;
  assign n979 = n382 & n531;
  assign n980 = n832 & n979;
  assign n981 = pi82 & ~n980;
  assign n982 = pi62 & ~n386;
  assign n983 = ~n981 & n982;
  assign n984 = ~pi129 & ~n972;
  assign n985 = ~n983 & n984;
  assign po63 = ~n978 & n985;
  assign n987 = ~pi24 & n379;
  assign n988 = n395 & n987;
  assign n989 = n576 & n988;
  assign n990 = pi49 & ~n989;
  assign n991 = n389 & ~n822;
  assign n992 = n579 & n991;
  assign n993 = ~n990 & ~n992;
  assign n994 = pi82 & ~n993;
  assign n995 = pi49 & n387;
  assign n996 = pi82 & ~n580;
  assign n997 = ~pi69 & ~n386;
  assign n998 = ~n996 & n997;
  assign n999 = ~n994 & ~n995;
  assign n1000 = ~n998 & n999;
  assign po64 = ~pi129 & ~n1000;
  assign n1002 = pi50 & pi82;
  assign n1003 = n577 & n1002;
  assign n1004 = pi82 & ~n577;
  assign n1005 = n575 & n902;
  assign n1006 = pi82 & ~n1005;
  assign n1007 = n386 & ~n1006;
  assign n1008 = ~n1004 & ~n1007;
  assign n1009 = ~pi50 & ~n1008;
  assign n1010 = n577 & n825;
  assign n1011 = pi82 & ~n1010;
  assign n1012 = pi66 & ~n386;
  assign n1013 = ~n1011 & n1012;
  assign n1014 = ~pi129 & ~n1003;
  assign n1015 = ~n1013 & n1014;
  assign po65 = ~n1009 & n1015;
  assign n1017 = pi51 & ~pi109;
  assign n1018 = ~pi106 & ~n845;
  assign n1019 = ~n1017 & n1018;
  assign po66 = ~pi129 & ~n1019;
  assign n1021 = pi52 & ~n845;
  assign n1022 = ~pi106 & ~n843;
  assign n1023 = ~n1021 & n1022;
  assign po67 = ~pi129 & ~n1023;
  assign n1025 = ~pi116 & n745;
  assign n1026 = pi58 & pi116;
  assign n1027 = ~pi58 & n629;
  assign n1028 = n637 & n1027;
  assign n1029 = ~n1026 & ~n1028;
  assign n1030 = ~pi53 & pi97;
  assign n1031 = ~n1029 & n1030;
  assign n1032 = ~n1025 & ~n1031;
  assign n1033 = n667 & n682;
  assign po68 = ~n1032 & n1033;
  assign n1035 = ~pi45 & n934;
  assign n1036 = pi82 & ~n1035;
  assign n1037 = ~n386 & ~n1036;
  assign po69 = pi129 | n1037;
  assign po129 = pi123 | pi129;
  assign n1040 = pi114 & ~pi122;
  assign po70 = ~po129 & n1040;
  assign n1042 = ~pi26 & pi58;
  assign n1043 = ~pi58 & n641;
  assign n1044 = ~n1042 & ~n1043;
  assign n1045 = pi94 & ~n1044;
  assign n1046 = pi58 & ~pi116;
  assign n1047 = pi37 & ~pi116;
  assign n1048 = ~n1042 & ~n1047;
  assign n1049 = ~n1046 & ~n1048;
  assign n1050 = ~n1045 & ~n1049;
  assign n1051 = ~pi53 & ~n1050;
  assign n1052 = ~pi26 & pi37;
  assign n1053 = ~pi58 & n1052;
  assign n1054 = ~n1051 & ~n1053;
  assign n1055 = ~pi85 & ~n1054;
  assign n1056 = n681 & n1052;
  assign n1057 = ~n1055 & ~n1056;
  assign n1058 = ~pi27 & ~n1057;
  assign n1059 = n757 & n1052;
  assign n1060 = ~n1058 & ~n1059;
  assign po71 = n338 & ~n1060;
  assign n1062 = ~pi26 & ~pi53;
  assign n1063 = ~pi85 & n1062;
  assign n1064 = ~pi116 & n1063;
  assign n1065 = pi26 & pi53;
  assign n1066 = pi85 & ~n1062;
  assign n1067 = ~pi58 & ~n1065;
  assign n1068 = ~n1066 & n1067;
  assign n1069 = ~n1064 & ~n1068;
  assign n1070 = pi57 & ~n1069;
  assign n1071 = pi60 & n1026;
  assign n1072 = n1063 & n1071;
  assign n1073 = ~n1070 & ~n1072;
  assign n1074 = ~pi27 & ~n1073;
  assign n1075 = pi57 & ~pi58;
  assign n1076 = n1063 & n1075;
  assign n1077 = ~n1074 & ~n1076;
  assign po72 = n338 & ~n1077;
  assign n1079 = n694 & n1046;
  assign n1080 = ~pi58 & ~n707;
  assign n1081 = n652 & n1080;
  assign n1082 = ~n1079 & ~n1081;
  assign n1083 = ~pi53 & ~pi85;
  assign n1084 = n338 & n1083;
  assign po73 = ~n1082 & n1084;
  assign n1086 = ~n668 & ~n745;
  assign n1087 = ~pi116 & ~n1086;
  assign n1088 = ~n639 & n681;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = pi59 & ~n1089;
  assign n1091 = pi96 & n681;
  assign n1092 = n639 & n1091;
  assign n1093 = ~n1090 & ~n1092;
  assign n1094 = ~pi85 & ~n1093;
  assign n1095 = pi59 & ~pi116;
  assign n1096 = pi85 & n681;
  assign n1097 = n1095 & n1096;
  assign n1098 = ~n1094 & ~n1097;
  assign n1099 = ~pi27 & ~n1098;
  assign n1100 = pi27 & n1095;
  assign n1101 = n757 & n1100;
  assign n1102 = ~n1099 & ~n1101;
  assign n1103 = ~pi26 & ~n1102;
  assign n1104 = n758 & n1095;
  assign n1105 = ~n1103 & ~n1104;
  assign po74 = n338 & ~n1105;
  assign n1107 = ~pi117 & ~pi122;
  assign n1108 = pi60 & ~n1107;
  assign n1109 = pi123 & n1107;
  assign po75 = n1108 | n1109;
  assign n1111 = ~pi114 & ~pi122;
  assign n1112 = pi123 & ~pi129;
  assign po76 = n1111 & n1112;
  assign n1114 = pi136 & ~pi137;
  assign n1115 = pi131 & pi132;
  assign n1116 = pi133 & n1115;
  assign n1117 = ~pi138 & n1116;
  assign n1118 = n1114 & n1117;
  assign n1119 = ~pi62 & ~n1118;
  assign n1120 = pi140 & n1118;
  assign n1121 = ~pi129 & ~n1119;
  assign po77 = n1120 | ~n1121;
  assign n1123 = ~pi63 & ~n1118;
  assign n1124 = pi142 & n1118;
  assign n1125 = ~pi129 & ~n1123;
  assign po78 = n1124 | ~n1125;
  assign n1127 = ~pi64 & ~n1118;
  assign n1128 = pi139 & n1118;
  assign n1129 = ~pi129 & ~n1127;
  assign po79 = n1128 | ~n1129;
  assign n1131 = ~pi65 & ~n1118;
  assign n1132 = pi146 & n1118;
  assign n1133 = ~pi129 & ~n1131;
  assign po80 = n1132 | ~n1133;
  assign n1135 = ~pi136 & ~pi137;
  assign n1136 = n1117 & n1135;
  assign n1137 = ~pi66 & ~n1136;
  assign n1138 = pi143 & n1136;
  assign n1139 = ~pi129 & ~n1137;
  assign po81 = n1138 | ~n1139;
  assign n1141 = ~pi67 & ~n1136;
  assign n1142 = pi139 & n1136;
  assign n1143 = ~pi129 & ~n1141;
  assign po82 = n1142 | ~n1143;
  assign n1145 = ~pi68 & ~n1118;
  assign n1146 = pi141 & n1118;
  assign n1147 = ~pi129 & ~n1145;
  assign po83 = n1146 | ~n1147;
  assign n1149 = ~pi69 & ~n1118;
  assign n1150 = pi143 & n1118;
  assign n1151 = ~pi129 & ~n1149;
  assign po84 = n1150 | ~n1151;
  assign n1153 = ~pi70 & ~n1118;
  assign n1154 = pi144 & n1118;
  assign n1155 = ~pi129 & ~n1153;
  assign po85 = n1154 | ~n1155;
  assign n1157 = ~pi71 & ~n1118;
  assign n1158 = pi145 & n1118;
  assign n1159 = ~pi129 & ~n1157;
  assign po86 = n1158 | ~n1159;
  assign n1161 = ~pi72 & ~n1136;
  assign n1162 = pi140 & n1136;
  assign n1163 = ~pi129 & ~n1161;
  assign po87 = n1162 | ~n1163;
  assign n1165 = ~pi73 & ~n1136;
  assign n1166 = pi141 & n1136;
  assign n1167 = ~pi129 & ~n1165;
  assign po88 = n1166 | ~n1167;
  assign n1169 = ~pi74 & ~n1136;
  assign n1170 = pi142 & n1136;
  assign n1171 = ~pi129 & ~n1169;
  assign po89 = n1170 | ~n1171;
  assign n1173 = ~pi75 & ~n1136;
  assign n1174 = pi144 & n1136;
  assign n1175 = ~pi129 & ~n1173;
  assign po90 = n1174 | ~n1175;
  assign n1177 = ~pi76 & ~n1136;
  assign n1178 = pi145 & n1136;
  assign n1179 = ~pi129 & ~n1177;
  assign po91 = n1178 | ~n1179;
  assign n1181 = ~pi77 & ~n1136;
  assign n1182 = pi146 & n1136;
  assign n1183 = ~pi129 & ~n1181;
  assign po92 = n1182 | ~n1183;
  assign n1185 = ~pi136 & pi137;
  assign n1186 = n1117 & n1185;
  assign n1187 = ~pi78 & ~n1186;
  assign n1188 = ~pi142 & n1186;
  assign n1189 = ~pi129 & ~n1187;
  assign po93 = ~n1188 & n1189;
  assign n1191 = ~pi79 & ~n1186;
  assign n1192 = ~pi143 & n1186;
  assign n1193 = ~pi129 & ~n1191;
  assign po94 = ~n1192 & n1193;
  assign n1195 = ~pi80 & ~n1186;
  assign n1196 = ~pi144 & n1186;
  assign n1197 = ~pi129 & ~n1195;
  assign po95 = ~n1196 & n1197;
  assign n1199 = ~pi81 & ~n1186;
  assign n1200 = ~pi145 & n1186;
  assign n1201 = ~pi129 & ~n1199;
  assign po96 = ~n1200 & n1201;
  assign n1203 = ~pi82 & ~n1186;
  assign n1204 = ~pi146 & n1186;
  assign n1205 = ~pi129 & ~n1203;
  assign po97 = ~n1204 & n1205;
  assign n1207 = ~pi89 & pi138;
  assign n1208 = pi62 & ~pi138;
  assign n1209 = pi136 & ~n1207;
  assign n1210 = ~n1208 & n1209;
  assign n1211 = ~pi119 & pi138;
  assign n1212 = pi72 & ~pi138;
  assign n1213 = ~pi136 & ~n1211;
  assign n1214 = ~n1212 & n1213;
  assign n1215 = ~n1210 & ~n1214;
  assign n1216 = ~pi137 & ~n1215;
  assign n1217 = pi136 & ~pi138;
  assign n1218 = pi31 & n1217;
  assign n1219 = ~pi87 & ~pi138;
  assign n1220 = pi115 & pi138;
  assign n1221 = ~pi136 & ~n1219;
  assign n1222 = ~n1220 & n1221;
  assign n1223 = ~n1218 & ~n1222;
  assign n1224 = pi137 & ~n1223;
  assign po98 = n1216 | n1224;
  assign n1226 = ~pi84 & ~n1186;
  assign n1227 = ~pi141 & n1186;
  assign n1228 = ~pi129 & ~n1226;
  assign po99 = ~n1227 & n1228;
  assign n1230 = ~pi85 & n639;
  assign n1231 = pi96 & n1230;
  assign n1232 = ~n627 & ~n1231;
  assign n1233 = n674 & n682;
  assign po100 = ~n1232 & n1233;
  assign n1235 = ~pi86 & ~n1186;
  assign n1236 = ~pi139 & n1186;
  assign n1237 = ~pi129 & ~n1235;
  assign po101 = ~n1236 & n1237;
  assign n1239 = ~pi87 & ~n1186;
  assign n1240 = ~pi140 & n1186;
  assign n1241 = ~pi129 & ~n1239;
  assign po102 = ~n1240 & n1241;
  assign n1243 = pi137 & n1217;
  assign n1244 = n1116 & n1243;
  assign n1245 = ~pi88 & ~n1244;
  assign n1246 = ~pi139 & n1244;
  assign n1247 = ~pi129 & ~n1245;
  assign po103 = ~n1246 & n1247;
  assign n1249 = ~pi89 & ~n1244;
  assign n1250 = ~pi140 & n1244;
  assign n1251 = ~pi129 & ~n1249;
  assign po104 = ~n1250 & n1251;
  assign n1253 = ~pi90 & ~n1244;
  assign n1254 = ~pi142 & n1244;
  assign n1255 = ~pi129 & ~n1253;
  assign po105 = ~n1254 & n1255;
  assign n1257 = ~pi91 & ~n1244;
  assign n1258 = ~pi143 & n1244;
  assign n1259 = ~pi129 & ~n1257;
  assign po106 = ~n1258 & n1259;
  assign n1261 = ~pi92 & ~n1244;
  assign n1262 = ~pi144 & n1244;
  assign n1263 = ~pi129 & ~n1261;
  assign po107 = ~n1262 & n1263;
  assign n1265 = ~pi93 & ~n1244;
  assign n1266 = ~pi146 & n1244;
  assign n1267 = ~pi129 & ~n1265;
  assign po108 = ~n1266 & n1267;
  assign n1269 = pi82 & pi138;
  assign n1270 = n1135 & n1269;
  assign n1271 = n1116 & n1270;
  assign n1272 = ~pi94 & ~n1271;
  assign n1273 = ~pi142 & n1271;
  assign n1274 = ~pi129 & ~n1272;
  assign po109 = ~n1273 & n1274;
  assign n1276 = ~pi3 & ~pi110;
  assign n1277 = ~n1116 & ~n1276;
  assign n1278 = ~n1271 & ~n1277;
  assign n1279 = pi95 & n1278;
  assign n1280 = pi143 & n1271;
  assign n1281 = ~n1279 & ~n1280;
  assign po110 = ~pi129 & ~n1281;
  assign n1283 = pi96 & n1278;
  assign n1284 = pi146 & n1271;
  assign n1285 = ~n1283 & ~n1284;
  assign po111 = ~pi129 & ~n1285;
  assign n1287 = pi97 & n1278;
  assign n1288 = pi145 & n1271;
  assign n1289 = ~n1287 & ~n1288;
  assign po112 = ~pi129 & ~n1289;
  assign n1291 = ~pi98 & ~n1244;
  assign n1292 = ~pi145 & n1244;
  assign n1293 = ~pi129 & ~n1291;
  assign po113 = ~n1292 & n1293;
  assign n1295 = ~pi99 & ~n1244;
  assign n1296 = ~pi141 & n1244;
  assign n1297 = ~pi129 & ~n1295;
  assign po114 = ~n1296 & n1297;
  assign n1299 = pi100 & n1278;
  assign n1300 = pi144 & n1271;
  assign n1301 = ~n1299 & ~n1300;
  assign po115 = ~pi129 & ~n1301;
  assign n1303 = ~pi124 & pi138;
  assign n1304 = pi77 & ~pi138;
  assign n1305 = ~pi136 & ~n1303;
  assign n1306 = ~n1304 & n1305;
  assign n1307 = ~pi93 & pi138;
  assign n1308 = pi65 & ~pi138;
  assign n1309 = pi136 & ~n1307;
  assign n1310 = ~n1308 & n1309;
  assign n1311 = ~n1306 & ~n1310;
  assign n1312 = ~pi137 & ~n1311;
  assign n1313 = pi37 & n1217;
  assign n1314 = ~pi82 & ~pi138;
  assign n1315 = ~pi96 & pi138;
  assign n1316 = ~pi136 & ~n1314;
  assign n1317 = ~n1315 & n1316;
  assign n1318 = ~n1313 & ~n1317;
  assign n1319 = pi137 & ~n1318;
  assign po116 = n1312 | n1319;
  assign n1321 = pi91 & n1114;
  assign n1322 = pi95 & n1185;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = pi138 & ~n1323;
  assign n1325 = ~pi79 & ~pi136;
  assign n1326 = ~pi34 & pi136;
  assign n1327 = pi137 & ~n1325;
  assign n1328 = ~n1326 & n1327;
  assign n1329 = pi66 & ~pi136;
  assign n1330 = pi69 & pi136;
  assign n1331 = ~pi137 & ~n1329;
  assign n1332 = ~n1330 & n1331;
  assign n1333 = ~n1328 & ~n1332;
  assign n1334 = ~pi138 & ~n1333;
  assign po117 = n1324 | n1334;
  assign n1336 = pi90 & n1114;
  assign n1337 = pi94 & n1185;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = pi138 & ~n1338;
  assign n1340 = ~pi78 & ~pi136;
  assign n1341 = ~pi33 & pi136;
  assign n1342 = pi137 & ~n1340;
  assign n1343 = ~n1341 & n1342;
  assign n1344 = pi74 & ~pi136;
  assign n1345 = pi63 & pi136;
  assign n1346 = ~pi137 & ~n1344;
  assign n1347 = ~n1345 & n1346;
  assign n1348 = ~n1343 & ~n1347;
  assign n1349 = ~pi138 & ~n1348;
  assign po118 = n1339 | n1349;
  assign n1351 = pi99 & n1114;
  assign n1352 = ~pi112 & n1185;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = pi138 & ~n1353;
  assign n1355 = pi73 & ~pi136;
  assign n1356 = pi68 & pi136;
  assign n1357 = ~pi137 & ~n1355;
  assign n1358 = ~n1356 & n1357;
  assign n1359 = ~pi84 & ~pi136;
  assign n1360 = ~pi32 & pi136;
  assign n1361 = pi137 & ~n1359;
  assign n1362 = ~n1360 & n1361;
  assign n1363 = ~n1358 & ~n1362;
  assign n1364 = ~pi138 & ~n1363;
  assign po119 = n1354 | n1364;
  assign n1366 = ~pi92 & pi138;
  assign n1367 = pi70 & ~pi138;
  assign n1368 = pi136 & ~n1366;
  assign n1369 = ~n1367 & n1368;
  assign n1370 = ~pi125 & pi138;
  assign n1371 = pi75 & ~pi138;
  assign n1372 = ~pi136 & ~n1370;
  assign n1373 = ~n1371 & n1372;
  assign n1374 = ~n1369 & ~n1373;
  assign n1375 = ~pi137 & ~n1374;
  assign n1376 = pi35 & n1217;
  assign n1377 = ~pi80 & ~pi138;
  assign n1378 = ~pi100 & pi138;
  assign n1379 = ~pi136 & ~n1377;
  assign n1380 = ~n1378 & n1379;
  assign n1381 = ~n1376 & ~n1380;
  assign n1382 = pi137 & ~n1381;
  assign po120 = n1375 | n1382;
  assign n1384 = ~pi26 & n674;
  assign n1385 = n1230 & n1384;
  assign n1386 = ~n685 & ~n1385;
  assign po121 = n338 & ~n1386;
  assign n1388 = ~pi98 & pi138;
  assign n1389 = pi71 & ~pi138;
  assign n1390 = pi136 & ~n1388;
  assign n1391 = ~n1389 & n1390;
  assign n1392 = ~pi23 & pi138;
  assign n1393 = pi76 & ~pi138;
  assign n1394 = ~pi136 & ~n1392;
  assign n1395 = ~n1393 & n1394;
  assign n1396 = ~n1391 & ~n1395;
  assign n1397 = ~pi137 & ~n1396;
  assign n1398 = pi36 & n1217;
  assign n1399 = ~pi81 & ~pi138;
  assign n1400 = ~pi97 & pi138;
  assign n1401 = ~pi136 & ~n1399;
  assign n1402 = ~n1400 & n1401;
  assign n1403 = ~n1398 & ~n1402;
  assign n1404 = pi137 & ~n1403;
  assign po122 = n1397 | n1404;
  assign n1406 = ~pi88 & pi138;
  assign n1407 = pi64 & ~pi138;
  assign n1408 = pi136 & ~n1406;
  assign n1409 = ~n1407 & n1408;
  assign n1410 = ~pi120 & pi138;
  assign n1411 = pi67 & ~pi138;
  assign n1412 = ~pi136 & ~n1410;
  assign n1413 = ~n1411 & n1412;
  assign n1414 = ~n1409 & ~n1413;
  assign n1415 = ~pi137 & ~n1414;
  assign n1416 = pi30 & n1217;
  assign n1417 = ~pi86 & ~pi138;
  assign n1418 = ~pi111 & pi138;
  assign n1419 = ~pi136 & ~n1417;
  assign n1420 = ~n1418 & n1419;
  assign n1421 = ~n1416 & ~n1420;
  assign n1422 = pi137 & ~n1421;
  assign po123 = n1415 | n1422;
  assign n1424 = ~pi26 & n644;
  assign n1425 = pi116 & n338;
  assign n1426 = ~n707 & n1425;
  assign po124 = ~n1424 & n1426;
  assign n1428 = ~pi97 & n668;
  assign n1429 = ~n745 & ~n1428;
  assign po125 = n1425 & ~n1429;
  assign n1431 = ~pi111 & ~n1270;
  assign n1432 = ~pi129 & n1116;
  assign n1433 = ~pi139 & n1270;
  assign n1434 = ~n1431 & n1432;
  assign po126 = ~n1433 & n1434;
  assign n1436 = ~pi141 & n1270;
  assign n1437 = pi112 & ~n1270;
  assign n1438 = n1432 & ~n1436;
  assign po127 = ~n1437 & n1438;
  assign n1440 = ~pi54 & pi113;
  assign n1441 = ~pi11 & ~pi22;
  assign n1442 = pi54 & n1441;
  assign n1443 = n338 & ~n1440;
  assign po128 = ~n1442 & n1443;
  assign n1445 = ~pi140 & n1270;
  assign n1446 = pi115 & ~n1270;
  assign n1447 = n1432 & ~n1445;
  assign po130 = ~n1446 & n1447;
  assign n1449 = ~pi4 & ~pi7;
  assign n1450 = ~pi9 & ~pi12;
  assign n1451 = n1449 & n1450;
  assign n1452 = pi54 & n338;
  assign po131 = ~n1451 & n1452;
  assign po132 = ~pi122 | pi129;
  assign n1455 = ~pi54 & pi118;
  assign n1456 = pi54 & ~pi59;
  assign n1457 = n503 & n1456;
  assign n1458 = ~n1455 & ~n1457;
  assign po133 = ~pi129 & ~n1458;
  assign po134 = ~pi129 & ~n637;
  assign n1461 = ~pi120 & n1276;
  assign n1462 = ~pi111 & ~pi129;
  assign po135 = ~n1461 & n1462;
  assign n1464 = pi81 & pi120;
  assign po136 = ~pi129 & n1464;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi57 & ~pi129;
  assign n1469 = ~pi96 & pi125;
  assign n1470 = ~pi3 & ~n1469;
  assign po140 = ~pi129 & ~n1470;
  assign n1472 = ~pi126 & pi132;
  assign po141 = pi133 & n1472;
  assign po12 = 1'b1;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
endmodule
