module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 ;
  wire n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102,
    n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396,
    n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426,
    n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894,
    n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924,
    n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170,
    n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182,
    n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200,
    n3201, n3202, n3203, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212,
    n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242,
    n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272,
    n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302,
    n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332,
    n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362,
    n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3390, n3391, n3392,
    n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416,
    n3417, n3418, n3419, n3420, n3421, n3422,
    n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3439, n3440,
    n3441, n3442, n3443, n3444, n3445, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476,
    n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722,
    n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782,
    n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052,
    n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292,
    n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334,
    n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346,
    n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382,
    n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412,
    n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430,
    n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442,
    n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466,
    n4467, n4468, n4469, n4470, n4471, n4472,
    n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496,
    n4497, n4498, n4499, n4500, n4501, n4502,
    n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526,
    n4527, n4528, n4529, n4530, n4531, n4532,
    n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562,
    n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586,
    n4587, n4588, n4589, n4590, n4591, n4592,
    n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622,
    n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700,
    n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708, n4709, n4710, n4711, n4712,
    n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5040, n5041, n5042,
    n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072,
    n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372,
    n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390,
    n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402,
    n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414,
    n5415, n5416, n5417, n5418, n5419, n5420,
    n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5436, n5437, n5438,
    n5439, n5440, n5441, n5442, n5443, n5444,
    n5445, n5446, n5447, n5448, n5449, n5450,
    n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5460, n5461, n5462,
    n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5470, n5471, n5472, n5473, n5474,
    n5475, n5476, n5477, n5478, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528,
    n5529, n5530, n5531, n5532, n5533, n5534,
    n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5542, n5543, n5544, n5545, n5546,
    n5547, n5548, n5549, n5550, n5551, n5552,
    n5553, n5554, n5555, n5556, n5557, n5558,
    n5559, n5560, n5561, n5562, n5563, n5564,
    n5565, n5566, n5567, n5568, n5569, n5570,
    n5571, n5572, n5573, n5574, n5575, n5576,
    n5577, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588,
    n5589, n5590, n5591, n5592, n5593, n5594,
    n5595, n5596, n5597, n5598, n5599, n5600,
    n5601, n5602, n5603, n5604, n5605, n5606,
    n5607, n5608, n5609, n5610, n5611, n5612,
    n5613, n5614, n5615, n5616, n5617, n5618,
    n5619, n5620, n5621, n5622, n5623, n5624,
    n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636,
    n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648,
    n5649, n5650, n5651, n5652, n5653, n5654,
    n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678,
    n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708,
    n5709, n5710, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5718, n5719, n5720,
    n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732,
    n5733, n5734, n5735, n5736, n5737, n5738,
    n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750,
    n5751, n5752, n5753, n5754, n5755, n5756,
    n5757, n5758, n5759, n5760, n5761, n5762,
    n5763, n5764, n5765, n5766, n5767, n5768,
    n5769, n5770, n5771, n5772, n5773, n5774,
    n5775, n5776, n5777, n5778, n5779, n5780,
    n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792,
    n5793, n5794, n5795, n5796, n5797, n5798,
    n5799, n5800, n5801, n5802, n5803, n5804,
    n5805, n5806, n5807, n5808, n5809, n5810,
    n5811, n5812, n5813, n5814, n5815, n5816,
    n5817, n5818, n5819, n5820, n5821, n5822,
    n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5834,
    n5835, n5836, n5837, n5838, n5839, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846,
    n5847, n5848, n5849, n5850, n5851, n5852,
    n5853, n5854, n5855, n5856, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864,
    n5865, n5866, n5867, n5868, n5869, n5870,
    n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882,
    n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894,
    n5895, n5896, n5897, n5898, n5899, n5900,
    n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912,
    n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924,
    n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954,
    n5955, n5956, n5957, n5958, n5959, n5960,
    n5961, n5962, n5963, n5964, n5965, n5966,
    n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5986, n5987, n5988, n5989, n5990,
    n5991, n5992, n5993, n5994, n5995, n5996,
    n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020,
    n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050,
    n6051, n6052, n6053, n6054, n6055, n6056,
    n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074,
    n6075, n6076, n6077, n6078, n6079, n6080,
    n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110,
    n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122,
    n6123, n6124, n6125, n6126, n6127, n6128,
    n6129, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140,
    n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236,
    n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266,
    n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278,
    n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296,
    n6297, n6298, n6299, n6300, n6301, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326,
    n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362,
    n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386,
    n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398,
    n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416,
    n6417, n6418, n6419, n6420, n6421, n6422,
    n6423, n6424, n6425, n6426, n6427, n6428,
    n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446,
    n6447, n6448, n6449, n6450, n6451, n6452,
    n6453, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470,
    n6471, n6472, n6473, n6474, n6475, n6476,
    n6477, n6478, n6479, n6480, n6481, n6482,
    n6483, n6484, n6485, n6486, n6487, n6488,
    n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500,
    n6501, n6502, n6503, n6504, n6505, n6506,
    n6507, n6508, n6509, n6510, n6511, n6512,
    n6513, n6514, n6515, n6516, n6517, n6518,
    n6519, n6520, n6521, n6522, n6523, n6524,
    n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6533, n6534, n6535, n6536,
    n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548,
    n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566,
    n6567, n6568, n6569, n6570, n6571, n6572,
    n6573, n6574, n6575, n6576, n6577, n6578,
    n6579, n6580, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6588, n6589, n6590,
    n6591, n6592, n6593, n6594, n6595, n6596,
    n6597, n6598, n6599, n6600, n6601, n6602,
    n6603, n6604, n6605, n6606, n6607, n6608,
    n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620,
    n6621, n6622, n6623, n6624, n6625, n6626,
    n6627, n6628, n6629, n6630, n6631, n6632,
    n6633, n6634, n6635, n6636, n6637, n6638,
    n6639, n6640, n6641, n6642, n6643, n6644,
    n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902,
    n6903, n6904, n6905, n6906, n6907, n6908,
    n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6937, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962,
    n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992,
    n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112,
    n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136,
    n7137, n7138, n7139, n7140, n7141, n7142,
    n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154,
    n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172,
    n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214,
    n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370,
    n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400,
    n7401, n7402, n7403, n7404, n7405, n7406,
    n7407, n7408, n7409, n7410, n7411, n7412,
    n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430,
    n7431, n7432, n7433, n7434, n7435, n7436,
    n7437, n7438, n7439, n7440, n7441, n7442,
    n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472,
    n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496,
    n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562,
    n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580,
    n7581, n7582, n7583, n7584, n7585, n7586,
    n7587, n7588, n7589, n7590, n7591, n7592,
    n7593, n7594, n7595, n7596, n7597, n7598,
    n7599, n7600, n7601, n7602, n7603, n7604,
    n7605, n7606, n7607, n7608, n7609, n7610,
    n7611, n7612, n7613, n7614, n7615, n7616,
    n7617, n7618, n7619, n7620, n7621, n7622,
    n7623, n7624, n7625, n7626, n7627, n7628,
    n7629, n7630, n7631, n7632, n7633, n7634,
    n7635, n7636, n7637, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7645, n7646,
    n7647, n7648, n7649, n7650, n7651, n7652,
    n7653, n7654, n7655, n7656, n7657, n7658,
    n7659, n7660, n7661, n7662, n7663, n7664,
    n7665, n7666, n7667, n7668, n7669, n7670,
    n7671, n7672, n7673, n7674, n7675, n7676,
    n7677, n7678, n7679, n7680, n7681, n7682,
    n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694,
    n7695, n7696, n7697, n7698, n7699, n7700,
    n7701, n7702, n7703, n7704, n7705, n7706,
    n7707, n7708, n7709, n7710, n7711, n7712,
    n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724,
    n7725, n7726, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7735, n7736,
    n7737, n7738, n7739, n7740, n7741, n7742,
    n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7760,
    n7761, n7762, n7763, n7764, n7765, n7766,
    n7767, n7768, n7769, n7770, n7771, n7772,
    n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790,
    n7791, n7792, n7793, n7794, n7795, n7796,
    n7797, n7798, n7799, n7800, n7801, n7802,
    n7803, n7804, n7805, n7806, n7807, n7808,
    n7809, n7810, n7811, n7812, n7813, n7814,
    n7815, n7816, n7817, n7818, n7819, n7820,
    n7821, n7822, n7823, n7824, n7825, n7826,
    n7827, n7828, n7829, n7830, n7831, n7832,
    n7833, n7834, n7835, n7836, n7837, n7838,
    n7839, n7840, n7841, n7842, n7843, n7844,
    n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7854, n7855, n7856,
    n7857, n7858, n7859, n7860, n7861, n7862,
    n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886,
    n7887, n7888, n7889, n7890, n7891, n7892,
    n7893, n7894, n7895, n7896, n7897, n7898,
    n7899, n7900, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922,
    n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7948, n7949, n7950, n7951, n7952,
    n7953, n7954, n7955, n7956, n7957, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976,
    n7977, n7978, n7979, n7980, n7981, n7982,
    n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012,
    n8013, n8014, n8015, n8016, n8017, n8018,
    n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042,
    n8043, n8044, n8045, n8046, n8047, n8048,
    n8049, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066,
    n8067, n8068, n8069, n8070, n8071, n8072,
    n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084,
    n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102,
    n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114,
    n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126,
    n8127, n8128, n8129, n8130, n8131, n8132,
    n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144,
    n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156,
    n8157, n8158, n8159, n8160, n8161, n8162,
    n8163, n8164, n8165, n8166, n8167, n8168,
    n8169, n8170, n8171, n8172, n8173, n8174,
    n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186,
    n8187, n8188, n8189, n8190, n8191, n8192,
    n8193, n8194, n8195, n8196, n8197, n8198,
    n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8219, n8220, n8221, n8222,
    n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246,
    n8247, n8248, n8249, n8250, n8251, n8252,
    n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8278, n8279, n8280, n8281, n8282,
    n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8290, n8291, n8292, n8293, n8294,
    n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306,
    n8307, n8308, n8309, n8310, n8311, n8312,
    n8313, n8314, n8315, n8316, n8317, n8318,
    n8319, n8320, n8321, n8322, n8323, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336,
    n8337, n8338, n8339, n8340, n8341, n8342,
    n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366,
    n8367, n8368, n8369, n8370, n8371, n8372,
    n8373, n8374, n8375, n8376, n8377, n8378,
    n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396,
    n8397, n8398, n8399, n8400, n8401, n8402,
    n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456,
    n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486,
    n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564,
    n8565, n8566, n8567, n8568, n8569, n8570,
    n8571, n8572, n8573, n8574, n8575, n8576,
    n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8593, n8594,
    n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606,
    n8607, n8608, n8609, n8610, n8611, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618,
    n8619, n8620, n8621, n8622, n8623, n8624,
    n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648,
    n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678,
    n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708,
    n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726,
    n8727, n8728, n8729, n8730, n8731, n8732,
    n8733, n8734, n8735, n8736, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756,
    n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768,
    n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786,
    n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816,
    n8817, n8818, n8819, n8820, n8821, n8822,
    n8823, n8824, n8825, n8826, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8834,
    n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846,
    n8847, n8848, n8849, n8850, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864,
    n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876,
    n8877, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888,
    n8889, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8902, n8903, n8904, n8905, n8906,
    n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936,
    n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966,
    n8967, n8968, n8969, n8970, n8971, n8972,
    n8973, n8974, n8975, n8976, n8977, n8978,
    n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n8993, n8994, n8995, n8996,
    n8997, n8998, n8999, n9000, n9001, n9002,
    n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9026,
    n9027, n9028, n9029, n9030, n9031, n9032,
    n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050,
    n9051, n9052, n9053, n9054, n9055, n9056,
    n9057, n9058, n9059, n9060, n9061, n9062,
    n9063, n9064, n9065, n9066, n9067, n9068,
    n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9080,
    n9081, n9082, n9083, n9084, n9085, n9086,
    n9087, n9088, n9089, n9090, n9091, n9092,
    n9093, n9094, n9095, n9096, n9097, n9098,
    n9099, n9100, n9101, n9102, n9103, n9104,
    n9105, n9106, n9107, n9108, n9109, n9110,
    n9111, n9112, n9113, n9114, n9115, n9116,
    n9117, n9118, n9119, n9120, n9121, n9122,
    n9123, n9124, n9125, n9126, n9127, n9128,
    n9129, n9130, n9131, n9132, n9133, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140,
    n9141, n9142, n9143, n9144, n9145, n9146,
    n9147, n9148, n9149, n9150, n9151, n9152,
    n9153, n9154, n9155, n9156, n9157, n9158,
    n9159, n9160, n9161, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170,
    n9171, n9172, n9173, n9174, n9175, n9176,
    n9177, n9178, n9179, n9180, n9181, n9182,
    n9183, n9184, n9185, n9186, n9187, n9188,
    n9189, n9190, n9191, n9192, n9193, n9194,
    n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206,
    n9207, n9208, n9209, n9210, n9211, n9212,
    n9213, n9214, n9215, n9216, n9217, n9218,
    n9219, n9220, n9221, n9222, n9223, n9224,
    n9225, n9226, n9227, n9228, n9229, n9230,
    n9231, n9232, n9233, n9234, n9235, n9236,
    n9237, n9238, n9239, n9240, n9241, n9242,
    n9243, n9244, n9245, n9246, n9247, n9248,
    n9249, n9250, n9251, n9252, n9253, n9254,
    n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266,
    n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296,
    n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326,
    n9327, n9328, n9329, n9330, n9331, n9332,
    n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386,
    n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416,
    n9417, n9418, n9419, n9420, n9421, n9422,
    n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446,
    n9447, n9448, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052,
    n10053, n10054, n10055, n10056, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064,
    n10065, n10066, n10067, n10068, n10069, n10070,
    n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10082,
    n10083, n10084, n10085, n10086, n10087, n10088,
    n10089, n10090, n10091, n10092, n10093, n10094,
    n10095, n10096, n10097, n10098, n10099, n10100,
    n10101, n10102, n10103, n10104, n10105, n10106,
    n10107, n10108, n10109, n10110, n10111, n10112,
    n10113, n10114, n10115, n10116, n10117, n10118,
    n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10128, n10129, n10130,
    n10131, n10132, n10133, n10134, n10135, n10136,
    n10137, n10138, n10139, n10140, n10141, n10142,
    n10143, n10144, n10145, n10146, n10147, n10148,
    n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10158, n10159, n10160,
    n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10169, n10170, n10171, n10172,
    n10173, n10174, n10175, n10176, n10177, n10178,
    n10179, n10180, n10181, n10182, n10183, n10184,
    n10185, n10186, n10187, n10188, n10189, n10190,
    n10191, n10192, n10193, n10194, n10195, n10196,
    n10197, n10198, n10199, n10200, n10201, n10202,
    n10203, n10204, n10205, n10206, n10207, n10208,
    n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10222, n10223, n10224, n10225, n10226,
    n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238,
    n10239, n10240, n10241, n10242, n10243, n10244,
    n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256,
    n10257, n10258, n10259, n10260, n10261, n10262,
    n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292,
    n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328,
    n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10370,
    n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382,
    n10383, n10384, n10385, n10386, n10387, n10388,
    n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406,
    n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424,
    n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442,
    n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460,
    n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472,
    n10473, n10474, n10475, n10476, n10477, n10478,
    n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490,
    n10491, n10492, n10493, n10494, n10495, n10496,
    n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514,
    n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532,
    n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10546, n10547, n10548, n10549, n10550,
    n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562,
    n10563, n10564, n10565, n10566, n10567, n10568,
    n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580,
    n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598,
    n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10651, n10652,
    n10653, n10654, n10655, n10656, n10657, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664,
    n10665, n10666, n10667, n10668, n10669, n10670,
    n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706,
    n10707, n10708, n10709, n10710, n10711, n10712,
    n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724,
    n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742,
    n10743, n10744, n10745, n10746, n10747, n10748,
    n10749, n10750, n10751, n10752, n10753, n10754,
    n10755, n10756, n10757, n10758, n10759, n10760,
    n10761, n10762, n10763, n10764, n10765, n10766,
    n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778,
    n10779, n10780, n10781, n10782, n10783, n10784,
    n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868,
    n10869, n10870, n10871, n10872, n10873, n10874,
    n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892,
    n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904,
    n10905, n10906, n10907, n10908, n10909, n10910,
    n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922,
    n10923, n10924, n10925, n10926, n10927, n10928,
    n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940,
    n10941, n10942, n10943, n10944, n10945, n10946,
    n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054,
    n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066,
    n11067, n11068, n11069, n11070, n11071, n11072,
    n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084,
    n11085, n11086, n11087, n11088, n11089, n11090,
    n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108,
    n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126,
    n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144,
    n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156,
    n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174,
    n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11189, n11190, n11191, n11192,
    n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204,
    n11205, n11206, n11207, n11208, n11209, n11210,
    n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222,
    n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11242, n11243, n11244, n11245, n11246,
    n11247, n11248, n11249, n11250, n11251, n11252,
    n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264,
    n11265, n11266, n11267, n11268, n11269, n11270,
    n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282,
    n11283, n11284, n11285, n11286, n11287, n11288,
    n11289, n11290, n11291, n11292, n11293, n11294,
    n11295, n11296, n11297, n11298, n11299, n11300,
    n11301, n11302, n11303, n11304, n11305, n11306,
    n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318,
    n11319, n11320, n11321, n11322, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336,
    n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354,
    n11355, n11356, n11357, n11358, n11359, n11360,
    n11361, n11362, n11363, n11364, n11365, n11366,
    n11367, n11368, n11369, n11370, n11371, n11372,
    n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11394, n11395, n11396,
    n11397, n11398, n11399, n11400, n11401, n11402,
    n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414,
    n11415, n11416, n11417, n11418, n11419, n11420,
    n11421, n11422, n11423, n11424, n11425, n11426,
    n11427, n11428, n11429, n11430, n11431, n11432,
    n11433, n11434, n11435, n11436, n11437, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444,
    n11445, n11446, n11447, n11448, n11449, n11450,
    n11451, n11452, n11453, n11454, n11455, n11456,
    n11457, n11458, n11459, n11460, n11461, n11462,
    n11463, n11464, n11465, n11466, n11467, n11468,
    n11469, n11470, n11471, n11472, n11473, n11474,
    n11475, n11476, n11477, n11478, n11479, n11480,
    n11481, n11482, n11483, n11484, n11485, n11486,
    n11487, n11488, n11489, n11490, n11491, n11492,
    n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504,
    n11505, n11506, n11507, n11508, n11509, n11510,
    n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11520, n11521, n11522,
    n11523, n11524, n11525, n11526, n11527, n11528,
    n11529, n11530, n11531, n11532, n11533, n11534,
    n11535, n11536, n11537, n11538, n11539, n11540,
    n11541, n11542, n11543, n11544, n11545, n11546,
    n11547, n11548, n11549, n11550, n11551, n11552,
    n11553, n11554, n11555, n11556, n11557, n11558,
    n11559, n11560, n11561, n11562, n11563, n11564,
    n11565, n11566, n11567, n11568, n11569, n11570,
    n11571, n11572, n11573, n11574, n11575, n11576,
    n11577, n11578, n11579, n11580, n11581, n11582,
    n11583, n11584, n11585, n11586, n11587, n11588,
    n11589, n11590, n11591, n11592, n11593, n11594,
    n11595, n11596, n11597, n11598, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618,
    n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630,
    n11631, n11632, n11633, n11634, n11635, n11636,
    n11637, n11638, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11648,
    n11649, n11650, n11651, n11652, n11653, n11654,
    n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666,
    n11667, n11668, n11669, n11670, n11671, n11672,
    n11673, n11674, n11675, n11676, n11677, n11678,
    n11679, n11680, n11681, n11682, n11683, n11684,
    n11685, n11686, n11687, n11688, n11689, n11690,
    n11691, n11692, n11693, n11694, n11695, n11696,
    n11697, n11698, n11699, n11700, n11701, n11702,
    n11703, n11704, n11705, n11706, n11707, n11708,
    n11709, n11710, n11711, n11712, n11713, n11714,
    n11715, n11716, n11717, n11718, n11719, n11720,
    n11721, n11722, n11723, n11724, n11725, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756,
    n11757, n11758, n11759, n11760, n11761, n11762,
    n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774,
    n11775, n11776, n11777, n11778, n11779, n11780,
    n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792,
    n11793, n11794, n11795, n11796, n11797, n11798,
    n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810,
    n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218,
    n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236,
    n12237, n12238, n12239, n12240, n12241, n12242,
    n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254,
    n12255, n12256, n12257, n12258, n12259, n12260,
    n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272,
    n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290,
    n12291, n12292, n12293, n12294, n12295, n12296,
    n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314,
    n12315, n12316, n12317, n12318, n12319, n12320,
    n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12340, n12341, n12342, n12343, n12344,
    n12345, n12346, n12347, n12348, n12349, n12350,
    n12351, n12352, n12353, n12354, n12355, n12356,
    n12357, n12358, n12359, n12360, n12361, n12362,
    n12363, n12364, n12365, n12366, n12367, n12368,
    n12369, n12370, n12371, n12372, n12373, n12374,
    n12375, n12376, n12377, n12378, n12379, n12380,
    n12381, n12382, n12383, n12384, n12385, n12386,
    n12387, n12388, n12389, n12390, n12391, n12392,
    n12393, n12394, n12395, n12396, n12397, n12398,
    n12399, n12400, n12401, n12402, n12403, n12404,
    n12405, n12406, n12407, n12408, n12409, n12410,
    n12411, n12412, n12413, n12414, n12415, n12416,
    n12417, n12418, n12419, n12420, n12421, n12422,
    n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434,
    n12435, n12436, n12437, n12438, n12439, n12440,
    n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452,
    n12453, n12454, n12455, n12456, n12457, n12458,
    n12459, n12460, n12461, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470,
    n12471, n12472, n12473, n12474, n12475, n12476,
    n12477, n12478, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488,
    n12489, n12490, n12491, n12492, n12493, n12494,
    n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506,
    n12507, n12508, n12509, n12510, n12511, n12512,
    n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524,
    n12525, n12526, n12527, n12528, n12529, n12530,
    n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542,
    n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560,
    n12561, n12562, n12563, n12564, n12565, n12566,
    n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578,
    n12579, n12580, n12581, n12582, n12583, n12584,
    n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596,
    n12597, n12598, n12599, n12600, n12601, n12602,
    n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614,
    n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632,
    n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650,
    n12651, n12652, n12653, n12654, n12655, n12656,
    n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668,
    n12669, n12670, n12671, n12672, n12673, n12674,
    n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12691, n12692,
    n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704,
    n12705, n12706, n12707, n12708, n12709, n12710,
    n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722,
    n12723, n12724, n12725, n12726, n12727, n12728,
    n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740,
    n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758,
    n12759, n12760, n12761, n12762, n12763, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776,
    n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794,
    n12795, n12796, n12797, n12798, n12799, n12800,
    n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812,
    n12813, n12814, n12815, n12816, n12817, n12818,
    n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12830,
    n12831, n12832, n12833, n12834, n12835, n12836,
    n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848,
    n12849, n12850, n12851, n12852, n12853, n12854,
    n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866,
    n12867, n12868, n12869, n12870, n12871, n12872,
    n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884,
    n12885, n12886, n12887, n12888, n12889, n12890,
    n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902,
    n12903, n12904, n12905, n12906, n12907, n12908,
    n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920,
    n12921, n12922, n12923, n12924, n12925, n12926,
    n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938,
    n12939, n12940, n12941, n12942, n12943, n12944,
    n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956,
    n12957, n12958, n12959, n12960, n12961, n12962,
    n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974,
    n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010,
    n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028,
    n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046,
    n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058,
    n13059, n13060, n13061, n13062, n13063, n13064,
    n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13073, n13074, n13075, n13076,
    n13077, n13078, n13079, n13080, n13081, n13082,
    n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100,
    n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112,
    n13113, n13114, n13115, n13116, n13117, n13118,
    n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130,
    n13131, n13132, n13133, n13134, n13135, n13136,
    n13137, n13138, n13139, n13140, n13141, n13142,
    n13143, n13144, n13145, n13146, n13147, n13148,
    n13149, n13150, n13151, n13152, n13153, n13154,
    n13155, n13156, n13157, n13158, n13159, n13160,
    n13161, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232,
    n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322,
    n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13354, n13355, n13356, n13357, n13358,
    n13359, n13360, n13361, n13362, n13363, n13364,
    n13365, n13366, n13367, n13368, n13369, n13370,
    n13371, n13372, n13373, n13374, n13375, n13376,
    n13377, n13378, n13379, n13380, n13381, n13382,
    n13383, n13384, n13385, n13386, n13387, n13388,
    n13389, n13390, n13391, n13392, n13393, n13394,
    n13395, n13396, n13397, n13398, n13399, n13400,
    n13401, n13402, n13403, n13404, n13405, n13406,
    n13407, n13408, n13409, n13410, n13411, n13412,
    n13413, n13414, n13415, n13416, n13417, n13418,
    n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430,
    n13431, n13432, n13433, n13434, n13435, n13436,
    n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448,
    n13449, n13450, n13451, n13452, n13453, n13454,
    n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13464, n13465, n13466,
    n13467, n13468, n13469, n13470, n13471, n13472,
    n13473, n13474, n13475, n13476, n13477, n13478,
    n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13486, n13487, n13488, n13489, n13490,
    n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502,
    n13503, n13504, n13505, n13506, n13507, n13508,
    n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13516, n13517, n13518, n13519, n13520,
    n13521, n13522, n13523, n13524, n13525, n13526,
    n13527, n13528, n13529, n13530, n13531, n13532,
    n13533, n13534, n13535, n13536, n13537, n13538,
    n13539, n13540, n13541, n13542, n13543, n13544,
    n13545, n13546, n13547, n13548, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562,
    n13563, n13564, n13565, n13566, n13567, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580,
    n13581, n13582, n13583, n13584, n13585, n13586,
    n13587, n13588, n13589, n13590, n13591, n13592,
    n13593, n13594, n13595, n13596, n13597, n13598,
    n13599, n13600, n13601, n13602, n13603, n13604,
    n13605, n13606, n13607, n13608, n13609, n13610,
    n13611, n13612, n13613, n13614, n13615, n13616,
    n13617, n13618, n13619, n13620, n13621, n13622,
    n13623, n13624, n13625, n13626, n13627, n13628,
    n13629, n13630, n13631, n13632, n13633, n13634,
    n13635, n13636, n13637, n13638, n13639, n13640,
    n13641, n13642, n13643, n13644, n13645, n13646,
    n13647, n13648, n13649, n13650, n13651, n13652,
    n13653, n13654, n13655, n13656, n13657, n13658,
    n13659, n13660, n13661, n13662, n13663, n13664,
    n13665, n13666, n13667, n13668, n13669, n13670,
    n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682,
    n13683, n13684, n13685, n13686, n13687, n13688,
    n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700,
    n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718,
    n13719, n13720, n13721, n13722, n13723, n13724,
    n13725, n13726, n13727, n13728, n13729, n13730,
    n13731, n13732, n13733, n13734, n13735, n13736,
    n13737, n13738, n13739, n13740, n13741, n13742,
    n13743, n13744, n13745, n13746, n13747, n13748,
    n13749, n13750, n13751, n13752, n13753, n13754,
    n13755, n13756, n13757, n13758, n13759, n13760,
    n13761, n13762, n13763, n13764, n13765, n13766,
    n13767, n13768, n13769, n13770, n13771, n13772,
    n13773, n13774, n13775, n13776, n13777, n13778,
    n13779, n13780, n13781, n13782, n13783, n13784,
    n13785, n13786, n13787, n13788, n13789, n13790,
    n13791, n13792, n13793, n13794, n13795, n13796,
    n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808,
    n13809, n13810, n13811, n13812, n13813, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826,
    n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844,
    n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862,
    n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880,
    n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898,
    n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916,
    n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934,
    n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952,
    n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970,
    n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988,
    n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006,
    n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060,
    n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078,
    n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144,
    n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330,
    n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348,
    n14349, n14350, n14351, n14352, n14353, n14354,
    n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372,
    n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14381, n14382, n14383, n14384,
    n14385, n14386, n14387, n14388, n14389, n14390,
    n14391, n14392, n14393, n14394, n14395, n14396,
    n14397, n14398, n14399, n14400, n14401, n14402,
    n14403, n14404, n14405, n14406, n14407, n14408,
    n14409, n14410, n14411, n14412, n14413, n14414,
    n14415, n14416, n14417, n14418, n14419, n14420,
    n14421, n14422, n14423, n14424, n14425, n14426,
    n14427, n14428, n14429, n14430, n14431, n14432,
    n14433, n14434, n14435, n14436, n14437, n14438,
    n14439, n14440, n14441, n14442, n14443, n14444,
    n14445, n14446, n14447, n14448, n14449, n14450,
    n14451, n14452, n14453, n14454, n14455, n14456,
    n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468,
    n14469, n14470, n14471, n14472, n14473, n14474,
    n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486,
    n14487, n14488, n14489, n14490, n14491, n14492,
    n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504,
    n14505, n14506, n14507, n14508, n14509, n14510,
    n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522,
    n14523, n14524, n14525, n14526, n14527, n14528,
    n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540,
    n14541, n14542, n14543, n14544, n14545, n14546,
    n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558,
    n14559, n14560, n14561, n14562, n14563, n14564,
    n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576,
    n14577, n14578, n14579, n14580, n14581, n14582,
    n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594,
    n14595, n14596, n14597, n14598, n14599, n14600,
    n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612,
    n14613, n14614, n14615, n14616, n14617, n14618,
    n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630,
    n14631, n14632, n14633, n14634, n14635, n14636,
    n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648,
    n14649, n14650, n14651, n14652, n14653, n14654,
    n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666,
    n14667, n14668, n14669, n14670, n14671, n14672,
    n14673, n14674, n14675, n14676, n14677, n14678,
    n14679, n14680, n14681, n14682, n14683, n14684,
    n14685, n14686, n14687, n14688, n14689, n14690,
    n14691, n14692, n14693, n14694, n14695, n14696,
    n14697, n14698, n14699, n14700, n14701, n14702,
    n14703, n14704, n14705, n14706, n14707, n14708,
    n14709, n14710, n14711, n14712, n14713, n14714,
    n14715, n14716, n14717, n14718, n14719, n14720,
    n14721, n14722, n14723, n14724, n14725, n14726,
    n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738,
    n14739, n14740, n14741, n14742, n14743, n14744,
    n14745, n14746, n14747, n14748, n14749, n14750,
    n14751, n14752, n14753, n14754, n14755, n14756,
    n14757, n14758, n14759, n14760, n14761, n14762,
    n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816,
    n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834,
    n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846,
    n14847, n14848, n14849, n14850, n14851, n14852,
    n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864,
    n14865, n14866, n14867, n14868, n14869, n14870,
    n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882,
    n14883, n14884, n14885, n14886, n14887, n14888,
    n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906,
    n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924,
    n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942,
    n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978,
    n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996,
    n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014,
    n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032,
    n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050,
    n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068,
    n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086,
    n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122,
    n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194,
    n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230,
    n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248,
    n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15281, n15282, n15283, n15284,
    n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302,
    n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314,
    n15315, n15316, n15317, n15318, n15319, n15320,
    n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338,
    n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15355, n15356,
    n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368,
    n15369, n15370, n15371, n15372, n15373, n15374,
    n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392,
    n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404,
    n15405, n15406, n15407, n15408, n15409, n15410,
    n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422,
    n15423, n15424, n15425, n15426, n15427, n15428,
    n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440,
    n15441, n15442, n15443, n15444, n15445, n15446,
    n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458,
    n15459, n15460, n15461, n15462, n15463, n15464,
    n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476,
    n15477, n15478, n15479, n15480, n15481, n15482,
    n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494,
    n15495, n15496, n15497, n15498, n15499, n15500,
    n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512,
    n15513, n15514, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530,
    n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15768, n15769, n15770,
    n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782,
    n15783, n15784, n15785, n15786, n15787, n15788,
    n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800,
    n15801, n15802, n15803, n15804, n15805, n15806,
    n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824,
    n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854,
    n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872,
    n15873, n15874, n15875, n15876, n15877, n15878,
    n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890,
    n15891, n15892, n15893, n15894, n15895, n15896,
    n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908,
    n15909, n15910, n15911, n15912, n15913, n15914,
    n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926,
    n15927, n15928, n15929, n15930, n15931, n15932,
    n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944,
    n15945, n15946, n15947, n15948, n15949, n15950,
    n15951, n15952, n15953, n15954, n15955, n15956,
    n15957, n15958, n15959, n15960, n15961, n15962,
    n15963, n15964, n15965, n15966, n15967, n15968,
    n15969, n15970, n15971, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980,
    n15981, n15982, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998,
    n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016,
    n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034,
    n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106,
    n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178,
    n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196,
    n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214,
    n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232,
    n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250,
    n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262,
    n16263, n16264, n16265, n16266, n16267, n16268,
    n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280,
    n16281, n16282, n16283, n16284, n16285, n16286,
    n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16302, n16303, n16304,
    n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316,
    n16317, n16318, n16319, n16320, n16321, n16322,
    n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334,
    n16335, n16336, n16337, n16338, n16339, n16340,
    n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352,
    n16353, n16354, n16355, n16356, n16357, n16358,
    n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370,
    n16371, n16372, n16373, n16374, n16375, n16376,
    n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388,
    n16389, n16390, n16391, n16392, n16393, n16394,
    n16395, n16396, n16397, n16398, n16399, n16400,
    n16401, n16402, n16403, n16404, n16405, n16406,
    n16407, n16408, n16409, n16410, n16411, n16412,
    n16413, n16414, n16415, n16416, n16417, n16418,
    n16419, n16420, n16421, n16422, n16423, n16424,
    n16425, n16426, n16427, n16428, n16429, n16430,
    n16431, n16432, n16433, n16434, n16435, n16436,
    n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448,
    n16449, n16450, n16451, n16452, n16453, n16454,
    n16455, n16456, n16457, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466,
    n16467, n16468, n16469, n16470, n16471, n16472,
    n16473, n16474, n16475, n16476, n16477, n16478,
    n16479, n16480, n16481, n16482, n16483, n16484,
    n16485, n16486, n16487, n16488, n16489, n16490,
    n16491, n16492, n16493, n16494, n16495, n16496,
    n16497, n16498, n16499, n16500, n16501, n16502,
    n16503, n16504, n16505, n16506, n16507, n16508,
    n16509, n16510, n16511, n16512, n16513, n16514,
    n16515, n16516, n16517, n16518, n16519, n16520,
    n16521, n16522, n16523, n16524, n16525, n16526,
    n16527, n16528, n16529, n16530, n16531, n16532,
    n16533, n16534, n16535, n16536, n16537, n16538,
    n16539, n16540, n16541, n16542, n16543, n16544,
    n16545, n16546, n16547, n16548, n16549, n16550,
    n16551, n16552, n16553, n16554, n16555, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562,
    n16563, n16564, n16565, n16566, n16567, n16568,
    n16569, n16570, n16571, n16572, n16573, n16574,
    n16575, n16576, n16577, n16578, n16579, n16580,
    n16581, n16582, n16583, n16584, n16585, n16586,
    n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598,
    n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652,
    n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670,
    n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16687, n16688,
    n16689, n16690, n16691, n16692, n16693, n16694,
    n16695, n16696, n16697, n16698, n16699, n16700,
    n16701, n16702, n16703, n16704, n16705, n16706,
    n16707, n16708, n16709, n16710, n16711, n16712,
    n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724,
    n16725, n16726, n16727, n16728, n16729, n16730,
    n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742,
    n16743, n16744, n16745, n16746, n16747, n16748,
    n16749, n16750, n16751, n16752, n16753, n16754,
    n16755, n16756, n16757, n16758, n16759, n16760,
    n16761, n16762, n16763, n16764, n16765, n16766,
    n16767, n16768, n16769, n16770, n16771, n16772,
    n16773, n16774, n16775, n16776, n16777, n16778,
    n16779, n16780, n16781, n16782, n16783, n16784,
    n16785, n16786, n16787, n16788, n16789, n16790,
    n16791, n16792, n16793, n16794, n16795, n16796,
    n16797, n16798, n16799, n16800, n16801, n16802,
    n16803, n16804, n16805, n16806, n16807, n16808,
    n16809, n16810, n16811, n16812, n16813, n16814,
    n16815, n16816, n16817, n16818, n16819, n16820,
    n16821, n16822, n16823, n16824, n16825, n16826,
    n16827, n16828, n16829, n16830, n16831, n16832,
    n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844,
    n16845, n16846, n16847, n16848, n16849, n16850,
    n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16868,
    n16869, n16870, n16871, n16872, n16873, n16874,
    n16875, n16876, n16877, n16878, n16879, n16880,
    n16881, n16882, n16883, n16884, n16885, n16886,
    n16887, n16888, n16889, n16890, n16891, n16892,
    n16893, n16894, n16895, n16896, n16897, n16898,
    n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16906, n16907, n16908, n16909, n16910,
    n16911, n16912, n16913, n16914, n16915, n16916,
    n16917, n16918, n16919, n16920, n16921, n16922,
    n16923, n16924, n16925, n16926, n16927, n16928,
    n16929, n16930, n16931, n16932, n16933, n16934,
    n16935, n16936, n16937, n16938, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16952,
    n16953, n16954, n16955, n16956, n16957, n16958,
    n16959, n16960, n16961, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976,
    n16977, n16978, n16979, n16980, n16981, n16982,
    n16983, n16984, n16985, n16986, n16987, n16988,
    n16989, n16990, n16991, n16992, n16993, n16994,
    n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17004, n17005, n17006,
    n17007, n17008, n17009, n17010, n17011, n17012,
    n17013, n17014, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024,
    n17025, n17026, n17027, n17028, n17029, n17030,
    n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042,
    n17043, n17044, n17045, n17046, n17047, n17048,
    n17049, n17050, n17051, n17052, n17053, n17054,
    n17055, n17056, n17057, n17058, n17059, n17060,
    n17061, n17062, n17063, n17064, n17065, n17066,
    n17067, n17068, n17069, n17070, n17071, n17072,
    n17073, n17074, n17075, n17076, n17077, n17078,
    n17079, n17080, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090,
    n17091, n17092, n17093, n17094, n17095, n17096,
    n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17114,
    n17115, n17116, n17117, n17118, n17119, n17120,
    n17121, n17122, n17123, n17124, n17125, n17126,
    n17127, n17128, n17129, n17130, n17131, n17132,
    n17133, n17134, n17135, n17136, n17137, n17138,
    n17139, n17140, n17141, n17142, n17143, n17144,
    n17145, n17146, n17147, n17148, n17149, n17150,
    n17151, n17152, n17153, n17154, n17155, n17156,
    n17157, n17158, n17159, n17160, n17161, n17162,
    n17163, n17164, n17165, n17166, n17167, n17168,
    n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180,
    n17181, n17182, n17183, n17184, n17185, n17186,
    n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204,
    n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222,
    n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240,
    n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258,
    n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276,
    n17277, n17278, n17279, n17280, n17281, n17282,
    n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294,
    n17295, n17296, n17297, n17298, n17299, n17300,
    n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312,
    n17313, n17314, n17315, n17316, n17317, n17318,
    n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330,
    n17331, n17332, n17333, n17334, n17335, n17336,
    n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348,
    n17349, n17350, n17351, n17352, n17353, n17354,
    n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366,
    n17367, n17368, n17369, n17370, n17371, n17372,
    n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384,
    n17385, n17386, n17387, n17388, n17389, n17390,
    n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402,
    n17403, n17404, n17405, n17406, n17407, n17408,
    n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420,
    n17421, n17422, n17423, n17424, n17425, n17426,
    n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438,
    n17439, n17440, n17441, n17442, n17443, n17444,
    n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456,
    n17457, n17458, n17459, n17460, n17461, n17462,
    n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474,
    n17475, n17476, n17477, n17478, n17479, n17480,
    n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492,
    n17493, n17494, n17495, n17496, n17497, n17498,
    n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510,
    n17511, n17512, n17513, n17514, n17515, n17516,
    n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528,
    n17529, n17530, n17531, n17532, n17533, n17534,
    n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546,
    n17547, n17548, n17549, n17550, n17551, n17552,
    n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564,
    n17565, n17566, n17567, n17568, n17569, n17570,
    n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582,
    n17583, n17584, n17585, n17586, n17587, n17588,
    n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624,
    n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672,
    n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696,
    n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708,
    n17709, n17710, n17711, n17712, n17713, n17714,
    n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726,
    n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744,
    n17745, n17746, n17747, n17748, n17749, n17750,
    n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762,
    n17763, n17764, n17765, n17766, n17767, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780,
    n17781, n17782, n17783, n17784, n17785, n17786,
    n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798,
    n17799, n17800, n17801, n17802, n17803, n17804,
    n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816,
    n17817, n17818, n17819, n17820, n17821, n17822,
    n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834,
    n17835, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852,
    n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888,
    n17889, n17890, n17891, n17892, n17893, n17894,
    n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906,
    n17907, n17908, n17909, n17910, n17911, n17912,
    n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17923, n17924,
    n17925, n17926, n17927, n17928, n17929, n17930,
    n17931, n17932, n17933, n17934, n17935, n17936,
    n17937, n17938, n17939, n17940, n17941, n17942,
    n17943, n17944, n17945, n17946, n17947, n17948,
    n17949, n17950, n17951, n17952, n17953, n17954,
    n17955, n17956, n17957, n17958, n17959, n17960,
    n17961, n17962, n17963, n17964, n17965, n17966,
    n17967, n17968, n17969, n17970, n17971, n17972,
    n17973, n17974, n17975, n17976, n17977, n17978,
    n17979, n17980, n17981, n17982, n17983, n17984,
    n17985, n17986, n17987, n17988, n17989, n17990,
    n17991, n17992, n17993, n17994, n17995, n17996,
    n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014,
    n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032,
    n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050,
    n18051, n18052, n18053, n18054, n18055, n18056,
    n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068,
    n18069, n18070, n18071, n18072, n18073, n18074,
    n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086,
    n18087, n18088, n18089, n18090, n18091, n18092,
    n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104,
    n18105, n18106, n18107, n18108, n18109, n18110,
    n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122,
    n18123, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140,
    n18141, n18142, n18143, n18144, n18145, n18146,
    n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158,
    n18159, n18160, n18161, n18162, n18163, n18164,
    n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176,
    n18177, n18178, n18179, n18180, n18181, n18182,
    n18183, n18184, n18185, n18186, n18187, n18188,
    n18189, n18190, n18191, n18192, n18193, n18194,
    n18195, n18196, n18197, n18198, n18199, n18200,
    n18201, n18202, n18203, n18204, n18205, n18206,
    n18207, n18208, n18209, n18210, n18211, n18212,
    n18213, n18214, n18215, n18216, n18217, n18218,
    n18219, n18220, n18221, n18222, n18223, n18224,
    n18225, n18226, n18227, n18228, n18229, n18230,
    n18231, n18232, n18233, n18234, n18235, n18236,
    n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18248,
    n18249, n18250, n18251, n18252, n18253, n18254,
    n18255, n18256, n18257, n18258, n18259, n18260,
    n18261, n18262, n18263, n18264, n18265, n18266,
    n18267, n18268, n18269, n18270, n18271, n18272,
    n18273, n18274, n18275, n18276, n18277, n18278,
    n18279, n18280, n18281, n18282, n18283, n18284,
    n18285, n18286, n18287, n18288, n18289, n18290,
    n18291, n18292, n18293, n18294, n18295, n18296,
    n18297, n18298, n18299, n18300, n18301, n18302,
    n18303, n18304, n18305, n18306, n18307, n18308,
    n18309, n18310, n18311, n18312, n18313, n18314,
    n18315, n18316, n18317, n18318, n18319, n18320,
    n18321, n18322, n18323, n18324, n18325, n18326,
    n18327, n18328, n18329, n18330, n18331, n18332,
    n18333, n18334, n18335, n18336, n18337, n18338,
    n18339, n18340, n18341, n18342, n18343, n18344,
    n18345, n18346, n18347, n18348, n18349, n18350,
    n18351, n18352, n18353, n18354, n18355, n18356,
    n18357, n18358, n18359, n18360, n18361, n18362,
    n18363, n18364, n18365, n18366, n18367, n18368,
    n18369, n18370, n18371, n18372, n18373, n18374,
    n18375, n18376, n18377, n18378, n18379, n18380,
    n18381, n18382, n18383, n18384, n18385, n18386,
    n18387, n18388, n18389, n18390, n18391, n18392,
    n18393, n18394, n18395, n18396, n18397, n18398,
    n18399, n18400, n18401, n18402, n18403, n18404,
    n18405, n18406, n18407, n18408, n18409, n18410,
    n18411, n18412, n18413, n18414, n18415, n18416,
    n18417, n18418, n18419, n18420, n18421, n18422,
    n18423, n18424, n18425, n18426, n18427, n18428,
    n18429, n18430, n18431, n18432, n18433, n18434,
    n18435, n18436, n18437, n18438, n18439, n18440,
    n18441, n18442, n18443, n18444, n18445, n18446,
    n18447, n18448, n18449, n18450, n18451, n18452,
    n18453, n18454, n18455, n18456, n18457, n18458,
    n18459, n18460, n18461, n18462, n18463, n18464,
    n18465, n18466, n18467, n18468, n18469, n18470,
    n18471, n18472, n18473, n18474, n18475, n18476,
    n18477, n18478, n18479, n18480, n18481, n18482,
    n18483, n18484, n18485, n18486, n18487, n18488,
    n18489, n18490, n18491, n18492, n18493, n18494,
    n18495, n18496, n18497, n18498, n18499, n18500,
    n18501, n18502, n18503, n18504, n18505, n18506,
    n18507, n18508, n18509, n18510, n18511, n18512,
    n18513, n18514, n18515, n18516, n18517, n18518,
    n18519, n18520, n18521, n18522, n18523, n18524,
    n18525, n18526, n18527, n18528, n18529, n18530,
    n18531, n18532, n18533, n18534, n18535, n18536,
    n18537, n18538, n18539, n18540, n18541, n18542,
    n18543, n18544, n18545, n18546, n18547, n18548,
    n18549, n18550, n18551, n18552, n18553, n18554,
    n18555, n18556, n18557, n18558, n18559, n18560,
    n18561, n18562, n18563, n18564, n18565, n18566,
    n18567, n18568, n18569, n18570, n18571, n18572,
    n18573, n18574, n18575, n18576, n18577, n18578,
    n18579, n18580, n18581, n18582, n18583, n18584,
    n18585, n18586, n18587, n18588, n18589, n18590,
    n18591, n18592, n18593, n18594, n18595, n18596,
    n18597, n18598, n18599, n18600, n18601, n18602,
    n18603, n18604, n18605, n18606, n18607, n18608,
    n18609, n18610, n18611, n18612, n18613, n18614,
    n18615, n18616, n18617, n18618, n18619, n18620,
    n18621, n18622, n18623, n18624, n18625, n18626,
    n18627, n18628, n18629, n18630, n18631, n18632,
    n18633, n18634, n18635, n18636, n18637, n18638,
    n18639, n18640, n18641, n18642, n18643, n18644,
    n18645, n18646, n18647, n18648, n18649, n18650,
    n18651, n18652, n18653, n18654, n18655, n18656,
    n18657, n18658, n18659, n18660, n18661, n18662,
    n18663, n18664, n18665, n18666, n18667, n18668,
    n18669, n18670, n18671, n18672, n18673, n18674,
    n18675, n18676, n18677, n18678, n18679, n18680,
    n18681, n18682, n18683, n18684, n18685, n18686,
    n18687, n18688, n18689, n18690, n18691, n18692,
    n18693, n18694, n18695, n18696, n18697, n18698,
    n18699, n18700, n18701, n18702, n18703, n18704,
    n18705, n18706, n18707, n18708, n18709, n18710,
    n18711, n18712, n18713, n18714, n18715, n18716,
    n18717, n18718, n18719, n18720, n18721, n18722,
    n18723, n18724, n18725, n18726, n18727, n18728,
    n18729, n18730, n18731, n18732, n18733, n18734,
    n18735, n18736, n18737, n18738, n18739, n18740,
    n18741, n18742, n18743, n18744, n18745, n18746,
    n18747, n18748, n18749, n18750, n18751, n18752,
    n18753, n18754, n18755, n18756, n18757, n18758,
    n18759, n18760, n18761, n18762, n18763, n18764,
    n18765, n18766, n18767, n18768, n18769, n18770,
    n18771, n18772, n18773, n18774, n18775, n18776,
    n18777, n18778, n18779, n18780, n18781, n18782,
    n18783, n18784, n18785, n18786, n18787, n18788,
    n18789, n18790, n18791, n18792, n18793, n18794,
    n18795, n18796, n18797, n18798, n18799, n18800,
    n18801, n18802, n18803, n18804, n18805, n18806,
    n18807, n18808, n18809, n18810, n18811, n18812,
    n18813, n18814, n18815, n18816, n18817, n18818,
    n18819, n18820, n18821, n18822, n18823, n18824,
    n18825, n18826, n18827, n18828, n18829, n18830,
    n18831, n18832, n18833, n18834, n18835, n18836,
    n18837, n18838, n18839, n18840, n18841, n18842,
    n18843, n18844, n18845, n18846, n18847, n18848,
    n18849, n18850, n18851, n18852, n18853, n18854,
    n18855, n18856, n18857, n18858, n18859, n18860,
    n18861, n18862, n18863, n18864, n18865, n18866,
    n18867, n18868, n18869, n18870, n18871, n18872,
    n18873, n18874, n18875, n18876, n18877, n18878,
    n18879, n18880, n18881, n18882, n18883, n18884,
    n18885, n18886, n18887, n18888, n18889, n18890,
    n18891, n18892, n18893, n18894, n18895, n18896,
    n18897, n18898, n18899, n18900, n18901, n18902,
    n18903, n18904, n18905, n18906, n18907, n18908,
    n18909, n18910, n18911, n18912, n18913, n18914,
    n18915, n18916, n18917, n18918, n18919, n18920,
    n18921, n18922, n18923, n18924, n18925, n18926,
    n18927, n18928, n18929, n18930, n18931, n18932,
    n18933, n18934, n18935, n18936, n18937, n18938,
    n18939, n18940, n18941, n18942, n18943, n18944,
    n18945, n18946, n18947, n18948, n18949, n18950,
    n18951, n18952, n18953, n18954, n18955, n18956,
    n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968,
    n18969, n18970, n18971, n18972, n18973, n18974,
    n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986,
    n18987, n18988, n18989, n18990, n18991, n18992,
    n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004,
    n19005, n19006, n19007, n19008, n19009, n19010,
    n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022,
    n19023, n19024, n19025, n19026, n19027, n19028,
    n19029, n19030, n19031, n19032, n19033, n19034,
    n19035, n19036, n19037, n19038, n19039, n19040,
    n19041, n19042, n19043, n19044, n19045, n19046,
    n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058,
    n19059, n19060, n19061, n19062, n19063, n19064,
    n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076,
    n19077, n19078, n19079, n19080, n19081, n19082,
    n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094,
    n19095, n19096, n19097, n19098, n19099, n19100,
    n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112,
    n19113, n19114, n19115, n19116, n19117, n19118,
    n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130,
    n19131, n19132, n19133, n19134, n19135, n19136,
    n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148,
    n19149, n19150, n19151, n19152, n19153, n19154,
    n19155, n19156, n19157, n19158, n19159, n19160,
    n19161, n19162, n19163, n19164, n19165, n19166,
    n19167, n19168, n19169, n19170, n19171, n19172,
    n19173, n19174, n19175, n19176, n19177, n19178,
    n19179, n19180, n19181, n19182, n19183, n19184,
    n19185, n19186, n19187, n19188, n19189, n19190,
    n19191, n19192, n19193, n19194, n19195, n19196,
    n19197, n19198, n19199, n19200, n19201, n19202,
    n19203, n19204, n19205, n19206, n19207, n19208,
    n19209, n19210, n19211, n19212, n19213, n19214,
    n19215, n19216, n19217, n19218, n19219, n19220,
    n19221, n19222, n19223, n19224, n19225, n19226,
    n19227, n19228, n19229, n19230, n19231, n19232,
    n19233, n19234, n19235, n19236, n19237, n19238,
    n19239, n19240, n19241, n19242, n19243, n19244,
    n19245, n19246, n19247, n19248, n19249, n19250,
    n19251, n19252, n19253, n19254, n19255, n19256,
    n19257, n19258, n19259, n19260, n19261, n19262,
    n19263, n19264, n19265, n19266, n19267, n19268,
    n19269, n19270, n19271, n19272, n19273, n19274,
    n19275, n19276, n19277, n19278, n19279, n19280,
    n19281, n19282, n19283, n19284, n19285, n19286,
    n19287, n19288, n19289, n19290, n19291, n19292,
    n19293, n19294, n19295, n19296, n19297, n19298,
    n19299, n19300, n19301, n19302, n19303, n19304,
    n19305, n19306, n19307, n19308, n19309, n19310,
    n19311, n19312, n19313, n19314, n19315, n19316,
    n19317, n19318, n19319, n19320, n19321, n19322,
    n19323, n19324, n19325, n19326, n19327, n19328,
    n19329, n19330, n19331, n19332, n19333, n19334,
    n19335, n19336, n19337, n19338, n19339, n19340,
    n19341, n19342, n19343, n19344, n19345, n19346,
    n19347, n19348, n19349, n19350, n19351, n19352,
    n19353, n19354, n19355, n19356, n19357, n19358,
    n19359, n19360, n19361, n19362, n19363, n19364,
    n19365, n19366, n19367, n19368, n19369, n19370,
    n19371, n19372, n19373, n19374, n19375, n19376,
    n19377, n19378, n19379, n19380, n19381, n19382,
    n19383, n19384, n19385, n19386, n19387, n19388,
    n19389, n19390, n19391, n19392, n19393, n19394,
    n19395, n19396, n19397, n19398, n19399, n19400,
    n19401, n19402, n19403, n19404, n19405, n19406,
    n19407, n19408, n19409, n19410, n19411, n19412,
    n19413, n19414, n19415, n19416, n19417, n19418,
    n19419, n19420, n19421, n19422, n19423, n19424,
    n19425, n19426, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19435, n19436,
    n19437, n19438, n19439, n19440, n19441, n19442,
    n19443, n19444, n19445, n19446, n19447, n19448,
    n19449, n19450, n19451, n19452, n19453, n19454,
    n19455, n19456, n19457, n19458, n19459, n19460,
    n19461, n19462, n19463, n19464, n19465, n19466,
    n19467, n19468, n19469, n19470, n19471, n19472,
    n19473, n19474, n19475, n19476, n19477, n19478,
    n19479, n19480, n19481, n19482, n19483, n19484,
    n19485, n19486, n19487, n19488, n19489, n19490,
    n19491, n19492, n19493, n19494, n19495, n19496,
    n19497, n19498, n19499, n19500, n19501, n19502,
    n19503, n19504, n19505, n19506, n19507, n19508,
    n19509, n19510, n19511, n19512, n19513, n19514,
    n19515, n19516, n19517, n19518, n19519, n19520,
    n19521, n19522, n19523, n19524, n19525, n19526,
    n19527, n19528, n19529, n19530, n19531, n19532,
    n19533, n19534, n19535, n19536, n19537, n19538,
    n19539, n19540, n19541, n19542, n19543, n19544,
    n19545, n19546, n19547, n19548, n19549, n19550,
    n19551, n19552, n19553, n19554, n19555, n19556,
    n19557, n19558, n19559, n19560, n19561, n19562,
    n19563, n19564, n19565, n19566, n19567, n19568,
    n19569, n19570, n19571, n19572, n19573, n19574,
    n19575, n19576, n19577, n19578, n19579, n19580,
    n19581, n19582, n19583, n19584, n19585, n19586,
    n19587, n19588, n19589, n19590, n19591, n19592,
    n19593, n19594, n19595, n19596, n19597, n19598,
    n19599, n19600, n19601, n19602, n19603, n19604,
    n19605, n19606, n19607, n19608, n19609, n19610,
    n19611, n19612, n19613, n19614, n19615, n19616,
    n19617, n19618, n19619, n19620, n19621, n19622,
    n19623, n19624, n19625, n19626, n19627, n19628,
    n19629, n19630, n19631, n19632, n19633, n19634,
    n19635, n19636, n19637, n19638, n19639, n19640,
    n19641, n19642, n19643, n19644, n19645, n19646,
    n19647, n19648, n19649, n19650, n19651, n19652,
    n19653, n19654, n19655, n19656, n19657, n19658,
    n19659, n19660, n19661, n19662, n19663, n19664,
    n19665, n19666, n19667, n19668, n19669, n19670,
    n19671, n19672, n19673, n19674, n19675, n19676,
    n19677, n19678, n19679, n19680, n19681, n19682,
    n19683, n19684, n19685, n19686, n19687, n19688,
    n19689, n19690, n19691, n19692, n19693, n19694,
    n19695, n19696, n19697, n19698, n19699, n19700,
    n19701, n19702, n19703, n19704, n19705, n19706,
    n19707, n19708, n19709, n19710, n19711, n19712,
    n19713, n19714, n19715, n19716, n19717, n19718,
    n19719, n19720, n19721, n19722, n19723, n19724,
    n19725, n19726, n19727, n19728, n19729, n19730,
    n19731, n19732, n19733, n19734, n19735, n19736,
    n19737, n19738, n19739, n19740, n19741, n19742,
    n19743, n19744, n19745, n19746, n19747, n19748,
    n19749, n19750, n19751, n19752, n19753, n19754,
    n19755, n19756, n19757, n19758, n19759, n19760,
    n19761, n19762, n19763, n19764, n19765, n19766,
    n19767, n19768, n19769, n19770, n19771, n19772,
    n19773, n19774, n19775, n19776, n19777, n19778,
    n19779, n19780, n19781, n19782, n19783, n19784,
    n19785, n19786, n19787, n19788, n19789, n19790,
    n19791, n19792, n19793, n19794, n19795, n19796,
    n19797, n19798, n19799, n19800, n19801, n19802,
    n19803, n19804, n19805, n19806, n19807, n19808,
    n19809, n19810, n19811, n19812, n19813, n19814,
    n19815, n19816, n19817, n19818, n19819, n19820,
    n19821, n19822, n19823, n19824, n19825, n19826,
    n19827, n19828, n19829, n19830, n19831, n19832,
    n19833, n19834, n19835, n19836, n19837, n19838,
    n19839, n19840, n19841, n19842, n19843, n19844,
    n19845, n19846, n19847, n19848, n19849, n19850,
    n19851, n19852, n19853, n19854, n19855, n19856,
    n19857, n19858, n19859, n19860, n19861, n19862,
    n19863, n19864, n19865, n19866, n19867, n19868,
    n19869, n19870, n19871, n19872, n19873, n19874,
    n19875, n19876, n19877, n19878, n19879, n19880,
    n19881, n19882, n19883, n19884, n19885, n19886,
    n19887, n19888, n19889, n19890, n19891, n19892,
    n19893, n19894, n19895, n19896, n19897, n19898,
    n19899, n19900, n19901, n19902, n19903, n19904,
    n19905, n19906, n19907, n19908, n19909, n19910,
    n19911, n19912, n19913, n19914, n19915, n19916,
    n19917, n19918, n19919, n19920, n19921, n19922,
    n19923, n19924, n19925, n19926, n19927, n19928,
    n19929, n19930, n19931, n19932, n19933, n19934,
    n19935, n19936, n19937, n19938, n19939, n19940,
    n19941, n19942, n19943, n19944, n19945, n19946,
    n19947, n19948, n19949, n19950, n19951, n19952,
    n19953, n19954, n19955, n19956, n19957, n19958,
    n19959, n19960, n19961, n19962, n19963, n19964,
    n19965, n19966, n19967, n19968, n19969, n19970,
    n19971, n19972, n19973, n19974, n19975, n19976,
    n19977, n19978, n19979, n19980, n19981, n19982,
    n19983, n19984, n19985, n19986, n19987, n19988,
    n19989, n19990, n19991, n19992, n19993, n19994,
    n19995, n19996, n19997, n19998, n19999, n20000,
    n20001, n20002, n20003, n20004, n20005, n20006,
    n20007, n20008, n20009, n20010, n20011, n20012,
    n20013, n20014, n20015, n20016, n20017, n20018,
    n20019, n20020, n20021, n20022, n20023, n20024,
    n20025, n20026, n20027, n20028, n20029, n20030,
    n20031, n20032, n20033, n20034, n20035, n20036,
    n20037, n20038, n20039, n20040, n20041, n20042,
    n20043, n20044, n20045, n20046, n20047, n20048,
    n20049, n20050, n20051, n20052, n20053, n20054,
    n20055, n20056, n20057, n20058, n20059, n20060,
    n20061, n20062, n20063, n20064, n20065, n20066,
    n20067, n20068, n20069, n20070, n20071, n20072,
    n20073, n20074, n20075, n20076, n20077, n20078,
    n20079, n20080, n20081, n20082, n20083, n20084,
    n20085, n20086, n20087, n20088, n20089, n20090,
    n20091, n20092, n20093, n20094, n20095, n20096,
    n20097, n20098, n20099, n20100, n20101, n20102,
    n20103, n20104, n20105, n20106, n20107, n20108,
    n20109, n20110, n20111, n20112, n20113, n20114,
    n20115, n20116, n20117, n20118, n20119, n20120,
    n20121, n20122, n20123, n20124, n20125, n20126,
    n20127, n20128, n20129, n20130, n20131, n20132,
    n20133, n20134, n20135, n20136, n20137, n20138,
    n20139, n20140, n20141, n20142, n20143, n20144,
    n20145, n20146, n20147, n20148, n20149, n20150,
    n20151, n20152, n20153, n20154, n20155, n20156,
    n20157, n20158, n20159, n20160, n20161, n20162,
    n20163, n20164, n20165, n20166, n20167, n20168,
    n20169, n20170, n20171, n20172, n20173, n20174,
    n20175, n20176, n20177, n20178, n20179, n20180,
    n20181, n20182, n20183, n20184, n20185, n20186,
    n20187, n20188, n20189, n20190, n20191, n20192,
    n20193, n20194, n20195, n20196, n20197, n20198,
    n20199, n20200, n20201, n20202, n20203, n20204,
    n20205, n20206, n20207, n20208, n20209, n20210,
    n20211, n20212, n20213, n20214, n20215, n20216,
    n20217, n20218, n20219, n20220, n20221, n20222,
    n20223, n20224, n20225, n20226, n20227, n20228,
    n20229, n20230, n20231, n20232, n20233, n20234,
    n20235, n20236, n20237, n20238, n20239, n20240,
    n20241, n20242, n20243, n20244, n20245, n20246,
    n20247, n20248, n20249, n20250, n20251, n20252,
    n20253, n20254, n20255, n20256, n20257, n20258,
    n20259, n20260, n20261, n20262, n20263, n20264,
    n20265, n20266, n20267, n20268, n20269, n20270,
    n20271, n20272, n20273, n20274, n20275, n20276,
    n20277, n20278, n20279, n20280, n20281, n20282,
    n20283, n20284, n20285, n20286, n20287, n20288,
    n20289, n20290, n20291, n20292, n20293, n20294,
    n20295, n20296, n20297, n20298, n20299, n20300,
    n20301, n20302, n20303, n20304, n20305, n20306,
    n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318,
    n20319, n20320, n20321, n20322, n20323, n20324,
    n20325, n20326, n20327, n20328, n20329, n20330,
    n20331, n20332, n20333, n20334, n20335, n20336,
    n20337, n20338, n20339, n20340, n20341, n20342,
    n20343, n20344, n20345, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354,
    n20355, n20356, n20357, n20358, n20359, n20360,
    n20361, n20362, n20363, n20364, n20365, n20366,
    n20367, n20368, n20369, n20370, n20371, n20372,
    n20373, n20374, n20375, n20376, n20377, n20378,
    n20379, n20380, n20381, n20382, n20383, n20384,
    n20385, n20386, n20387, n20388, n20389, n20390,
    n20391, n20392, n20393, n20394, n20395, n20396,
    n20397, n20398, n20399, n20400, n20401, n20402,
    n20403, n20404, n20405, n20406, n20407, n20408,
    n20409, n20410, n20411, n20412, n20413, n20414,
    n20415, n20416, n20417, n20418, n20419, n20420,
    n20421, n20422, n20423, n20424, n20425, n20426,
    n20427, n20428, n20429, n20430, n20431, n20432,
    n20433, n20434, n20435, n20436, n20437, n20438,
    n20439, n20440, n20441, n20442, n20443, n20444,
    n20445, n20446, n20447, n20448, n20449, n20450,
    n20451, n20452, n20453, n20454, n20455, n20456,
    n20457, n20458, n20459, n20460, n20461, n20462,
    n20463, n20464, n20465, n20466, n20467, n20468,
    n20469, n20470, n20471, n20472, n20473, n20474,
    n20475, n20476, n20477, n20478, n20479, n20480,
    n20481, n20482, n20483, n20484, n20485, n20486,
    n20487, n20488, n20489, n20490, n20491, n20492,
    n20493, n20494, n20495, n20496, n20497, n20498,
    n20499, n20500, n20501, n20502, n20503, n20504,
    n20505, n20506, n20507, n20508, n20509, n20510,
    n20511, n20512, n20513, n20514, n20515, n20516,
    n20517, n20518, n20519, n20520, n20521, n20522,
    n20523, n20524, n20525, n20526, n20527, n20528,
    n20529, n20530, n20531, n20532, n20533, n20534,
    n20535, n20536, n20537, n20538, n20539, n20540,
    n20541, n20542, n20543, n20544, n20545, n20546,
    n20547, n20548, n20549, n20550, n20551, n20552,
    n20553, n20554, n20555, n20556, n20557, n20558,
    n20559, n20560, n20561, n20562, n20563, n20564,
    n20565, n20566, n20567, n20568, n20569, n20570,
    n20571, n20572, n20573, n20574, n20575, n20576,
    n20577, n20578, n20579, n20580, n20581, n20582,
    n20583, n20584, n20585, n20586, n20587, n20588,
    n20589, n20590, n20591, n20592, n20593, n20594,
    n20595, n20596, n20597, n20598, n20599, n20600,
    n20601, n20602, n20603, n20604, n20605, n20606,
    n20607, n20608, n20609, n20610, n20611, n20612,
    n20613, n20614, n20615, n20616, n20617, n20618,
    n20619, n20620, n20621, n20622, n20623, n20624,
    n20625, n20626, n20627, n20628, n20629, n20630,
    n20631, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20645, n20646, n20647, n20648,
    n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660,
    n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20675, n20676, n20677, n20678,
    n20679, n20680, n20681, n20682, n20683, n20684,
    n20685, n20686, n20687, n20688, n20689, n20690,
    n20691, n20692, n20693, n20694, n20695, n20696,
    n20697, n20698, n20699, n20700, n20701, n20702,
    n20703, n20704, n20705, n20706, n20707, n20708,
    n20709, n20710, n20711, n20712, n20713, n20714,
    n20715, n20716, n20717, n20718, n20719, n20720,
    n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732,
    n20733, n20734, n20735, n20736, n20737, n20738,
    n20739, n20740, n20741, n20742, n20743, n20744,
    n20745, n20746, n20747, n20748, n20749, n20750,
    n20751, n20752, n20753, n20754, n20755, n20756,
    n20757, n20758, n20759, n20760, n20761, n20762,
    n20763, n20764, n20765, n20766, n20767, n20768,
    n20769, n20770, n20771, n20772, n20773, n20774,
    n20775, n20776, n20777, n20778, n20779, n20780,
    n20781, n20782, n20783, n20784, n20785, n20786,
    n20787, n20788, n20789, n20790, n20791, n20792,
    n20793, n20794, n20795, n20796, n20797, n20798,
    n20799, n20800, n20801, n20802, n20803, n20804,
    n20805, n20806, n20807, n20808, n20809, n20810,
    n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822,
    n20823, n20824, n20825, n20826, n20827, n20828,
    n20829, n20830, n20831, n20832, n20833, n20834,
    n20835, n20836, n20837, n20838, n20839, n20840,
    n20841, n20842, n20843, n20844, n20845, n20846,
    n20847, n20848, n20849, n20850, n20851, n20852,
    n20853, n20854, n20855, n20856, n20857, n20858,
    n20859, n20860, n20861, n20862, n20863, n20864,
    n20865, n20866, n20867, n20868, n20869, n20870,
    n20871, n20872, n20873, n20874, n20875, n20876,
    n20877, n20878, n20879, n20880, n20881, n20882,
    n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20892, n20893, n20894,
    n20895, n20896, n20897, n20898, n20899, n20900,
    n20901, n20902, n20903, n20904, n20905, n20906,
    n20907, n20908, n20909, n20910, n20911, n20912,
    n20913, n20914, n20915, n20916, n20917, n20918,
    n20919, n20920, n20921, n20922, n20923, n20924,
    n20925, n20926, n20927, n20928, n20929, n20930,
    n20931, n20932, n20933, n20934, n20935, n20936,
    n20937, n20938, n20939, n20940, n20941, n20942,
    n20943, n20944, n20945, n20946, n20947, n20948,
    n20949, n20950, n20951, n20952, n20953, n20954,
    n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972,
    n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984,
    n20985, n20986, n20987, n20988, n20989, n20990,
    n20991, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008,
    n21009, n21010, n21011, n21012, n21013, n21014,
    n21015, n21016, n21017, n21018, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026,
    n21027, n21028, n21029, n21030, n21031, n21032,
    n21033, n21034, n21035, n21036, n21037, n21038,
    n21039, n21040, n21041, n21042, n21043, n21044,
    n21045, n21046, n21047, n21048, n21049, n21050,
    n21051, n21052, n21053, n21054, n21055, n21056,
    n21057, n21058, n21059, n21060, n21061, n21062,
    n21063, n21064, n21065, n21066, n21067, n21068,
    n21069, n21070, n21071, n21072, n21073, n21074,
    n21075, n21076, n21077, n21078, n21079, n21080,
    n21081, n21082, n21083, n21084, n21085, n21086,
    n21087, n21088, n21089, n21090, n21091, n21092,
    n21093, n21094, n21095, n21096, n21097, n21098,
    n21099, n21100, n21101, n21102, n21103, n21104,
    n21105, n21106, n21107, n21108, n21109, n21110,
    n21111, n21112, n21113, n21114, n21115, n21116,
    n21117, n21118, n21119, n21120, n21121, n21122,
    n21123, n21124, n21125, n21126, n21127, n21128,
    n21129, n21130, n21131, n21132, n21133, n21134,
    n21135, n21136, n21137, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21145, n21146,
    n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158,
    n21159, n21160, n21161, n21162, n21163, n21164,
    n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176,
    n21177, n21178, n21179, n21180, n21181, n21182,
    n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200,
    n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218,
    n21219, n21220, n21221, n21222, n21223, n21224,
    n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236,
    n21237, n21238, n21239, n21240, n21241, n21242,
    n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260,
    n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21278,
    n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290,
    n21291, n21292, n21293, n21294, n21295, n21296,
    n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314,
    n21315, n21316, n21317, n21318, n21319, n21320,
    n21321, n21322, n21323, n21324, n21325, n21326,
    n21327, n21328, n21329, n21330, n21331, n21332,
    n21333, n21334, n21335, n21336, n21337, n21338,
    n21339, n21340, n21341, n21342, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350,
    n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368,
    n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428,
    n21429, n21430, n21431, n21432, n21433, n21434,
    n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21446,
    n21447, n21448, n21449, n21450, n21451, n21452,
    n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464,
    n21465, n21466, n21467, n21468, n21469, n21470,
    n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482,
    n21483, n21484, n21485, n21486, n21487, n21488,
    n21489, n21490, n21491, n21492, n21493, n21494,
    n21495, n21496, n21497, n21498, n21499, n21500,
    n21501, n21502, n21503, n21504, n21505, n21506,
    n21507, n21508, n21509, n21510, n21511, n21512,
    n21513, n21514, n21515, n21516, n21517, n21518,
    n21519, n21520, n21521, n21522, n21523, n21524,
    n21525, n21526, n21527, n21528, n21529, n21530,
    n21531, n21532, n21533, n21534, n21535, n21536,
    n21537, n21538, n21539, n21540, n21541, n21542,
    n21543, n21544, n21545, n21546, n21547, n21548,
    n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560,
    n21561, n21562, n21563, n21564, n21565, n21566,
    n21567, n21568, n21569, n21570, n21571, n21572,
    n21573, n21574, n21575, n21576, n21577, n21578,
    n21579, n21580, n21581, n21582, n21583, n21584,
    n21585, n21586, n21587, n21588, n21589, n21590,
    n21591, n21592, n21593, n21594, n21595, n21596,
    n21597, n21598, n21599, n21600, n21601, n21602,
    n21603, n21604, n21605, n21606, n21607, n21608,
    n21609, n21610, n21611, n21612, n21613, n21614,
    n21615, n21616, n21617, n21618, n21619, n21620,
    n21621, n21622, n21623, n21624, n21625, n21626,
    n21627, n21628, n21629, n21630, n21631, n21632,
    n21633, n21634, n21635, n21636, n21637, n21638,
    n21639, n21640, n21641, n21642, n21643, n21644,
    n21645, n21646, n21647, n21648, n21649, n21650,
    n21651, n21652, n21653, n21654, n21655, n21656,
    n21657, n21658, n21659, n21660, n21661, n21662,
    n21663, n21664, n21665, n21666, n21667, n21668,
    n21669, n21670, n21671, n21672, n21673, n21674,
    n21675, n21676, n21677, n21678, n21679, n21680,
    n21681, n21682, n21683, n21684, n21685, n21686,
    n21687, n21688, n21689, n21690, n21691, n21692,
    n21693, n21694, n21695, n21696, n21697, n21698,
    n21699, n21700, n21701, n21702, n21703, n21704,
    n21705, n21706, n21707, n21708, n21709, n21710,
    n21711, n21712, n21713, n21714, n21715, n21716,
    n21717, n21718, n21719, n21720, n21721, n21722,
    n21723, n21724, n21725, n21726, n21727, n21728,
    n21729, n21730, n21731, n21732, n21733, n21734,
    n21735, n21736, n21737, n21738, n21739, n21740,
    n21741, n21742, n21743, n21744, n21745, n21746,
    n21747, n21748, n21749, n21750, n21751, n21752,
    n21753, n21754, n21755, n21756, n21757, n21758,
    n21759, n21760, n21761, n21762, n21763, n21764,
    n21765, n21766, n21767, n21768, n21769, n21770,
    n21771, n21772, n21773, n21774, n21775, n21776,
    n21777, n21778, n21779, n21780, n21781, n21782,
    n21783, n21784, n21785, n21786, n21787, n21788,
    n21789, n21790, n21791, n21792, n21793, n21794,
    n21795, n21796, n21797, n21798, n21799, n21800,
    n21801, n21802, n21803, n21804, n21805, n21806,
    n21807, n21808, n21809, n21810, n21811, n21812,
    n21813, n21814, n21815, n21816, n21817, n21818,
    n21819, n21820, n21821, n21822, n21823, n21824,
    n21825, n21826, n21827, n21828, n21829, n21830,
    n21831, n21832, n21833, n21834, n21835, n21836,
    n21837, n21838, n21839, n21840, n21841, n21842,
    n21843, n21844, n21845, n21846, n21847, n21848,
    n21849, n21850, n21851, n21852, n21853, n21854,
    n21855, n21856, n21857, n21858, n21859, n21860,
    n21861, n21862, n21863, n21864, n21865, n21866,
    n21867, n21868, n21869, n21870, n21871, n21872,
    n21873, n21874, n21875, n21876, n21877, n21878,
    n21879, n21880, n21881, n21882, n21883, n21884,
    n21885, n21886, n21887, n21888, n21889, n21890,
    n21891, n21892, n21893, n21894, n21895, n21896,
    n21897, n21898, n21899, n21900, n21901, n21902,
    n21903, n21904, n21905, n21906, n21907, n21908,
    n21909, n21910, n21911, n21912, n21913, n21914,
    n21915, n21916, n21917, n21918, n21919, n21920,
    n21921, n21922, n21923, n21924, n21925, n21926,
    n21927, n21928, n21929, n21930, n21931, n21932,
    n21933, n21934, n21935, n21936, n21937, n21938,
    n21939, n21940, n21941, n21942, n21943, n21944,
    n21945, n21946, n21947, n21948, n21949, n21950,
    n21951, n21952, n21953, n21954, n21955, n21956,
    n21957, n21958, n21959, n21960, n21961, n21962,
    n21963, n21964, n21965, n21966, n21967, n21968,
    n21969, n21970, n21971, n21972, n21973, n21974,
    n21975, n21976, n21977, n21978, n21979, n21980,
    n21981, n21982, n21983, n21984, n21985, n21986,
    n21987, n21988, n21989, n21990, n21991, n21992,
    n21993, n21994, n21995, n21996, n21997, n21998,
    n21999, n22000, n22001, n22002, n22003, n22004,
    n22005, n22006, n22007, n22008, n22009, n22010,
    n22011, n22012, n22013, n22014, n22015, n22016,
    n22017, n22018, n22019, n22020, n22021, n22022,
    n22023, n22024, n22025, n22026, n22027, n22028,
    n22029, n22030, n22031, n22032, n22033, n22034,
    n22035, n22036, n22037, n22038, n22039, n22040,
    n22041, n22042, n22043, n22044, n22045, n22046,
    n22047, n22048, n22049, n22050, n22051, n22052,
    n22053, n22054, n22055, n22056, n22057, n22058,
    n22059, n22060, n22061, n22062, n22063, n22064,
    n22065, n22066, n22067, n22068, n22069, n22070,
    n22071, n22072, n22073, n22074, n22075, n22076,
    n22077, n22078, n22079, n22080, n22081, n22082,
    n22083, n22084, n22085, n22086, n22087, n22088,
    n22089, n22090, n22091, n22092, n22093, n22094,
    n22095, n22096, n22097, n22098, n22099, n22100,
    n22101, n22102, n22103, n22104, n22105, n22106,
    n22107, n22108, n22109, n22110, n22111, n22112,
    n22113, n22114, n22115, n22116, n22117, n22118,
    n22119, n22120, n22121, n22122, n22123, n22124,
    n22125, n22126, n22127, n22128, n22129, n22130,
    n22131, n22132, n22133, n22134, n22135, n22136,
    n22137, n22138, n22139, n22140, n22141, n22142,
    n22143, n22144, n22145, n22146, n22147, n22148,
    n22149, n22150, n22151, n22152, n22153, n22154,
    n22155, n22156, n22157, n22158, n22159, n22160,
    n22161, n22162, n22163, n22164, n22165, n22166,
    n22167, n22168, n22169, n22170, n22171, n22172,
    n22173, n22174, n22175, n22176, n22177, n22178,
    n22179, n22180, n22181, n22182, n22183, n22184,
    n22185, n22186, n22187, n22188, n22189, n22190,
    n22191, n22192, n22193, n22194, n22195, n22196,
    n22197, n22198, n22199, n22200, n22201, n22202,
    n22203, n22204, n22205, n22206, n22207, n22208,
    n22209, n22210, n22211, n22212, n22213, n22214,
    n22215, n22216, n22217, n22218, n22219, n22220,
    n22221, n22222, n22223, n22224, n22225, n22226,
    n22227, n22228, n22229, n22230, n22231, n22232,
    n22233, n22234, n22235, n22236, n22237, n22238,
    n22239, n22240, n22241, n22242, n22243, n22244,
    n22245, n22246, n22247, n22248, n22249, n22250,
    n22251, n22252, n22253, n22254, n22255, n22256,
    n22257, n22258, n22259, n22260, n22261, n22262,
    n22263, n22264, n22265, n22266, n22267, n22268,
    n22269, n22270, n22271, n22272, n22273, n22274,
    n22275, n22276, n22277, n22278, n22279, n22280,
    n22281, n22282, n22283, n22284, n22285, n22286,
    n22287, n22288, n22289, n22290, n22291, n22292,
    n22293, n22294, n22295, n22296, n22297, n22298,
    n22299, n22300, n22301, n22302, n22303, n22304,
    n22305, n22306, n22307, n22308, n22309, n22310,
    n22311, n22312, n22313, n22314, n22315, n22316,
    n22317, n22318, n22319, n22320, n22321, n22322,
    n22323, n22324, n22325, n22326, n22327, n22328,
    n22329, n22330, n22331, n22332, n22333, n22334,
    n22335, n22336, n22337, n22338, n22339, n22340,
    n22341, n22342, n22343, n22344, n22345, n22346,
    n22347, n22348, n22349, n22350, n22351, n22352,
    n22353, n22354, n22355, n22356, n22357, n22358,
    n22359, n22360, n22361, n22362, n22363, n22364,
    n22365, n22366, n22367, n22368, n22369, n22370,
    n22371, n22372, n22373, n22374, n22375, n22376,
    n22377, n22378, n22379, n22380, n22381, n22382,
    n22383, n22384, n22385, n22386, n22387, n22388,
    n22389, n22390, n22391, n22392, n22393, n22394,
    n22395, n22396, n22397, n22398, n22399, n22400,
    n22401, n22402, n22403, n22404, n22405, n22406,
    n22407, n22408, n22409, n22410, n22411, n22412,
    n22413, n22414, n22415, n22416, n22417, n22418,
    n22419, n22420, n22421, n22422, n22423, n22424,
    n22425, n22426, n22427, n22428, n22429, n22430,
    n22431, n22432, n22433, n22434, n22435, n22436,
    n22437, n22438, n22439, n22440, n22441, n22442,
    n22443, n22444, n22445, n22446, n22447, n22448,
    n22449, n22450, n22451, n22452, n22453, n22454,
    n22455, n22456, n22457, n22458, n22459, n22460,
    n22461, n22462, n22463, n22464, n22465, n22466,
    n22467, n22468, n22469, n22470, n22471, n22472,
    n22473, n22474, n22475, n22476, n22477, n22478,
    n22479, n22480, n22481, n22482, n22483, n22484,
    n22485, n22486, n22487, n22488, n22489, n22490,
    n22491, n22492, n22493, n22494, n22495, n22496,
    n22497, n22498, n22499, n22500, n22501, n22502,
    n22503, n22504, n22505, n22506, n22507, n22508,
    n22509, n22510, n22511, n22512, n22513, n22514,
    n22515, n22516, n22517, n22518, n22519, n22520,
    n22521, n22522, n22523, n22524, n22525, n22526,
    n22527, n22528, n22529, n22530, n22531, n22532,
    n22533, n22534, n22535, n22536, n22537, n22538,
    n22539, n22540, n22541, n22542, n22543, n22544,
    n22545, n22546, n22547, n22548, n22549, n22550,
    n22551, n22552, n22553, n22554, n22555, n22556,
    n22557, n22558, n22559, n22560, n22561, n22562,
    n22563, n22564, n22565, n22566, n22567, n22568,
    n22569, n22570, n22571, n22572, n22573, n22574,
    n22575, n22576, n22577, n22578, n22579, n22580,
    n22581, n22582, n22583, n22584, n22585, n22586,
    n22587, n22588, n22589, n22590, n22591, n22592,
    n22593, n22594, n22595, n22596, n22597, n22598,
    n22599, n22600, n22601, n22602, n22603, n22604,
    n22605, n22606, n22607, n22608, n22609, n22610,
    n22611, n22612, n22613, n22614, n22615, n22616,
    n22617, n22618, n22619, n22620, n22621, n22622,
    n22623, n22624, n22625, n22626, n22627, n22628,
    n22629, n22630, n22631, n22632, n22633, n22634,
    n22635, n22636, n22637, n22638, n22639, n22640,
    n22641, n22642, n22643, n22644, n22645, n22646,
    n22647, n22648, n22649, n22650, n22651, n22652,
    n22653, n22654, n22655, n22656, n22657, n22658,
    n22659, n22660, n22661, n22662, n22663, n22664,
    n22665, n22666, n22667, n22668, n22669, n22670,
    n22671, n22672, n22673, n22674, n22675, n22676,
    n22677, n22678, n22679, n22680, n22681, n22682,
    n22683, n22684, n22685, n22686, n22687, n22688,
    n22689, n22690, n22691, n22692, n22693, n22694,
    n22695, n22696, n22697, n22698, n22699, n22700,
    n22701, n22702, n22703, n22704, n22705, n22706,
    n22707, n22708, n22709, n22710, n22711, n22712,
    n22713, n22714, n22715, n22716, n22717, n22718,
    n22719, n22720, n22721, n22722, n22723, n22724,
    n22725, n22726, n22727, n22728, n22729, n22730,
    n22731, n22732, n22733, n22734, n22735, n22736,
    n22737, n22738, n22739, n22740, n22741, n22742,
    n22743, n22744, n22745, n22746, n22747, n22748,
    n22749, n22750, n22751, n22752, n22753, n22754,
    n22755, n22756, n22757, n22758, n22759, n22760,
    n22761, n22762, n22763, n22764, n22765, n22766,
    n22767, n22768, n22769, n22770, n22771, n22772,
    n22773, n22774, n22775, n22776, n22777, n22778,
    n22779, n22780, n22781, n22782, n22783, n22784,
    n22785, n22786, n22787, n22788, n22789, n22790,
    n22791, n22792, n22793, n22794, n22795, n22796,
    n22797, n22798, n22799, n22800, n22801, n22802,
    n22803, n22804, n22805, n22806, n22807, n22808,
    n22809, n22810, n22811, n22812, n22813, n22814,
    n22815, n22816, n22817, n22818, n22819, n22820,
    n22821, n22822, n22823, n22824, n22825, n22826,
    n22827, n22828, n22829, n22830, n22831, n22832,
    n22833, n22834, n22835, n22836, n22837, n22838,
    n22839, n22840, n22841, n22842, n22843, n22844,
    n22845, n22846, n22847, n22848, n22849, n22850,
    n22851, n22852, n22853, n22854, n22855, n22856,
    n22857, n22858, n22859, n22860, n22861, n22862,
    n22863, n22864, n22865, n22866, n22867, n22868,
    n22869, n22870, n22871, n22872, n22873, n22874,
    n22875, n22876, n22877, n22878, n22879, n22880,
    n22881, n22882, n22883, n22884, n22885, n22886,
    n22887, n22888, n22889, n22890, n22891, n22892,
    n22893, n22894, n22895, n22896, n22897, n22898,
    n22899, n22900, n22901, n22902, n22903, n22904,
    n22905, n22906, n22907, n22908, n22909, n22910,
    n22911, n22912, n22913, n22914, n22915, n22916,
    n22917, n22918, n22919, n22920, n22921, n22922,
    n22923, n22924, n22925, n22926, n22927, n22928,
    n22929, n22930, n22931, n22932, n22933, n22934,
    n22935, n22936, n22937, n22938, n22939, n22940,
    n22941, n22942, n22943, n22944, n22945, n22946,
    n22947, n22948, n22949, n22950, n22951, n22952,
    n22953, n22954, n22955, n22956, n22957, n22958,
    n22959, n22960, n22961, n22962, n22963, n22964,
    n22965, n22966, n22967, n22968, n22969, n22970,
    n22971, n22972, n22973, n22974, n22975, n22976,
    n22977, n22978, n22979, n22980, n22981, n22982,
    n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994,
    n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012,
    n23013, n23014, n23015, n23016, n23017, n23018,
    n23019, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n23028, n23029, n23030,
    n23031, n23032, n23033, n23034, n23035, n23036,
    n23037, n23038, n23039, n23040, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048,
    n23049, n23050, n23051, n23052, n23053, n23054,
    n23055, n23056, n23057, n23058, n23059, n23060,
    n23061, n23062, n23063, n23064, n23065, n23066,
    n23067, n23068, n23069, n23070, n23071, n23072,
    n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084,
    n23085, n23086, n23087, n23088, n23089, n23090,
    n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102,
    n23103, n23104, n23105, n23106, n23107, n23108,
    n23109, n23110, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120,
    n23121, n23122, n23123, n23124, n23125, n23126,
    n23127, n23128, n23129, n23130, n23131, n23132,
    n23133, n23134, n23135, n23136, n23137, n23138,
    n23139, n23140, n23141, n23142, n23143, n23144,
    n23145, n23146, n23147, n23148, n23149, n23150,
    n23151, n23152, n23153, n23154, n23155, n23156,
    n23157, n23158, n23159, n23160, n23161, n23162,
    n23163, n23164, n23165, n23166, n23167, n23168,
    n23169, n23170, n23171, n23172, n23173, n23174,
    n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186,
    n23187, n23188, n23189, n23190, n23191, n23192,
    n23193, n23194, n23195, n23196, n23197, n23198,
    n23199, n23200, n23201, n23202, n23203, n23204,
    n23205, n23206, n23207, n23208, n23209, n23210,
    n23211, n23212, n23213, n23214, n23215, n23216,
    n23217, n23218, n23219, n23220, n23221, n23222,
    n23223, n23224, n23225, n23226, n23227, n23228,
    n23229, n23230, n23231, n23232, n23233, n23234,
    n23235, n23236, n23237, n23238, n23239, n23240,
    n23241, n23242, n23243, n23244, n23245, n23246,
    n23247, n23248, n23249, n23250, n23251, n23252,
    n23253, n23254, n23255, n23256, n23257, n23258,
    n23259, n23260, n23261, n23262, n23263, n23264,
    n23265, n23266, n23267, n23268, n23269, n23270,
    n23271, n23272, n23273, n23274, n23275, n23276,
    n23277, n23278, n23279, n23280, n23281, n23282,
    n23283, n23284, n23285, n23286, n23287, n23288,
    n23289, n23290, n23291, n23292, n23293, n23294,
    n23295, n23296, n23297, n23298, n23299, n23300,
    n23301, n23302, n23303, n23304, n23305, n23306,
    n23307, n23308, n23309, n23310, n23311, n23312,
    n23313, n23314, n23315, n23316, n23317, n23318,
    n23319, n23320, n23321, n23322, n23323, n23324,
    n23325, n23326, n23327, n23328, n23329, n23330,
    n23331, n23332, n23333, n23334, n23335, n23336,
    n23337, n23338, n23339, n23340, n23341, n23342,
    n23343, n23344, n23345, n23346, n23347, n23348,
    n23349, n23350, n23351, n23352, n23353, n23354,
    n23355, n23356, n23357, n23358, n23359, n23360,
    n23361, n23362, n23363, n23364, n23365, n23366,
    n23367, n23368, n23369, n23370, n23371, n23372,
    n23373, n23374, n23375, n23376, n23377, n23378,
    n23379, n23380, n23381, n23382, n23383, n23384,
    n23385, n23386, n23387, n23388, n23389, n23390,
    n23391, n23392, n23393, n23394, n23395, n23396,
    n23397, n23398, n23399, n23400, n23401, n23402,
    n23403, n23404, n23405, n23406, n23407, n23408,
    n23409, n23410, n23411, n23412, n23413, n23414,
    n23415, n23416, n23417, n23418, n23419, n23420,
    n23421, n23422, n23423, n23424, n23425, n23426,
    n23427, n23428, n23429, n23430, n23431, n23432,
    n23433, n23434, n23435, n23436, n23437, n23438,
    n23439, n23440, n23441, n23442, n23443, n23444,
    n23445, n23446, n23447, n23448, n23449, n23450,
    n23451, n23452, n23453, n23454, n23455, n23456,
    n23457, n23458, n23459, n23460, n23461, n23462,
    n23463, n23464, n23465, n23466, n23467, n23468,
    n23469, n23470, n23471, n23472, n23473, n23474,
    n23475, n23476, n23477, n23478, n23479, n23480,
    n23481, n23482, n23483, n23484, n23485, n23486,
    n23487, n23488, n23489, n23490, n23491, n23492,
    n23493, n23494, n23495, n23496, n23497, n23498,
    n23499, n23500, n23501, n23502, n23503, n23504,
    n23505, n23506, n23507, n23508, n23509, n23510,
    n23511, n23512, n23513, n23514, n23515, n23516,
    n23517, n23518, n23519, n23520, n23521, n23522,
    n23523, n23524, n23525, n23526, n23527, n23528,
    n23529, n23530, n23531, n23532, n23533, n23534,
    n23535, n23536, n23537, n23538, n23539, n23540,
    n23541, n23542, n23543, n23544, n23545, n23546,
    n23547, n23548, n23549, n23550, n23551, n23552,
    n23553, n23554, n23555, n23556, n23557, n23558,
    n23559, n23560, n23561, n23562, n23563, n23564,
    n23565, n23566, n23567, n23568, n23569, n23570,
    n23571, n23572, n23573, n23574, n23575, n23576,
    n23577, n23578, n23579, n23580, n23581, n23582,
    n23583, n23584, n23585, n23586, n23587, n23588,
    n23589, n23590, n23591, n23592, n23593, n23594,
    n23595, n23596, n23597, n23598, n23599, n23600,
    n23601, n23602, n23603, n23604, n23605, n23606,
    n23607, n23608, n23609, n23610, n23611, n23612,
    n23613, n23614, n23615, n23616, n23617, n23618,
    n23619, n23620, n23621, n23622, n23623, n23624,
    n23625, n23626, n23627, n23628, n23629, n23630,
    n23631, n23632, n23633, n23634, n23635, n23636,
    n23637, n23638, n23639, n23640, n23641, n23642,
    n23643, n23644, n23645, n23646, n23647, n23648,
    n23649, n23650, n23651, n23652, n23653, n23654,
    n23655, n23656, n23657, n23658, n23659, n23660,
    n23661, n23662, n23663, n23664, n23665, n23666,
    n23667, n23668, n23669, n23670, n23671, n23672,
    n23673, n23674, n23675, n23676, n23677, n23678,
    n23679, n23680, n23681, n23682, n23683, n23684,
    n23685, n23686, n23687, n23688, n23689, n23690,
    n23691, n23692, n23693, n23694, n23695, n23696,
    n23697, n23698, n23699, n23700, n23701, n23702,
    n23703, n23704, n23705, n23706, n23707, n23708,
    n23709, n23710, n23711, n23712, n23713, n23714,
    n23715, n23716, n23717, n23718, n23719, n23720,
    n23721, n23722, n23723, n23724, n23725, n23726,
    n23727, n23728, n23729, n23730, n23731, n23732,
    n23733, n23734, n23735, n23736, n23737, n23738,
    n23739, n23740, n23741, n23742, n23743, n23744,
    n23745, n23746, n23747, n23748, n23749, n23750,
    n23751, n23752, n23753, n23754, n23755, n23756,
    n23757, n23758, n23759, n23760, n23761, n23762,
    n23763, n23764, n23765, n23766, n23767, n23768,
    n23769, n23770, n23771, n23772, n23773, n23774,
    n23775, n23776, n23777, n23778, n23779, n23780,
    n23781, n23782, n23783, n23784, n23785, n23786,
    n23787, n23788, n23789, n23790, n23791, n23792,
    n23793, n23794, n23795, n23796, n23797, n23798,
    n23799, n23800, n23801, n23802, n23803, n23804,
    n23805, n23806, n23807, n23808, n23809, n23810,
    n23811, n23812, n23813, n23814, n23815, n23816,
    n23817, n23818, n23819, n23820, n23821, n23822,
    n23823, n23824, n23825, n23826, n23827, n23828,
    n23829, n23830, n23831, n23832, n23833, n23834,
    n23835, n23836, n23837, n23838, n23839, n23840,
    n23841, n23842, n23843, n23844, n23845, n23846,
    n23847, n23848, n23849, n23850, n23851, n23852,
    n23853, n23854, n23855, n23856, n23857, n23858,
    n23859, n23860, n23861, n23862, n23863, n23864,
    n23865, n23866, n23867, n23868, n23869, n23870,
    n23871, n23872, n23873, n23874, n23875, n23876,
    n23877, n23878, n23879, n23880, n23881, n23882,
    n23883, n23884, n23885, n23886, n23887, n23888,
    n23889, n23890, n23891, n23892, n23893, n23894,
    n23895, n23896, n23897, n23898, n23899, n23900,
    n23901, n23902, n23903, n23904, n23905, n23906,
    n23907, n23908, n23909, n23910, n23911, n23912,
    n23913, n23914, n23915, n23916, n23917, n23918,
    n23919, n23920, n23921, n23922, n23923, n23924,
    n23925, n23926, n23927, n23928, n23929, n23930,
    n23931, n23932, n23933, n23934, n23935, n23936,
    n23937, n23938, n23939, n23940, n23941, n23942,
    n23943, n23944, n23945, n23946, n23947, n23948,
    n23949, n23950, n23951, n23952, n23953, n23954,
    n23955, n23956, n23957, n23958, n23959, n23960,
    n23961, n23962, n23963, n23964, n23965, n23966,
    n23967, n23968, n23969, n23970, n23971, n23972,
    n23973, n23974, n23975, n23976, n23977, n23978,
    n23979, n23980, n23981, n23982, n23983, n23984,
    n23985, n23986, n23987, n23988, n23989, n23990,
    n23991, n23992, n23993, n23994, n23995, n23996,
    n23997, n23998, n23999, n24000, n24001, n24002,
    n24003, n24004, n24005, n24006, n24007, n24008,
    n24009, n24010, n24011, n24012, n24013, n24014,
    n24015, n24016, n24017, n24018, n24019, n24020,
    n24021, n24022, n24023, n24024, n24025, n24026,
    n24027, n24028, n24029, n24030, n24031, n24032,
    n24033, n24034, n24035, n24036, n24037, n24038,
    n24039, n24040, n24041, n24042, n24043, n24044,
    n24045, n24046, n24047, n24048, n24049, n24050,
    n24051, n24052, n24053, n24054, n24055, n24056,
    n24057, n24058, n24059, n24060, n24061, n24062,
    n24063, n24064, n24065, n24066, n24067, n24068,
    n24069, n24070, n24071, n24072, n24073, n24074,
    n24075, n24076, n24077, n24078, n24079, n24080,
    n24081, n24082, n24083, n24084, n24085, n24086,
    n24087, n24088, n24089, n24090, n24091, n24092,
    n24093, n24094, n24095, n24096, n24097, n24098,
    n24099, n24100, n24101, n24102, n24103, n24104,
    n24105, n24106, n24107, n24108, n24109, n24110,
    n24111, n24112, n24113, n24114, n24115, n24116,
    n24117, n24118, n24119, n24120, n24121, n24122,
    n24123, n24124, n24125, n24126, n24127, n24128,
    n24129, n24130, n24131, n24132, n24133, n24134,
    n24135, n24136, n24137, n24138, n24139, n24140,
    n24141, n24142, n24143, n24144, n24145, n24146,
    n24147, n24148, n24149, n24150, n24151, n24152,
    n24153, n24154, n24155, n24156, n24157, n24158,
    n24159, n24160, n24161, n24162, n24163, n24164,
    n24165, n24166, n24167, n24168, n24169, n24170,
    n24171, n24172, n24173, n24174, n24175, n24176,
    n24177, n24178, n24179, n24180, n24181, n24182,
    n24183, n24184, n24185, n24186, n24187, n24188,
    n24189, n24190, n24191, n24192, n24193, n24194,
    n24195, n24196, n24197, n24198, n24199, n24200,
    n24201, n24202, n24203, n24204, n24205, n24206,
    n24207, n24208, n24209, n24210, n24211, n24212,
    n24213, n24214, n24215, n24216, n24217, n24218,
    n24219, n24220, n24221, n24222, n24223, n24224,
    n24225, n24226, n24227, n24228, n24229, n24230,
    n24231, n24232, n24233, n24234, n24235, n24236,
    n24237, n24238, n24239, n24240, n24241, n24242,
    n24243, n24244, n24245, n24246, n24247, n24248,
    n24249, n24250, n24251, n24252, n24253, n24254,
    n24255, n24256, n24257, n24258, n24259, n24260,
    n24261, n24262, n24263, n24264, n24265, n24266,
    n24267, n24268, n24269, n24270, n24271, n24272,
    n24273, n24274, n24275, n24276, n24277, n24278,
    n24279, n24280, n24281, n24282, n24283, n24284,
    n24285, n24286, n24287, n24288, n24289, n24290,
    n24291, n24292, n24293, n24294, n24295, n24296,
    n24297, n24298, n24299, n24300, n24301, n24302,
    n24303, n24304, n24305, n24306, n24307, n24308,
    n24309, n24310, n24311, n24312, n24313, n24314,
    n24315, n24316, n24317, n24318, n24319, n24320,
    n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332,
    n24333, n24334, n24335, n24336, n24337, n24338,
    n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350,
    n24351, n24352, n24353, n24354, n24355, n24356,
    n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368,
    n24369, n24370, n24371, n24372, n24373, n24374,
    n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386,
    n24387, n24388, n24389, n24390, n24391, n24392,
    n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404,
    n24405, n24406, n24407, n24408, n24409, n24410,
    n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422,
    n24423, n24424, n24425, n24426, n24427, n24428,
    n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440,
    n24441, n24442, n24443, n24444, n24445, n24446,
    n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24458,
    n24459, n24460, n24461, n24462, n24463, n24464,
    n24465, n24466, n24467, n24468, n24469, n24470,
    n24471, n24472, n24473, n24474, n24475, n24476,
    n24477, n24478, n24479, n24480, n24481, n24482,
    n24483, n24484, n24485, n24486, n24487, n24488,
    n24489, n24490, n24491, n24492, n24493, n24494,
    n24495, n24496, n24497, n24498, n24499, n24500,
    n24501, n24502, n24503, n24504, n24505, n24506,
    n24507, n24508, n24509, n24510, n24511, n24512,
    n24513, n24514, n24515, n24516, n24517, n24518,
    n24519, n24520, n24521, n24522, n24523, n24524,
    n24525, n24526, n24527, n24528, n24529, n24530,
    n24531, n24532, n24533, n24534, n24535, n24536,
    n24537, n24538, n24539, n24540, n24541, n24542,
    n24543, n24544, n24545, n24546, n24547, n24548,
    n24549, n24550, n24551, n24552, n24553, n24554,
    n24555, n24556, n24557, n24558, n24559, n24560,
    n24561, n24562, n24563, n24564, n24565, n24566,
    n24567, n24568, n24569, n24570, n24571, n24572,
    n24573, n24574, n24575, n24576, n24577, n24578,
    n24579, n24580, n24581, n24582, n24583, n24584,
    n24585, n24586, n24587, n24588, n24589, n24590,
    n24591, n24592, n24593, n24594, n24595, n24596,
    n24597, n24598, n24599, n24600, n24601, n24602,
    n24603, n24604, n24605, n24606, n24607, n24608,
    n24609, n24610, n24611, n24612, n24613, n24614,
    n24615, n24616, n24617, n24618, n24619, n24620,
    n24621, n24622, n24623, n24624, n24625, n24626,
    n24627, n24628, n24629, n24630, n24631, n24632,
    n24633, n24634, n24635, n24636, n24637, n24638,
    n24639, n24640, n24641, n24642, n24643, n24644,
    n24645, n24646, n24647, n24648, n24649, n24650,
    n24651, n24652, n24653, n24654, n24655, n24656,
    n24657, n24658, n24659, n24660, n24661, n24662,
    n24663, n24664, n24665, n24666, n24667, n24668,
    n24669, n24670, n24671, n24672, n24673, n24674,
    n24675, n24676, n24677, n24678, n24679, n24680,
    n24681, n24682, n24683, n24684, n24685, n24686,
    n24687, n24688, n24689, n24690, n24691, n24692,
    n24693, n24694, n24695, n24696, n24697, n24698,
    n24699, n24700, n24701, n24702, n24703, n24704,
    n24705, n24706, n24707, n24708, n24709, n24710,
    n24711, n24712, n24713, n24714, n24715, n24716,
    n24717, n24718, n24719, n24720, n24721, n24722,
    n24723, n24724, n24725, n24726, n24727, n24728,
    n24729, n24730, n24731, n24732, n24733, n24734,
    n24735, n24736, n24737, n24738, n24739, n24740,
    n24741, n24742, n24743, n24744, n24745, n24746,
    n24747, n24748, n24749, n24750, n24751, n24752,
    n24753, n24754, n24755, n24756, n24757, n24758,
    n24759, n24760, n24761, n24762, n24763, n24764,
    n24765, n24766, n24767, n24768, n24769, n24770,
    n24771, n24772, n24773, n24774, n24775, n24776,
    n24777, n24778, n24779, n24780, n24781, n24782,
    n24783, n24784, n24785, n24786, n24787, n24788,
    n24789, n24790, n24791, n24792, n24793, n24794,
    n24795, n24796, n24797, n24798, n24799, n24800,
    n24801, n24802, n24803, n24804, n24805, n24806,
    n24807, n24808, n24809, n24810, n24811, n24812,
    n24813, n24814, n24815, n24816, n24817, n24818,
    n24819, n24820, n24821, n24822, n24823, n24824,
    n24825, n24826, n24827, n24828, n24829, n24830,
    n24831, n24832, n24833, n24834, n24835, n24836,
    n24837, n24838, n24839, n24840, n24841, n24842,
    n24843, n24844, n24845, n24846, n24847, n24848,
    n24849, n24850, n24851, n24852, n24853, n24854,
    n24855, n24856, n24857, n24858, n24859, n24860,
    n24861, n24862, n24863, n24864, n24865, n24866,
    n24867, n24868, n24869, n24870, n24871, n24872,
    n24873, n24874, n24875, n24876, n24877, n24878,
    n24879, n24880, n24881, n24882, n24883, n24884,
    n24885, n24886, n24887, n24888, n24889, n24890,
    n24891, n24892, n24893, n24894, n24895, n24896,
    n24897, n24898, n24899, n24900, n24901, n24902,
    n24903, n24904, n24905, n24906, n24907, n24908,
    n24909, n24910, n24911, n24912, n24913, n24914,
    n24915, n24916, n24917, n24918, n24919, n24920,
    n24921, n24922, n24923, n24924, n24925, n24926,
    n24927, n24928, n24929, n24930, n24931, n24932,
    n24933, n24934, n24935, n24936, n24937, n24938,
    n24939, n24940, n24941, n24942, n24943, n24944,
    n24945, n24946, n24947, n24948, n24949, n24950,
    n24951, n24952, n24953, n24954, n24955, n24956,
    n24957, n24958, n24959, n24960, n24961, n24962,
    n24963, n24964, n24965, n24966, n24967, n24968,
    n24969, n24970, n24971, n24972, n24973, n24974,
    n24975, n24976, n24977, n24978, n24979, n24980,
    n24981, n24982, n24983, n24984, n24985, n24986,
    n24987, n24988, n24989, n24990, n24991, n24992,
    n24993, n24994, n24995, n24996, n24997, n24998,
    n24999, n25000, n25001, n25002, n25003, n25004,
    n25005, n25006, n25007, n25008, n25009, n25010,
    n25011, n25012, n25013, n25014, n25015, n25016,
    n25017, n25018, n25019, n25020, n25021, n25022,
    n25023, n25024, n25025, n25026, n25027, n25028,
    n25029, n25030, n25031, n25032, n25033, n25034,
    n25035, n25036, n25037, n25038, n25039, n25040,
    n25041, n25042, n25043, n25044, n25045, n25046,
    n25047, n25048, n25049, n25050, n25051, n25052,
    n25053, n25054, n25055, n25056, n25057, n25058,
    n25059, n25060, n25061, n25062, n25063, n25064,
    n25065, n25066, n25067, n25068, n25069, n25070,
    n25071, n25072, n25073, n25074, n25075, n25076,
    n25077, n25078, n25079, n25080, n25081, n25082,
    n25083, n25084, n25085, n25086, n25087, n25088,
    n25089, n25090, n25091, n25092, n25093, n25094,
    n25095, n25096, n25097, n25098, n25099, n25100,
    n25101, n25102, n25103, n25104, n25105, n25106,
    n25107, n25108, n25109, n25110, n25111, n25112,
    n25113, n25114, n25115, n25116, n25117, n25118,
    n25119, n25120, n25121, n25122, n25123, n25124,
    n25125, n25126, n25127, n25128, n25129, n25130,
    n25131, n25132, n25133, n25134, n25135, n25136,
    n25137, n25138, n25139, n25140, n25141, n25142,
    n25143, n25144, n25145, n25146, n25147, n25148,
    n25149, n25150, n25151, n25152, n25153, n25154,
    n25155, n25156, n25157, n25158, n25159, n25160,
    n25161, n25162, n25163, n25164, n25165, n25166,
    n25167, n25168, n25169, n25170, n25171, n25172,
    n25173, n25174, n25175, n25176, n25177, n25178,
    n25179, n25180, n25181, n25182, n25183, n25184,
    n25185, n25186, n25187, n25188, n25189, n25190,
    n25191, n25192, n25193, n25194, n25195, n25196,
    n25197, n25198, n25199, n25200, n25201, n25202,
    n25203, n25204, n25205, n25206, n25207, n25208,
    n25209, n25210, n25211, n25212, n25213, n25214,
    n25215, n25216, n25217, n25218, n25219, n25220,
    n25221, n25222, n25223, n25224, n25225, n25226,
    n25227, n25228, n25229, n25230, n25231, n25232,
    n25233, n25234, n25235, n25236, n25237, n25238,
    n25239, n25240, n25241, n25242, n25243, n25244,
    n25245, n25246, n25247, n25248, n25249, n25250,
    n25251, n25252, n25253, n25254, n25255, n25256,
    n25257, n25258, n25259, n25260, n25261, n25262,
    n25263, n25264, n25265, n25266, n25267, n25268,
    n25269, n25270, n25271, n25272, n25273, n25274,
    n25275, n25276, n25277, n25278, n25279, n25280,
    n25281, n25282, n25283, n25284, n25285, n25286,
    n25287, n25288, n25289, n25290, n25291, n25292,
    n25293, n25294, n25295, n25296, n25297, n25298,
    n25299, n25300, n25301, n25302, n25303, n25304,
    n25305, n25306, n25307, n25308, n25309, n25310,
    n25311, n25312, n25313, n25314, n25315, n25316,
    n25317, n25318, n25319, n25320, n25321, n25322,
    n25323, n25324, n25325, n25326, n25327, n25328,
    n25329, n25330, n25331, n25332, n25333, n25334,
    n25335, n25336, n25337, n25338, n25339, n25340,
    n25341, n25342, n25343, n25344, n25345, n25346,
    n25347, n25348, n25349, n25350, n25351, n25352,
    n25353, n25354, n25355, n25356, n25357, n25358,
    n25359, n25360, n25361, n25362, n25364, n25365,
    n25366, n25367, n25368, n25369, n25370, n25371,
    n25372, n25373, n25374, n25375, n25376, n25377,
    n25378, n25379, n25380, n25381, n25382, n25383,
    n25384, n25385, n25386, n25387, n25388, n25389,
    n25390, n25391, n25392, n25393, n25394, n25395,
    n25396, n25397, n25398, n25399, n25400, n25401,
    n25402, n25403, n25404, n25405, n25406, n25407,
    n25408, n25409, n25410, n25411, n25412, n25413,
    n25414, n25415, n25416, n25417, n25418, n25419,
    n25420, n25421, n25422, n25423, n25424, n25425,
    n25426, n25427, n25428, n25429, n25430, n25431,
    n25432, n25433, n25434, n25435, n25436, n25437,
    n25438, n25439, n25440, n25441, n25442, n25443,
    n25444, n25445, n25446, n25447, n25448, n25449,
    n25450, n25451, n25452, n25453, n25454, n25455,
    n25456, n25457, n25458, n25459, n25460, n25461,
    n25462, n25463, n25464, n25465, n25466, n25467,
    n25468, n25469, n25470, n25471, n25472, n25473,
    n25474, n25475, n25476, n25477, n25478, n25479,
    n25480, n25481, n25482, n25483, n25484, n25485,
    n25486, n25487, n25488, n25489, n25490, n25491,
    n25492, n25493, n25494, n25495, n25496, n25497,
    n25498, n25499, n25500, n25501, n25502, n25503,
    n25504, n25505, n25506, n25507, n25508, n25509,
    n25510, n25511, n25512, n25513, n25514, n25515,
    n25516, n25517, n25518, n25519, n25520, n25521,
    n25522, n25523, n25524, n25525, n25526, n25527,
    n25528, n25529, n25530, n25531, n25532, n25533,
    n25534, n25535, n25536, n25537, n25538, n25539,
    n25540, n25541, n25542, n25543, n25544, n25545,
    n25546, n25547, n25548, n25549, n25550, n25551,
    n25552, n25553, n25554, n25555, n25556, n25557,
    n25558, n25559, n25560, n25561, n25562, n25563,
    n25564, n25565, n25566, n25567, n25568, n25569,
    n25570, n25571, n25572, n25573, n25574, n25575,
    n25576, n25577, n25578, n25579, n25580, n25581,
    n25582, n25583, n25584, n25585, n25586, n25587,
    n25588, n25589, n25590, n25591, n25592, n25593,
    n25594, n25595, n25596, n25597, n25598, n25599,
    n25600, n25601, n25602, n25603, n25604, n25605,
    n25606, n25607, n25608, n25609, n25610, n25611,
    n25612, n25613, n25614, n25615, n25616, n25617,
    n25618, n25619, n25620, n25621, n25622, n25624,
    n25625, n25626, n25627, n25628, n25629, n25630,
    n25631, n25632, n25633, n25634, n25635, n25636,
    n25637, n25638, n25639, n25640, n25641, n25642,
    n25643, n25644, n25645, n25646, n25647, n25648,
    n25649, n25650, n25651, n25652, n25653, n25654,
    n25655, n25656, n25657, n25658, n25659, n25660,
    n25661, n25662, n25663, n25664, n25665, n25666,
    n25667, n25668, n25669, n25670, n25671, n25672,
    n25673, n25674, n25675, n25676, n25677, n25678,
    n25679, n25680, n25681, n25682, n25683, n25684,
    n25685, n25686, n25687, n25688, n25689, n25690,
    n25691, n25692, n25693, n25694, n25695, n25696,
    n25697, n25698, n25699, n25700, n25701, n25702,
    n25703, n25704, n25705, n25706, n25707, n25708,
    n25709, n25710, n25711, n25712, n25713, n25714,
    n25715, n25716, n25717, n25718, n25719, n25720,
    n25721, n25722, n25723, n25724, n25725, n25726,
    n25727, n25728, n25729, n25730, n25731, n25732,
    n25733, n25734, n25735, n25736, n25737, n25738,
    n25739, n25740, n25741, n25742, n25743, n25744,
    n25745, n25746, n25747, n25748, n25749, n25750,
    n25751, n25752, n25753, n25754, n25755, n25756,
    n25757, n25758, n25759, n25760, n25761, n25762,
    n25763, n25764, n25765, n25766, n25767, n25768,
    n25769, n25770, n25771, n25772, n25773, n25774,
    n25775, n25776, n25777, n25778, n25779, n25780,
    n25781, n25782, n25783, n25784, n25785, n25786,
    n25787, n25788, n25789, n25790, n25791, n25792,
    n25793, n25794, n25795, n25796, n25797, n25798,
    n25799, n25800, n25801, n25802, n25803, n25804,
    n25805, n25806, n25807, n25808, n25809, n25810,
    n25811, n25812, n25813, n25814, n25815, n25816,
    n25817, n25818, n25819, n25820, n25821, n25822,
    n25823, n25824, n25825, n25826, n25827, n25828,
    n25829, n25830, n25831, n25832, n25833, n25834,
    n25835, n25836, n25837, n25838, n25839, n25840,
    n25841, n25842, n25843, n25844, n25845, n25846,
    n25847, n25848, n25849, n25850, n25851, n25852,
    n25853, n25854, n25855, n25856, n25857, n25858,
    n25859, n25860, n25861, n25862, n25863, n25864,
    n25865, n25866, n25867, n25868, n25869, n25870,
    n25871, n25872, n25873, n25874, n25875, n25876,
    n25878, n25879, n25880, n25881, n25882, n25883,
    n25884, n25885, n25886, n25887, n25888, n25889,
    n25890, n25891, n25892, n25893, n25894, n25895,
    n25896, n25897, n25898, n25899, n25900, n25901,
    n25902, n25903, n25904, n25905, n25906, n25907,
    n25908, n25909, n25910, n25911, n25912, n25913,
    n25914, n25915, n25916, n25917, n25918, n25919,
    n25920, n25921, n25922, n25923, n25924, n25925,
    n25926, n25927, n25928, n25929, n25930, n25931,
    n25932, n25933, n25934, n25935, n25936, n25937,
    n25938, n25939, n25940, n25941, n25942, n25943,
    n25944, n25945, n25946, n25947, n25948, n25949,
    n25950, n25951, n25952, n25953, n25954, n25955,
    n25956, n25957, n25958, n25959, n25960, n25961,
    n25962, n25963, n25964, n25965, n25966, n25967,
    n25968, n25969, n25970, n25971, n25972, n25973,
    n25974, n25975, n25976, n25977, n25978, n25979,
    n25980, n25981, n25982, n25983, n25984, n25985,
    n25986, n25987, n25988, n25989, n25990, n25991,
    n25992, n25993, n25994, n25995, n25996, n25997,
    n25998, n25999, n26000, n26001, n26002, n26003,
    n26004, n26005, n26006, n26007, n26008, n26009,
    n26010, n26011, n26012, n26013, n26014, n26015,
    n26016, n26017, n26018, n26019, n26020, n26021,
    n26022, n26023, n26024, n26025, n26026, n26027,
    n26028, n26029, n26030, n26031, n26032, n26033,
    n26034, n26035, n26036, n26037, n26038, n26039,
    n26040, n26041, n26042, n26043, n26044, n26045,
    n26046, n26047, n26048, n26049, n26050, n26051,
    n26052, n26053, n26054, n26055, n26056, n26057,
    n26058, n26059, n26060, n26061, n26062, n26063,
    n26064, n26065, n26066, n26067, n26068, n26069,
    n26070, n26071, n26072, n26073, n26074, n26075,
    n26076, n26077, n26078, n26079, n26080, n26081,
    n26082, n26083, n26084, n26085, n26086, n26087,
    n26088, n26089, n26090, n26091, n26092, n26093,
    n26094, n26095, n26096, n26097, n26098, n26099,
    n26100, n26101, n26102, n26103, n26104, n26105,
    n26106, n26107, n26108, n26109, n26110, n26111,
    n26112, n26113, n26114, n26115, n26116, n26117,
    n26119, n26120, n26121, n26122, n26123, n26124,
    n26125, n26126, n26127, n26128, n26129, n26130,
    n26131, n26132, n26133, n26134, n26135, n26136,
    n26137, n26138, n26139, n26140, n26141, n26142,
    n26143, n26144, n26145, n26146, n26147, n26148,
    n26149, n26150, n26151, n26152, n26153, n26154,
    n26155, n26156, n26157, n26158, n26159, n26160,
    n26161, n26162, n26163, n26164, n26165, n26166,
    n26167, n26168, n26169, n26170, n26171, n26172,
    n26173, n26174, n26175, n26176, n26177, n26178,
    n26179, n26180, n26181, n26182, n26183, n26184,
    n26185, n26186, n26187, n26188, n26189, n26190,
    n26191, n26192, n26193, n26194, n26195, n26196,
    n26197, n26198, n26199, n26200, n26201, n26202,
    n26203, n26204, n26205, n26206, n26207, n26208,
    n26209, n26210, n26211, n26212, n26213, n26214,
    n26215, n26216, n26217, n26218, n26219, n26220,
    n26221, n26222, n26223, n26224, n26225, n26226,
    n26227, n26228, n26229, n26230, n26231, n26232,
    n26233, n26234, n26235, n26236, n26237, n26238,
    n26239, n26240, n26241, n26242, n26243, n26244,
    n26245, n26246, n26247, n26248, n26249, n26250,
    n26251, n26252, n26253, n26254, n26255, n26256,
    n26257, n26258, n26259, n26260, n26261, n26262,
    n26263, n26264, n26265, n26266, n26267, n26268,
    n26269, n26270, n26271, n26272, n26273, n26274,
    n26275, n26276, n26277, n26278, n26279, n26280,
    n26281, n26282, n26283, n26284, n26285, n26286,
    n26287, n26288, n26289, n26290, n26291, n26292,
    n26293, n26294, n26295, n26296, n26297, n26298,
    n26299, n26300, n26301, n26302, n26303, n26304,
    n26305, n26306, n26307, n26308, n26309, n26310,
    n26311, n26312, n26313, n26314, n26315, n26316,
    n26317, n26318, n26319, n26320, n26321, n26322,
    n26323, n26324, n26325, n26326, n26327, n26328,
    n26329, n26330, n26331, n26332, n26333, n26334,
    n26335, n26336, n26337, n26338, n26339, n26340,
    n26341, n26342, n26343, n26344, n26345, n26346,
    n26347, n26348, n26349, n26350, n26351, n26352,
    n26353, n26354, n26355, n26356, n26357, n26358,
    n26359, n26360, n26361, n26362, n26363, n26364,
    n26366, n26367, n26368, n26369, n26370, n26371,
    n26372, n26373, n26374, n26375, n26376, n26377,
    n26378, n26379, n26380, n26381, n26382, n26383,
    n26384, n26385, n26386, n26387, n26388, n26389,
    n26390, n26391, n26392, n26393, n26394, n26395,
    n26396, n26397, n26398, n26399, n26400, n26401,
    n26402, n26403, n26404, n26405, n26406, n26407,
    n26408, n26409, n26410, n26411, n26412, n26413,
    n26414, n26415, n26416, n26417, n26418, n26419,
    n26420, n26421, n26422, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26431,
    n26432, n26433, n26434, n26435, n26436, n26437,
    n26438, n26439, n26440, n26441, n26442, n26443,
    n26444, n26445, n26446, n26447, n26448, n26449,
    n26450, n26451, n26452, n26453, n26454, n26455,
    n26456, n26457, n26458, n26459, n26460, n26461,
    n26462, n26463, n26464, n26465, n26466, n26467,
    n26468, n26469, n26470, n26471, n26472, n26473,
    n26474, n26475, n26476, n26477, n26478, n26479,
    n26480, n26481, n26482, n26483, n26484, n26485,
    n26486, n26487, n26488, n26489, n26490, n26491,
    n26492, n26493, n26494, n26495, n26496, n26497,
    n26498, n26499, n26500, n26501, n26502, n26503,
    n26504, n26505, n26506, n26507, n26508, n26509,
    n26510, n26511, n26512, n26513, n26514, n26515,
    n26516, n26517, n26518, n26519, n26520, n26521,
    n26522, n26523, n26524, n26525, n26526, n26527,
    n26528, n26529, n26530, n26531, n26532, n26533,
    n26534, n26535, n26536, n26537, n26538, n26539,
    n26540, n26541, n26542, n26543, n26544, n26545,
    n26546, n26547, n26548, n26549, n26550, n26551,
    n26552, n26553, n26554, n26555, n26556, n26557,
    n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26571, n26572, n26573, n26574, n26575,
    n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587,
    n26588, n26589, n26590, n26591, n26592, n26594,
    n26595, n26596, n26597, n26598, n26599, n26600,
    n26601, n26602, n26603, n26604, n26605, n26606,
    n26607, n26608, n26609, n26610, n26611, n26612,
    n26613, n26614, n26615, n26616, n26617, n26618,
    n26619, n26620, n26621, n26622, n26623, n26624,
    n26625, n26626, n26627, n26628, n26629, n26630,
    n26631, n26632, n26633, n26634, n26635, n26636,
    n26637, n26638, n26639, n26640, n26641, n26642,
    n26643, n26644, n26645, n26646, n26647, n26648,
    n26649, n26650, n26651, n26652, n26653, n26654,
    n26655, n26656, n26657, n26658, n26659, n26660,
    n26661, n26662, n26663, n26664, n26665, n26666,
    n26667, n26668, n26669, n26670, n26671, n26672,
    n26673, n26674, n26675, n26676, n26677, n26678,
    n26679, n26680, n26681, n26682, n26683, n26684,
    n26685, n26686, n26687, n26688, n26689, n26690,
    n26691, n26692, n26693, n26694, n26695, n26696,
    n26697, n26698, n26699, n26700, n26701, n26702,
    n26703, n26704, n26705, n26706, n26707, n26708,
    n26709, n26710, n26711, n26712, n26713, n26714,
    n26715, n26716, n26717, n26718, n26719, n26720,
    n26721, n26722, n26723, n26724, n26725, n26726,
    n26727, n26728, n26729, n26730, n26731, n26732,
    n26733, n26734, n26735, n26736, n26737, n26738,
    n26739, n26740, n26741, n26742, n26743, n26744,
    n26745, n26746, n26747, n26748, n26749, n26750,
    n26751, n26752, n26753, n26754, n26755, n26756,
    n26757, n26758, n26759, n26760, n26761, n26762,
    n26763, n26764, n26765, n26766, n26767, n26768,
    n26769, n26770, n26771, n26772, n26773, n26774,
    n26775, n26776, n26777, n26778, n26779, n26780,
    n26781, n26782, n26783, n26784, n26785, n26786,
    n26787, n26788, n26789, n26790, n26791, n26792,
    n26793, n26794, n26795, n26796, n26797, n26798,
    n26799, n26800, n26801, n26802, n26803, n26804,
    n26805, n26806, n26807, n26808, n26809, n26810,
    n26811, n26813, n26814, n26815, n26816, n26817,
    n26818, n26819, n26820, n26821, n26822, n26823,
    n26824, n26825, n26826, n26827, n26828, n26829,
    n26830, n26831, n26832, n26833, n26834, n26835,
    n26836, n26837, n26838, n26839, n26840, n26841,
    n26842, n26843, n26844, n26845, n26846, n26847,
    n26848, n26849, n26850, n26851, n26852, n26853,
    n26854, n26855, n26856, n26857, n26858, n26859,
    n26860, n26861, n26862, n26863, n26864, n26865,
    n26866, n26867, n26868, n26869, n26870, n26871,
    n26872, n26873, n26874, n26875, n26876, n26877,
    n26878, n26879, n26880, n26881, n26882, n26883,
    n26884, n26885, n26886, n26887, n26888, n26889,
    n26890, n26891, n26892, n26893, n26894, n26895,
    n26896, n26897, n26898, n26899, n26900, n26901,
    n26902, n26903, n26904, n26905, n26906, n26907,
    n26908, n26909, n26910, n26911, n26912, n26913,
    n26914, n26915, n26916, n26917, n26918, n26919,
    n26920, n26921, n26922, n26923, n26924, n26925,
    n26926, n26927, n26928, n26929, n26930, n26931,
    n26932, n26933, n26934, n26935, n26936, n26937,
    n26938, n26939, n26940, n26941, n26942, n26943,
    n26944, n26945, n26946, n26947, n26948, n26949,
    n26950, n26951, n26952, n26953, n26954, n26955,
    n26956, n26957, n26958, n26959, n26960, n26961,
    n26962, n26963, n26964, n26965, n26966, n26967,
    n26968, n26969, n26970, n26971, n26972, n26973,
    n26974, n26975, n26976, n26977, n26978, n26979,
    n26980, n26981, n26982, n26983, n26984, n26985,
    n26986, n26987, n26988, n26989, n26990, n26991,
    n26992, n26993, n26994, n26995, n26996, n26997,
    n26998, n26999, n27000, n27001, n27002, n27003,
    n27004, n27005, n27006, n27007, n27008, n27009,
    n27010, n27011, n27012, n27014, n27015, n27016,
    n27017, n27018, n27019, n27020, n27021, n27022,
    n27023, n27024, n27025, n27026, n27027, n27028,
    n27029, n27030, n27031, n27032, n27033, n27034,
    n27035, n27036, n27037, n27038, n27039, n27040,
    n27041, n27042, n27043, n27044, n27045, n27046,
    n27047, n27048, n27049, n27050, n27051, n27052,
    n27053, n27054, n27055, n27056, n27057, n27058,
    n27059, n27060, n27061, n27062, n27063, n27064,
    n27065, n27066, n27067, n27068, n27069, n27070,
    n27071, n27072, n27073, n27074, n27075, n27076,
    n27077, n27078, n27079, n27080, n27081, n27082,
    n27083, n27084, n27085, n27086, n27087, n27088,
    n27089, n27090, n27091, n27092, n27093, n27094,
    n27095, n27096, n27097, n27098, n27099, n27100,
    n27101, n27102, n27103, n27104, n27105, n27106,
    n27107, n27108, n27109, n27110, n27111, n27112,
    n27113, n27114, n27115, n27116, n27117, n27118,
    n27119, n27120, n27121, n27122, n27123, n27124,
    n27125, n27126, n27127, n27128, n27129, n27130,
    n27131, n27132, n27133, n27134, n27135, n27136,
    n27137, n27138, n27139, n27140, n27141, n27142,
    n27143, n27144, n27145, n27146, n27147, n27148,
    n27149, n27150, n27151, n27152, n27153, n27154,
    n27155, n27156, n27157, n27158, n27159, n27160,
    n27161, n27162, n27163, n27164, n27165, n27166,
    n27167, n27168, n27169, n27170, n27171, n27172,
    n27173, n27174, n27175, n27176, n27177, n27178,
    n27179, n27180, n27181, n27182, n27183, n27184,
    n27185, n27186, n27187, n27188, n27189, n27190,
    n27191, n27192, n27193, n27194, n27195, n27196,
    n27197, n27198, n27199, n27200, n27201, n27202,
    n27203, n27204, n27205, n27206, n27207, n27208,
    n27209, n27210, n27211, n27212, n27213, n27214,
    n27215, n27216, n27217, n27218, n27219, n27220,
    n27222, n27223, n27224, n27225, n27226, n27227,
    n27228, n27229, n27230, n27231, n27232, n27233,
    n27234, n27235, n27236, n27237, n27238, n27239,
    n27240, n27241, n27242, n27243, n27244, n27245,
    n27246, n27247, n27248, n27249, n27250, n27251,
    n27252, n27253, n27254, n27255, n27256, n27257,
    n27258, n27259, n27260, n27261, n27262, n27263,
    n27264, n27265, n27266, n27267, n27268, n27269,
    n27270, n27271, n27272, n27273, n27274, n27275,
    n27276, n27277, n27278, n27279, n27280, n27281,
    n27282, n27283, n27284, n27285, n27286, n27287,
    n27288, n27289, n27290, n27291, n27292, n27293,
    n27294, n27295, n27296, n27297, n27298, n27299,
    n27300, n27301, n27302, n27303, n27304, n27305,
    n27306, n27307, n27308, n27309, n27310, n27311,
    n27312, n27313, n27314, n27315, n27316, n27317,
    n27318, n27319, n27320, n27321, n27322, n27323,
    n27324, n27325, n27326, n27327, n27328, n27329,
    n27330, n27331, n27332, n27333, n27334, n27335,
    n27336, n27337, n27338, n27339, n27340, n27341,
    n27342, n27343, n27344, n27345, n27346, n27347,
    n27348, n27349, n27350, n27351, n27352, n27353,
    n27354, n27355, n27356, n27357, n27358, n27359,
    n27360, n27361, n27362, n27363, n27364, n27365,
    n27366, n27367, n27368, n27369, n27370, n27371,
    n27372, n27373, n27374, n27375, n27376, n27377,
    n27378, n27379, n27380, n27381, n27382, n27383,
    n27384, n27385, n27386, n27387, n27388, n27389,
    n27390, n27391, n27392, n27393, n27394, n27395,
    n27396, n27397, n27398, n27399, n27400, n27401,
    n27402, n27403, n27404, n27405, n27406, n27407,
    n27408, n27409, n27410, n27411, n27412, n27413,
    n27414, n27415, n27416, n27417, n27418, n27419,
    n27420, n27421, n27423, n27424, n27425, n27426,
    n27427, n27428, n27429, n27430, n27431, n27432,
    n27433, n27434, n27435, n27436, n27437, n27438,
    n27439, n27440, n27441, n27442, n27443, n27444,
    n27445, n27446, n27447, n27448, n27449, n27450,
    n27451, n27452, n27453, n27454, n27455, n27456,
    n27457, n27458, n27459, n27460, n27461, n27462,
    n27463, n27464, n27465, n27466, n27467, n27468,
    n27469, n27470, n27471, n27472, n27473, n27474,
    n27475, n27476, n27477, n27478, n27479, n27480,
    n27481, n27482, n27483, n27484, n27485, n27486,
    n27487, n27488, n27489, n27490, n27491, n27492,
    n27493, n27494, n27495, n27496, n27497, n27498,
    n27499, n27500, n27501, n27502, n27503, n27504,
    n27505, n27506, n27507, n27508, n27509, n27510,
    n27511, n27512, n27513, n27514, n27515, n27516,
    n27517, n27518, n27519, n27520, n27521, n27522,
    n27523, n27524, n27525, n27526, n27527, n27528,
    n27529, n27530, n27531, n27532, n27533, n27534,
    n27535, n27536, n27537, n27538, n27539, n27540,
    n27541, n27542, n27543, n27544, n27545, n27546,
    n27547, n27548, n27549, n27550, n27551, n27552,
    n27553, n27554, n27555, n27556, n27557, n27558,
    n27559, n27560, n27561, n27562, n27563, n27564,
    n27565, n27566, n27567, n27568, n27569, n27570,
    n27571, n27572, n27573, n27574, n27575, n27576,
    n27577, n27578, n27579, n27580, n27581, n27582,
    n27583, n27584, n27585, n27586, n27587, n27588,
    n27589, n27590, n27591, n27592, n27593, n27594,
    n27595, n27596, n27597, n27598, n27599, n27600,
    n27601, n27602, n27603, n27604, n27605, n27606,
    n27607, n27608, n27609, n27610, n27611, n27612,
    n27613, n27614, n27615, n27616, n27618, n27619,
    n27620, n27621, n27622, n27623, n27624, n27625,
    n27626, n27627, n27628, n27629, n27630, n27631,
    n27632, n27633, n27634, n27635, n27636, n27637,
    n27638, n27639, n27640, n27641, n27642, n27643,
    n27644, n27645, n27646, n27647, n27648, n27649,
    n27650, n27651, n27652, n27653, n27654, n27655,
    n27656, n27657, n27658, n27659, n27660, n27661,
    n27662, n27663, n27664, n27665, n27666, n27667,
    n27668, n27669, n27670, n27671, n27672, n27673,
    n27674, n27675, n27676, n27677, n27678, n27679,
    n27680, n27681, n27682, n27683, n27684, n27685,
    n27686, n27687, n27688, n27689, n27690, n27691,
    n27692, n27693, n27694, n27695, n27696, n27697,
    n27698, n27699, n27700, n27701, n27702, n27703,
    n27704, n27705, n27706, n27707, n27708, n27709,
    n27710, n27711, n27712, n27713, n27714, n27715,
    n27716, n27717, n27718, n27719, n27720, n27721,
    n27722, n27723, n27724, n27725, n27726, n27727,
    n27728, n27729, n27730, n27731, n27732, n27733,
    n27734, n27735, n27736, n27737, n27738, n27739,
    n27740, n27741, n27742, n27743, n27744, n27745,
    n27746, n27747, n27748, n27749, n27750, n27751,
    n27752, n27753, n27754, n27755, n27756, n27757,
    n27758, n27759, n27760, n27761, n27762, n27763,
    n27764, n27765, n27766, n27767, n27768, n27769,
    n27770, n27771, n27772, n27773, n27774, n27775,
    n27776, n27777, n27778, n27779, n27780, n27781,
    n27782, n27783, n27784, n27785, n27786, n27787,
    n27788, n27789, n27790, n27791, n27792, n27793,
    n27794, n27795, n27796, n27797, n27798, n27799,
    n27800, n27801, n27802, n27803, n27804, n27805,
    n27806, n27807, n27808, n27809, n27810, n27811,
    n27812, n27813, n27815, n27816, n27817, n27818,
    n27819, n27820, n27821, n27822, n27823, n27824,
    n27825, n27826, n27827, n27828, n27829, n27830,
    n27831, n27832, n27833, n27834, n27835, n27836,
    n27837, n27838, n27839, n27840, n27841, n27842,
    n27843, n27844, n27845, n27846, n27847, n27848,
    n27849, n27850, n27851, n27852, n27853, n27854,
    n27855, n27856, n27857, n27858, n27859, n27860,
    n27861, n27862, n27863, n27864, n27865, n27866,
    n27867, n27868, n27869, n27870, n27871, n27872,
    n27873, n27874, n27875, n27876, n27877, n27878,
    n27879, n27880, n27881, n27882, n27883, n27884,
    n27885, n27886, n27887, n27888, n27889, n27890,
    n27891, n27892, n27893, n27894, n27895, n27896,
    n27897, n27898, n27899, n27900, n27901, n27902,
    n27903, n27904, n27905, n27906, n27907, n27908,
    n27909, n27910, n27911, n27912, n27913, n27914,
    n27915, n27916, n27917, n27918, n27919, n27920,
    n27921, n27922, n27923, n27924, n27925, n27926,
    n27927, n27928, n27929, n27930, n27931, n27932,
    n27933, n27934, n27935, n27936, n27937, n27938,
    n27939, n27940, n27941, n27942, n27943, n27944,
    n27945, n27946, n27947, n27948, n27949, n27950,
    n27951, n27952, n27953, n27954, n27955, n27956,
    n27957, n27958, n27959, n27960, n27961, n27962,
    n27963, n27964, n27965, n27966, n27967, n27968,
    n27969, n27970, n27971, n27972, n27973, n27974,
    n27975, n27976, n27977, n27978, n27979, n27980,
    n27981, n27982, n27983, n27984, n27985, n27986,
    n27987, n27988, n27989, n27990, n27991, n27992,
    n27993, n27994, n27995, n27996, n27997, n27998,
    n27999, n28000, n28001, n28002, n28003, n28004,
    n28005, n28006, n28007, n28008, n28009, n28010,
    n28011, n28012, n28014, n28015, n28016, n28017,
    n28018, n28019, n28020, n28021, n28022, n28023,
    n28024, n28025, n28026, n28027, n28028, n28029,
    n28030, n28031, n28032, n28033, n28034, n28035,
    n28036, n28037, n28038, n28039, n28040, n28041,
    n28042, n28043, n28044, n28045, n28046, n28047,
    n28048, n28049, n28050, n28051, n28052, n28053,
    n28054, n28055, n28056, n28057, n28058, n28059,
    n28060, n28061, n28062, n28063, n28064, n28065,
    n28066, n28067, n28068, n28069, n28070, n28071,
    n28072, n28073, n28074, n28075, n28076, n28077,
    n28078, n28079, n28080, n28081, n28082, n28083,
    n28084, n28085, n28086, n28087, n28088, n28089,
    n28090, n28091, n28092, n28093, n28094, n28095,
    n28096, n28097, n28098, n28099, n28100, n28101,
    n28102, n28103, n28104, n28105, n28106, n28107,
    n28108, n28109, n28110, n28111, n28112, n28113,
    n28114, n28115, n28116, n28117, n28118, n28119,
    n28120, n28121, n28122, n28123, n28124, n28125,
    n28126, n28127, n28128, n28129, n28130, n28131,
    n28132, n28133, n28134, n28135, n28136, n28137,
    n28138, n28139, n28140, n28141, n28142, n28143,
    n28144, n28145, n28146, n28147, n28148, n28149,
    n28150, n28151, n28152, n28153, n28154, n28155,
    n28156, n28157, n28158, n28159, n28160, n28161,
    n28162, n28163, n28164, n28165, n28166, n28167,
    n28168, n28169, n28170, n28171, n28172, n28173,
    n28174, n28175, n28176, n28177, n28178, n28179,
    n28180, n28181, n28182, n28183, n28184, n28185,
    n28186, n28187, n28188, n28190, n28191, n28192,
    n28193, n28194, n28195, n28196, n28197, n28198,
    n28199, n28200, n28201, n28202, n28203, n28204,
    n28205, n28206, n28207, n28208, n28209, n28210,
    n28211, n28212, n28213, n28214, n28215, n28216,
    n28217, n28218, n28219, n28220, n28221, n28222,
    n28223, n28224, n28225, n28226, n28227, n28228,
    n28229, n28230, n28231, n28232, n28233, n28234,
    n28235, n28236, n28237, n28238, n28239, n28240,
    n28241, n28242, n28243, n28244, n28245, n28246,
    n28247, n28248, n28249, n28250, n28251, n28252,
    n28253, n28254, n28255, n28256, n28257, n28258,
    n28259, n28260, n28261, n28262, n28263, n28264,
    n28265, n28266, n28267, n28268, n28269, n28270,
    n28271, n28272, n28273, n28274, n28275, n28276,
    n28277, n28278, n28279, n28280, n28281, n28282,
    n28283, n28284, n28285, n28286, n28287, n28288,
    n28289, n28290, n28291, n28292, n28293, n28294,
    n28295, n28296, n28297, n28298, n28299, n28300,
    n28301, n28302, n28303, n28304, n28305, n28306,
    n28307, n28308, n28309, n28310, n28311, n28312,
    n28313, n28314, n28315, n28316, n28317, n28318,
    n28319, n28320, n28321, n28322, n28323, n28324,
    n28325, n28326, n28327, n28328, n28329, n28330,
    n28331, n28332, n28333, n28334, n28335, n28336,
    n28337, n28338, n28339, n28340, n28341, n28342,
    n28343, n28344, n28345, n28346, n28347, n28348,
    n28349, n28350, n28351, n28352, n28354, n28355,
    n28356, n28357, n28358, n28359, n28360, n28361,
    n28362, n28363, n28364, n28365, n28366, n28367,
    n28368, n28369, n28370, n28371, n28372, n28373,
    n28374, n28375, n28376, n28377, n28378, n28379,
    n28380, n28381, n28382, n28383, n28384, n28385,
    n28386, n28387, n28388, n28389, n28390, n28391,
    n28392, n28393, n28394, n28395, n28396, n28397,
    n28398, n28399, n28400, n28401, n28402, n28403,
    n28404, n28405, n28406, n28407, n28408, n28409,
    n28410, n28411, n28412, n28413, n28414, n28415,
    n28416, n28417, n28418, n28419, n28420, n28421,
    n28422, n28423, n28424, n28425, n28426, n28427,
    n28428, n28429, n28430, n28431, n28432, n28433,
    n28434, n28435, n28436, n28437, n28438, n28439,
    n28440, n28441, n28442, n28443, n28444, n28445,
    n28446, n28447, n28448, n28449, n28450, n28451,
    n28452, n28453, n28454, n28455, n28456, n28457,
    n28458, n28459, n28460, n28461, n28462, n28463,
    n28464, n28465, n28466, n28467, n28468, n28469,
    n28470, n28471, n28472, n28473, n28474, n28475,
    n28476, n28477, n28478, n28479, n28480, n28481,
    n28482, n28483, n28484, n28485, n28486, n28487,
    n28488, n28489, n28490, n28491, n28492, n28493,
    n28494, n28495, n28496, n28497, n28498, n28499,
    n28500, n28501, n28502, n28503, n28504, n28505,
    n28506, n28507, n28508, n28509, n28510, n28511,
    n28512, n28513, n28514, n28515, n28516, n28518,
    n28519, n28520, n28521, n28522, n28523, n28524,
    n28525, n28526, n28527, n28528, n28529, n28530,
    n28531, n28532, n28533, n28534, n28535, n28536,
    n28537, n28538, n28539, n28540, n28541, n28542,
    n28543, n28544, n28545, n28546, n28547, n28548,
    n28549, n28550, n28551, n28552, n28553, n28554,
    n28555, n28556, n28557, n28558, n28559, n28560,
    n28561, n28562, n28563, n28564, n28565, n28566,
    n28567, n28568, n28569, n28570, n28571, n28572,
    n28573, n28574, n28575, n28576, n28577, n28578,
    n28579, n28580, n28581, n28582, n28583, n28584,
    n28585, n28586, n28587, n28588, n28589, n28590,
    n28591, n28592, n28593, n28594, n28595, n28596,
    n28597, n28598, n28599, n28600, n28601, n28602,
    n28603, n28604, n28605, n28606, n28607, n28608,
    n28609, n28610, n28611, n28612, n28613, n28614,
    n28615, n28616, n28617, n28618, n28619, n28620,
    n28621, n28622, n28623, n28624, n28625, n28626,
    n28627, n28628, n28629, n28630, n28631, n28632,
    n28633, n28634, n28635, n28636, n28637, n28638,
    n28639, n28640, n28641, n28642, n28643, n28644,
    n28645, n28646, n28647, n28648, n28649, n28650,
    n28651, n28652, n28653, n28654, n28655, n28656,
    n28657, n28658, n28659, n28660, n28661, n28662,
    n28663, n28664, n28665, n28666, n28667, n28668,
    n28669, n28670, n28671, n28672, n28673, n28674,
    n28675, n28677, n28678, n28679, n28680, n28681,
    n28682, n28683, n28684, n28685, n28686, n28687,
    n28688, n28689, n28690, n28691, n28692, n28693,
    n28694, n28695, n28696, n28697, n28698, n28699,
    n28700, n28701, n28702, n28703, n28704, n28705,
    n28706, n28707, n28708, n28709, n28710, n28711,
    n28712, n28713, n28714, n28715, n28716, n28717,
    n28718, n28719, n28720, n28721, n28722, n28723,
    n28724, n28725, n28726, n28727, n28728, n28729,
    n28730, n28731, n28732, n28733, n28734, n28735,
    n28736, n28737, n28738, n28739, n28740, n28741,
    n28742, n28743, n28744, n28745, n28746, n28747,
    n28748, n28749, n28750, n28751, n28752, n28753,
    n28754, n28755, n28756, n28757, n28758, n28759,
    n28760, n28761, n28762, n28763, n28764, n28765,
    n28766, n28767, n28768, n28769, n28770, n28771,
    n28772, n28773, n28774, n28775, n28776, n28777,
    n28778, n28779, n28780, n28781, n28782, n28783,
    n28784, n28785, n28786, n28787, n28788, n28789,
    n28790, n28791, n28792, n28793, n28794, n28795,
    n28796, n28797, n28798, n28799, n28800, n28801,
    n28802, n28803, n28804, n28805, n28806, n28807,
    n28808, n28809, n28810, n28811, n28812, n28813,
    n28814, n28815, n28816, n28817, n28818, n28819,
    n28820, n28821, n28822, n28823, n28824, n28826,
    n28827, n28828, n28829, n28830, n28831, n28832,
    n28833, n28834, n28835, n28836, n28837, n28838,
    n28839, n28840, n28841, n28842, n28843, n28844,
    n28845, n28846, n28847, n28848, n28849, n28850,
    n28851, n28852, n28853, n28854, n28855, n28856,
    n28857, n28858, n28859, n28860, n28861, n28862,
    n28863, n28864, n28865, n28866, n28867, n28868,
    n28869, n28870, n28871, n28872, n28873, n28874,
    n28875, n28876, n28877, n28878, n28879, n28880,
    n28881, n28882, n28883, n28884, n28885, n28886,
    n28887, n28888, n28889, n28890, n28891, n28892,
    n28893, n28894, n28895, n28896, n28897, n28898,
    n28899, n28900, n28901, n28902, n28903, n28904,
    n28905, n28906, n28907, n28908, n28909, n28910,
    n28911, n28912, n28913, n28914, n28915, n28916,
    n28917, n28918, n28919, n28920, n28921, n28922,
    n28923, n28924, n28925, n28926, n28927, n28928,
    n28929, n28930, n28931, n28932, n28933, n28934,
    n28935, n28936, n28937, n28938, n28939, n28940,
    n28941, n28942, n28943, n28944, n28945, n28946,
    n28947, n28948, n28949, n28950, n28951, n28952,
    n28953, n28954, n28955, n28956, n28957, n28958,
    n28959, n28960, n28961, n28962, n28963, n28964,
    n28965, n28966, n28967, n28968, n28969, n28970,
    n28971, n28973, n28974, n28975, n28976, n28977,
    n28978, n28979, n28980, n28981, n28982, n28983,
    n28984, n28985, n28986, n28987, n28988, n28989,
    n28990, n28991, n28992, n28993, n28994, n28995,
    n28996, n28997, n28998, n28999, n29000, n29001,
    n29002, n29003, n29004, n29005, n29006, n29007,
    n29008, n29009, n29010, n29011, n29012, n29013,
    n29014, n29015, n29016, n29017, n29018, n29019,
    n29020, n29021, n29022, n29023, n29024, n29025,
    n29026, n29027, n29028, n29029, n29030, n29031,
    n29032, n29033, n29034, n29035, n29036, n29037,
    n29038, n29039, n29040, n29041, n29042, n29043,
    n29044, n29045, n29046, n29047, n29048, n29049,
    n29050, n29051, n29052, n29053, n29054, n29055,
    n29056, n29057, n29058, n29059, n29060, n29061,
    n29062, n29063, n29064, n29065, n29066, n29067,
    n29068, n29069, n29070, n29071, n29072, n29073,
    n29074, n29075, n29076, n29077, n29078, n29079,
    n29080, n29081, n29082, n29083, n29084, n29085,
    n29086, n29087, n29088, n29089, n29090, n29091,
    n29092, n29093, n29094, n29095, n29096, n29097,
    n29098, n29099, n29100, n29101, n29102, n29103,
    n29104, n29105, n29106, n29107, n29109, n29110,
    n29111, n29112, n29113, n29114, n29115, n29116,
    n29117, n29118, n29119, n29120, n29121, n29122,
    n29123, n29124, n29125, n29126, n29127, n29128,
    n29129, n29130, n29131, n29132, n29133, n29134,
    n29135, n29136, n29137, n29138, n29139, n29140,
    n29141, n29142, n29143, n29144, n29145, n29146,
    n29147, n29148, n29149, n29150, n29151, n29152,
    n29153, n29154, n29155, n29156, n29157, n29158,
    n29159, n29160, n29161, n29162, n29163, n29164,
    n29165, n29166, n29167, n29168, n29169, n29170,
    n29171, n29172, n29173, n29174, n29175, n29176,
    n29177, n29178, n29179, n29180, n29181, n29182,
    n29183, n29184, n29185, n29186, n29187, n29188,
    n29189, n29190, n29191, n29192, n29193, n29194,
    n29195, n29196, n29197, n29198, n29199, n29200,
    n29201, n29202, n29203, n29204, n29205, n29206,
    n29207, n29208, n29209, n29210, n29211, n29212,
    n29213, n29214, n29215, n29216, n29217, n29218,
    n29219, n29220, n29221, n29222, n29223, n29224,
    n29225, n29226, n29227, n29228, n29229, n29230,
    n29231, n29232, n29233, n29234, n29235, n29236,
    n29238, n29239, n29240, n29241, n29242, n29243,
    n29244, n29245, n29246, n29247, n29248, n29249,
    n29250, n29251, n29252, n29253, n29254, n29255,
    n29256, n29257, n29258, n29259, n29260, n29261,
    n29262, n29263, n29264, n29265, n29266, n29267,
    n29268, n29269, n29270, n29271, n29272, n29273,
    n29274, n29275, n29276, n29277, n29278, n29279,
    n29280, n29281, n29282, n29283, n29284, n29285,
    n29286, n29287, n29288, n29289, n29290, n29291,
    n29292, n29293, n29294, n29295, n29296, n29297,
    n29298, n29299, n29300, n29301, n29302, n29303,
    n29304, n29305, n29306, n29307, n29308, n29309,
    n29310, n29311, n29312, n29313, n29314, n29315,
    n29316, n29317, n29318, n29319, n29320, n29321,
    n29322, n29323, n29324, n29325, n29326, n29327,
    n29328, n29329, n29330, n29331, n29332, n29333,
    n29334, n29335, n29336, n29337, n29338, n29339,
    n29340, n29341, n29342, n29343, n29344, n29345,
    n29346, n29347, n29348, n29349, n29350, n29351,
    n29352, n29353, n29354, n29355, n29356, n29357,
    n29358, n29359, n29360, n29361, n29362, n29363,
    n29364, n29365, n29367, n29368, n29369, n29370,
    n29371, n29372, n29373, n29374, n29375, n29376,
    n29377, n29378, n29379, n29380, n29381, n29382,
    n29383, n29384, n29385, n29386, n29387, n29388,
    n29389, n29390, n29391, n29392, n29393, n29394,
    n29395, n29396, n29397, n29398, n29399, n29400,
    n29401, n29402, n29403, n29404, n29405, n29406,
    n29407, n29408, n29409, n29410, n29411, n29412,
    n29413, n29414, n29415, n29416, n29417, n29418,
    n29419, n29420, n29421, n29422, n29423, n29424,
    n29425, n29426, n29427, n29428, n29429, n29430,
    n29431, n29432, n29433, n29434, n29435, n29436,
    n29437, n29438, n29439, n29440, n29441, n29442,
    n29443, n29444, n29445, n29446, n29447, n29448,
    n29449, n29450, n29451, n29452, n29453, n29454,
    n29455, n29456, n29457, n29458, n29459, n29460,
    n29461, n29462, n29463, n29464, n29465, n29466,
    n29467, n29468, n29469, n29470, n29471, n29472,
    n29473, n29474, n29475, n29476, n29477, n29478,
    n29479, n29480, n29481, n29482, n29483, n29484,
    n29485, n29487, n29488, n29489, n29490, n29491,
    n29492, n29493, n29494, n29495, n29496, n29497,
    n29498, n29499, n29500, n29501, n29502, n29503,
    n29504, n29505, n29506, n29507, n29508, n29509,
    n29510, n29511, n29512, n29513, n29514, n29515,
    n29516, n29517, n29518, n29519, n29520, n29521,
    n29522, n29523, n29524, n29525, n29526, n29527,
    n29528, n29529, n29530, n29531, n29532, n29533,
    n29534, n29535, n29536, n29537, n29538, n29539,
    n29540, n29541, n29542, n29543, n29544, n29545,
    n29546, n29547, n29548, n29549, n29550, n29551,
    n29552, n29553, n29554, n29555, n29556, n29557,
    n29558, n29559, n29560, n29561, n29562, n29563,
    n29564, n29565, n29566, n29567, n29568, n29569,
    n29570, n29571, n29572, n29573, n29574, n29575,
    n29576, n29577, n29578, n29579, n29580, n29581,
    n29582, n29583, n29584, n29585, n29586, n29587,
    n29588, n29589, n29590, n29591, n29592, n29593,
    n29594, n29595, n29596, n29597, n29599, n29600,
    n29601, n29602, n29603, n29604, n29605, n29606,
    n29607, n29608, n29609, n29610, n29611, n29612,
    n29613, n29614, n29615, n29616, n29617, n29618,
    n29619, n29620, n29621, n29622, n29623, n29624,
    n29625, n29626, n29627, n29628, n29629, n29630,
    n29631, n29632, n29633, n29634, n29635, n29636,
    n29637, n29638, n29639, n29640, n29641, n29642,
    n29643, n29644, n29645, n29646, n29647, n29648,
    n29649, n29650, n29651, n29652, n29653, n29654,
    n29655, n29656, n29657, n29658, n29659, n29660,
    n29661, n29662, n29663, n29664, n29665, n29666,
    n29667, n29668, n29669, n29670, n29671, n29672,
    n29673, n29674, n29675, n29676, n29677, n29678,
    n29679, n29680, n29681, n29682, n29683, n29684,
    n29685, n29686, n29687, n29688, n29689, n29690,
    n29691, n29692, n29693, n29694, n29695, n29696,
    n29697, n29698, n29699, n29700, n29701, n29702,
    n29703, n29704, n29706, n29707, n29708, n29709,
    n29710, n29711, n29712, n29713, n29714, n29715,
    n29716, n29717, n29718, n29719, n29720, n29721,
    n29722, n29723, n29724, n29725, n29726, n29727,
    n29728, n29729, n29730, n29731, n29732, n29733,
    n29734, n29735, n29736, n29737, n29738, n29739,
    n29740, n29741, n29742, n29743, n29744, n29745,
    n29746, n29747, n29748, n29749, n29750, n29751,
    n29752, n29753, n29754, n29755, n29756, n29757,
    n29758, n29759, n29760, n29761, n29762, n29763,
    n29764, n29765, n29766, n29767, n29768, n29769,
    n29770, n29771, n29772, n29773, n29774, n29775,
    n29776, n29777, n29778, n29779, n29780, n29781,
    n29782, n29783, n29784, n29785, n29786, n29787,
    n29788, n29789, n29790, n29791, n29792, n29793,
    n29794, n29795, n29796, n29797, n29798, n29799,
    n29800, n29801, n29802, n29803, n29804, n29805,
    n29806, n29807, n29808, n29809, n29811, n29812,
    n29813, n29814, n29815, n29816, n29817, n29818,
    n29819, n29820, n29821, n29822, n29823, n29824,
    n29825, n29826, n29827, n29828, n29829, n29830,
    n29831, n29832, n29833, n29834, n29835, n29836,
    n29837, n29838, n29839, n29840, n29841, n29842,
    n29843, n29844, n29845, n29846, n29847, n29848,
    n29849, n29850, n29851, n29852, n29853, n29854,
    n29855, n29856, n29857, n29858, n29859, n29860,
    n29861, n29862, n29863, n29864, n29865, n29866,
    n29867, n29868, n29869, n29870, n29871, n29872,
    n29873, n29874, n29875, n29876, n29877, n29878,
    n29879, n29880, n29881, n29882, n29883, n29884,
    n29885, n29886, n29887, n29888, n29889, n29890,
    n29891, n29892, n29893, n29894, n29895, n29896,
    n29897, n29898, n29899, n29900, n29901, n29902,
    n29903, n29905, n29906, n29907, n29908, n29909,
    n29910, n29911, n29912, n29913, n29914, n29915,
    n29916, n29917, n29918, n29919, n29920, n29921,
    n29922, n29923, n29924, n29925, n29926, n29927,
    n29928, n29929, n29930, n29931, n29932, n29933,
    n29934, n29935, n29936, n29937, n29938, n29939,
    n29940, n29941, n29942, n29943, n29944, n29945,
    n29946, n29947, n29948, n29949, n29950, n29951,
    n29952, n29953, n29954, n29955, n29956, n29957,
    n29958, n29959, n29960, n29961, n29962, n29963,
    n29964, n29965, n29966, n29967, n29968, n29969,
    n29970, n29971, n29972, n29973, n29974, n29975,
    n29976, n29977, n29978, n29979, n29980, n29981,
    n29982, n29983, n29984, n29985, n29986, n29987,
    n29988, n29989, n29990, n29991, n29992, n29993,
    n29994, n29995, n29997, n29998, n29999, n30000,
    n30001, n30002, n30003, n30004, n30005, n30006,
    n30007, n30008, n30009, n30010, n30011, n30012,
    n30013, n30014, n30015, n30016, n30017, n30018,
    n30019, n30020, n30021, n30022, n30023, n30024,
    n30025, n30026, n30027, n30028, n30029, n30030,
    n30031, n30032, n30033, n30034, n30035, n30036,
    n30037, n30038, n30039, n30040, n30041, n30042,
    n30043, n30044, n30045, n30046, n30047, n30048,
    n30049, n30050, n30051, n30052, n30053, n30054,
    n30055, n30056, n30057, n30058, n30059, n30060,
    n30061, n30062, n30063, n30064, n30065, n30066,
    n30067, n30068, n30069, n30070, n30071, n30072,
    n30073, n30074, n30075, n30076, n30077, n30078,
    n30079, n30081, n30082, n30083, n30084, n30085,
    n30086, n30087, n30088, n30089, n30090, n30091,
    n30092, n30093, n30094, n30095, n30096, n30097,
    n30098, n30099, n30100, n30101, n30102, n30103,
    n30104, n30105, n30106, n30107, n30108, n30109,
    n30110, n30111, n30112, n30113, n30114, n30115,
    n30116, n30117, n30118, n30119, n30120, n30121,
    n30122, n30123, n30124, n30125, n30126, n30127,
    n30128, n30129, n30130, n30131, n30132, n30133,
    n30134, n30135, n30136, n30137, n30138, n30139,
    n30140, n30141, n30142, n30143, n30144, n30145,
    n30146, n30147, n30148, n30149, n30150, n30151,
    n30152, n30153, n30154, n30155, n30156, n30158,
    n30159, n30160, n30161, n30162, n30163, n30164,
    n30165, n30166, n30167, n30168, n30169, n30170,
    n30171, n30172, n30173, n30174, n30175, n30176,
    n30177, n30178, n30179, n30180, n30181, n30182,
    n30183, n30184, n30185, n30186, n30187, n30188,
    n30189, n30190, n30191, n30192, n30193, n30194,
    n30195, n30196, n30197, n30198, n30199, n30200,
    n30201, n30202, n30203, n30204, n30205, n30206,
    n30207, n30208, n30209, n30210, n30211, n30212,
    n30213, n30214, n30215, n30216, n30217, n30218,
    n30219, n30220, n30222, n30223, n30224, n30225,
    n30226, n30227, n30228, n30229, n30230, n30231,
    n30232, n30233, n30234, n30235, n30236, n30237,
    n30238, n30239, n30240, n30241, n30242, n30243,
    n30244, n30245, n30246, n30247, n30248, n30249,
    n30250, n30251, n30252, n30253, n30254, n30255,
    n30256, n30257, n30258, n30259, n30260, n30261,
    n30262, n30263, n30264, n30265, n30266, n30267,
    n30268, n30269, n30270, n30271, n30272, n30273,
    n30274, n30275;
  assign n65 = ~pi3  & pi4 ;
  assign n66 = pi3  & ~pi4 ;
  assign n67 = ~n65 & ~n66;
  assign n68 = pi2  & ~pi3 ;
  assign n69 = ~pi2  & pi3 ;
  assign n70 = ~n68 & ~n69;
  assign n71 = pi4  & ~pi5 ;
  assign n72 = ~pi4  & pi5 ;
  assign n73 = ~n71 & ~n72;
  assign n74 = n70 & ~n73;
  assign n75 = n67 & n74;
  assign n76 = pi25  & ~pi26 ;
  assign n77 = ~pi25  & pi26 ;
  assign n78 = ~n76 & ~n77;
  assign n79 = pi23  & ~pi24 ;
  assign n80 = ~pi23  & pi24 ;
  assign n81 = ~n79 & ~n80;
  assign n82 = pi24  & pi25 ;
  assign n83 = ~pi24  & ~pi25 ;
  assign n84 = ~n82 & ~n83;
  assign n85 = n81 & ~n84;
  assign n86 = ~n78 & n85;
  assign n87 = ~pi27  & pi28 ;
  assign n88 = pi29  & pi30 ;
  assign n89 = n87 & n88;
  assign n90 = ~pi24  & pi25 ;
  assign n91 = ~pi23  & ~pi26 ;
  assign n92 = n90 & n91;
  assign n93 = n89 & n92;
  assign n94 = ~pi29  & ~pi30 ;
  assign n95 = n87 & n94;
  assign n96 = pi23  & pi26 ;
  assign n97 = n83 & n96;
  assign n98 = n95 & n97;
  assign n99 = ~n93 & ~n98;
  assign n100 = pi29  & ~pi30 ;
  assign n101 = pi27  & ~pi28 ;
  assign n102 = n100 & n101;
  assign n103 = ~pi23  & pi26 ;
  assign n104 = pi24  & ~pi25 ;
  assign n105 = n103 & n104;
  assign n106 = n102 & n105;
  assign n107 = pi27  & pi28 ;
  assign n108 = ~pi29  & pi30 ;
  assign n109 = n107 & n108;
  assign n110 = n83 & n91;
  assign n111 = n109 & n110;
  assign n112 = ~pi27  & ~pi28 ;
  assign n113 = n100 & n112;
  assign n114 = pi23  & ~pi26 ;
  assign n115 = n104 & n114;
  assign n116 = n113 & n115;
  assign n117 = ~n111 & ~n116;
  assign n118 = ~n106 & n117;
  assign n119 = n82 & n103;
  assign n120 = n89 & n119;
  assign n121 = n96 & n104;
  assign n122 = n88 & n101;
  assign n123 = n121 & n122;
  assign n124 = ~n120 & ~n123;
  assign n125 = n82 & n91;
  assign n126 = n113 & n125;
  assign n127 = n90 & n103;
  assign n128 = n94 & n101;
  assign n129 = n127 & n128;
  assign n130 = n92 & n95;
  assign n131 = ~n126 & ~n129;
  assign n132 = ~n130 & n131;
  assign n133 = n124 & n132;
  assign n134 = n100 & n107;
  assign n135 = n127 & n134;
  assign n136 = n119 & n134;
  assign n137 = ~n135 & ~n136;
  assign n138 = n82 & n96;
  assign n139 = n134 & n138;
  assign n140 = n88 & n112;
  assign n141 = n138 & n140;
  assign n142 = ~n139 & ~n141;
  assign n143 = n105 & n140;
  assign n144 = n94 & n112;
  assign n145 = n125 & n144;
  assign n146 = ~n143 & ~n145;
  assign n147 = n87 & n100;
  assign n148 = n119 & n147;
  assign n149 = n110 & n128;
  assign n150 = ~n148 & ~n149;
  assign n151 = n122 & n125;
  assign n152 = n83 & n103;
  assign n153 = n140 & n152;
  assign n154 = ~n151 & ~n153;
  assign n155 = n115 & n128;
  assign n156 = n125 & n134;
  assign n157 = n87 & n108;
  assign n158 = n90 & n114;
  assign n159 = n157 & n158;
  assign n160 = ~n156 & ~n159;
  assign n161 = n82 & n114;
  assign n162 = n113 & n161;
  assign n163 = n113 & n138;
  assign n164 = ~n162 & ~n163;
  assign n165 = ~n155 & n160;
  assign n166 = n164 & n165;
  assign n167 = n128 & n161;
  assign n168 = n138 & n147;
  assign n169 = n83 & n114;
  assign n170 = n157 & n169;
  assign n171 = n102 & n127;
  assign n172 = ~n170 & ~n171;
  assign n173 = n91 & n104;
  assign n174 = n102 & n173;
  assign n175 = n147 & n173;
  assign n176 = ~n174 & ~n175;
  assign n177 = n144 & n152;
  assign n178 = n89 & n158;
  assign n179 = ~n177 & ~n178;
  assign n180 = n121 & n134;
  assign n181 = n90 & n96;
  assign n182 = n94 & n107;
  assign n183 = n181 & n182;
  assign n184 = n97 & n113;
  assign n185 = n88 & n107;
  assign n186 = n97 & n185;
  assign n187 = ~n184 & ~n186;
  assign n188 = n121 & n185;
  assign n189 = n95 & n121;
  assign n190 = n95 & n152;
  assign n191 = ~n188 & ~n189;
  assign n192 = ~n190 & n191;
  assign n193 = n119 & n122;
  assign n194 = n109 & n173;
  assign n195 = n113 & n127;
  assign n196 = n134 & n152;
  assign n197 = n92 & n109;
  assign n198 = ~n196 & ~n197;
  assign n199 = n125 & n147;
  assign n200 = n138 & n144;
  assign n201 = ~n199 & ~n200;
  assign n202 = ~n180 & ~n183;
  assign n203 = ~n193 & ~n194;
  assign n204 = ~n195 & n203;
  assign n205 = n179 & n202;
  assign n206 = n187 & n198;
  assign n207 = n201 & n206;
  assign n208 = n204 & n205;
  assign n209 = n192 & n208;
  assign n210 = n207 & n209;
  assign n211 = n110 & n147;
  assign n212 = n134 & n173;
  assign n213 = n138 & n185;
  assign n214 = n108 & n112;
  assign n215 = n125 & n214;
  assign n216 = n122 & n152;
  assign n217 = ~n215 & ~n216;
  assign n218 = ~n212 & ~n213;
  assign n219 = n217 & n218;
  assign n220 = ~n167 & ~n168;
  assign n221 = ~n211 & n220;
  assign n222 = n99 & n137;
  assign n223 = n142 & n146;
  assign n224 = n150 & n154;
  assign n225 = n172 & n176;
  assign n226 = n224 & n225;
  assign n227 = n222 & n223;
  assign n228 = n118 & n221;
  assign n229 = n219 & n228;
  assign n230 = n226 & n227;
  assign n231 = n133 & n166;
  assign n232 = n230 & n231;
  assign n233 = n229 & n232;
  assign n234 = n210 & n233;
  assign n235 = n97 & n134;
  assign n236 = n109 & n121;
  assign n237 = n102 & n121;
  assign n238 = n121 & n214;
  assign n239 = n95 & n119;
  assign n240 = ~n238 & ~n239;
  assign n241 = ~n237 & n240;
  assign n242 = n147 & n169;
  assign n243 = n125 & n128;
  assign n244 = ~n242 & ~n243;
  assign n245 = n109 & n181;
  assign n246 = n119 & n128;
  assign n247 = n140 & n173;
  assign n248 = n125 & n182;
  assign n249 = n97 & n128;
  assign n250 = n89 & n169;
  assign n251 = ~n249 & ~n250;
  assign n252 = n110 & n122;
  assign n253 = n92 & n128;
  assign n254 = ~n252 & ~n253;
  assign n255 = n161 & n182;
  assign n256 = n89 & n152;
  assign n257 = ~n255 & ~n256;
  assign n258 = n152 & n185;
  assign n259 = n121 & n182;
  assign n260 = ~n258 & ~n259;
  assign n261 = ~n245 & ~n246;
  assign n262 = ~n247 & ~n248;
  assign n263 = n261 & n262;
  assign n264 = n244 & n251;
  assign n265 = n254 & n257;
  assign n266 = n260 & n265;
  assign n267 = n263 & n264;
  assign n268 = n266 & n267;
  assign n269 = n147 & n161;
  assign n270 = n113 & n152;
  assign n271 = n92 & n113;
  assign n272 = ~n270 & ~n271;
  assign n273 = n169 & n185;
  assign n274 = n92 & n185;
  assign n275 = ~n273 & ~n274;
  assign n276 = n115 & n140;
  assign n277 = n121 & n157;
  assign n278 = n173 & n185;
  assign n279 = ~n277 & ~n278;
  assign n280 = n101 & n108;
  assign n281 = n97 & n280;
  assign n282 = n95 & n110;
  assign n283 = n134 & n158;
  assign n284 = n97 & n102;
  assign n285 = ~n282 & ~n283;
  assign n286 = ~n284 & n285;
  assign n287 = ~n276 & ~n281;
  assign n288 = n279 & n287;
  assign n289 = n286 & n288;
  assign n290 = n113 & n158;
  assign n291 = n144 & n161;
  assign n292 = ~n290 & ~n291;
  assign n293 = n97 & n157;
  assign n294 = n92 & n214;
  assign n295 = ~n293 & ~n294;
  assign n296 = n119 & n214;
  assign n297 = n157 & n181;
  assign n298 = ~n296 & ~n297;
  assign n299 = n102 & n110;
  assign n300 = n122 & n158;
  assign n301 = ~n299 & ~n300;
  assign n302 = n161 & n214;
  assign n303 = n89 & n121;
  assign n304 = n110 & n280;
  assign n305 = ~n302 & ~n303;
  assign n306 = ~n304 & n305;
  assign n307 = n109 & n125;
  assign n308 = n144 & n158;
  assign n309 = n121 & n280;
  assign n310 = n158 & n185;
  assign n311 = ~n309 & ~n310;
  assign n312 = n138 & n157;
  assign n313 = n113 & n121;
  assign n314 = n105 & n128;
  assign n315 = ~n312 & ~n313;
  assign n316 = ~n314 & n315;
  assign n317 = n113 & n119;
  assign n318 = n140 & n181;
  assign n319 = n105 & n113;
  assign n320 = ~n307 & ~n308;
  assign n321 = ~n317 & ~n318;
  assign n322 = ~n319 & n321;
  assign n323 = n311 & n320;
  assign n324 = n322 & n323;
  assign n325 = n306 & n316;
  assign n326 = n324 & n325;
  assign n327 = n169 & n214;
  assign n328 = n89 & n161;
  assign n329 = n95 & n125;
  assign n330 = n110 & n140;
  assign n331 = ~n329 & ~n330;
  assign n332 = n181 & n280;
  assign n333 = n138 & n280;
  assign n334 = n173 & n280;
  assign n335 = ~n332 & ~n333;
  assign n336 = ~n334 & n335;
  assign n337 = n121 & n147;
  assign n338 = n173 & n182;
  assign n339 = n122 & n173;
  assign n340 = ~n327 & ~n328;
  assign n341 = ~n337 & ~n338;
  assign n342 = ~n339 & n341;
  assign n343 = n292 & n340;
  assign n344 = n295 & n298;
  assign n345 = n301 & n331;
  assign n346 = n344 & n345;
  assign n347 = n342 & n343;
  assign n348 = n336 & n347;
  assign n349 = n289 & n346;
  assign n350 = n348 & n349;
  assign n351 = n326 & n350;
  assign n352 = n115 & n280;
  assign n353 = n157 & n161;
  assign n354 = ~n352 & ~n353;
  assign n355 = n95 & n173;
  assign n356 = n102 & n169;
  assign n357 = ~n355 & ~n356;
  assign n358 = n115 & n122;
  assign n359 = n158 & n280;
  assign n360 = ~n358 & ~n359;
  assign n361 = n119 & n144;
  assign n362 = n127 & n182;
  assign n363 = ~n361 & ~n362;
  assign n364 = n105 & n147;
  assign n365 = n127 & n185;
  assign n366 = ~n364 & ~n365;
  assign n367 = n113 & n181;
  assign n368 = n140 & n158;
  assign n369 = ~n367 & ~n368;
  assign n370 = n97 & n109;
  assign n371 = n95 & n138;
  assign n372 = ~n370 & ~n371;
  assign n373 = n127 & n214;
  assign n374 = n97 & n214;
  assign n375 = ~n373 & ~n374;
  assign n376 = n89 & n105;
  assign n377 = n95 & n127;
  assign n378 = n102 & n115;
  assign n379 = n140 & n161;
  assign n380 = n147 & n158;
  assign n381 = n109 & n119;
  assign n382 = n161 & n280;
  assign n383 = n115 & n157;
  assign n384 = ~n382 & ~n383;
  assign n385 = ~n376 & ~n377;
  assign n386 = ~n378 & ~n379;
  assign n387 = ~n380 & ~n381;
  assign n388 = n386 & n387;
  assign n389 = n384 & n385;
  assign n390 = n388 & n389;
  assign n391 = ~n235 & ~n236;
  assign n392 = ~n269 & n391;
  assign n393 = n272 & n275;
  assign n394 = n354 & n357;
  assign n395 = n360 & n363;
  assign n396 = n366 & n369;
  assign n397 = n372 & n375;
  assign n398 = n396 & n397;
  assign n399 = n394 & n395;
  assign n400 = n392 & n393;
  assign n401 = n241 & n400;
  assign n402 = n398 & n399;
  assign n403 = n390 & n402;
  assign n404 = n268 & n401;
  assign n405 = n403 & n404;
  assign n406 = n351 & n405;
  assign n407 = n234 & n406;
  assign n408 = n109 & n169;
  assign n409 = n121 & n140;
  assign n410 = ~n408 & ~n409;
  assign n411 = n110 & n134;
  assign n412 = n115 & n144;
  assign n413 = ~n411 & ~n412;
  assign n414 = n144 & n181;
  assign n415 = n125 & n157;
  assign n416 = n102 & n152;
  assign n417 = ~n415 & ~n416;
  assign n418 = ~n414 & n417;
  assign n419 = ~n249 & ~n378;
  assign n420 = n418 & n419;
  assign n421 = ~n129 & ~n329;
  assign n422 = n92 & n102;
  assign n423 = ~n304 & ~n422;
  assign n424 = ~n216 & ~n377;
  assign n425 = n295 & ~n368;
  assign n426 = n424 & n425;
  assign n427 = n109 & n161;
  assign n428 = ~n175 & ~n427;
  assign n429 = ~n252 & n428;
  assign n430 = n110 & n185;
  assign n431 = ~n167 & ~n430;
  assign n432 = n97 & n144;
  assign n433 = ~n199 & ~n432;
  assign n434 = ~n196 & ~n328;
  assign n435 = n109 & n152;
  assign n436 = ~n370 & ~n435;
  assign n437 = n115 & n214;
  assign n438 = n89 & n115;
  assign n439 = n134 & n161;
  assign n440 = ~n213 & ~n281;
  assign n441 = ~n374 & ~n439;
  assign n442 = n440 & n441;
  assign n443 = n89 & n125;
  assign n444 = ~n178 & ~n443;
  assign n445 = n102 & n181;
  assign n446 = n169 & n280;
  assign n447 = ~n334 & ~n446;
  assign n448 = ~n270 & ~n337;
  assign n449 = ~n141 & ~n149;
  assign n450 = ~n273 & ~n437;
  assign n451 = ~n438 & ~n445;
  assign n452 = n450 & n451;
  assign n453 = n444 & n449;
  assign n454 = n447 & n448;
  assign n455 = n453 & n454;
  assign n456 = n442 & n452;
  assign n457 = n455 & n456;
  assign n458 = n125 & n280;
  assign n459 = n140 & n169;
  assign n460 = n128 & n173;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n248 & ~n458;
  assign n463 = n410 & n462;
  assign n464 = n413 & n421;
  assign n465 = n423 & n431;
  assign n466 = n433 & n434;
  assign n467 = n436 & n461;
  assign n468 = n466 & n467;
  assign n469 = n464 & n465;
  assign n470 = n429 & n463;
  assign n471 = n469 & n470;
  assign n472 = n420 & n468;
  assign n473 = n426 & n472;
  assign n474 = n457 & n471;
  assign n475 = n473 & n474;
  assign n476 = n138 & n182;
  assign n477 = n134 & n181;
  assign n478 = ~n476 & ~n477;
  assign n479 = ~n247 & ~n312;
  assign n480 = n89 & n173;
  assign n481 = n158 & n182;
  assign n482 = n134 & n169;
  assign n483 = ~n276 & ~n482;
  assign n484 = ~n308 & ~n481;
  assign n485 = n483 & n484;
  assign n486 = n97 & n182;
  assign n487 = ~n246 & ~n486;
  assign n488 = n122 & n161;
  assign n489 = ~n98 & ~n361;
  assign n490 = ~n488 & n489;
  assign n491 = n487 & n490;
  assign n492 = ~n212 & ~n271;
  assign n493 = ~n338 & ~n480;
  assign n494 = n492 & n493;
  assign n495 = n478 & n479;
  assign n496 = n494 & n495;
  assign n497 = n485 & n496;
  assign n498 = n491 & n497;
  assign n499 = n127 & n140;
  assign n500 = ~n236 & ~n499;
  assign n501 = ~n284 & ~n291;
  assign n502 = n152 & n280;
  assign n503 = n121 & n144;
  assign n504 = ~n502 & ~n503;
  assign n505 = ~n163 & ~n274;
  assign n506 = ~n130 & ~n353;
  assign n507 = n505 & n506;
  assign n508 = n152 & n182;
  assign n509 = n89 & n138;
  assign n510 = n152 & n157;
  assign n511 = n119 & n280;
  assign n512 = n110 & n157;
  assign n513 = ~n382 & ~n512;
  assign n514 = ~n256 & ~n318;
  assign n515 = n173 & n214;
  assign n516 = ~n123 & ~n313;
  assign n517 = ~n515 & n516;
  assign n518 = n152 & n214;
  assign n519 = ~n93 & ~n518;
  assign n520 = n181 & n185;
  assign n521 = ~n310 & ~n520;
  assign n522 = n119 & n157;
  assign n523 = n121 & n128;
  assign n524 = ~n522 & ~n523;
  assign n525 = n127 & n147;
  assign n526 = n115 & n185;
  assign n527 = ~n525 & ~n526;
  assign n528 = ~n183 & ~n299;
  assign n529 = n105 & n122;
  assign n530 = ~n333 & ~n529;
  assign n531 = n105 & n214;
  assign n532 = n144 & n169;
  assign n533 = ~n531 & ~n532;
  assign n534 = n95 & n115;
  assign n535 = n92 & n140;
  assign n536 = n119 & n140;
  assign n537 = n97 & n122;
  assign n538 = ~n242 & ~n537;
  assign n539 = n119 & n185;
  assign n540 = ~n278 & ~n539;
  assign n541 = ~n194 & ~n534;
  assign n542 = ~n535 & ~n536;
  assign n543 = n541 & n542;
  assign n544 = n172 & n538;
  assign n545 = n540 & n544;
  assign n546 = n543 & n545;
  assign n547 = ~n162 & ~n253;
  assign n548 = ~n510 & ~n511;
  assign n549 = n547 & n548;
  assign n550 = n513 & n514;
  assign n551 = n519 & n521;
  assign n552 = n524 & n527;
  assign n553 = n528 & n530;
  assign n554 = n533 & n553;
  assign n555 = n551 & n552;
  assign n556 = n549 & n550;
  assign n557 = n517 & n556;
  assign n558 = n554 & n555;
  assign n559 = n557 & n558;
  assign n560 = n546 & n559;
  assign n561 = n95 & n169;
  assign n562 = ~n371 & ~n561;
  assign n563 = n110 & n113;
  assign n564 = n105 & n109;
  assign n565 = ~n563 & ~n564;
  assign n566 = n138 & n214;
  assign n567 = ~n269 & ~n566;
  assign n568 = n102 & n161;
  assign n569 = ~n156 & ~n195;
  assign n570 = ~n568 & n569;
  assign n571 = n137 & n570;
  assign n572 = ~n238 & ~n362;
  assign n573 = ~n508 & ~n509;
  assign n574 = n572 & n573;
  assign n575 = n117 & n500;
  assign n576 = n501 & n504;
  assign n577 = n562 & n565;
  assign n578 = n567 & n577;
  assign n579 = n575 & n576;
  assign n580 = n507 & n574;
  assign n581 = n579 & n580;
  assign n582 = n571 & n578;
  assign n583 = n581 & n582;
  assign n584 = n498 & n583;
  assign n585 = n475 & n584;
  assign n586 = n560 & n585;
  assign n587 = ~n407 & ~n586;
  assign n588 = n407 & n586;
  assign n589 = ~pi26  & ~n587;
  assign n590 = ~n588 & n589;
  assign n591 = ~n587 & ~n590;
  assign n592 = n128 & n169;
  assign n593 = ~n310 & ~n592;
  assign n594 = n105 & n157;
  assign n595 = ~n312 & ~n594;
  assign n596 = n109 & n127;
  assign n597 = n89 & n181;
  assign n598 = ~n278 & ~n597;
  assign n599 = n102 & n158;
  assign n600 = ~n568 & ~n599;
  assign n601 = n110 & n214;
  assign n602 = ~n211 & ~n601;
  assign n603 = n97 & n147;
  assign n604 = n92 & n122;
  assign n605 = n105 & n280;
  assign n606 = ~n377 & ~n459;
  assign n607 = ~n486 & ~n605;
  assign n608 = n606 & n607;
  assign n609 = ~n126 & ~n361;
  assign n610 = ~n526 & n609;
  assign n611 = ~n167 & ~n255;
  assign n612 = ~n290 & ~n308;
  assign n613 = ~n373 & ~n596;
  assign n614 = ~n603 & ~n604;
  assign n615 = n613 & n614;
  assign n616 = n611 & n612;
  assign n617 = n593 & n595;
  assign n618 = n598 & n600;
  assign n619 = n602 & n618;
  assign n620 = n616 & n617;
  assign n621 = n608 & n615;
  assign n622 = n610 & n621;
  assign n623 = n619 & n620;
  assign n624 = n622 & n623;
  assign n625 = n109 & n138;
  assign n626 = ~n332 & ~n625;
  assign n627 = n89 & n97;
  assign n628 = ~n120 & ~n627;
  assign n629 = ~n303 & ~n364;
  assign n630 = ~n414 & n629;
  assign n631 = ~n337 & ~n439;
  assign n632 = ~n522 & n631;
  assign n633 = ~n216 & ~n314;
  assign n634 = n128 & n158;
  assign n635 = ~n317 & ~n634;
  assign n636 = n102 & n119;
  assign n637 = ~n432 & ~n636;
  assign n638 = n102 & n138;
  assign n639 = n127 & n144;
  assign n640 = ~n638 & ~n639;
  assign n641 = ~n297 & ~n339;
  assign n642 = n637 & n641;
  assign n643 = n640 & n642;
  assign n644 = ~n408 & ~n509;
  assign n645 = ~n123 & ~n151;
  assign n646 = n147 & n152;
  assign n647 = ~n525 & ~n646;
  assign n648 = n127 & n280;
  assign n649 = ~n111 & ~n488;
  assign n650 = ~n648 & n649;
  assign n651 = n645 & n647;
  assign n652 = n650 & n651;
  assign n653 = n169 & n182;
  assign n654 = ~n512 & ~n653;
  assign n655 = ~n194 & ~n330;
  assign n656 = n127 & n157;
  assign n657 = ~n381 & ~n535;
  assign n658 = ~n368 & n657;
  assign n659 = ~n656 & n658;
  assign n660 = ~n338 & ~n376;
  assign n661 = n110 & n182;
  assign n662 = ~n276 & ~n661;
  assign n663 = n95 & n158;
  assign n664 = ~n170 & ~n663;
  assign n665 = n530 & ~n566;
  assign n666 = n654 & n655;
  assign n667 = n660 & n662;
  assign n668 = n664 & n667;
  assign n669 = n665 & n666;
  assign n670 = n668 & n669;
  assign n671 = n659 & n670;
  assign n672 = ~n277 & ~n416;
  assign n673 = ~n511 & n672;
  assign n674 = n301 & n626;
  assign n675 = n628 & n633;
  assign n676 = n635 & n644;
  assign n677 = n675 & n676;
  assign n678 = n673 & n674;
  assign n679 = n630 & n632;
  assign n680 = n678 & n679;
  assign n681 = n643 & n677;
  assign n682 = n652 & n681;
  assign n683 = n680 & n682;
  assign n684 = n671 & n683;
  assign n685 = n110 & n144;
  assign n686 = ~n446 & ~n685;
  assign n687 = n128 & n138;
  assign n688 = ~n274 & ~n687;
  assign n689 = n122 & n169;
  assign n690 = ~n156 & ~n270;
  assign n691 = ~n189 & ~n689;
  assign n692 = n690 & n691;
  assign n693 = ~n175 & ~n532;
  assign n694 = n538 & n693;
  assign n695 = n686 & n688;
  assign n696 = n694 & n695;
  assign n697 = n692 & n696;
  assign n698 = n115 & n134;
  assign n699 = ~n561 & ~n698;
  assign n700 = n102 & n125;
  assign n701 = ~n334 & ~n700;
  assign n702 = ~n367 & ~n563;
  assign n703 = n89 & n127;
  assign n704 = ~n327 & ~n703;
  assign n705 = ~n245 & ~n523;
  assign n706 = ~n247 & ~n304;
  assign n707 = ~n358 & ~n430;
  assign n708 = ~n515 & n707;
  assign n709 = n699 & n706;
  assign n710 = n701 & n702;
  assign n711 = n704 & n705;
  assign n712 = n710 & n711;
  assign n713 = n708 & n709;
  assign n714 = n712 & n713;
  assign n715 = n119 & n182;
  assign n716 = ~n508 & ~n715;
  assign n717 = ~n177 & n716;
  assign n718 = n92 & n134;
  assign n719 = ~n196 & ~n718;
  assign n720 = ~n309 & n719;
  assign n721 = n181 & n214;
  assign n722 = ~n139 & ~n721;
  assign n723 = n95 & n105;
  assign n724 = n92 & n144;
  assign n725 = ~n294 & ~n437;
  assign n726 = ~n243 & ~n273;
  assign n727 = ~n296 & ~n460;
  assign n728 = ~n476 & ~n723;
  assign n729 = ~n724 & n728;
  assign n730 = n726 & n727;
  assign n731 = n164 & n421;
  assign n732 = n722 & n725;
  assign n733 = n731 & n732;
  assign n734 = n729 & n730;
  assign n735 = n286 & n717;
  assign n736 = n720 & n735;
  assign n737 = n733 & n734;
  assign n738 = n736 & n737;
  assign n739 = n697 & n714;
  assign n740 = n738 & n739;
  assign n741 = n624 & n740;
  assign n742 = n684 & n741;
  assign n743 = ~n591 & n742;
  assign n744 = n591 & ~n742;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~n100 & ~n108;
  assign n747 = pi30  & pi31 ;
  assign n748 = n746 & n747;
  assign n749 = ~n149 & ~n367;
  assign n750 = ~n592 & ~n724;
  assign n751 = n144 & n173;
  assign n752 = ~n412 & ~n751;
  assign n753 = n115 & n182;
  assign n754 = n92 & n182;
  assign n755 = ~n753 & ~n754;
  assign n756 = ~n200 & ~n255;
  assign n757 = ~n338 & n756;
  assign n758 = ~n246 & ~n317;
  assign n759 = ~n282 & ~n687;
  assign n760 = ~n174 & ~n299;
  assign n761 = ~n378 & ~n422;
  assign n762 = ~n561 & n761;
  assign n763 = n357 & n760;
  assign n764 = n758 & n759;
  assign n765 = n763 & n764;
  assign n766 = n762 & n765;
  assign n767 = ~n248 & ~n358;
  assign n768 = n92 & n147;
  assign n769 = ~n327 & ~n768;
  assign n770 = n115 & n147;
  assign n771 = ~n199 & ~n380;
  assign n772 = ~n481 & ~n646;
  assign n773 = ~n770 & n772;
  assign n774 = n767 & n771;
  assign n775 = n769 & n774;
  assign n776 = n773 & n775;
  assign n777 = ~n190 & ~n276;
  assign n778 = ~n339 & ~n368;
  assign n779 = n137 & n778;
  assign n780 = n777 & n779;
  assign n781 = n720 & n780;
  assign n782 = ~n236 & ~n459;
  assign n783 = ~n511 & n782;
  assign n784 = ~n235 & ~n636;
  assign n785 = ~n98 & ~n186;
  assign n786 = ~n283 & ~n439;
  assign n787 = n125 & n140;
  assign n788 = ~n180 & ~n536;
  assign n789 = ~n252 & ~n359;
  assign n790 = ~n381 & ~n432;
  assign n791 = ~n143 & ~n520;
  assign n792 = n92 & n280;
  assign n793 = ~n332 & ~n352;
  assign n794 = ~n792 & n793;
  assign n795 = n790 & n791;
  assign n796 = n794 & n795;
  assign n797 = ~n189 & ~n723;
  assign n798 = n113 & n169;
  assign n799 = ~n715 & ~n798;
  assign n800 = ~n596 & ~n625;
  assign n801 = ~n177 & ~n330;
  assign n802 = ~n141 & ~n512;
  assign n803 = ~n601 & ~n638;
  assign n804 = n800 & n803;
  assign n805 = n801 & n802;
  assign n806 = n804 & n805;
  assign n807 = ~n167 & ~n188;
  assign n808 = n157 & n173;
  assign n809 = ~n477 & ~n808;
  assign n810 = n128 & n152;
  assign n811 = ~n213 & ~n535;
  assign n812 = ~n810 & n811;
  assign n813 = ~n139 & ~n605;
  assign n814 = n105 & n134;
  assign n815 = ~n409 & ~n814;
  assign n816 = ~n116 & ~n247;
  assign n817 = ~n379 & n816;
  assign n818 = n813 & n815;
  assign n819 = n817 & n818;
  assign n820 = n812 & n819;
  assign n821 = ~n648 & n807;
  assign n822 = n809 & n821;
  assign n823 = n820 & n822;
  assign n824 = ~n153 & ~n249;
  assign n825 = ~n281 & ~n382;
  assign n826 = ~n787 & n825;
  assign n827 = n784 & n824;
  assign n828 = n785 & n786;
  assign n829 = n788 & n789;
  assign n830 = n797 & n799;
  assign n831 = n829 & n830;
  assign n832 = n827 & n828;
  assign n833 = n826 & n832;
  assign n834 = n796 & n831;
  assign n835 = n806 & n834;
  assign n836 = n833 & n835;
  assign n837 = n823 & n836;
  assign n838 = n105 & n144;
  assign n839 = n105 & n185;
  assign n840 = ~n365 & ~n839;
  assign n841 = n113 & n173;
  assign n842 = ~n242 & ~n838;
  assign n843 = ~n841 & n842;
  assign n844 = n840 & n843;
  assign n845 = ~n245 & ~n476;
  assign n846 = n97 & n140;
  assign n847 = ~n689 & ~n846;
  assign n848 = ~n243 & ~n502;
  assign n849 = ~n175 & n845;
  assign n850 = n847 & n848;
  assign n851 = n849 & n850;
  assign n852 = ~n458 & ~n539;
  assign n853 = ~n211 & ~n499;
  assign n854 = n852 & n853;
  assign n855 = ~n156 & ~n170;
  assign n856 = ~n271 & ~n318;
  assign n857 = ~n333 & ~n377;
  assign n858 = ~n563 & n857;
  assign n859 = n855 & n856;
  assign n860 = n858 & n859;
  assign n861 = n783 & n854;
  assign n862 = n860 & n861;
  assign n863 = n844 & n851;
  assign n864 = n862 & n863;
  assign n865 = n781 & n864;
  assign n866 = n837 & n865;
  assign n867 = ~n163 & ~n269;
  assign n868 = ~n564 & ~n604;
  assign n869 = n867 & n868;
  assign n870 = n447 & n749;
  assign n871 = n750 & n752;
  assign n872 = n755 & n871;
  assign n873 = n869 & n870;
  assign n874 = n757 & n873;
  assign n875 = n872 & n874;
  assign n876 = n766 & n776;
  assign n877 = n875 & n876;
  assign n878 = n866 & n877;
  assign n879 = n748 & ~n878;
  assign n880 = pi31  & ~n746;
  assign n881 = ~n333 & ~n648;
  assign n882 = ~n502 & n881;
  assign n883 = ~n359 & ~n458;
  assign n884 = ~n170 & ~n281;
  assign n885 = ~n309 & ~n511;
  assign n886 = ~n605 & n885;
  assign n887 = n513 & n884;
  assign n888 = n883 & n887;
  assign n889 = n794 & n886;
  assign n890 = n882 & n889;
  assign n891 = n888 & n890;
  assign n892 = ~n361 & ~n532;
  assign n893 = n128 & n181;
  assign n894 = n109 & n115;
  assign n895 = ~n482 & ~n698;
  assign n896 = ~n212 & n895;
  assign n897 = ~n685 & n896;
  assign n898 = ~n211 & ~n242;
  assign n899 = ~n638 & n898;
  assign n900 = ~n129 & ~n523;
  assign n901 = ~n168 & ~n838;
  assign n902 = n109 & n158;
  assign n903 = ~n307 & n436;
  assign n904 = ~n902 & n903;
  assign n905 = ~n503 & ~n639;
  assign n906 = ~n411 & ~n414;
  assign n907 = ~n432 & ~n476;
  assign n908 = ~n563 & n907;
  assign n909 = n901 & n906;
  assign n910 = n905 & n909;
  assign n911 = n908 & n910;
  assign n912 = n904 & n911;
  assign n913 = ~n270 & ~n377;
  assign n914 = ~n167 & ~n190;
  assign n915 = ~n353 & n914;
  assign n916 = n913 & n915;
  assign n917 = ~n162 & ~n290;
  assign n918 = ~n126 & ~n314;
  assign n919 = ~n383 & ~n653;
  assign n920 = n918 & n919;
  assign n921 = n917 & n920;
  assign n922 = n95 & n181;
  assign n923 = ~n380 & ~n603;
  assign n924 = n785 & n923;
  assign n925 = ~n277 & ~n415;
  assign n926 = ~n159 & ~n297;
  assign n927 = ~n408 & ~n510;
  assign n928 = ~n522 & n927;
  assign n929 = n925 & n926;
  assign n930 = n928 & n929;
  assign n931 = n595 & ~n656;
  assign n932 = n930 & n931;
  assign n933 = ~n188 & ~n213;
  assign n934 = n840 & n933;
  assign n935 = ~n271 & ~n337;
  assign n936 = ~n243 & ~n371;
  assign n937 = n92 & n157;
  assign n938 = ~n810 & ~n937;
  assign n939 = ~n646 & ~n661;
  assign n940 = ~n239 & ~n808;
  assign n941 = ~n195 & ~n319;
  assign n942 = ~n269 & ~n313;
  assign n943 = n941 & n942;
  assign n944 = n147 & n181;
  assign n945 = ~n111 & ~n184;
  assign n946 = ~n194 & ~n199;
  assign n947 = ~n539 & ~n723;
  assign n948 = ~n770 & ~n944;
  assign n949 = n947 & n948;
  assign n950 = n945 & n946;
  assign n951 = n935 & n936;
  assign n952 = n938 & n939;
  assign n953 = n940 & n952;
  assign n954 = n950 & n951;
  assign n955 = n943 & n949;
  assign n956 = n954 & n955;
  assign n957 = n953 & n956;
  assign n958 = ~n148 & ~n768;
  assign n959 = ~n189 & ~n525;
  assign n960 = ~n293 & ~n364;
  assign n961 = ~n116 & ~n249;
  assign n962 = ~n520 & ~n841;
  assign n963 = ~n922 & n962;
  assign n964 = n958 & n961;
  assign n965 = n959 & n960;
  assign n966 = n964 & n965;
  assign n967 = n924 & n963;
  assign n968 = n934 & n967;
  assign n969 = n916 & n966;
  assign n970 = n921 & n969;
  assign n971 = n932 & n968;
  assign n972 = n970 & n971;
  assign n973 = n957 & n972;
  assign n974 = ~n177 & ~n197;
  assign n975 = ~n636 & ~n893;
  assign n976 = ~n894 & n975;
  assign n977 = n428 & n974;
  assign n978 = n447 & n799;
  assign n979 = n892 & n900;
  assign n980 = n978 & n979;
  assign n981 = n976 & n977;
  assign n982 = n899 & n981;
  assign n983 = n897 & n980;
  assign n984 = n982 & n983;
  assign n985 = n891 & n984;
  assign n986 = n912 & n985;
  assign n987 = n973 & n986;
  assign n988 = ~n878 & ~n987;
  assign n989 = n122 & n138;
  assign n990 = ~n250 & ~n412;
  assign n991 = ~n989 & n990;
  assign n992 = ~n383 & ~n937;
  assign n993 = ~n159 & ~n178;
  assign n994 = ~n242 & n993;
  assign n995 = ~n93 & ~n239;
  assign n996 = ~n432 & ~n508;
  assign n997 = n995 & n996;
  assign n998 = n366 & n992;
  assign n999 = n997 & n998;
  assign n1000 = n991 & n994;
  assign n1001 = n999 & n1000;
  assign n1002 = n89 & n110;
  assign n1003 = ~n638 & ~n1002;
  assign n1004 = ~n314 & ~n438;
  assign n1005 = ~n523 & ~n639;
  assign n1006 = ~n126 & ~n520;
  assign n1007 = ~n283 & ~n563;
  assign n1008 = n600 & n1007;
  assign n1009 = ~n300 & ~n537;
  assign n1010 = ~n330 & ~n839;
  assign n1011 = ~n382 & ~n754;
  assign n1012 = ~n196 & ~n518;
  assign n1013 = n658 & n800;
  assign n1014 = ~n167 & ~n294;
  assign n1015 = ~n502 & n749;
  assign n1016 = n1014 & n1015;
  assign n1017 = ~n437 & ~n439;
  assign n1018 = ~n700 & ~n753;
  assign n1019 = ~n193 & ~n415;
  assign n1020 = ~n123 & ~n156;
  assign n1021 = ~n177 & n1020;
  assign n1022 = ~n246 & ~n281;
  assign n1023 = n1018 & n1022;
  assign n1024 = n1019 & n1023;
  assign n1025 = n1021 & n1024;
  assign n1026 = ~n236 & ~n247;
  assign n1027 = ~n510 & n1026;
  assign n1028 = n845 & n1027;
  assign n1029 = ~n594 & ~n603;
  assign n1030 = ~n685 & n1029;
  assign n1031 = ~n151 & ~n293;
  assign n1032 = n122 & n181;
  assign n1033 = ~n270 & ~n1032;
  assign n1034 = n158 & n214;
  assign n1035 = ~n488 & ~n1034;
  assign n1036 = ~n284 & ~n718;
  assign n1037 = n777 & n1036;
  assign n1038 = n1017 & n1031;
  assign n1039 = n1033 & n1035;
  assign n1040 = n1038 & n1039;
  assign n1041 = n1030 & n1037;
  assign n1042 = n1040 & n1041;
  assign n1043 = n1016 & n1028;
  assign n1044 = n1042 & n1043;
  assign n1045 = n1025 & n1044;
  assign n1046 = n354 & n785;
  assign n1047 = ~n338 & ~n515;
  assign n1048 = ~n243 & n1047;
  assign n1049 = ~n302 & ~n792;
  assign n1050 = ~n277 & n1049;
  assign n1051 = n122 & n127;
  assign n1052 = ~n145 & ~n459;
  assign n1053 = ~n297 & ~n308;
  assign n1054 = ~n200 & ~n416;
  assign n1055 = ~n656 & ~n1051;
  assign n1056 = n1054 & n1055;
  assign n1057 = n883 & n1052;
  assign n1058 = n1053 & n1057;
  assign n1059 = n1056 & n1058;
  assign n1060 = n217 & ~n529;
  assign n1061 = n759 & n799;
  assign n1062 = n1009 & n1010;
  assign n1063 = n1011 & n1012;
  assign n1064 = n1062 & n1063;
  assign n1065 = n1060 & n1061;
  assign n1066 = n1008 & n1046;
  assign n1067 = n1048 & n1050;
  assign n1068 = n1066 & n1067;
  assign n1069 = n1064 & n1065;
  assign n1070 = n1013 & n1069;
  assign n1071 = n1059 & n1068;
  assign n1072 = n1070 & n1071;
  assign n1073 = n1045 & n1072;
  assign n1074 = ~n486 & ~n944;
  assign n1075 = ~n290 & ~n337;
  assign n1076 = ~n534 & ~n814;
  assign n1077 = ~n922 & n1076;
  assign n1078 = n164 & n1075;
  assign n1079 = n1074 & n1078;
  assign n1080 = n1077 & n1079;
  assign n1081 = ~n130 & ~n480;
  assign n1082 = ~n751 & n784;
  assign n1083 = n1081 & n1082;
  assign n1084 = ~n155 & ~n460;
  assign n1085 = ~n503 & n1084;
  assign n1086 = n105 & n182;
  assign n1087 = ~n317 & ~n1086;
  assign n1088 = ~n175 & ~n564;
  assign n1089 = ~n211 & ~n299;
  assign n1090 = ~n525 & ~n539;
  assign n1091 = n1089 & n1090;
  assign n1092 = n447 & n933;
  assign n1093 = n1003 & n1004;
  assign n1094 = n1005 & n1006;
  assign n1095 = n1087 & n1088;
  assign n1096 = n1094 & n1095;
  assign n1097 = n1092 & n1093;
  assign n1098 = n1085 & n1091;
  assign n1099 = n1097 & n1098;
  assign n1100 = n1083 & n1096;
  assign n1101 = n1099 & n1100;
  assign n1102 = n1001 & n1080;
  assign n1103 = n1101 & n1102;
  assign n1104 = n1073 & n1103;
  assign n1105 = ~n878 & ~n1104;
  assign n1106 = ~n213 & ~n314;
  assign n1107 = ~n328 & ~n460;
  assign n1108 = ~n510 & ~n838;
  assign n1109 = n1107 & n1108;
  assign n1110 = n354 & n1106;
  assign n1111 = n1109 & n1110;
  assign n1112 = ~n126 & ~n522;
  assign n1113 = ~n290 & ~n408;
  assign n1114 = n117 & ~n184;
  assign n1115 = n478 & n1113;
  assign n1116 = n1114 & n1115;
  assign n1117 = ~n238 & ~n486;
  assign n1118 = ~n511 & ~n596;
  assign n1119 = n1117 & n1118;
  assign n1120 = ~n174 & ~n259;
  assign n1121 = ~n180 & n1120;
  assign n1122 = ~n529 & ~n1051;
  assign n1123 = ~n365 & ~n415;
  assign n1124 = ~n312 & ~n409;
  assign n1125 = ~n488 & ~n846;
  assign n1126 = n1124 & n1125;
  assign n1127 = n1122 & n1123;
  assign n1128 = n1126 & n1127;
  assign n1129 = n1121 & n1128;
  assign n1130 = ~n374 & ~n605;
  assign n1131 = ~n216 & ~n599;
  assign n1132 = n1130 & n1131;
  assign n1133 = ~n319 & ~n663;
  assign n1134 = ~n481 & ~n839;
  assign n1135 = n1133 & n1134;
  assign n1136 = ~n200 & ~n253;
  assign n1137 = ~n135 & n1136;
  assign n1138 = ~n194 & ~n332;
  assign n1139 = ~n383 & n1138;
  assign n1140 = n1137 & n1139;
  assign n1141 = ~n446 & ~n723;
  assign n1142 = ~n597 & ~n661;
  assign n1143 = ~n787 & n1142;
  assign n1144 = ~n129 & ~n309;
  assign n1145 = ~n362 & ~n371;
  assign n1146 = n387 & ~n715;
  assign n1147 = n1144 & n1145;
  assign n1148 = n1141 & n1147;
  assign n1149 = n1143 & n1146;
  assign n1150 = n1148 & n1149;
  assign n1151 = ~n237 & ~n700;
  assign n1152 = ~n303 & n1151;
  assign n1153 = ~n123 & ~n143;
  assign n1154 = ~n153 & ~n294;
  assign n1155 = ~n334 & ~n338;
  assign n1156 = ~n503 & ~n508;
  assign n1157 = ~n648 & n1156;
  assign n1158 = n1154 & n1155;
  assign n1159 = n500 & n1153;
  assign n1160 = n1158 & n1159;
  assign n1161 = n1135 & n1157;
  assign n1162 = n1152 & n1161;
  assign n1163 = n1140 & n1160;
  assign n1164 = n1162 & n1163;
  assign n1165 = n1150 & n1164;
  assign n1166 = ~n120 & ~n186;
  assign n1167 = ~n520 & ~n539;
  assign n1168 = ~n703 & n1167;
  assign n1169 = n1166 & n1168;
  assign n1170 = ~n156 & n786;
  assign n1171 = ~n168 & ~n356;
  assign n1172 = ~n106 & n958;
  assign n1173 = n1171 & n1172;
  assign n1174 = ~n636 & ~n718;
  assign n1175 = ~n770 & ~n894;
  assign n1176 = ~n308 & ~n922;
  assign n1177 = ~n177 & ~n246;
  assign n1178 = ~n561 & ~n564;
  assign n1179 = n1177 & n1178;
  assign n1180 = n1174 & n1175;
  assign n1181 = n1176 & n1180;
  assign n1182 = n1170 & n1179;
  assign n1183 = n1181 & n1182;
  assign n1184 = n1169 & n1173;
  assign n1185 = n1183 & n1184;
  assign n1186 = ~n364 & ~n531;
  assign n1187 = ~n300 & ~n337;
  assign n1188 = ~n243 & ~n751;
  assign n1189 = ~n151 & ~n534;
  assign n1190 = ~n625 & n1189;
  assign n1191 = n1188 & n1190;
  assign n1192 = ~n190 & ~n414;
  assign n1193 = ~n515 & ~n603;
  assign n1194 = ~n841 & n1193;
  assign n1195 = n1192 & n1194;
  assign n1196 = ~n159 & ~n188;
  assign n1197 = ~n367 & n1196;
  assign n1198 = ~n245 & ~n379;
  assign n1199 = ~n373 & ~n443;
  assign n1200 = ~n638 & n1199;
  assign n1201 = n514 & n938;
  assign n1202 = n1186 & n1187;
  assign n1203 = n1198 & n1202;
  assign n1204 = n1200 & n1201;
  assign n1205 = n1197 & n1204;
  assign n1206 = n1191 & n1203;
  assign n1207 = n1195 & n1206;
  assign n1208 = n1205 & n1207;
  assign n1209 = ~n211 & ~n317;
  assign n1210 = ~n376 & ~n411;
  assign n1211 = ~n437 & ~n537;
  assign n1212 = ~n627 & ~n753;
  assign n1213 = ~n792 & n1212;
  assign n1214 = n1210 & n1211;
  assign n1215 = n1112 & n1209;
  assign n1216 = n1214 & n1215;
  assign n1217 = n1119 & n1213;
  assign n1218 = n1132 & n1217;
  assign n1219 = n1111 & n1216;
  assign n1220 = n1116 & n1219;
  assign n1221 = n1129 & n1218;
  assign n1222 = n1220 & n1221;
  assign n1223 = n1185 & n1222;
  assign n1224 = n1165 & n1208;
  assign n1225 = n1223 & n1224;
  assign n1226 = ~n1104 & ~n1225;
  assign n1227 = ~n159 & ~n768;
  assign n1228 = n479 & n1227;
  assign n1229 = ~n309 & ~n414;
  assign n1230 = ~n283 & ~n512;
  assign n1231 = ~n168 & ~n376;
  assign n1232 = ~n634 & ~n638;
  assign n1233 = ~n893 & n1232;
  assign n1234 = n1229 & n1231;
  assign n1235 = n1230 & n1234;
  assign n1236 = n1233 & n1235;
  assign n1237 = ~n515 & ~n627;
  assign n1238 = ~n687 & ~n724;
  assign n1239 = n1237 & n1238;
  assign n1240 = ~n236 & ~n246;
  assign n1241 = ~n596 & n1240;
  assign n1242 = ~n334 & ~n509;
  assign n1243 = ~n460 & ~n841;
  assign n1244 = ~n259 & ~n503;
  assign n1245 = ~n522 & ~n787;
  assign n1246 = ~n171 & ~n278;
  assign n1247 = ~n199 & ~n846;
  assign n1248 = ~n256 & ~n526;
  assign n1249 = ~n365 & ~n715;
  assign n1250 = ~n902 & n1249;
  assign n1251 = n788 & n900;
  assign n1252 = n1242 & n1243;
  assign n1253 = n1244 & n1245;
  assign n1254 = n1246 & n1247;
  assign n1255 = n1248 & n1254;
  assign n1256 = n1252 & n1253;
  assign n1257 = n1250 & n1251;
  assign n1258 = n1228 & n1239;
  assign n1259 = n1241 & n1258;
  assign n1260 = n1256 & n1257;
  assign n1261 = n1255 & n1260;
  assign n1262 = n1236 & n1259;
  assign n1263 = n1261 & n1262;
  assign n1264 = ~n330 & ~n508;
  assign n1265 = ~n636 & n1264;
  assign n1266 = ~n136 & ~n481;
  assign n1267 = n431 & n1266;
  assign n1268 = ~n141 & ~n313;
  assign n1269 = n722 & n1268;
  assign n1270 = ~n188 & ~n378;
  assign n1271 = ~n592 & ~n603;
  assign n1272 = ~n383 & ~n520;
  assign n1273 = ~n177 & ~n242;
  assign n1274 = ~n416 & ~n458;
  assign n1275 = ~n810 & n1274;
  assign n1276 = n702 & n1273;
  assign n1277 = n1275 & n1276;
  assign n1278 = ~n314 & ~n338;
  assign n1279 = ~n382 & n1278;
  assign n1280 = n251 & n719;
  assign n1281 = ~n273 & ~n605;
  assign n1282 = ~n989 & n1281;
  assign n1283 = ~n197 & ~n300;
  assign n1284 = ~n106 & ~n374;
  assign n1285 = ~n531 & ~n539;
  assign n1286 = ~n839 & n1285;
  assign n1287 = n164 & n789;
  assign n1288 = n1283 & n1284;
  assign n1289 = n1287 & n1288;
  assign n1290 = n1286 & n1289;
  assign n1291 = ~n155 & ~n371;
  assign n1292 = ~n293 & ~n568;
  assign n1293 = ~n663 & ~n1002;
  assign n1294 = ~n333 & ~n1032;
  assign n1295 = ~n239 & ~n248;
  assign n1296 = ~n130 & ~n329;
  assign n1297 = ~n183 & ~n356;
  assign n1298 = ~n459 & ~n599;
  assign n1299 = ~n770 & n1298;
  assign n1300 = n187 & n1297;
  assign n1301 = n1294 & n1295;
  assign n1302 = n1296 & n1301;
  assign n1303 = n1299 & n1300;
  assign n1304 = n1302 & n1303;
  assign n1305 = ~n189 & ~n328;
  assign n1306 = ~n212 & ~n594;
  assign n1307 = ~n153 & ~n525;
  assign n1308 = ~n291 & ~n482;
  assign n1309 = ~n296 & ~n379;
  assign n1310 = n1035 & n1309;
  assign n1311 = n1188 & n1291;
  assign n1312 = n1292 & n1293;
  assign n1313 = n1305 & n1306;
  assign n1314 = n1307 & n1308;
  assign n1315 = n1313 & n1314;
  assign n1316 = n1311 & n1312;
  assign n1317 = n1310 & n1316;
  assign n1318 = n1315 & n1317;
  assign n1319 = n1290 & n1304;
  assign n1320 = n1318 & n1319;
  assign n1321 = ~n290 & ~n937;
  assign n1322 = ~n111 & ~n308;
  assign n1323 = ~n639 & n1322;
  assign n1324 = n1141 & n1321;
  assign n1325 = n1323 & n1324;
  assign n1326 = n1280 & n1282;
  assign n1327 = n1325 & n1326;
  assign n1328 = n1320 & n1327;
  assign n1329 = ~n151 & ~n193;
  assign n1330 = ~n532 & ~n564;
  assign n1331 = n1329 & n1330;
  assign n1332 = ~n148 & ~n253;
  assign n1333 = ~n443 & n1332;
  assign n1334 = n217 & n1270;
  assign n1335 = n1271 & n1272;
  assign n1336 = n1334 & n1335;
  assign n1337 = n1265 & n1333;
  assign n1338 = n1267 & n1269;
  assign n1339 = n1279 & n1331;
  assign n1340 = n1338 & n1339;
  assign n1341 = n1336 & n1337;
  assign n1342 = n1277 & n1341;
  assign n1343 = n1340 & n1342;
  assign n1344 = n1263 & n1343;
  assign n1345 = n1328 & n1344;
  assign n1346 = ~n1225 & ~n1345;
  assign n1347 = ~n238 & ~n566;
  assign n1348 = ~n302 & ~n515;
  assign n1349 = n1347 & n1348;
  assign n1350 = ~n151 & ~n522;
  assign n1351 = ~n339 & ~n536;
  assign n1352 = ~n235 & ~n427;
  assign n1353 = ~n476 & n1352;
  assign n1354 = ~n430 & ~n715;
  assign n1355 = ~n171 & ~n409;
  assign n1356 = ~n293 & ~n721;
  assign n1357 = ~n364 & ~n770;
  assign n1358 = ~n564 & ~n893;
  assign n1359 = ~n438 & ~n937;
  assign n1360 = n433 & n1358;
  assign n1361 = n1359 & n1360;
  assign n1362 = ~n126 & ~n162;
  assign n1363 = ~n482 & ~n599;
  assign n1364 = n1362 & n1363;
  assign n1365 = n530 & n593;
  assign n1366 = n1291 & n1350;
  assign n1367 = n1351 & n1354;
  assign n1368 = n1355 & n1356;
  assign n1369 = n1357 & n1368;
  assign n1370 = n1366 & n1367;
  assign n1371 = n1364 & n1365;
  assign n1372 = n1349 & n1353;
  assign n1373 = n1371 & n1372;
  assign n1374 = n1369 & n1370;
  assign n1375 = n1361 & n1374;
  assign n1376 = n1373 & n1375;
  assign n1377 = ~n148 & ~n700;
  assign n1378 = ~n480 & ~n636;
  assign n1379 = n1198 & n1378;
  assign n1380 = ~n330 & ~n787;
  assign n1381 = ~n352 & ~n408;
  assign n1382 = n1380 & n1381;
  assign n1383 = ~n143 & ~n291;
  assign n1384 = ~n534 & ~n568;
  assign n1385 = ~n460 & n1383;
  assign n1386 = n1384 & n1385;
  assign n1387 = ~n273 & ~n1032;
  assign n1388 = ~n170 & ~n653;
  assign n1389 = ~n269 & ~n271;
  assign n1390 = ~n255 & ~n329;
  assign n1391 = ~n698 & ~n839;
  assign n1392 = ~n509 & ~n922;
  assign n1393 = n1391 & n1392;
  assign n1394 = ~n98 & ~n411;
  assign n1395 = ~n535 & ~n601;
  assign n1396 = ~n605 & ~n656;
  assign n1397 = ~n718 & ~n944;
  assign n1398 = n1396 & n1397;
  assign n1399 = n1394 & n1395;
  assign n1400 = n504 & n1399;
  assign n1401 = n1393 & n1398;
  assign n1402 = n1400 & n1401;
  assign n1403 = ~n378 & ~n437;
  assign n1404 = n125 & n185;
  assign n1405 = ~n383 & ~n703;
  assign n1406 = ~n1404 & n1405;
  assign n1407 = ~n188 & ~n259;
  assign n1408 = ~n359 & ~n374;
  assign n1409 = ~n415 & ~n1086;
  assign n1410 = n1408 & n1409;
  assign n1411 = n1387 & n1407;
  assign n1412 = n1388 & n1389;
  assign n1413 = n1390 & n1403;
  assign n1414 = n1412 & n1413;
  assign n1415 = n1410 & n1411;
  assign n1416 = n1406 & n1415;
  assign n1417 = n1386 & n1414;
  assign n1418 = n1416 & n1417;
  assign n1419 = n1402 & n1418;
  assign n1420 = ~n248 & ~n307;
  assign n1421 = ~n186 & ~n213;
  assign n1422 = ~n174 & ~n290;
  assign n1423 = ~n276 & ~n443;
  assign n1424 = ~n361 & ~n724;
  assign n1425 = ~n246 & n1422;
  assign n1426 = n1423 & n1424;
  assign n1427 = n1425 & n1426;
  assign n1428 = ~n193 & ~n303;
  assign n1429 = ~n180 & ~n754;
  assign n1430 = ~n445 & ~n648;
  assign n1431 = ~n422 & ~n1034;
  assign n1432 = n1429 & n1431;
  assign n1433 = n1430 & n1432;
  assign n1434 = ~n277 & ~n328;
  assign n1435 = ~n355 & n1434;
  assign n1436 = n137 & n1283;
  assign n1437 = n1377 & n1420;
  assign n1438 = n1421 & n1428;
  assign n1439 = n1437 & n1438;
  assign n1440 = n1435 & n1436;
  assign n1441 = n1379 & n1382;
  assign n1442 = n1440 & n1441;
  assign n1443 = n1427 & n1439;
  assign n1444 = n1433 & n1443;
  assign n1445 = n697 & n1442;
  assign n1446 = n1444 & n1445;
  assign n1447 = n1376 & n1446;
  assign n1448 = n1419 & n1447;
  assign n1449 = ~n1345 & ~n1448;
  assign n1450 = ~n482 & ~n989;
  assign n1451 = ~n458 & ~n721;
  assign n1452 = ~n278 & ~n435;
  assign n1453 = ~n536 & ~n1086;
  assign n1454 = ~n238 & ~n477;
  assign n1455 = ~n256 & n1454;
  assign n1456 = ~n445 & ~n798;
  assign n1457 = ~n106 & ~n522;
  assign n1458 = ~n136 & ~n141;
  assign n1459 = ~n296 & n1458;
  assign n1460 = n301 & n1005;
  assign n1461 = n1420 & n1450;
  assign n1462 = n1451 & n1452;
  assign n1463 = n1453 & n1456;
  assign n1464 = n1457 & n1463;
  assign n1465 = n1461 & n1462;
  assign n1466 = n1459 & n1460;
  assign n1467 = n1455 & n1466;
  assign n1468 = n1464 & n1465;
  assign n1469 = n1467 & n1468;
  assign n1470 = ~n274 & ~n1032;
  assign n1471 = ~n148 & ~n685;
  assign n1472 = ~n358 & ~n412;
  assign n1473 = ~n568 & n1472;
  assign n1474 = ~n359 & ~n443;
  assign n1475 = ~n603 & ~n687;
  assign n1476 = ~n93 & ~n770;
  assign n1477 = n1174 & n1476;
  assign n1478 = ~n271 & ~n509;
  assign n1479 = ~n213 & ~n304;
  assign n1480 = ~n518 & ~n902;
  assign n1481 = n1479 & n1480;
  assign n1482 = n1474 & n1475;
  assign n1483 = n1478 & n1482;
  assign n1484 = n1477 & n1481;
  assign n1485 = n1483 & n1484;
  assign n1486 = ~n283 & ~n312;
  assign n1487 = n161 & n185;
  assign n1488 = ~n190 & ~n1487;
  assign n1489 = ~n163 & ~n689;
  assign n1490 = ~n98 & ~n211;
  assign n1491 = ~n537 & n1490;
  assign n1492 = ~n525 & ~n634;
  assign n1493 = ~n189 & ~n235;
  assign n1494 = ~n276 & ~n356;
  assign n1495 = ~n563 & n1494;
  assign n1496 = n533 & n1493;
  assign n1497 = n567 & n593;
  assign n1498 = n1035 & n1049;
  assign n1499 = n1052 & n1123;
  assign n1500 = n1388 & n1489;
  assign n1501 = n1492 & n1500;
  assign n1502 = n1498 & n1499;
  assign n1503 = n1496 & n1497;
  assign n1504 = n1491 & n1495;
  assign n1505 = n1503 & n1504;
  assign n1506 = n1501 & n1502;
  assign n1507 = n1505 & n1506;
  assign n1508 = ~n195 & ~n313;
  assign n1509 = ~n534 & ~n561;
  assign n1510 = ~n277 & ~n437;
  assign n1511 = ~n330 & ~n808;
  assign n1512 = n1508 & n1511;
  assign n1513 = n1509 & n1510;
  assign n1514 = n1512 & n1513;
  assign n1515 = ~n196 & ~n430;
  assign n1516 = ~n215 & ~n480;
  assign n1517 = n187 & n375;
  assign n1518 = n1516 & n1517;
  assign n1519 = n292 & ~n317;
  assign n1520 = n354 & n369;
  assign n1521 = n1470 & n1471;
  assign n1522 = n1486 & n1488;
  assign n1523 = n1515 & n1522;
  assign n1524 = n1520 & n1521;
  assign n1525 = n1473 & n1519;
  assign n1526 = n1524 & n1525;
  assign n1527 = n1514 & n1523;
  assign n1528 = n1518 & n1527;
  assign n1529 = n1485 & n1526;
  assign n1530 = n1528 & n1529;
  assign n1531 = n1469 & n1507;
  assign n1532 = n1530 & n1531;
  assign n1533 = n1165 & n1532;
  assign n1534 = ~n1448 & ~n1533;
  assign n1535 = ~n177 & n752;
  assign n1536 = ~n145 & ~n184;
  assign n1537 = n1535 & n1536;
  assign n1538 = ~n197 & ~n437;
  assign n1539 = ~n281 & ~n989;
  assign n1540 = ~n339 & ~n352;
  assign n1541 = ~n537 & n1540;
  assign n1542 = ~n627 & ~n653;
  assign n1543 = ~n1051 & n1542;
  assign n1544 = n428 & n1543;
  assign n1545 = n924 & n1544;
  assign n1546 = ~n422 & ~n636;
  assign n1547 = n1357 & n1546;
  assign n1548 = ~n153 & ~n167;
  assign n1549 = ~n381 & ~n476;
  assign n1550 = ~n639 & n1549;
  assign n1551 = n434 & n1548;
  assign n1552 = n1171 & n1268;
  assign n1553 = n1423 & n1470;
  assign n1554 = n1538 & n1539;
  assign n1555 = n1553 & n1554;
  assign n1556 = n1551 & n1552;
  assign n1557 = n1541 & n1550;
  assign n1558 = n1547 & n1557;
  assign n1559 = n1555 & n1556;
  assign n1560 = n1537 & n1559;
  assign n1561 = n1545 & n1558;
  assign n1562 = n1560 & n1561;
  assign n1563 = ~n120 & ~n810;
  assign n1564 = ~n477 & ~n488;
  assign n1565 = ~n243 & ~n307;
  assign n1566 = ~n332 & n1565;
  assign n1567 = n421 & n1563;
  assign n1568 = n1564 & n1567;
  assign n1569 = n1566 & n1568;
  assign n1570 = ~n841 & ~n1002;
  assign n1571 = ~n460 & n1570;
  assign n1572 = ~n432 & n1571;
  assign n1573 = ~n159 & ~n922;
  assign n1574 = n600 & n1573;
  assign n1575 = ~n123 & ~n838;
  assign n1576 = ~n135 & ~n768;
  assign n1577 = n1575 & n1576;
  assign n1578 = ~n212 & ~n563;
  assign n1579 = ~n299 & ~n689;
  assign n1580 = ~n284 & ~n592;
  assign n1581 = ~n1034 & n1580;
  assign n1582 = n1424 & n1579;
  assign n1583 = n1581 & n1582;
  assign n1584 = ~n156 & ~n237;
  assign n1585 = ~n814 & n1584;
  assign n1586 = n1278 & n1585;
  assign n1587 = ~n249 & ~n358;
  assign n1588 = ~n383 & ~n594;
  assign n1589 = ~n605 & ~n754;
  assign n1590 = ~n792 & n1589;
  assign n1591 = n1587 & n1588;
  assign n1592 = n150 & n1247;
  assign n1593 = n1591 & n1592;
  assign n1594 = n1590 & n1593;
  assign n1595 = n1586 & n1594;
  assign n1596 = ~n258 & ~n458;
  assign n1597 = ~n718 & n1596;
  assign n1598 = n257 & n479;
  assign n1599 = n1133 & n1198;
  assign n1600 = n1578 & n1599;
  assign n1601 = n1597 & n1598;
  assign n1602 = n1331 & n1574;
  assign n1603 = n1577 & n1602;
  assign n1604 = n1600 & n1601;
  assign n1605 = n1583 & n1604;
  assign n1606 = n1603 & n1605;
  assign n1607 = n1595 & n1606;
  assign n1608 = ~n190 & ~n529;
  assign n1609 = ~n604 & n1608;
  assign n1610 = ~n163 & ~n216;
  assign n1611 = ~n271 & ~n297;
  assign n1612 = ~n353 & ~n459;
  assign n1613 = ~n526 & ~n787;
  assign n1614 = n1612 & n1613;
  assign n1615 = n1610 & n1611;
  assign n1616 = n644 & n789;
  assign n1617 = n1615 & n1616;
  assign n1618 = n1609 & n1614;
  assign n1619 = n1617 & n1618;
  assign n1620 = ~n139 & ~n246;
  assign n1621 = ~n646 & n1620;
  assign n1622 = ~n269 & ~n512;
  assign n1623 = ~n300 & ~n601;
  assign n1624 = n1622 & n1623;
  assign n1625 = ~n294 & ~n365;
  assign n1626 = ~n377 & ~n482;
  assign n1627 = n1625 & n1626;
  assign n1628 = n1006 & n1136;
  assign n1629 = n1295 & n1628;
  assign n1630 = n1621 & n1627;
  assign n1631 = n1624 & n1630;
  assign n1632 = n1572 & n1629;
  assign n1633 = n1631 & n1632;
  assign n1634 = n1569 & n1619;
  assign n1635 = n1633 & n1634;
  assign n1636 = n1562 & n1635;
  assign n1637 = n1607 & n1636;
  assign n1638 = ~n1533 & ~n1637;
  assign n1639 = ~n141 & ~n143;
  assign n1640 = ~n236 & ~n252;
  assign n1641 = n1429 & n1640;
  assign n1642 = ~n168 & ~n597;
  assign n1643 = ~n317 & ~n638;
  assign n1644 = ~n715 & ~n989;
  assign n1645 = ~n359 & ~n364;
  assign n1646 = ~n648 & n1645;
  assign n1647 = n725 & n1643;
  assign n1648 = n1644 & n1647;
  assign n1649 = n1646 & n1648;
  assign n1650 = ~n293 & ~n446;
  assign n1651 = ~n535 & ~n1002;
  assign n1652 = ~n274 & ~n307;
  assign n1653 = ~n408 & n704;
  assign n1654 = n807 & n848;
  assign n1655 = n1639 & n1642;
  assign n1656 = n1650 & n1651;
  assign n1657 = n1652 & n1656;
  assign n1658 = n1654 & n1655;
  assign n1659 = n1641 & n1653;
  assign n1660 = n1658 & n1659;
  assign n1661 = n1657 & n1660;
  assign n1662 = n1649 & n1661;
  assign n1663 = ~n409 & ~n481;
  assign n1664 = ~n277 & ~n367;
  assign n1665 = ~n377 & ~n787;
  assign n1666 = n1664 & n1665;
  assign n1667 = n1246 & n1663;
  assign n1668 = n1666 & n1667;
  assign n1669 = ~n194 & ~n753;
  assign n1670 = ~n139 & ~n193;
  assign n1671 = ~n379 & ~n723;
  assign n1672 = ~n338 & ~n460;
  assign n1673 = ~n361 & ~n378;
  assign n1674 = ~n605 & ~n689;
  assign n1675 = ~n178 & ~n215;
  assign n1676 = ~n594 & ~n698;
  assign n1677 = n1675 & n1676;
  assign n1678 = n1673 & n1674;
  assign n1679 = n1677 & n1678;
  assign n1680 = ~n162 & ~n175;
  assign n1681 = ~n302 & ~n314;
  assign n1682 = ~n625 & n1681;
  assign n1683 = n1680 & n1682;
  assign n1684 = ~n432 & ~n532;
  assign n1685 = ~n195 & ~n808;
  assign n1686 = ~n339 & ~n838;
  assign n1687 = ~n902 & n1686;
  assign n1688 = n1074 & n1578;
  assign n1689 = n1670 & n1671;
  assign n1690 = n1672 & n1684;
  assign n1691 = n1685 & n1690;
  assign n1692 = n1688 & n1689;
  assign n1693 = n1687 & n1692;
  assign n1694 = n1679 & n1691;
  assign n1695 = n1683 & n1694;
  assign n1696 = n1693 & n1695;
  assign n1697 = ~n458 & ~n508;
  assign n1698 = n137 & n1697;
  assign n1699 = n95 & n161;
  assign n1700 = ~n435 & n1488;
  assign n1701 = ~n177 & ~n245;
  assign n1702 = ~n922 & n1701;
  assign n1703 = ~n213 & ~n627;
  assign n1704 = ~n1699 & n1703;
  assign n1705 = n519 & n1151;
  assign n1706 = n1242 & n1272;
  assign n1707 = n1475 & n1669;
  assign n1708 = n1706 & n1707;
  assign n1709 = n1704 & n1705;
  assign n1710 = n1698 & n1700;
  assign n1711 = n1702 & n1710;
  assign n1712 = n1708 & n1709;
  assign n1713 = n1668 & n1712;
  assign n1714 = n1304 & n1711;
  assign n1715 = n1713 & n1714;
  assign n1716 = n1662 & n1715;
  assign n1717 = n1696 & n1716;
  assign n1718 = ~n1637 & ~n1717;
  assign n1719 = ~n190 & ~n243;
  assign n1720 = ~n634 & ~n838;
  assign n1721 = n1719 & n1720;
  assign n1722 = ~n330 & ~n1404;
  assign n1723 = n647 & n705;
  assign n1724 = n1722 & n1723;
  assign n1725 = ~n162 & ~n502;
  assign n1726 = ~n638 & n1725;
  assign n1727 = ~n327 & ~n381;
  assign n1728 = ~n944 & n1727;
  assign n1729 = ~n531 & ~n648;
  assign n1730 = ~n143 & ~n247;
  assign n1731 = ~n139 & ~n248;
  assign n1732 = ~n278 & ~n568;
  assign n1733 = n1731 & n1732;
  assign n1734 = n1004 & n1729;
  assign n1735 = n1730 & n1734;
  assign n1736 = n1726 & n1733;
  assign n1737 = n1728 & n1736;
  assign n1738 = n1735 & n1737;
  assign n1739 = ~n197 & ~n364;
  assign n1740 = ~n382 & ~n458;
  assign n1741 = ~n601 & ~n792;
  assign n1742 = n1740 & n1741;
  assign n1743 = n257 & n1739;
  assign n1744 = n440 & n628;
  assign n1745 = n1743 & n1744;
  assign n1746 = n1353 & n1742;
  assign n1747 = n1721 & n1746;
  assign n1748 = n1724 & n1745;
  assign n1749 = n1747 & n1748;
  assign n1750 = n1738 & n1749;
  assign n1751 = ~n304 & ~n566;
  assign n1752 = ~n184 & ~n604;
  assign n1753 = ~n186 & ~n563;
  assign n1754 = ~n194 & ~n1086;
  assign n1755 = ~n539 & ~n718;
  assign n1756 = ~n258 & ~n488;
  assign n1757 = ~n685 & n1756;
  assign n1758 = n595 & n1751;
  assign n1759 = n1752 & n1753;
  assign n1760 = n1754 & n1755;
  assign n1761 = n1759 & n1760;
  assign n1762 = n1757 & n1758;
  assign n1763 = n1761 & n1762;
  assign n1764 = ~n111 & ~n215;
  assign n1765 = ~n293 & n802;
  assign n1766 = n1764 & n1765;
  assign n1767 = ~n284 & ~n411;
  assign n1768 = ~n106 & ~n211;
  assign n1769 = ~n520 & n1768;
  assign n1770 = n1136 & n1769;
  assign n1771 = ~n123 & ~n592;
  assign n1772 = ~n159 & ~n499;
  assign n1773 = ~n1487 & n1772;
  assign n1774 = ~n239 & ~n374;
  assign n1775 = n154 & n1774;
  assign n1776 = n637 & n1771;
  assign n1777 = n1775 & n1776;
  assign n1778 = n1773 & n1777;
  assign n1779 = ~n508 & ~n1002;
  assign n1780 = ~n175 & ~n319;
  assign n1781 = ~n661 & n1780;
  assign n1782 = ~n377 & ~n724;
  assign n1783 = ~n283 & ~n290;
  assign n1784 = ~n307 & ~n537;
  assign n1785 = ~n989 & ~n1034;
  assign n1786 = n1784 & n1785;
  assign n1787 = n179 & n958;
  assign n1788 = n1782 & n1783;
  assign n1789 = n1787 & n1788;
  assign n1790 = n1781 & n1786;
  assign n1791 = n1789 & n1790;
  assign n1792 = ~n155 & ~n358;
  assign n1793 = ~n564 & n1792;
  assign n1794 = n1510 & n1793;
  assign n1795 = ~n171 & ~n249;
  assign n1796 = ~n291 & ~n937;
  assign n1797 = n1795 & n1796;
  assign n1798 = n840 & n1797;
  assign n1799 = ~n259 & ~n273;
  assign n1800 = ~n303 & ~n362;
  assign n1801 = ~n814 & n1800;
  assign n1802 = n301 & n1799;
  assign n1803 = n799 & n1779;
  assign n1804 = n1802 & n1803;
  assign n1805 = n1241 & n1801;
  assign n1806 = n1804 & n1805;
  assign n1807 = n1770 & n1794;
  assign n1808 = n1798 & n1807;
  assign n1809 = n1778 & n1806;
  assign n1810 = n1791 & n1809;
  assign n1811 = n1808 & n1810;
  assign n1812 = ~n599 & ~n625;
  assign n1813 = ~n380 & ~n639;
  assign n1814 = ~n317 & ~n329;
  assign n1815 = ~n212 & ~n216;
  assign n1816 = ~n269 & ~n787;
  assign n1817 = n1815 & n1816;
  assign n1818 = n1122 & n1229;
  assign n1819 = n1642 & n1812;
  assign n1820 = n1813 & n1814;
  assign n1821 = n1819 & n1820;
  assign n1822 = n1817 & n1818;
  assign n1823 = n1821 & n1822;
  assign n1824 = ~n332 & n369;
  assign n1825 = n1685 & n1824;
  assign n1826 = ~n188 & ~n459;
  assign n1827 = ~n126 & ~n135;
  assign n1828 = ~n334 & ~n416;
  assign n1829 = ~n503 & ~n515;
  assign n1830 = ~n810 & ~n922;
  assign n1831 = n1829 & n1830;
  assign n1832 = n1827 & n1828;
  assign n1833 = n1767 & n1826;
  assign n1834 = n1832 & n1833;
  assign n1835 = n1831 & n1834;
  assign n1836 = n1766 & n1825;
  assign n1837 = n1835 & n1836;
  assign n1838 = n1763 & n1823;
  assign n1839 = n1837 & n1838;
  assign n1840 = n1750 & n1839;
  assign n1841 = n1811 & n1840;
  assign n1842 = ~n1717 & ~n1841;
  assign n1843 = ~n359 & ~n411;
  assign n1844 = ~n307 & n1843;
  assign n1845 = ~n332 & ~n526;
  assign n1846 = ~n438 & ~n721;
  assign n1847 = ~n180 & ~n383;
  assign n1848 = ~n534 & ~n1699;
  assign n1849 = n1847 & n1848;
  assign n1850 = ~n193 & ~n304;
  assign n1851 = ~n508 & ~n798;
  assign n1852 = n1850 & n1851;
  assign n1853 = n1845 & n1846;
  assign n1854 = n1852 & n1853;
  assign n1855 = n1143 & n1844;
  assign n1856 = n1849 & n1855;
  assign n1857 = n1854 & n1856;
  assign n1858 = ~n248 & ~n296;
  assign n1859 = ~n199 & ~n282;
  assign n1860 = ~n503 & n1424;
  assign n1861 = n1859 & n1860;
  assign n1862 = n1455 & n1861;
  assign n1863 = ~n594 & ~n636;
  assign n1864 = ~n126 & ~n249;
  assign n1865 = ~n318 & ~n687;
  assign n1866 = ~n239 & ~n373;
  assign n1867 = n1794 & n1866;
  assign n1868 = ~n435 & ~n703;
  assign n1869 = ~n1404 & n1868;
  assign n1870 = n434 & n635;
  assign n1871 = n644 & n690;
  assign n1872 = n1508 & n1863;
  assign n1873 = n1864 & n1865;
  assign n1874 = n1872 & n1873;
  assign n1875 = n1870 & n1871;
  assign n1876 = n1535 & n1869;
  assign n1877 = n1571 & n1876;
  assign n1878 = n1874 & n1875;
  assign n1879 = n1766 & n1878;
  assign n1880 = n820 & n1877;
  assign n1881 = n1867 & n1880;
  assign n1882 = n1879 & n1881;
  assign n1883 = ~n415 & ~n1051;
  assign n1884 = ~n273 & ~n902;
  assign n1885 = ~n271 & ~n333;
  assign n1886 = ~n439 & ~n481;
  assign n1887 = n1885 & n1886;
  assign n1888 = n1883 & n1884;
  assign n1889 = n1887 & n1888;
  assign n1890 = ~n356 & ~n522;
  assign n1891 = ~n302 & ~n480;
  assign n1892 = ~n638 & n1891;
  assign n1893 = n749 & n1892;
  assign n1894 = ~n252 & ~n319;
  assign n1895 = ~n374 & ~n937;
  assign n1896 = ~n1487 & n1895;
  assign n1897 = n1307 & n1894;
  assign n1898 = n1858 & n1890;
  assign n1899 = n1897 & n1898;
  assign n1900 = n854 & n1896;
  assign n1901 = n1048 & n1577;
  assign n1902 = n1900 & n1901;
  assign n1903 = n1889 & n1899;
  assign n1904 = n1893 & n1903;
  assign n1905 = n1862 & n1902;
  assign n1906 = n1904 & n1905;
  assign n1907 = n1857 & n1906;
  assign n1908 = n1882 & n1907;
  assign n1909 = ~n1841 & ~n1908;
  assign n1910 = ~n247 & n1489;
  assign n1911 = ~n143 & ~n293;
  assign n1912 = ~n1404 & n1911;
  assign n1913 = ~n215 & ~n327;
  assign n1914 = ~n199 & ~n1699;
  assign n1915 = ~n253 & ~n661;
  assign n1916 = n99 & ~n186;
  assign n1917 = ~n303 & ~n568;
  assign n1918 = ~n592 & n1917;
  assign n1919 = ~n368 & ~n893;
  assign n1920 = n1915 & n1919;
  assign n1921 = n1916 & n1920;
  assign n1922 = n1918 & n1921;
  assign n1923 = ~n195 & ~n312;
  assign n1924 = ~n636 & ~n715;
  assign n1925 = ~n753 & ~n787;
  assign n1926 = ~n937 & n1925;
  assign n1927 = n1923 & n1924;
  assign n1928 = n301 & n933;
  assign n1929 = n1390 & n1457;
  assign n1930 = n1538 & n1913;
  assign n1931 = n1914 & n1930;
  assign n1932 = n1928 & n1929;
  assign n1933 = n1926 & n1927;
  assign n1934 = n1910 & n1912;
  assign n1935 = n1933 & n1934;
  assign n1936 = n1931 & n1932;
  assign n1937 = n1935 & n1936;
  assign n1938 = n1922 & n1937;
  assign n1939 = ~n170 & ~n270;
  assign n1940 = ~n126 & ~n362;
  assign n1941 = ~n414 & ~n422;
  assign n1942 = ~n459 & ~n1051;
  assign n1943 = n1941 & n1942;
  assign n1944 = n719 & n1940;
  assign n1945 = n1939 & n1944;
  assign n1946 = n1943 & n1945;
  assign n1947 = ~n377 & ~n814;
  assign n1948 = ~n353 & ~n458;
  assign n1949 = ~n274 & ~n318;
  assign n1950 = ~n480 & ~n1086;
  assign n1951 = n1949 & n1950;
  assign n1952 = n1053 & n1948;
  assign n1953 = n1951 & n1952;
  assign n1954 = ~n111 & ~n294;
  assign n1955 = ~n446 & n1954;
  assign n1956 = n602 & n1243;
  assign n1957 = n1955 & n1956;
  assign n1958 = ~n194 & ~n296;
  assign n1959 = ~n256 & ~n482;
  assign n1960 = ~n520 & n1959;
  assign n1961 = n1958 & n1960;
  assign n1962 = ~n252 & ~n944;
  assign n1963 = ~n242 & ~n282;
  assign n1964 = ~n534 & ~n594;
  assign n1965 = ~n638 & ~n646;
  assign n1966 = ~n846 & ~n894;
  assign n1967 = n1965 & n1966;
  assign n1968 = n1963 & n1964;
  assign n1969 = n1962 & n1968;
  assign n1970 = n1967 & n1969;
  assign n1971 = ~n189 & ~n236;
  assign n1972 = ~n258 & ~n503;
  assign n1973 = ~n605 & ~n798;
  assign n1974 = ~n808 & ~n838;
  assign n1975 = n1973 & n1974;
  assign n1976 = n840 & n1972;
  assign n1977 = n1420 & n1430;
  assign n1978 = n1971 & n1977;
  assign n1979 = n1975 & n1976;
  assign n1980 = n1279 & n1609;
  assign n1981 = n1979 & n1980;
  assign n1982 = n1961 & n1978;
  assign n1983 = n1981 & n1982;
  assign n1984 = n1970 & n1983;
  assign n1985 = ~n371 & n900;
  assign n1986 = ~n249 & ~n328;
  assign n1987 = ~n333 & ~n663;
  assign n1988 = n1986 & n1987;
  assign n1989 = n635 & n1642;
  assign n1990 = n1947 & n1989;
  assign n1991 = n1050 & n1988;
  assign n1992 = n1985 & n1991;
  assign n1993 = n1953 & n1990;
  assign n1994 = n1957 & n1993;
  assign n1995 = n1946 & n1992;
  assign n1996 = n1994 & n1995;
  assign n1997 = n1938 & n1996;
  assign n1998 = n1984 & n1997;
  assign n1999 = ~n1908 & ~n1998;
  assign n2000 = ~n328 & ~n334;
  assign n2001 = ~n601 & n2000;
  assign n2002 = ~n276 & ~n371;
  assign n2003 = n784 & n2002;
  assign n2004 = ~n162 & ~n170;
  assign n2005 = ~n330 & ~n520;
  assign n2006 = n2004 & n2005;
  assign n2007 = ~n481 & ~n689;
  assign n2008 = ~n646 & n2007;
  assign n2009 = ~n358 & ~n535;
  assign n2010 = n160 & n2009;
  assign n2011 = n448 & n1011;
  assign n2012 = n1685 & n2011;
  assign n2013 = n608 & n2010;
  assign n2014 = n2001 & n2003;
  assign n2015 = n2006 & n2008;
  assign n2016 = n2014 & n2015;
  assign n2017 = n2012 & n2013;
  assign n2018 = n2016 & n2017;
  assign n2019 = n1862 & n2018;
  assign n2020 = ~n446 & ~n596;
  assign n2021 = ~n416 & n2020;
  assign n2022 = ~n130 & ~n411;
  assign n2023 = n176 & n2022;
  assign n2024 = ~n255 & ~n511;
  assign n2025 = ~n111 & ~n277;
  assign n2026 = ~n297 & ~n313;
  assign n2027 = ~n376 & ~n526;
  assign n2028 = ~n564 & ~n846;
  assign n2029 = n2027 & n2028;
  assign n2030 = n2025 & n2026;
  assign n2031 = n2024 & n2030;
  assign n2032 = n2021 & n2029;
  assign n2033 = n2023 & n2032;
  assign n2034 = n2031 & n2033;
  assign n2035 = ~n163 & ~n291;
  assign n2036 = ~n537 & n2035;
  assign n2037 = ~n200 & ~n922;
  assign n2038 = ~n259 & ~n302;
  assign n2039 = n2037 & n2038;
  assign n2040 = ~n258 & ~n787;
  assign n2041 = ~n145 & ~n250;
  assign n2042 = ~n499 & ~n656;
  assign n2043 = ~n197 & ~n445;
  assign n2044 = ~n106 & ~n362;
  assign n2045 = ~n143 & ~n415;
  assign n2046 = ~n502 & ~n661;
  assign n2047 = ~n1032 & n2046;
  assign n2048 = n2042 & n2045;
  assign n2049 = n2043 & n2044;
  assign n2050 = n2048 & n2049;
  assign n2051 = n2047 & n2050;
  assign n2052 = ~n422 & ~n653;
  assign n2053 = ~n379 & ~n718;
  assign n2054 = ~n894 & n2053;
  assign n2055 = ~n129 & ~n252;
  assign n2056 = ~n408 & ~n439;
  assign n2057 = n2055 & n2056;
  assign n2058 = n2054 & n2057;
  assign n2059 = ~n284 & ~n332;
  assign n2060 = ~n751 & n1720;
  assign n2061 = n2059 & n2060;
  assign n2062 = ~n148 & ~n352;
  assign n2063 = ~n563 & ~n568;
  assign n2064 = ~n770 & ~n1699;
  assign n2065 = n2063 & n2064;
  assign n2066 = n1133 & n2062;
  assign n2067 = n1243 & n1451;
  assign n2068 = n2040 & n2041;
  assign n2069 = n2052 & n2068;
  assign n2070 = n2066 & n2067;
  assign n2071 = n2065 & n2070;
  assign n2072 = n2058 & n2069;
  assign n2073 = n2061 & n2072;
  assign n2074 = n2051 & n2071;
  assign n2075 = n2073 & n2074;
  assign n2076 = ~n189 & ~n523;
  assign n2077 = ~n536 & n2076;
  assign n2078 = ~n155 & ~n237;
  assign n2079 = ~n338 & ~n603;
  assign n2080 = ~n604 & n2079;
  assign n2081 = n2078 & n2080;
  assign n2082 = n2077 & n2081;
  assign n2083 = n699 & n1754;
  assign n2084 = n1913 & n2083;
  assign n2085 = ~n120 & ~n139;
  assign n2086 = n749 & n2085;
  assign n2087 = n898 & n1031;
  assign n2088 = n1684 & n1751;
  assign n2089 = n1864 & n2088;
  assign n2090 = n2086 & n2087;
  assign n2091 = n2036 & n2039;
  assign n2092 = n2090 & n2091;
  assign n2093 = n2084 & n2089;
  assign n2094 = n2092 & n2093;
  assign n2095 = n2082 & n2094;
  assign n2096 = n2034 & n2095;
  assign n2097 = n2019 & n2075;
  assign n2098 = n2096 & n2097;
  assign n2099 = ~n1998 & ~n2098;
  assign n2100 = ~n458 & ~n1699;
  assign n2101 = n688 & n2100;
  assign n2102 = n1640 & n2101;
  assign n2103 = ~n98 & ~n129;
  assign n2104 = ~n246 & ~n798;
  assign n2105 = n2103 & n2104;
  assign n2106 = ~n136 & ~n178;
  assign n2107 = ~n838 & n2106;
  assign n2108 = ~n379 & ~n846;
  assign n2109 = ~n383 & n749;
  assign n2110 = n1457 & n2109;
  assign n2111 = ~n177 & ~n296;
  assign n2112 = ~n318 & ~n373;
  assign n2113 = ~n661 & ~n698;
  assign n2114 = ~n715 & n2113;
  assign n2115 = n2111 & n2112;
  assign n2116 = n506 & n898;
  assign n2117 = n925 & n1012;
  assign n2118 = n1672 & n2108;
  assign n2119 = n2117 & n2118;
  assign n2120 = n2115 & n2116;
  assign n2121 = n2114 & n2120;
  assign n2122 = n1798 & n2119;
  assign n2123 = n2110 & n2122;
  assign n2124 = n1763 & n2121;
  assign n2125 = n2123 & n2124;
  assign n2126 = ~n841 & ~n893;
  assign n2127 = ~n339 & ~n439;
  assign n2128 = ~n770 & n2127;
  assign n2129 = ~n278 & ~n355;
  assign n2130 = n1478 & n2129;
  assign n2131 = n2126 & n2130;
  assign n2132 = n2128 & n2131;
  assign n2133 = ~n183 & ~n427;
  assign n2134 = ~n525 & ~n700;
  assign n2135 = ~n1487 & n2134;
  assign n2136 = n1014 & n2133;
  assign n2137 = n1403 & n2136;
  assign n2138 = n1918 & n2135;
  assign n2139 = n2105 & n2107;
  assign n2140 = n2138 & n2139;
  assign n2141 = n2102 & n2137;
  assign n2142 = n2140 & n2141;
  assign n2143 = n1823 & n2132;
  assign n2144 = n2142 & n2143;
  assign n2145 = n2019 & n2144;
  assign n2146 = n2125 & n2145;
  assign n2147 = ~n2098 & ~n2146;
  assign n2148 = ~n93 & ~n718;
  assign n2149 = ~n284 & n424;
  assign n2150 = ~n123 & ~n211;
  assign n2151 = ~n243 & ~n259;
  assign n2152 = ~n902 & n2151;
  assign n2153 = n2007 & n2150;
  assign n2154 = n2148 & n2153;
  assign n2155 = n2149 & n2152;
  assign n2156 = n2154 & n2155;
  assign n2157 = ~n536 & ~n937;
  assign n2158 = ~n380 & ~n700;
  assign n2159 = ~n459 & n2158;
  assign n2160 = ~n526 & ~n724;
  assign n2161 = ~n753 & n2160;
  assign n2162 = ~n235 & ~n488;
  assign n2163 = ~n510 & ~n687;
  assign n2164 = ~n703 & n2163;
  assign n2165 = n2162 & n2164;
  assign n2166 = n2161 & n2165;
  assign n2167 = ~n143 & ~n333;
  assign n2168 = ~n427 & ~n460;
  assign n2169 = ~n599 & ~n663;
  assign n2170 = ~n156 & ~n378;
  assign n2171 = n2168 & n2169;
  assign n2172 = n2170 & n2171;
  assign n2173 = ~n300 & ~n302;
  assign n2174 = ~n352 & ~n359;
  assign n2175 = n2173 & n2174;
  assign n2176 = n1779 & n2157;
  assign n2177 = n2167 & n2176;
  assign n2178 = n118 & n2175;
  assign n2179 = n2159 & n2178;
  assign n2180 = n2172 & n2177;
  assign n2181 = n2179 & n2180;
  assign n2182 = n2156 & n2166;
  assign n2183 = n2181 & n2182;
  assign n2184 = ~n247 & ~n537;
  assign n2185 = ~n648 & ~n1487;
  assign n2186 = n2184 & n2185;
  assign n2187 = ~n269 & ~n604;
  assign n2188 = ~n754 & ~n810;
  assign n2189 = n2187 & n2188;
  assign n2190 = n137 & n2189;
  assign n2191 = n2186 & n2190;
  assign n2192 = ~n368 & ~n373;
  assign n2193 = ~n318 & ~n518;
  assign n2194 = n1306 & n2193;
  assign n2195 = ~n293 & ~n408;
  assign n2196 = n1357 & n2195;
  assign n2197 = ~n253 & ~n798;
  assign n2198 = ~n486 & n1123;
  assign n2199 = n2197 & n2198;
  assign n2200 = ~n282 & ~n605;
  assign n2201 = ~n236 & ~n627;
  assign n2202 = ~n317 & ~n723;
  assign n2203 = ~n751 & ~n893;
  assign n2204 = n2202 & n2203;
  assign n2205 = n1420 & n2204;
  assign n2206 = ~n376 & ~n480;
  assign n2207 = ~n159 & ~n653;
  assign n2208 = ~n148 & ~n476;
  assign n2209 = ~n120 & ~n308;
  assign n2210 = ~n432 & ~n634;
  assign n2211 = n2209 & n2210;
  assign n2212 = n413 & n722;
  assign n2213 = n1308 & n2208;
  assign n2214 = n2212 & n2213;
  assign n2215 = n1726 & n2211;
  assign n2216 = n1781 & n2215;
  assign n2217 = n2214 & n2216;
  assign n2218 = ~n151 & ~n310;
  assign n2219 = ~n332 & ~n370;
  assign n2220 = ~n841 & n2219;
  assign n2221 = n533 & n2218;
  assign n2222 = n2024 & n2200;
  assign n2223 = n2201 & n2206;
  assign n2224 = n2207 & n2223;
  assign n2225 = n2221 & n2222;
  assign n2226 = n1455 & n2220;
  assign n2227 = n2194 & n2196;
  assign n2228 = n2226 & n2227;
  assign n2229 = n2224 & n2225;
  assign n2230 = n2199 & n2205;
  assign n2231 = n2229 & n2230;
  assign n2232 = n2228 & n2231;
  assign n2233 = n2217 & n2232;
  assign n2234 = ~n252 & ~n358;
  assign n2235 = ~n568 & ~n597;
  assign n2236 = ~n838 & ~n922;
  assign n2237 = n2235 & n2236;
  assign n2238 = n298 & n423;
  assign n2239 = n513 & ~n535;
  assign n2240 = n2192 & n2234;
  assign n2241 = n2239 & n2240;
  assign n2242 = n2237 & n2238;
  assign n2243 = n2109 & n2242;
  assign n2244 = n1724 & n2241;
  assign n2245 = n2243 & n2244;
  assign n2246 = n2191 & n2245;
  assign n2247 = n210 & n2246;
  assign n2248 = n2183 & n2247;
  assign n2249 = n2233 & n2248;
  assign n2250 = ~n2146 & ~n2249;
  assign n2251 = ~n511 & ~n529;
  assign n2252 = ~n700 & n2251;
  assign n2253 = ~n518 & ~n768;
  assign n2254 = ~n373 & ~n634;
  assign n2255 = ~n435 & ~n1699;
  assign n2256 = n2253 & n2255;
  assign n2257 = n2254 & n2256;
  assign n2258 = ~n422 & ~n510;
  assign n2259 = n448 & n2258;
  assign n2260 = ~n382 & ~n414;
  assign n2261 = ~n685 & ~n902;
  assign n2262 = n2260 & n2261;
  assign n2263 = ~n175 & ~n327;
  assign n2264 = n1428 & n2263;
  assign n2265 = ~n141 & ~n238;
  assign n2266 = ~n564 & ~n638;
  assign n2267 = n2265 & n2266;
  assign n2268 = n759 & n777;
  assign n2269 = n1403 & n2268;
  assign n2270 = n2252 & n2267;
  assign n2271 = n2259 & n2262;
  assign n2272 = n2264 & n2271;
  assign n2273 = n2269 & n2270;
  assign n2274 = n1825 & n2257;
  assign n2275 = n2273 & n2274;
  assign n2276 = n2272 & n2275;
  assign n2277 = ~n294 & ~n380;
  assign n2278 = ~n432 & n2277;
  assign n2279 = ~n250 & ~n1034;
  assign n2280 = ~n247 & ~n290;
  assign n2281 = ~n753 & ~n814;
  assign n2282 = n172 & n2281;
  assign n2283 = ~n120 & ~n362;
  assign n2284 = ~n411 & ~n703;
  assign n2285 = ~n274 & ~n339;
  assign n2286 = ~n477 & n2285;
  assign n2287 = n2040 & n2283;
  assign n2288 = n2284 & n2287;
  assign n2289 = n2105 & n2286;
  assign n2290 = n2282 & n2289;
  assign n2291 = n2288 & n2290;
  assign n2292 = ~n526 & ~n1002;
  assign n2293 = ~n1404 & n2292;
  assign n2294 = ~n111 & ~n278;
  assign n2295 = ~n525 & ~n661;
  assign n2296 = n2294 & n2295;
  assign n2297 = n298 & n1296;
  assign n2298 = n1864 & n2279;
  assign n2299 = n2280 & n2298;
  assign n2300 = n2296 & n2297;
  assign n2301 = n882 & n2008;
  assign n2302 = n2054 & n2293;
  assign n2303 = n2301 & n2302;
  assign n2304 = n2299 & n2300;
  assign n2305 = n2303 & n2304;
  assign n2306 = n2291 & n2305;
  assign n2307 = ~n188 & n1424;
  assign n2308 = n2306 & n2307;
  assign n2309 = ~n180 & ~n308;
  assign n2310 = ~n213 & ~n291;
  assign n2311 = ~n508 & ~n520;
  assign n2312 = ~n563 & ~n566;
  assign n2313 = ~n596 & ~n944;
  assign n2314 = n2312 & n2313;
  assign n2315 = n2310 & n2311;
  assign n2316 = n1387 & n1812;
  assign n2317 = n2309 & n2316;
  assign n2318 = n2314 & n2315;
  assign n2319 = n2317 & n2318;
  assign n2320 = ~n153 & ~n353;
  assign n2321 = ~n200 & ~n356;
  assign n2322 = ~n480 & n2321;
  assign n2323 = ~n523 & ~n537;
  assign n2324 = ~n328 & ~n416;
  assign n2325 = n2323 & n2324;
  assign n2326 = ~n318 & ~n365;
  assign n2327 = n797 & n2326;
  assign n2328 = n2320 & n2327;
  assign n2329 = n2322 & n2325;
  assign n2330 = n2328 & n2329;
  assign n2331 = ~n317 & ~n358;
  assign n2332 = ~n486 & ~n810;
  assign n2333 = n2331 & n2332;
  assign n2334 = ~n143 & ~n197;
  assign n2335 = ~n512 & ~n539;
  assign n2336 = ~n561 & ~n604;
  assign n2337 = n2335 & n2336;
  assign n2338 = n528 & n2334;
  assign n2339 = n1306 & n1354;
  assign n2340 = n2338 & n2339;
  assign n2341 = n2278 & n2337;
  assign n2342 = n2333 & n2341;
  assign n2343 = n2340 & n2342;
  assign n2344 = n2319 & n2330;
  assign n2345 = n2343 & n2344;
  assign n2346 = n2276 & n2345;
  assign n2347 = n2308 & n2346;
  assign n2348 = ~n2249 & ~n2347;
  assign n2349 = ~n723 & ~n894;
  assign n2350 = ~n313 & ~n525;
  assign n2351 = ~n663 & ~n846;
  assign n2352 = ~n1032 & n2351;
  assign n2353 = n1865 & n2349;
  assign n2354 = n2350 & n2353;
  assign n2355 = n2352 & n2354;
  assign n2356 = ~n249 & ~n596;
  assign n2357 = ~n1051 & n2356;
  assign n2358 = ~n438 & ~n499;
  assign n2359 = ~n333 & ~n661;
  assign n2360 = ~n242 & ~n561;
  assign n2361 = ~n273 & ~n319;
  assign n2362 = ~n377 & ~n531;
  assign n2363 = ~n599 & n2362;
  assign n2364 = n1456 & n2360;
  assign n2365 = n2361 & n2364;
  assign n2366 = n2363 & n2365;
  assign n2367 = n2257 & n2366;
  assign n2368 = ~n258 & ~n526;
  assign n2369 = ~n1487 & n2368;
  assign n2370 = ~n443 & ~n841;
  assign n2371 = ~n235 & ~n378;
  assign n2372 = n895 & n2371;
  assign n2373 = n938 & n2358;
  assign n2374 = n2359 & n2370;
  assign n2375 = n2373 & n2374;
  assign n2376 = n2357 & n2372;
  assign n2377 = n2369 & n2376;
  assign n2378 = n2375 & n2377;
  assign n2379 = n2355 & n2378;
  assign n2380 = n2367 & n2379;
  assign n2381 = ~n312 & ~n411;
  assign n2382 = ~n509 & ~n515;
  assign n2383 = ~n787 & ~n808;
  assign n2384 = ~n1086 & ~n1404;
  assign n2385 = n2383 & n2384;
  assign n2386 = n2381 & n2382;
  assign n2387 = n1494 & n1948;
  assign n2388 = n2386 & n2387;
  assign n2389 = n2385 & n2388;
  assign n2390 = ~n269 & ~n724;
  assign n2391 = ~n893 & n2390;
  assign n2392 = n654 & n1049;
  assign n2393 = n1151 & n2392;
  assign n2394 = n2391 & n2393;
  assign n2395 = ~n532 & ~n594;
  assign n2396 = ~n460 & n2395;
  assign n2397 = ~n238 & ~n603;
  assign n2398 = n593 & ~n814;
  assign n2399 = ~n481 & ~n751;
  assign n2400 = ~n380 & ~n754;
  assign n2401 = n565 & n2400;
  assign n2402 = n1384 & n2258;
  assign n2403 = n2397 & n2399;
  assign n2404 = n2402 & n2403;
  assign n2405 = n2396 & n2401;
  assign n2406 = n2398 & n2405;
  assign n2407 = n2404 & n2406;
  assign n2408 = n1649 & n2389;
  assign n2409 = n2394 & n2408;
  assign n2410 = n2407 & n2409;
  assign n2411 = n234 & n2410;
  assign n2412 = n2380 & n2411;
  assign n2413 = ~n2347 & ~n2412;
  assign n2414 = ~n237 & ~n476;
  assign n2415 = ~n653 & n2414;
  assign n2416 = ~n361 & n1767;
  assign n2417 = ~n276 & ~n293;
  assign n2418 = ~n317 & n2417;
  assign n2419 = n357 & n1014;
  assign n2420 = n1047 & n2419;
  assign n2421 = n1455 & n2418;
  assign n2422 = n2416 & n2421;
  assign n2423 = n2420 & n2422;
  assign n2424 = ~n310 & ~n446;
  assign n2425 = ~n458 & ~n502;
  assign n2426 = n2424 & n2425;
  assign n2427 = n369 & n500;
  assign n2428 = n895 & n1244;
  assign n2429 = n1270 & n1779;
  assign n2430 = n2428 & n2429;
  assign n2431 = n2426 & n2427;
  assign n2432 = n2282 & n2415;
  assign n2433 = n2431 & n2432;
  assign n2434 = n2430 & n2433;
  assign n2435 = n2423 & n2434;
  assign n2436 = ~n93 & ~n189;
  assign n2437 = ~n416 & ~n594;
  assign n2438 = n2436 & n2437;
  assign n2439 = ~n141 & ~n687;
  assign n2440 = n722 & n2439;
  assign n2441 = ~n212 & ~n327;
  assign n2442 = ~n518 & ~n718;
  assign n2443 = ~n893 & n2442;
  assign n2444 = n2441 & n2443;
  assign n2445 = ~n149 & ~n509;
  assign n2446 = ~n370 & ~n535;
  assign n2447 = n244 & n2446;
  assign n2448 = n2445 & n2447;
  assign n2449 = ~n183 & ~n353;
  assign n2450 = ~n944 & n2449;
  assign n2451 = ~n130 & ~n894;
  assign n2452 = ~n194 & ~n792;
  assign n2453 = ~n252 & ~n274;
  assign n2454 = ~n523 & ~n810;
  assign n2455 = n2453 & n2454;
  assign n2456 = n1489 & n2451;
  assign n2457 = n2452 & n2456;
  assign n2458 = n2455 & n2457;
  assign n2459 = ~n258 & ~n412;
  assign n2460 = ~n373 & ~n380;
  assign n2461 = ~n126 & ~n430;
  assign n2462 = ~n638 & ~n922;
  assign n2463 = n2461 & n2462;
  assign n2464 = n1019 & n1622;
  assign n2465 = n2459 & n2460;
  assign n2466 = n2464 & n2465;
  assign n2467 = n2450 & n2463;
  assign n2468 = n2466 & n2467;
  assign n2469 = n2444 & n2448;
  assign n2470 = n2468 & n2469;
  assign n2471 = n2458 & n2470;
  assign n2472 = ~n334 & ~n592;
  assign n2473 = ~n304 & ~n723;
  assign n2474 = ~n510 & ~n754;
  assign n2475 = ~n566 & ~n703;
  assign n2476 = ~n798 & ~n1487;
  assign n2477 = n2475 & n2476;
  assign n2478 = n2474 & n2477;
  assign n2479 = ~n174 & ~n213;
  assign n2480 = ~n432 & ~n460;
  assign n2481 = ~n563 & n2480;
  assign n2482 = n187 & n2479;
  assign n2483 = n540 & n1186;
  assign n2484 = n1245 & n1575;
  assign n2485 = n2206 & n2472;
  assign n2486 = n2473 & n2485;
  assign n2487 = n2483 & n2484;
  assign n2488 = n2481 & n2482;
  assign n2489 = n2438 & n2440;
  assign n2490 = n2488 & n2489;
  assign n2491 = n2486 & n2487;
  assign n2492 = n2478 & n2491;
  assign n2493 = n1791 & n2490;
  assign n2494 = n2492 & n2493;
  assign n2495 = n2435 & n2494;
  assign n2496 = n2471 & n2495;
  assign n2497 = ~n2412 & ~n2496;
  assign n2498 = ~n520 & ~n798;
  assign n2499 = n2452 & n2498;
  assign n2500 = ~n432 & ~n446;
  assign n2501 = ~n248 & ~n535;
  assign n2502 = ~n120 & ~n367;
  assign n2503 = ~n215 & ~n656;
  assign n2504 = ~n212 & ~n297;
  assign n2505 = ~n371 & n2504;
  assign n2506 = n2503 & n2505;
  assign n2507 = ~n376 & ~n605;
  assign n2508 = ~n787 & ~n902;
  assign n2509 = n2507 & n2508;
  assign n2510 = n301 & n598;
  assign n2511 = n1033 & n2500;
  assign n2512 = n2501 & n2502;
  assign n2513 = n2511 & n2512;
  assign n2514 = n2509 & n2510;
  assign n2515 = n2325 & n2499;
  assign n2516 = n2514 & n2515;
  assign n2517 = n921 & n2513;
  assign n2518 = n2506 & n2517;
  assign n2519 = n2516 & n2518;
  assign n2520 = ~n175 & ~n361;
  assign n2521 = ~n700 & n2520;
  assign n2522 = ~n370 & ~n374;
  assign n2523 = ~n808 & n2522;
  assign n2524 = n192 & n2523;
  assign n2525 = n2521 & n2524;
  assign n2526 = ~n159 & ~n296;
  assign n2527 = n755 & n2526;
  assign n2528 = ~n427 & ~n814;
  assign n2529 = ~n482 & ~n561;
  assign n2530 = ~n183 & ~n239;
  assign n2531 = ~n381 & n2530;
  assign n2532 = n1845 & n2531;
  assign n2533 = ~n156 & n1814;
  assign n2534 = ~n430 & ~n564;
  assign n2535 = ~n111 & ~n155;
  assign n2536 = ~n249 & ~n353;
  assign n2537 = ~n422 & ~n477;
  assign n2538 = ~n1699 & n2537;
  assign n2539 = n2535 & n2536;
  assign n2540 = n802 & n1859;
  assign n2541 = n2534 & n2540;
  assign n2542 = n2538 & n2539;
  assign n2543 = n2396 & n2533;
  assign n2544 = n2542 & n2543;
  assign n2545 = n2541 & n2544;
  assign n2546 = ~n283 & ~n412;
  assign n2547 = ~n499 & n2546;
  assign n2548 = ~n277 & ~n459;
  assign n2549 = ~n768 & ~n989;
  assign n2550 = n2548 & n2549;
  assign n2551 = ~n685 & ~n770;
  assign n2552 = n311 & n2551;
  assign n2553 = n1755 & n2528;
  assign n2554 = n2529 & n2553;
  assign n2555 = n2547 & n2552;
  assign n2556 = n2550 & n2555;
  assign n2557 = n2532 & n2554;
  assign n2558 = n2556 & n2557;
  assign n2559 = n1129 & n2558;
  assign n2560 = n2545 & n2559;
  assign n2561 = ~n177 & ~n255;
  assign n2562 = ~n123 & ~n294;
  assign n2563 = ~n639 & ~n839;
  assign n2564 = ~n1034 & n2563;
  assign n2565 = n2037 & n2562;
  assign n2566 = n2167 & n2361;
  assign n2567 = n2561 & n2566;
  assign n2568 = n2564 & n2565;
  assign n2569 = n2567 & n2568;
  assign n2570 = n2560 & n2569;
  assign n2571 = ~n256 & ~n596;
  assign n2572 = ~n338 & ~n414;
  assign n2573 = ~n698 & ~n944;
  assign n2574 = n2572 & n2573;
  assign n2575 = n2571 & n2574;
  assign n2576 = ~n246 & ~n252;
  assign n2577 = ~n271 & ~n476;
  assign n2578 = ~n715 & n2577;
  assign n2579 = n1012 & n2576;
  assign n2580 = n1017 & n1347;
  assign n2581 = n1752 & n2580;
  assign n2582 = n2578 & n2579;
  assign n2583 = n1698 & n2527;
  assign n2584 = n2582 & n2583;
  assign n2585 = n2575 & n2581;
  assign n2586 = n2584 & n2585;
  assign n2587 = n2525 & n2586;
  assign n2588 = n2519 & n2587;
  assign n2589 = n2570 & n2588;
  assign n2590 = ~n2496 & ~n2589;
  assign n2591 = ~n480 & ~n627;
  assign n2592 = ~n141 & ~n283;
  assign n2593 = ~n1051 & n2592;
  assign n2594 = n2591 & n2593;
  assign n2595 = ~n149 & ~n359;
  assign n2596 = ~n703 & n2595;
  assign n2597 = ~n277 & ~n653;
  assign n2598 = ~n634 & n816;
  assign n2599 = n421 & n686;
  assign n2600 = n785 & n1387;
  assign n2601 = n2597 & n2600;
  assign n2602 = n2598 & n2599;
  assign n2603 = n1137 & n2596;
  assign n2604 = n2602 & n2603;
  assign n2605 = n2594 & n2601;
  assign n2606 = n2604 & n2605;
  assign n2607 = n1970 & n2606;
  assign n2608 = ~n171 & ~n332;
  assign n2609 = ~n687 & ~n753;
  assign n2610 = ~n355 & ~n371;
  assign n2611 = ~n151 & ~n328;
  assign n2612 = ~n339 & n2611;
  assign n2613 = n1864 & n2571;
  assign n2614 = n2608 & n2609;
  assign n2615 = n2610 & n2614;
  assign n2616 = n2612 & n2613;
  assign n2617 = n783 & n2616;
  assign n2618 = n2615 & n2617;
  assign n2619 = ~n130 & ~n374;
  assign n2620 = ~n379 & ~n648;
  assign n2621 = n801 & n2620;
  assign n2622 = n1053 & n2619;
  assign n2623 = n2621 & n2622;
  assign n2624 = ~n300 & ~n376;
  assign n2625 = ~n255 & ~n539;
  assign n2626 = ~n148 & ~n167;
  assign n2627 = ~n250 & ~n422;
  assign n2628 = ~n488 & ~n718;
  assign n2629 = ~n841 & n2628;
  assign n2630 = n2626 & n2627;
  assign n2631 = n1272 & n2529;
  assign n2632 = n2624 & n2625;
  assign n2633 = n2631 & n2632;
  assign n2634 = n2629 & n2630;
  assign n2635 = n2633 & n2634;
  assign n2636 = ~n111 & ~n120;
  assign n2637 = ~n382 & ~n518;
  assign n2638 = ~n700 & ~n1002;
  assign n2639 = n2637 & n2638;
  assign n2640 = n428 & n2636;
  assign n2641 = n478 & n530;
  assign n2642 = n705 & n941;
  assign n2643 = n1244 & n2642;
  assign n2644 = n2640 & n2641;
  assign n2645 = n2639 & n2644;
  assign n2646 = n2623 & n2643;
  assign n2647 = n2645 & n2646;
  assign n2648 = n2635 & n2647;
  assign n2649 = ~n188 & ~n243;
  assign n2650 = n2648 & n2649;
  assign n2651 = ~n159 & ~n303;
  assign n2652 = ~n439 & ~n502;
  assign n2653 = ~n537 & ~n563;
  assign n2654 = n2652 & n2653;
  assign n2655 = n2651 & n2654;
  assign n2656 = ~n358 & ~n435;
  assign n2657 = ~n768 & n2656;
  assign n2658 = ~n698 & ~n1404;
  assign n2659 = ~n294 & ~n310;
  assign n2660 = ~n536 & ~n798;
  assign n2661 = n2659 & n2660;
  assign n2662 = n164 & n602;
  assign n2663 = n644 & n1049;
  assign n2664 = n1357 & n1751;
  assign n2665 = n2658 & n2664;
  assign n2666 = n2662 & n2663;
  assign n2667 = n2657 & n2661;
  assign n2668 = n2666 & n2667;
  assign n2669 = n1427 & n2665;
  assign n2670 = n2655 & n2669;
  assign n2671 = n2668 & n2670;
  assign n2672 = n2618 & n2671;
  assign n2673 = n2607 & n2672;
  assign n2674 = n2650 & n2673;
  assign n2675 = ~n2589 & ~n2674;
  assign n2676 = ~n318 & ~n438;
  assign n2677 = ~n566 & ~n639;
  assign n2678 = n2676 & n2677;
  assign n2679 = ~n313 & ~n532;
  assign n2680 = ~n539 & n2679;
  assign n2681 = n2678 & n2680;
  assign n2682 = ~n625 & ~n792;
  assign n2683 = ~n153 & n1650;
  assign n2684 = n2682 & n2683;
  assign n2685 = ~n145 & ~n277;
  assign n2686 = ~n237 & ~n310;
  assign n2687 = n2685 & n2686;
  assign n2688 = ~n163 & ~n281;
  assign n2689 = ~n319 & n2688;
  assign n2690 = ~n408 & ~n416;
  assign n2691 = ~n291 & n363;
  assign n2692 = n2207 & n2279;
  assign n2693 = n2690 & n2692;
  assign n2694 = n2691 & n2693;
  assign n2695 = ~n273 & ~n379;
  assign n2696 = ~n511 & n2695;
  assign n2697 = n1245 & n1355;
  assign n2698 = n2397 & n2697;
  assign n2699 = n2547 & n2696;
  assign n2700 = n2687 & n2689;
  assign n2701 = n2699 & n2700;
  assign n2702 = n2681 & n2698;
  assign n2703 = n2684 & n2702;
  assign n2704 = n2132 & n2701;
  assign n2705 = n2694 & n2704;
  assign n2706 = n2703 & n2705;
  assign n2707 = n1984 & n2183;
  assign n2708 = n2706 & n2707;
  assign n2709 = ~n2674 & ~n2708;
  assign n2710 = ~n93 & ~n627;
  assign n2711 = ~n193 & ~n605;
  assign n2712 = ~n685 & n1420;
  assign n2713 = n2711 & n2712;
  assign n2714 = ~n189 & ~n502;
  assign n2715 = n172 & n2714;
  assign n2716 = n565 & n1389;
  assign n2717 = n1890 & n2710;
  assign n2718 = n2716 & n2717;
  assign n2719 = n2715 & n2718;
  assign n2720 = n2713 & n2719;
  assign n2721 = ~n174 & ~n459;
  assign n2722 = ~n534 & n2721;
  assign n2723 = ~n318 & ~n415;
  assign n2724 = ~n1487 & n2723;
  assign n2725 = ~n136 & ~n196;
  assign n2726 = ~n242 & ~n355;
  assign n2727 = ~n368 & ~n414;
  assign n2728 = ~n532 & ~n1086;
  assign n2729 = n2727 & n2728;
  assign n2730 = n2725 & n2726;
  assign n2731 = n752 & n1914;
  assign n2732 = n1947 & n2731;
  assign n2733 = n2729 & n2730;
  assign n2734 = n1119 & n2722;
  assign n2735 = n2724 & n2734;
  assign n2736 = n2732 & n2733;
  assign n2737 = n2735 & n2736;
  assign n2738 = n2720 & n2737;
  assign n2739 = ~n155 & ~n211;
  assign n2740 = ~n365 & ~n438;
  assign n2741 = ~n445 & ~n515;
  assign n2742 = ~n518 & ~n561;
  assign n2743 = ~n656 & n2742;
  assign n2744 = n2740 & n2741;
  assign n2745 = n2739 & n2744;
  assign n2746 = n2743 & n2745;
  assign n2747 = n331 & n1165;
  assign n2748 = n1539 & n2108;
  assign n2749 = ~n168 & ~n184;
  assign n2750 = ~n293 & ~n358;
  assign n2751 = ~n526 & n2750;
  assign n2752 = n1767 & n2749;
  assign n2753 = n1864 & n2752;
  assign n2754 = n1197 & n2751;
  assign n2755 = n2748 & n2754;
  assign n2756 = n2753 & n2755;
  assign n2757 = ~n296 & ~n422;
  assign n2758 = ~n312 & n2206;
  assign n2759 = n2280 & n2758;
  assign n2760 = ~n163 & ~n167;
  assign n2761 = ~n235 & ~n258;
  assign n2762 = ~n512 & ~n634;
  assign n2763 = ~n754 & ~n792;
  assign n2764 = n2762 & n2763;
  assign n2765 = n2760 & n2761;
  assign n2766 = n785 & n1003;
  assign n2767 = n1186 & n1351;
  assign n2768 = n1673 & n1884;
  assign n2769 = n2757 & n2768;
  assign n2770 = n2766 & n2767;
  assign n2771 = n2764 & n2765;
  assign n2772 = n2770 & n2771;
  assign n2773 = n2759 & n2769;
  assign n2774 = n2772 & n2773;
  assign n2775 = n2746 & n2774;
  assign n2776 = n2756 & n2775;
  assign n2777 = n2738 & n2776;
  assign n2778 = n2747 & n2777;
  assign n2779 = ~n2708 & ~n2778;
  assign n2780 = ~n297 & ~n309;
  assign n2781 = ~n1699 & n2780;
  assign n2782 = ~n126 & ~n200;
  assign n2783 = ~n365 & ~n511;
  assign n2784 = ~n376 & ~n481;
  assign n2785 = n631 & n2784;
  assign n2786 = n1492 & n1813;
  assign n2787 = n2782 & n2783;
  assign n2788 = n2786 & n2787;
  assign n2789 = n2689 & n2785;
  assign n2790 = n2781 & n2789;
  assign n2791 = n2788 & n2790;
  assign n2792 = ~n153 & ~n197;
  assign n2793 = ~n148 & ~n374;
  assign n2794 = n2792 & n2793;
  assign n2795 = ~n685 & n1474;
  assign n2796 = n1913 & n2795;
  assign n2797 = ~n362 & ~n1086;
  assign n2798 = n176 & ~n724;
  assign n2799 = n1175 & n2797;
  assign n2800 = n2798 & n2799;
  assign n2801 = ~n136 & ~n149;
  assign n2802 = ~n312 & ~n838;
  assign n2803 = ~n568 & ~n839;
  assign n2804 = n2802 & n2803;
  assign n2805 = ~n199 & ~n253;
  assign n2806 = ~n703 & ~n841;
  assign n2807 = ~n922 & n2806;
  assign n2808 = n117 & n2805;
  assign n2809 = n1291 & n1321;
  assign n2810 = n1430 & n2167;
  assign n2811 = n2534 & n2801;
  assign n2812 = n2810 & n2811;
  assign n2813 = n2808 & n2809;
  assign n2814 = n1541 & n2807;
  assign n2815 = n2804 & n2814;
  assign n2816 = n2812 & n2813;
  assign n2817 = n2532 & n2816;
  assign n2818 = n2815 & n2817;
  assign n2819 = ~n139 & ~n274;
  assign n2820 = ~n303 & ~n488;
  assign n2821 = ~n512 & ~n531;
  assign n2822 = ~n599 & ~n754;
  assign n2823 = n2821 & n2822;
  assign n2824 = n2819 & n2820;
  assign n2825 = n799 & n2108;
  assign n2826 = n2591 & n2825;
  assign n2827 = n2823 & n2824;
  assign n2828 = n2794 & n2827;
  assign n2829 = n1191 & n2826;
  assign n2830 = n2796 & n2800;
  assign n2831 = n2829 & n2830;
  assign n2832 = n2828 & n2831;
  assign n2833 = n2791 & n2832;
  assign n2834 = n2435 & n2818;
  assign n2835 = n2833 & n2834;
  assign n2836 = ~n2778 & ~n2835;
  assign n2837 = ~n841 & ~n846;
  assign n2838 = ~n250 & ~n1051;
  assign n2839 = ~n194 & ~n294;
  assign n2840 = ~n145 & ~n180;
  assign n2841 = ~n238 & ~n338;
  assign n2842 = ~n438 & ~n718;
  assign n2843 = ~n810 & n2842;
  assign n2844 = n2840 & n2841;
  assign n2845 = n179 & n1272;
  assign n2846 = n2839 & n2845;
  assign n2847 = n2843 & n2844;
  assign n2848 = n2846 & n2847;
  assign n2849 = ~n174 & ~n989;
  assign n2850 = n657 & n2849;
  assign n2851 = ~n126 & ~n721;
  assign n2852 = ~n1034 & n2851;
  assign n2853 = n2206 & n2208;
  assign n2854 = n2852 & n2853;
  assign n2855 = ~n183 & ~n216;
  assign n2856 = ~n379 & ~n601;
  assign n2857 = n2855 & n2856;
  assign n2858 = n785 & n1011;
  assign n2859 = n1134 & n1730;
  assign n2860 = n2052 & n2859;
  assign n2861 = n2857 & n2858;
  assign n2862 = n783 & n1844;
  assign n2863 = n2850 & n2862;
  assign n2864 = n2860 & n2861;
  assign n2865 = n2854 & n2864;
  assign n2866 = n2848 & n2863;
  assign n2867 = n2865 & n2866;
  assign n2868 = ~n333 & ~n723;
  assign n2869 = ~n352 & ~n435;
  assign n2870 = ~n443 & ~n523;
  assign n2871 = ~n605 & ~n625;
  assign n2872 = n2870 & n2871;
  assign n2873 = n2868 & n2869;
  assign n2874 = n2872 & n2873;
  assign n2875 = ~n123 & ~n656;
  assign n2876 = n448 & n2875;
  assign n2877 = ~n303 & ~n310;
  assign n2878 = ~n409 & n2877;
  assign n2879 = n363 & n1237;
  assign n2880 = n1283 & n1291;
  assign n2881 = n1470 & n1962;
  assign n2882 = n2040 & n2881;
  assign n2883 = n2879 & n2880;
  assign n2884 = n2438 & n2878;
  assign n2885 = n2876 & n2884;
  assign n2886 = n2882 & n2883;
  assign n2887 = n2874 & n2886;
  assign n2888 = n2885 & n2887;
  assign n2889 = ~n129 & ~n328;
  assign n2890 = n160 & ~n312;
  assign n2891 = ~n141 & ~n291;
  assign n2892 = ~n168 & ~n685;
  assign n2893 = ~n239 & ~n648;
  assign n2894 = ~n715 & n2893;
  assign n2895 = n504 & n1230;
  assign n2896 = n2193 & n2889;
  assign n2897 = n2891 & n2892;
  assign n2898 = n2896 & n2897;
  assign n2899 = n2894 & n2895;
  assign n2900 = n2890 & n2899;
  assign n2901 = n2898 & n2900;
  assign n2902 = ~n193 & ~n213;
  assign n2903 = ~n334 & ~n412;
  assign n2904 = ~n427 & ~n499;
  assign n2905 = ~n534 & ~n698;
  assign n2906 = n2904 & n2905;
  assign n2907 = n2902 & n2903;
  assign n2908 = n369 & n375;
  assign n2909 = n1175 & n1576;
  assign n2910 = n2837 & n2838;
  assign n2911 = n2909 & n2910;
  assign n2912 = n2907 & n2908;
  assign n2913 = n2906 & n2912;
  assign n2914 = n643 & n2911;
  assign n2915 = n2199 & n2914;
  assign n2916 = n2913 & n2915;
  assign n2917 = n2901 & n2916;
  assign n2918 = n2867 & n2888;
  assign n2919 = n2917 & n2918;
  assign n2920 = ~n2835 & ~n2919;
  assign n2921 = ~n370 & ~n503;
  assign n2922 = n384 & ~n846;
  assign n2923 = n1476 & n1753;
  assign n2924 = n2921 & n2923;
  assign n2925 = n2259 & n2922;
  assign n2926 = n2924 & n2925;
  assign n2927 = n659 & n2172;
  assign n2928 = n2681 & n2927;
  assign n2929 = n2926 & n2928;
  assign n2930 = n784 & n840;
  assign n2931 = n1754 & n2930;
  assign n2932 = ~n168 & ~n243;
  assign n2933 = ~n627 & n2932;
  assign n2934 = ~n239 & ~n893;
  assign n2935 = ~n151 & n375;
  assign n2936 = n2934 & n2935;
  assign n2937 = n500 & ~n597;
  assign n2938 = n2687 & n2937;
  assign n2939 = ~n248 & ~n515;
  assign n2940 = n1423 & n2939;
  assign n2941 = n1575 & n2207;
  assign n2942 = n2534 & n2941;
  assign n2943 = n2933 & n2940;
  assign n2944 = n2942 & n2943;
  assign n2945 = n1683 & n1770;
  assign n2946 = n2931 & n2936;
  assign n2947 = n2938 & n2946;
  assign n2948 = n2944 & n2945;
  assign n2949 = n2947 & n2948;
  assign n2950 = n2929 & n2949;
  assign n2951 = n2308 & n2950;
  assign n2952 = ~n2919 & ~n2951;
  assign n2953 = ~n380 & ~n944;
  assign n2954 = n1151 & n2953;
  assign n2955 = ~n199 & ~n416;
  assign n2956 = n899 & n2955;
  assign n2957 = n1547 & n2954;
  assign n2958 = n2956 & n2957;
  assign n2959 = n1173 & n2958;
  assign n2960 = ~n299 & ~n319;
  assign n2961 = n2959 & n2960;
  assign n2962 = ~n116 & ~n184;
  assign n2963 = ~n290 & ~n476;
  assign n2964 = ~n563 & n2963;
  assign n2965 = n164 & n799;
  assign n2966 = n2962 & n2965;
  assign n2967 = n2964 & n2966;
  assign n2968 = ~n536 & ~n814;
  assign n2969 = ~n1051 & n2968;
  assign n2970 = n1650 & n2625;
  assign n2971 = n2969 & n2970;
  assign n2972 = ~n247 & ~n332;
  assign n2973 = ~n596 & n1350;
  assign n2974 = n1509 & n1782;
  assign n2975 = n2972 & n2974;
  assign n2976 = n2724 & n2973;
  assign n2977 = n2975 & n2976;
  assign n2978 = ~n246 & ~n1032;
  assign n2979 = n1428 & n2978;
  assign n2980 = ~n167 & ~n245;
  assign n2981 = ~n371 & ~n480;
  assign n2982 = n2980 & n2981;
  assign n2983 = ~n358 & ~n373;
  assign n2984 = ~n382 & ~n639;
  assign n2985 = n1305 & n2984;
  assign n2986 = n1663 & n1771;
  assign n2987 = n2891 & n2983;
  assign n2988 = n2986 & n2987;
  assign n2989 = n2985 & n2988;
  assign n2990 = n2058 & n2989;
  assign n2991 = ~n216 & ~n277;
  assign n2992 = ~n432 & ~n488;
  assign n2993 = ~n502 & ~n515;
  assign n2994 = ~n689 & ~n989;
  assign n2995 = n2993 & n2994;
  assign n2996 = n2991 & n2992;
  assign n2997 = n354 & n2783;
  assign n2998 = n2996 & n2997;
  assign n2999 = n1406 & n2995;
  assign n3000 = n1721 & n2527;
  assign n3001 = n2979 & n2982;
  assign n3002 = n3000 & n3001;
  assign n3003 = n2998 & n2999;
  assign n3004 = n3002 & n3003;
  assign n3005 = n2977 & n3004;
  assign n3006 = n2990 & n3005;
  assign n3007 = ~n259 & ~n308;
  assign n3008 = ~n153 & ~n253;
  assign n3009 = ~n155 & ~n278;
  assign n3010 = ~n302 & ~n601;
  assign n3011 = ~n1002 & n3010;
  assign n3012 = n813 & n3009;
  assign n3013 = n3007 & n3008;
  assign n3014 = n3012 & n3013;
  assign n3015 = n3011 & n3014;
  assign n3016 = ~n183 & ~n810;
  assign n3017 = ~n186 & ~n294;
  assign n3018 = n3016 & n3017;
  assign n3019 = ~n327 & ~n374;
  assign n3020 = ~n721 & n3019;
  assign n3021 = n1359 & n1486;
  assign n3022 = n1538 & n3021;
  assign n3023 = n3018 & n3020;
  assign n3024 = n3022 & n3023;
  assign n3025 = n2205 & n2971;
  assign n3026 = n3024 & n3025;
  assign n3027 = n2967 & n3015;
  assign n3028 = n3026 & n3027;
  assign n3029 = n671 & n3028;
  assign n3030 = n2961 & n3029;
  assign n3031 = n3006 & n3030;
  assign n3032 = ~n2951 & ~n3031;
  assign n3033 = ~n370 & ~n1699;
  assign n3034 = n487 & ~n597;
  assign n3035 = ~n314 & ~n355;
  assign n3036 = ~n409 & ~n509;
  assign n3037 = ~n511 & ~n768;
  assign n3038 = n3036 & n3037;
  assign n3039 = n1033 & n3035;
  assign n3040 = n1176 & n1453;
  assign n3041 = n2474 & n3033;
  assign n3042 = n3040 & n3041;
  assign n3043 = n3038 & n3039;
  assign n3044 = n3034 & n3043;
  assign n3045 = n3042 & n3044;
  assign n3046 = ~n427 & ~n430;
  assign n3047 = ~n503 & n3046;
  assign n3048 = ~n153 & ~n184;
  assign n3049 = ~n302 & ~n329;
  assign n3050 = ~n414 & ~n439;
  assign n3051 = n3049 & n3050;
  assign n3052 = n366 & n3048;
  assign n3053 = n3051 & n3052;
  assign n3054 = n3047 & n3053;
  assign n3055 = ~n937 & n2397;
  assign n3056 = n2001 & n3055;
  assign n3057 = ~n278 & ~n599;
  assign n3058 = ~n751 & n3057;
  assign n3059 = n767 & n3058;
  assign n3060 = ~n130 & ~n174;
  assign n3061 = ~n310 & ~n435;
  assign n3062 = ~n539 & n3061;
  assign n3063 = n530 & n3060;
  assign n3064 = n1134 & n1230;
  assign n3065 = n1971 & n3064;
  assign n3066 = n3062 & n3063;
  assign n3067 = n1728 & n2933;
  assign n3068 = n3066 & n3067;
  assign n3069 = n166 & n3065;
  assign n3070 = n652 & n3056;
  assign n3071 = n3059 & n3070;
  assign n3072 = n3068 & n3069;
  assign n3073 = n3071 & n3072;
  assign n3074 = ~n93 & ~n135;
  assign n3075 = ~n186 & ~n378;
  assign n3076 = ~n415 & n3075;
  assign n3077 = n1247 & n3074;
  assign n3078 = n3076 & n3077;
  assign n3079 = ~n253 & ~n258;
  assign n3080 = ~n276 & ~n373;
  assign n3081 = ~n689 & ~n715;
  assign n3082 = ~n792 & n3081;
  assign n3083 = n3079 & n3080;
  assign n3084 = n2500 & n3083;
  assign n3085 = n3082 & n3084;
  assign n3086 = ~n129 & ~n445;
  assign n3087 = ~n687 & n3086;
  assign n3088 = ~n183 & ~n625;
  assign n3089 = ~n718 & n3088;
  assign n3090 = ~n215 & ~n245;
  assign n3091 = ~n337 & ~n499;
  assign n3092 = n3090 & n3091;
  assign n3093 = n813 & n1457;
  assign n3094 = n1652 & n1864;
  assign n3095 = n3093 & n3094;
  assign n3096 = n3087 & n3092;
  assign n3097 = n3089 & n3096;
  assign n3098 = n3078 & n3095;
  assign n3099 = n3097 & n3098;
  assign n3100 = n3085 & n3099;
  assign n3101 = ~n304 & ~n841;
  assign n3102 = ~n116 & ~n271;
  assign n3103 = ~n273 & ~n477;
  assign n3104 = ~n564 & ~n663;
  assign n3105 = n3103 & n3104;
  assign n3106 = n749 & n3102;
  assign n3107 = n801 & n1813;
  assign n3108 = n1958 & n2208;
  assign n3109 = n2529 & n3101;
  assign n3110 = n3108 & n3109;
  assign n3111 = n3106 & n3107;
  assign n3112 = n1491 & n3105;
  assign n3113 = n3111 & n3112;
  assign n3114 = n3110 & n3113;
  assign n3115 = n3054 & n3114;
  assign n3116 = n3045 & n3115;
  assign n3117 = n3073 & n3100;
  assign n3118 = n3116 & n3117;
  assign n3119 = ~n3031 & ~n3118;
  assign n3120 = ~n282 & n500;
  assign n3121 = ~n367 & ~n503;
  assign n3122 = ~n141 & ~n379;
  assign n3123 = ~n511 & ~n599;
  assign n3124 = ~n171 & ~n355;
  assign n3125 = ~n481 & ~n535;
  assign n3126 = n3124 & n3125;
  assign n3127 = n3123 & n3126;
  assign n3128 = ~n153 & ~n563;
  assign n3129 = ~n188 & ~n508;
  assign n3130 = ~n685 & ~n1086;
  assign n3131 = ~n1404 & ~n1699;
  assign n3132 = n3130 & n3131;
  assign n3133 = n2168 & n3129;
  assign n3134 = n3128 & n3133;
  assign n3135 = n3132 & n3134;
  assign n3136 = ~n212 & ~n307;
  assign n3137 = ~n522 & ~n531;
  assign n3138 = ~n534 & n3137;
  assign n3139 = n2207 & n3136;
  assign n3140 = n3121 & n3122;
  assign n3141 = n3139 & n3140;
  assign n3142 = n991 & n3138;
  assign n3143 = n2001 & n3120;
  assign n3144 = n3142 & n3143;
  assign n3145 = n3127 & n3141;
  assign n3146 = n3144 & n3145;
  assign n3147 = n3135 & n3146;
  assign n3148 = n2398 & n3147;
  assign n3149 = ~n247 & ~n281;
  assign n3150 = ~n337 & ~n356;
  assign n3151 = ~n368 & ~n488;
  assign n3152 = ~n539 & ~n700;
  assign n3153 = ~n751 & ~n808;
  assign n3154 = n3152 & n3153;
  assign n3155 = n3150 & n3151;
  assign n3156 = n363 & n3149;
  assign n3157 = n755 & n939;
  assign n3158 = n2020 & n2253;
  assign n3159 = n3157 & n3158;
  assign n3160 = n3155 & n3156;
  assign n3161 = n3154 & n3160;
  assign n3162 = n1518 & n3159;
  assign n3163 = n3161 & n3162;
  assign n3164 = ~n162 & ~n193;
  assign n3165 = ~n256 & ~n364;
  assign n3166 = ~n515 & ~n636;
  assign n3167 = ~n638 & ~n663;
  assign n3168 = n3166 & n3167;
  assign n3169 = n3164 & n3165;
  assign n3170 = n501 & n644;
  assign n3171 = n1122 & n1296;
  assign n3172 = n1684 & n2529;
  assign n3173 = n3171 & n3172;
  assign n3174 = n3169 & n3170;
  assign n3175 = n692 & n3168;
  assign n3176 = n3174 & n3175;
  assign n3177 = n420 & n3173;
  assign n3178 = n3176 & n3177;
  assign n3179 = n2848 & n3178;
  assign n3180 = n3163 & n3179;
  assign n3181 = n2818 & n3180;
  assign n3182 = n3148 & n3181;
  assign n3183 = ~n3118 & ~n3182;
  assign n3184 = ~n130 & ~n520;
  assign n3185 = ~n627 & ~n1487;
  assign n3186 = n3184 & n3185;
  assign n3187 = ~n242 & ~n330;
  assign n3188 = ~n353 & ~n411;
  assign n3189 = ~n438 & ~n656;
  assign n3190 = n3188 & n3189;
  assign n3191 = n635 & n3187;
  assign n3192 = n704 & n1052;
  assign n3193 = n1486 & n1864;
  assign n3194 = n2126 & n2757;
  assign n3195 = n3193 & n3194;
  assign n3196 = n3191 & n3192;
  assign n3197 = n3186 & n3190;
  assign n3198 = n3196 & n3197;
  assign n3199 = n3195 & n3198;
  assign n3200 = ~n792 & n1348;
  assign n3201 = n1454 & n3200;
  assign n3202 = ~n120 & ~n445;
  assign n3203 = n1151 & n3202;
  assign n3204 = ~n568 & ~n753;
  assign n3205 = ~n284 & ~n537;
  assign n3206 = ~n168 & ~n216;
  assign n3207 = ~n319 & ~n488;
  assign n3208 = ~n532 & ~n698;
  assign n3209 = n3207 & n3208;
  assign n3210 = n1136 & n3206;
  assign n3211 = n1176 & n1356;
  assign n3212 = n1390 & n3204;
  assign n3213 = n3205 & n3212;
  assign n3214 = n3210 & n3211;
  assign n3215 = n3203 & n3209;
  assign n3216 = n3214 & n3215;
  assign n3217 = n3213 & n3216;
  assign n3218 = n1867 & n3217;
  assign n3219 = ~n151 & ~n378;
  assign n3220 = ~n248 & ~n409;
  assign n3221 = ~n839 & n3220;
  assign n3222 = n2953 & n3219;
  assign n3223 = n3221 & n3222;
  assign n3224 = ~n129 & ~n314;
  assign n3225 = ~n300 & ~n525;
  assign n3226 = ~n149 & ~n163;
  assign n3227 = ~n246 & ~n414;
  assign n3228 = ~n536 & n3227;
  assign n3229 = n372 & n3226;
  assign n3230 = n799 & n2972;
  assign n3231 = n3224 & n3225;
  assign n3232 = n3230 & n3231;
  assign n3233 = n3228 & n3229;
  assign n3234 = n3232 & n3233;
  assign n3235 = n851 & n3201;
  assign n3236 = n3223 & n3235;
  assign n3237 = n1485 & n3234;
  assign n3238 = n3236 & n3237;
  assign n3239 = n3199 & n3238;
  assign n3240 = n3147 & n3218;
  assign n3241 = n3239 & n3240;
  assign n3242 = ~n3182 & ~n3241;
  assign n3243 = ~n167 & ~n307;
  assign n3244 = ~n663 & n3243;
  assign n3245 = ~n310 & ~n721;
  assign n3246 = ~n98 & ~n148;
  assign n3247 = ~n477 & ~n703;
  assign n3248 = n3246 & n3247;
  assign n3249 = n410 & n2934;
  assign n3250 = n3245 & n3249;
  assign n3251 = n3120 & n3248;
  assign n3252 = n3244 & n3251;
  assign n3253 = n3250 & n3252;
  assign n3254 = ~n430 & ~n509;
  assign n3255 = ~n189 & ~n989;
  assign n3256 = n3254 & n3255;
  assign n3257 = ~n299 & ~n445;
  assign n3258 = ~n534 & n3257;
  assign n3259 = n612 & n725;
  assign n3260 = n3258 & n3259;
  assign n3261 = n3256 & n3260;
  assign n3262 = ~n155 & ~n596;
  assign n3263 = ~n297 & ~n1032;
  assign n3264 = n363 & n3263;
  assign n3265 = n788 & n1428;
  assign n3266 = n1651 & n1914;
  assign n3267 = n2258 & n2370;
  assign n3268 = n3262 & n3267;
  assign n3269 = n3265 & n3266;
  assign n3270 = n3264 & n3269;
  assign n3271 = n3268 & n3270;
  assign n3272 = n3261 & n3271;
  assign n3273 = n3253 & n3272;
  assign n3274 = n1750 & n2125;
  assign n3275 = n3273 & n3274;
  assign n3276 = ~n3241 & ~n3275;
  assign n3277 = ~n139 & ~n698;
  assign n3278 = ~n237 & ~n445;
  assign n3279 = ~n787 & n3278;
  assign n3280 = ~n184 & ~n839;
  assign n3281 = n3279 & n3280;
  assign n3282 = ~n106 & ~n274;
  assign n3283 = ~n297 & n3282;
  assign n3284 = n940 & n1729;
  assign n3285 = n1859 & n2501;
  assign n3286 = n2624 & n3224;
  assign n3287 = n3277 & n3286;
  assign n3288 = n3284 & n3285;
  assign n3289 = n2416 & n3283;
  assign n3290 = n3288 & n3289;
  assign n3291 = n3281 & n3287;
  assign n3292 = n3290 & n3291;
  assign n3293 = n2319 & n3292;
  assign n3294 = ~n278 & ~n382;
  assign n3295 = ~n458 & n3294;
  assign n3296 = n1292 & n2395;
  assign n3297 = n2782 & n3296;
  assign n3298 = n3295 & n3297;
  assign n3299 = ~n339 & n431;
  assign n3300 = n1049 & n3299;
  assign n3301 = ~n408 & ~n922;
  assign n3302 = ~n111 & ~n460;
  assign n3303 = ~n141 & ~n337;
  assign n3304 = ~n597 & ~n770;
  assign n3305 = n3303 & n3304;
  assign n3306 = n504 & n3301;
  assign n3307 = n3302 & n3306;
  assign n3308 = n3305 & n3307;
  assign n3309 = ~n355 & ~n639;
  assign n3310 = ~n1086 & n3309;
  assign n3311 = ~n290 & n1047;
  assign n3312 = n1403 & n3311;
  assign n3313 = ~n196 & ~n299;
  assign n3314 = ~n352 & ~n364;
  assign n3315 = ~n627 & ~n846;
  assign n3316 = n3314 & n3315;
  assign n3317 = n801 & n3313;
  assign n3318 = n1947 & n3033;
  assign n3319 = n3317 & n3318;
  assign n3320 = n3310 & n3316;
  assign n3321 = n3319 & n3320;
  assign n3322 = n3312 & n3321;
  assign n3323 = ~n168 & ~n381;
  assign n3324 = ~n751 & n3323;
  assign n3325 = ~n197 & ~n638;
  assign n3326 = ~n193 & ~n476;
  assign n3327 = ~n368 & ~n480;
  assign n3328 = ~n309 & ~n312;
  assign n3329 = ~n486 & ~n754;
  assign n3330 = n3328 & n3329;
  assign n3331 = n786 & n1122;
  assign n3332 = n1663 & n2460;
  assign n3333 = n3325 & n3326;
  assign n3334 = n3327 & n3333;
  assign n3335 = n3331 & n3332;
  assign n3336 = n2596 & n3330;
  assign n3337 = n3324 & n3336;
  assign n3338 = n3334 & n3335;
  assign n3339 = n3337 & n3338;
  assign n3340 = n3308 & n3339;
  assign n3341 = n3322 & n3340;
  assign n3342 = ~n259 & ~n383;
  assign n3343 = ~n512 & n3342;
  assign n3344 = ~n186 & ~n307;
  assign n3345 = ~n281 & ~n534;
  assign n3346 = n1700 & n3345;
  assign n3347 = ~n416 & n3101;
  assign n3348 = n3344 & n3347;
  assign n3349 = n3343 & n3348;
  assign n3350 = n3346 & n3349;
  assign n3351 = ~n245 & ~n329;
  assign n3352 = n2359 & n3351;
  assign n3353 = ~n135 & ~n148;
  assign n3354 = ~n159 & ~n269;
  assign n3355 = ~n427 & ~n477;
  assign n3356 = ~n646 & ~n656;
  assign n3357 = ~n893 & n3356;
  assign n3358 = n3354 & n3355;
  assign n3359 = n272 & n3353;
  assign n3360 = n799 & n1133;
  assign n3361 = n1913 & n3360;
  assign n3362 = n3358 & n3359;
  assign n3363 = n3352 & n3357;
  assign n3364 = n3362 & n3363;
  assign n3365 = n3300 & n3361;
  assign n3366 = n3364 & n3365;
  assign n3367 = n3298 & n3366;
  assign n3368 = n3350 & n3367;
  assign n3369 = n3293 & n3368;
  assign n3370 = n3341 & n3369;
  assign n3371 = ~n3275 & ~n3370;
  assign n3372 = n3275 & n3370;
  assign n3373 = ~n3371 & ~n3372;
  assign n3374 = ~n604 & ~n1404;
  assign n3375 = ~n148 & ~n537;
  assign n3376 = ~n894 & ~n937;
  assign n3377 = ~n944 & n3376;
  assign n3378 = n3374 & n3375;
  assign n3379 = n3377 & n3378;
  assign n3380 = ~n358 & ~n508;
  assign n3381 = ~n605 & n3380;
  assign n3382 = n917 & n3381;
  assign n3383 = n1621 & n3382;
  assign n3384 = ~n243 & ~n639;
  assign n3385 = n479 & n3384;
  assign n3386 = ~n126 & ~n239;
  assign n3387 = n260 & n3386;
  assign n3388 = n298 & n785;
  assign n3389 = n1429 & n1652;
  assign n3390 = n2783 & n3389;
  assign n3391 = n3387 & n3388;
  assign n3392 = n1152 & n3385;
  assign n3393 = n3391 & n3392;
  assign n3394 = n3379 & n3390;
  assign n3395 = n3393 & n3394;
  assign n3396 = n3383 & n3395;
  assign n3397 = ~n269 & ~n715;
  assign n3398 = n657 & n3397;
  assign n3399 = ~n168 & ~n313;
  assign n3400 = ~n656 & n2905;
  assign n3401 = n172 & n3399;
  assign n3402 = n1685 & n1971;
  assign n3403 = n2460 & n2792;
  assign n3404 = n3402 & n3403;
  assign n3405 = n3400 & n3401;
  assign n3406 = n3404 & n3405;
  assign n3407 = ~n163 & ~n685;
  assign n3408 = ~n116 & ~n383;
  assign n3409 = ~n271 & ~n561;
  assign n3410 = ~n123 & ~n531;
  assign n3411 = ~n653 & ~n687;
  assign n3412 = n3410 & n3411;
  assign n3413 = n357 & n1003;
  assign n3414 = n1198 & n1357;
  assign n3415 = n1812 & n2561;
  assign n3416 = n2624 & n3016;
  assign n3417 = n3407 & n3408;
  assign n3418 = n3409 & n3417;
  assign n3419 = n3415 & n3416;
  assign n3420 = n3413 & n3414;
  assign n3421 = n3398 & n3412;
  assign n3422 = n3420 & n3421;
  assign n3423 = n3418 & n3419;
  assign n3424 = n3422 & n3423;
  assign n3425 = n3406 & n3424;
  assign n3426 = n475 & n3425;
  assign n3427 = n3396 & n3426;
  assign n3428 = n3370 & n3427;
  assign n3429 = ~n211 & ~n374;
  assign n3430 = ~n476 & ~n1086;
  assign n3431 = n3429 & n3430;
  assign n3432 = ~n188 & ~n700;
  assign n3433 = ~n98 & ~n482;
  assign n3434 = ~n724 & n3433;
  assign n3435 = n2608 & n3434;
  assign n3436 = ~n256 & ~n438;
  assign n3437 = ~n989 & ~n1002;
  assign n3438 = n3436 & n3437;
  assign n3439 = n2710 & n3438;
  assign n3440 = ~n130 & ~n355;
  assign n3441 = ~n422 & n3440;
  assign n3442 = n1508 & n3441;
  assign n3443 = n2077 & n3442;
  assign n3444 = ~n136 & ~n310;
  assign n3445 = ~n352 & n3444;
  assign n3446 = ~n216 & ~n270;
  assign n3447 = ~n381 & n3446;
  assign n3448 = n939 & n1012;
  assign n3449 = n1422 & n1913;
  assign n3450 = n2838 & n3325;
  assign n3451 = n3449 & n3450;
  assign n3452 = n3447 & n3448;
  assign n3453 = n2262 & n3445;
  assign n3454 = n3452 & n3453;
  assign n3455 = n3451 & n3454;
  assign n3456 = n3085 & n3443;
  assign n3457 = n3455 & n3456;
  assign n3458 = ~n116 & ~n120;
  assign n3459 = ~n183 & ~n439;
  assign n3460 = ~n525 & ~n597;
  assign n3461 = ~n235 & ~n252;
  assign n3462 = ~n368 & ~n377;
  assign n3463 = ~n539 & ~n894;
  assign n3464 = n3462 & n3463;
  assign n3465 = n372 & n3461;
  assign n3466 = n2474 & n3458;
  assign n3467 = n3459 & n3460;
  assign n3468 = n3466 & n3467;
  assign n3469 = n3464 & n3465;
  assign n3470 = n3468 & n3469;
  assign n3471 = ~n721 & n758;
  assign n3472 = ~n242 & ~n703;
  assign n3473 = n749 & n3472;
  assign n3474 = n901 & n1350;
  assign n3475 = n2108 & n3432;
  assign n3476 = n3474 & n3475;
  assign n3477 = n3431 & n3473;
  assign n3478 = n3471 & n3477;
  assign n3479 = n3056 & n3476;
  assign n3480 = n3435 & n3439;
  assign n3481 = n3479 & n3480;
  assign n3482 = n3470 & n3478;
  assign n3483 = n3481 & n3482;
  assign n3484 = n3293 & n3483;
  assign n3485 = n3457 & n3484;
  assign n3486 = ~n3428 & ~n3485;
  assign n3487 = n3373 & n3486;
  assign n3488 = ~n3371 & ~n3487;
  assign n3489 = n3241 & n3275;
  assign n3490 = ~n3276 & ~n3489;
  assign n3491 = ~n3488 & n3490;
  assign n3492 = ~n3276 & ~n3491;
  assign n3493 = n3182 & n3241;
  assign n3494 = ~n3242 & ~n3493;
  assign n3495 = ~n3492 & n3494;
  assign n3496 = ~n3242 & ~n3495;
  assign n3497 = n3118 & n3182;
  assign n3498 = ~n3183 & ~n3497;
  assign n3499 = ~n3496 & n3498;
  assign n3500 = ~n3183 & ~n3499;
  assign n3501 = n3031 & n3118;
  assign n3502 = ~n3119 & ~n3501;
  assign n3503 = ~n3500 & n3502;
  assign n3504 = ~n3119 & ~n3503;
  assign n3505 = n2951 & n3031;
  assign n3506 = ~n3032 & ~n3505;
  assign n3507 = ~n3504 & n3506;
  assign n3508 = ~n3032 & ~n3507;
  assign n3509 = n2919 & n2951;
  assign n3510 = ~n2952 & ~n3509;
  assign n3511 = ~n3508 & n3510;
  assign n3512 = ~n2952 & ~n3511;
  assign n3513 = n2835 & n2919;
  assign n3514 = ~n2920 & ~n3513;
  assign n3515 = ~n3512 & n3514;
  assign n3516 = ~n2920 & ~n3515;
  assign n3517 = n2778 & n2835;
  assign n3518 = ~n2836 & ~n3517;
  assign n3519 = ~n3516 & n3518;
  assign n3520 = ~n2836 & ~n3519;
  assign n3521 = n2708 & n2778;
  assign n3522 = ~n2779 & ~n3521;
  assign n3523 = ~n3520 & n3522;
  assign n3524 = ~n2779 & ~n3523;
  assign n3525 = n2674 & n2708;
  assign n3526 = ~n2709 & ~n3525;
  assign n3527 = ~n3524 & n3526;
  assign n3528 = ~n2709 & ~n3527;
  assign n3529 = n2589 & n2674;
  assign n3530 = ~n2675 & ~n3529;
  assign n3531 = ~n3528 & n3530;
  assign n3532 = ~n2675 & ~n3531;
  assign n3533 = n2496 & n2589;
  assign n3534 = ~n2590 & ~n3533;
  assign n3535 = ~n3532 & n3534;
  assign n3536 = ~n2590 & ~n3535;
  assign n3537 = n2412 & n2496;
  assign n3538 = ~n2497 & ~n3537;
  assign n3539 = ~n3536 & n3538;
  assign n3540 = ~n2497 & ~n3539;
  assign n3541 = n2347 & n2412;
  assign n3542 = ~n2413 & ~n3541;
  assign n3543 = ~n3540 & n3542;
  assign n3544 = ~n2413 & ~n3543;
  assign n3545 = n2249 & n2347;
  assign n3546 = ~n2348 & ~n3545;
  assign n3547 = ~n3544 & n3546;
  assign n3548 = ~n2348 & ~n3547;
  assign n3549 = n2146 & n2249;
  assign n3550 = ~n2250 & ~n3549;
  assign n3551 = ~n3548 & n3550;
  assign n3552 = ~n2250 & ~n3551;
  assign n3553 = n2098 & n2146;
  assign n3554 = ~n2147 & ~n3553;
  assign n3555 = ~n3552 & n3554;
  assign n3556 = ~n2147 & ~n3555;
  assign n3557 = n1998 & n2098;
  assign n3558 = ~n2099 & ~n3557;
  assign n3559 = ~n3556 & n3558;
  assign n3560 = ~n2099 & ~n3559;
  assign n3561 = n1908 & n1998;
  assign n3562 = ~n1999 & ~n3561;
  assign n3563 = ~n3560 & n3562;
  assign n3564 = ~n1999 & ~n3563;
  assign n3565 = n1841 & n1908;
  assign n3566 = ~n1909 & ~n3565;
  assign n3567 = ~n3564 & n3566;
  assign n3568 = ~n1909 & ~n3567;
  assign n3569 = n1717 & n1841;
  assign n3570 = ~n1842 & ~n3569;
  assign n3571 = ~n3568 & n3570;
  assign n3572 = ~n1842 & ~n3571;
  assign n3573 = n1637 & n1717;
  assign n3574 = ~n1718 & ~n3573;
  assign n3575 = ~n3572 & n3574;
  assign n3576 = ~n1718 & ~n3575;
  assign n3577 = n1533 & n1637;
  assign n3578 = ~n1638 & ~n3577;
  assign n3579 = ~n3576 & n3578;
  assign n3580 = ~n1638 & ~n3579;
  assign n3581 = n1448 & n1533;
  assign n3582 = ~n1534 & ~n3581;
  assign n3583 = ~n3580 & n3582;
  assign n3584 = ~n1534 & ~n3583;
  assign n3585 = n1345 & n1448;
  assign n3586 = ~n1449 & ~n3585;
  assign n3587 = ~n3584 & n3586;
  assign n3588 = ~n1449 & ~n3587;
  assign n3589 = n1225 & n1345;
  assign n3590 = ~n1346 & ~n3589;
  assign n3591 = ~n3588 & n3590;
  assign n3592 = ~n1346 & ~n3591;
  assign n3593 = n1104 & n1225;
  assign n3594 = ~n1226 & ~n3593;
  assign n3595 = ~n3592 & n3594;
  assign n3596 = ~n1226 & ~n3595;
  assign n3597 = n878 & n1104;
  assign n3598 = ~n1105 & ~n3597;
  assign n3599 = ~n3596 & n3598;
  assign n3600 = ~n1105 & ~n3599;
  assign n3601 = n878 & n987;
  assign n3602 = ~n988 & ~n3601;
  assign n3603 = ~n3600 & n3602;
  assign n3604 = ~n988 & ~n3603;
  assign n3605 = ~n126 & ~n367;
  assign n3606 = n272 & n3605;
  assign n3607 = n1508 & n3606;
  assign n3608 = n2967 & n3607;
  assign n3609 = ~n534 & n900;
  assign n3610 = n1133 & n1296;
  assign n3611 = n2126 & n3610;
  assign n3612 = n3609 & n3611;
  assign n3613 = n766 & n3612;
  assign n3614 = n3608 & n3613;
  assign n3615 = ~n167 & ~n243;
  assign n3616 = ~n249 & ~n314;
  assign n3617 = ~n810 & n3616;
  assign n3618 = n3615 & n3617;
  assign n3619 = ~n145 & ~n308;
  assign n3620 = ~n106 & ~n171;
  assign n3621 = ~n284 & ~n416;
  assign n3622 = ~n703 & n3621;
  assign n3623 = n3619 & n3620;
  assign n3624 = n3622 & n3623;
  assign n3625 = n3203 & n3624;
  assign n3626 = n275 & ~n310;
  assign n3627 = n598 & n3254;
  assign n3628 = n3626 & n3627;
  assign n3629 = n2369 & n3628;
  assign n3630 = ~n1404 & n3629;
  assign n3631 = ~n247 & ~n276;
  assign n3632 = n1380 & n3631;
  assign n3633 = ~n328 & ~n1032;
  assign n3634 = n444 & n3633;
  assign n3635 = n1428 & n2206;
  assign n3636 = n2838 & n3635;
  assign n3637 = n3634 & n3636;
  assign n3638 = n3439 & n3637;
  assign n3639 = ~n409 & ~n604;
  assign n3640 = n645 & n3639;
  assign n3641 = n1009 & n1351;
  assign n3642 = n1639 & n3641;
  assign n3643 = n3640 & n3642;
  assign n3644 = ~n318 & ~n488;
  assign n3645 = ~n153 & ~n529;
  assign n3646 = n3644 & n3645;
  assign n3647 = ~n216 & ~n499;
  assign n3648 = n2234 & n3647;
  assign n3649 = n3646 & n3648;
  assign n3650 = ~n532 & ~n685;
  assign n3651 = n752 & n3650;
  assign n3652 = n847 & n3651;
  assign n3653 = n3649 & n3652;
  assign n3654 = n3643 & n3653;
  assign n3655 = ~n724 & n782;
  assign n3656 = n1198 & n3655;
  assign n3657 = n3632 & n3656;
  assign n3658 = n1013 & n3657;
  assign n3659 = n3638 & n3658;
  assign n3660 = n3654 & n3659;
  assign n3661 = ~n111 & n1650;
  assign n3662 = ~n334 & ~n564;
  assign n3663 = ~n427 & ~n808;
  assign n3664 = ~n197 & ~n894;
  assign n3665 = ~n194 & ~n353;
  assign n3666 = n992 & n3665;
  assign n3667 = n3662 & n3663;
  assign n3668 = n3664 & n3667;
  assign n3669 = n3661 & n3666;
  assign n3670 = n3668 & n3669;
  assign n3671 = n904 & n3670;
  assign n3672 = n932 & n3671;
  assign n3673 = n891 & n3672;
  assign n3674 = ~n291 & n3630;
  assign n3675 = n3660 & n3674;
  assign n3676 = n3673 & n3675;
  assign n3677 = n600 & ~n1699;
  assign n3678 = n3618 & n3677;
  assign n3679 = n3625 & n3678;
  assign n3680 = n3614 & n3679;
  assign n3681 = n3676 & n3680;
  assign n3682 = ~n987 & ~n3681;
  assign n3683 = n987 & n3681;
  assign n3684 = ~n3682 & ~n3683;
  assign n3685 = ~n3604 & n3684;
  assign n3686 = n3604 & ~n3684;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = n880 & n3687;
  assign n3689 = pi30  & ~pi31 ;
  assign n3690 = ~pi30  & pi31 ;
  assign n3691 = ~n3689 & ~n3690;
  assign n3692 = n746 & ~n3691;
  assign n3693 = ~n987 & n3692;
  assign n3694 = ~pi31  & ~n746;
  assign n3695 = ~n3681 & n3694;
  assign n3696 = ~n879 & ~n3693;
  assign n3697 = ~n3695 & n3696;
  assign n3698 = ~n3688 & n3697;
  assign n3699 = n745 & ~n3698;
  assign n3700 = ~n745 & n3698;
  assign n3701 = ~n3699 & ~n3700;
  assign n3702 = ~n149 & ~n592;
  assign n3703 = ~n443 & ~n445;
  assign n3704 = ~n846 & n3703;
  assign n3705 = ~n151 & ~n477;
  assign n3706 = ~n259 & ~n296;
  assign n3707 = ~n537 & n3706;
  assign n3708 = ~n170 & ~n189;
  assign n3709 = ~n282 & ~n299;
  assign n3710 = ~n416 & n3709;
  assign n3711 = n272 & n3708;
  assign n3712 = n786 & n3705;
  assign n3713 = n3711 & n3712;
  assign n3714 = n3707 & n3710;
  assign n3715 = n3713 & n3714;
  assign n3716 = n1662 & n3715;
  assign n3717 = ~n195 & ~n250;
  assign n3718 = ~n284 & ~n625;
  assign n3719 = n3662 & n3718;
  assign n3720 = n3717 & n3719;
  assign n3721 = ~n183 & ~n328;
  assign n3722 = ~n529 & n3721;
  assign n3723 = ~n368 & ~n656;
  assign n3724 = ~n190 & ~n211;
  assign n3725 = ~n281 & n3724;
  assign n3726 = ~n380 & ~n510;
  assign n3727 = ~n256 & ~n297;
  assign n3728 = ~n332 & n3727;
  assign n3729 = n3723 & n3726;
  assign n3730 = n3728 & n3729;
  assign n3731 = n3725 & n3730;
  assign n3732 = ~n136 & ~n212;
  assign n3733 = ~n902 & n3732;
  assign n3734 = ~n174 & ~n422;
  assign n3735 = ~n486 & ~n839;
  assign n3736 = n3734 & n3735;
  assign n3737 = n719 & n1049;
  assign n3738 = n2207 & n2397;
  assign n3739 = n2934 & n3738;
  assign n3740 = n3736 & n3737;
  assign n3741 = n1624 & n3733;
  assign n3742 = n3740 & n3741;
  assign n3743 = n3739 & n3742;
  assign n3744 = ~n175 & ~n248;
  assign n3745 = ~n365 & ~n536;
  assign n3746 = ~n563 & ~n604;
  assign n3747 = ~n814 & n3746;
  assign n3748 = n655 & n3745;
  assign n3749 = n1151 & n3245;
  assign n3750 = n3744 & n3749;
  assign n3751 = n3747 & n3748;
  assign n3752 = n3722 & n3751;
  assign n3753 = n133 & n3750;
  assign n3754 = n3720 & n3753;
  assign n3755 = n3731 & n3752;
  assign n3756 = n3754 & n3755;
  assign n3757 = n3743 & n3756;
  assign n3758 = ~n200 & ~n361;
  assign n3759 = ~n531 & ~n768;
  assign n3760 = n3758 & n3759;
  assign n3761 = n527 & n938;
  assign n3762 = n1133 & n1243;
  assign n3763 = n2529 & n3702;
  assign n3764 = n3762 & n3763;
  assign n3765 = n3760 & n3761;
  assign n3766 = n3704 & n3765;
  assign n3767 = n3764 & n3766;
  assign n3768 = n3716 & n3767;
  assign n3769 = n3757 & n3768;
  assign n3770 = n407 & ~n3769;
  assign n3771 = ~n407 & n3769;
  assign n3772 = ~n3770 & ~n3771;
  assign n3773 = ~n1104 & n3692;
  assign n3774 = n3596 & ~n3598;
  assign n3775 = ~n3599 & ~n3774;
  assign n3776 = n880 & n3775;
  assign n3777 = n748 & ~n1225;
  assign n3778 = ~n878 & n3694;
  assign n3779 = ~n3773 & ~n3777;
  assign n3780 = ~n3778 & n3779;
  assign n3781 = ~n3776 & n3780;
  assign n3782 = n3772 & ~n3781;
  assign n3783 = ~n3770 & ~n3782;
  assign n3784 = ~pi26  & ~n590;
  assign n3785 = ~n588 & n591;
  assign n3786 = ~n3784 & ~n3785;
  assign n3787 = ~n3783 & ~n3786;
  assign n3788 = n3783 & n3786;
  assign n3789 = ~n987 & n3694;
  assign n3790 = n3600 & ~n3602;
  assign n3791 = ~n3603 & ~n3790;
  assign n3792 = n880 & n3791;
  assign n3793 = n748 & ~n1104;
  assign n3794 = ~n878 & n3692;
  assign n3795 = ~n3789 & ~n3793;
  assign n3796 = ~n3794 & n3795;
  assign n3797 = ~n3792 & n3796;
  assign n3798 = ~n3788 & ~n3797;
  assign n3799 = ~n3787 & ~n3798;
  assign n3800 = n3701 & ~n3799;
  assign n3801 = ~n3701 & n3799;
  assign n3802 = pi28  & ~pi29 ;
  assign n3803 = ~pi28  & pi29 ;
  assign n3804 = ~n3802 & ~n3803;
  assign n3805 = pi26  & ~pi27 ;
  assign n3806 = ~pi26  & pi27 ;
  assign n3807 = ~n3805 & ~n3806;
  assign n3808 = ~n107 & ~n112;
  assign n3809 = n3807 & ~n3808;
  assign n3810 = ~n3804 & n3809;
  assign n3811 = ~n414 & ~n639;
  assign n3812 = ~n838 & n3811;
  assign n3813 = n3702 & n3812;
  assign n3814 = n1085 & n3813;
  assign n3815 = ~n291 & ~n685;
  assign n3816 = n1136 & n3815;
  assign n3817 = n1424 & n1684;
  assign n3818 = n3619 & n3817;
  assign n3819 = n1535 & n3816;
  assign n3820 = n3818 & n3819;
  assign n3821 = n3814 & n3820;
  assign n3822 = n600 & n647;
  assign n3823 = ~n171 & ~n269;
  assign n3824 = ~n337 & ~n378;
  assign n3825 = ~n445 & ~n603;
  assign n3826 = n3824 & n3825;
  assign n3827 = n176 & n3823;
  assign n3828 = n1767 & n3827;
  assign n3829 = n3822 & n3826;
  assign n3830 = n3828 & n3829;
  assign n3831 = ~n317 & ~n841;
  assign n3832 = n3830 & n3831;
  assign n3833 = n3608 & n3832;
  assign n3834 = n2961 & n3833;
  assign n3835 = ~n477 & ~n814;
  assign n3836 = n137 & n3835;
  assign n3837 = ~n296 & ~n518;
  assign n3838 = ~n531 & ~n601;
  assign n3839 = ~n1034 & n3838;
  assign n3840 = n375 & n722;
  assign n3841 = n725 & n1913;
  assign n3842 = n3837 & n3841;
  assign n3843 = n3839 & n3840;
  assign n3844 = n1349 & n3843;
  assign n3845 = n3842 & n3844;
  assign n3846 = ~n180 & ~n235;
  assign n3847 = n3836 & n3846;
  assign n3848 = n3845 & n3847;
  assign n3849 = n719 & n896;
  assign n3850 = n1170 & n3849;
  assign n3851 = n3848 & n3850;
  assign n3852 = n3834 & n3851;
  assign n3853 = ~n304 & ~n634;
  assign n3854 = n3821 & n3853;
  assign n3855 = n3852 & n3854;
  assign n3856 = n3810 & ~n3855;
  assign n3857 = ~n634 & n3618;
  assign n3858 = ~n922 & ~n1699;
  assign n3859 = ~n98 & ~n190;
  assign n3860 = ~n338 & ~n377;
  assign n3861 = ~n661 & ~n663;
  assign n3862 = n3860 & n3861;
  assign n3863 = n759 & n3859;
  assign n3864 = n1296 & n2610;
  assign n3865 = n2934 & n3864;
  assign n3866 = n3862 & n3863;
  assign n3867 = n3865 & n3866;
  assign n3868 = ~n248 & ~n255;
  assign n3869 = ~n259 & ~n481;
  assign n3870 = ~n508 & n3869;
  assign n3871 = n2797 & n3868;
  assign n3872 = n3870 & n3871;
  assign n3873 = n487 & ~n653;
  assign n3874 = n755 & n797;
  assign n3875 = n900 & n1509;
  assign n3876 = n3858 & n3875;
  assign n3877 = n3873 & n3874;
  assign n3878 = n3876 & n3877;
  assign n3879 = n3872 & n3878;
  assign n3880 = n3867 & n3879;
  assign n3881 = ~n183 & n3880;
  assign n3882 = n3857 & n3881;
  assign n3883 = n3821 & n3882;
  assign n3884 = n3807 & n3808;
  assign n3885 = ~n3883 & n3884;
  assign n3886 = ~n3804 & ~n3807;
  assign n3887 = ~n3681 & ~n3855;
  assign n3888 = ~n3682 & ~n3685;
  assign n3889 = n3681 & n3855;
  assign n3890 = ~n3887 & ~n3889;
  assign n3891 = ~n3888 & n3890;
  assign n3892 = ~n3887 & ~n3891;
  assign n3893 = ~n3855 & ~n3883;
  assign n3894 = n3855 & n3882;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = ~n3892 & n3895;
  assign n3897 = n3855 & ~n3896;
  assign n3898 = ~n3883 & n3897;
  assign n3899 = n3883 & n3896;
  assign n3900 = ~n3898 & ~n3899;
  assign n3901 = n3886 & ~n3900;
  assign n3902 = ~n3856 & ~n3885;
  assign n3903 = ~n3901 & n3902;
  assign n3904 = pi29  & n3903;
  assign n3905 = ~pi29  & ~n3903;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = ~n3801 & ~n3906;
  assign n3908 = ~n3800 & ~n3907;
  assign n3909 = ~n482 & ~n510;
  assign n3910 = ~n532 & n3909;
  assign n3911 = ~n252 & ~n355;
  assign n3912 = ~n163 & ~n175;
  assign n3913 = ~n195 & ~n529;
  assign n3914 = n3912 & n3913;
  assign n3915 = n633 & n1351;
  assign n3916 = n2323 & n3911;
  assign n3917 = n3915 & n3916;
  assign n3918 = n3910 & n3914;
  assign n3919 = n3917 & n3918;
  assign n3920 = ~n653 & ~n689;
  assign n3921 = ~n238 & ~n300;
  assign n3922 = ~n411 & ~n663;
  assign n3923 = ~n810 & ~n1034;
  assign n3924 = n3922 & n3923;
  assign n3925 = n447 & n3921;
  assign n3926 = n791 & n1268;
  assign n3927 = n1643 & n3926;
  assign n3928 = n3924 & n3925;
  assign n3929 = n1170 & n3928;
  assign n3930 = n3927 & n3929;
  assign n3931 = ~n129 & ~n319;
  assign n3932 = ~n362 & n3931;
  assign n3933 = n3930 & n3932;
  assign n3934 = ~n145 & ~n534;
  assign n3935 = ~n329 & ~n1404;
  assign n3936 = n3934 & n3935;
  assign n3937 = ~n111 & ~n168;
  assign n3938 = ~n358 & ~n531;
  assign n3939 = ~n808 & ~n944;
  assign n3940 = n3938 & n3939;
  assign n3941 = n410 & n3937;
  assign n3942 = n528 & n933;
  assign n3943 = n1356 & n2208;
  assign n3944 = n3920 & n3943;
  assign n3945 = n3941 & n3942;
  assign n3946 = n2039 & n3940;
  assign n3947 = n3279 & n3936;
  assign n3948 = n3946 & n3947;
  assign n3949 = n3944 & n3945;
  assign n3950 = n2506 & n3949;
  assign n3951 = n1778 & n3948;
  assign n3952 = n3919 & n3951;
  assign n3953 = n3950 & n3952;
  assign n3954 = n2125 & n3933;
  assign n3955 = n3953 & n3954;
  assign n3956 = ~n742 & n3955;
  assign n3957 = n742 & ~n3955;
  assign n3958 = ~n3956 & ~n3957;
  assign n3959 = ~n744 & ~n3698;
  assign n3960 = ~n743 & ~n3959;
  assign n3961 = n3958 & ~n3960;
  assign n3962 = ~n3958 & n3960;
  assign n3963 = ~n3961 & ~n3962;
  assign n3964 = n3886 & ~n3897;
  assign n3965 = ~n3810 & ~n3964;
  assign n3966 = ~n3883 & ~n3965;
  assign n3967 = ~pi29  & n3966;
  assign n3968 = pi29  & ~n3966;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = n3694 & ~n3855;
  assign n3971 = n3888 & ~n3890;
  assign n3972 = ~n3891 & ~n3971;
  assign n3973 = n880 & n3972;
  assign n3974 = n748 & ~n987;
  assign n3975 = ~n3681 & n3692;
  assign n3976 = ~n3970 & ~n3974;
  assign n3977 = ~n3975 & n3976;
  assign n3978 = ~n3973 & n3977;
  assign n3979 = ~n3969 & ~n3978;
  assign n3980 = n3969 & n3978;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = n3963 & ~n3981;
  assign n3983 = ~n3963 & n3981;
  assign n3984 = ~n3982 & ~n3983;
  assign n3985 = ~n3908 & ~n3984;
  assign n3986 = ~n3772 & n3781;
  assign n3987 = ~n3782 & ~n3986;
  assign n3988 = ~n258 & ~n435;
  assign n3989 = ~n193 & ~n276;
  assign n3990 = ~n355 & ~n445;
  assign n3991 = ~n656 & n3990;
  assign n3992 = n900 & n3989;
  assign n3993 = n3988 & n3992;
  assign n3994 = n3991 & n3993;
  assign n3995 = ~n242 & ~n329;
  assign n3996 = n2253 & n3995;
  assign n3997 = ~n601 & ~n841;
  assign n3998 = ~n215 & ~n248;
  assign n3999 = ~n597 & n3998;
  assign n4000 = n562 & n1151;
  assign n4001 = n3997 & n4000;
  assign n4002 = n3999 & n4001;
  assign n4003 = ~n238 & ~n459;
  assign n4004 = ~n300 & ~n661;
  assign n4005 = ~n180 & ~n186;
  assign n4006 = ~n412 & ~n446;
  assign n4007 = ~n1487 & n4006;
  assign n4008 = n1113 & n4005;
  assign n4009 = n1387 & n4003;
  assign n4010 = n4004 & n4009;
  assign n4011 = n4007 & n4008;
  assign n4012 = n1239 & n2278;
  assign n4013 = n4011 & n4012;
  assign n4014 = n4010 & n4013;
  assign n4015 = ~n281 & ~n358;
  assign n4016 = ~n143 & ~n178;
  assign n4017 = ~n250 & ~n639;
  assign n4018 = n4016 & n4017;
  assign n4019 = n198 & n1248;
  assign n4020 = n4015 & n4019;
  assign n4021 = n4018 & n4020;
  assign n4022 = n164 & ~n703;
  assign n4023 = ~n249 & ~n255;
  assign n4024 = ~n636 & ~n698;
  assign n4025 = ~n838 & n4024;
  assign n4026 = n1453 & n4023;
  assign n4027 = n2597 & n4026;
  assign n4028 = n4022 & n4025;
  assign n4029 = n4027 & n4028;
  assign n4030 = n3298 & n4029;
  assign n4031 = n4002 & n4021;
  assign n4032 = n4030 & n4031;
  assign n4033 = n4014 & n4032;
  assign n4034 = ~n98 & ~n356;
  assign n4035 = ~n136 & ~n476;
  assign n4036 = ~n502 & n4035;
  assign n4037 = n4034 & n4036;
  assign n4038 = ~n111 & ~n334;
  assign n4039 = ~n361 & ~n368;
  assign n4040 = ~n381 & ~n839;
  assign n4041 = n4039 & n4040;
  assign n4042 = n154 & n4038;
  assign n4043 = n528 & n2757;
  assign n4044 = n4042 & n4043;
  assign n4045 = n3120 & n4041;
  assign n4046 = n3996 & n4045;
  assign n4047 = n4037 & n4044;
  assign n4048 = n4046 & n4047;
  assign n4049 = n2156 & n3994;
  assign n4050 = n4048 & n4049;
  assign n4051 = n4033 & n4050;
  assign n4052 = n593 & n809;
  assign n4053 = n3016 & n4052;
  assign n4054 = ~n120 & ~n358;
  assign n4055 = ~n481 & n4054;
  assign n4056 = n1423 & n4055;
  assign n4057 = ~n330 & ~n371;
  assign n4058 = ~n446 & n4057;
  assign n4059 = n786 & n3301;
  assign n4060 = n4058 & n4059;
  assign n4061 = n4053 & n4060;
  assign n4062 = n4056 & n4061;
  assign n4063 = ~n249 & ~n309;
  assign n4064 = ~n136 & ~n211;
  assign n4065 = ~n380 & ~n422;
  assign n4066 = n4064 & n4065;
  assign n4067 = ~n212 & ~n597;
  assign n4068 = ~n724 & n4067;
  assign n4069 = ~n130 & ~n155;
  assign n4070 = ~n838 & n4069;
  assign n4071 = n257 & n436;
  assign n4072 = n657 & n913;
  assign n4073 = n941 & n1047;
  assign n4074 = n1751 & n4073;
  assign n4075 = n4071 & n4072;
  assign n4076 = n336 & n4070;
  assign n4077 = n4066 & n4068;
  assign n4078 = n4076 & n4077;
  assign n4079 = n4074 & n4075;
  assign n4080 = n1191 & n4079;
  assign n4081 = n4078 & n4080;
  assign n4082 = ~n303 & ~n383;
  assign n4083 = n1357 & n4082;
  assign n4084 = n2044 & n3645;
  assign n4085 = n4083 & n4084;
  assign n4086 = ~n111 & ~n170;
  assign n4087 = ~n284 & ~n374;
  assign n4088 = ~n754 & n4087;
  assign n4089 = n413 & n4086;
  assign n4090 = n540 & n635;
  assign n4091 = n1515 & n1729;
  assign n4092 = n1752 & n2783;
  assign n4093 = n4091 & n4092;
  assign n4094 = n4089 & n4090;
  assign n4095 = n4088 & n4094;
  assign n4096 = n491 & n4093;
  assign n4097 = n1361 & n4085;
  assign n4098 = n4096 & n4097;
  assign n4099 = n2355 & n4095;
  assign n4100 = n4098 & n4099;
  assign n4101 = n4081 & n4100;
  assign n4102 = ~n563 & ~n599;
  assign n4103 = ~n353 & ~n1034;
  assign n4104 = n654 & n4103;
  assign n4105 = n2200 & n3911;
  assign n4106 = n4102 & n4105;
  assign n4107 = n4104 & n4106;
  assign n4108 = ~n180 & ~n415;
  assign n4109 = ~n503 & ~n646;
  assign n4110 = n4108 & n4109;
  assign n4111 = ~n148 & ~n178;
  assign n4112 = ~n186 & ~n238;
  assign n4113 = ~n367 & ~n510;
  assign n4114 = ~n814 & n4113;
  assign n4115 = n4111 & n4112;
  assign n4116 = n1456 & n1570;
  assign n4117 = n4063 & n4116;
  assign n4118 = n4114 & n4115;
  assign n4119 = n1773 & n4110;
  assign n4120 = n4118 & n4119;
  assign n4121 = n2084 & n4117;
  assign n4122 = n4120 & n4121;
  assign n4123 = n4107 & n4122;
  assign n4124 = n4062 & n4123;
  assign n4125 = n4101 & n4124;
  assign n4126 = ~n4051 & ~n4125;
  assign n4127 = n4051 & n4125;
  assign n4128 = ~pi23  & ~n4126;
  assign n4129 = ~n4127 & n4128;
  assign n4130 = ~n4126 & ~n4129;
  assign n4131 = ~n407 & n4130;
  assign n4132 = n407 & ~n4130;
  assign n4133 = ~n1225 & n3692;
  assign n4134 = n3592 & ~n3594;
  assign n4135 = ~n3595 & ~n4134;
  assign n4136 = n880 & n4135;
  assign n4137 = n748 & ~n1345;
  assign n4138 = ~n1104 & n3694;
  assign n4139 = ~n4133 & ~n4137;
  assign n4140 = ~n4138 & n4139;
  assign n4141 = ~n4136 & n4140;
  assign n4142 = ~n4132 & n4141;
  assign n4143 = ~n4131 & ~n4142;
  assign n4144 = n3987 & n4143;
  assign n4145 = ~n3987 & ~n4143;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = ~pi23  & ~n4129;
  assign n4148 = ~n4127 & n4130;
  assign n4149 = ~n4147 & ~n4148;
  assign n4150 = n748 & ~n1448;
  assign n4151 = n3588 & ~n3590;
  assign n4152 = ~n3591 & ~n4151;
  assign n4153 = n880 & n4152;
  assign n4154 = ~n1345 & n3692;
  assign n4155 = ~n1225 & n3694;
  assign n4156 = ~n4150 & ~n4154;
  assign n4157 = ~n4155 & n4156;
  assign n4158 = ~n4153 & n4157;
  assign n4159 = ~n4149 & ~n4158;
  assign n4160 = ~n139 & ~n370;
  assign n4161 = ~n437 & n4160;
  assign n4162 = n940 & n4161;
  assign n4163 = ~n194 & ~n339;
  assign n4164 = ~n135 & ~n178;
  assign n4165 = ~n200 & ~n252;
  assign n4166 = ~n515 & n4165;
  assign n4167 = ~n186 & ~n276;
  assign n4168 = ~n126 & n640;
  assign n4169 = n3920 & n4167;
  assign n4170 = n4168 & n4169;
  assign n4171 = n426 & n4170;
  assign n4172 = ~n197 & ~n246;
  assign n4173 = ~n625 & n4172;
  assign n4174 = n533 & n750;
  assign n4175 = n784 & n935;
  assign n4176 = n1357 & n2658;
  assign n4177 = n4163 & n4164;
  assign n4178 = n4176 & n4177;
  assign n4179 = n4174 & n4175;
  assign n4180 = n4166 & n4173;
  assign n4181 = n4179 & n4180;
  assign n4182 = n4178 & n4181;
  assign n4183 = n4171 & n4182;
  assign n4184 = ~n502 & ~n535;
  assign n4185 = ~n596 & n4184;
  assign n4186 = ~n170 & ~n242;
  assign n4187 = ~n297 & ~n520;
  assign n4188 = n4186 & n4187;
  assign n4189 = n2158 & n4188;
  assign n4190 = n4185 & n4189;
  assign n4191 = ~n215 & ~n303;
  assign n4192 = ~n511 & ~n594;
  assign n4193 = ~n1086 & n4192;
  assign n4194 = n421 & n4191;
  assign n4195 = n431 & n440;
  assign n4196 = n1471 & n2279;
  assign n4197 = n4195 & n4196;
  assign n4198 = n4193 & n4194;
  assign n4199 = n4197 & n4198;
  assign n4200 = n1572 & n4162;
  assign n4201 = n4199 & n4200;
  assign n4202 = n4190 & n4201;
  assign n4203 = n1857 & n4202;
  assign n4204 = n3073 & n4183;
  assign n4205 = n4203 & n4204;
  assign n4206 = n4051 & ~n4205;
  assign n4207 = ~n4051 & n4205;
  assign n4208 = ~n4206 & ~n4207;
  assign n4209 = ~n276 & n3034;
  assign n4210 = ~n355 & ~n564;
  assign n4211 = ~n661 & n4210;
  assign n4212 = n664 & n1348;
  assign n4213 = n4211 & n4212;
  assign n4214 = ~n200 & ~n307;
  assign n4215 = ~n313 & n4214;
  assign n4216 = n528 & n1003;
  assign n4217 = n1011 & n2206;
  assign n4218 = n2658 & n4217;
  assign n4219 = n4215 & n4216;
  assign n4220 = n720 & n2159;
  assign n4221 = n3431 & n4220;
  assign n4222 = n4218 & n4219;
  assign n4223 = n4209 & n4213;
  assign n4224 = n4222 & n4223;
  assign n4225 = n4221 & n4224;
  assign n4226 = ~n184 & ~n304;
  assign n4227 = ~n308 & ~n437;
  assign n4228 = ~n488 & n4227;
  assign n4229 = n154 & n4226;
  assign n4230 = n1242 & n2921;
  assign n4231 = n4229 & n4230;
  assign n4232 = n630 & n4228;
  assign n4233 = n4231 & n4232;
  assign n4234 = ~n162 & ~n167;
  assign n4235 = ~n310 & ~n368;
  assign n4236 = ~n723 & ~n787;
  assign n4237 = n4235 & n4236;
  assign n4238 = n272 & n4234;
  assign n4239 = n279 & n901;
  assign n4240 = n1563 & n2625;
  assign n4241 = n4239 & n4240;
  assign n4242 = n4237 & n4238;
  assign n4243 = n4185 & n4242;
  assign n4244 = n4241 & n4243;
  assign n4245 = n2694 & n4233;
  assign n4246 = n4244 & n4245;
  assign n4247 = ~n193 & ~n510;
  assign n4248 = ~n529 & ~n563;
  assign n4249 = n4247 & n4248;
  assign n4250 = n150 & n298;
  assign n4251 = n936 & n1230;
  assign n4252 = n1476 & n1539;
  assign n4253 = n1669 & n1863;
  assign n4254 = n2783 & n4253;
  assign n4255 = n4251 & n4252;
  assign n4256 = n4249 & n4250;
  assign n4257 = n3661 & n4256;
  assign n4258 = n4254 & n4255;
  assign n4259 = n4257 & n4258;
  assign n4260 = n2082 & n4259;
  assign n4261 = n2367 & n4260;
  assign n4262 = n4225 & n4246;
  assign n4263 = n4261 & n4262;
  assign n4264 = ~n178 & ~n247;
  assign n4265 = ~n242 & ~n416;
  assign n4266 = n840 & n4265;
  assign n4267 = ~n136 & ~n768;
  assign n4268 = n4063 & n4267;
  assign n4269 = ~n271 & ~n382;
  assign n4270 = ~n145 & ~n151;
  assign n4271 = ~n604 & n4270;
  assign n4272 = n1883 & n3408;
  assign n4273 = n4271 & n4272;
  assign n4274 = ~n277 & ~n721;
  assign n4275 = n440 & n4274;
  assign n4276 = n940 & n1004;
  assign n4277 = n1476 & n1684;
  assign n4278 = n2007 & n2040;
  assign n4279 = n3033 & n4264;
  assign n4280 = n4269 & n4279;
  assign n4281 = n4277 & n4278;
  assign n4282 = n4275 & n4276;
  assign n4283 = n4266 & n4268;
  assign n4284 = n4282 & n4283;
  assign n4285 = n4280 & n4281;
  assign n4286 = n4273 & n4285;
  assign n4287 = n4284 & n4286;
  assign n4288 = ~n129 & ~n135;
  assign n4289 = ~n171 & ~n245;
  assign n4290 = ~n274 & ~n293;
  assign n4291 = ~n376 & ~n414;
  assign n4292 = ~n522 & ~n596;
  assign n4293 = ~n636 & ~n989;
  assign n4294 = ~n1404 & n4293;
  assign n4295 = n4291 & n4292;
  assign n4296 = n4289 & n4290;
  assign n4297 = n3837 & n4288;
  assign n4298 = n4296 & n4297;
  assign n4299 = n4294 & n4295;
  assign n4300 = n4298 & n4299;
  assign n4301 = ~n170 & ~n294;
  assign n4302 = ~n902 & n4301;
  assign n4303 = ~n106 & ~n235;
  assign n4304 = ~n299 & ~n303;
  assign n4305 = ~n353 & ~n371;
  assign n4306 = ~n412 & n4305;
  assign n4307 = n4303 & n4304;
  assign n4308 = n789 & n959;
  assign n4309 = n1136 & n1538;
  assign n4310 = n4308 & n4309;
  assign n4311 = n4306 & n4307;
  assign n4312 = n4310 & n4311;
  assign n4313 = n434 & ~n894;
  assign n4314 = ~n291 & ~n503;
  assign n4315 = ~n509 & ~n627;
  assign n4316 = n4314 & n4315;
  assign n4317 = n530 & n1354;
  assign n4318 = n1779 & n2208;
  assign n4319 = n4317 & n4318;
  assign n4320 = n4302 & n4316;
  assign n4321 = n4313 & n4320;
  assign n4322 = n4319 & n4321;
  assign n4323 = n2394 & n4312;
  assign n4324 = n4322 & n4323;
  assign n4325 = ~n255 & ~n798;
  assign n4326 = ~n422 & ~n443;
  assign n4327 = ~n167 & ~n283;
  assign n4328 = n1088 & n4327;
  assign n4329 = n1508 & n3205;
  assign n4330 = n4325 & n4326;
  assign n4331 = n4329 & n4330;
  assign n4332 = n4328 & n4331;
  assign n4333 = ~n184 & ~n319;
  assign n4334 = ~n482 & ~n515;
  assign n4335 = n4333 & n4334;
  assign n4336 = n369 & n704;
  assign n4337 = n1186 & n1248;
  assign n4338 = n4336 & n4337;
  assign n4339 = n3089 & n4335;
  assign n4340 = n4338 & n4339;
  assign n4341 = n1080 & n4340;
  assign n4342 = n4300 & n4332;
  assign n4343 = n4341 & n4342;
  assign n4344 = n4287 & n4343;
  assign n4345 = n4324 & n4344;
  assign n4346 = ~n4263 & ~n4345;
  assign n4347 = n4263 & n4345;
  assign n4348 = ~pi20  & ~n4346;
  assign n4349 = ~n4347 & n4348;
  assign n4350 = ~n4346 & ~n4349;
  assign n4351 = ~n4205 & n4350;
  assign n4352 = n4205 & ~n4350;
  assign n4353 = ~n1533 & n3692;
  assign n4354 = n3580 & ~n3582;
  assign n4355 = ~n3583 & ~n4354;
  assign n4356 = n880 & n4355;
  assign n4357 = n748 & ~n1637;
  assign n4358 = ~n1448 & n3694;
  assign n4359 = ~n4353 & ~n4357;
  assign n4360 = ~n4358 & n4359;
  assign n4361 = ~n4356 & n4360;
  assign n4362 = ~n4352 & n4361;
  assign n4363 = ~n4351 & ~n4362;
  assign n4364 = n4208 & n4363;
  assign n4365 = ~n4206 & ~n4364;
  assign n4366 = n4149 & n4158;
  assign n4367 = ~n4159 & ~n4366;
  assign n4368 = ~n4365 & n4367;
  assign n4369 = ~n4159 & ~n4368;
  assign n4370 = ~n4131 & ~n4132;
  assign n4371 = ~n4141 & n4370;
  assign n4372 = n4141 & ~n4370;
  assign n4373 = ~n4371 & ~n4372;
  assign n4374 = ~n4369 & n4373;
  assign n4375 = n4369 & ~n4373;
  assign n4376 = ~n4374 & ~n4375;
  assign n4377 = ~n878 & n3810;
  assign n4378 = n3687 & n3886;
  assign n4379 = ~n987 & n3884;
  assign n4380 = n3804 & ~n3807;
  assign n4381 = ~n3681 & n4380;
  assign n4382 = ~n4377 & ~n4379;
  assign n4383 = ~n4381 & n4382;
  assign n4384 = ~n4378 & n4383;
  assign n4385 = pi29  & n4384;
  assign n4386 = ~pi29  & ~n4384;
  assign n4387 = ~n4385 & ~n4386;
  assign n4388 = n4376 & ~n4387;
  assign n4389 = ~n4374 & ~n4388;
  assign n4390 = n4146 & ~n4389;
  assign n4391 = ~n4144 & ~n4390;
  assign n4392 = ~n3787 & ~n3788;
  assign n4393 = ~n3797 & n4392;
  assign n4394 = n3797 & ~n4392;
  assign n4395 = ~n4393 & ~n4394;
  assign n4396 = ~n4391 & n4395;
  assign n4397 = ~n3883 & n4380;
  assign n4398 = n3892 & ~n3895;
  assign n4399 = ~n3896 & ~n4398;
  assign n4400 = n3886 & n4399;
  assign n4401 = ~n3855 & n3884;
  assign n4402 = ~n3681 & n3810;
  assign n4403 = ~n4397 & ~n4401;
  assign n4404 = ~n4402 & n4403;
  assign n4405 = ~n4400 & n4404;
  assign n4406 = pi29  & n4405;
  assign n4407 = ~pi29  & ~n4405;
  assign n4408 = ~n4406 & ~n4407;
  assign n4409 = n4391 & ~n4395;
  assign n4410 = ~n4396 & ~n4409;
  assign n4411 = ~n4408 & n4410;
  assign n4412 = ~n4396 & ~n4411;
  assign n4413 = ~n3800 & ~n3801;
  assign n4414 = ~n3906 & n4413;
  assign n4415 = n3906 & ~n4413;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = ~n4412 & n4416;
  assign n4418 = n4412 & ~n4416;
  assign n4419 = ~n4417 & ~n4418;
  assign n4420 = ~n78 & ~n81;
  assign n4421 = ~n3897 & n4420;
  assign n4422 = ~n86 & ~n4421;
  assign n4423 = ~n3883 & ~n4422;
  assign n4424 = ~pi26  & n4423;
  assign n4425 = pi26  & ~n4423;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = ~n3855 & n4380;
  assign n4428 = n3886 & n3972;
  assign n4429 = ~n987 & n3810;
  assign n4430 = ~n3681 & n3884;
  assign n4431 = ~n4427 & ~n4429;
  assign n4432 = ~n4430 & n4431;
  assign n4433 = ~n4428 & n4432;
  assign n4434 = pi29  & n4433;
  assign n4435 = ~pi29  & ~n4433;
  assign n4436 = ~n4434 & ~n4435;
  assign n4437 = ~n4426 & ~n4436;
  assign n4438 = ~n4146 & n4389;
  assign n4439 = ~n4390 & ~n4438;
  assign n4440 = n4426 & n4436;
  assign n4441 = ~n4437 & ~n4440;
  assign n4442 = n4439 & n4441;
  assign n4443 = ~n4437 & ~n4442;
  assign n4444 = n4408 & ~n4410;
  assign n4445 = ~n4411 & ~n4444;
  assign n4446 = ~n4443 & n4445;
  assign n4447 = ~n4376 & n4387;
  assign n4448 = ~n4388 & ~n4447;
  assign n4449 = ~n4208 & ~n4363;
  assign n4450 = ~n4364 & ~n4449;
  assign n4451 = n748 & ~n1533;
  assign n4452 = n3584 & ~n3586;
  assign n4453 = ~n3587 & ~n4452;
  assign n4454 = n880 & n4453;
  assign n4455 = ~n1448 & n3692;
  assign n4456 = ~n1345 & n3694;
  assign n4457 = ~n4451 & ~n4455;
  assign n4458 = ~n4456 & n4457;
  assign n4459 = ~n4454 & n4458;
  assign n4460 = n4450 & ~n4459;
  assign n4461 = ~n4351 & ~n4352;
  assign n4462 = ~n4361 & n4461;
  assign n4463 = n4361 & ~n4461;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = ~n236 & ~n414;
  assign n4466 = ~n178 & ~n253;
  assign n4467 = ~n302 & ~n408;
  assign n4468 = ~n535 & n4467;
  assign n4469 = n3460 & n4466;
  assign n4470 = n4465 & n4469;
  assign n4471 = n4468 & n4470;
  assign n4472 = ~n189 & ~n721;
  assign n4473 = n2252 & n4472;
  assign n4474 = ~n162 & ~n296;
  assign n4475 = ~n373 & n4474;
  assign n4476 = n1535 & n4475;
  assign n4477 = ~n299 & n448;
  assign n4478 = n2040 & n4477;
  assign n4479 = ~n135 & ~n180;
  assign n4480 = ~n246 & ~n502;
  assign n4481 = n4479 & n4480;
  assign n4482 = n1035 & n1516;
  assign n4483 = n1754 & n1962;
  assign n4484 = n4482 & n4483;
  assign n4485 = n1008 & n4481;
  assign n4486 = n1393 & n4485;
  assign n4487 = n4473 & n4484;
  assign n4488 = n4476 & n4478;
  assign n4489 = n4487 & n4488;
  assign n4490 = n4471 & n4486;
  assign n4491 = n4489 & n4490;
  assign n4492 = ~n149 & ~n297;
  assign n4493 = ~n846 & n4492;
  assign n4494 = n1575 & n1779;
  assign n4495 = ~n273 & ~n282;
  assign n4496 = ~n308 & ~n422;
  assign n4497 = ~n503 & ~n792;
  assign n4498 = n4496 & n4497;
  assign n4499 = n799 & n4495;
  assign n4500 = n4498 & n4499;
  assign n4501 = ~n339 & ~n443;
  assign n4502 = ~n168 & ~n235;
  assign n4503 = ~n370 & ~n382;
  assign n4504 = ~n601 & n4503;
  assign n4505 = n1826 & n4502;
  assign n4506 = n4501 & n4505;
  assign n4507 = n4504 & n4506;
  assign n4508 = ~n239 & ~n284;
  assign n4509 = ~n477 & n4508;
  assign n4510 = n146 & n434;
  assign n4511 = n938 & n1508;
  assign n4512 = n4510 & n4511;
  assign n4513 = n610 & n4509;
  assign n4514 = n1267 & n4494;
  assign n4515 = n4513 & n4514;
  assign n4516 = n4500 & n4512;
  assign n4517 = n4515 & n4516;
  assign n4518 = n4507 & n4517;
  assign n4519 = ~n256 & ~n319;
  assign n4520 = ~n409 & n4519;
  assign n4521 = n440 & n1243;
  assign n4522 = n2044 & n4004;
  assign n4523 = n4521 & n4522;
  assign n4524 = n854 & n4520;
  assign n4525 = n4493 & n4524;
  assign n4526 = n2713 & n4523;
  assign n4527 = n4525 & n4526;
  assign n4528 = n1545 & n2977;
  assign n4529 = n4527 & n4528;
  assign n4530 = n4491 & n4529;
  assign n4531 = n4518 & n4530;
  assign n4532 = n4263 & ~n4531;
  assign n4533 = ~n4263 & n4531;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = ~n1717 & n3692;
  assign n4536 = n3572 & ~n3574;
  assign n4537 = ~n3575 & ~n4536;
  assign n4538 = n880 & n4537;
  assign n4539 = n748 & ~n1841;
  assign n4540 = ~n1637 & n3694;
  assign n4541 = ~n4535 & ~n4539;
  assign n4542 = ~n4540 & n4541;
  assign n4543 = ~n4538 & n4542;
  assign n4544 = n4534 & ~n4543;
  assign n4545 = ~n4532 & ~n4544;
  assign n4546 = ~pi20  & ~n4349;
  assign n4547 = ~n4347 & n4350;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = ~n4545 & ~n4548;
  assign n4550 = n4545 & n4548;
  assign n4551 = ~n1637 & n3692;
  assign n4552 = n3576 & ~n3578;
  assign n4553 = ~n3579 & ~n4552;
  assign n4554 = n880 & n4553;
  assign n4555 = n748 & ~n1717;
  assign n4556 = ~n1533 & n3694;
  assign n4557 = ~n4551 & ~n4555;
  assign n4558 = ~n4556 & n4557;
  assign n4559 = ~n4554 & n4558;
  assign n4560 = ~n4550 & ~n4559;
  assign n4561 = ~n4549 & ~n4560;
  assign n4562 = n4464 & ~n4561;
  assign n4563 = ~n4464 & n4561;
  assign n4564 = ~n4562 & ~n4563;
  assign n4565 = ~n1225 & n3884;
  assign n4566 = n3886 & n4135;
  assign n4567 = ~n1345 & n3810;
  assign n4568 = ~n1104 & n4380;
  assign n4569 = ~n4565 & ~n4567;
  assign n4570 = ~n4568 & n4569;
  assign n4571 = ~n4566 & n4570;
  assign n4572 = pi29  & n4571;
  assign n4573 = ~pi29  & ~n4571;
  assign n4574 = ~n4572 & ~n4573;
  assign n4575 = n4564 & ~n4574;
  assign n4576 = ~n4562 & ~n4575;
  assign n4577 = n4450 & n4459;
  assign n4578 = ~n4450 & ~n4459;
  assign n4579 = ~n4577 & ~n4578;
  assign n4580 = ~n4576 & ~n4579;
  assign n4581 = ~n4460 & ~n4580;
  assign n4582 = n4365 & ~n4367;
  assign n4583 = ~n4368 & ~n4582;
  assign n4584 = n4581 & ~n4583;
  assign n4585 = ~n4581 & n4583;
  assign n4586 = ~n987 & n4380;
  assign n4587 = n3791 & n3886;
  assign n4588 = ~n1104 & n3810;
  assign n4589 = ~n878 & n3884;
  assign n4590 = ~n4586 & ~n4588;
  assign n4591 = ~n4589 & n4590;
  assign n4592 = ~n4587 & n4591;
  assign n4593 = pi29  & n4592;
  assign n4594 = ~pi29  & ~n4592;
  assign n4595 = ~n4593 & ~n4594;
  assign n4596 = ~n4585 & n4595;
  assign n4597 = ~n4584 & ~n4596;
  assign n4598 = n4448 & n4597;
  assign n4599 = n86 & ~n3855;
  assign n4600 = n81 & n84;
  assign n4601 = ~n3883 & n4600;
  assign n4602 = ~n3900 & n4420;
  assign n4603 = ~n4599 & ~n4601;
  assign n4604 = ~n4602 & n4603;
  assign n4605 = ~pi26  & ~n4604;
  assign n4606 = pi26  & n4604;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = ~n4448 & ~n4597;
  assign n4609 = ~n4598 & ~n4608;
  assign n4610 = ~n4607 & n4609;
  assign n4611 = ~n4598 & ~n4610;
  assign n4612 = ~n4439 & ~n4441;
  assign n4613 = ~n4442 & ~n4612;
  assign n4614 = ~n4611 & n4613;
  assign n4615 = n78 & ~n81;
  assign n4616 = ~n3883 & n4615;
  assign n4617 = n4399 & n4420;
  assign n4618 = ~n3855 & n4600;
  assign n4619 = n86 & ~n3681;
  assign n4620 = ~n4616 & ~n4618;
  assign n4621 = ~n4619 & n4620;
  assign n4622 = ~n4617 & n4621;
  assign n4623 = pi26  & n4622;
  assign n4624 = ~pi26  & ~n4622;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = ~n1104 & n3884;
  assign n4627 = n3775 & n3886;
  assign n4628 = ~n1225 & n3810;
  assign n4629 = ~n878 & n4380;
  assign n4630 = ~n4626 & ~n4628;
  assign n4631 = ~n4629 & n4630;
  assign n4632 = ~n4627 & n4631;
  assign n4633 = pi29  & n4632;
  assign n4634 = ~pi29  & ~n4632;
  assign n4635 = ~n4633 & ~n4634;
  assign n4636 = n4576 & n4579;
  assign n4637 = ~n4580 & ~n4636;
  assign n4638 = n4635 & ~n4637;
  assign n4639 = ~n4635 & n4637;
  assign n4640 = ~n3855 & n4615;
  assign n4641 = n3972 & n4420;
  assign n4642 = n86 & ~n987;
  assign n4643 = ~n3681 & n4600;
  assign n4644 = ~n4640 & ~n4642;
  assign n4645 = ~n4643 & n4644;
  assign n4646 = ~n4641 & n4645;
  assign n4647 = pi26  & n4646;
  assign n4648 = ~pi26  & ~n4646;
  assign n4649 = ~n4647 & ~n4648;
  assign n4650 = ~n4639 & n4649;
  assign n4651 = ~n4638 & ~n4650;
  assign n4652 = ~n4625 & n4651;
  assign n4653 = n4625 & n4651;
  assign n4654 = ~n4625 & ~n4651;
  assign n4655 = ~n4653 & ~n4654;
  assign n4656 = ~n4584 & ~n4585;
  assign n4657 = ~n4595 & ~n4656;
  assign n4658 = n4595 & n4656;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = ~n4655 & ~n4659;
  assign n4661 = ~n4652 & ~n4660;
  assign n4662 = n4607 & ~n4609;
  assign n4663 = ~n4610 & ~n4662;
  assign n4664 = ~n4661 & n4663;
  assign n4665 = n4655 & n4659;
  assign n4666 = ~n4660 & ~n4665;
  assign n4667 = ~n1345 & n3884;
  assign n4668 = n3886 & n4152;
  assign n4669 = ~n1448 & n3810;
  assign n4670 = ~n1225 & n4380;
  assign n4671 = ~n4667 & ~n4669;
  assign n4672 = ~n4670 & n4671;
  assign n4673 = ~n4668 & n4672;
  assign n4674 = ~pi29  & ~n4673;
  assign n4675 = pi29  & n4673;
  assign n4676 = ~n4674 & ~n4675;
  assign n4677 = ~n4549 & ~n4550;
  assign n4678 = ~n4559 & n4677;
  assign n4679 = n4559 & ~n4677;
  assign n4680 = ~n4678 & ~n4679;
  assign n4681 = ~n4676 & n4680;
  assign n4682 = ~n4676 & ~n4680;
  assign n4683 = n4676 & n4680;
  assign n4684 = ~n4682 & ~n4683;
  assign n4685 = ~n4534 & n4543;
  assign n4686 = ~n4544 & ~n4685;
  assign n4687 = ~n409 & ~n526;
  assign n4688 = ~n787 & ~n894;
  assign n4689 = n2983 & n4688;
  assign n4690 = ~n174 & ~n509;
  assign n4691 = ~n592 & ~n689;
  assign n4692 = n4690 & n4691;
  assign n4693 = n434 & n660;
  assign n4694 = n1229 & n1347;
  assign n4695 = n1450 & n1884;
  assign n4696 = n2108 & n4687;
  assign n4697 = n4695 & n4696;
  assign n4698 = n4693 & n4694;
  assign n4699 = n4689 & n4692;
  assign n4700 = n4698 & n4699;
  assign n4701 = n1386 & n4697;
  assign n4702 = n4700 & n4701;
  assign n4703 = n3015 & n4702;
  assign n4704 = n957 & n3199;
  assign n4705 = n4703 & n4704;
  assign n4706 = n1045 & n4705;
  assign n4707 = ~n258 & ~n604;
  assign n4708 = n1014 & n4707;
  assign n4709 = ~n317 & ~n526;
  assign n4710 = ~n190 & ~n282;
  assign n4711 = ~n362 & ~n893;
  assign n4712 = n4710 & n4711;
  assign n4713 = n2042 & n4709;
  assign n4714 = n4712 & n4713;
  assign n4715 = ~n139 & ~n307;
  assign n4716 = n2007 & n4715;
  assign n4717 = n2658 & n4716;
  assign n4718 = ~n174 & ~n376;
  assign n4719 = ~n409 & ~n808;
  assign n4720 = n4718 & n4719;
  assign n4721 = n784 & n1006;
  assign n4722 = n1018 & n1730;
  assign n4723 = n2528 & n4501;
  assign n4724 = n4722 & n4723;
  assign n4725 = n4720 & n4721;
  assign n4726 = n1050 & n4708;
  assign n4727 = n4725 & n4726;
  assign n4728 = n2199 & n4724;
  assign n4729 = n4714 & n4717;
  assign n4730 = n4728 & n4729;
  assign n4731 = n4727 & n4730;
  assign n4732 = ~n377 & ~n1699;
  assign n4733 = n567 & n4732;
  assign n4734 = ~n116 & ~n135;
  assign n4735 = ~n309 & ~n355;
  assign n4736 = n4734 & n4735;
  assign n4737 = ~n213 & ~n237;
  assign n4738 = ~n297 & ~n373;
  assign n4739 = n4737 & n4738;
  assign n4740 = n124 & n602;
  assign n4741 = n1424 & n1754;
  assign n4742 = n2251 & n2445;
  assign n4743 = n3101 & n4742;
  assign n4744 = n4740 & n4741;
  assign n4745 = n1455 & n4739;
  assign n4746 = n4733 & n4736;
  assign n4747 = n4745 & n4746;
  assign n4748 = n4743 & n4744;
  assign n4749 = n1013 & n4748;
  assign n4750 = n4747 & n4749;
  assign n4751 = n4731 & n4750;
  assign n4752 = n1328 & n4751;
  assign n4753 = ~n4706 & ~n4752;
  assign n4754 = n4706 & n4752;
  assign n4755 = ~pi17  & ~n4753;
  assign n4756 = ~n4754 & n4755;
  assign n4757 = ~n4753 & ~n4756;
  assign n4758 = n4263 & ~n4757;
  assign n4759 = ~n4263 & n4757;
  assign n4760 = ~n1841 & n3692;
  assign n4761 = n3568 & ~n3570;
  assign n4762 = ~n3571 & ~n4761;
  assign n4763 = n880 & n4762;
  assign n4764 = n748 & ~n1908;
  assign n4765 = ~n1717 & n3694;
  assign n4766 = ~n4760 & ~n4764;
  assign n4767 = ~n4765 & n4766;
  assign n4768 = ~n4763 & n4767;
  assign n4769 = ~n4759 & ~n4768;
  assign n4770 = ~n4758 & ~n4769;
  assign n4771 = n4686 & ~n4770;
  assign n4772 = ~n4686 & n4770;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = ~pi17  & ~n4756;
  assign n4775 = ~n4754 & n4757;
  assign n4776 = ~n4774 & ~n4775;
  assign n4777 = n748 & ~n1998;
  assign n4778 = n3564 & ~n3566;
  assign n4779 = ~n3567 & ~n4778;
  assign n4780 = n880 & n4779;
  assign n4781 = ~n1908 & n3692;
  assign n4782 = ~n1841 & n3694;
  assign n4783 = ~n4777 & ~n4781;
  assign n4784 = ~n4782 & n4783;
  assign n4785 = ~n4780 & n4784;
  assign n4786 = ~n4776 & ~n4785;
  assign n4787 = ~n270 & ~n810;
  assign n4788 = n3204 & n4787;
  assign n4789 = ~n98 & ~n188;
  assign n4790 = ~n215 & ~n249;
  assign n4791 = ~n256 & ~n291;
  assign n4792 = ~n352 & ~n808;
  assign n4793 = n4791 & n4792;
  assign n4794 = n4789 & n4790;
  assign n4795 = n447 & n500;
  assign n4796 = n1755 & n3702;
  assign n4797 = n4795 & n4796;
  assign n4798 = n4793 & n4794;
  assign n4799 = n4788 & n4798;
  assign n4800 = n2800 & n4797;
  assign n4801 = n4799 & n4800;
  assign n4802 = ~n116 & ~n213;
  assign n4803 = ~n212 & n504;
  assign n4804 = n1176 & n1783;
  assign n4805 = n1947 & n4804;
  assign n4806 = n4803 & n4805;
  assign n4807 = n3201 & n4806;
  assign n4808 = ~n211 & ~n259;
  assign n4809 = ~n278 & ~n411;
  assign n4810 = ~n526 & ~n594;
  assign n4811 = n4809 & n4810;
  assign n4812 = n3164 & n4808;
  assign n4813 = n372 & n2658;
  assign n4814 = n2978 & n4802;
  assign n4815 = n4813 & n4814;
  assign n4816 = n4811 & n4812;
  assign n4817 = n3279 & n4816;
  assign n4818 = n1537 & n4815;
  assign n4819 = n3078 & n4818;
  assign n4820 = n3443 & n4817;
  assign n4821 = n4819 & n4820;
  assign n4822 = n4801 & n4807;
  assign n4823 = n4821 & n4822;
  assign n4824 = n684 & n4823;
  assign n4825 = n4706 & ~n4824;
  assign n4826 = ~n4706 & n4824;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = ~n93 & ~n1487;
  assign n4829 = ~n636 & n4828;
  assign n4830 = ~n291 & ~n902;
  assign n4831 = n2169 & n4830;
  assign n4832 = ~n143 & ~n189;
  assign n4833 = ~n339 & ~n476;
  assign n4834 = ~n512 & ~n646;
  assign n4835 = ~n808 & n4834;
  assign n4836 = n4832 & n4833;
  assign n4837 = n436 & n4836;
  assign n4838 = n632 & n4835;
  assign n4839 = n1985 & n4829;
  assign n4840 = n4831 & n4839;
  assign n4841 = n4837 & n4838;
  assign n4842 = n1277 & n3281;
  assign n4843 = n4841 & n4842;
  assign n4844 = n4840 & n4843;
  assign n4845 = ~n437 & n892;
  assign n4846 = ~n145 & ~n213;
  assign n4847 = ~n216 & ~n249;
  assign n4848 = ~n330 & ~n409;
  assign n4849 = ~n539 & ~n703;
  assign n4850 = n4848 & n4849;
  assign n4851 = n4846 & n4847;
  assign n4852 = n1307 & n2460;
  assign n4853 = n4465 & n4852;
  assign n4854 = n4850 & n4851;
  assign n4855 = n4845 & n4854;
  assign n4856 = n4853 & n4855;
  assign n4857 = ~n256 & ~n273;
  assign n4858 = ~n499 & ~n648;
  assign n4859 = ~n156 & ~n314;
  assign n4860 = ~n596 & ~n604;
  assign n4861 = n4859 & n4860;
  assign n4862 = n1450 & n4858;
  assign n4863 = n4861 & n4862;
  assign n4864 = ~n282 & ~n566;
  assign n4865 = ~n529 & ~n754;
  assign n4866 = n1671 & n4865;
  assign n4867 = n1939 & n4866;
  assign n4868 = ~n123 & ~n274;
  assign n4869 = ~n537 & n4868;
  assign n4870 = n298 & n1003;
  assign n4871 = n1377 & n1754;
  assign n4872 = n4864 & n4871;
  assign n4873 = n4869 & n4870;
  assign n4874 = n2722 & n3445;
  assign n4875 = n4873 & n4874;
  assign n4876 = n4863 & n4872;
  assign n4877 = n4867 & n4876;
  assign n4878 = n4875 & n4877;
  assign n4879 = n4807 & n4878;
  assign n4880 = ~n180 & ~n605;
  assign n4881 = ~n653 & n4880;
  assign n4882 = ~n178 & ~n281;
  assign n4883 = ~n378 & n4882;
  assign n4884 = n657 & n3101;
  assign n4885 = n4883 & n4884;
  assign n4886 = n4881 & n4885;
  assign n4887 = ~n269 & ~n753;
  assign n4888 = ~n197 & ~n253;
  assign n4889 = ~n770 & n4888;
  assign n4890 = ~n135 & ~n317;
  assign n4891 = ~n368 & ~n944;
  assign n4892 = n4890 & n4891;
  assign n4893 = n447 & n1006;
  assign n4894 = n1012 & n4857;
  assign n4895 = n4887 & n4894;
  assign n4896 = n4892 & n4893;
  assign n4897 = n2933 & n4889;
  assign n4898 = n4896 & n4897;
  assign n4899 = n4209 & n4895;
  assign n4900 = n4898 & n4899;
  assign n4901 = n4886 & n4900;
  assign n4902 = n4856 & n4901;
  assign n4903 = n4844 & n4902;
  assign n4904 = n4879 & n4903;
  assign n4905 = ~n625 & ~n636;
  assign n4906 = n117 & n647;
  assign n4907 = ~n183 & ~n281;
  assign n4908 = ~n294 & ~n409;
  assign n4909 = ~n535 & ~n1032;
  assign n4910 = n4908 & n4909;
  assign n4911 = n137 & n4907;
  assign n4912 = n933 & n1242;
  assign n4913 = n1813 & n2619;
  assign n4914 = n4905 & n4913;
  assign n4915 = n4911 & n4912;
  assign n4916 = n4906 & n4910;
  assign n4917 = n4915 & n4916;
  assign n4918 = n3059 & n4914;
  assign n4919 = n4500 & n4918;
  assign n4920 = n4917 & n4919;
  assign n4921 = ~n283 & ~n370;
  assign n4922 = ~n1034 & n4921;
  assign n4923 = n1670 & n4922;
  assign n4924 = n2533 & n4923;
  assign n4925 = ~n238 & ~n303;
  assign n4926 = ~n486 & ~n510;
  assign n4927 = ~n536 & ~n685;
  assign n4928 = n602 & n4927;
  assign n4929 = n1846 & n4925;
  assign n4930 = n4926 & n4929;
  assign n4931 = n2006 & n4928;
  assign n4932 = n3087 & n4931;
  assign n4933 = n4930 & n4932;
  assign n4934 = ~n245 & ~n893;
  assign n4935 = ~n194 & ~n381;
  assign n4936 = ~n846 & n4935;
  assign n4937 = n505 & n1175;
  assign n4938 = n1883 & n3008;
  assign n4939 = n3409 & n4938;
  assign n4940 = n4936 & n4937;
  assign n4941 = n4733 & n4940;
  assign n4942 = n4939 & n4941;
  assign n4943 = ~n123 & ~n237;
  assign n4944 = ~n482 & ~n563;
  assign n4945 = ~n594 & ~n634;
  assign n4946 = n4944 & n4945;
  assign n4947 = n150 & n4943;
  assign n4948 = n654 & n2201;
  assign n4949 = n4934 & n4948;
  assign n4950 = n4946 & n4947;
  assign n4951 = n4788 & n4950;
  assign n4952 = n4949 & n4951;
  assign n4953 = n1001 & n4952;
  assign n4954 = n4942 & n4953;
  assign n4955 = n1752 & n2192;
  assign n4956 = ~n246 & ~n297;
  assign n4957 = ~n359 & n4956;
  assign n4958 = n533 & n901;
  assign n4959 = n1112 & n2610;
  assign n4960 = n2797 & n4959;
  assign n4961 = n4957 & n4958;
  assign n4962 = n1046 & n1912;
  assign n4963 = n4955 & n4962;
  assign n4964 = n4960 & n4961;
  assign n4965 = n4963 & n4964;
  assign n4966 = n4924 & n4965;
  assign n4967 = n4933 & n4966;
  assign n4968 = n4920 & n4967;
  assign n4969 = n4954 & n4968;
  assign n4970 = ~n4904 & ~n4969;
  assign n4971 = n4904 & n4969;
  assign n4972 = ~pi14  & ~n4970;
  assign n4973 = ~n4971 & n4972;
  assign n4974 = ~n4970 & ~n4973;
  assign n4975 = n4824 & ~n4974;
  assign n4976 = ~n4824 & n4974;
  assign n4977 = ~n2098 & n3692;
  assign n4978 = n3556 & ~n3558;
  assign n4979 = ~n3559 & ~n4978;
  assign n4980 = n880 & n4979;
  assign n4981 = n748 & ~n2146;
  assign n4982 = ~n1998 & n3694;
  assign n4983 = ~n4977 & ~n4981;
  assign n4984 = ~n4982 & n4983;
  assign n4985 = ~n4980 & n4984;
  assign n4986 = ~n4976 & ~n4985;
  assign n4987 = ~n4975 & ~n4986;
  assign n4988 = n4827 & ~n4987;
  assign n4989 = ~n4825 & ~n4988;
  assign n4990 = n4776 & n4785;
  assign n4991 = ~n4786 & ~n4990;
  assign n4992 = ~n4989 & n4991;
  assign n4993 = ~n4786 & ~n4992;
  assign n4994 = ~n4758 & ~n4759;
  assign n4995 = ~n4768 & n4994;
  assign n4996 = n4768 & ~n4994;
  assign n4997 = ~n4995 & ~n4996;
  assign n4998 = ~n4993 & n4997;
  assign n4999 = n4993 & ~n4997;
  assign n5000 = ~n4998 & ~n4999;
  assign n5001 = ~n1533 & n3884;
  assign n5002 = n3886 & n4355;
  assign n5003 = ~n1637 & n3810;
  assign n5004 = ~n1448 & n4380;
  assign n5005 = ~n5001 & ~n5003;
  assign n5006 = ~n5004 & n5005;
  assign n5007 = ~n5002 & n5006;
  assign n5008 = pi29  & n5007;
  assign n5009 = ~pi29  & ~n5007;
  assign n5010 = ~n5008 & ~n5009;
  assign n5011 = n5000 & ~n5010;
  assign n5012 = ~n4998 & ~n5011;
  assign n5013 = n4773 & ~n5012;
  assign n5014 = ~n4771 & ~n5013;
  assign n5015 = ~n4684 & ~n5014;
  assign n5016 = ~n4681 & ~n5015;
  assign n5017 = ~n4564 & n4574;
  assign n5018 = ~n4575 & ~n5017;
  assign n5019 = ~n5016 & n5018;
  assign n5020 = n86 & ~n878;
  assign n5021 = n3687 & n4420;
  assign n5022 = ~n987 & n4600;
  assign n5023 = ~n3681 & n4615;
  assign n5024 = ~n5020 & ~n5022;
  assign n5025 = ~n5023 & n5024;
  assign n5026 = ~n5021 & n5025;
  assign n5027 = ~pi26  & ~n5026;
  assign n5028 = pi26  & n5026;
  assign n5029 = ~n5027 & ~n5028;
  assign n5030 = n5016 & ~n5018;
  assign n5031 = ~n5019 & ~n5030;
  assign n5032 = ~n5029 & n5031;
  assign n5033 = ~n5019 & ~n5032;
  assign n5034 = ~pi22  & pi23 ;
  assign n5035 = pi22  & ~pi23 ;
  assign n5036 = ~n5034 & ~n5035;
  assign n5037 = ~pi21  & pi22 ;
  assign n5038 = pi21  & ~pi22 ;
  assign n5039 = ~n5037 & ~n5038;
  assign n5040 = pi20  & ~pi21 ;
  assign n5041 = ~pi20  & pi21 ;
  assign n5042 = ~n5040 & ~n5041;
  assign n5043 = n5039 & n5042;
  assign n5044 = ~n5036 & n5043;
  assign n5045 = ~n5036 & ~n5042;
  assign n5046 = ~n3897 & n5045;
  assign n5047 = ~n5044 & ~n5046;
  assign n5048 = ~n3883 & ~n5047;
  assign n5049 = pi23  & ~n5048;
  assign n5050 = ~pi23  & n5048;
  assign n5051 = ~n5049 & ~n5050;
  assign n5052 = n5033 & n5051;
  assign n5053 = ~n5033 & ~n5051;
  assign n5054 = ~n4638 & ~n4639;
  assign n5055 = ~n4649 & ~n5054;
  assign n5056 = n4649 & n5054;
  assign n5057 = ~n5055 & ~n5056;
  assign n5058 = ~n5053 & n5057;
  assign n5059 = ~n5052 & ~n5058;
  assign n5060 = n4666 & n5059;
  assign n5061 = n4684 & n5014;
  assign n5062 = ~n5015 & ~n5061;
  assign n5063 = ~n987 & n4615;
  assign n5064 = n3791 & n4420;
  assign n5065 = n86 & ~n1104;
  assign n5066 = ~n878 & n4600;
  assign n5067 = ~n5063 & ~n5065;
  assign n5068 = ~n5066 & n5067;
  assign n5069 = ~n5064 & n5068;
  assign n5070 = pi26  & n5069;
  assign n5071 = ~pi26  & ~n5069;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = n5062 & ~n5072;
  assign n5074 = n5062 & n5072;
  assign n5075 = ~n5062 & ~n5072;
  assign n5076 = ~n5074 & ~n5075;
  assign n5077 = ~n4773 & n5012;
  assign n5078 = ~n5013 & ~n5077;
  assign n5079 = ~n1448 & n3884;
  assign n5080 = n3886 & n4453;
  assign n5081 = ~n1533 & n3810;
  assign n5082 = ~n1345 & n4380;
  assign n5083 = ~n5079 & ~n5081;
  assign n5084 = ~n5082 & n5083;
  assign n5085 = ~n5080 & n5084;
  assign n5086 = pi29  & n5085;
  assign n5087 = ~pi29  & ~n5085;
  assign n5088 = ~n5086 & ~n5087;
  assign n5089 = n5078 & ~n5088;
  assign n5090 = ~n1104 & n4600;
  assign n5091 = n3775 & n4420;
  assign n5092 = n86 & ~n1225;
  assign n5093 = ~n878 & n4615;
  assign n5094 = ~n5090 & ~n5092;
  assign n5095 = ~n5093 & n5094;
  assign n5096 = ~n5091 & n5095;
  assign n5097 = pi26  & n5096;
  assign n5098 = ~pi26  & ~n5096;
  assign n5099 = ~n5097 & ~n5098;
  assign n5100 = ~n5078 & n5088;
  assign n5101 = ~n5099 & ~n5100;
  assign n5102 = ~n5089 & ~n5101;
  assign n5103 = ~n5076 & ~n5102;
  assign n5104 = ~n5073 & ~n5103;
  assign n5105 = n5029 & ~n5031;
  assign n5106 = ~n5032 & ~n5105;
  assign n5107 = ~n5104 & n5106;
  assign n5108 = ~n3855 & n5044;
  assign n5109 = ~n5039 & n5042;
  assign n5110 = ~n3883 & n5109;
  assign n5111 = ~n3900 & n5045;
  assign n5112 = ~n5108 & ~n5110;
  assign n5113 = ~n5111 & n5112;
  assign n5114 = ~pi23  & ~n5113;
  assign n5115 = pi23  & n5113;
  assign n5116 = ~n5114 & ~n5115;
  assign n5117 = n5104 & ~n5106;
  assign n5118 = ~n5107 & ~n5117;
  assign n5119 = ~n5116 & n5118;
  assign n5120 = ~n5107 & ~n5119;
  assign n5121 = ~n5052 & ~n5053;
  assign n5122 = ~n5057 & n5121;
  assign n5123 = n5057 & ~n5121;
  assign n5124 = ~n5122 & ~n5123;
  assign n5125 = ~n5120 & n5124;
  assign n5126 = n5120 & ~n5124;
  assign n5127 = ~n5125 & ~n5126;
  assign n5128 = n5116 & ~n5118;
  assign n5129 = ~n5119 & ~n5128;
  assign n5130 = n5036 & ~n5042;
  assign n5131 = ~n3883 & n5130;
  assign n5132 = n4399 & n5045;
  assign n5133 = ~n3855 & n5109;
  assign n5134 = ~n3681 & n5044;
  assign n5135 = ~n5131 & ~n5133;
  assign n5136 = ~n5134 & n5135;
  assign n5137 = ~n5132 & n5136;
  assign n5138 = pi23  & n5137;
  assign n5139 = ~pi23  & ~n5137;
  assign n5140 = ~n5138 & ~n5139;
  assign n5141 = ~n5089 & ~n5100;
  assign n5142 = n5099 & ~n5141;
  assign n5143 = ~n5099 & n5141;
  assign n5144 = ~n5142 & ~n5143;
  assign n5145 = ~n5000 & n5010;
  assign n5146 = ~n5011 & ~n5145;
  assign n5147 = ~n4827 & n4987;
  assign n5148 = ~n4988 & ~n5147;
  assign n5149 = n748 & ~n2098;
  assign n5150 = n3560 & ~n3562;
  assign n5151 = ~n3563 & ~n5150;
  assign n5152 = n880 & n5151;
  assign n5153 = ~n1998 & n3692;
  assign n5154 = ~n1908 & n3694;
  assign n5155 = ~n5149 & ~n5153;
  assign n5156 = ~n5154 & n5155;
  assign n5157 = ~n5152 & n5156;
  assign n5158 = n5148 & ~n5157;
  assign n5159 = ~n1717 & n3884;
  assign n5160 = n3886 & n4537;
  assign n5161 = ~n1841 & n3810;
  assign n5162 = ~n1637 & n4380;
  assign n5163 = ~n5159 & ~n5161;
  assign n5164 = ~n5162 & n5163;
  assign n5165 = ~n5160 & n5164;
  assign n5166 = ~pi29  & ~n5165;
  assign n5167 = pi29  & n5165;
  assign n5168 = ~n5166 & ~n5167;
  assign n5169 = n5148 & n5157;
  assign n5170 = ~n5148 & ~n5157;
  assign n5171 = ~n5169 & ~n5170;
  assign n5172 = ~n5168 & ~n5171;
  assign n5173 = ~n5158 & ~n5172;
  assign n5174 = n4989 & ~n4991;
  assign n5175 = ~n4992 & ~n5174;
  assign n5176 = ~n5173 & n5175;
  assign n5177 = ~n1637 & n3884;
  assign n5178 = n3886 & n4553;
  assign n5179 = ~n1717 & n3810;
  assign n5180 = ~n1533 & n4380;
  assign n5181 = ~n5177 & ~n5179;
  assign n5182 = ~n5180 & n5181;
  assign n5183 = ~n5178 & n5182;
  assign n5184 = pi29  & n5183;
  assign n5185 = ~pi29  & ~n5183;
  assign n5186 = ~n5184 & ~n5185;
  assign n5187 = n5173 & ~n5175;
  assign n5188 = ~n5186 & ~n5187;
  assign n5189 = ~n5176 & ~n5188;
  assign n5190 = n5146 & ~n5189;
  assign n5191 = ~n5146 & n5189;
  assign n5192 = ~n1225 & n4600;
  assign n5193 = n4135 & n4420;
  assign n5194 = n86 & ~n1345;
  assign n5195 = ~n1104 & n4615;
  assign n5196 = ~n5192 & ~n5194;
  assign n5197 = ~n5195 & n5196;
  assign n5198 = ~n5193 & n5197;
  assign n5199 = pi26  & n5198;
  assign n5200 = ~pi26  & ~n5198;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = ~n5191 & ~n5201;
  assign n5203 = ~n5190 & ~n5202;
  assign n5204 = n5144 & ~n5203;
  assign n5205 = ~n5144 & n5203;
  assign n5206 = ~n3855 & n5130;
  assign n5207 = n3972 & n5045;
  assign n5208 = ~n987 & n5044;
  assign n5209 = ~n3681 & n5109;
  assign n5210 = ~n5206 & ~n5208;
  assign n5211 = ~n5209 & n5210;
  assign n5212 = ~n5207 & n5211;
  assign n5213 = pi23  & n5212;
  assign n5214 = ~pi23  & ~n5212;
  assign n5215 = ~n5213 & ~n5214;
  assign n5216 = ~n5205 & ~n5215;
  assign n5217 = ~n5204 & ~n5216;
  assign n5218 = ~n5140 & ~n5217;
  assign n5219 = n5140 & n5217;
  assign n5220 = n5076 & ~n5102;
  assign n5221 = ~n5076 & n5102;
  assign n5222 = ~n5220 & ~n5221;
  assign n5223 = ~n5219 & ~n5222;
  assign n5224 = ~n5218 & ~n5223;
  assign n5225 = n5129 & ~n5224;
  assign n5226 = ~n5218 & ~n5219;
  assign n5227 = ~n5222 & n5226;
  assign n5228 = n5222 & ~n5226;
  assign n5229 = ~n5227 & ~n5228;
  assign n5230 = pi19  & ~pi20 ;
  assign n5231 = ~pi19  & pi20 ;
  assign n5232 = ~n5230 & ~n5231;
  assign n5233 = pi17  & ~pi18 ;
  assign n5234 = ~pi17  & pi18 ;
  assign n5235 = ~n5233 & ~n5234;
  assign n5236 = ~pi18  & pi19 ;
  assign n5237 = pi18  & ~pi19 ;
  assign n5238 = ~n5236 & ~n5237;
  assign n5239 = n5235 & n5238;
  assign n5240 = ~n5232 & n5239;
  assign n5241 = ~n5232 & ~n5235;
  assign n5242 = ~n3897 & n5241;
  assign n5243 = ~n5240 & ~n5242;
  assign n5244 = ~n3883 & ~n5243;
  assign n5245 = pi20  & ~n5244;
  assign n5246 = ~pi20  & n5244;
  assign n5247 = ~n5245 & ~n5246;
  assign n5248 = ~n1345 & n4600;
  assign n5249 = n4152 & n4420;
  assign n5250 = n86 & ~n1448;
  assign n5251 = ~n1225 & n4615;
  assign n5252 = ~n5248 & ~n5250;
  assign n5253 = ~n5251 & n5252;
  assign n5254 = ~n5249 & n5253;
  assign n5255 = pi26  & n5254;
  assign n5256 = ~pi26  & ~n5254;
  assign n5257 = ~n5255 & ~n5256;
  assign n5258 = ~n5176 & ~n5187;
  assign n5259 = n5186 & ~n5258;
  assign n5260 = ~n5186 & n5258;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = ~n5257 & n5261;
  assign n5263 = n5257 & ~n5261;
  assign n5264 = ~n5262 & ~n5263;
  assign n5265 = ~n4975 & ~n4976;
  assign n5266 = ~n4985 & n5265;
  assign n5267 = n4985 & ~n5265;
  assign n5268 = ~n5266 & ~n5267;
  assign n5269 = ~n116 & ~n646;
  assign n5270 = n1293 & n5269;
  assign n5271 = ~n381 & ~n592;
  assign n5272 = ~n212 & n1428;
  assign n5273 = n1475 & n5272;
  assign n5274 = ~n445 & ~n1699;
  assign n5275 = n366 & n5274;
  assign n5276 = n719 & n1014;
  assign n5277 = n1890 & n2625;
  assign n5278 = n3325 & n4004;
  assign n5279 = n4687 & n5271;
  assign n5280 = n5278 & n5279;
  assign n5281 = n5276 & n5277;
  assign n5282 = n5270 & n5275;
  assign n5283 = n5281 & n5282;
  assign n5284 = n1514 & n5280;
  assign n5285 = n5273 & n5284;
  assign n5286 = n5283 & n5285;
  assign n5287 = ~n512 & ~n700;
  assign n5288 = ~n715 & ~n751;
  assign n5289 = ~n944 & n5288;
  assign n5290 = n5287 & n5289;
  assign n5291 = ~n239 & ~n488;
  assign n5292 = ~n523 & ~n894;
  assign n5293 = n5291 & n5292;
  assign n5294 = n598 & n1243;
  assign n5295 = n3301 & n5294;
  assign n5296 = n3471 & n5293;
  assign n5297 = n5295 & n5296;
  assign n5298 = n5290 & n5297;
  assign n5299 = ~n318 & ~n810;
  assign n5300 = ~n430 & ~n625;
  assign n5301 = ~n236 & ~n293;
  assign n5302 = ~n304 & ~n377;
  assign n5303 = n5301 & n5302;
  assign n5304 = n1725 & n4163;
  assign n5305 = n5303 & n5304;
  assign n5306 = ~n273 & n505;
  assign n5307 = n755 & n5306;
  assign n5308 = ~n159 & ~n170;
  assign n5309 = ~n200 & ~n258;
  assign n5310 = ~n414 & ~n601;
  assign n5311 = n5309 & n5310;
  assign n5312 = n150 & n5308;
  assign n5313 = n360 & n881;
  assign n5314 = n1476 & n1492;
  assign n5315 = n1859 & n5314;
  assign n5316 = n5312 & n5313;
  assign n5317 = n485 & n5311;
  assign n5318 = n1406 & n5317;
  assign n5319 = n5315 & n5316;
  assign n5320 = n5307 & n5319;
  assign n5321 = n3731 & n5318;
  assign n5322 = n5320 & n5321;
  assign n5323 = ~n106 & ~n177;
  assign n5324 = ~n248 & ~n532;
  assign n5325 = ~n563 & n5324;
  assign n5326 = n1244 & n5323;
  assign n5327 = n1575 & n3205;
  assign n5328 = n5299 & n5300;
  assign n5329 = n5327 & n5328;
  assign n5330 = n5325 & n5326;
  assign n5331 = n1119 & n5330;
  assign n5332 = n2759 & n5329;
  assign n5333 = n5305 & n5332;
  assign n5334 = n5331 & n5333;
  assign n5335 = n5298 & n5334;
  assign n5336 = n5286 & n5322;
  assign n5337 = n5335 & n5336;
  assign n5338 = n4904 & ~n5337;
  assign n5339 = ~n4904 & n5337;
  assign n5340 = ~n5338 & ~n5339;
  assign n5341 = ~n2146 & n3694;
  assign n5342 = n3548 & ~n3550;
  assign n5343 = ~n3551 & ~n5342;
  assign n5344 = n880 & n5343;
  assign n5345 = n748 & ~n2347;
  assign n5346 = ~n2249 & n3692;
  assign n5347 = ~n5341 & ~n5345;
  assign n5348 = ~n5346 & n5347;
  assign n5349 = ~n5344 & n5348;
  assign n5350 = n5340 & ~n5349;
  assign n5351 = ~n5338 & ~n5350;
  assign n5352 = ~pi14  & ~n4973;
  assign n5353 = ~n4971 & n4974;
  assign n5354 = ~n5352 & ~n5353;
  assign n5355 = ~n5351 & ~n5354;
  assign n5356 = n5351 & n5354;
  assign n5357 = ~n2098 & n3694;
  assign n5358 = n3552 & ~n3554;
  assign n5359 = ~n3555 & ~n5358;
  assign n5360 = n880 & n5359;
  assign n5361 = ~n2146 & n3692;
  assign n5362 = n748 & ~n2249;
  assign n5363 = ~n5357 & ~n5361;
  assign n5364 = ~n5362 & n5363;
  assign n5365 = ~n5360 & n5364;
  assign n5366 = ~n5356 & ~n5365;
  assign n5367 = ~n5355 & ~n5366;
  assign n5368 = n5268 & ~n5367;
  assign n5369 = ~n5268 & n5367;
  assign n5370 = ~n5368 & ~n5369;
  assign n5371 = ~n1841 & n3884;
  assign n5372 = n3886 & n4762;
  assign n5373 = ~n1908 & n3810;
  assign n5374 = ~n1717 & n4380;
  assign n5375 = ~n5371 & ~n5373;
  assign n5376 = ~n5374 & n5375;
  assign n5377 = ~n5372 & n5376;
  assign n5378 = pi29  & n5377;
  assign n5379 = ~pi29  & ~n5377;
  assign n5380 = ~n5378 & ~n5379;
  assign n5381 = n5370 & ~n5380;
  assign n5382 = ~n5368 & ~n5381;
  assign n5383 = n5168 & n5171;
  assign n5384 = ~n5172 & ~n5383;
  assign n5385 = ~n5382 & n5384;
  assign n5386 = n5382 & ~n5384;
  assign n5387 = ~n1448 & n4600;
  assign n5388 = n4420 & n4453;
  assign n5389 = n86 & ~n1533;
  assign n5390 = ~n1345 & n4615;
  assign n5391 = ~n5387 & ~n5389;
  assign n5392 = ~n5390 & n5391;
  assign n5393 = ~n5388 & n5392;
  assign n5394 = pi26  & n5393;
  assign n5395 = ~pi26  & ~n5393;
  assign n5396 = ~n5394 & ~n5395;
  assign n5397 = ~n5386 & ~n5396;
  assign n5398 = ~n5385 & ~n5397;
  assign n5399 = n5264 & ~n5398;
  assign n5400 = ~n5262 & ~n5399;
  assign n5401 = ~n5190 & ~n5191;
  assign n5402 = ~n5201 & n5401;
  assign n5403 = n5201 & ~n5401;
  assign n5404 = ~n5402 & ~n5403;
  assign n5405 = ~n5400 & n5404;
  assign n5406 = n5400 & ~n5404;
  assign n5407 = ~n878 & n5044;
  assign n5408 = n3687 & n5045;
  assign n5409 = ~n987 & n5109;
  assign n5410 = ~n3681 & n5130;
  assign n5411 = ~n5407 & ~n5409;
  assign n5412 = ~n5410 & n5411;
  assign n5413 = ~n5408 & n5412;
  assign n5414 = pi23  & n5413;
  assign n5415 = ~pi23  & ~n5413;
  assign n5416 = ~n5414 & ~n5415;
  assign n5417 = ~n5406 & ~n5416;
  assign n5418 = ~n5405 & ~n5417;
  assign n5419 = ~n5247 & ~n5418;
  assign n5420 = n5247 & n5418;
  assign n5421 = ~n5204 & ~n5205;
  assign n5422 = ~n5215 & n5421;
  assign n5423 = n5215 & ~n5421;
  assign n5424 = ~n5422 & ~n5423;
  assign n5425 = ~n5420 & n5424;
  assign n5426 = ~n5419 & ~n5425;
  assign n5427 = n5229 & ~n5426;
  assign n5428 = ~n5229 & n5426;
  assign n5429 = ~n5427 & ~n5428;
  assign n5430 = ~n5419 & ~n5420;
  assign n5431 = n5424 & n5430;
  assign n5432 = ~n5424 & ~n5430;
  assign n5433 = ~n5431 & ~n5432;
  assign n5434 = ~n987 & n5130;
  assign n5435 = n3791 & n5045;
  assign n5436 = ~n1104 & n5044;
  assign n5437 = ~n878 & n5109;
  assign n5438 = ~n5434 & ~n5436;
  assign n5439 = ~n5437 & n5438;
  assign n5440 = ~n5435 & n5439;
  assign n5441 = ~pi23  & ~n5440;
  assign n5442 = pi23  & n5440;
  assign n5443 = ~n5441 & ~n5442;
  assign n5444 = ~n5264 & n5398;
  assign n5445 = ~n5399 & ~n5444;
  assign n5446 = ~n5443 & n5445;
  assign n5447 = ~n5443 & ~n5445;
  assign n5448 = n5443 & n5445;
  assign n5449 = ~n5447 & ~n5448;
  assign n5450 = ~n5385 & ~n5386;
  assign n5451 = ~n5396 & n5450;
  assign n5452 = n5396 & ~n5450;
  assign n5453 = ~n5451 & ~n5452;
  assign n5454 = ~n1908 & n3884;
  assign n5455 = n3886 & n4779;
  assign n5456 = ~n1998 & n3810;
  assign n5457 = ~n1841 & n4380;
  assign n5458 = ~n5454 & ~n5456;
  assign n5459 = ~n5457 & n5458;
  assign n5460 = ~n5455 & n5459;
  assign n5461 = ~pi29  & ~n5460;
  assign n5462 = pi29  & n5460;
  assign n5463 = ~n5461 & ~n5462;
  assign n5464 = ~n5355 & ~n5356;
  assign n5465 = ~n5365 & n5464;
  assign n5466 = n5365 & ~n5464;
  assign n5467 = ~n5465 & ~n5466;
  assign n5468 = ~n5463 & n5467;
  assign n5469 = ~n5463 & ~n5467;
  assign n5470 = n5463 & n5467;
  assign n5471 = ~n5469 & ~n5470;
  assign n5472 = ~n5340 & n5349;
  assign n5473 = ~n5350 & ~n5472;
  assign n5474 = ~n250 & ~n377;
  assign n5475 = n942 & n4926;
  assign n5476 = ~n270 & ~n365;
  assign n5477 = ~n537 & n5476;
  assign n5478 = n298 & n1087;
  assign n5479 = n1198 & n3858;
  assign n5480 = n5474 & n5479;
  assign n5481 = n5477 & n5478;
  assign n5482 = n3244 & n5475;
  assign n5483 = n5481 & n5482;
  assign n5484 = n5480 & n5483;
  assign n5485 = n501 & ~n656;
  assign n5486 = n1913 & n5485;
  assign n5487 = ~n211 & ~n798;
  assign n5488 = ~n1051 & n5487;
  assign n5489 = ~n604 & ~n1487;
  assign n5490 = ~n271 & ~n319;
  assign n5491 = ~n330 & ~n534;
  assign n5492 = n2561 & n5491;
  assign n5493 = n2802 & n5490;
  assign n5494 = n5492 & n5493;
  assign n5495 = ~n175 & ~n1404;
  assign n5496 = ~n723 & n5495;
  assign n5497 = ~n236 & ~n437;
  assign n5498 = ~n511 & ~n753;
  assign n5499 = n5497 & n5498;
  assign n5500 = n1564 & n1729;
  assign n5501 = n4063 & n5489;
  assign n5502 = n5500 & n5501;
  assign n5503 = n118 & n5499;
  assign n5504 = n2657 & n5496;
  assign n5505 = n5503 & n5504;
  assign n5506 = n5494 & n5502;
  assign n5507 = n5505 & n5506;
  assign n5508 = ~n93 & ~n408;
  assign n5509 = ~n532 & n5508;
  assign n5510 = ~n139 & ~n237;
  assign n5511 = ~n376 & ~n596;
  assign n5512 = n5510 & n5511;
  assign n5513 = n633 & n1730;
  assign n5514 = n5512 & n5513;
  assign n5515 = n5488 & n5509;
  assign n5516 = n5514 & n5515;
  assign n5517 = n5486 & n5516;
  assign n5518 = n2458 & n4886;
  assign n5519 = n5517 & n5518;
  assign n5520 = n5484 & n5507;
  assign n5521 = n5519 & n5520;
  assign n5522 = n1376 & n5521;
  assign n5523 = ~n155 & ~n299;
  assign n5524 = ~n139 & ~n281;
  assign n5525 = ~n532 & ~n937;
  assign n5526 = n5524 & n5525;
  assign n5527 = ~n258 & ~n338;
  assign n5528 = ~n529 & n5527;
  assign n5529 = n704 & n1864;
  assign n5530 = n3326 & n4163;
  assign n5531 = n5529 & n5530;
  assign n5532 = n5526 & n5528;
  assign n5533 = n5531 & n5532;
  assign n5534 = ~n111 & ~n604;
  assign n5535 = ~n792 & n5534;
  assign n5536 = ~n190 & ~n293;
  assign n5537 = ~n319 & ~n355;
  assign n5538 = ~n359 & ~n381;
  assign n5539 = n2637 & n5538;
  assign n5540 = n5536 & n5537;
  assign n5541 = n375 & n602;
  assign n5542 = n2197 & n2529;
  assign n5543 = n2534 & n5523;
  assign n5544 = n5542 & n5543;
  assign n5545 = n5540 & n5541;
  assign n5546 = n5535 & n5539;
  assign n5547 = n5545 & n5546;
  assign n5548 = n1679 & n5544;
  assign n5549 = n5547 & n5548;
  assign n5550 = n5533 & n5549;
  assign n5551 = ~n328 & ~n592;
  assign n5552 = ~n718 & ~n754;
  assign n5553 = ~n770 & n5552;
  assign n5554 = n354 & n5551;
  assign n5555 = n479 & n815;
  assign n5556 = n1423 & n1729;
  assign n5557 = n1812 & n1962;
  assign n5558 = n2934 & n4864;
  assign n5559 = n5557 & n5558;
  assign n5560 = n5555 & n5556;
  assign n5561 = n5553 & n5554;
  assign n5562 = n2023 & n3936;
  assign n5563 = n5561 & n5562;
  assign n5564 = n5559 & n5560;
  assign n5565 = n5563 & n5564;
  assign n5566 = n4233 & n5565;
  assign n5567 = n4014 & n5484;
  assign n5568 = n5566 & n5567;
  assign n5569 = n5550 & n5568;
  assign n5570 = ~n5522 & ~n5569;
  assign n5571 = n5522 & n5569;
  assign n5572 = ~pi11  & ~n5570;
  assign n5573 = ~n5571 & n5572;
  assign n5574 = ~n5570 & ~n5573;
  assign n5575 = n4904 & ~n5574;
  assign n5576 = ~n4904 & n5574;
  assign n5577 = n748 & ~n2412;
  assign n5578 = n3544 & ~n3546;
  assign n5579 = ~n3547 & ~n5578;
  assign n5580 = n880 & n5579;
  assign n5581 = ~n2347 & n3692;
  assign n5582 = ~n2249 & n3694;
  assign n5583 = ~n5577 & ~n5581;
  assign n5584 = ~n5582 & n5583;
  assign n5585 = ~n5580 & n5584;
  assign n5586 = ~n5576 & ~n5585;
  assign n5587 = ~n5575 & ~n5586;
  assign n5588 = n5473 & ~n5587;
  assign n5589 = ~n5473 & n5587;
  assign n5590 = ~n5588 & ~n5589;
  assign n5591 = ~pi11  & ~n5573;
  assign n5592 = ~n5571 & n5574;
  assign n5593 = ~n5591 & ~n5592;
  assign n5594 = ~n2347 & n3694;
  assign n5595 = n3540 & ~n3542;
  assign n5596 = ~n3543 & ~n5595;
  assign n5597 = n880 & n5596;
  assign n5598 = n748 & ~n2496;
  assign n5599 = ~n2412 & n3692;
  assign n5600 = ~n5594 & ~n5598;
  assign n5601 = ~n5599 & n5600;
  assign n5602 = ~n5597 & n5601;
  assign n5603 = ~n5593 & ~n5602;
  assign n5604 = ~n646 & ~n1032;
  assign n5605 = ~n352 & ~n481;
  assign n5606 = n2108 & n5605;
  assign n5607 = n5604 & n5606;
  assign n5608 = ~n156 & ~n235;
  assign n5609 = n146 & n5608;
  assign n5610 = ~n309 & ~n445;
  assign n5611 = n117 & n5610;
  assign n5612 = ~n271 & ~n486;
  assign n5613 = ~n488 & ~n627;
  assign n5614 = ~n656 & ~n751;
  assign n5615 = ~n1404 & n5614;
  assign n5616 = n5612 & n5613;
  assign n5617 = n2757 & n3224;
  assign n5618 = n5616 & n5617;
  assign n5619 = n1849 & n5615;
  assign n5620 = n5609 & n5611;
  assign n5621 = n5619 & n5620;
  assign n5622 = n5607 & n5618;
  assign n5623 = n5621 & n5622;
  assign n5624 = n4002 & n5623;
  assign n5625 = n2423 & n5624;
  assign n5626 = n2471 & n5625;
  assign n5627 = n1811 & n5626;
  assign n5628 = n5522 & ~n5627;
  assign n5629 = ~n5522 & n5627;
  assign n5630 = ~n5628 & ~n5629;
  assign n5631 = ~n304 & ~n310;
  assign n5632 = n448 & n5631;
  assign n5633 = ~n216 & ~n356;
  assign n5634 = ~n893 & ~n1002;
  assign n5635 = n5633 & n5634;
  assign n5636 = n375 & n1539;
  assign n5637 = n1685 & n1863;
  assign n5638 = n3225 & n3432;
  assign n5639 = n4063 & n5638;
  assign n5640 = n5636 & n5637;
  assign n5641 = n3018 & n5635;
  assign n5642 = n5632 & n5641;
  assign n5643 = n5639 & n5640;
  assign n5644 = n5642 & n5643;
  assign n5645 = n4924 & n5644;
  assign n5646 = ~n564 & n5271;
  assign n5647 = ~n509 & ~n894;
  assign n5648 = n3121 & n5647;
  assign n5649 = n5646 & n5648;
  assign n5650 = ~n376 & ~n515;
  assign n5651 = ~n149 & ~n248;
  assign n5652 = ~n435 & ~n522;
  assign n5653 = ~n648 & ~n685;
  assign n5654 = ~n698 & ~n937;
  assign n5655 = n5653 & n5654;
  assign n5656 = n5651 & n5652;
  assign n5657 = n5655 & n5656;
  assign n5658 = n4068 & n5657;
  assign n5659 = ~n130 & ~n308;
  assign n5660 = ~n486 & ~n568;
  assign n5661 = n5659 & n5660;
  assign n5662 = n4802 & n5661;
  assign n5663 = n2982 & n5662;
  assign n5664 = ~n129 & ~n174;
  assign n5665 = ~n247 & ~n353;
  assign n5666 = ~n638 & ~n661;
  assign n5667 = ~n841 & n5666;
  assign n5668 = n5664 & n5665;
  assign n5669 = n645 & n769;
  assign n5670 = n1246 & n5669;
  assign n5671 = n5667 & n5668;
  assign n5672 = n2001 & n4845;
  assign n5673 = n5671 & n5672;
  assign n5674 = n1961 & n5670;
  assign n5675 = n5673 & n5674;
  assign n5676 = n5658 & n5663;
  assign n5677 = n5675 & n5676;
  assign n5678 = ~n333 & ~n508;
  assign n5679 = ~n196 & ~n364;
  assign n5680 = ~n416 & ~n902;
  assign n5681 = n5679 & n5680;
  assign n5682 = n433 & n797;
  assign n5683 = n898 & n2052;
  assign n5684 = n3934 & n5683;
  assign n5685 = n5681 & n5682;
  assign n5686 = n5684 & n5685;
  assign n5687 = ~n319 & ~n339;
  assign n5688 = ~n721 & n5687;
  assign n5689 = n2503 & n2838;
  assign n5690 = n4003 & n5689;
  assign n5691 = n5688 & n5690;
  assign n5692 = ~n162 & ~n237;
  assign n5693 = ~n814 & n5692;
  assign n5694 = n2148 & n5650;
  assign n5695 = n5678 & n5694;
  assign n5696 = n1641 & n5693;
  assign n5697 = n5535 & n5696;
  assign n5698 = n2655 & n5695;
  assign n5699 = n5649 & n5698;
  assign n5700 = n5686 & n5697;
  assign n5701 = n5691 & n5700;
  assign n5702 = n5699 & n5701;
  assign n5703 = n5645 & n5677;
  assign n5704 = n5702 & n5703;
  assign n5705 = ~n190 & ~n269;
  assign n5706 = ~n537 & ~n808;
  assign n5707 = ~n1032 & n5706;
  assign n5708 = n521 & n5705;
  assign n5709 = n845 & n1684;
  assign n5710 = n2024 & n2451;
  assign n5711 = n5709 & n5710;
  assign n5712 = n5707 & n5708;
  assign n5713 = n5711 & n5712;
  assign n5714 = ~n135 & ~n1086;
  assign n5715 = n483 & n5714;
  assign n5716 = n749 & n1429;
  assign n5717 = n5715 & n5716;
  assign n5718 = ~n156 & ~n1051;
  assign n5719 = n1151 & n5718;
  assign n5720 = ~n212 & ~n318;
  assign n5721 = ~n174 & ~n200;
  assign n5722 = ~n294 & ~n312;
  assign n5723 = ~n352 & ~n374;
  assign n5724 = n5722 & n5723;
  assign n5725 = n750 & n5721;
  assign n5726 = n1291 & n3122;
  assign n5727 = n5720 & n5726;
  assign n5728 = n5724 & n5725;
  assign n5729 = n5727 & n5728;
  assign n5730 = ~n98 & ~n175;
  assign n5731 = ~n249 & ~n510;
  assign n5732 = ~n531 & ~n663;
  assign n5733 = n5731 & n5732;
  assign n5734 = n487 & n5730;
  assign n5735 = n704 & n1047;
  assign n5736 = n1246 & n2473;
  assign n5737 = n5735 & n5736;
  assign n5738 = n5733 & n5734;
  assign n5739 = n854 & n5719;
  assign n5740 = n5738 & n5739;
  assign n5741 = n4478 & n5737;
  assign n5742 = n5717 & n5741;
  assign n5743 = n5729 & n5740;
  assign n5744 = n5742 & n5743;
  assign n5745 = ~n184 & ~n236;
  assign n5746 = ~n416 & ~n566;
  assign n5747 = ~n646 & ~n1699;
  assign n5748 = n5746 & n5747;
  assign n5749 = n2206 & n5745;
  assign n5750 = n4905 & n5749;
  assign n5751 = n5748 & n5750;
  assign n5752 = ~n253 & ~n359;
  assign n5753 = ~n634 & ~n814;
  assign n5754 = n5752 & n5753;
  assign n5755 = n292 & n357;
  assign n5756 = n722 & n1005;
  assign n5757 = n1242 & n3374;
  assign n5758 = n5756 & n5757;
  assign n5759 = n5754 & n5755;
  assign n5760 = n3343 & n5759;
  assign n5761 = n4476 & n5758;
  assign n5762 = n5760 & n5761;
  assign n5763 = n5713 & n5751;
  assign n5764 = n5762 & n5763;
  assign n5765 = n4518 & n5764;
  assign n5766 = n5744 & n5765;
  assign n5767 = ~n5704 & ~n5766;
  assign n5768 = n5704 & n5766;
  assign n5769 = ~pi8  & ~n5767;
  assign n5770 = ~n5768 & n5769;
  assign n5771 = ~n5767 & ~n5770;
  assign n5772 = n5522 & ~n5771;
  assign n5773 = ~n5522 & n5771;
  assign n5774 = ~n2496 & n3694;
  assign n5775 = n3532 & ~n3534;
  assign n5776 = ~n3535 & ~n5775;
  assign n5777 = n880 & n5776;
  assign n5778 = n748 & ~n2674;
  assign n5779 = ~n2589 & n3692;
  assign n5780 = ~n5774 & ~n5778;
  assign n5781 = ~n5779 & n5780;
  assign n5782 = ~n5777 & n5781;
  assign n5783 = ~n5773 & ~n5782;
  assign n5784 = ~n5772 & ~n5783;
  assign n5785 = n5630 & ~n5784;
  assign n5786 = ~n5628 & ~n5785;
  assign n5787 = n5593 & n5602;
  assign n5788 = ~n5603 & ~n5787;
  assign n5789 = ~n5786 & n5788;
  assign n5790 = ~n5603 & ~n5789;
  assign n5791 = ~n5575 & ~n5576;
  assign n5792 = ~n5585 & n5791;
  assign n5793 = n5585 & ~n5791;
  assign n5794 = ~n5792 & ~n5793;
  assign n5795 = ~n5790 & n5794;
  assign n5796 = n5790 & ~n5794;
  assign n5797 = ~n5795 & ~n5796;
  assign n5798 = ~n2098 & n3884;
  assign n5799 = n3886 & n4979;
  assign n5800 = ~n2146 & n3810;
  assign n5801 = ~n1998 & n4380;
  assign n5802 = ~n5798 & ~n5800;
  assign n5803 = ~n5801 & n5802;
  assign n5804 = ~n5799 & n5803;
  assign n5805 = pi29  & n5804;
  assign n5806 = ~pi29  & ~n5804;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = n5797 & ~n5807;
  assign n5809 = ~n5795 & ~n5808;
  assign n5810 = n5590 & ~n5809;
  assign n5811 = ~n5588 & ~n5810;
  assign n5812 = ~n5471 & ~n5811;
  assign n5813 = ~n5468 & ~n5812;
  assign n5814 = ~n5370 & n5380;
  assign n5815 = ~n5381 & ~n5814;
  assign n5816 = ~n5813 & n5815;
  assign n5817 = n5813 & ~n5815;
  assign n5818 = ~n1533 & n4600;
  assign n5819 = n4355 & n4420;
  assign n5820 = n86 & ~n1637;
  assign n5821 = ~n1448 & n4615;
  assign n5822 = ~n5818 & ~n5820;
  assign n5823 = ~n5821 & n5822;
  assign n5824 = ~n5819 & n5823;
  assign n5825 = pi26  & n5824;
  assign n5826 = ~pi26  & ~n5824;
  assign n5827 = ~n5825 & ~n5826;
  assign n5828 = ~n5817 & ~n5827;
  assign n5829 = ~n5816 & ~n5828;
  assign n5830 = n5453 & ~n5829;
  assign n5831 = ~n5453 & n5829;
  assign n5832 = ~n1104 & n5109;
  assign n5833 = n3775 & n5045;
  assign n5834 = ~n1225 & n5044;
  assign n5835 = ~n878 & n5130;
  assign n5836 = ~n5832 & ~n5834;
  assign n5837 = ~n5835 & n5836;
  assign n5838 = ~n5833 & n5837;
  assign n5839 = pi23  & n5838;
  assign n5840 = ~pi23  & ~n5838;
  assign n5841 = ~n5839 & ~n5840;
  assign n5842 = ~n5831 & ~n5841;
  assign n5843 = ~n5830 & ~n5842;
  assign n5844 = ~n5449 & ~n5843;
  assign n5845 = ~n5446 & ~n5844;
  assign n5846 = ~n5405 & ~n5406;
  assign n5847 = ~n5416 & n5846;
  assign n5848 = n5416 & ~n5846;
  assign n5849 = ~n5847 & ~n5848;
  assign n5850 = ~n5845 & n5849;
  assign n5851 = n5845 & ~n5849;
  assign n5852 = ~n3855 & n5240;
  assign n5853 = n5235 & ~n5238;
  assign n5854 = ~n3883 & n5853;
  assign n5855 = ~n3900 & n5241;
  assign n5856 = ~n5852 & ~n5854;
  assign n5857 = ~n5855 & n5856;
  assign n5858 = pi20  & n5857;
  assign n5859 = ~pi20  & ~n5857;
  assign n5860 = ~n5858 & ~n5859;
  assign n5861 = ~n5851 & ~n5860;
  assign n5862 = ~n5850 & ~n5861;
  assign n5863 = n5433 & ~n5862;
  assign n5864 = ~n5433 & n5862;
  assign n5865 = ~n5863 & ~n5864;
  assign n5866 = n5232 & ~n5235;
  assign n5867 = ~n3883 & n5866;
  assign n5868 = n4399 & n5241;
  assign n5869 = ~n3855 & n5853;
  assign n5870 = ~n3681 & n5240;
  assign n5871 = ~n5867 & ~n5869;
  assign n5872 = ~n5870 & n5871;
  assign n5873 = ~n5868 & n5872;
  assign n5874 = pi20  & n5873;
  assign n5875 = ~pi20  & ~n5873;
  assign n5876 = ~n5874 & ~n5875;
  assign n5877 = ~n5830 & ~n5831;
  assign n5878 = ~n5841 & n5877;
  assign n5879 = n5841 & ~n5877;
  assign n5880 = ~n5878 & ~n5879;
  assign n5881 = n5471 & n5811;
  assign n5882 = ~n5812 & ~n5881;
  assign n5883 = ~n1637 & n4600;
  assign n5884 = n4420 & n4553;
  assign n5885 = n86 & ~n1717;
  assign n5886 = ~n1533 & n4615;
  assign n5887 = ~n5883 & ~n5885;
  assign n5888 = ~n5886 & n5887;
  assign n5889 = ~n5884 & n5888;
  assign n5890 = pi26  & n5889;
  assign n5891 = ~pi26  & ~n5889;
  assign n5892 = ~n5890 & ~n5891;
  assign n5893 = n5882 & ~n5892;
  assign n5894 = ~n5882 & n5892;
  assign n5895 = ~n5893 & ~n5894;
  assign n5896 = ~n5590 & n5809;
  assign n5897 = ~n5810 & ~n5896;
  assign n5898 = ~n1998 & n3884;
  assign n5899 = n3886 & n5151;
  assign n5900 = ~n2098 & n3810;
  assign n5901 = ~n1908 & n4380;
  assign n5902 = ~n5898 & ~n5900;
  assign n5903 = ~n5901 & n5902;
  assign n5904 = ~n5899 & n5903;
  assign n5905 = pi29  & n5904;
  assign n5906 = ~pi29  & ~n5904;
  assign n5907 = ~n5905 & ~n5906;
  assign n5908 = n5897 & ~n5907;
  assign n5909 = ~n1717 & n4600;
  assign n5910 = n4420 & n4537;
  assign n5911 = n86 & ~n1841;
  assign n5912 = ~n1637 & n4615;
  assign n5913 = ~n5909 & ~n5911;
  assign n5914 = ~n5912 & n5913;
  assign n5915 = ~n5910 & n5914;
  assign n5916 = pi26  & n5915;
  assign n5917 = ~pi26  & ~n5915;
  assign n5918 = ~n5916 & ~n5917;
  assign n5919 = ~n5897 & n5907;
  assign n5920 = ~n5918 & ~n5919;
  assign n5921 = ~n5908 & ~n5920;
  assign n5922 = n5895 & ~n5921;
  assign n5923 = ~n5893 & ~n5922;
  assign n5924 = ~n5816 & ~n5817;
  assign n5925 = ~n5827 & n5924;
  assign n5926 = n5827 & ~n5924;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = ~n5923 & n5927;
  assign n5929 = n5923 & ~n5927;
  assign n5930 = ~n1225 & n5109;
  assign n5931 = n4135 & n5045;
  assign n5932 = ~n1345 & n5044;
  assign n5933 = ~n1104 & n5130;
  assign n5934 = ~n5930 & ~n5932;
  assign n5935 = ~n5933 & n5934;
  assign n5936 = ~n5931 & n5935;
  assign n5937 = pi23  & n5936;
  assign n5938 = ~pi23  & ~n5936;
  assign n5939 = ~n5937 & ~n5938;
  assign n5940 = ~n5929 & ~n5939;
  assign n5941 = ~n5928 & ~n5940;
  assign n5942 = n5880 & ~n5941;
  assign n5943 = ~n5880 & n5941;
  assign n5944 = ~n3855 & n5866;
  assign n5945 = n3972 & n5241;
  assign n5946 = ~n987 & n5240;
  assign n5947 = ~n3681 & n5853;
  assign n5948 = ~n5944 & ~n5946;
  assign n5949 = ~n5947 & n5948;
  assign n5950 = ~n5945 & n5949;
  assign n5951 = pi20  & n5950;
  assign n5952 = ~pi20  & ~n5950;
  assign n5953 = ~n5951 & ~n5952;
  assign n5954 = ~n5943 & ~n5953;
  assign n5955 = ~n5942 & ~n5954;
  assign n5956 = ~n5876 & ~n5955;
  assign n5957 = n5449 & n5843;
  assign n5958 = ~n5844 & ~n5957;
  assign n5959 = n5876 & n5955;
  assign n5960 = ~n5956 & ~n5959;
  assign n5961 = n5958 & n5960;
  assign n5962 = ~n5956 & ~n5961;
  assign n5963 = ~n5850 & ~n5851;
  assign n5964 = ~n5860 & n5963;
  assign n5965 = n5860 & ~n5963;
  assign n5966 = ~n5964 & ~n5965;
  assign n5967 = ~n5962 & n5966;
  assign n5968 = n5962 & ~n5966;
  assign n5969 = ~n5967 & ~n5968;
  assign n5970 = ~n5958 & ~n5960;
  assign n5971 = ~n5961 & ~n5970;
  assign n5972 = pi16  & ~pi17 ;
  assign n5973 = ~pi16  & pi17 ;
  assign n5974 = ~n5972 & ~n5973;
  assign n5975 = ~pi15  & pi16 ;
  assign n5976 = pi15  & ~pi16 ;
  assign n5977 = ~n5975 & ~n5976;
  assign n5978 = pi14  & ~pi15 ;
  assign n5979 = ~pi14  & pi15 ;
  assign n5980 = ~n5978 & ~n5979;
  assign n5981 = n5977 & n5980;
  assign n5982 = ~n5974 & n5981;
  assign n5983 = ~n5974 & ~n5980;
  assign n5984 = ~n3897 & n5983;
  assign n5985 = ~n5982 & ~n5984;
  assign n5986 = ~n3883 & ~n5985;
  assign n5987 = pi17  & ~n5986;
  assign n5988 = ~pi17  & n5986;
  assign n5989 = ~n5987 & ~n5988;
  assign n5990 = ~n1345 & n5109;
  assign n5991 = n4152 & n5045;
  assign n5992 = ~n1448 & n5044;
  assign n5993 = ~n1225 & n5130;
  assign n5994 = ~n5990 & ~n5992;
  assign n5995 = ~n5993 & n5994;
  assign n5996 = ~n5991 & n5995;
  assign n5997 = ~pi23  & ~n5996;
  assign n5998 = pi23  & n5996;
  assign n5999 = ~n5997 & ~n5998;
  assign n6000 = ~n5895 & n5921;
  assign n6001 = ~n5922 & ~n6000;
  assign n6002 = ~n5999 & n6001;
  assign n6003 = ~n5999 & ~n6001;
  assign n6004 = n5999 & n6001;
  assign n6005 = ~n6003 & ~n6004;
  assign n6006 = ~n5908 & ~n5919;
  assign n6007 = n5918 & ~n6006;
  assign n6008 = ~n5918 & n6006;
  assign n6009 = ~n6007 & ~n6008;
  assign n6010 = ~n5797 & n5807;
  assign n6011 = ~n5808 & ~n6010;
  assign n6012 = ~n5630 & n5784;
  assign n6013 = ~n5785 & ~n6012;
  assign n6014 = n748 & ~n2589;
  assign n6015 = n3536 & ~n3538;
  assign n6016 = ~n3539 & ~n6015;
  assign n6017 = n880 & n6016;
  assign n6018 = ~n2496 & n3692;
  assign n6019 = ~n2412 & n3694;
  assign n6020 = ~n6014 & ~n6018;
  assign n6021 = ~n6019 & n6020;
  assign n6022 = ~n6017 & n6021;
  assign n6023 = n6013 & ~n6022;
  assign n6024 = ~n2146 & n4380;
  assign n6025 = n3886 & n5343;
  assign n6026 = ~n2347 & n3810;
  assign n6027 = ~n2249 & n3884;
  assign n6028 = ~n6024 & ~n6026;
  assign n6029 = ~n6027 & n6028;
  assign n6030 = ~n6025 & n6029;
  assign n6031 = ~pi29  & ~n6030;
  assign n6032 = pi29  & n6030;
  assign n6033 = ~n6031 & ~n6032;
  assign n6034 = n6013 & n6022;
  assign n6035 = ~n6013 & ~n6022;
  assign n6036 = ~n6034 & ~n6035;
  assign n6037 = ~n6033 & ~n6036;
  assign n6038 = ~n6023 & ~n6037;
  assign n6039 = n5786 & ~n5788;
  assign n6040 = ~n5789 & ~n6039;
  assign n6041 = ~n6038 & n6040;
  assign n6042 = ~n2098 & n4380;
  assign n6043 = n3886 & n5359;
  assign n6044 = ~n2146 & n3884;
  assign n6045 = ~n2249 & n3810;
  assign n6046 = ~n6042 & ~n6044;
  assign n6047 = ~n6045 & n6046;
  assign n6048 = ~n6043 & n6047;
  assign n6049 = pi29  & n6048;
  assign n6050 = ~pi29  & ~n6048;
  assign n6051 = ~n6049 & ~n6050;
  assign n6052 = n6038 & ~n6040;
  assign n6053 = ~n6051 & ~n6052;
  assign n6054 = ~n6041 & ~n6053;
  assign n6055 = n6011 & ~n6054;
  assign n6056 = ~n6011 & n6054;
  assign n6057 = ~n1841 & n4600;
  assign n6058 = n4420 & n4762;
  assign n6059 = n86 & ~n1908;
  assign n6060 = ~n1717 & n4615;
  assign n6061 = ~n6057 & ~n6059;
  assign n6062 = ~n6060 & n6061;
  assign n6063 = ~n6058 & n6062;
  assign n6064 = pi26  & n6063;
  assign n6065 = ~pi26  & ~n6063;
  assign n6066 = ~n6064 & ~n6065;
  assign n6067 = ~n6056 & ~n6066;
  assign n6068 = ~n6055 & ~n6067;
  assign n6069 = n6009 & ~n6068;
  assign n6070 = ~n6009 & n6068;
  assign n6071 = ~n1448 & n5109;
  assign n6072 = n4453 & n5045;
  assign n6073 = ~n1533 & n5044;
  assign n6074 = ~n1345 & n5130;
  assign n6075 = ~n6071 & ~n6073;
  assign n6076 = ~n6074 & n6075;
  assign n6077 = ~n6072 & n6076;
  assign n6078 = pi23  & n6077;
  assign n6079 = ~pi23  & ~n6077;
  assign n6080 = ~n6078 & ~n6079;
  assign n6081 = ~n6070 & ~n6080;
  assign n6082 = ~n6069 & ~n6081;
  assign n6083 = ~n6005 & ~n6082;
  assign n6084 = ~n6002 & ~n6083;
  assign n6085 = ~n5928 & ~n5929;
  assign n6086 = ~n5939 & n6085;
  assign n6087 = n5939 & ~n6085;
  assign n6088 = ~n6086 & ~n6087;
  assign n6089 = ~n6084 & n6088;
  assign n6090 = n6084 & ~n6088;
  assign n6091 = ~n878 & n5240;
  assign n6092 = n3687 & n5241;
  assign n6093 = ~n987 & n5853;
  assign n6094 = ~n3681 & n5866;
  assign n6095 = ~n6091 & ~n6093;
  assign n6096 = ~n6094 & n6095;
  assign n6097 = ~n6092 & n6096;
  assign n6098 = pi20  & n6097;
  assign n6099 = ~pi20  & ~n6097;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = ~n6090 & ~n6100;
  assign n6102 = ~n6089 & ~n6101;
  assign n6103 = ~n5989 & ~n6102;
  assign n6104 = n5989 & n6102;
  assign n6105 = ~n5942 & ~n5943;
  assign n6106 = ~n5953 & n6105;
  assign n6107 = n5953 & ~n6105;
  assign n6108 = ~n6106 & ~n6107;
  assign n6109 = ~n6104 & n6108;
  assign n6110 = ~n6103 & ~n6109;
  assign n6111 = n5971 & ~n6110;
  assign n6112 = ~n6103 & ~n6104;
  assign n6113 = n6108 & n6112;
  assign n6114 = ~n6108 & ~n6112;
  assign n6115 = ~n6113 & ~n6114;
  assign n6116 = n6005 & n6082;
  assign n6117 = ~n6083 & ~n6116;
  assign n6118 = ~n987 & n5866;
  assign n6119 = n3791 & n5241;
  assign n6120 = ~n1104 & n5240;
  assign n6121 = ~n878 & n5853;
  assign n6122 = ~n6118 & ~n6120;
  assign n6123 = ~n6121 & n6122;
  assign n6124 = ~n6119 & n6123;
  assign n6125 = pi20  & n6124;
  assign n6126 = ~pi20  & ~n6124;
  assign n6127 = ~n6125 & ~n6126;
  assign n6128 = n6117 & ~n6127;
  assign n6129 = ~n6117 & n6127;
  assign n6130 = ~n6128 & ~n6129;
  assign n6131 = ~n6069 & ~n6070;
  assign n6132 = ~n6080 & n6131;
  assign n6133 = n6080 & ~n6131;
  assign n6134 = ~n6132 & ~n6133;
  assign n6135 = ~n1908 & n4600;
  assign n6136 = n4420 & n4779;
  assign n6137 = n86 & ~n1998;
  assign n6138 = ~n1841 & n4615;
  assign n6139 = ~n6135 & ~n6137;
  assign n6140 = ~n6138 & n6139;
  assign n6141 = ~n6136 & n6140;
  assign n6142 = pi26  & n6141;
  assign n6143 = ~pi26  & ~n6141;
  assign n6144 = ~n6142 & ~n6143;
  assign n6145 = ~n6041 & ~n6052;
  assign n6146 = n6051 & ~n6145;
  assign n6147 = ~n6051 & n6145;
  assign n6148 = ~n6146 & ~n6147;
  assign n6149 = ~n6144 & n6148;
  assign n6150 = n6144 & ~n6148;
  assign n6151 = ~n6149 & ~n6150;
  assign n6152 = ~n5772 & ~n5773;
  assign n6153 = ~n5782 & n6152;
  assign n6154 = n5782 & ~n6152;
  assign n6155 = ~n6153 & ~n6154;
  assign n6156 = ~n634 & n1272;
  assign n6157 = n1357 & n6156;
  assign n6158 = ~n159 & ~n355;
  assign n6159 = ~n698 & ~n751;
  assign n6160 = n6158 & n6159;
  assign n6161 = n1947 & n2283;
  assign n6162 = n2473 & n4269;
  assign n6163 = n5720 & n6162;
  assign n6164 = n6160 & n6161;
  assign n6165 = n1132 & n3996;
  assign n6166 = n6164 & n6165;
  assign n6167 = n6157 & n6163;
  assign n6168 = n6166 & n6167;
  assign n6169 = ~n310 & ~n312;
  assign n6170 = ~n1034 & n6169;
  assign n6171 = ~n183 & ~n661;
  assign n6172 = ~n186 & ~n246;
  assign n6173 = ~n352 & ~n373;
  assign n6174 = ~n532 & ~n787;
  assign n6175 = n6173 & n6174;
  assign n6176 = n940 & n6172;
  assign n6177 = n1243 & n1470;
  assign n6178 = n1673 & n6171;
  assign n6179 = n6177 & n6178;
  assign n6180 = n6175 & n6176;
  assign n6181 = n6170 & n6180;
  assign n6182 = n5717 & n6179;
  assign n6183 = n6181 & n6182;
  assign n6184 = n5691 & n6183;
  assign n6185 = n1738 & n6168;
  assign n6186 = n6184 & n6185;
  assign n6187 = n4324 & n6186;
  assign n6188 = n5704 & ~n6187;
  assign n6189 = ~n5704 & n6187;
  assign n6190 = ~n6188 & ~n6189;
  assign n6191 = ~n162 & ~n476;
  assign n6192 = ~n522 & n6191;
  assign n6193 = n1271 & n2358;
  assign n6194 = n2399 & n6193;
  assign n6195 = n6192 & n6194;
  assign n6196 = ~n111 & ~n687;
  assign n6197 = ~n196 & ~n446;
  assign n6198 = ~n515 & ~n523;
  assign n6199 = ~n638 & n6198;
  assign n6200 = n428 & n6197;
  assign n6201 = n431 & n3705;
  assign n6202 = n6196 & n6201;
  assign n6203 = n6199 & n6200;
  assign n6204 = n1700 & n3733;
  assign n6205 = n6203 & n6204;
  assign n6206 = n1433 & n6202;
  assign n6207 = n6205 & n6206;
  assign n6208 = n1402 & n6195;
  assign n6209 = n6207 & n6208;
  assign n6210 = n351 & n6209;
  assign n6211 = n4954 & n6210;
  assign n6212 = ~pi2  & ~n6211;
  assign n6213 = pi2  & ~n6211;
  assign n6214 = ~pi2  & n6211;
  assign n6215 = ~n6213 & ~n6214;
  assign n6216 = ~pi5  & ~n6215;
  assign n6217 = ~n6212 & ~n6216;
  assign n6218 = n5704 & ~n6217;
  assign n6219 = ~n5704 & n6217;
  assign n6220 = ~n2708 & n3694;
  assign n6221 = n3520 & ~n3522;
  assign n6222 = ~n3523 & ~n6221;
  assign n6223 = n880 & n6222;
  assign n6224 = n748 & ~n2835;
  assign n6225 = ~n2778 & n3692;
  assign n6226 = ~n6220 & ~n6224;
  assign n6227 = ~n6225 & n6226;
  assign n6228 = ~n6223 & n6227;
  assign n6229 = ~n6219 & ~n6228;
  assign n6230 = ~n6218 & ~n6229;
  assign n6231 = n6190 & ~n6230;
  assign n6232 = ~n6188 & ~n6231;
  assign n6233 = ~pi8  & ~n5770;
  assign n6234 = ~n5768 & n5771;
  assign n6235 = ~n6233 & ~n6234;
  assign n6236 = ~n6232 & ~n6235;
  assign n6237 = n6232 & n6235;
  assign n6238 = ~n2674 & n3692;
  assign n6239 = n3528 & ~n3530;
  assign n6240 = ~n3531 & ~n6239;
  assign n6241 = n880 & n6240;
  assign n6242 = n748 & ~n2708;
  assign n6243 = ~n2589 & n3694;
  assign n6244 = ~n6238 & ~n6242;
  assign n6245 = ~n6243 & n6244;
  assign n6246 = ~n6241 & n6245;
  assign n6247 = ~n6237 & ~n6246;
  assign n6248 = ~n6236 & ~n6247;
  assign n6249 = n6155 & ~n6248;
  assign n6250 = ~n6155 & n6248;
  assign n6251 = ~n6249 & ~n6250;
  assign n6252 = ~n2412 & n3810;
  assign n6253 = n3886 & n5579;
  assign n6254 = ~n2347 & n3884;
  assign n6255 = ~n2249 & n4380;
  assign n6256 = ~n6252 & ~n6254;
  assign n6257 = ~n6255 & n6256;
  assign n6258 = ~n6253 & n6257;
  assign n6259 = pi29  & n6258;
  assign n6260 = ~pi29  & ~n6258;
  assign n6261 = ~n6259 & ~n6260;
  assign n6262 = n6251 & ~n6261;
  assign n6263 = ~n6249 & ~n6262;
  assign n6264 = n6033 & n6036;
  assign n6265 = ~n6037 & ~n6264;
  assign n6266 = ~n6263 & n6265;
  assign n6267 = n6263 & ~n6265;
  assign n6268 = ~n1998 & n4600;
  assign n6269 = n4420 & n5151;
  assign n6270 = n86 & ~n2098;
  assign n6271 = ~n1908 & n4615;
  assign n6272 = ~n6268 & ~n6270;
  assign n6273 = ~n6271 & n6272;
  assign n6274 = ~n6269 & n6273;
  assign n6275 = pi26  & n6274;
  assign n6276 = ~pi26  & ~n6274;
  assign n6277 = ~n6275 & ~n6276;
  assign n6278 = ~n6267 & ~n6277;
  assign n6279 = ~n6266 & ~n6278;
  assign n6280 = n6151 & ~n6279;
  assign n6281 = ~n6149 & ~n6280;
  assign n6282 = ~n6055 & ~n6056;
  assign n6283 = ~n6066 & n6282;
  assign n6284 = n6066 & ~n6282;
  assign n6285 = ~n6283 & ~n6284;
  assign n6286 = ~n6281 & n6285;
  assign n6287 = n6281 & ~n6285;
  assign n6288 = ~n1533 & n5109;
  assign n6289 = n4355 & n5045;
  assign n6290 = ~n1637 & n5044;
  assign n6291 = ~n1448 & n5130;
  assign n6292 = ~n6288 & ~n6290;
  assign n6293 = ~n6291 & n6292;
  assign n6294 = ~n6289 & n6293;
  assign n6295 = pi23  & n6294;
  assign n6296 = ~pi23  & ~n6294;
  assign n6297 = ~n6295 & ~n6296;
  assign n6298 = ~n6287 & ~n6297;
  assign n6299 = ~n6286 & ~n6298;
  assign n6300 = n6134 & ~n6299;
  assign n6301 = ~n6134 & n6299;
  assign n6302 = ~n1104 & n5853;
  assign n6303 = n3775 & n5241;
  assign n6304 = ~n1225 & n5240;
  assign n6305 = ~n878 & n5866;
  assign n6306 = ~n6302 & ~n6304;
  assign n6307 = ~n6305 & n6306;
  assign n6308 = ~n6303 & n6307;
  assign n6309 = pi20  & n6308;
  assign n6310 = ~pi20  & ~n6308;
  assign n6311 = ~n6309 & ~n6310;
  assign n6312 = ~n6301 & ~n6311;
  assign n6313 = ~n6300 & ~n6312;
  assign n6314 = n6130 & ~n6313;
  assign n6315 = ~n6128 & ~n6314;
  assign n6316 = ~n6089 & ~n6090;
  assign n6317 = ~n6100 & n6316;
  assign n6318 = n6100 & ~n6316;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = ~n6315 & n6319;
  assign n6321 = n6315 & ~n6319;
  assign n6322 = ~n3855 & n5982;
  assign n6323 = ~n5977 & n5980;
  assign n6324 = ~n3883 & n6323;
  assign n6325 = ~n3900 & n5983;
  assign n6326 = ~n6322 & ~n6324;
  assign n6327 = ~n6325 & n6326;
  assign n6328 = pi17  & n6327;
  assign n6329 = ~pi17  & ~n6327;
  assign n6330 = ~n6328 & ~n6329;
  assign n6331 = ~n6321 & ~n6330;
  assign n6332 = ~n6320 & ~n6331;
  assign n6333 = n6115 & ~n6332;
  assign n6334 = ~n6115 & n6332;
  assign n6335 = ~n6333 & ~n6334;
  assign n6336 = n5974 & ~n5980;
  assign n6337 = ~n3883 & n6336;
  assign n6338 = n4399 & n5983;
  assign n6339 = ~n3855 & n6323;
  assign n6340 = ~n3681 & n5982;
  assign n6341 = ~n6337 & ~n6339;
  assign n6342 = ~n6340 & n6341;
  assign n6343 = ~n6338 & n6342;
  assign n6344 = pi17  & n6343;
  assign n6345 = ~pi17  & ~n6343;
  assign n6346 = ~n6344 & ~n6345;
  assign n6347 = ~n6300 & ~n6301;
  assign n6348 = ~n6311 & n6347;
  assign n6349 = n6311 & ~n6347;
  assign n6350 = ~n6348 & ~n6349;
  assign n6351 = ~n1637 & n5109;
  assign n6352 = n4553 & n5045;
  assign n6353 = ~n1717 & n5044;
  assign n6354 = ~n1533 & n5130;
  assign n6355 = ~n6351 & ~n6353;
  assign n6356 = ~n6354 & n6355;
  assign n6357 = ~n6352 & n6356;
  assign n6358 = ~pi23  & ~n6357;
  assign n6359 = pi23  & n6357;
  assign n6360 = ~n6358 & ~n6359;
  assign n6361 = ~n6151 & n6279;
  assign n6362 = ~n6280 & ~n6361;
  assign n6363 = ~n6360 & n6362;
  assign n6364 = ~n6360 & ~n6362;
  assign n6365 = n6360 & n6362;
  assign n6366 = ~n6364 & ~n6365;
  assign n6367 = ~n6266 & ~n6267;
  assign n6368 = ~n6277 & n6367;
  assign n6369 = n6277 & ~n6367;
  assign n6370 = ~n6368 & ~n6369;
  assign n6371 = ~n2347 & n4380;
  assign n6372 = n3886 & n5596;
  assign n6373 = ~n2496 & n3810;
  assign n6374 = ~n2412 & n3884;
  assign n6375 = ~n6371 & ~n6373;
  assign n6376 = ~n6374 & n6375;
  assign n6377 = ~n6372 & n6376;
  assign n6378 = ~pi29  & ~n6377;
  assign n6379 = pi29  & n6377;
  assign n6380 = ~n6378 & ~n6379;
  assign n6381 = ~n6236 & ~n6237;
  assign n6382 = ~n6246 & n6381;
  assign n6383 = n6246 & ~n6381;
  assign n6384 = ~n6382 & ~n6383;
  assign n6385 = ~n6380 & n6384;
  assign n6386 = ~n6380 & ~n6384;
  assign n6387 = n6380 & n6384;
  assign n6388 = ~n6386 & ~n6387;
  assign n6389 = ~n6190 & n6230;
  assign n6390 = ~n6231 & ~n6389;
  assign n6391 = n748 & ~n2778;
  assign n6392 = n3524 & ~n3526;
  assign n6393 = ~n3527 & ~n6392;
  assign n6394 = n880 & n6393;
  assign n6395 = ~n2708 & n3692;
  assign n6396 = ~n2674 & n3694;
  assign n6397 = ~n6391 & ~n6395;
  assign n6398 = ~n6396 & n6397;
  assign n6399 = ~n6394 & n6398;
  assign n6400 = n6390 & ~n6399;
  assign n6401 = ~n6218 & ~n6219;
  assign n6402 = ~n6228 & n6401;
  assign n6403 = n6228 & ~n6401;
  assign n6404 = ~n6402 & ~n6403;
  assign n6405 = ~n235 & ~n255;
  assign n6406 = ~n902 & n6405;
  assign n6407 = n788 & n917;
  assign n6408 = n1120 & n3460;
  assign n6409 = n6407 & n6408;
  assign n6410 = n6406 & n6409;
  assign n6411 = ~n327 & ~n377;
  assign n6412 = ~n1034 & n6411;
  assign n6413 = n1081 & n2839;
  assign n6414 = n6412 & n6413;
  assign n6415 = ~n196 & ~n313;
  assign n6416 = n360 & n6415;
  assign n6417 = n1650 & n3744;
  assign n6418 = n4857 & n6417;
  assign n6419 = n1279 & n6416;
  assign n6420 = n5526 & n5611;
  assign n6421 = n6419 & n6420;
  assign n6422 = n2061 & n6418;
  assign n6423 = n6414 & n6422;
  assign n6424 = n6410 & n6421;
  assign n6425 = n6423 & n6424;
  assign n6426 = n1185 & n6425;
  assign n6427 = n2888 & n3147;
  assign n6428 = n6426 & n6427;
  assign n6429 = pi2  & ~n6428;
  assign n6430 = ~n116 & ~n414;
  assign n6431 = n1650 & n1669;
  assign n6432 = n4004 & n6431;
  assign n6433 = ~n143 & ~n171;
  assign n6434 = ~n212 & ~n523;
  assign n6435 = n6433 & n6434;
  assign n6436 = n1296 & n1424;
  assign n6437 = n2258 & n5299;
  assign n6438 = n6430 & n6437;
  assign n6439 = n6435 & n6436;
  assign n6440 = n1152 & n4494;
  assign n6441 = n6439 & n6440;
  assign n6442 = n1361 & n6438;
  assign n6443 = n4863 & n6432;
  assign n6444 = n6442 & n6443;
  assign n6445 = n268 & n6441;
  assign n6446 = n6444 & n6445;
  assign n6447 = n1507 & n6446;
  assign n6448 = n3341 & n6447;
  assign n6449 = pi2  & ~n6448;
  assign n6450 = ~n276 & ~n284;
  assign n6451 = ~n296 & ~n300;
  assign n6452 = ~n596 & n6451;
  assign n6453 = n527 & n6450;
  assign n6454 = n1245 & n1424;
  assign n6455 = n1913 & n2279;
  assign n6456 = n6454 & n6455;
  assign n6457 = n6452 & n6453;
  assign n6458 = n1279 & n3310;
  assign n6459 = n5609 & n6458;
  assign n6460 = n6456 & n6457;
  assign n6461 = n5649 & n6460;
  assign n6462 = n6459 & n6461;
  assign n6463 = ~n259 & ~n656;
  assign n6464 = ~n753 & ~n768;
  assign n6465 = ~n839 & n6464;
  assign n6466 = n137 & n6463;
  assign n6467 = n6465 & n6466;
  assign n6468 = ~n126 & ~n237;
  assign n6469 = n360 & n6468;
  assign n6470 = n1475 & n2978;
  assign n6471 = n3409 & n4858;
  assign n6472 = n5269 & n6471;
  assign n6473 = n6469 & n6470;
  assign n6474 = n507 & n6473;
  assign n6475 = n6467 & n6472;
  assign n6476 = n6474 & n6475;
  assign n6477 = n457 & n546;
  assign n6478 = n6476 & n6477;
  assign n6479 = n6462 & n6478;
  assign n6480 = n2233 & n6479;
  assign n6481 = pi2  & ~n6480;
  assign n6482 = ~pi2  & n6480;
  assign n6483 = ~n6481 & ~n6482;
  assign n6484 = ~n2951 & n3694;
  assign n6485 = n3504 & ~n3506;
  assign n6486 = ~n3507 & ~n6485;
  assign n6487 = n880 & n6486;
  assign n6488 = n748 & ~n3118;
  assign n6489 = ~n3031 & n3692;
  assign n6490 = ~n6484 & ~n6488;
  assign n6491 = ~n6489 & n6490;
  assign n6492 = ~n6487 & n6491;
  assign n6493 = n6483 & ~n6492;
  assign n6494 = ~n6481 & ~n6493;
  assign n6495 = ~pi2  & n6448;
  assign n6496 = ~n6449 & ~n6495;
  assign n6497 = ~n6494 & n6496;
  assign n6498 = ~n6449 & ~n6497;
  assign n6499 = ~pi2  & n6428;
  assign n6500 = ~n6429 & ~n6499;
  assign n6501 = ~n6498 & n6500;
  assign n6502 = ~n6429 & ~n6501;
  assign n6503 = pi5  & n6215;
  assign n6504 = ~n6216 & ~n6503;
  assign n6505 = ~n6502 & n6504;
  assign n6506 = n6502 & ~n6504;
  assign n6507 = n748 & ~n2919;
  assign n6508 = n3516 & ~n3518;
  assign n6509 = ~n3519 & ~n6508;
  assign n6510 = n880 & n6509;
  assign n6511 = ~n2835 & n3692;
  assign n6512 = ~n2778 & n3694;
  assign n6513 = ~n6507 & ~n6511;
  assign n6514 = ~n6512 & n6513;
  assign n6515 = ~n6510 & n6514;
  assign n6516 = ~n6506 & ~n6515;
  assign n6517 = ~n6505 & ~n6516;
  assign n6518 = n6404 & ~n6517;
  assign n6519 = ~n6404 & n6517;
  assign n6520 = ~n6518 & ~n6519;
  assign n6521 = ~n2496 & n4380;
  assign n6522 = n3886 & n5776;
  assign n6523 = ~n2674 & n3810;
  assign n6524 = ~n2589 & n3884;
  assign n6525 = ~n6521 & ~n6523;
  assign n6526 = ~n6524 & n6525;
  assign n6527 = ~n6522 & n6526;
  assign n6528 = pi29  & n6527;
  assign n6529 = ~pi29  & ~n6527;
  assign n6530 = ~n6528 & ~n6529;
  assign n6531 = n6520 & ~n6530;
  assign n6532 = ~n6518 & ~n6531;
  assign n6533 = n6390 & n6399;
  assign n6534 = ~n6390 & ~n6399;
  assign n6535 = ~n6533 & ~n6534;
  assign n6536 = ~n6532 & ~n6535;
  assign n6537 = ~n6400 & ~n6536;
  assign n6538 = ~n6388 & ~n6537;
  assign n6539 = ~n6385 & ~n6538;
  assign n6540 = ~n6251 & n6261;
  assign n6541 = ~n6262 & ~n6540;
  assign n6542 = ~n6539 & n6541;
  assign n6543 = n6539 & ~n6541;
  assign n6544 = ~n2098 & n4600;
  assign n6545 = n4420 & n4979;
  assign n6546 = n86 & ~n2146;
  assign n6547 = ~n1998 & n4615;
  assign n6548 = ~n6544 & ~n6546;
  assign n6549 = ~n6547 & n6548;
  assign n6550 = ~n6545 & n6549;
  assign n6551 = pi26  & n6550;
  assign n6552 = ~pi26  & ~n6550;
  assign n6553 = ~n6551 & ~n6552;
  assign n6554 = ~n6543 & ~n6553;
  assign n6555 = ~n6542 & ~n6554;
  assign n6556 = n6370 & ~n6555;
  assign n6557 = ~n6370 & n6555;
  assign n6558 = ~n1717 & n5109;
  assign n6559 = n4537 & n5045;
  assign n6560 = ~n1841 & n5044;
  assign n6561 = ~n1637 & n5130;
  assign n6562 = ~n6558 & ~n6560;
  assign n6563 = ~n6561 & n6562;
  assign n6564 = ~n6559 & n6563;
  assign n6565 = pi23  & n6564;
  assign n6566 = ~pi23  & ~n6564;
  assign n6567 = ~n6565 & ~n6566;
  assign n6568 = ~n6557 & ~n6567;
  assign n6569 = ~n6556 & ~n6568;
  assign n6570 = ~n6366 & ~n6569;
  assign n6571 = ~n6363 & ~n6570;
  assign n6572 = ~n6286 & ~n6287;
  assign n6573 = ~n6297 & n6572;
  assign n6574 = n6297 & ~n6572;
  assign n6575 = ~n6573 & ~n6574;
  assign n6576 = ~n6571 & n6575;
  assign n6577 = n6571 & ~n6575;
  assign n6578 = ~n1225 & n5853;
  assign n6579 = n4135 & n5241;
  assign n6580 = ~n1345 & n5240;
  assign n6581 = ~n1104 & n5866;
  assign n6582 = ~n6578 & ~n6580;
  assign n6583 = ~n6581 & n6582;
  assign n6584 = ~n6579 & n6583;
  assign n6585 = pi20  & n6584;
  assign n6586 = ~pi20  & ~n6584;
  assign n6587 = ~n6585 & ~n6586;
  assign n6588 = ~n6577 & ~n6587;
  assign n6589 = ~n6576 & ~n6588;
  assign n6590 = n6350 & ~n6589;
  assign n6591 = ~n6350 & n6589;
  assign n6592 = ~n3855 & n6336;
  assign n6593 = n3972 & n5983;
  assign n6594 = ~n987 & n5982;
  assign n6595 = ~n3681 & n6323;
  assign n6596 = ~n6592 & ~n6594;
  assign n6597 = ~n6595 & n6596;
  assign n6598 = ~n6593 & n6597;
  assign n6599 = pi17  & n6598;
  assign n6600 = ~pi17  & ~n6598;
  assign n6601 = ~n6599 & ~n6600;
  assign n6602 = ~n6591 & ~n6601;
  assign n6603 = ~n6590 & ~n6602;
  assign n6604 = ~n6346 & ~n6603;
  assign n6605 = n6346 & n6603;
  assign n6606 = ~n6604 & ~n6605;
  assign n6607 = ~n6130 & n6313;
  assign n6608 = ~n6314 & ~n6607;
  assign n6609 = n6606 & n6608;
  assign n6610 = ~n6604 & ~n6609;
  assign n6611 = ~n6320 & ~n6321;
  assign n6612 = ~n6330 & n6611;
  assign n6613 = n6330 & ~n6611;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = ~n6610 & n6614;
  assign n6616 = n6610 & ~n6614;
  assign n6617 = ~n6615 & ~n6616;
  assign n6618 = ~n6606 & ~n6608;
  assign n6619 = ~n6609 & ~n6618;
  assign n6620 = pi13  & ~pi14 ;
  assign n6621 = ~pi13  & pi14 ;
  assign n6622 = ~n6620 & ~n6621;
  assign n6623 = ~pi12  & pi13 ;
  assign n6624 = pi12  & ~pi13 ;
  assign n6625 = ~n6623 & ~n6624;
  assign n6626 = pi11  & ~pi12 ;
  assign n6627 = ~pi11  & pi12 ;
  assign n6628 = ~n6626 & ~n6627;
  assign n6629 = n6625 & n6628;
  assign n6630 = ~n6622 & n6629;
  assign n6631 = ~n6622 & ~n6628;
  assign n6632 = ~n3897 & n6631;
  assign n6633 = ~n6630 & ~n6632;
  assign n6634 = ~n3883 & ~n6633;
  assign n6635 = pi14  & ~n6634;
  assign n6636 = ~pi14  & n6634;
  assign n6637 = ~n6635 & ~n6636;
  assign n6638 = n6366 & n6569;
  assign n6639 = ~n6570 & ~n6638;
  assign n6640 = ~n1345 & n5853;
  assign n6641 = n4152 & n5241;
  assign n6642 = ~n1448 & n5240;
  assign n6643 = ~n1225 & n5866;
  assign n6644 = ~n6640 & ~n6642;
  assign n6645 = ~n6643 & n6644;
  assign n6646 = ~n6641 & n6645;
  assign n6647 = pi20  & n6646;
  assign n6648 = ~pi20  & ~n6646;
  assign n6649 = ~n6647 & ~n6648;
  assign n6650 = n6639 & ~n6649;
  assign n6651 = ~n6639 & n6649;
  assign n6652 = ~n6650 & ~n6651;
  assign n6653 = ~n6556 & ~n6557;
  assign n6654 = ~n6567 & n6653;
  assign n6655 = n6567 & ~n6653;
  assign n6656 = ~n6654 & ~n6655;
  assign n6657 = n6388 & n6537;
  assign n6658 = ~n6538 & ~n6657;
  assign n6659 = ~n2098 & n4615;
  assign n6660 = n4420 & n5359;
  assign n6661 = ~n2146 & n4600;
  assign n6662 = n86 & ~n2249;
  assign n6663 = ~n6659 & ~n6661;
  assign n6664 = ~n6662 & n6663;
  assign n6665 = ~n6660 & n6664;
  assign n6666 = pi26  & n6665;
  assign n6667 = ~pi26  & ~n6665;
  assign n6668 = ~n6666 & ~n6667;
  assign n6669 = n6658 & ~n6668;
  assign n6670 = ~n6658 & n6668;
  assign n6671 = ~n6669 & ~n6670;
  assign n6672 = ~n2589 & n3810;
  assign n6673 = n3886 & n6016;
  assign n6674 = ~n2496 & n3884;
  assign n6675 = ~n2412 & n4380;
  assign n6676 = ~n6672 & ~n6674;
  assign n6677 = ~n6675 & n6676;
  assign n6678 = ~n6673 & n6677;
  assign n6679 = pi29  & n6678;
  assign n6680 = ~pi29  & ~n6678;
  assign n6681 = ~n6679 & ~n6680;
  assign n6682 = n6532 & n6535;
  assign n6683 = ~n6536 & ~n6682;
  assign n6684 = ~n6681 & n6683;
  assign n6685 = n6681 & ~n6683;
  assign n6686 = ~n2146 & n4615;
  assign n6687 = n4420 & n5343;
  assign n6688 = n86 & ~n2347;
  assign n6689 = ~n2249 & n4600;
  assign n6690 = ~n6686 & ~n6688;
  assign n6691 = ~n6689 & n6690;
  assign n6692 = ~n6687 & n6691;
  assign n6693 = pi26  & n6692;
  assign n6694 = ~pi26  & ~n6692;
  assign n6695 = ~n6693 & ~n6694;
  assign n6696 = ~n6685 & ~n6695;
  assign n6697 = ~n6684 & ~n6696;
  assign n6698 = n6671 & ~n6697;
  assign n6699 = ~n6669 & ~n6698;
  assign n6700 = ~n6542 & ~n6543;
  assign n6701 = ~n6553 & n6700;
  assign n6702 = n6553 & ~n6700;
  assign n6703 = ~n6701 & ~n6702;
  assign n6704 = ~n6699 & n6703;
  assign n6705 = n6699 & ~n6703;
  assign n6706 = ~n1841 & n5109;
  assign n6707 = n4762 & n5045;
  assign n6708 = ~n1908 & n5044;
  assign n6709 = ~n1717 & n5130;
  assign n6710 = ~n6706 & ~n6708;
  assign n6711 = ~n6709 & n6710;
  assign n6712 = ~n6707 & n6711;
  assign n6713 = pi23  & n6712;
  assign n6714 = ~pi23  & ~n6712;
  assign n6715 = ~n6713 & ~n6714;
  assign n6716 = ~n6705 & ~n6715;
  assign n6717 = ~n6704 & ~n6716;
  assign n6718 = n6656 & ~n6717;
  assign n6719 = ~n6656 & n6717;
  assign n6720 = ~n1448 & n5853;
  assign n6721 = n4453 & n5241;
  assign n6722 = ~n1533 & n5240;
  assign n6723 = ~n1345 & n5866;
  assign n6724 = ~n6720 & ~n6722;
  assign n6725 = ~n6723 & n6724;
  assign n6726 = ~n6721 & n6725;
  assign n6727 = pi20  & n6726;
  assign n6728 = ~pi20  & ~n6726;
  assign n6729 = ~n6727 & ~n6728;
  assign n6730 = ~n6719 & ~n6729;
  assign n6731 = ~n6718 & ~n6730;
  assign n6732 = n6652 & ~n6731;
  assign n6733 = ~n6650 & ~n6732;
  assign n6734 = ~n6576 & ~n6577;
  assign n6735 = ~n6587 & n6734;
  assign n6736 = n6587 & ~n6734;
  assign n6737 = ~n6735 & ~n6736;
  assign n6738 = ~n6733 & n6737;
  assign n6739 = n6733 & ~n6737;
  assign n6740 = ~n878 & n5982;
  assign n6741 = n3687 & n5983;
  assign n6742 = ~n987 & n6323;
  assign n6743 = ~n3681 & n6336;
  assign n6744 = ~n6740 & ~n6742;
  assign n6745 = ~n6743 & n6744;
  assign n6746 = ~n6741 & n6745;
  assign n6747 = pi17  & n6746;
  assign n6748 = ~pi17  & ~n6746;
  assign n6749 = ~n6747 & ~n6748;
  assign n6750 = ~n6739 & ~n6749;
  assign n6751 = ~n6738 & ~n6750;
  assign n6752 = ~n6637 & ~n6751;
  assign n6753 = n6637 & n6751;
  assign n6754 = ~n6590 & ~n6591;
  assign n6755 = ~n6601 & n6754;
  assign n6756 = n6601 & ~n6754;
  assign n6757 = ~n6755 & ~n6756;
  assign n6758 = ~n6753 & n6757;
  assign n6759 = ~n6752 & ~n6758;
  assign n6760 = n6619 & ~n6759;
  assign n6761 = ~n6619 & n6759;
  assign n6762 = ~n6760 & ~n6761;
  assign n6763 = ~n987 & n6336;
  assign n6764 = n3791 & n5983;
  assign n6765 = ~n1104 & n5982;
  assign n6766 = ~n878 & n6323;
  assign n6767 = ~n6763 & ~n6765;
  assign n6768 = ~n6766 & n6767;
  assign n6769 = ~n6764 & n6768;
  assign n6770 = ~pi17  & ~n6769;
  assign n6771 = pi17  & n6769;
  assign n6772 = ~n6770 & ~n6771;
  assign n6773 = ~n6652 & n6731;
  assign n6774 = ~n6732 & ~n6773;
  assign n6775 = ~n6772 & n6774;
  assign n6776 = ~n6772 & ~n6774;
  assign n6777 = n6772 & n6774;
  assign n6778 = ~n6776 & ~n6777;
  assign n6779 = ~n6718 & ~n6719;
  assign n6780 = ~n6729 & n6779;
  assign n6781 = n6729 & ~n6779;
  assign n6782 = ~n6780 & ~n6781;
  assign n6783 = ~n1908 & n5109;
  assign n6784 = n4779 & n5045;
  assign n6785 = ~n1998 & n5044;
  assign n6786 = ~n1841 & n5130;
  assign n6787 = ~n6783 & ~n6785;
  assign n6788 = ~n6786 & n6787;
  assign n6789 = ~n6784 & n6788;
  assign n6790 = ~pi23  & ~n6789;
  assign n6791 = pi23  & n6789;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = ~n6671 & n6697;
  assign n6794 = ~n6698 & ~n6793;
  assign n6795 = ~n6792 & n6794;
  assign n6796 = ~n6792 & ~n6794;
  assign n6797 = n6792 & n6794;
  assign n6798 = ~n6796 & ~n6797;
  assign n6799 = ~n6684 & ~n6685;
  assign n6800 = ~n6695 & n6799;
  assign n6801 = n6695 & ~n6799;
  assign n6802 = ~n6800 & ~n6801;
  assign n6803 = ~n6520 & n6530;
  assign n6804 = ~n6531 & ~n6803;
  assign n6805 = n6498 & ~n6500;
  assign n6806 = ~n6501 & ~n6805;
  assign n6807 = n748 & ~n2951;
  assign n6808 = n3512 & ~n3514;
  assign n6809 = ~n3515 & ~n6808;
  assign n6810 = n880 & n6809;
  assign n6811 = ~n2919 & n3692;
  assign n6812 = ~n2835 & n3694;
  assign n6813 = ~n6807 & ~n6811;
  assign n6814 = ~n6812 & n6813;
  assign n6815 = ~n6810 & n6814;
  assign n6816 = n6806 & ~n6815;
  assign n6817 = n6494 & ~n6496;
  assign n6818 = ~n6497 & ~n6817;
  assign n6819 = ~n2919 & n3694;
  assign n6820 = n3508 & ~n3510;
  assign n6821 = ~n3511 & ~n6820;
  assign n6822 = n880 & n6821;
  assign n6823 = ~n2951 & n3692;
  assign n6824 = n748 & ~n3031;
  assign n6825 = ~n6819 & ~n6823;
  assign n6826 = ~n6824 & n6825;
  assign n6827 = ~n6822 & n6826;
  assign n6828 = n6818 & ~n6827;
  assign n6829 = ~n293 & ~n412;
  assign n6830 = ~n414 & ~n438;
  assign n6831 = ~n458 & n6830;
  assign n6832 = n354 & n6829;
  assign n6833 = n513 & n1380;
  assign n6834 = n1890 & n2007;
  assign n6835 = n3326 & n4926;
  assign n6836 = n5299 & n6835;
  assign n6837 = n6833 & n6834;
  assign n6838 = n6831 & n6832;
  assign n6839 = n6837 & n6838;
  assign n6840 = n4867 & n6836;
  assign n6841 = n6839 & n6840;
  assign n6842 = n2618 & n6841;
  assign n6843 = ~n235 & ~n663;
  assign n6844 = n3663 & n6843;
  assign n6845 = ~n597 & n1391;
  assign n6846 = n5650 & n6845;
  assign n6847 = ~n199 & n519;
  assign n6848 = n1271 & n1424;
  assign n6849 = n1779 & n2561;
  assign n6850 = n2685 & n3255;
  assign n6851 = n6849 & n6850;
  assign n6852 = n6847 & n6848;
  assign n6853 = n316 & n2369;
  assign n6854 = n6844 & n6853;
  assign n6855 = n6851 & n6852;
  assign n6856 = n6846 & n6855;
  assign n6857 = n6854 & n6856;
  assign n6858 = n4942 & n6857;
  assign n6859 = n4920 & n6842;
  assign n6860 = n6858 & n6859;
  assign n6861 = n748 & ~n3182;
  assign n6862 = n3500 & ~n3502;
  assign n6863 = ~n3503 & ~n6862;
  assign n6864 = n880 & n6863;
  assign n6865 = ~n3118 & n3692;
  assign n6866 = ~n3031 & n3694;
  assign n6867 = ~n6861 & ~n6865;
  assign n6868 = ~n6866 & n6867;
  assign n6869 = ~n6864 & n6868;
  assign n6870 = ~n6860 & ~n6869;
  assign n6871 = ~n151 & ~n531;
  assign n6872 = n448 & n6871;
  assign n6873 = ~n216 & ~n364;
  assign n6874 = ~n566 & n6873;
  assign n6875 = ~n196 & ~n502;
  assign n6876 = ~n539 & n6875;
  assign n6877 = n292 & n626;
  assign n6878 = n1270 & n2610;
  assign n6879 = n3325 & n5604;
  assign n6880 = n6878 & n6879;
  assign n6881 = n6876 & n6877;
  assign n6882 = n5496 & n6874;
  assign n6883 = n6881 & n6882;
  assign n6884 = n4714 & n6880;
  assign n6885 = n6883 & n6884;
  assign n6886 = ~n168 & ~n318;
  assign n6887 = n1575 & n6886;
  assign n6888 = n2041 & n6887;
  assign n6889 = ~n329 & ~n383;
  assign n6890 = n505 & n6889;
  assign n6891 = n662 & n701;
  assign n6892 = n755 & n1305;
  assign n6893 = n1578 & n1884;
  assign n6894 = n2502 & n2528;
  assign n6895 = n2561 & n6894;
  assign n6896 = n6892 & n6893;
  assign n6897 = n6890 & n6891;
  assign n6898 = n1046 & n6872;
  assign n6899 = n6897 & n6898;
  assign n6900 = n6895 & n6896;
  assign n6901 = n6888 & n6900;
  assign n6902 = n5533 & n6899;
  assign n6903 = n6901 & n6902;
  assign n6904 = n1469 & n6885;
  assign n6905 = n6903 & n6904;
  assign n6906 = ~n3118 & n3694;
  assign n6907 = n3496 & ~n3498;
  assign n6908 = ~n3499 & ~n6907;
  assign n6909 = n880 & n6908;
  assign n6910 = n748 & ~n3241;
  assign n6911 = ~n3182 & n3692;
  assign n6912 = ~n6906 & ~n6910;
  assign n6913 = ~n6911 & n6912;
  assign n6914 = ~n6909 & n6913;
  assign n6915 = ~n6905 & ~n6914;
  assign n6916 = ~n255 & ~n382;
  assign n6917 = ~n523 & ~n944;
  assign n6918 = ~n1034 & n6917;
  assign n6919 = n292 & n6916;
  assign n6920 = n567 & n664;
  assign n6921 = n6919 & n6920;
  assign n6922 = n1844 & n6918;
  assign n6923 = n6921 & n6922;
  assign n6924 = ~n126 & n941;
  assign n6925 = n3262 & n6924;
  assign n6926 = ~n216 & ~n304;
  assign n6927 = ~n922 & n6926;
  assign n6928 = n785 & n6927;
  assign n6929 = ~n282 & ~n294;
  assign n6930 = ~n356 & ~n373;
  assign n6931 = ~n539 & n6930;
  assign n6932 = n799 & n6929;
  assign n6933 = n1429 & n2283;
  assign n6934 = n2459 & n2690;
  assign n6935 = n6933 & n6934;
  assign n6936 = n6931 & n6932;
  assign n6937 = n2415 & n6936;
  assign n6938 = n5607 & n6935;
  assign n6939 = n6925 & n6928;
  assign n6940 = n6938 & n6939;
  assign n6941 = n6937 & n6940;
  assign n6942 = ~n93 & ~n509;
  assign n6943 = ~n512 & n6942;
  assign n6944 = n2933 & n6943;
  assign n6945 = ~n215 & ~n299;
  assign n6946 = ~n358 & ~n1404;
  assign n6947 = n6945 & n6946;
  assign n6948 = n201 & n1141;
  assign n6949 = n2358 & n6948;
  assign n6950 = n6947 & n6949;
  assign n6951 = n6944 & n6950;
  assign n6952 = n781 & n3054;
  assign n6953 = n6923 & n6952;
  assign n6954 = n6951 & n6953;
  assign n6955 = n5677 & n6941;
  assign n6956 = n6954 & n6955;
  assign n6957 = ~n3241 & n3692;
  assign n6958 = n3492 & ~n3494;
  assign n6959 = ~n3495 & ~n6958;
  assign n6960 = n880 & n6959;
  assign n6961 = n748 & ~n3275;
  assign n6962 = ~n3182 & n3694;
  assign n6963 = ~n6957 & ~n6961;
  assign n6964 = ~n6962 & n6963;
  assign n6965 = ~n6960 & n6964;
  assign n6966 = ~n6956 & ~n6965;
  assign n6967 = ~n98 & ~n319;
  assign n6968 = ~n156 & ~n184;
  assign n6969 = ~n427 & n6968;
  assign n6970 = n647 & n6967;
  assign n6971 = n6969 & n6970;
  assign n6972 = ~n304 & ~n314;
  assign n6973 = ~n518 & ~n594;
  assign n6974 = ~n604 & ~n770;
  assign n6975 = ~n808 & n6974;
  assign n6976 = n6972 & n6973;
  assign n6977 = n146 & n176;
  assign n6978 = n883 & n1187;
  assign n6979 = n6977 & n6978;
  assign n6980 = n6975 & n6976;
  assign n6981 = n4493 & n6980;
  assign n6982 = n6979 & n6981;
  assign n6983 = ~n603 & ~n792;
  assign n6984 = n1296 & n6983;
  assign n6985 = ~n215 & ~n520;
  assign n6986 = ~n638 & ~n715;
  assign n6987 = n6985 & n6986;
  assign n6988 = n164 & n272;
  assign n6989 = n461 & n628;
  assign n6990 = n784 & n933;
  assign n6991 = n2037 & n4858;
  assign n6992 = n6990 & n6991;
  assign n6993 = n6988 & n6989;
  assign n6994 = n2416 & n6987;
  assign n6995 = n4066 & n6984;
  assign n6996 = n6994 & n6995;
  assign n6997 = n6992 & n6993;
  assign n6998 = n6971 & n6997;
  assign n6999 = n6996 & n6998;
  assign n7000 = n6982 & n6999;
  assign n7001 = n3006 & n7000;
  assign n7002 = ~n3241 & n3694;
  assign n7003 = n3488 & ~n3490;
  assign n7004 = ~n3491 & ~n7003;
  assign n7005 = n880 & n7004;
  assign n7006 = ~n3275 & n3692;
  assign n7007 = n748 & ~n3370;
  assign n7008 = ~n7002 & ~n7006;
  assign n7009 = ~n7007 & n7008;
  assign n7010 = ~n7005 & n7009;
  assign n7011 = ~n7001 & ~n7010;
  assign n7012 = ~n7001 & n7010;
  assign n7013 = n7001 & ~n7010;
  assign n7014 = ~n7012 & ~n7013;
  assign n7015 = ~n180 & ~n337;
  assign n7016 = n4022 & n7015;
  assign n7017 = n179 & n1004;
  assign n7018 = ~n148 & ~n246;
  assign n7019 = ~n353 & ~n510;
  assign n7020 = ~n687 & ~n1487;
  assign n7021 = n7019 & n7020;
  assign n7022 = n1052 & n7018;
  assign n7023 = n3459 & n7022;
  assign n7024 = n7021 & n7023;
  assign n7025 = ~n303 & ~n1034;
  assign n7026 = n524 & n7025;
  assign n7027 = n593 & n852;
  assign n7028 = n1270 & n1356;
  assign n7029 = n1538 & n1858;
  assign n7030 = n2534 & n4015;
  assign n7031 = n7029 & n7030;
  assign n7032 = n7027 & n7028;
  assign n7033 = n7017 & n7026;
  assign n7034 = n7032 & n7033;
  assign n7035 = n7016 & n7031;
  assign n7036 = n7034 & n7035;
  assign n7037 = n7024 & n7036;
  assign n7038 = n2901 & n7037;
  assign n7039 = n4081 & n4731;
  assign n7040 = n7038 & n7039;
  assign n7041 = ~n3485 & n3692;
  assign n7042 = n3427 & ~n3485;
  assign n7043 = n3370 & ~n7042;
  assign n7044 = ~n3370 & n7042;
  assign n7045 = ~n7043 & ~n7044;
  assign n7046 = n880 & n7045;
  assign n7047 = n748 & ~n3427;
  assign n7048 = ~n3370 & n3694;
  assign n7049 = ~n7041 & ~n7047;
  assign n7050 = ~n7048 & n7049;
  assign n7051 = ~n7046 & n7050;
  assign n7052 = ~n7040 & ~n7051;
  assign n7053 = ~n213 & ~n303;
  assign n7054 = ~n310 & ~n415;
  assign n7055 = ~n511 & n7054;
  assign n7056 = n1052 & n7053;
  assign n7057 = n7055 & n7056;
  assign n7058 = ~n601 & n2890;
  assign n7059 = ~n237 & ~n561;
  assign n7060 = n1130 & n7059;
  assign n7061 = ~n180 & ~n273;
  assign n7062 = ~n568 & ~n685;
  assign n7063 = n7061 & n7062;
  assign n7064 = n217 & n940;
  assign n7065 = n942 & n7064;
  assign n7066 = n2450 & n7063;
  assign n7067 = n7065 & n7066;
  assign n7068 = ~n253 & ~n282;
  assign n7069 = ~n364 & ~n376;
  assign n7070 = ~n427 & ~n768;
  assign n7071 = n7069 & n7070;
  assign n7072 = n164 & n7068;
  assign n7073 = n301 & n705;
  assign n7074 = n1684 & n1863;
  assign n7075 = n2397 & n3121;
  assign n7076 = n7074 & n7075;
  assign n7077 = n7072 & n7073;
  assign n7078 = n7060 & n7071;
  assign n7079 = n7077 & n7078;
  assign n7080 = n7058 & n7076;
  assign n7081 = n7079 & n7080;
  assign n7082 = n7067 & n7081;
  assign n7083 = ~n338 & n635;
  assign n7084 = ~n256 & n7083;
  assign n7085 = ~n174 & ~n284;
  assign n7086 = ~n356 & ~n687;
  assign n7087 = n7085 & n7086;
  assign n7088 = n1291 & n3277;
  assign n7089 = n7087 & n7088;
  assign n7090 = n717 & n2107;
  assign n7091 = n7089 & n7090;
  assign n7092 = n2448 & n7057;
  assign n7093 = n7084 & n7092;
  assign n7094 = n7091 & n7093;
  assign n7095 = n3350 & n7094;
  assign n7096 = n2306 & n7082;
  assign n7097 = n7095 & n7096;
  assign n7098 = n7052 & ~n7097;
  assign n7099 = ~n7052 & n7097;
  assign n7100 = ~n3275 & n3694;
  assign n7101 = ~n3373 & ~n3486;
  assign n7102 = ~n3487 & ~n7101;
  assign n7103 = n880 & n7102;
  assign n7104 = n748 & ~n3485;
  assign n7105 = ~n3370 & n3692;
  assign n7106 = ~n7100 & ~n7104;
  assign n7107 = ~n7105 & n7106;
  assign n7108 = ~n7103 & n7107;
  assign n7109 = ~n7099 & ~n7108;
  assign n7110 = ~n7098 & ~n7109;
  assign n7111 = ~n7014 & ~n7110;
  assign n7112 = ~n7011 & ~n7111;
  assign n7113 = ~n6956 & n6965;
  assign n7114 = n6956 & ~n6965;
  assign n7115 = ~n7113 & ~n7114;
  assign n7116 = ~n7112 & ~n7115;
  assign n7117 = ~n6966 & ~n7116;
  assign n7118 = ~n6905 & n6914;
  assign n7119 = n6905 & ~n6914;
  assign n7120 = ~n7118 & ~n7119;
  assign n7121 = ~n7117 & ~n7120;
  assign n7122 = ~n6915 & ~n7121;
  assign n7123 = ~n6860 & n6869;
  assign n7124 = n6860 & ~n6869;
  assign n7125 = ~n7123 & ~n7124;
  assign n7126 = ~n7122 & ~n7125;
  assign n7127 = ~n6870 & ~n7126;
  assign n7128 = ~n6483 & n6492;
  assign n7129 = ~n6493 & ~n7128;
  assign n7130 = ~n7127 & n7129;
  assign n7131 = n7127 & ~n7129;
  assign n7132 = ~n7130 & ~n7131;
  assign n7133 = ~n2919 & n3810;
  assign n7134 = n3886 & n6509;
  assign n7135 = ~n2835 & n3884;
  assign n7136 = ~n2778 & n4380;
  assign n7137 = ~n7133 & ~n7135;
  assign n7138 = ~n7136 & n7137;
  assign n7139 = ~n7134 & n7138;
  assign n7140 = pi29  & n7139;
  assign n7141 = ~pi29  & ~n7139;
  assign n7142 = ~n7140 & ~n7141;
  assign n7143 = n7132 & ~n7142;
  assign n7144 = ~n7130 & ~n7143;
  assign n7145 = n6818 & n6827;
  assign n7146 = ~n6818 & ~n6827;
  assign n7147 = ~n7145 & ~n7146;
  assign n7148 = ~n7144 & ~n7147;
  assign n7149 = ~n6828 & ~n7148;
  assign n7150 = n6806 & n6815;
  assign n7151 = ~n6806 & ~n6815;
  assign n7152 = ~n7150 & ~n7151;
  assign n7153 = ~n7149 & ~n7152;
  assign n7154 = ~n6816 & ~n7153;
  assign n7155 = ~n6505 & ~n6506;
  assign n7156 = ~n6515 & n7155;
  assign n7157 = n6515 & ~n7155;
  assign n7158 = ~n7156 & ~n7157;
  assign n7159 = ~n7154 & n7158;
  assign n7160 = n7154 & ~n7158;
  assign n7161 = ~n2674 & n3884;
  assign n7162 = n3886 & n6240;
  assign n7163 = ~n2708 & n3810;
  assign n7164 = ~n2589 & n4380;
  assign n7165 = ~n7161 & ~n7163;
  assign n7166 = ~n7164 & n7165;
  assign n7167 = ~n7162 & n7166;
  assign n7168 = pi29  & n7167;
  assign n7169 = ~pi29  & ~n7167;
  assign n7170 = ~n7168 & ~n7169;
  assign n7171 = ~n7160 & ~n7170;
  assign n7172 = ~n7159 & ~n7171;
  assign n7173 = n6804 & ~n7172;
  assign n7174 = ~n6804 & n7172;
  assign n7175 = n86 & ~n2412;
  assign n7176 = n4420 & n5579;
  assign n7177 = ~n2347 & n4600;
  assign n7178 = ~n2249 & n4615;
  assign n7179 = ~n7175 & ~n7177;
  assign n7180 = ~n7178 & n7179;
  assign n7181 = ~n7176 & n7180;
  assign n7182 = pi26  & n7181;
  assign n7183 = ~pi26  & ~n7181;
  assign n7184 = ~n7182 & ~n7183;
  assign n7185 = ~n7174 & ~n7184;
  assign n7186 = ~n7173 & ~n7185;
  assign n7187 = n6802 & ~n7186;
  assign n7188 = ~n6802 & n7186;
  assign n7189 = ~n1998 & n5109;
  assign n7190 = n5045 & n5151;
  assign n7191 = ~n2098 & n5044;
  assign n7192 = ~n1908 & n5130;
  assign n7193 = ~n7189 & ~n7191;
  assign n7194 = ~n7192 & n7193;
  assign n7195 = ~n7190 & n7194;
  assign n7196 = pi23  & n7195;
  assign n7197 = ~pi23  & ~n7195;
  assign n7198 = ~n7196 & ~n7197;
  assign n7199 = ~n7188 & ~n7198;
  assign n7200 = ~n7187 & ~n7199;
  assign n7201 = ~n6798 & ~n7200;
  assign n7202 = ~n6795 & ~n7201;
  assign n7203 = ~n6704 & ~n6705;
  assign n7204 = ~n6715 & n7203;
  assign n7205 = n6715 & ~n7203;
  assign n7206 = ~n7204 & ~n7205;
  assign n7207 = ~n7202 & n7206;
  assign n7208 = n7202 & ~n7206;
  assign n7209 = ~n1533 & n5853;
  assign n7210 = n4355 & n5241;
  assign n7211 = ~n1637 & n5240;
  assign n7212 = ~n1448 & n5866;
  assign n7213 = ~n7209 & ~n7211;
  assign n7214 = ~n7212 & n7213;
  assign n7215 = ~n7210 & n7214;
  assign n7216 = pi20  & n7215;
  assign n7217 = ~pi20  & ~n7215;
  assign n7218 = ~n7216 & ~n7217;
  assign n7219 = ~n7208 & ~n7218;
  assign n7220 = ~n7207 & ~n7219;
  assign n7221 = n6782 & ~n7220;
  assign n7222 = ~n6782 & n7220;
  assign n7223 = ~n1104 & n6323;
  assign n7224 = n3775 & n5983;
  assign n7225 = ~n1225 & n5982;
  assign n7226 = ~n878 & n6336;
  assign n7227 = ~n7223 & ~n7225;
  assign n7228 = ~n7226 & n7227;
  assign n7229 = ~n7224 & n7228;
  assign n7230 = pi17  & n7229;
  assign n7231 = ~pi17  & ~n7229;
  assign n7232 = ~n7230 & ~n7231;
  assign n7233 = ~n7222 & ~n7232;
  assign n7234 = ~n7221 & ~n7233;
  assign n7235 = ~n6778 & ~n7234;
  assign n7236 = ~n6775 & ~n7235;
  assign n7237 = ~n3855 & n6630;
  assign n7238 = ~n6625 & n6628;
  assign n7239 = ~n3883 & n7238;
  assign n7240 = ~n3900 & n6631;
  assign n7241 = ~n7237 & ~n7239;
  assign n7242 = ~n7240 & n7241;
  assign n7243 = pi14  & n7242;
  assign n7244 = ~pi14  & ~n7242;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = ~n7236 & ~n7245;
  assign n7247 = n7236 & n7245;
  assign n7248 = ~n7246 & ~n7247;
  assign n7249 = ~n6738 & ~n6739;
  assign n7250 = ~n6749 & n7249;
  assign n7251 = n6749 & ~n7249;
  assign n7252 = ~n7250 & ~n7251;
  assign n7253 = n7248 & n7252;
  assign n7254 = ~n7246 & ~n7253;
  assign n7255 = ~n6752 & ~n6753;
  assign n7256 = n6757 & n7255;
  assign n7257 = ~n6757 & ~n7255;
  assign n7258 = ~n7256 & ~n7257;
  assign n7259 = ~n7254 & n7258;
  assign n7260 = n7254 & ~n7258;
  assign n7261 = ~n7259 & ~n7260;
  assign n7262 = n6622 & ~n6628;
  assign n7263 = ~n3883 & n7262;
  assign n7264 = n4399 & n6631;
  assign n7265 = ~n3855 & n7238;
  assign n7266 = ~n3681 & n6630;
  assign n7267 = ~n7263 & ~n7265;
  assign n7268 = ~n7266 & n7267;
  assign n7269 = ~n7264 & n7268;
  assign n7270 = pi14  & n7269;
  assign n7271 = ~pi14  & ~n7269;
  assign n7272 = ~n7270 & ~n7271;
  assign n7273 = ~n7221 & ~n7222;
  assign n7274 = ~n7232 & n7273;
  assign n7275 = n7232 & ~n7273;
  assign n7276 = ~n7274 & ~n7275;
  assign n7277 = n6798 & n7200;
  assign n7278 = ~n7201 & ~n7277;
  assign n7279 = ~n1637 & n5853;
  assign n7280 = n4553 & n5241;
  assign n7281 = ~n1717 & n5240;
  assign n7282 = ~n1533 & n5866;
  assign n7283 = ~n7279 & ~n7281;
  assign n7284 = ~n7282 & n7283;
  assign n7285 = ~n7280 & n7284;
  assign n7286 = pi20  & n7285;
  assign n7287 = ~pi20  & ~n7285;
  assign n7288 = ~n7286 & ~n7287;
  assign n7289 = n7278 & ~n7288;
  assign n7290 = ~n7278 & n7288;
  assign n7291 = ~n7289 & ~n7290;
  assign n7292 = ~n7187 & ~n7188;
  assign n7293 = ~n7198 & n7292;
  assign n7294 = n7198 & ~n7292;
  assign n7295 = ~n7293 & ~n7294;
  assign n7296 = ~n2347 & n4615;
  assign n7297 = n4420 & n5596;
  assign n7298 = n86 & ~n2496;
  assign n7299 = ~n2412 & n4600;
  assign n7300 = ~n7296 & ~n7298;
  assign n7301 = ~n7299 & n7300;
  assign n7302 = ~n7297 & n7301;
  assign n7303 = pi26  & n7302;
  assign n7304 = ~pi26  & ~n7302;
  assign n7305 = ~n7303 & ~n7304;
  assign n7306 = ~n7159 & ~n7160;
  assign n7307 = ~n7170 & n7306;
  assign n7308 = n7170 & ~n7306;
  assign n7309 = ~n7307 & ~n7308;
  assign n7310 = ~n7305 & n7309;
  assign n7311 = n7305 & ~n7309;
  assign n7312 = ~n7310 & ~n7311;
  assign n7313 = ~n2778 & n3810;
  assign n7314 = n3886 & n6393;
  assign n7315 = ~n2708 & n3884;
  assign n7316 = ~n2674 & n4380;
  assign n7317 = ~n7313 & ~n7315;
  assign n7318 = ~n7316 & n7317;
  assign n7319 = ~n7314 & n7318;
  assign n7320 = pi29  & n7319;
  assign n7321 = ~pi29  & ~n7319;
  assign n7322 = ~n7320 & ~n7321;
  assign n7323 = n7149 & n7152;
  assign n7324 = ~n7153 & ~n7323;
  assign n7325 = ~n7322 & n7324;
  assign n7326 = n7322 & ~n7324;
  assign n7327 = n86 & ~n2589;
  assign n7328 = n4420 & n6016;
  assign n7329 = ~n2496 & n4600;
  assign n7330 = ~n2412 & n4615;
  assign n7331 = ~n7327 & ~n7329;
  assign n7332 = ~n7330 & n7331;
  assign n7333 = ~n7328 & n7332;
  assign n7334 = pi26  & n7333;
  assign n7335 = ~pi26  & ~n7333;
  assign n7336 = ~n7334 & ~n7335;
  assign n7337 = ~n7326 & ~n7336;
  assign n7338 = ~n7325 & ~n7337;
  assign n7339 = n7312 & ~n7338;
  assign n7340 = ~n7310 & ~n7339;
  assign n7341 = ~n7173 & ~n7174;
  assign n7342 = ~n7184 & n7341;
  assign n7343 = n7184 & ~n7341;
  assign n7344 = ~n7342 & ~n7343;
  assign n7345 = ~n7340 & n7344;
  assign n7346 = n7340 & ~n7344;
  assign n7347 = ~n2098 & n5109;
  assign n7348 = n4979 & n5045;
  assign n7349 = ~n2146 & n5044;
  assign n7350 = ~n1998 & n5130;
  assign n7351 = ~n7347 & ~n7349;
  assign n7352 = ~n7350 & n7351;
  assign n7353 = ~n7348 & n7352;
  assign n7354 = pi23  & n7353;
  assign n7355 = ~pi23  & ~n7353;
  assign n7356 = ~n7354 & ~n7355;
  assign n7357 = ~n7346 & ~n7356;
  assign n7358 = ~n7345 & ~n7357;
  assign n7359 = n7295 & ~n7358;
  assign n7360 = ~n7295 & n7358;
  assign n7361 = ~n1717 & n5853;
  assign n7362 = n4537 & n5241;
  assign n7363 = ~n1841 & n5240;
  assign n7364 = ~n1637 & n5866;
  assign n7365 = ~n7361 & ~n7363;
  assign n7366 = ~n7364 & n7365;
  assign n7367 = ~n7362 & n7366;
  assign n7368 = pi20  & n7367;
  assign n7369 = ~pi20  & ~n7367;
  assign n7370 = ~n7368 & ~n7369;
  assign n7371 = ~n7360 & ~n7370;
  assign n7372 = ~n7359 & ~n7371;
  assign n7373 = n7291 & ~n7372;
  assign n7374 = ~n7289 & ~n7373;
  assign n7375 = ~n7207 & ~n7208;
  assign n7376 = ~n7218 & n7375;
  assign n7377 = n7218 & ~n7375;
  assign n7378 = ~n7376 & ~n7377;
  assign n7379 = ~n7374 & n7378;
  assign n7380 = n7374 & ~n7378;
  assign n7381 = ~n1225 & n6323;
  assign n7382 = n4135 & n5983;
  assign n7383 = ~n1345 & n5982;
  assign n7384 = ~n1104 & n6336;
  assign n7385 = ~n7381 & ~n7383;
  assign n7386 = ~n7384 & n7385;
  assign n7387 = ~n7382 & n7386;
  assign n7388 = pi17  & n7387;
  assign n7389 = ~pi17  & ~n7387;
  assign n7390 = ~n7388 & ~n7389;
  assign n7391 = ~n7380 & ~n7390;
  assign n7392 = ~n7379 & ~n7391;
  assign n7393 = n7276 & ~n7392;
  assign n7394 = ~n7276 & n7392;
  assign n7395 = ~n3855 & n7262;
  assign n7396 = n3972 & n6631;
  assign n7397 = ~n987 & n6630;
  assign n7398 = ~n3681 & n7238;
  assign n7399 = ~n7395 & ~n7397;
  assign n7400 = ~n7398 & n7399;
  assign n7401 = ~n7396 & n7400;
  assign n7402 = pi14  & n7401;
  assign n7403 = ~pi14  & ~n7401;
  assign n7404 = ~n7402 & ~n7403;
  assign n7405 = ~n7394 & ~n7404;
  assign n7406 = ~n7393 & ~n7405;
  assign n7407 = ~n7272 & ~n7406;
  assign n7408 = n6778 & n7234;
  assign n7409 = ~n7235 & ~n7408;
  assign n7410 = n7272 & ~n7406;
  assign n7411 = ~n7272 & n7406;
  assign n7412 = ~n7410 & ~n7411;
  assign n7413 = n7409 & ~n7412;
  assign n7414 = ~n7407 & ~n7413;
  assign n7415 = ~n7248 & ~n7252;
  assign n7416 = ~n7253 & ~n7415;
  assign n7417 = ~n7414 & n7416;
  assign n7418 = ~n7409 & n7412;
  assign n7419 = ~n7413 & ~n7418;
  assign n7420 = pi10  & ~pi11 ;
  assign n7421 = ~pi10  & pi11 ;
  assign n7422 = ~n7420 & ~n7421;
  assign n7423 = pi8  & ~pi9 ;
  assign n7424 = ~pi8  & pi9 ;
  assign n7425 = ~n7423 & ~n7424;
  assign n7426 = ~pi9  & pi10 ;
  assign n7427 = pi9  & ~pi10 ;
  assign n7428 = ~n7426 & ~n7427;
  assign n7429 = n7425 & n7428;
  assign n7430 = ~n7422 & n7429;
  assign n7431 = ~n7422 & ~n7425;
  assign n7432 = ~n3897 & n7431;
  assign n7433 = ~n7430 & ~n7432;
  assign n7434 = ~n3883 & ~n7433;
  assign n7435 = pi11  & ~n7434;
  assign n7436 = ~pi11  & n7434;
  assign n7437 = ~n7435 & ~n7436;
  assign n7438 = ~n1345 & n6323;
  assign n7439 = n4152 & n5983;
  assign n7440 = ~n1448 & n5982;
  assign n7441 = ~n1225 & n6336;
  assign n7442 = ~n7438 & ~n7440;
  assign n7443 = ~n7441 & n7442;
  assign n7444 = ~n7439 & n7443;
  assign n7445 = ~pi17  & ~n7444;
  assign n7446 = pi17  & n7444;
  assign n7447 = ~n7445 & ~n7446;
  assign n7448 = ~n7291 & n7372;
  assign n7449 = ~n7373 & ~n7448;
  assign n7450 = ~n7447 & n7449;
  assign n7451 = ~n7447 & ~n7449;
  assign n7452 = n7447 & n7449;
  assign n7453 = ~n7451 & ~n7452;
  assign n7454 = ~n7359 & ~n7360;
  assign n7455 = ~n7370 & n7454;
  assign n7456 = n7370 & ~n7454;
  assign n7457 = ~n7455 & ~n7456;
  assign n7458 = ~n2098 & n5130;
  assign n7459 = n5045 & n5359;
  assign n7460 = ~n2146 & n5109;
  assign n7461 = ~n2249 & n5044;
  assign n7462 = ~n7458 & ~n7460;
  assign n7463 = ~n7461 & n7462;
  assign n7464 = ~n7459 & n7463;
  assign n7465 = ~pi23  & ~n7464;
  assign n7466 = pi23  & n7464;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = ~n7312 & n7338;
  assign n7469 = ~n7339 & ~n7468;
  assign n7470 = ~n7467 & n7469;
  assign n7471 = ~n7467 & ~n7469;
  assign n7472 = n7467 & n7469;
  assign n7473 = ~n7471 & ~n7472;
  assign n7474 = ~n7325 & ~n7326;
  assign n7475 = ~n7336 & n7474;
  assign n7476 = n7336 & ~n7474;
  assign n7477 = ~n7475 & ~n7476;
  assign n7478 = ~n2708 & n4380;
  assign n7479 = n3886 & n6222;
  assign n7480 = ~n2835 & n3810;
  assign n7481 = ~n2778 & n3884;
  assign n7482 = ~n7478 & ~n7480;
  assign n7483 = ~n7481 & n7482;
  assign n7484 = ~n7479 & n7483;
  assign n7485 = pi29  & n7484;
  assign n7486 = ~pi29  & ~n7484;
  assign n7487 = ~n7485 & ~n7486;
  assign n7488 = n7144 & n7147;
  assign n7489 = ~n7148 & ~n7488;
  assign n7490 = ~n7487 & n7489;
  assign n7491 = n7487 & ~n7489;
  assign n7492 = ~n2496 & n4615;
  assign n7493 = n4420 & n5776;
  assign n7494 = n86 & ~n2674;
  assign n7495 = ~n2589 & n4600;
  assign n7496 = ~n7492 & ~n7494;
  assign n7497 = ~n7495 & n7496;
  assign n7498 = ~n7493 & n7497;
  assign n7499 = pi26  & n7498;
  assign n7500 = ~pi26  & ~n7498;
  assign n7501 = ~n7499 & ~n7500;
  assign n7502 = ~n7491 & ~n7501;
  assign n7503 = ~n7490 & ~n7502;
  assign n7504 = n7477 & ~n7503;
  assign n7505 = ~n7477 & n7503;
  assign n7506 = ~n2146 & n5130;
  assign n7507 = n5045 & n5343;
  assign n7508 = ~n2347 & n5044;
  assign n7509 = ~n2249 & n5109;
  assign n7510 = ~n7506 & ~n7508;
  assign n7511 = ~n7509 & n7510;
  assign n7512 = ~n7507 & n7511;
  assign n7513 = pi23  & n7512;
  assign n7514 = ~pi23  & ~n7512;
  assign n7515 = ~n7513 & ~n7514;
  assign n7516 = ~n7505 & ~n7515;
  assign n7517 = ~n7504 & ~n7516;
  assign n7518 = ~n7473 & ~n7517;
  assign n7519 = ~n7470 & ~n7518;
  assign n7520 = ~n7345 & ~n7346;
  assign n7521 = ~n7356 & n7520;
  assign n7522 = n7356 & ~n7520;
  assign n7523 = ~n7521 & ~n7522;
  assign n7524 = ~n7519 & n7523;
  assign n7525 = n7519 & ~n7523;
  assign n7526 = ~n1841 & n5853;
  assign n7527 = n4762 & n5241;
  assign n7528 = ~n1908 & n5240;
  assign n7529 = ~n1717 & n5866;
  assign n7530 = ~n7526 & ~n7528;
  assign n7531 = ~n7529 & n7530;
  assign n7532 = ~n7527 & n7531;
  assign n7533 = pi20  & n7532;
  assign n7534 = ~pi20  & ~n7532;
  assign n7535 = ~n7533 & ~n7534;
  assign n7536 = ~n7525 & ~n7535;
  assign n7537 = ~n7524 & ~n7536;
  assign n7538 = n7457 & ~n7537;
  assign n7539 = ~n7457 & n7537;
  assign n7540 = ~n1448 & n6323;
  assign n7541 = n4453 & n5983;
  assign n7542 = ~n1533 & n5982;
  assign n7543 = ~n1345 & n6336;
  assign n7544 = ~n7540 & ~n7542;
  assign n7545 = ~n7543 & n7544;
  assign n7546 = ~n7541 & n7545;
  assign n7547 = pi17  & n7546;
  assign n7548 = ~pi17  & ~n7546;
  assign n7549 = ~n7547 & ~n7548;
  assign n7550 = ~n7539 & ~n7549;
  assign n7551 = ~n7538 & ~n7550;
  assign n7552 = ~n7453 & ~n7551;
  assign n7553 = ~n7450 & ~n7552;
  assign n7554 = ~n7379 & ~n7380;
  assign n7555 = ~n7390 & n7554;
  assign n7556 = n7390 & ~n7554;
  assign n7557 = ~n7555 & ~n7556;
  assign n7558 = ~n7553 & n7557;
  assign n7559 = n7553 & ~n7557;
  assign n7560 = ~n878 & n6630;
  assign n7561 = n3687 & n6631;
  assign n7562 = ~n987 & n7238;
  assign n7563 = ~n3681 & n7262;
  assign n7564 = ~n7560 & ~n7562;
  assign n7565 = ~n7563 & n7564;
  assign n7566 = ~n7561 & n7565;
  assign n7567 = pi14  & n7566;
  assign n7568 = ~pi14  & ~n7566;
  assign n7569 = ~n7567 & ~n7568;
  assign n7570 = ~n7559 & ~n7569;
  assign n7571 = ~n7558 & ~n7570;
  assign n7572 = ~n7437 & ~n7571;
  assign n7573 = n7437 & n7571;
  assign n7574 = ~n7393 & ~n7394;
  assign n7575 = ~n7404 & n7574;
  assign n7576 = n7404 & ~n7574;
  assign n7577 = ~n7575 & ~n7576;
  assign n7578 = ~n7573 & n7577;
  assign n7579 = ~n7572 & ~n7578;
  assign n7580 = n7419 & ~n7579;
  assign n7581 = n7453 & n7551;
  assign n7582 = ~n7552 & ~n7581;
  assign n7583 = ~n987 & n7262;
  assign n7584 = n3791 & n6631;
  assign n7585 = ~n1104 & n6630;
  assign n7586 = ~n878 & n7238;
  assign n7587 = ~n7583 & ~n7585;
  assign n7588 = ~n7586 & n7587;
  assign n7589 = ~n7584 & n7588;
  assign n7590 = pi14  & n7589;
  assign n7591 = ~pi14  & ~n7589;
  assign n7592 = ~n7590 & ~n7591;
  assign n7593 = n7582 & ~n7592;
  assign n7594 = n7582 & n7592;
  assign n7595 = ~n7582 & ~n7592;
  assign n7596 = ~n7594 & ~n7595;
  assign n7597 = ~n7538 & ~n7539;
  assign n7598 = ~n7549 & n7597;
  assign n7599 = n7549 & ~n7597;
  assign n7600 = ~n7598 & ~n7599;
  assign n7601 = n7473 & n7517;
  assign n7602 = ~n7518 & ~n7601;
  assign n7603 = ~n1908 & n5853;
  assign n7604 = n4779 & n5241;
  assign n7605 = ~n1998 & n5240;
  assign n7606 = ~n1841 & n5866;
  assign n7607 = ~n7603 & ~n7605;
  assign n7608 = ~n7606 & n7607;
  assign n7609 = ~n7604 & n7608;
  assign n7610 = pi20  & n7609;
  assign n7611 = ~pi20  & ~n7609;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = n7602 & ~n7612;
  assign n7614 = ~n7602 & n7612;
  assign n7615 = ~n7613 & ~n7614;
  assign n7616 = ~n7504 & ~n7505;
  assign n7617 = ~n7515 & n7616;
  assign n7618 = n7515 & ~n7616;
  assign n7619 = ~n7617 & ~n7618;
  assign n7620 = ~n2919 & n3884;
  assign n7621 = n3886 & n6809;
  assign n7622 = ~n2951 & n3810;
  assign n7623 = ~n2835 & n4380;
  assign n7624 = ~n7620 & ~n7622;
  assign n7625 = ~n7623 & n7624;
  assign n7626 = ~n7621 & n7625;
  assign n7627 = pi29  & n7626;
  assign n7628 = ~pi29  & ~n7626;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = n7122 & n7125;
  assign n7631 = ~n7126 & ~n7630;
  assign n7632 = ~n7629 & n7631;
  assign n7633 = ~n2919 & n4380;
  assign n7634 = n3886 & n6821;
  assign n7635 = ~n2951 & n3884;
  assign n7636 = ~n3031 & n3810;
  assign n7637 = ~n7633 & ~n7635;
  assign n7638 = ~n7636 & n7637;
  assign n7639 = ~n7634 & n7638;
  assign n7640 = pi29  & n7639;
  assign n7641 = ~pi29  & ~n7639;
  assign n7642 = ~n7640 & ~n7641;
  assign n7643 = n7117 & n7120;
  assign n7644 = ~n7121 & ~n7643;
  assign n7645 = ~n7642 & n7644;
  assign n7646 = ~n2951 & n4380;
  assign n7647 = n3886 & n6486;
  assign n7648 = ~n3118 & n3810;
  assign n7649 = ~n3031 & n3884;
  assign n7650 = ~n7646 & ~n7648;
  assign n7651 = ~n7649 & n7650;
  assign n7652 = ~n7647 & n7651;
  assign n7653 = ~pi29  & ~n7652;
  assign n7654 = pi29  & n7652;
  assign n7655 = ~n7653 & ~n7654;
  assign n7656 = n7112 & n7115;
  assign n7657 = ~n7116 & ~n7656;
  assign n7658 = ~n7655 & n7657;
  assign n7659 = ~n7655 & ~n7657;
  assign n7660 = n7655 & n7657;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = ~n3182 & n3810;
  assign n7663 = n3886 & n6863;
  assign n7664 = ~n3118 & n3884;
  assign n7665 = ~n3031 & n4380;
  assign n7666 = ~n7662 & ~n7664;
  assign n7667 = ~n7665 & n7666;
  assign n7668 = ~n7663 & n7667;
  assign n7669 = ~pi29  & ~n7668;
  assign n7670 = pi29  & n7668;
  assign n7671 = ~n7669 & ~n7670;
  assign n7672 = n7014 & n7110;
  assign n7673 = ~n7111 & ~n7672;
  assign n7674 = ~n7671 & n7673;
  assign n7675 = ~n7671 & ~n7673;
  assign n7676 = n7671 & n7673;
  assign n7677 = ~n7675 & ~n7676;
  assign n7678 = ~n3118 & n4380;
  assign n7679 = n3886 & n6908;
  assign n7680 = ~n3241 & n3810;
  assign n7681 = ~n3182 & n3884;
  assign n7682 = ~n7678 & ~n7680;
  assign n7683 = ~n7681 & n7682;
  assign n7684 = ~n7679 & n7683;
  assign n7685 = ~pi29  & ~n7684;
  assign n7686 = pi29  & n7684;
  assign n7687 = ~n7685 & ~n7686;
  assign n7688 = ~n7098 & ~n7099;
  assign n7689 = ~n7108 & n7688;
  assign n7690 = n7108 & ~n7688;
  assign n7691 = ~n7689 & ~n7690;
  assign n7692 = ~n7687 & n7691;
  assign n7693 = ~n3275 & n3810;
  assign n7694 = n3886 & n6959;
  assign n7695 = ~n3241 & n3884;
  assign n7696 = ~n3182 & n4380;
  assign n7697 = ~n7693 & ~n7695;
  assign n7698 = ~n7696 & n7697;
  assign n7699 = ~n7694 & n7698;
  assign n7700 = ~pi29  & ~n7699;
  assign n7701 = pi29  & n7699;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = ~n7040 & n7051;
  assign n7704 = n7040 & ~n7051;
  assign n7705 = ~n7703 & ~n7704;
  assign n7706 = ~n7702 & ~n7705;
  assign n7707 = ~n3241 & n4380;
  assign n7708 = n3886 & n7004;
  assign n7709 = ~n3275 & n3884;
  assign n7710 = ~n3370 & n3810;
  assign n7711 = ~n7707 & ~n7709;
  assign n7712 = ~n7710 & n7711;
  assign n7713 = ~n7708 & n7712;
  assign n7714 = ~pi29  & ~n7713;
  assign n7715 = pi29  & n7713;
  assign n7716 = ~n7714 & ~n7715;
  assign n7717 = ~n3427 & n3692;
  assign n7718 = ~n3485 & n3694;
  assign n7719 = ~n3427 & n3485;
  assign n7720 = ~n7042 & ~n7719;
  assign n7721 = n880 & ~n7720;
  assign n7722 = ~n7717 & ~n7718;
  assign n7723 = ~n7721 & n7722;
  assign n7724 = ~n7716 & ~n7723;
  assign n7725 = ~n7716 & n7723;
  assign n7726 = n7716 & ~n7723;
  assign n7727 = ~n7725 & ~n7726;
  assign n7728 = ~n746 & ~n3427;
  assign n7729 = ~n3427 & ~n3807;
  assign n7730 = ~n3427 & n3884;
  assign n7731 = ~n3485 & n4380;
  assign n7732 = n3886 & ~n7720;
  assign n7733 = ~n7730 & ~n7731;
  assign n7734 = ~n7732 & n7733;
  assign n7735 = pi29  & ~n7729;
  assign n7736 = n7734 & n7735;
  assign n7737 = ~n3427 & n3810;
  assign n7738 = n3886 & n7045;
  assign n7739 = ~n3485 & n3884;
  assign n7740 = ~n3370 & n4380;
  assign n7741 = ~n7737 & ~n7739;
  assign n7742 = ~n7740 & n7741;
  assign n7743 = ~n7738 & n7742;
  assign n7744 = n7736 & n7743;
  assign n7745 = n7728 & n7744;
  assign n7746 = ~n3275 & n4380;
  assign n7747 = n3886 & n7102;
  assign n7748 = ~n3485 & n3810;
  assign n7749 = ~n3370 & n3884;
  assign n7750 = ~n7746 & ~n7748;
  assign n7751 = ~n7749 & n7750;
  assign n7752 = ~n7747 & n7751;
  assign n7753 = ~pi29  & ~n7752;
  assign n7754 = pi29  & n7752;
  assign n7755 = ~n7753 & ~n7754;
  assign n7756 = ~n7728 & n7744;
  assign n7757 = n7728 & ~n7744;
  assign n7758 = ~n7756 & ~n7757;
  assign n7759 = ~n7755 & ~n7758;
  assign n7760 = ~n7745 & ~n7759;
  assign n7761 = ~n7727 & ~n7760;
  assign n7762 = ~n7724 & ~n7761;
  assign n7763 = n7702 & n7705;
  assign n7764 = ~n7706 & ~n7763;
  assign n7765 = ~n7762 & n7764;
  assign n7766 = ~n7706 & ~n7765;
  assign n7767 = n7687 & ~n7691;
  assign n7768 = ~n7692 & ~n7767;
  assign n7769 = ~n7766 & n7768;
  assign n7770 = ~n7692 & ~n7769;
  assign n7771 = ~n7677 & ~n7770;
  assign n7772 = ~n7674 & ~n7771;
  assign n7773 = ~n7661 & ~n7772;
  assign n7774 = ~n7658 & ~n7773;
  assign n7775 = n7642 & ~n7644;
  assign n7776 = ~n7645 & ~n7775;
  assign n7777 = ~n7774 & n7776;
  assign n7778 = ~n7645 & ~n7777;
  assign n7779 = n7629 & ~n7631;
  assign n7780 = ~n7632 & ~n7779;
  assign n7781 = ~n7778 & n7780;
  assign n7782 = ~n7632 & ~n7781;
  assign n7783 = ~n7132 & n7142;
  assign n7784 = ~n7143 & ~n7783;
  assign n7785 = ~n7782 & n7784;
  assign n7786 = ~n2674 & n4600;
  assign n7787 = n4420 & n6240;
  assign n7788 = n86 & ~n2708;
  assign n7789 = ~n2589 & n4615;
  assign n7790 = ~n7786 & ~n7788;
  assign n7791 = ~n7789 & n7790;
  assign n7792 = ~n7787 & n7791;
  assign n7793 = ~pi26  & ~n7792;
  assign n7794 = pi26  & n7792;
  assign n7795 = ~n7793 & ~n7794;
  assign n7796 = n7782 & ~n7784;
  assign n7797 = ~n7785 & ~n7796;
  assign n7798 = ~n7795 & n7797;
  assign n7799 = ~n7785 & ~n7798;
  assign n7800 = ~n7490 & ~n7491;
  assign n7801 = ~n7501 & n7800;
  assign n7802 = n7501 & ~n7800;
  assign n7803 = ~n7801 & ~n7802;
  assign n7804 = ~n7799 & n7803;
  assign n7805 = n7799 & ~n7803;
  assign n7806 = ~n2412 & n5044;
  assign n7807 = n5045 & n5579;
  assign n7808 = ~n2347 & n5109;
  assign n7809 = ~n2249 & n5130;
  assign n7810 = ~n7806 & ~n7808;
  assign n7811 = ~n7809 & n7810;
  assign n7812 = ~n7807 & n7811;
  assign n7813 = pi23  & n7812;
  assign n7814 = ~pi23  & ~n7812;
  assign n7815 = ~n7813 & ~n7814;
  assign n7816 = ~n7805 & ~n7815;
  assign n7817 = ~n7804 & ~n7816;
  assign n7818 = n7619 & ~n7817;
  assign n7819 = ~n7619 & n7817;
  assign n7820 = ~n1998 & n5853;
  assign n7821 = n5151 & n5241;
  assign n7822 = ~n2098 & n5240;
  assign n7823 = ~n1908 & n5866;
  assign n7824 = ~n7820 & ~n7822;
  assign n7825 = ~n7823 & n7824;
  assign n7826 = ~n7821 & n7825;
  assign n7827 = pi20  & n7826;
  assign n7828 = ~pi20  & ~n7826;
  assign n7829 = ~n7827 & ~n7828;
  assign n7830 = ~n7819 & ~n7829;
  assign n7831 = ~n7818 & ~n7830;
  assign n7832 = n7615 & ~n7831;
  assign n7833 = ~n7613 & ~n7832;
  assign n7834 = ~n7524 & ~n7525;
  assign n7835 = ~n7535 & n7834;
  assign n7836 = n7535 & ~n7834;
  assign n7837 = ~n7835 & ~n7836;
  assign n7838 = ~n7833 & n7837;
  assign n7839 = n7833 & ~n7837;
  assign n7840 = ~n1533 & n6323;
  assign n7841 = n4355 & n5983;
  assign n7842 = ~n1637 & n5982;
  assign n7843 = ~n1448 & n6336;
  assign n7844 = ~n7840 & ~n7842;
  assign n7845 = ~n7843 & n7844;
  assign n7846 = ~n7841 & n7845;
  assign n7847 = pi17  & n7846;
  assign n7848 = ~pi17  & ~n7846;
  assign n7849 = ~n7847 & ~n7848;
  assign n7850 = ~n7839 & ~n7849;
  assign n7851 = ~n7838 & ~n7850;
  assign n7852 = n7600 & ~n7851;
  assign n7853 = ~n7600 & n7851;
  assign n7854 = ~n1104 & n7238;
  assign n7855 = n3775 & n6631;
  assign n7856 = ~n1225 & n6630;
  assign n7857 = ~n878 & n7262;
  assign n7858 = ~n7854 & ~n7856;
  assign n7859 = ~n7857 & n7858;
  assign n7860 = ~n7855 & n7859;
  assign n7861 = pi14  & n7860;
  assign n7862 = ~pi14  & ~n7860;
  assign n7863 = ~n7861 & ~n7862;
  assign n7864 = ~n7853 & ~n7863;
  assign n7865 = ~n7852 & ~n7864;
  assign n7866 = ~n7596 & ~n7865;
  assign n7867 = ~n7593 & ~n7866;
  assign n7868 = ~n3855 & n7430;
  assign n7869 = n7425 & ~n7428;
  assign n7870 = ~n3883 & n7869;
  assign n7871 = ~n3900 & n7431;
  assign n7872 = ~n7868 & ~n7870;
  assign n7873 = ~n7871 & n7872;
  assign n7874 = pi11  & n7873;
  assign n7875 = ~pi11  & ~n7873;
  assign n7876 = ~n7874 & ~n7875;
  assign n7877 = ~n7867 & ~n7876;
  assign n7878 = n7867 & n7876;
  assign n7879 = ~n7877 & ~n7878;
  assign n7880 = ~n7558 & ~n7559;
  assign n7881 = ~n7569 & n7880;
  assign n7882 = n7569 & ~n7880;
  assign n7883 = ~n7881 & ~n7882;
  assign n7884 = n7879 & n7883;
  assign n7885 = ~n7877 & ~n7884;
  assign n7886 = ~n7572 & ~n7573;
  assign n7887 = n7577 & n7886;
  assign n7888 = ~n7577 & ~n7886;
  assign n7889 = ~n7887 & ~n7888;
  assign n7890 = ~n7885 & n7889;
  assign n7891 = n7885 & ~n7889;
  assign n7892 = ~n7890 & ~n7891;
  assign n7893 = ~n7879 & ~n7883;
  assign n7894 = ~n7884 & ~n7893;
  assign n7895 = n7422 & ~n7425;
  assign n7896 = ~n3883 & n7895;
  assign n7897 = n4399 & n7431;
  assign n7898 = ~n3855 & n7869;
  assign n7899 = ~n3681 & n7430;
  assign n7900 = ~n7896 & ~n7898;
  assign n7901 = ~n7899 & n7900;
  assign n7902 = ~n7897 & n7901;
  assign n7903 = pi11  & n7902;
  assign n7904 = ~pi11  & ~n7902;
  assign n7905 = ~n7903 & ~n7904;
  assign n7906 = ~n7852 & ~n7853;
  assign n7907 = ~n7863 & n7906;
  assign n7908 = n7863 & ~n7906;
  assign n7909 = ~n7907 & ~n7908;
  assign n7910 = ~n1637 & n6323;
  assign n7911 = n4553 & n5983;
  assign n7912 = ~n1717 & n5982;
  assign n7913 = ~n1533 & n6336;
  assign n7914 = ~n7910 & ~n7912;
  assign n7915 = ~n7913 & n7914;
  assign n7916 = ~n7911 & n7915;
  assign n7917 = ~pi17  & ~n7916;
  assign n7918 = pi17  & n7916;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = ~n7615 & n7831;
  assign n7921 = ~n7832 & ~n7920;
  assign n7922 = ~n7919 & n7921;
  assign n7923 = ~n7919 & ~n7921;
  assign n7924 = n7919 & n7921;
  assign n7925 = ~n7923 & ~n7924;
  assign n7926 = ~n7818 & ~n7819;
  assign n7927 = ~n7829 & n7926;
  assign n7928 = n7829 & ~n7926;
  assign n7929 = ~n7927 & ~n7928;
  assign n7930 = n7778 & ~n7780;
  assign n7931 = ~n7781 & ~n7930;
  assign n7932 = n86 & ~n2778;
  assign n7933 = n4420 & n6393;
  assign n7934 = ~n2708 & n4600;
  assign n7935 = ~n2674 & n4615;
  assign n7936 = ~n7932 & ~n7934;
  assign n7937 = ~n7935 & n7936;
  assign n7938 = ~n7933 & n7937;
  assign n7939 = pi26  & n7938;
  assign n7940 = ~pi26  & ~n7938;
  assign n7941 = ~n7939 & ~n7940;
  assign n7942 = n7931 & ~n7941;
  assign n7943 = n7774 & ~n7776;
  assign n7944 = ~n7777 & ~n7943;
  assign n7945 = ~n2708 & n4615;
  assign n7946 = n4420 & n6222;
  assign n7947 = n86 & ~n2835;
  assign n7948 = ~n2778 & n4600;
  assign n7949 = ~n7945 & ~n7947;
  assign n7950 = ~n7948 & n7949;
  assign n7951 = ~n7946 & n7950;
  assign n7952 = pi26  & n7951;
  assign n7953 = ~pi26  & ~n7951;
  assign n7954 = ~n7952 & ~n7953;
  assign n7955 = n7944 & ~n7954;
  assign n7956 = n7661 & n7772;
  assign n7957 = ~n7773 & ~n7956;
  assign n7958 = n86 & ~n2919;
  assign n7959 = n4420 & n6509;
  assign n7960 = ~n2835 & n4600;
  assign n7961 = ~n2778 & n4615;
  assign n7962 = ~n7958 & ~n7960;
  assign n7963 = ~n7961 & n7962;
  assign n7964 = ~n7959 & n7963;
  assign n7965 = pi26  & n7964;
  assign n7966 = ~pi26  & ~n7964;
  assign n7967 = ~n7965 & ~n7966;
  assign n7968 = n7957 & ~n7967;
  assign n7969 = n7677 & n7770;
  assign n7970 = ~n7771 & ~n7969;
  assign n7971 = ~n2919 & n4600;
  assign n7972 = n4420 & n6809;
  assign n7973 = n86 & ~n2951;
  assign n7974 = ~n2835 & n4615;
  assign n7975 = ~n7971 & ~n7973;
  assign n7976 = ~n7974 & n7975;
  assign n7977 = ~n7972 & n7976;
  assign n7978 = pi26  & n7977;
  assign n7979 = ~pi26  & ~n7977;
  assign n7980 = ~n7978 & ~n7979;
  assign n7981 = n7970 & ~n7980;
  assign n7982 = n7766 & ~n7768;
  assign n7983 = ~n7769 & ~n7982;
  assign n7984 = ~n2919 & n4615;
  assign n7985 = n4420 & n6821;
  assign n7986 = ~n2951 & n4600;
  assign n7987 = n86 & ~n3031;
  assign n7988 = ~n7984 & ~n7986;
  assign n7989 = ~n7987 & n7988;
  assign n7990 = ~n7985 & n7989;
  assign n7991 = pi26  & n7990;
  assign n7992 = ~pi26  & ~n7990;
  assign n7993 = ~n7991 & ~n7992;
  assign n7994 = n7983 & ~n7993;
  assign n7995 = n7762 & ~n7764;
  assign n7996 = ~n7765 & ~n7995;
  assign n7997 = ~n2951 & n4615;
  assign n7998 = n4420 & n6486;
  assign n7999 = n86 & ~n3118;
  assign n8000 = ~n3031 & n4600;
  assign n8001 = ~n7997 & ~n7999;
  assign n8002 = ~n8000 & n8001;
  assign n8003 = ~n7998 & n8002;
  assign n8004 = pi26  & n8003;
  assign n8005 = ~pi26  & ~n8003;
  assign n8006 = ~n8004 & ~n8005;
  assign n8007 = n7996 & ~n8006;
  assign n8008 = n86 & ~n3182;
  assign n8009 = n4420 & n6863;
  assign n8010 = ~n3118 & n4600;
  assign n8011 = ~n3031 & n4615;
  assign n8012 = ~n8008 & ~n8010;
  assign n8013 = ~n8011 & n8012;
  assign n8014 = ~n8009 & n8013;
  assign n8015 = pi26  & n8014;
  assign n8016 = ~pi26  & ~n8014;
  assign n8017 = ~n8015 & ~n8016;
  assign n8018 = n7727 & n7760;
  assign n8019 = ~n7761 & ~n8018;
  assign n8020 = ~n8017 & n8019;
  assign n8021 = ~n3118 & n4615;
  assign n8022 = n4420 & n6908;
  assign n8023 = n86 & ~n3241;
  assign n8024 = ~n3182 & n4600;
  assign n8025 = ~n8021 & ~n8023;
  assign n8026 = ~n8024 & n8025;
  assign n8027 = ~n8022 & n8026;
  assign n8028 = ~pi26  & ~n8027;
  assign n8029 = pi26  & n8027;
  assign n8030 = ~n8028 & ~n8029;
  assign n8031 = n7755 & n7758;
  assign n8032 = ~n7759 & ~n8031;
  assign n8033 = ~n8030 & n8032;
  assign n8034 = ~n8030 & ~n8032;
  assign n8035 = n8030 & n8032;
  assign n8036 = ~n8034 & ~n8035;
  assign n8037 = n86 & ~n3275;
  assign n8038 = n4420 & n6959;
  assign n8039 = ~n3241 & n4600;
  assign n8040 = ~n3182 & n4615;
  assign n8041 = ~n8037 & ~n8039;
  assign n8042 = ~n8040 & n8041;
  assign n8043 = ~n8038 & n8042;
  assign n8044 = ~pi26  & ~n8043;
  assign n8045 = pi26  & n8043;
  assign n8046 = ~n8044 & ~n8045;
  assign n8047 = pi29  & ~n7736;
  assign n8048 = n7743 & ~n8047;
  assign n8049 = ~n7743 & n8047;
  assign n8050 = ~n8048 & ~n8049;
  assign n8051 = ~n8046 & n8050;
  assign n8052 = ~n8046 & ~n8050;
  assign n8053 = n8046 & n8050;
  assign n8054 = ~n8052 & ~n8053;
  assign n8055 = ~n3241 & n4615;
  assign n8056 = n4420 & n7004;
  assign n8057 = ~n3275 & n4600;
  assign n8058 = n86 & ~n3370;
  assign n8059 = ~n8055 & ~n8057;
  assign n8060 = ~n8058 & n8059;
  assign n8061 = ~n8056 & n8060;
  assign n8062 = pi26  & n8061;
  assign n8063 = ~pi26  & ~n8061;
  assign n8064 = ~n8062 & ~n8063;
  assign n8065 = pi29  & n7729;
  assign n8066 = ~n7734 & n8065;
  assign n8067 = n7734 & ~n8065;
  assign n8068 = ~n8066 & ~n8067;
  assign n8069 = ~n8064 & n8068;
  assign n8070 = ~n81 & ~n3427;
  assign n8071 = ~n3427 & n4600;
  assign n8072 = ~n3485 & n4615;
  assign n8073 = n4420 & ~n7720;
  assign n8074 = ~n8071 & ~n8072;
  assign n8075 = ~n8073 & n8074;
  assign n8076 = pi26  & ~n8070;
  assign n8077 = n8075 & n8076;
  assign n8078 = n86 & ~n3427;
  assign n8079 = n4420 & n7045;
  assign n8080 = ~n3485 & n4600;
  assign n8081 = ~n3370 & n4615;
  assign n8082 = ~n8078 & ~n8080;
  assign n8083 = ~n8081 & n8082;
  assign n8084 = ~n8079 & n8083;
  assign n8085 = n8077 & n8084;
  assign n8086 = n7729 & n8085;
  assign n8087 = ~n7729 & n8085;
  assign n8088 = n7729 & ~n8085;
  assign n8089 = ~n8087 & ~n8088;
  assign n8090 = ~n3275 & n4615;
  assign n8091 = n4420 & n7102;
  assign n8092 = n86 & ~n3485;
  assign n8093 = ~n3370 & n4600;
  assign n8094 = ~n8090 & ~n8092;
  assign n8095 = ~n8093 & n8094;
  assign n8096 = ~n8091 & n8095;
  assign n8097 = pi26  & n8096;
  assign n8098 = ~pi26  & ~n8096;
  assign n8099 = ~n8097 & ~n8098;
  assign n8100 = ~n8089 & ~n8099;
  assign n8101 = ~n8086 & ~n8100;
  assign n8102 = n8064 & ~n8068;
  assign n8103 = ~n8069 & ~n8102;
  assign n8104 = ~n8101 & n8103;
  assign n8105 = ~n8069 & ~n8104;
  assign n8106 = ~n8054 & ~n8105;
  assign n8107 = ~n8051 & ~n8106;
  assign n8108 = ~n8036 & ~n8107;
  assign n8109 = ~n8033 & ~n8108;
  assign n8110 = n8017 & n8019;
  assign n8111 = ~n8017 & ~n8019;
  assign n8112 = ~n8110 & ~n8111;
  assign n8113 = ~n8109 & ~n8112;
  assign n8114 = ~n8020 & ~n8113;
  assign n8115 = n7996 & n8006;
  assign n8116 = ~n7996 & ~n8006;
  assign n8117 = ~n8115 & ~n8116;
  assign n8118 = ~n8114 & ~n8117;
  assign n8119 = ~n8007 & ~n8118;
  assign n8120 = n7983 & n7993;
  assign n8121 = ~n7983 & ~n7993;
  assign n8122 = ~n8120 & ~n8121;
  assign n8123 = ~n8119 & ~n8122;
  assign n8124 = ~n7994 & ~n8123;
  assign n8125 = n7970 & n7980;
  assign n8126 = ~n7970 & ~n7980;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = ~n8124 & ~n8127;
  assign n8129 = ~n7981 & ~n8128;
  assign n8130 = n7957 & n7967;
  assign n8131 = ~n7957 & ~n7967;
  assign n8132 = ~n8130 & ~n8131;
  assign n8133 = ~n8129 & ~n8132;
  assign n8134 = ~n7968 & ~n8133;
  assign n8135 = n7944 & n7954;
  assign n8136 = ~n7944 & ~n7954;
  assign n8137 = ~n8135 & ~n8136;
  assign n8138 = ~n8134 & ~n8137;
  assign n8139 = ~n7955 & ~n8138;
  assign n8140 = n7931 & n7941;
  assign n8141 = ~n7931 & ~n7941;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = ~n8139 & ~n8142;
  assign n8144 = ~n7942 & ~n8143;
  assign n8145 = n7795 & ~n7797;
  assign n8146 = ~n7798 & ~n8145;
  assign n8147 = ~n8144 & n8146;
  assign n8148 = ~n2347 & n5130;
  assign n8149 = n5045 & n5596;
  assign n8150 = ~n2496 & n5044;
  assign n8151 = ~n2412 & n5109;
  assign n8152 = ~n8148 & ~n8150;
  assign n8153 = ~n8151 & n8152;
  assign n8154 = ~n8149 & n8153;
  assign n8155 = ~pi23  & ~n8154;
  assign n8156 = pi23  & n8154;
  assign n8157 = ~n8155 & ~n8156;
  assign n8158 = n8144 & ~n8146;
  assign n8159 = ~n8147 & ~n8158;
  assign n8160 = ~n8157 & n8159;
  assign n8161 = ~n8147 & ~n8160;
  assign n8162 = ~n7804 & ~n7805;
  assign n8163 = ~n7815 & n8162;
  assign n8164 = n7815 & ~n8162;
  assign n8165 = ~n8163 & ~n8164;
  assign n8166 = ~n8161 & n8165;
  assign n8167 = n8161 & ~n8165;
  assign n8168 = ~n2098 & n5853;
  assign n8169 = n4979 & n5241;
  assign n8170 = ~n2146 & n5240;
  assign n8171 = ~n1998 & n5866;
  assign n8172 = ~n8168 & ~n8170;
  assign n8173 = ~n8171 & n8172;
  assign n8174 = ~n8169 & n8173;
  assign n8175 = pi20  & n8174;
  assign n8176 = ~pi20  & ~n8174;
  assign n8177 = ~n8175 & ~n8176;
  assign n8178 = ~n8167 & ~n8177;
  assign n8179 = ~n8166 & ~n8178;
  assign n8180 = n7929 & ~n8179;
  assign n8181 = ~n7929 & n8179;
  assign n8182 = ~n1717 & n6323;
  assign n8183 = n4537 & n5983;
  assign n8184 = ~n1841 & n5982;
  assign n8185 = ~n1637 & n6336;
  assign n8186 = ~n8182 & ~n8184;
  assign n8187 = ~n8185 & n8186;
  assign n8188 = ~n8183 & n8187;
  assign n8189 = pi17  & n8188;
  assign n8190 = ~pi17  & ~n8188;
  assign n8191 = ~n8189 & ~n8190;
  assign n8192 = ~n8181 & ~n8191;
  assign n8193 = ~n8180 & ~n8192;
  assign n8194 = ~n7925 & ~n8193;
  assign n8195 = ~n7922 & ~n8194;
  assign n8196 = ~n7838 & ~n7839;
  assign n8197 = ~n7849 & n8196;
  assign n8198 = n7849 & ~n8196;
  assign n8199 = ~n8197 & ~n8198;
  assign n8200 = ~n8195 & n8199;
  assign n8201 = n8195 & ~n8199;
  assign n8202 = ~n1225 & n7238;
  assign n8203 = n4135 & n6631;
  assign n8204 = ~n1345 & n6630;
  assign n8205 = ~n1104 & n7262;
  assign n8206 = ~n8202 & ~n8204;
  assign n8207 = ~n8205 & n8206;
  assign n8208 = ~n8203 & n8207;
  assign n8209 = pi14  & n8208;
  assign n8210 = ~pi14  & ~n8208;
  assign n8211 = ~n8209 & ~n8210;
  assign n8212 = ~n8201 & ~n8211;
  assign n8213 = ~n8200 & ~n8212;
  assign n8214 = n7909 & ~n8213;
  assign n8215 = ~n7909 & n8213;
  assign n8216 = ~n3855 & n7895;
  assign n8217 = n3972 & n7431;
  assign n8218 = ~n987 & n7430;
  assign n8219 = ~n3681 & n7869;
  assign n8220 = ~n8216 & ~n8218;
  assign n8221 = ~n8219 & n8220;
  assign n8222 = ~n8217 & n8221;
  assign n8223 = pi11  & n8222;
  assign n8224 = ~pi11  & ~n8222;
  assign n8225 = ~n8223 & ~n8224;
  assign n8226 = ~n8215 & ~n8225;
  assign n8227 = ~n8214 & ~n8226;
  assign n8228 = ~n7905 & ~n8227;
  assign n8229 = n7905 & n8227;
  assign n8230 = n7596 & ~n7865;
  assign n8231 = ~n7596 & n7865;
  assign n8232 = ~n8230 & ~n8231;
  assign n8233 = ~n8229 & ~n8232;
  assign n8234 = ~n8228 & ~n8233;
  assign n8235 = n7894 & ~n8234;
  assign n8236 = ~n8228 & ~n8229;
  assign n8237 = ~n8232 & n8236;
  assign n8238 = n8232 & ~n8236;
  assign n8239 = ~n8237 & ~n8238;
  assign n8240 = pi7  & ~pi8 ;
  assign n8241 = ~pi7  & pi8 ;
  assign n8242 = ~n8240 & ~n8241;
  assign n8243 = pi5  & ~pi6 ;
  assign n8244 = ~pi5  & pi6 ;
  assign n8245 = ~n8243 & ~n8244;
  assign n8246 = ~pi6  & pi7 ;
  assign n8247 = pi6  & ~pi7 ;
  assign n8248 = ~n8246 & ~n8247;
  assign n8249 = n8245 & n8248;
  assign n8250 = ~n8242 & n8249;
  assign n8251 = ~n8242 & ~n8245;
  assign n8252 = ~n3897 & n8251;
  assign n8253 = ~n8250 & ~n8252;
  assign n8254 = ~n3883 & ~n8253;
  assign n8255 = pi8  & ~n8254;
  assign n8256 = ~pi8  & n8254;
  assign n8257 = ~n8255 & ~n8256;
  assign n8258 = n7925 & n8193;
  assign n8259 = ~n8194 & ~n8258;
  assign n8260 = ~n1345 & n7238;
  assign n8261 = n4152 & n6631;
  assign n8262 = ~n1448 & n6630;
  assign n8263 = ~n1225 & n7262;
  assign n8264 = ~n8260 & ~n8262;
  assign n8265 = ~n8263 & n8264;
  assign n8266 = ~n8261 & n8265;
  assign n8267 = pi14  & n8266;
  assign n8268 = ~pi14  & ~n8266;
  assign n8269 = ~n8267 & ~n8268;
  assign n8270 = n8259 & ~n8269;
  assign n8271 = ~n8259 & n8269;
  assign n8272 = ~n8270 & ~n8271;
  assign n8273 = ~n8180 & ~n8181;
  assign n8274 = ~n8191 & n8273;
  assign n8275 = n8191 & ~n8273;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = ~n2589 & n5044;
  assign n8278 = n5045 & n6016;
  assign n8279 = ~n2496 & n5109;
  assign n8280 = ~n2412 & n5130;
  assign n8281 = ~n8277 & ~n8279;
  assign n8282 = ~n8280 & n8281;
  assign n8283 = ~n8278 & n8282;
  assign n8284 = ~pi23  & ~n8283;
  assign n8285 = pi23  & n8283;
  assign n8286 = ~n8284 & ~n8285;
  assign n8287 = n8139 & n8142;
  assign n8288 = ~n8143 & ~n8287;
  assign n8289 = ~n8286 & n8288;
  assign n8290 = ~n8286 & ~n8288;
  assign n8291 = n8286 & n8288;
  assign n8292 = ~n8290 & ~n8291;
  assign n8293 = ~n2496 & n5130;
  assign n8294 = n5045 & n5776;
  assign n8295 = ~n2674 & n5044;
  assign n8296 = ~n2589 & n5109;
  assign n8297 = ~n8293 & ~n8295;
  assign n8298 = ~n8296 & n8297;
  assign n8299 = ~n8294 & n8298;
  assign n8300 = ~pi23  & ~n8299;
  assign n8301 = pi23  & n8299;
  assign n8302 = ~n8300 & ~n8301;
  assign n8303 = n8134 & n8137;
  assign n8304 = ~n8138 & ~n8303;
  assign n8305 = ~n8302 & n8304;
  assign n8306 = ~n8302 & ~n8304;
  assign n8307 = n8302 & n8304;
  assign n8308 = ~n8306 & ~n8307;
  assign n8309 = ~n2674 & n5109;
  assign n8310 = n5045 & n6240;
  assign n8311 = ~n2708 & n5044;
  assign n8312 = ~n2589 & n5130;
  assign n8313 = ~n8309 & ~n8311;
  assign n8314 = ~n8312 & n8313;
  assign n8315 = ~n8310 & n8314;
  assign n8316 = ~pi23  & ~n8315;
  assign n8317 = pi23  & n8315;
  assign n8318 = ~n8316 & ~n8317;
  assign n8319 = ~n8129 & n8132;
  assign n8320 = n8129 & ~n8132;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = ~n8318 & ~n8321;
  assign n8323 = ~n2778 & n5044;
  assign n8324 = n5045 & n6393;
  assign n8325 = ~n2708 & n5109;
  assign n8326 = ~n2674 & n5130;
  assign n8327 = ~n8323 & ~n8325;
  assign n8328 = ~n8326 & n8327;
  assign n8329 = ~n8324 & n8328;
  assign n8330 = ~pi23  & ~n8329;
  assign n8331 = pi23  & n8329;
  assign n8332 = ~n8330 & ~n8331;
  assign n8333 = ~n8124 & n8127;
  assign n8334 = n8124 & ~n8127;
  assign n8335 = ~n8333 & ~n8334;
  assign n8336 = ~n8332 & ~n8335;
  assign n8337 = ~n2708 & n5130;
  assign n8338 = n5045 & n6222;
  assign n8339 = ~n2835 & n5044;
  assign n8340 = ~n2778 & n5109;
  assign n8341 = ~n8337 & ~n8339;
  assign n8342 = ~n8340 & n8341;
  assign n8343 = ~n8338 & n8342;
  assign n8344 = ~pi23  & ~n8343;
  assign n8345 = pi23  & n8343;
  assign n8346 = ~n8344 & ~n8345;
  assign n8347 = n8119 & n8122;
  assign n8348 = ~n8123 & ~n8347;
  assign n8349 = ~n8346 & n8348;
  assign n8350 = ~n8346 & ~n8348;
  assign n8351 = n8346 & n8348;
  assign n8352 = ~n8350 & ~n8351;
  assign n8353 = ~n2919 & n5044;
  assign n8354 = n5045 & n6509;
  assign n8355 = ~n2835 & n5109;
  assign n8356 = ~n2778 & n5130;
  assign n8357 = ~n8353 & ~n8355;
  assign n8358 = ~n8356 & n8357;
  assign n8359 = ~n8354 & n8358;
  assign n8360 = ~pi23  & ~n8359;
  assign n8361 = pi23  & n8359;
  assign n8362 = ~n8360 & ~n8361;
  assign n8363 = n8114 & n8117;
  assign n8364 = ~n8118 & ~n8363;
  assign n8365 = ~n8362 & n8364;
  assign n8366 = ~n8362 & ~n8364;
  assign n8367 = n8362 & n8364;
  assign n8368 = ~n8366 & ~n8367;
  assign n8369 = ~n2919 & n5109;
  assign n8370 = n5045 & n6809;
  assign n8371 = ~n2951 & n5044;
  assign n8372 = ~n2835 & n5130;
  assign n8373 = ~n8369 & ~n8371;
  assign n8374 = ~n8372 & n8373;
  assign n8375 = ~n8370 & n8374;
  assign n8376 = ~pi23  & ~n8375;
  assign n8377 = pi23  & n8375;
  assign n8378 = ~n8376 & ~n8377;
  assign n8379 = ~n8109 & n8112;
  assign n8380 = n8109 & ~n8112;
  assign n8381 = ~n8379 & ~n8380;
  assign n8382 = ~n8378 & ~n8381;
  assign n8383 = n8036 & n8107;
  assign n8384 = ~n8108 & ~n8383;
  assign n8385 = ~n2919 & n5130;
  assign n8386 = n5045 & n6821;
  assign n8387 = ~n2951 & n5109;
  assign n8388 = ~n3031 & n5044;
  assign n8389 = ~n8385 & ~n8387;
  assign n8390 = ~n8388 & n8389;
  assign n8391 = ~n8386 & n8390;
  assign n8392 = pi23  & n8391;
  assign n8393 = ~pi23  & ~n8391;
  assign n8394 = ~n8392 & ~n8393;
  assign n8395 = n8384 & ~n8394;
  assign n8396 = n8054 & n8105;
  assign n8397 = ~n8106 & ~n8396;
  assign n8398 = ~n2951 & n5130;
  assign n8399 = n5045 & n6486;
  assign n8400 = ~n3118 & n5044;
  assign n8401 = ~n3031 & n5109;
  assign n8402 = ~n8398 & ~n8400;
  assign n8403 = ~n8401 & n8402;
  assign n8404 = ~n8399 & n8403;
  assign n8405 = pi23  & n8404;
  assign n8406 = ~pi23  & ~n8404;
  assign n8407 = ~n8405 & ~n8406;
  assign n8408 = n8397 & ~n8407;
  assign n8409 = ~n3182 & n5044;
  assign n8410 = n5045 & n6863;
  assign n8411 = ~n3118 & n5109;
  assign n8412 = ~n3031 & n5130;
  assign n8413 = ~n8409 & ~n8411;
  assign n8414 = ~n8412 & n8413;
  assign n8415 = ~n8410 & n8414;
  assign n8416 = ~pi23  & ~n8415;
  assign n8417 = pi23  & n8415;
  assign n8418 = ~n8416 & ~n8417;
  assign n8419 = n8101 & ~n8103;
  assign n8420 = ~n8104 & ~n8419;
  assign n8421 = ~n8418 & n8420;
  assign n8422 = ~n8418 & ~n8420;
  assign n8423 = n8418 & n8420;
  assign n8424 = ~n8422 & ~n8423;
  assign n8425 = ~n3118 & n5130;
  assign n8426 = n5045 & n6908;
  assign n8427 = ~n3241 & n5044;
  assign n8428 = ~n3182 & n5109;
  assign n8429 = ~n8425 & ~n8427;
  assign n8430 = ~n8428 & n8429;
  assign n8431 = ~n8426 & n8430;
  assign n8432 = pi23  & n8431;
  assign n8433 = ~pi23  & ~n8431;
  assign n8434 = ~n8432 & ~n8433;
  assign n8435 = n8089 & n8099;
  assign n8436 = ~n8100 & ~n8435;
  assign n8437 = ~n8434 & n8436;
  assign n8438 = ~n3275 & n5044;
  assign n8439 = n5045 & n6959;
  assign n8440 = ~n3241 & n5109;
  assign n8441 = ~n3182 & n5130;
  assign n8442 = ~n8438 & ~n8440;
  assign n8443 = ~n8441 & n8442;
  assign n8444 = ~n8439 & n8443;
  assign n8445 = ~pi23  & ~n8444;
  assign n8446 = pi23  & n8444;
  assign n8447 = ~n8445 & ~n8446;
  assign n8448 = pi26  & ~n8077;
  assign n8449 = n8084 & ~n8448;
  assign n8450 = ~n8084 & n8448;
  assign n8451 = ~n8449 & ~n8450;
  assign n8452 = ~n8447 & n8451;
  assign n8453 = ~n8447 & ~n8451;
  assign n8454 = n8447 & n8451;
  assign n8455 = ~n8453 & ~n8454;
  assign n8456 = ~n3241 & n5130;
  assign n8457 = n5045 & n7004;
  assign n8458 = ~n3275 & n5109;
  assign n8459 = ~n3370 & n5044;
  assign n8460 = ~n8456 & ~n8458;
  assign n8461 = ~n8459 & n8460;
  assign n8462 = ~n8457 & n8461;
  assign n8463 = pi23  & n8462;
  assign n8464 = ~pi23  & ~n8462;
  assign n8465 = ~n8463 & ~n8464;
  assign n8466 = pi26  & n8070;
  assign n8467 = ~n8075 & n8466;
  assign n8468 = n8075 & ~n8466;
  assign n8469 = ~n8467 & ~n8468;
  assign n8470 = ~n8465 & n8469;
  assign n8471 = ~n3427 & ~n5042;
  assign n8472 = ~n3427 & n5109;
  assign n8473 = ~n3485 & n5130;
  assign n8474 = n5045 & ~n7720;
  assign n8475 = ~n8472 & ~n8473;
  assign n8476 = ~n8474 & n8475;
  assign n8477 = pi23  & ~n8471;
  assign n8478 = n8476 & n8477;
  assign n8479 = ~n3427 & n5044;
  assign n8480 = n5045 & n7045;
  assign n8481 = ~n3485 & n5109;
  assign n8482 = ~n3370 & n5130;
  assign n8483 = ~n8479 & ~n8481;
  assign n8484 = ~n8482 & n8483;
  assign n8485 = ~n8480 & n8484;
  assign n8486 = n8478 & n8485;
  assign n8487 = n8070 & n8486;
  assign n8488 = ~n8070 & n8486;
  assign n8489 = n8070 & ~n8486;
  assign n8490 = ~n8488 & ~n8489;
  assign n8491 = ~n3275 & n5130;
  assign n8492 = n5045 & n7102;
  assign n8493 = ~n3485 & n5044;
  assign n8494 = ~n3370 & n5109;
  assign n8495 = ~n8491 & ~n8493;
  assign n8496 = ~n8494 & n8495;
  assign n8497 = ~n8492 & n8496;
  assign n8498 = pi23  & n8497;
  assign n8499 = ~pi23  & ~n8497;
  assign n8500 = ~n8498 & ~n8499;
  assign n8501 = ~n8490 & ~n8500;
  assign n8502 = ~n8487 & ~n8501;
  assign n8503 = n8465 & ~n8469;
  assign n8504 = ~n8470 & ~n8503;
  assign n8505 = ~n8502 & n8504;
  assign n8506 = ~n8470 & ~n8505;
  assign n8507 = ~n8455 & ~n8506;
  assign n8508 = ~n8452 & ~n8507;
  assign n8509 = n8434 & ~n8436;
  assign n8510 = ~n8437 & ~n8509;
  assign n8511 = ~n8508 & n8510;
  assign n8512 = ~n8437 & ~n8511;
  assign n8513 = ~n8424 & ~n8512;
  assign n8514 = ~n8421 & ~n8513;
  assign n8515 = n8397 & n8407;
  assign n8516 = ~n8397 & ~n8407;
  assign n8517 = ~n8515 & ~n8516;
  assign n8518 = ~n8514 & ~n8517;
  assign n8519 = ~n8408 & ~n8518;
  assign n8520 = ~n8384 & n8394;
  assign n8521 = ~n8395 & ~n8520;
  assign n8522 = ~n8519 & n8521;
  assign n8523 = ~n8395 & ~n8522;
  assign n8524 = n8378 & n8381;
  assign n8525 = ~n8382 & ~n8524;
  assign n8526 = ~n8523 & n8525;
  assign n8527 = ~n8382 & ~n8526;
  assign n8528 = ~n8368 & ~n8527;
  assign n8529 = ~n8365 & ~n8528;
  assign n8530 = ~n8352 & ~n8529;
  assign n8531 = ~n8349 & ~n8530;
  assign n8532 = n8332 & n8335;
  assign n8533 = ~n8336 & ~n8532;
  assign n8534 = ~n8531 & n8533;
  assign n8535 = ~n8336 & ~n8534;
  assign n8536 = n8318 & n8321;
  assign n8537 = ~n8322 & ~n8536;
  assign n8538 = ~n8535 & n8537;
  assign n8539 = ~n8322 & ~n8538;
  assign n8540 = ~n8308 & ~n8539;
  assign n8541 = ~n8305 & ~n8540;
  assign n8542 = ~n8292 & ~n8541;
  assign n8543 = ~n8289 & ~n8542;
  assign n8544 = n8157 & ~n8159;
  assign n8545 = ~n8160 & ~n8544;
  assign n8546 = ~n8543 & n8545;
  assign n8547 = ~n2098 & n5866;
  assign n8548 = n5241 & n5359;
  assign n8549 = ~n2146 & n5853;
  assign n8550 = ~n2249 & n5240;
  assign n8551 = ~n8547 & ~n8549;
  assign n8552 = ~n8550 & n8551;
  assign n8553 = ~n8548 & n8552;
  assign n8554 = ~pi20  & ~n8553;
  assign n8555 = pi20  & n8553;
  assign n8556 = ~n8554 & ~n8555;
  assign n8557 = n8543 & ~n8545;
  assign n8558 = ~n8546 & ~n8557;
  assign n8559 = ~n8556 & n8558;
  assign n8560 = ~n8546 & ~n8559;
  assign n8561 = ~n8166 & ~n8167;
  assign n8562 = ~n8177 & n8561;
  assign n8563 = n8177 & ~n8561;
  assign n8564 = ~n8562 & ~n8563;
  assign n8565 = ~n8560 & n8564;
  assign n8566 = n8560 & ~n8564;
  assign n8567 = ~n1841 & n6323;
  assign n8568 = n4762 & n5983;
  assign n8569 = ~n1908 & n5982;
  assign n8570 = ~n1717 & n6336;
  assign n8571 = ~n8567 & ~n8569;
  assign n8572 = ~n8570 & n8571;
  assign n8573 = ~n8568 & n8572;
  assign n8574 = pi17  & n8573;
  assign n8575 = ~pi17  & ~n8573;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = ~n8566 & ~n8576;
  assign n8578 = ~n8565 & ~n8577;
  assign n8579 = n8276 & ~n8578;
  assign n8580 = ~n8276 & n8578;
  assign n8581 = ~n1448 & n7238;
  assign n8582 = n4453 & n6631;
  assign n8583 = ~n1533 & n6630;
  assign n8584 = ~n1345 & n7262;
  assign n8585 = ~n8581 & ~n8583;
  assign n8586 = ~n8584 & n8585;
  assign n8587 = ~n8582 & n8586;
  assign n8588 = pi14  & n8587;
  assign n8589 = ~pi14  & ~n8587;
  assign n8590 = ~n8588 & ~n8589;
  assign n8591 = ~n8580 & ~n8590;
  assign n8592 = ~n8579 & ~n8591;
  assign n8593 = n8272 & ~n8592;
  assign n8594 = ~n8270 & ~n8593;
  assign n8595 = ~n8200 & ~n8201;
  assign n8596 = ~n8211 & n8595;
  assign n8597 = n8211 & ~n8595;
  assign n8598 = ~n8596 & ~n8597;
  assign n8599 = ~n8594 & n8598;
  assign n8600 = n8594 & ~n8598;
  assign n8601 = ~n878 & n7430;
  assign n8602 = n3687 & n7431;
  assign n8603 = ~n987 & n7869;
  assign n8604 = ~n3681 & n7895;
  assign n8605 = ~n8601 & ~n8603;
  assign n8606 = ~n8604 & n8605;
  assign n8607 = ~n8602 & n8606;
  assign n8608 = pi11  & n8607;
  assign n8609 = ~pi11  & ~n8607;
  assign n8610 = ~n8608 & ~n8609;
  assign n8611 = ~n8600 & ~n8610;
  assign n8612 = ~n8599 & ~n8611;
  assign n8613 = ~n8257 & ~n8612;
  assign n8614 = n8257 & n8612;
  assign n8615 = ~n8214 & ~n8215;
  assign n8616 = ~n8225 & n8615;
  assign n8617 = n8225 & ~n8615;
  assign n8618 = ~n8616 & ~n8617;
  assign n8619 = ~n8614 & n8618;
  assign n8620 = ~n8613 & ~n8619;
  assign n8621 = n8239 & ~n8620;
  assign n8622 = ~n8239 & n8620;
  assign n8623 = ~n8621 & ~n8622;
  assign n8624 = ~n987 & n7895;
  assign n8625 = n3791 & n7431;
  assign n8626 = ~n1104 & n7430;
  assign n8627 = ~n878 & n7869;
  assign n8628 = ~n8624 & ~n8626;
  assign n8629 = ~n8627 & n8628;
  assign n8630 = ~n8625 & n8629;
  assign n8631 = pi11  & n8630;
  assign n8632 = ~pi11  & ~n8630;
  assign n8633 = ~n8631 & ~n8632;
  assign n8634 = ~n8579 & ~n8580;
  assign n8635 = ~n8590 & n8634;
  assign n8636 = n8590 & ~n8634;
  assign n8637 = ~n8635 & ~n8636;
  assign n8638 = n8292 & n8541;
  assign n8639 = ~n8542 & ~n8638;
  assign n8640 = ~n2146 & n5866;
  assign n8641 = n5241 & n5343;
  assign n8642 = ~n2347 & n5240;
  assign n8643 = ~n2249 & n5853;
  assign n8644 = ~n8640 & ~n8642;
  assign n8645 = ~n8643 & n8644;
  assign n8646 = ~n8641 & n8645;
  assign n8647 = pi20  & n8646;
  assign n8648 = ~pi20  & ~n8646;
  assign n8649 = ~n8647 & ~n8648;
  assign n8650 = n8639 & ~n8649;
  assign n8651 = n8308 & n8539;
  assign n8652 = ~n8540 & ~n8651;
  assign n8653 = ~n2412 & n5240;
  assign n8654 = n5241 & n5579;
  assign n8655 = ~n2347 & n5853;
  assign n8656 = ~n2249 & n5866;
  assign n8657 = ~n8653 & ~n8655;
  assign n8658 = ~n8656 & n8657;
  assign n8659 = ~n8654 & n8658;
  assign n8660 = pi20  & n8659;
  assign n8661 = ~pi20  & ~n8659;
  assign n8662 = ~n8660 & ~n8661;
  assign n8663 = n8652 & ~n8662;
  assign n8664 = n8535 & ~n8537;
  assign n8665 = ~n8538 & ~n8664;
  assign n8666 = ~n2347 & n5866;
  assign n8667 = n5241 & n5596;
  assign n8668 = ~n2496 & n5240;
  assign n8669 = ~n2412 & n5853;
  assign n8670 = ~n8666 & ~n8668;
  assign n8671 = ~n8669 & n8670;
  assign n8672 = ~n8667 & n8671;
  assign n8673 = pi20  & n8672;
  assign n8674 = ~pi20  & ~n8672;
  assign n8675 = ~n8673 & ~n8674;
  assign n8676 = n8665 & ~n8675;
  assign n8677 = n8531 & ~n8533;
  assign n8678 = ~n8534 & ~n8677;
  assign n8679 = ~n2589 & n5240;
  assign n8680 = n5241 & n6016;
  assign n8681 = ~n2496 & n5853;
  assign n8682 = ~n2412 & n5866;
  assign n8683 = ~n8679 & ~n8681;
  assign n8684 = ~n8682 & n8683;
  assign n8685 = ~n8680 & n8684;
  assign n8686 = pi20  & n8685;
  assign n8687 = ~pi20  & ~n8685;
  assign n8688 = ~n8686 & ~n8687;
  assign n8689 = n8678 & ~n8688;
  assign n8690 = n8352 & n8529;
  assign n8691 = ~n8530 & ~n8690;
  assign n8692 = ~n2496 & n5866;
  assign n8693 = n5241 & n5776;
  assign n8694 = ~n2674 & n5240;
  assign n8695 = ~n2589 & n5853;
  assign n8696 = ~n8692 & ~n8694;
  assign n8697 = ~n8695 & n8696;
  assign n8698 = ~n8693 & n8697;
  assign n8699 = pi20  & n8698;
  assign n8700 = ~pi20  & ~n8698;
  assign n8701 = ~n8699 & ~n8700;
  assign n8702 = n8691 & ~n8701;
  assign n8703 = n8368 & n8527;
  assign n8704 = ~n8528 & ~n8703;
  assign n8705 = ~n2674 & n5853;
  assign n8706 = n5241 & n6240;
  assign n8707 = ~n2708 & n5240;
  assign n8708 = ~n2589 & n5866;
  assign n8709 = ~n8705 & ~n8707;
  assign n8710 = ~n8708 & n8709;
  assign n8711 = ~n8706 & n8710;
  assign n8712 = pi20  & n8711;
  assign n8713 = ~pi20  & ~n8711;
  assign n8714 = ~n8712 & ~n8713;
  assign n8715 = n8704 & ~n8714;
  assign n8716 = n8523 & ~n8525;
  assign n8717 = ~n8526 & ~n8716;
  assign n8718 = ~n2778 & n5240;
  assign n8719 = n5241 & n6393;
  assign n8720 = ~n2708 & n5853;
  assign n8721 = ~n2674 & n5866;
  assign n8722 = ~n8718 & ~n8720;
  assign n8723 = ~n8721 & n8722;
  assign n8724 = ~n8719 & n8723;
  assign n8725 = pi20  & n8724;
  assign n8726 = ~pi20  & ~n8724;
  assign n8727 = ~n8725 & ~n8726;
  assign n8728 = n8717 & ~n8727;
  assign n8729 = ~n2708 & n5866;
  assign n8730 = n5241 & n6222;
  assign n8731 = ~n2835 & n5240;
  assign n8732 = ~n2778 & n5853;
  assign n8733 = ~n8729 & ~n8731;
  assign n8734 = ~n8732 & n8733;
  assign n8735 = ~n8730 & n8734;
  assign n8736 = ~pi20  & ~n8735;
  assign n8737 = pi20  & n8735;
  assign n8738 = ~n8736 & ~n8737;
  assign n8739 = n8519 & ~n8521;
  assign n8740 = ~n8522 & ~n8739;
  assign n8741 = ~n8738 & n8740;
  assign n8742 = ~n8738 & ~n8740;
  assign n8743 = n8738 & n8740;
  assign n8744 = ~n8742 & ~n8743;
  assign n8745 = ~n2919 & n5240;
  assign n8746 = n5241 & n6509;
  assign n8747 = ~n2835 & n5853;
  assign n8748 = ~n2778 & n5866;
  assign n8749 = ~n8745 & ~n8747;
  assign n8750 = ~n8748 & n8749;
  assign n8751 = ~n8746 & n8750;
  assign n8752 = ~pi20  & ~n8751;
  assign n8753 = pi20  & n8751;
  assign n8754 = ~n8752 & ~n8753;
  assign n8755 = ~n8514 & n8517;
  assign n8756 = n8514 & ~n8517;
  assign n8757 = ~n8755 & ~n8756;
  assign n8758 = ~n8754 & ~n8757;
  assign n8759 = n8424 & n8512;
  assign n8760 = ~n8513 & ~n8759;
  assign n8761 = ~n2919 & n5853;
  assign n8762 = n5241 & n6809;
  assign n8763 = ~n2951 & n5240;
  assign n8764 = ~n2835 & n5866;
  assign n8765 = ~n8761 & ~n8763;
  assign n8766 = ~n8764 & n8765;
  assign n8767 = ~n8762 & n8766;
  assign n8768 = pi20  & n8767;
  assign n8769 = ~pi20  & ~n8767;
  assign n8770 = ~n8768 & ~n8769;
  assign n8771 = n8760 & ~n8770;
  assign n8772 = n8508 & ~n8510;
  assign n8773 = ~n8511 & ~n8772;
  assign n8774 = ~n2919 & n5866;
  assign n8775 = n5241 & n6821;
  assign n8776 = ~n2951 & n5853;
  assign n8777 = ~n3031 & n5240;
  assign n8778 = ~n8774 & ~n8776;
  assign n8779 = ~n8777 & n8778;
  assign n8780 = ~n8775 & n8779;
  assign n8781 = pi20  & n8780;
  assign n8782 = ~pi20  & ~n8780;
  assign n8783 = ~n8781 & ~n8782;
  assign n8784 = n8773 & ~n8783;
  assign n8785 = n8455 & n8506;
  assign n8786 = ~n8507 & ~n8785;
  assign n8787 = ~n2951 & n5866;
  assign n8788 = n5241 & n6486;
  assign n8789 = ~n3118 & n5240;
  assign n8790 = ~n3031 & n5853;
  assign n8791 = ~n8787 & ~n8789;
  assign n8792 = ~n8790 & n8791;
  assign n8793 = ~n8788 & n8792;
  assign n8794 = pi20  & n8793;
  assign n8795 = ~pi20  & ~n8793;
  assign n8796 = ~n8794 & ~n8795;
  assign n8797 = n8786 & ~n8796;
  assign n8798 = ~n3182 & n5240;
  assign n8799 = n5241 & n6863;
  assign n8800 = ~n3118 & n5853;
  assign n8801 = ~n3031 & n5866;
  assign n8802 = ~n8798 & ~n8800;
  assign n8803 = ~n8801 & n8802;
  assign n8804 = ~n8799 & n8803;
  assign n8805 = ~pi20  & ~n8804;
  assign n8806 = pi20  & n8804;
  assign n8807 = ~n8805 & ~n8806;
  assign n8808 = n8502 & ~n8504;
  assign n8809 = ~n8505 & ~n8808;
  assign n8810 = ~n8807 & n8809;
  assign n8811 = ~n8807 & ~n8809;
  assign n8812 = n8807 & n8809;
  assign n8813 = ~n8811 & ~n8812;
  assign n8814 = ~n3118 & n5866;
  assign n8815 = n5241 & n6908;
  assign n8816 = ~n3241 & n5240;
  assign n8817 = ~n3182 & n5853;
  assign n8818 = ~n8814 & ~n8816;
  assign n8819 = ~n8817 & n8818;
  assign n8820 = ~n8815 & n8819;
  assign n8821 = pi20  & n8820;
  assign n8822 = ~pi20  & ~n8820;
  assign n8823 = ~n8821 & ~n8822;
  assign n8824 = n8490 & n8500;
  assign n8825 = ~n8501 & ~n8824;
  assign n8826 = ~n8823 & n8825;
  assign n8827 = ~n3275 & n5240;
  assign n8828 = n5241 & n6959;
  assign n8829 = ~n3241 & n5853;
  assign n8830 = ~n3182 & n5866;
  assign n8831 = ~n8827 & ~n8829;
  assign n8832 = ~n8830 & n8831;
  assign n8833 = ~n8828 & n8832;
  assign n8834 = ~pi20  & ~n8833;
  assign n8835 = pi20  & n8833;
  assign n8836 = ~n8834 & ~n8835;
  assign n8837 = pi23  & ~n8478;
  assign n8838 = n8485 & ~n8837;
  assign n8839 = ~n8485 & n8837;
  assign n8840 = ~n8838 & ~n8839;
  assign n8841 = ~n8836 & n8840;
  assign n8842 = ~n8836 & ~n8840;
  assign n8843 = n8836 & n8840;
  assign n8844 = ~n8842 & ~n8843;
  assign n8845 = ~n3241 & n5866;
  assign n8846 = n5241 & n7004;
  assign n8847 = ~n3275 & n5853;
  assign n8848 = ~n3370 & n5240;
  assign n8849 = ~n8845 & ~n8847;
  assign n8850 = ~n8848 & n8849;
  assign n8851 = ~n8846 & n8850;
  assign n8852 = pi20  & n8851;
  assign n8853 = ~pi20  & ~n8851;
  assign n8854 = ~n8852 & ~n8853;
  assign n8855 = pi23  & n8471;
  assign n8856 = ~n8476 & n8855;
  assign n8857 = n8476 & ~n8855;
  assign n8858 = ~n8856 & ~n8857;
  assign n8859 = ~n8854 & n8858;
  assign n8860 = ~n3427 & ~n5235;
  assign n8861 = ~n3427 & n5853;
  assign n8862 = ~n3485 & n5866;
  assign n8863 = n5241 & ~n7720;
  assign n8864 = ~n8861 & ~n8862;
  assign n8865 = ~n8863 & n8864;
  assign n8866 = pi20  & ~n8860;
  assign n8867 = n8865 & n8866;
  assign n8868 = ~n3427 & n5240;
  assign n8869 = n5241 & n7045;
  assign n8870 = ~n3485 & n5853;
  assign n8871 = ~n3370 & n5866;
  assign n8872 = ~n8868 & ~n8870;
  assign n8873 = ~n8871 & n8872;
  assign n8874 = ~n8869 & n8873;
  assign n8875 = n8867 & n8874;
  assign n8876 = n8471 & n8875;
  assign n8877 = ~n8471 & n8875;
  assign n8878 = n8471 & ~n8875;
  assign n8879 = ~n8877 & ~n8878;
  assign n8880 = ~n3275 & n5866;
  assign n8881 = n5241 & n7102;
  assign n8882 = ~n3485 & n5240;
  assign n8883 = ~n3370 & n5853;
  assign n8884 = ~n8880 & ~n8882;
  assign n8885 = ~n8883 & n8884;
  assign n8886 = ~n8881 & n8885;
  assign n8887 = pi20  & n8886;
  assign n8888 = ~pi20  & ~n8886;
  assign n8889 = ~n8887 & ~n8888;
  assign n8890 = ~n8879 & ~n8889;
  assign n8891 = ~n8876 & ~n8890;
  assign n8892 = n8854 & ~n8858;
  assign n8893 = ~n8859 & ~n8892;
  assign n8894 = ~n8891 & n8893;
  assign n8895 = ~n8859 & ~n8894;
  assign n8896 = ~n8844 & ~n8895;
  assign n8897 = ~n8841 & ~n8896;
  assign n8898 = n8823 & ~n8825;
  assign n8899 = ~n8826 & ~n8898;
  assign n8900 = ~n8897 & n8899;
  assign n8901 = ~n8826 & ~n8900;
  assign n8902 = ~n8813 & ~n8901;
  assign n8903 = ~n8810 & ~n8902;
  assign n8904 = n8786 & n8796;
  assign n8905 = ~n8786 & ~n8796;
  assign n8906 = ~n8904 & ~n8905;
  assign n8907 = ~n8903 & ~n8906;
  assign n8908 = ~n8797 & ~n8907;
  assign n8909 = n8773 & n8783;
  assign n8910 = ~n8773 & ~n8783;
  assign n8911 = ~n8909 & ~n8910;
  assign n8912 = ~n8908 & ~n8911;
  assign n8913 = ~n8784 & ~n8912;
  assign n8914 = ~n8760 & n8770;
  assign n8915 = ~n8771 & ~n8914;
  assign n8916 = ~n8913 & n8915;
  assign n8917 = ~n8771 & ~n8916;
  assign n8918 = n8754 & n8757;
  assign n8919 = ~n8758 & ~n8918;
  assign n8920 = ~n8917 & n8919;
  assign n8921 = ~n8758 & ~n8920;
  assign n8922 = ~n8744 & ~n8921;
  assign n8923 = ~n8741 & ~n8922;
  assign n8924 = n8717 & n8727;
  assign n8925 = ~n8717 & ~n8727;
  assign n8926 = ~n8924 & ~n8925;
  assign n8927 = ~n8923 & ~n8926;
  assign n8928 = ~n8728 & ~n8927;
  assign n8929 = n8704 & n8714;
  assign n8930 = ~n8704 & ~n8714;
  assign n8931 = ~n8929 & ~n8930;
  assign n8932 = ~n8928 & ~n8931;
  assign n8933 = ~n8715 & ~n8932;
  assign n8934 = n8691 & n8701;
  assign n8935 = ~n8691 & ~n8701;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = ~n8933 & ~n8936;
  assign n8938 = ~n8702 & ~n8937;
  assign n8939 = n8678 & n8688;
  assign n8940 = ~n8678 & ~n8688;
  assign n8941 = ~n8939 & ~n8940;
  assign n8942 = ~n8938 & ~n8941;
  assign n8943 = ~n8689 & ~n8942;
  assign n8944 = n8665 & n8675;
  assign n8945 = ~n8665 & ~n8675;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = ~n8943 & ~n8946;
  assign n8948 = ~n8676 & ~n8947;
  assign n8949 = n8652 & n8662;
  assign n8950 = ~n8652 & ~n8662;
  assign n8951 = ~n8949 & ~n8950;
  assign n8952 = ~n8948 & ~n8951;
  assign n8953 = ~n8663 & ~n8952;
  assign n8954 = n8639 & n8649;
  assign n8955 = ~n8639 & ~n8649;
  assign n8956 = ~n8954 & ~n8955;
  assign n8957 = ~n8953 & ~n8956;
  assign n8958 = ~n8650 & ~n8957;
  assign n8959 = n8556 & ~n8558;
  assign n8960 = ~n8559 & ~n8959;
  assign n8961 = ~n8958 & n8960;
  assign n8962 = ~n1908 & n6323;
  assign n8963 = n4779 & n5983;
  assign n8964 = ~n1998 & n5982;
  assign n8965 = ~n1841 & n6336;
  assign n8966 = ~n8962 & ~n8964;
  assign n8967 = ~n8965 & n8966;
  assign n8968 = ~n8963 & n8967;
  assign n8969 = ~pi17  & ~n8968;
  assign n8970 = pi17  & n8968;
  assign n8971 = ~n8969 & ~n8970;
  assign n8972 = n8958 & ~n8960;
  assign n8973 = ~n8961 & ~n8972;
  assign n8974 = ~n8971 & n8973;
  assign n8975 = ~n8961 & ~n8974;
  assign n8976 = ~n8565 & ~n8566;
  assign n8977 = ~n8576 & n8976;
  assign n8978 = n8576 & ~n8976;
  assign n8979 = ~n8977 & ~n8978;
  assign n8980 = ~n8975 & n8979;
  assign n8981 = n8975 & ~n8979;
  assign n8982 = ~n1533 & n7238;
  assign n8983 = n4355 & n6631;
  assign n8984 = ~n1637 & n6630;
  assign n8985 = ~n1448 & n7262;
  assign n8986 = ~n8982 & ~n8984;
  assign n8987 = ~n8985 & n8986;
  assign n8988 = ~n8983 & n8987;
  assign n8989 = pi14  & n8988;
  assign n8990 = ~pi14  & ~n8988;
  assign n8991 = ~n8989 & ~n8990;
  assign n8992 = ~n8981 & ~n8991;
  assign n8993 = ~n8980 & ~n8992;
  assign n8994 = n8637 & ~n8993;
  assign n8995 = ~n8637 & n8993;
  assign n8996 = ~n1104 & n7869;
  assign n8997 = n3775 & n7431;
  assign n8998 = ~n1225 & n7430;
  assign n8999 = ~n878 & n7895;
  assign n9000 = ~n8996 & ~n8998;
  assign n9001 = ~n8999 & n9000;
  assign n9002 = ~n8997 & n9001;
  assign n9003 = pi11  & n9002;
  assign n9004 = ~pi11  & ~n9002;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = ~n8995 & ~n9005;
  assign n9007 = ~n8994 & ~n9006;
  assign n9008 = ~n8633 & ~n9007;
  assign n9009 = n8633 & n9007;
  assign n9010 = ~n9008 & ~n9009;
  assign n9011 = ~n8272 & n8592;
  assign n9012 = ~n8593 & ~n9011;
  assign n9013 = n9010 & n9012;
  assign n9014 = ~n9008 & ~n9013;
  assign n9015 = ~n3855 & n8250;
  assign n9016 = n8245 & ~n8248;
  assign n9017 = ~n3883 & n9016;
  assign n9018 = ~n3900 & n8251;
  assign n9019 = ~n9015 & ~n9017;
  assign n9020 = ~n9018 & n9019;
  assign n9021 = pi8  & n9020;
  assign n9022 = ~pi8  & ~n9020;
  assign n9023 = ~n9021 & ~n9022;
  assign n9024 = ~n9014 & ~n9023;
  assign n9025 = n9014 & n9023;
  assign n9026 = ~n9024 & ~n9025;
  assign n9027 = ~n8599 & ~n8600;
  assign n9028 = ~n8610 & n9027;
  assign n9029 = n8610 & ~n9027;
  assign n9030 = ~n9028 & ~n9029;
  assign n9031 = n9026 & n9030;
  assign n9032 = ~n9024 & ~n9031;
  assign n9033 = ~n8613 & ~n8614;
  assign n9034 = n8618 & n9033;
  assign n9035 = ~n8618 & ~n9033;
  assign n9036 = ~n9034 & ~n9035;
  assign n9037 = ~n9032 & n9036;
  assign n9038 = n9032 & ~n9036;
  assign n9039 = ~n9037 & ~n9038;
  assign n9040 = n8242 & ~n8245;
  assign n9041 = ~n3883 & n9040;
  assign n9042 = n4399 & n8251;
  assign n9043 = ~n3855 & n9016;
  assign n9044 = ~n3681 & n8250;
  assign n9045 = ~n9041 & ~n9043;
  assign n9046 = ~n9044 & n9045;
  assign n9047 = ~n9042 & n9046;
  assign n9048 = pi8  & n9047;
  assign n9049 = ~pi8  & ~n9047;
  assign n9050 = ~n9048 & ~n9049;
  assign n9051 = ~n8994 & ~n8995;
  assign n9052 = ~n9005 & n9051;
  assign n9053 = n9005 & ~n9051;
  assign n9054 = ~n9052 & ~n9053;
  assign n9055 = ~n1998 & n6323;
  assign n9056 = n5151 & n5983;
  assign n9057 = ~n2098 & n5982;
  assign n9058 = ~n1908 & n6336;
  assign n9059 = ~n9055 & ~n9057;
  assign n9060 = ~n9058 & n9059;
  assign n9061 = ~n9056 & n9060;
  assign n9062 = ~pi17  & ~n9061;
  assign n9063 = pi17  & n9061;
  assign n9064 = ~n9062 & ~n9063;
  assign n9065 = ~n8953 & n8956;
  assign n9066 = n8953 & ~n8956;
  assign n9067 = ~n9065 & ~n9066;
  assign n9068 = ~n9064 & ~n9067;
  assign n9069 = ~n2098 & n6323;
  assign n9070 = n4979 & n5983;
  assign n9071 = ~n2146 & n5982;
  assign n9072 = ~n1998 & n6336;
  assign n9073 = ~n9069 & ~n9071;
  assign n9074 = ~n9072 & n9073;
  assign n9075 = ~n9070 & n9074;
  assign n9076 = ~pi17  & ~n9075;
  assign n9077 = pi17  & n9075;
  assign n9078 = ~n9076 & ~n9077;
  assign n9079 = ~n8948 & n8951;
  assign n9080 = n8948 & ~n8951;
  assign n9081 = ~n9079 & ~n9080;
  assign n9082 = ~n9078 & ~n9081;
  assign n9083 = ~n2098 & n6336;
  assign n9084 = n5359 & n5983;
  assign n9085 = ~n2146 & n6323;
  assign n9086 = ~n2249 & n5982;
  assign n9087 = ~n9083 & ~n9085;
  assign n9088 = ~n9086 & n9087;
  assign n9089 = ~n9084 & n9088;
  assign n9090 = ~pi17  & ~n9089;
  assign n9091 = pi17  & n9089;
  assign n9092 = ~n9090 & ~n9091;
  assign n9093 = n8943 & n8946;
  assign n9094 = ~n8947 & ~n9093;
  assign n9095 = ~n9092 & n9094;
  assign n9096 = ~n9092 & ~n9094;
  assign n9097 = n9092 & n9094;
  assign n9098 = ~n9096 & ~n9097;
  assign n9099 = ~n2146 & n6336;
  assign n9100 = n5343 & n5983;
  assign n9101 = ~n2347 & n5982;
  assign n9102 = ~n2249 & n6323;
  assign n9103 = ~n9099 & ~n9101;
  assign n9104 = ~n9102 & n9103;
  assign n9105 = ~n9100 & n9104;
  assign n9106 = ~pi17  & ~n9105;
  assign n9107 = pi17  & n9105;
  assign n9108 = ~n9106 & ~n9107;
  assign n9109 = n8938 & n8941;
  assign n9110 = ~n8942 & ~n9109;
  assign n9111 = ~n9108 & n9110;
  assign n9112 = ~n9108 & ~n9110;
  assign n9113 = n9108 & n9110;
  assign n9114 = ~n9112 & ~n9113;
  assign n9115 = ~n2412 & n5982;
  assign n9116 = n5579 & n5983;
  assign n9117 = ~n2347 & n6323;
  assign n9118 = ~n2249 & n6336;
  assign n9119 = ~n9115 & ~n9117;
  assign n9120 = ~n9118 & n9119;
  assign n9121 = ~n9116 & n9120;
  assign n9122 = ~pi17  & ~n9121;
  assign n9123 = pi17  & n9121;
  assign n9124 = ~n9122 & ~n9123;
  assign n9125 = ~n8933 & n8936;
  assign n9126 = n8933 & ~n8936;
  assign n9127 = ~n9125 & ~n9126;
  assign n9128 = ~n9124 & ~n9127;
  assign n9129 = ~n2347 & n6336;
  assign n9130 = n5596 & n5983;
  assign n9131 = ~n2496 & n5982;
  assign n9132 = ~n2412 & n6323;
  assign n9133 = ~n9129 & ~n9131;
  assign n9134 = ~n9132 & n9133;
  assign n9135 = ~n9130 & n9134;
  assign n9136 = ~pi17  & ~n9135;
  assign n9137 = pi17  & n9135;
  assign n9138 = ~n9136 & ~n9137;
  assign n9139 = ~n8928 & n8931;
  assign n9140 = n8928 & ~n8931;
  assign n9141 = ~n9139 & ~n9140;
  assign n9142 = ~n9138 & ~n9141;
  assign n9143 = ~n2589 & n5982;
  assign n9144 = n5983 & n6016;
  assign n9145 = ~n2496 & n6323;
  assign n9146 = ~n2412 & n6336;
  assign n9147 = ~n9143 & ~n9145;
  assign n9148 = ~n9146 & n9147;
  assign n9149 = ~n9144 & n9148;
  assign n9150 = ~pi17  & ~n9149;
  assign n9151 = pi17  & n9149;
  assign n9152 = ~n9150 & ~n9151;
  assign n9153 = n8923 & n8926;
  assign n9154 = ~n8927 & ~n9153;
  assign n9155 = ~n9152 & n9154;
  assign n9156 = ~n9152 & ~n9154;
  assign n9157 = n9152 & n9154;
  assign n9158 = ~n9156 & ~n9157;
  assign n9159 = n8744 & n8921;
  assign n9160 = ~n8922 & ~n9159;
  assign n9161 = ~n2496 & n6336;
  assign n9162 = n5776 & n5983;
  assign n9163 = ~n2674 & n5982;
  assign n9164 = ~n2589 & n6323;
  assign n9165 = ~n9161 & ~n9163;
  assign n9166 = ~n9164 & n9165;
  assign n9167 = ~n9162 & n9166;
  assign n9168 = pi17  & n9167;
  assign n9169 = ~pi17  & ~n9167;
  assign n9170 = ~n9168 & ~n9169;
  assign n9171 = n9160 & ~n9170;
  assign n9172 = n8917 & ~n8919;
  assign n9173 = ~n8920 & ~n9172;
  assign n9174 = ~n2674 & n6323;
  assign n9175 = n5983 & n6240;
  assign n9176 = ~n2708 & n5982;
  assign n9177 = ~n2589 & n6336;
  assign n9178 = ~n9174 & ~n9176;
  assign n9179 = ~n9177 & n9178;
  assign n9180 = ~n9175 & n9179;
  assign n9181 = pi17  & n9180;
  assign n9182 = ~pi17  & ~n9180;
  assign n9183 = ~n9181 & ~n9182;
  assign n9184 = n9173 & ~n9183;
  assign n9185 = ~n2778 & n5982;
  assign n9186 = n5983 & n6393;
  assign n9187 = ~n2708 & n6323;
  assign n9188 = ~n2674 & n6336;
  assign n9189 = ~n9185 & ~n9187;
  assign n9190 = ~n9188 & n9189;
  assign n9191 = ~n9186 & n9190;
  assign n9192 = ~pi17  & ~n9191;
  assign n9193 = pi17  & n9191;
  assign n9194 = ~n9192 & ~n9193;
  assign n9195 = n8913 & ~n8915;
  assign n9196 = ~n8916 & ~n9195;
  assign n9197 = ~n9194 & n9196;
  assign n9198 = ~n9194 & ~n9196;
  assign n9199 = n9194 & n9196;
  assign n9200 = ~n9198 & ~n9199;
  assign n9201 = ~n2708 & n6336;
  assign n9202 = n5983 & n6222;
  assign n9203 = ~n2835 & n5982;
  assign n9204 = ~n2778 & n6323;
  assign n9205 = ~n9201 & ~n9203;
  assign n9206 = ~n9204 & n9205;
  assign n9207 = ~n9202 & n9206;
  assign n9208 = ~pi17  & ~n9207;
  assign n9209 = pi17  & n9207;
  assign n9210 = ~n9208 & ~n9209;
  assign n9211 = n8908 & n8911;
  assign n9212 = ~n8912 & ~n9211;
  assign n9213 = ~n9210 & n9212;
  assign n9214 = ~n9210 & ~n9212;
  assign n9215 = n9210 & n9212;
  assign n9216 = ~n9214 & ~n9215;
  assign n9217 = ~n2919 & n5982;
  assign n9218 = n5983 & n6509;
  assign n9219 = ~n2835 & n6323;
  assign n9220 = ~n2778 & n6336;
  assign n9221 = ~n9217 & ~n9219;
  assign n9222 = ~n9220 & n9221;
  assign n9223 = ~n9218 & n9222;
  assign n9224 = ~pi17  & ~n9223;
  assign n9225 = pi17  & n9223;
  assign n9226 = ~n9224 & ~n9225;
  assign n9227 = ~n8903 & n8906;
  assign n9228 = n8903 & ~n8906;
  assign n9229 = ~n9227 & ~n9228;
  assign n9230 = ~n9226 & ~n9229;
  assign n9231 = n8813 & n8901;
  assign n9232 = ~n8902 & ~n9231;
  assign n9233 = ~n2919 & n6323;
  assign n9234 = n5983 & n6809;
  assign n9235 = ~n2951 & n5982;
  assign n9236 = ~n2835 & n6336;
  assign n9237 = ~n9233 & ~n9235;
  assign n9238 = ~n9236 & n9237;
  assign n9239 = ~n9234 & n9238;
  assign n9240 = pi17  & n9239;
  assign n9241 = ~pi17  & ~n9239;
  assign n9242 = ~n9240 & ~n9241;
  assign n9243 = n9232 & ~n9242;
  assign n9244 = n8897 & ~n8899;
  assign n9245 = ~n8900 & ~n9244;
  assign n9246 = ~n2919 & n6336;
  assign n9247 = n5983 & n6821;
  assign n9248 = ~n2951 & n6323;
  assign n9249 = ~n3031 & n5982;
  assign n9250 = ~n9246 & ~n9248;
  assign n9251 = ~n9249 & n9250;
  assign n9252 = ~n9247 & n9251;
  assign n9253 = pi17  & n9252;
  assign n9254 = ~pi17  & ~n9252;
  assign n9255 = ~n9253 & ~n9254;
  assign n9256 = n9245 & ~n9255;
  assign n9257 = n8844 & n8895;
  assign n9258 = ~n8896 & ~n9257;
  assign n9259 = ~n2951 & n6336;
  assign n9260 = n5983 & n6486;
  assign n9261 = ~n3118 & n5982;
  assign n9262 = ~n3031 & n6323;
  assign n9263 = ~n9259 & ~n9261;
  assign n9264 = ~n9262 & n9263;
  assign n9265 = ~n9260 & n9264;
  assign n9266 = pi17  & n9265;
  assign n9267 = ~pi17  & ~n9265;
  assign n9268 = ~n9266 & ~n9267;
  assign n9269 = n9258 & ~n9268;
  assign n9270 = ~n3182 & n5982;
  assign n9271 = n5983 & n6863;
  assign n9272 = ~n3118 & n6323;
  assign n9273 = ~n3031 & n6336;
  assign n9274 = ~n9270 & ~n9272;
  assign n9275 = ~n9273 & n9274;
  assign n9276 = ~n9271 & n9275;
  assign n9277 = ~pi17  & ~n9276;
  assign n9278 = pi17  & n9276;
  assign n9279 = ~n9277 & ~n9278;
  assign n9280 = n8891 & ~n8893;
  assign n9281 = ~n8894 & ~n9280;
  assign n9282 = ~n9279 & n9281;
  assign n9283 = ~n9279 & ~n9281;
  assign n9284 = n9279 & n9281;
  assign n9285 = ~n9283 & ~n9284;
  assign n9286 = ~n3118 & n6336;
  assign n9287 = n5983 & n6908;
  assign n9288 = ~n3241 & n5982;
  assign n9289 = ~n3182 & n6323;
  assign n9290 = ~n9286 & ~n9288;
  assign n9291 = ~n9289 & n9290;
  assign n9292 = ~n9287 & n9291;
  assign n9293 = pi17  & n9292;
  assign n9294 = ~pi17  & ~n9292;
  assign n9295 = ~n9293 & ~n9294;
  assign n9296 = n8879 & n8889;
  assign n9297 = ~n8890 & ~n9296;
  assign n9298 = ~n9295 & n9297;
  assign n9299 = ~n3275 & n5982;
  assign n9300 = n5983 & n6959;
  assign n9301 = ~n3241 & n6323;
  assign n9302 = ~n3182 & n6336;
  assign n9303 = ~n9299 & ~n9301;
  assign n9304 = ~n9302 & n9303;
  assign n9305 = ~n9300 & n9304;
  assign n9306 = ~pi17  & ~n9305;
  assign n9307 = pi17  & n9305;
  assign n9308 = ~n9306 & ~n9307;
  assign n9309 = pi20  & ~n8867;
  assign n9310 = n8874 & ~n9309;
  assign n9311 = ~n8874 & n9309;
  assign n9312 = ~n9310 & ~n9311;
  assign n9313 = ~n9308 & n9312;
  assign n9314 = ~n9308 & ~n9312;
  assign n9315 = n9308 & n9312;
  assign n9316 = ~n9314 & ~n9315;
  assign n9317 = ~n3241 & n6336;
  assign n9318 = n5983 & n7004;
  assign n9319 = ~n3275 & n6323;
  assign n9320 = ~n3370 & n5982;
  assign n9321 = ~n9317 & ~n9319;
  assign n9322 = ~n9320 & n9321;
  assign n9323 = ~n9318 & n9322;
  assign n9324 = pi17  & n9323;
  assign n9325 = ~pi17  & ~n9323;
  assign n9326 = ~n9324 & ~n9325;
  assign n9327 = pi20  & n8860;
  assign n9328 = ~n8865 & n9327;
  assign n9329 = n8865 & ~n9327;
  assign n9330 = ~n9328 & ~n9329;
  assign n9331 = ~n9326 & n9330;
  assign n9332 = ~n3427 & ~n5980;
  assign n9333 = ~n3427 & n6323;
  assign n9334 = ~n3485 & n6336;
  assign n9335 = n5983 & ~n7720;
  assign n9336 = ~n9333 & ~n9334;
  assign n9337 = ~n9335 & n9336;
  assign n9338 = pi17  & ~n9332;
  assign n9339 = n9337 & n9338;
  assign n9340 = ~n3427 & n5982;
  assign n9341 = n5983 & n7045;
  assign n9342 = ~n3485 & n6323;
  assign n9343 = ~n3370 & n6336;
  assign n9344 = ~n9340 & ~n9342;
  assign n9345 = ~n9343 & n9344;
  assign n9346 = ~n9341 & n9345;
  assign n9347 = n9339 & n9346;
  assign n9348 = n8860 & n9347;
  assign n9349 = ~n8860 & n9347;
  assign n9350 = n8860 & ~n9347;
  assign n9351 = ~n9349 & ~n9350;
  assign n9352 = ~n3275 & n6336;
  assign n9353 = n5983 & n7102;
  assign n9354 = ~n3485 & n5982;
  assign n9355 = ~n3370 & n6323;
  assign n9356 = ~n9352 & ~n9354;
  assign n9357 = ~n9355 & n9356;
  assign n9358 = ~n9353 & n9357;
  assign n9359 = pi17  & n9358;
  assign n9360 = ~pi17  & ~n9358;
  assign n9361 = ~n9359 & ~n9360;
  assign n9362 = ~n9351 & ~n9361;
  assign n9363 = ~n9348 & ~n9362;
  assign n9364 = n9326 & ~n9330;
  assign n9365 = ~n9331 & ~n9364;
  assign n9366 = ~n9363 & n9365;
  assign n9367 = ~n9331 & ~n9366;
  assign n9368 = ~n9316 & ~n9367;
  assign n9369 = ~n9313 & ~n9368;
  assign n9370 = n9295 & ~n9297;
  assign n9371 = ~n9298 & ~n9370;
  assign n9372 = ~n9369 & n9371;
  assign n9373 = ~n9298 & ~n9372;
  assign n9374 = ~n9285 & ~n9373;
  assign n9375 = ~n9282 & ~n9374;
  assign n9376 = n9258 & n9268;
  assign n9377 = ~n9258 & ~n9268;
  assign n9378 = ~n9376 & ~n9377;
  assign n9379 = ~n9375 & ~n9378;
  assign n9380 = ~n9269 & ~n9379;
  assign n9381 = n9245 & n9255;
  assign n9382 = ~n9245 & ~n9255;
  assign n9383 = ~n9381 & ~n9382;
  assign n9384 = ~n9380 & ~n9383;
  assign n9385 = ~n9256 & ~n9384;
  assign n9386 = ~n9232 & n9242;
  assign n9387 = ~n9243 & ~n9386;
  assign n9388 = ~n9385 & n9387;
  assign n9389 = ~n9243 & ~n9388;
  assign n9390 = n9226 & n9229;
  assign n9391 = ~n9230 & ~n9390;
  assign n9392 = ~n9389 & n9391;
  assign n9393 = ~n9230 & ~n9392;
  assign n9394 = ~n9216 & ~n9393;
  assign n9395 = ~n9213 & ~n9394;
  assign n9396 = ~n9200 & ~n9395;
  assign n9397 = ~n9197 & ~n9396;
  assign n9398 = n9173 & n9183;
  assign n9399 = ~n9173 & ~n9183;
  assign n9400 = ~n9398 & ~n9399;
  assign n9401 = ~n9397 & ~n9400;
  assign n9402 = ~n9184 & ~n9401;
  assign n9403 = ~n9160 & n9170;
  assign n9404 = ~n9171 & ~n9403;
  assign n9405 = ~n9402 & n9404;
  assign n9406 = ~n9171 & ~n9405;
  assign n9407 = ~n9158 & ~n9406;
  assign n9408 = ~n9155 & ~n9407;
  assign n9409 = n9138 & n9141;
  assign n9410 = ~n9142 & ~n9409;
  assign n9411 = ~n9408 & n9410;
  assign n9412 = ~n9142 & ~n9411;
  assign n9413 = n9124 & n9127;
  assign n9414 = ~n9128 & ~n9413;
  assign n9415 = ~n9412 & n9414;
  assign n9416 = ~n9128 & ~n9415;
  assign n9417 = ~n9114 & ~n9416;
  assign n9418 = ~n9111 & ~n9417;
  assign n9419 = ~n9098 & ~n9418;
  assign n9420 = ~n9095 & ~n9419;
  assign n9421 = n9078 & n9081;
  assign n9422 = ~n9082 & ~n9421;
  assign n9423 = ~n9420 & n9422;
  assign n9424 = ~n9082 & ~n9423;
  assign n9425 = n9064 & n9067;
  assign n9426 = ~n9068 & ~n9425;
  assign n9427 = ~n9424 & n9426;
  assign n9428 = ~n9068 & ~n9427;
  assign n9429 = n8971 & ~n8973;
  assign n9430 = ~n8974 & ~n9429;
  assign n9431 = ~n9428 & n9430;
  assign n9432 = ~n1637 & n7238;
  assign n9433 = n4553 & n6631;
  assign n9434 = ~n1717 & n6630;
  assign n9435 = ~n1533 & n7262;
  assign n9436 = ~n9432 & ~n9434;
  assign n9437 = ~n9435 & n9436;
  assign n9438 = ~n9433 & n9437;
  assign n9439 = ~pi14  & ~n9438;
  assign n9440 = pi14  & n9438;
  assign n9441 = ~n9439 & ~n9440;
  assign n9442 = n9428 & ~n9430;
  assign n9443 = ~n9431 & ~n9442;
  assign n9444 = ~n9441 & n9443;
  assign n9445 = ~n9431 & ~n9444;
  assign n9446 = ~n8980 & ~n8981;
  assign n9447 = ~n8991 & n9446;
  assign n9448 = n8991 & ~n9446;
  assign n9449 = ~n9447 & ~n9448;
  assign n9450 = ~n9445 & n9449;
  assign n9451 = n9445 & ~n9449;
  assign n9452 = ~n1225 & n7869;
  assign n9453 = n4135 & n7431;
  assign n9454 = ~n1345 & n7430;
  assign n9455 = ~n1104 & n7895;
  assign n9456 = ~n9452 & ~n9454;
  assign n9457 = ~n9455 & n9456;
  assign n9458 = ~n9453 & n9457;
  assign n9459 = pi11  & n9458;
  assign n9460 = ~pi11  & ~n9458;
  assign n9461 = ~n9459 & ~n9460;
  assign n9462 = ~n9451 & ~n9461;
  assign n9463 = ~n9450 & ~n9462;
  assign n9464 = n9054 & ~n9463;
  assign n9465 = ~n9054 & n9463;
  assign n9466 = ~n3855 & n9040;
  assign n9467 = n3972 & n8251;
  assign n9468 = ~n987 & n8250;
  assign n9469 = ~n3681 & n9016;
  assign n9470 = ~n9466 & ~n9468;
  assign n9471 = ~n9469 & n9470;
  assign n9472 = ~n9467 & n9471;
  assign n9473 = pi8  & n9472;
  assign n9474 = ~pi8  & ~n9472;
  assign n9475 = ~n9473 & ~n9474;
  assign n9476 = ~n9465 & ~n9475;
  assign n9477 = ~n9464 & ~n9476;
  assign n9478 = ~n9050 & ~n9477;
  assign n9479 = n9050 & ~n9477;
  assign n9480 = ~n9050 & n9477;
  assign n9481 = ~n9479 & ~n9480;
  assign n9482 = ~n9010 & ~n9012;
  assign n9483 = ~n9013 & ~n9482;
  assign n9484 = ~n9481 & n9483;
  assign n9485 = ~n9478 & ~n9484;
  assign n9486 = ~n9026 & ~n9030;
  assign n9487 = ~n9031 & ~n9486;
  assign n9488 = ~n9485 & n9487;
  assign n9489 = n9481 & ~n9483;
  assign n9490 = ~n9484 & ~n9489;
  assign n9491 = ~n70 & ~n73;
  assign n9492 = ~n3897 & n9491;
  assign n9493 = ~n75 & ~n9492;
  assign n9494 = ~n3883 & ~n9493;
  assign n9495 = pi5  & ~n9494;
  assign n9496 = ~pi5  & n9494;
  assign n9497 = ~n9495 & ~n9496;
  assign n9498 = n9424 & ~n9426;
  assign n9499 = ~n9427 & ~n9498;
  assign n9500 = ~n1717 & n7238;
  assign n9501 = n4537 & n6631;
  assign n9502 = ~n1841 & n6630;
  assign n9503 = ~n1637 & n7262;
  assign n9504 = ~n9500 & ~n9502;
  assign n9505 = ~n9503 & n9504;
  assign n9506 = ~n9501 & n9505;
  assign n9507 = pi14  & n9506;
  assign n9508 = ~pi14  & ~n9506;
  assign n9509 = ~n9507 & ~n9508;
  assign n9510 = n9499 & ~n9509;
  assign n9511 = n9420 & ~n9422;
  assign n9512 = ~n9423 & ~n9511;
  assign n9513 = ~n1841 & n7238;
  assign n9514 = n4762 & n6631;
  assign n9515 = ~n1908 & n6630;
  assign n9516 = ~n1717 & n7262;
  assign n9517 = ~n9513 & ~n9515;
  assign n9518 = ~n9516 & n9517;
  assign n9519 = ~n9514 & n9518;
  assign n9520 = pi14  & n9519;
  assign n9521 = ~pi14  & ~n9519;
  assign n9522 = ~n9520 & ~n9521;
  assign n9523 = n9512 & ~n9522;
  assign n9524 = n9098 & n9418;
  assign n9525 = ~n9419 & ~n9524;
  assign n9526 = ~n1908 & n7238;
  assign n9527 = n4779 & n6631;
  assign n9528 = ~n1998 & n6630;
  assign n9529 = ~n1841 & n7262;
  assign n9530 = ~n9526 & ~n9528;
  assign n9531 = ~n9529 & n9530;
  assign n9532 = ~n9527 & n9531;
  assign n9533 = pi14  & n9532;
  assign n9534 = ~pi14  & ~n9532;
  assign n9535 = ~n9533 & ~n9534;
  assign n9536 = n9525 & ~n9535;
  assign n9537 = n9114 & n9416;
  assign n9538 = ~n9417 & ~n9537;
  assign n9539 = ~n1998 & n7238;
  assign n9540 = n5151 & n6631;
  assign n9541 = ~n2098 & n6630;
  assign n9542 = ~n1908 & n7262;
  assign n9543 = ~n9539 & ~n9541;
  assign n9544 = ~n9542 & n9543;
  assign n9545 = ~n9540 & n9544;
  assign n9546 = pi14  & n9545;
  assign n9547 = ~pi14  & ~n9545;
  assign n9548 = ~n9546 & ~n9547;
  assign n9549 = n9538 & ~n9548;
  assign n9550 = n9412 & ~n9414;
  assign n9551 = ~n9415 & ~n9550;
  assign n9552 = ~n2098 & n7238;
  assign n9553 = n4979 & n6631;
  assign n9554 = ~n2146 & n6630;
  assign n9555 = ~n1998 & n7262;
  assign n9556 = ~n9552 & ~n9554;
  assign n9557 = ~n9555 & n9556;
  assign n9558 = ~n9553 & n9557;
  assign n9559 = pi14  & n9558;
  assign n9560 = ~pi14  & ~n9558;
  assign n9561 = ~n9559 & ~n9560;
  assign n9562 = n9551 & ~n9561;
  assign n9563 = n9408 & ~n9410;
  assign n9564 = ~n9411 & ~n9563;
  assign n9565 = ~n2098 & n7262;
  assign n9566 = n5359 & n6631;
  assign n9567 = ~n2146 & n7238;
  assign n9568 = ~n2249 & n6630;
  assign n9569 = ~n9565 & ~n9567;
  assign n9570 = ~n9568 & n9569;
  assign n9571 = ~n9566 & n9570;
  assign n9572 = pi14  & n9571;
  assign n9573 = ~pi14  & ~n9571;
  assign n9574 = ~n9572 & ~n9573;
  assign n9575 = n9564 & ~n9574;
  assign n9576 = n9158 & n9406;
  assign n9577 = ~n9407 & ~n9576;
  assign n9578 = ~n2146 & n7262;
  assign n9579 = n5343 & n6631;
  assign n9580 = ~n2347 & n6630;
  assign n9581 = ~n2249 & n7238;
  assign n9582 = ~n9578 & ~n9580;
  assign n9583 = ~n9581 & n9582;
  assign n9584 = ~n9579 & n9583;
  assign n9585 = pi14  & n9584;
  assign n9586 = ~pi14  & ~n9584;
  assign n9587 = ~n9585 & ~n9586;
  assign n9588 = n9577 & ~n9587;
  assign n9589 = ~n2412 & n6630;
  assign n9590 = n5579 & n6631;
  assign n9591 = ~n2347 & n7238;
  assign n9592 = ~n2249 & n7262;
  assign n9593 = ~n9589 & ~n9591;
  assign n9594 = ~n9592 & n9593;
  assign n9595 = ~n9590 & n9594;
  assign n9596 = ~pi14  & ~n9595;
  assign n9597 = pi14  & n9595;
  assign n9598 = ~n9596 & ~n9597;
  assign n9599 = n9402 & ~n9404;
  assign n9600 = ~n9405 & ~n9599;
  assign n9601 = ~n9598 & n9600;
  assign n9602 = ~n9598 & ~n9600;
  assign n9603 = n9598 & n9600;
  assign n9604 = ~n9602 & ~n9603;
  assign n9605 = ~n2347 & n7262;
  assign n9606 = n5596 & n6631;
  assign n9607 = ~n2496 & n6630;
  assign n9608 = ~n2412 & n7238;
  assign n9609 = ~n9605 & ~n9607;
  assign n9610 = ~n9608 & n9609;
  assign n9611 = ~n9606 & n9610;
  assign n9612 = ~pi14  & ~n9611;
  assign n9613 = pi14  & n9611;
  assign n9614 = ~n9612 & ~n9613;
  assign n9615 = n9397 & n9400;
  assign n9616 = ~n9401 & ~n9615;
  assign n9617 = ~n9614 & n9616;
  assign n9618 = ~n9614 & ~n9616;
  assign n9619 = n9614 & n9616;
  assign n9620 = ~n9618 & ~n9619;
  assign n9621 = n9200 & n9395;
  assign n9622 = ~n9396 & ~n9621;
  assign n9623 = ~n2589 & n6630;
  assign n9624 = n6016 & n6631;
  assign n9625 = ~n2496 & n7238;
  assign n9626 = ~n2412 & n7262;
  assign n9627 = ~n9623 & ~n9625;
  assign n9628 = ~n9626 & n9627;
  assign n9629 = ~n9624 & n9628;
  assign n9630 = pi14  & n9629;
  assign n9631 = ~pi14  & ~n9629;
  assign n9632 = ~n9630 & ~n9631;
  assign n9633 = n9622 & ~n9632;
  assign n9634 = n9216 & n9393;
  assign n9635 = ~n9394 & ~n9634;
  assign n9636 = ~n2496 & n7262;
  assign n9637 = n5776 & n6631;
  assign n9638 = ~n2674 & n6630;
  assign n9639 = ~n2589 & n7238;
  assign n9640 = ~n9636 & ~n9638;
  assign n9641 = ~n9639 & n9640;
  assign n9642 = ~n9637 & n9641;
  assign n9643 = pi14  & n9642;
  assign n9644 = ~pi14  & ~n9642;
  assign n9645 = ~n9643 & ~n9644;
  assign n9646 = n9635 & ~n9645;
  assign n9647 = n9389 & ~n9391;
  assign n9648 = ~n9392 & ~n9647;
  assign n9649 = ~n2674 & n7238;
  assign n9650 = n6240 & n6631;
  assign n9651 = ~n2708 & n6630;
  assign n9652 = ~n2589 & n7262;
  assign n9653 = ~n9649 & ~n9651;
  assign n9654 = ~n9652 & n9653;
  assign n9655 = ~n9650 & n9654;
  assign n9656 = pi14  & n9655;
  assign n9657 = ~pi14  & ~n9655;
  assign n9658 = ~n9656 & ~n9657;
  assign n9659 = n9648 & ~n9658;
  assign n9660 = ~n2778 & n6630;
  assign n9661 = n6393 & n6631;
  assign n9662 = ~n2708 & n7238;
  assign n9663 = ~n2674 & n7262;
  assign n9664 = ~n9660 & ~n9662;
  assign n9665 = ~n9663 & n9664;
  assign n9666 = ~n9661 & n9665;
  assign n9667 = ~pi14  & ~n9666;
  assign n9668 = pi14  & n9666;
  assign n9669 = ~n9667 & ~n9668;
  assign n9670 = n9385 & ~n9387;
  assign n9671 = ~n9388 & ~n9670;
  assign n9672 = ~n9669 & n9671;
  assign n9673 = ~n9669 & ~n9671;
  assign n9674 = n9669 & n9671;
  assign n9675 = ~n9673 & ~n9674;
  assign n9676 = ~n2708 & n7262;
  assign n9677 = n6222 & n6631;
  assign n9678 = ~n2835 & n6630;
  assign n9679 = ~n2778 & n7238;
  assign n9680 = ~n9676 & ~n9678;
  assign n9681 = ~n9679 & n9680;
  assign n9682 = ~n9677 & n9681;
  assign n9683 = ~pi14  & ~n9682;
  assign n9684 = pi14  & n9682;
  assign n9685 = ~n9683 & ~n9684;
  assign n9686 = n9380 & n9383;
  assign n9687 = ~n9384 & ~n9686;
  assign n9688 = ~n9685 & n9687;
  assign n9689 = ~n9685 & ~n9687;
  assign n9690 = n9685 & n9687;
  assign n9691 = ~n9689 & ~n9690;
  assign n9692 = ~n2919 & n6630;
  assign n9693 = n6509 & n6631;
  assign n9694 = ~n2835 & n7238;
  assign n9695 = ~n2778 & n7262;
  assign n9696 = ~n9692 & ~n9694;
  assign n9697 = ~n9695 & n9696;
  assign n9698 = ~n9693 & n9697;
  assign n9699 = ~pi14  & ~n9698;
  assign n9700 = pi14  & n9698;
  assign n9701 = ~n9699 & ~n9700;
  assign n9702 = ~n9375 & n9378;
  assign n9703 = n9375 & ~n9378;
  assign n9704 = ~n9702 & ~n9703;
  assign n9705 = ~n9701 & ~n9704;
  assign n9706 = n9285 & n9373;
  assign n9707 = ~n9374 & ~n9706;
  assign n9708 = ~n2919 & n7238;
  assign n9709 = n6631 & n6809;
  assign n9710 = ~n2951 & n6630;
  assign n9711 = ~n2835 & n7262;
  assign n9712 = ~n9708 & ~n9710;
  assign n9713 = ~n9711 & n9712;
  assign n9714 = ~n9709 & n9713;
  assign n9715 = pi14  & n9714;
  assign n9716 = ~pi14  & ~n9714;
  assign n9717 = ~n9715 & ~n9716;
  assign n9718 = n9707 & ~n9717;
  assign n9719 = n9369 & ~n9371;
  assign n9720 = ~n9372 & ~n9719;
  assign n9721 = ~n2919 & n7262;
  assign n9722 = n6631 & n6821;
  assign n9723 = ~n2951 & n7238;
  assign n9724 = ~n3031 & n6630;
  assign n9725 = ~n9721 & ~n9723;
  assign n9726 = ~n9724 & n9725;
  assign n9727 = ~n9722 & n9726;
  assign n9728 = pi14  & n9727;
  assign n9729 = ~pi14  & ~n9727;
  assign n9730 = ~n9728 & ~n9729;
  assign n9731 = n9720 & ~n9730;
  assign n9732 = n9316 & n9367;
  assign n9733 = ~n9368 & ~n9732;
  assign n9734 = ~n2951 & n7262;
  assign n9735 = n6486 & n6631;
  assign n9736 = ~n3118 & n6630;
  assign n9737 = ~n3031 & n7238;
  assign n9738 = ~n9734 & ~n9736;
  assign n9739 = ~n9737 & n9738;
  assign n9740 = ~n9735 & n9739;
  assign n9741 = pi14  & n9740;
  assign n9742 = ~pi14  & ~n9740;
  assign n9743 = ~n9741 & ~n9742;
  assign n9744 = n9733 & ~n9743;
  assign n9745 = ~n3182 & n6630;
  assign n9746 = n6631 & n6863;
  assign n9747 = ~n3118 & n7238;
  assign n9748 = ~n3031 & n7262;
  assign n9749 = ~n9745 & ~n9747;
  assign n9750 = ~n9748 & n9749;
  assign n9751 = ~n9746 & n9750;
  assign n9752 = ~pi14  & ~n9751;
  assign n9753 = pi14  & n9751;
  assign n9754 = ~n9752 & ~n9753;
  assign n9755 = n9363 & ~n9365;
  assign n9756 = ~n9366 & ~n9755;
  assign n9757 = ~n9754 & n9756;
  assign n9758 = ~n9754 & ~n9756;
  assign n9759 = n9754 & n9756;
  assign n9760 = ~n9758 & ~n9759;
  assign n9761 = ~n3118 & n7262;
  assign n9762 = n6631 & n6908;
  assign n9763 = ~n3241 & n6630;
  assign n9764 = ~n3182 & n7238;
  assign n9765 = ~n9761 & ~n9763;
  assign n9766 = ~n9764 & n9765;
  assign n9767 = ~n9762 & n9766;
  assign n9768 = pi14  & n9767;
  assign n9769 = ~pi14  & ~n9767;
  assign n9770 = ~n9768 & ~n9769;
  assign n9771 = n9351 & n9361;
  assign n9772 = ~n9362 & ~n9771;
  assign n9773 = ~n9770 & n9772;
  assign n9774 = ~n3275 & n6630;
  assign n9775 = n6631 & n6959;
  assign n9776 = ~n3241 & n7238;
  assign n9777 = ~n3182 & n7262;
  assign n9778 = ~n9774 & ~n9776;
  assign n9779 = ~n9777 & n9778;
  assign n9780 = ~n9775 & n9779;
  assign n9781 = ~pi14  & ~n9780;
  assign n9782 = pi14  & n9780;
  assign n9783 = ~n9781 & ~n9782;
  assign n9784 = pi17  & ~n9339;
  assign n9785 = n9346 & ~n9784;
  assign n9786 = ~n9346 & n9784;
  assign n9787 = ~n9785 & ~n9786;
  assign n9788 = ~n9783 & n9787;
  assign n9789 = ~n9783 & ~n9787;
  assign n9790 = n9783 & n9787;
  assign n9791 = ~n9789 & ~n9790;
  assign n9792 = ~n3241 & n7262;
  assign n9793 = n6631 & n7004;
  assign n9794 = ~n3275 & n7238;
  assign n9795 = ~n3370 & n6630;
  assign n9796 = ~n9792 & ~n9794;
  assign n9797 = ~n9795 & n9796;
  assign n9798 = ~n9793 & n9797;
  assign n9799 = pi14  & n9798;
  assign n9800 = ~pi14  & ~n9798;
  assign n9801 = ~n9799 & ~n9800;
  assign n9802 = pi17  & n9332;
  assign n9803 = ~n9337 & n9802;
  assign n9804 = n9337 & ~n9802;
  assign n9805 = ~n9803 & ~n9804;
  assign n9806 = ~n9801 & n9805;
  assign n9807 = ~n3427 & ~n6628;
  assign n9808 = ~n3427 & n7238;
  assign n9809 = ~n3485 & n7262;
  assign n9810 = n6631 & ~n7720;
  assign n9811 = ~n9808 & ~n9809;
  assign n9812 = ~n9810 & n9811;
  assign n9813 = pi14  & ~n9807;
  assign n9814 = n9812 & n9813;
  assign n9815 = ~n3427 & n6630;
  assign n9816 = n6631 & n7045;
  assign n9817 = ~n3485 & n7238;
  assign n9818 = ~n3370 & n7262;
  assign n9819 = ~n9815 & ~n9817;
  assign n9820 = ~n9818 & n9819;
  assign n9821 = ~n9816 & n9820;
  assign n9822 = n9814 & n9821;
  assign n9823 = n9332 & n9822;
  assign n9824 = ~n9332 & n9822;
  assign n9825 = n9332 & ~n9822;
  assign n9826 = ~n9824 & ~n9825;
  assign n9827 = ~n3275 & n7262;
  assign n9828 = n6631 & n7102;
  assign n9829 = ~n3485 & n6630;
  assign n9830 = ~n3370 & n7238;
  assign n9831 = ~n9827 & ~n9829;
  assign n9832 = ~n9830 & n9831;
  assign n9833 = ~n9828 & n9832;
  assign n9834 = pi14  & n9833;
  assign n9835 = ~pi14  & ~n9833;
  assign n9836 = ~n9834 & ~n9835;
  assign n9837 = ~n9826 & ~n9836;
  assign n9838 = ~n9823 & ~n9837;
  assign n9839 = n9801 & ~n9805;
  assign n9840 = ~n9806 & ~n9839;
  assign n9841 = ~n9838 & n9840;
  assign n9842 = ~n9806 & ~n9841;
  assign n9843 = ~n9791 & ~n9842;
  assign n9844 = ~n9788 & ~n9843;
  assign n9845 = n9770 & ~n9772;
  assign n9846 = ~n9773 & ~n9845;
  assign n9847 = ~n9844 & n9846;
  assign n9848 = ~n9773 & ~n9847;
  assign n9849 = ~n9760 & ~n9848;
  assign n9850 = ~n9757 & ~n9849;
  assign n9851 = n9733 & n9743;
  assign n9852 = ~n9733 & ~n9743;
  assign n9853 = ~n9851 & ~n9852;
  assign n9854 = ~n9850 & ~n9853;
  assign n9855 = ~n9744 & ~n9854;
  assign n9856 = n9720 & n9730;
  assign n9857 = ~n9720 & ~n9730;
  assign n9858 = ~n9856 & ~n9857;
  assign n9859 = ~n9855 & ~n9858;
  assign n9860 = ~n9731 & ~n9859;
  assign n9861 = ~n9707 & n9717;
  assign n9862 = ~n9718 & ~n9861;
  assign n9863 = ~n9860 & n9862;
  assign n9864 = ~n9718 & ~n9863;
  assign n9865 = n9701 & n9704;
  assign n9866 = ~n9705 & ~n9865;
  assign n9867 = ~n9864 & n9866;
  assign n9868 = ~n9705 & ~n9867;
  assign n9869 = ~n9691 & ~n9868;
  assign n9870 = ~n9688 & ~n9869;
  assign n9871 = ~n9675 & ~n9870;
  assign n9872 = ~n9672 & ~n9871;
  assign n9873 = n9648 & n9658;
  assign n9874 = ~n9648 & ~n9658;
  assign n9875 = ~n9873 & ~n9874;
  assign n9876 = ~n9872 & ~n9875;
  assign n9877 = ~n9659 & ~n9876;
  assign n9878 = n9635 & n9645;
  assign n9879 = ~n9635 & ~n9645;
  assign n9880 = ~n9878 & ~n9879;
  assign n9881 = ~n9877 & ~n9880;
  assign n9882 = ~n9646 & ~n9881;
  assign n9883 = ~n9622 & n9632;
  assign n9884 = ~n9633 & ~n9883;
  assign n9885 = ~n9882 & n9884;
  assign n9886 = ~n9633 & ~n9885;
  assign n9887 = ~n9620 & ~n9886;
  assign n9888 = ~n9617 & ~n9887;
  assign n9889 = ~n9604 & ~n9888;
  assign n9890 = ~n9601 & ~n9889;
  assign n9891 = n9577 & n9587;
  assign n9892 = ~n9577 & ~n9587;
  assign n9893 = ~n9891 & ~n9892;
  assign n9894 = ~n9890 & ~n9893;
  assign n9895 = ~n9588 & ~n9894;
  assign n9896 = n9564 & n9574;
  assign n9897 = ~n9564 & ~n9574;
  assign n9898 = ~n9896 & ~n9897;
  assign n9899 = ~n9895 & ~n9898;
  assign n9900 = ~n9575 & ~n9899;
  assign n9901 = n9551 & n9561;
  assign n9902 = ~n9551 & ~n9561;
  assign n9903 = ~n9901 & ~n9902;
  assign n9904 = ~n9900 & ~n9903;
  assign n9905 = ~n9562 & ~n9904;
  assign n9906 = n9538 & n9548;
  assign n9907 = ~n9538 & ~n9548;
  assign n9908 = ~n9906 & ~n9907;
  assign n9909 = ~n9905 & ~n9908;
  assign n9910 = ~n9549 & ~n9909;
  assign n9911 = n9525 & n9535;
  assign n9912 = ~n9525 & ~n9535;
  assign n9913 = ~n9911 & ~n9912;
  assign n9914 = ~n9910 & ~n9913;
  assign n9915 = ~n9536 & ~n9914;
  assign n9916 = n9512 & n9522;
  assign n9917 = ~n9512 & ~n9522;
  assign n9918 = ~n9916 & ~n9917;
  assign n9919 = ~n9915 & ~n9918;
  assign n9920 = ~n9523 & ~n9919;
  assign n9921 = n9499 & n9509;
  assign n9922 = ~n9499 & ~n9509;
  assign n9923 = ~n9921 & ~n9922;
  assign n9924 = ~n9920 & ~n9923;
  assign n9925 = ~n9510 & ~n9924;
  assign n9926 = n9441 & ~n9443;
  assign n9927 = ~n9444 & ~n9926;
  assign n9928 = ~n9925 & n9927;
  assign n9929 = ~n1345 & n7869;
  assign n9930 = n4152 & n7431;
  assign n9931 = ~n1448 & n7430;
  assign n9932 = ~n1225 & n7895;
  assign n9933 = ~n9929 & ~n9931;
  assign n9934 = ~n9932 & n9933;
  assign n9935 = ~n9930 & n9934;
  assign n9936 = ~pi11  & ~n9935;
  assign n9937 = pi11  & n9935;
  assign n9938 = ~n9936 & ~n9937;
  assign n9939 = n9925 & ~n9927;
  assign n9940 = ~n9928 & ~n9939;
  assign n9941 = ~n9938 & n9940;
  assign n9942 = ~n9928 & ~n9941;
  assign n9943 = ~n9450 & ~n9451;
  assign n9944 = ~n9461 & n9943;
  assign n9945 = n9461 & ~n9943;
  assign n9946 = ~n9944 & ~n9945;
  assign n9947 = ~n9942 & n9946;
  assign n9948 = n9942 & ~n9946;
  assign n9949 = ~n878 & n8250;
  assign n9950 = n3687 & n8251;
  assign n9951 = ~n987 & n9016;
  assign n9952 = ~n3681 & n9040;
  assign n9953 = ~n9949 & ~n9951;
  assign n9954 = ~n9952 & n9953;
  assign n9955 = ~n9950 & n9954;
  assign n9956 = pi8  & n9955;
  assign n9957 = ~pi8  & ~n9955;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = ~n9948 & ~n9958;
  assign n9960 = ~n9947 & ~n9959;
  assign n9961 = ~n9497 & ~n9960;
  assign n9962 = n9497 & n9960;
  assign n9963 = ~n9464 & ~n9465;
  assign n9964 = ~n9475 & n9963;
  assign n9965 = n9475 & ~n9963;
  assign n9966 = ~n9964 & ~n9965;
  assign n9967 = ~n9962 & n9966;
  assign n9968 = ~n9961 & ~n9967;
  assign n9969 = n9490 & ~n9968;
  assign n9970 = ~n1448 & n7869;
  assign n9971 = n4453 & n7431;
  assign n9972 = ~n1533 & n7430;
  assign n9973 = ~n1345 & n7895;
  assign n9974 = ~n9970 & ~n9972;
  assign n9975 = ~n9973 & n9974;
  assign n9976 = ~n9971 & n9975;
  assign n9977 = ~pi11  & ~n9976;
  assign n9978 = pi11  & n9976;
  assign n9979 = ~n9977 & ~n9978;
  assign n9980 = n9920 & n9923;
  assign n9981 = ~n9924 & ~n9980;
  assign n9982 = ~n9979 & n9981;
  assign n9983 = ~n9979 & ~n9981;
  assign n9984 = n9979 & n9981;
  assign n9985 = ~n9983 & ~n9984;
  assign n9986 = ~n1533 & n7869;
  assign n9987 = n4355 & n7431;
  assign n9988 = ~n1637 & n7430;
  assign n9989 = ~n1448 & n7895;
  assign n9990 = ~n9986 & ~n9988;
  assign n9991 = ~n9989 & n9990;
  assign n9992 = ~n9987 & n9991;
  assign n9993 = ~pi11  & ~n9992;
  assign n9994 = pi11  & n9992;
  assign n9995 = ~n9993 & ~n9994;
  assign n9996 = n9915 & n9918;
  assign n9997 = ~n9919 & ~n9996;
  assign n9998 = ~n9995 & n9997;
  assign n9999 = ~n9995 & ~n9997;
  assign n10000 = n9995 & n9997;
  assign n10001 = ~n9999 & ~n10000;
  assign n10002 = ~n1637 & n7869;
  assign n10003 = n4553 & n7431;
  assign n10004 = ~n1717 & n7430;
  assign n10005 = ~n1533 & n7895;
  assign n10006 = ~n10002 & ~n10004;
  assign n10007 = ~n10005 & n10006;
  assign n10008 = ~n10003 & n10007;
  assign n10009 = ~pi11  & ~n10008;
  assign n10010 = pi11  & n10008;
  assign n10011 = ~n10009 & ~n10010;
  assign n10012 = ~n9910 & n9913;
  assign n10013 = n9910 & ~n9913;
  assign n10014 = ~n10012 & ~n10013;
  assign n10015 = ~n10011 & ~n10014;
  assign n10016 = ~n1717 & n7869;
  assign n10017 = n4537 & n7431;
  assign n10018 = ~n1841 & n7430;
  assign n10019 = ~n1637 & n7895;
  assign n10020 = ~n10016 & ~n10018;
  assign n10021 = ~n10019 & n10020;
  assign n10022 = ~n10017 & n10021;
  assign n10023 = ~pi11  & ~n10022;
  assign n10024 = pi11  & n10022;
  assign n10025 = ~n10023 & ~n10024;
  assign n10026 = ~n9905 & n9908;
  assign n10027 = n9905 & ~n9908;
  assign n10028 = ~n10026 & ~n10027;
  assign n10029 = ~n10025 & ~n10028;
  assign n10030 = ~n1841 & n7869;
  assign n10031 = n4762 & n7431;
  assign n10032 = ~n1908 & n7430;
  assign n10033 = ~n1717 & n7895;
  assign n10034 = ~n10030 & ~n10032;
  assign n10035 = ~n10033 & n10034;
  assign n10036 = ~n10031 & n10035;
  assign n10037 = ~pi11  & ~n10036;
  assign n10038 = pi11  & n10036;
  assign n10039 = ~n10037 & ~n10038;
  assign n10040 = n9900 & n9903;
  assign n10041 = ~n9904 & ~n10040;
  assign n10042 = ~n10039 & n10041;
  assign n10043 = ~n10039 & ~n10041;
  assign n10044 = n10039 & n10041;
  assign n10045 = ~n10043 & ~n10044;
  assign n10046 = ~n1908 & n7869;
  assign n10047 = n4779 & n7431;
  assign n10048 = ~n1998 & n7430;
  assign n10049 = ~n1841 & n7895;
  assign n10050 = ~n10046 & ~n10048;
  assign n10051 = ~n10049 & n10050;
  assign n10052 = ~n10047 & n10051;
  assign n10053 = ~pi11  & ~n10052;
  assign n10054 = pi11  & n10052;
  assign n10055 = ~n10053 & ~n10054;
  assign n10056 = n9895 & n9898;
  assign n10057 = ~n9899 & ~n10056;
  assign n10058 = ~n10055 & n10057;
  assign n10059 = ~n10055 & ~n10057;
  assign n10060 = n10055 & n10057;
  assign n10061 = ~n10059 & ~n10060;
  assign n10062 = ~n1998 & n7869;
  assign n10063 = n5151 & n7431;
  assign n10064 = ~n2098 & n7430;
  assign n10065 = ~n1908 & n7895;
  assign n10066 = ~n10062 & ~n10064;
  assign n10067 = ~n10065 & n10066;
  assign n10068 = ~n10063 & n10067;
  assign n10069 = ~pi11  & ~n10068;
  assign n10070 = pi11  & n10068;
  assign n10071 = ~n10069 & ~n10070;
  assign n10072 = ~n9890 & n9893;
  assign n10073 = n9890 & ~n9893;
  assign n10074 = ~n10072 & ~n10073;
  assign n10075 = ~n10071 & ~n10074;
  assign n10076 = n9604 & n9888;
  assign n10077 = ~n9889 & ~n10076;
  assign n10078 = ~n2098 & n7869;
  assign n10079 = n4979 & n7431;
  assign n10080 = ~n2146 & n7430;
  assign n10081 = ~n1998 & n7895;
  assign n10082 = ~n10078 & ~n10080;
  assign n10083 = ~n10081 & n10082;
  assign n10084 = ~n10079 & n10083;
  assign n10085 = pi11  & n10084;
  assign n10086 = ~pi11  & ~n10084;
  assign n10087 = ~n10085 & ~n10086;
  assign n10088 = n10077 & ~n10087;
  assign n10089 = n9620 & n9886;
  assign n10090 = ~n9887 & ~n10089;
  assign n10091 = ~n2098 & n7895;
  assign n10092 = n5359 & n7431;
  assign n10093 = ~n2146 & n7869;
  assign n10094 = ~n2249 & n7430;
  assign n10095 = ~n10091 & ~n10093;
  assign n10096 = ~n10094 & n10095;
  assign n10097 = ~n10092 & n10096;
  assign n10098 = pi11  & n10097;
  assign n10099 = ~pi11  & ~n10097;
  assign n10100 = ~n10098 & ~n10099;
  assign n10101 = n10090 & ~n10100;
  assign n10102 = ~n2146 & n7895;
  assign n10103 = n5343 & n7431;
  assign n10104 = ~n2347 & n7430;
  assign n10105 = ~n2249 & n7869;
  assign n10106 = ~n10102 & ~n10104;
  assign n10107 = ~n10105 & n10106;
  assign n10108 = ~n10103 & n10107;
  assign n10109 = ~pi11  & ~n10108;
  assign n10110 = pi11  & n10108;
  assign n10111 = ~n10109 & ~n10110;
  assign n10112 = n9882 & ~n9884;
  assign n10113 = ~n9885 & ~n10112;
  assign n10114 = ~n10111 & n10113;
  assign n10115 = ~n10111 & ~n10113;
  assign n10116 = n10111 & n10113;
  assign n10117 = ~n10115 & ~n10116;
  assign n10118 = ~n2412 & n7430;
  assign n10119 = n5579 & n7431;
  assign n10120 = ~n2347 & n7869;
  assign n10121 = ~n2249 & n7895;
  assign n10122 = ~n10118 & ~n10120;
  assign n10123 = ~n10121 & n10122;
  assign n10124 = ~n10119 & n10123;
  assign n10125 = ~pi11  & ~n10124;
  assign n10126 = pi11  & n10124;
  assign n10127 = ~n10125 & ~n10126;
  assign n10128 = ~n9877 & n9880;
  assign n10129 = n9877 & ~n9880;
  assign n10130 = ~n10128 & ~n10129;
  assign n10131 = ~n10127 & ~n10130;
  assign n10132 = ~n2347 & n7895;
  assign n10133 = n5596 & n7431;
  assign n10134 = ~n2496 & n7430;
  assign n10135 = ~n2412 & n7869;
  assign n10136 = ~n10132 & ~n10134;
  assign n10137 = ~n10135 & n10136;
  assign n10138 = ~n10133 & n10137;
  assign n10139 = ~pi11  & ~n10138;
  assign n10140 = pi11  & n10138;
  assign n10141 = ~n10139 & ~n10140;
  assign n10142 = n9872 & n9875;
  assign n10143 = ~n9876 & ~n10142;
  assign n10144 = ~n10141 & n10143;
  assign n10145 = ~n10141 & ~n10143;
  assign n10146 = n10141 & n10143;
  assign n10147 = ~n10145 & ~n10146;
  assign n10148 = n9675 & n9870;
  assign n10149 = ~n9871 & ~n10148;
  assign n10150 = ~n2589 & n7430;
  assign n10151 = n6016 & n7431;
  assign n10152 = ~n2496 & n7869;
  assign n10153 = ~n2412 & n7895;
  assign n10154 = ~n10150 & ~n10152;
  assign n10155 = ~n10153 & n10154;
  assign n10156 = ~n10151 & n10155;
  assign n10157 = pi11  & n10156;
  assign n10158 = ~pi11  & ~n10156;
  assign n10159 = ~n10157 & ~n10158;
  assign n10160 = n10149 & ~n10159;
  assign n10161 = n9691 & n9868;
  assign n10162 = ~n9869 & ~n10161;
  assign n10163 = ~n2496 & n7895;
  assign n10164 = n5776 & n7431;
  assign n10165 = ~n2674 & n7430;
  assign n10166 = ~n2589 & n7869;
  assign n10167 = ~n10163 & ~n10165;
  assign n10168 = ~n10166 & n10167;
  assign n10169 = ~n10164 & n10168;
  assign n10170 = pi11  & n10169;
  assign n10171 = ~pi11  & ~n10169;
  assign n10172 = ~n10170 & ~n10171;
  assign n10173 = n10162 & ~n10172;
  assign n10174 = n9864 & ~n9866;
  assign n10175 = ~n9867 & ~n10174;
  assign n10176 = ~n2674 & n7869;
  assign n10177 = n6240 & n7431;
  assign n10178 = ~n2708 & n7430;
  assign n10179 = ~n2589 & n7895;
  assign n10180 = ~n10176 & ~n10178;
  assign n10181 = ~n10179 & n10180;
  assign n10182 = ~n10177 & n10181;
  assign n10183 = pi11  & n10182;
  assign n10184 = ~pi11  & ~n10182;
  assign n10185 = ~n10183 & ~n10184;
  assign n10186 = n10175 & ~n10185;
  assign n10187 = ~n2778 & n7430;
  assign n10188 = n6393 & n7431;
  assign n10189 = ~n2708 & n7869;
  assign n10190 = ~n2674 & n7895;
  assign n10191 = ~n10187 & ~n10189;
  assign n10192 = ~n10190 & n10191;
  assign n10193 = ~n10188 & n10192;
  assign n10194 = ~pi11  & ~n10193;
  assign n10195 = pi11  & n10193;
  assign n10196 = ~n10194 & ~n10195;
  assign n10197 = n9860 & ~n9862;
  assign n10198 = ~n9863 & ~n10197;
  assign n10199 = ~n10196 & n10198;
  assign n10200 = ~n10196 & ~n10198;
  assign n10201 = n10196 & n10198;
  assign n10202 = ~n10200 & ~n10201;
  assign n10203 = ~n2708 & n7895;
  assign n10204 = n6222 & n7431;
  assign n10205 = ~n2835 & n7430;
  assign n10206 = ~n2778 & n7869;
  assign n10207 = ~n10203 & ~n10205;
  assign n10208 = ~n10206 & n10207;
  assign n10209 = ~n10204 & n10208;
  assign n10210 = ~pi11  & ~n10209;
  assign n10211 = pi11  & n10209;
  assign n10212 = ~n10210 & ~n10211;
  assign n10213 = n9855 & n9858;
  assign n10214 = ~n9859 & ~n10213;
  assign n10215 = ~n10212 & n10214;
  assign n10216 = ~n10212 & ~n10214;
  assign n10217 = n10212 & n10214;
  assign n10218 = ~n10216 & ~n10217;
  assign n10219 = ~n2919 & n7430;
  assign n10220 = n6509 & n7431;
  assign n10221 = ~n2835 & n7869;
  assign n10222 = ~n2778 & n7895;
  assign n10223 = ~n10219 & ~n10221;
  assign n10224 = ~n10222 & n10223;
  assign n10225 = ~n10220 & n10224;
  assign n10226 = ~pi11  & ~n10225;
  assign n10227 = pi11  & n10225;
  assign n10228 = ~n10226 & ~n10227;
  assign n10229 = ~n9850 & n9853;
  assign n10230 = n9850 & ~n9853;
  assign n10231 = ~n10229 & ~n10230;
  assign n10232 = ~n10228 & ~n10231;
  assign n10233 = n9760 & n9848;
  assign n10234 = ~n9849 & ~n10233;
  assign n10235 = ~n2919 & n7869;
  assign n10236 = n6809 & n7431;
  assign n10237 = ~n2951 & n7430;
  assign n10238 = ~n2835 & n7895;
  assign n10239 = ~n10235 & ~n10237;
  assign n10240 = ~n10238 & n10239;
  assign n10241 = ~n10236 & n10240;
  assign n10242 = pi11  & n10241;
  assign n10243 = ~pi11  & ~n10241;
  assign n10244 = ~n10242 & ~n10243;
  assign n10245 = n10234 & ~n10244;
  assign n10246 = n9844 & ~n9846;
  assign n10247 = ~n9847 & ~n10246;
  assign n10248 = ~n2919 & n7895;
  assign n10249 = n6821 & n7431;
  assign n10250 = ~n2951 & n7869;
  assign n10251 = ~n3031 & n7430;
  assign n10252 = ~n10248 & ~n10250;
  assign n10253 = ~n10251 & n10252;
  assign n10254 = ~n10249 & n10253;
  assign n10255 = pi11  & n10254;
  assign n10256 = ~pi11  & ~n10254;
  assign n10257 = ~n10255 & ~n10256;
  assign n10258 = n10247 & ~n10257;
  assign n10259 = n9791 & n9842;
  assign n10260 = ~n9843 & ~n10259;
  assign n10261 = ~n2951 & n7895;
  assign n10262 = n6486 & n7431;
  assign n10263 = ~n3118 & n7430;
  assign n10264 = ~n3031 & n7869;
  assign n10265 = ~n10261 & ~n10263;
  assign n10266 = ~n10264 & n10265;
  assign n10267 = ~n10262 & n10266;
  assign n10268 = pi11  & n10267;
  assign n10269 = ~pi11  & ~n10267;
  assign n10270 = ~n10268 & ~n10269;
  assign n10271 = n10260 & ~n10270;
  assign n10272 = ~n3182 & n7430;
  assign n10273 = n6863 & n7431;
  assign n10274 = ~n3118 & n7869;
  assign n10275 = ~n3031 & n7895;
  assign n10276 = ~n10272 & ~n10274;
  assign n10277 = ~n10275 & n10276;
  assign n10278 = ~n10273 & n10277;
  assign n10279 = ~pi11  & ~n10278;
  assign n10280 = pi11  & n10278;
  assign n10281 = ~n10279 & ~n10280;
  assign n10282 = n9838 & ~n9840;
  assign n10283 = ~n9841 & ~n10282;
  assign n10284 = ~n10281 & n10283;
  assign n10285 = ~n10281 & ~n10283;
  assign n10286 = n10281 & n10283;
  assign n10287 = ~n10285 & ~n10286;
  assign n10288 = ~n3118 & n7895;
  assign n10289 = n6908 & n7431;
  assign n10290 = ~n3241 & n7430;
  assign n10291 = ~n3182 & n7869;
  assign n10292 = ~n10288 & ~n10290;
  assign n10293 = ~n10291 & n10292;
  assign n10294 = ~n10289 & n10293;
  assign n10295 = pi11  & n10294;
  assign n10296 = ~pi11  & ~n10294;
  assign n10297 = ~n10295 & ~n10296;
  assign n10298 = n9826 & n9836;
  assign n10299 = ~n9837 & ~n10298;
  assign n10300 = ~n10297 & n10299;
  assign n10301 = ~n3275 & n7430;
  assign n10302 = n6959 & n7431;
  assign n10303 = ~n3241 & n7869;
  assign n10304 = ~n3182 & n7895;
  assign n10305 = ~n10301 & ~n10303;
  assign n10306 = ~n10304 & n10305;
  assign n10307 = ~n10302 & n10306;
  assign n10308 = ~pi11  & ~n10307;
  assign n10309 = pi11  & n10307;
  assign n10310 = ~n10308 & ~n10309;
  assign n10311 = pi14  & ~n9814;
  assign n10312 = n9821 & ~n10311;
  assign n10313 = ~n9821 & n10311;
  assign n10314 = ~n10312 & ~n10313;
  assign n10315 = ~n10310 & n10314;
  assign n10316 = ~n10310 & ~n10314;
  assign n10317 = n10310 & n10314;
  assign n10318 = ~n10316 & ~n10317;
  assign n10319 = ~n3241 & n7895;
  assign n10320 = n7004 & n7431;
  assign n10321 = ~n3275 & n7869;
  assign n10322 = ~n3370 & n7430;
  assign n10323 = ~n10319 & ~n10321;
  assign n10324 = ~n10322 & n10323;
  assign n10325 = ~n10320 & n10324;
  assign n10326 = pi11  & n10325;
  assign n10327 = ~pi11  & ~n10325;
  assign n10328 = ~n10326 & ~n10327;
  assign n10329 = pi14  & n9807;
  assign n10330 = ~n9812 & n10329;
  assign n10331 = n9812 & ~n10329;
  assign n10332 = ~n10330 & ~n10331;
  assign n10333 = ~n10328 & n10332;
  assign n10334 = ~n3427 & ~n7425;
  assign n10335 = ~n3427 & n7869;
  assign n10336 = ~n3485 & n7895;
  assign n10337 = n7431 & ~n7720;
  assign n10338 = ~n10335 & ~n10336;
  assign n10339 = ~n10337 & n10338;
  assign n10340 = pi11  & ~n10334;
  assign n10341 = n10339 & n10340;
  assign n10342 = ~n3427 & n7430;
  assign n10343 = n7045 & n7431;
  assign n10344 = ~n3485 & n7869;
  assign n10345 = ~n3370 & n7895;
  assign n10346 = ~n10342 & ~n10344;
  assign n10347 = ~n10345 & n10346;
  assign n10348 = ~n10343 & n10347;
  assign n10349 = n10341 & n10348;
  assign n10350 = n9807 & n10349;
  assign n10351 = ~n9807 & n10349;
  assign n10352 = n9807 & ~n10349;
  assign n10353 = ~n10351 & ~n10352;
  assign n10354 = ~n3275 & n7895;
  assign n10355 = n7102 & n7431;
  assign n10356 = ~n3485 & n7430;
  assign n10357 = ~n3370 & n7869;
  assign n10358 = ~n10354 & ~n10356;
  assign n10359 = ~n10357 & n10358;
  assign n10360 = ~n10355 & n10359;
  assign n10361 = pi11  & n10360;
  assign n10362 = ~pi11  & ~n10360;
  assign n10363 = ~n10361 & ~n10362;
  assign n10364 = ~n10353 & ~n10363;
  assign n10365 = ~n10350 & ~n10364;
  assign n10366 = n10328 & ~n10332;
  assign n10367 = ~n10333 & ~n10366;
  assign n10368 = ~n10365 & n10367;
  assign n10369 = ~n10333 & ~n10368;
  assign n10370 = ~n10318 & ~n10369;
  assign n10371 = ~n10315 & ~n10370;
  assign n10372 = n10297 & ~n10299;
  assign n10373 = ~n10300 & ~n10372;
  assign n10374 = ~n10371 & n10373;
  assign n10375 = ~n10300 & ~n10374;
  assign n10376 = ~n10287 & ~n10375;
  assign n10377 = ~n10284 & ~n10376;
  assign n10378 = n10260 & n10270;
  assign n10379 = ~n10260 & ~n10270;
  assign n10380 = ~n10378 & ~n10379;
  assign n10381 = ~n10377 & ~n10380;
  assign n10382 = ~n10271 & ~n10381;
  assign n10383 = n10247 & n10257;
  assign n10384 = ~n10247 & ~n10257;
  assign n10385 = ~n10383 & ~n10384;
  assign n10386 = ~n10382 & ~n10385;
  assign n10387 = ~n10258 & ~n10386;
  assign n10388 = ~n10234 & n10244;
  assign n10389 = ~n10245 & ~n10388;
  assign n10390 = ~n10387 & n10389;
  assign n10391 = ~n10245 & ~n10390;
  assign n10392 = n10228 & n10231;
  assign n10393 = ~n10232 & ~n10392;
  assign n10394 = ~n10391 & n10393;
  assign n10395 = ~n10232 & ~n10394;
  assign n10396 = ~n10218 & ~n10395;
  assign n10397 = ~n10215 & ~n10396;
  assign n10398 = ~n10202 & ~n10397;
  assign n10399 = ~n10199 & ~n10398;
  assign n10400 = n10175 & n10185;
  assign n10401 = ~n10175 & ~n10185;
  assign n10402 = ~n10400 & ~n10401;
  assign n10403 = ~n10399 & ~n10402;
  assign n10404 = ~n10186 & ~n10403;
  assign n10405 = n10162 & n10172;
  assign n10406 = ~n10162 & ~n10172;
  assign n10407 = ~n10405 & ~n10406;
  assign n10408 = ~n10404 & ~n10407;
  assign n10409 = ~n10173 & ~n10408;
  assign n10410 = ~n10149 & n10159;
  assign n10411 = ~n10160 & ~n10410;
  assign n10412 = ~n10409 & n10411;
  assign n10413 = ~n10160 & ~n10412;
  assign n10414 = ~n10147 & ~n10413;
  assign n10415 = ~n10144 & ~n10414;
  assign n10416 = n10127 & n10130;
  assign n10417 = ~n10131 & ~n10416;
  assign n10418 = ~n10415 & n10417;
  assign n10419 = ~n10131 & ~n10418;
  assign n10420 = ~n10117 & ~n10419;
  assign n10421 = ~n10114 & ~n10420;
  assign n10422 = n10090 & n10100;
  assign n10423 = ~n10090 & ~n10100;
  assign n10424 = ~n10422 & ~n10423;
  assign n10425 = ~n10421 & ~n10424;
  assign n10426 = ~n10101 & ~n10425;
  assign n10427 = ~n10077 & n10087;
  assign n10428 = ~n10088 & ~n10427;
  assign n10429 = ~n10426 & n10428;
  assign n10430 = ~n10088 & ~n10429;
  assign n10431 = n10071 & n10074;
  assign n10432 = ~n10075 & ~n10431;
  assign n10433 = ~n10430 & n10432;
  assign n10434 = ~n10075 & ~n10433;
  assign n10435 = ~n10061 & ~n10434;
  assign n10436 = ~n10058 & ~n10435;
  assign n10437 = ~n10045 & ~n10436;
  assign n10438 = ~n10042 & ~n10437;
  assign n10439 = n10025 & n10028;
  assign n10440 = ~n10029 & ~n10439;
  assign n10441 = ~n10438 & n10440;
  assign n10442 = ~n10029 & ~n10441;
  assign n10443 = n10011 & n10014;
  assign n10444 = ~n10015 & ~n10443;
  assign n10445 = ~n10442 & n10444;
  assign n10446 = ~n10015 & ~n10445;
  assign n10447 = ~n10001 & ~n10446;
  assign n10448 = ~n9998 & ~n10447;
  assign n10449 = ~n9985 & ~n10448;
  assign n10450 = ~n9982 & ~n10449;
  assign n10451 = n9938 & ~n9940;
  assign n10452 = ~n9941 & ~n10451;
  assign n10453 = ~n10450 & n10452;
  assign n10454 = ~n987 & n9040;
  assign n10455 = n3791 & n8251;
  assign n10456 = ~n1104 & n8250;
  assign n10457 = ~n878 & n9016;
  assign n10458 = ~n10454 & ~n10456;
  assign n10459 = ~n10457 & n10458;
  assign n10460 = ~n10455 & n10459;
  assign n10461 = ~pi8  & ~n10460;
  assign n10462 = pi8  & n10460;
  assign n10463 = ~n10461 & ~n10462;
  assign n10464 = n10450 & ~n10452;
  assign n10465 = ~n10453 & ~n10464;
  assign n10466 = ~n10463 & n10465;
  assign n10467 = ~n10453 & ~n10466;
  assign n10468 = n75 & ~n3855;
  assign n10469 = ~n67 & n70;
  assign n10470 = ~n3883 & n10469;
  assign n10471 = ~n3900 & n9491;
  assign n10472 = ~n10468 & ~n10470;
  assign n10473 = ~n10471 & n10472;
  assign n10474 = pi5  & n10473;
  assign n10475 = ~pi5  & ~n10473;
  assign n10476 = ~n10474 & ~n10475;
  assign n10477 = ~n10467 & ~n10476;
  assign n10478 = n10467 & n10476;
  assign n10479 = ~n10477 & ~n10478;
  assign n10480 = ~n9947 & ~n9948;
  assign n10481 = ~n9958 & n10480;
  assign n10482 = n9958 & ~n10480;
  assign n10483 = ~n10481 & ~n10482;
  assign n10484 = n10479 & n10483;
  assign n10485 = ~n10477 & ~n10484;
  assign n10486 = ~n9961 & ~n9962;
  assign n10487 = n9966 & n10486;
  assign n10488 = ~n9966 & ~n10486;
  assign n10489 = ~n10487 & ~n10488;
  assign n10490 = ~n10485 & n10489;
  assign n10491 = n10485 & ~n10489;
  assign n10492 = ~n10490 & ~n10491;
  assign n10493 = n9985 & n10448;
  assign n10494 = ~n10449 & ~n10493;
  assign n10495 = ~n1104 & n9016;
  assign n10496 = n3775 & n8251;
  assign n10497 = ~n1225 & n8250;
  assign n10498 = ~n878 & n9040;
  assign n10499 = ~n10495 & ~n10497;
  assign n10500 = ~n10498 & n10499;
  assign n10501 = ~n10496 & n10500;
  assign n10502 = pi8  & n10501;
  assign n10503 = ~pi8  & ~n10501;
  assign n10504 = ~n10502 & ~n10503;
  assign n10505 = n10494 & ~n10504;
  assign n10506 = n10001 & n10446;
  assign n10507 = ~n10447 & ~n10506;
  assign n10508 = ~n1225 & n9016;
  assign n10509 = n4135 & n8251;
  assign n10510 = ~n1345 & n8250;
  assign n10511 = ~n1104 & n9040;
  assign n10512 = ~n10508 & ~n10510;
  assign n10513 = ~n10511 & n10512;
  assign n10514 = ~n10509 & n10513;
  assign n10515 = pi8  & n10514;
  assign n10516 = ~pi8  & ~n10514;
  assign n10517 = ~n10515 & ~n10516;
  assign n10518 = n10507 & ~n10517;
  assign n10519 = n10442 & ~n10444;
  assign n10520 = ~n10445 & ~n10519;
  assign n10521 = ~n1345 & n9016;
  assign n10522 = n4152 & n8251;
  assign n10523 = ~n1448 & n8250;
  assign n10524 = ~n1225 & n9040;
  assign n10525 = ~n10521 & ~n10523;
  assign n10526 = ~n10524 & n10525;
  assign n10527 = ~n10522 & n10526;
  assign n10528 = pi8  & n10527;
  assign n10529 = ~pi8  & ~n10527;
  assign n10530 = ~n10528 & ~n10529;
  assign n10531 = n10520 & ~n10530;
  assign n10532 = n10438 & ~n10440;
  assign n10533 = ~n10441 & ~n10532;
  assign n10534 = ~n1448 & n9016;
  assign n10535 = n4453 & n8251;
  assign n10536 = ~n1533 & n8250;
  assign n10537 = ~n1345 & n9040;
  assign n10538 = ~n10534 & ~n10536;
  assign n10539 = ~n10537 & n10538;
  assign n10540 = ~n10535 & n10539;
  assign n10541 = pi8  & n10540;
  assign n10542 = ~pi8  & ~n10540;
  assign n10543 = ~n10541 & ~n10542;
  assign n10544 = n10533 & ~n10543;
  assign n10545 = n10045 & n10436;
  assign n10546 = ~n10437 & ~n10545;
  assign n10547 = ~n1533 & n9016;
  assign n10548 = n4355 & n8251;
  assign n10549 = ~n1637 & n8250;
  assign n10550 = ~n1448 & n9040;
  assign n10551 = ~n10547 & ~n10549;
  assign n10552 = ~n10550 & n10551;
  assign n10553 = ~n10548 & n10552;
  assign n10554 = pi8  & n10553;
  assign n10555 = ~pi8  & ~n10553;
  assign n10556 = ~n10554 & ~n10555;
  assign n10557 = n10546 & ~n10556;
  assign n10558 = n10061 & n10434;
  assign n10559 = ~n10435 & ~n10558;
  assign n10560 = ~n1637 & n9016;
  assign n10561 = n4553 & n8251;
  assign n10562 = ~n1717 & n8250;
  assign n10563 = ~n1533 & n9040;
  assign n10564 = ~n10560 & ~n10562;
  assign n10565 = ~n10563 & n10564;
  assign n10566 = ~n10561 & n10565;
  assign n10567 = pi8  & n10566;
  assign n10568 = ~pi8  & ~n10566;
  assign n10569 = ~n10567 & ~n10568;
  assign n10570 = n10559 & ~n10569;
  assign n10571 = n10430 & ~n10432;
  assign n10572 = ~n10433 & ~n10571;
  assign n10573 = ~n1717 & n9016;
  assign n10574 = n4537 & n8251;
  assign n10575 = ~n1841 & n8250;
  assign n10576 = ~n1637 & n9040;
  assign n10577 = ~n10573 & ~n10575;
  assign n10578 = ~n10576 & n10577;
  assign n10579 = ~n10574 & n10578;
  assign n10580 = pi8  & n10579;
  assign n10581 = ~pi8  & ~n10579;
  assign n10582 = ~n10580 & ~n10581;
  assign n10583 = n10572 & ~n10582;
  assign n10584 = ~n1841 & n9016;
  assign n10585 = n4762 & n8251;
  assign n10586 = ~n1908 & n8250;
  assign n10587 = ~n1717 & n9040;
  assign n10588 = ~n10584 & ~n10586;
  assign n10589 = ~n10587 & n10588;
  assign n10590 = ~n10585 & n10589;
  assign n10591 = ~pi8  & ~n10590;
  assign n10592 = pi8  & n10590;
  assign n10593 = ~n10591 & ~n10592;
  assign n10594 = n10426 & ~n10428;
  assign n10595 = ~n10429 & ~n10594;
  assign n10596 = ~n10593 & n10595;
  assign n10597 = ~n10593 & ~n10595;
  assign n10598 = n10593 & n10595;
  assign n10599 = ~n10597 & ~n10598;
  assign n10600 = ~n1908 & n9016;
  assign n10601 = n4779 & n8251;
  assign n10602 = ~n1998 & n8250;
  assign n10603 = ~n1841 & n9040;
  assign n10604 = ~n10600 & ~n10602;
  assign n10605 = ~n10603 & n10604;
  assign n10606 = ~n10601 & n10605;
  assign n10607 = ~pi8  & ~n10606;
  assign n10608 = pi8  & n10606;
  assign n10609 = ~n10607 & ~n10608;
  assign n10610 = ~n10421 & n10424;
  assign n10611 = n10421 & ~n10424;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = ~n10609 & ~n10612;
  assign n10614 = n10117 & n10419;
  assign n10615 = ~n10420 & ~n10614;
  assign n10616 = ~n1998 & n9016;
  assign n10617 = n5151 & n8251;
  assign n10618 = ~n2098 & n8250;
  assign n10619 = ~n1908 & n9040;
  assign n10620 = ~n10616 & ~n10618;
  assign n10621 = ~n10619 & n10620;
  assign n10622 = ~n10617 & n10621;
  assign n10623 = pi8  & n10622;
  assign n10624 = ~pi8  & ~n10622;
  assign n10625 = ~n10623 & ~n10624;
  assign n10626 = n10615 & ~n10625;
  assign n10627 = n10415 & ~n10417;
  assign n10628 = ~n10418 & ~n10627;
  assign n10629 = ~n2098 & n9016;
  assign n10630 = n4979 & n8251;
  assign n10631 = ~n2146 & n8250;
  assign n10632 = ~n1998 & n9040;
  assign n10633 = ~n10629 & ~n10631;
  assign n10634 = ~n10632 & n10633;
  assign n10635 = ~n10630 & n10634;
  assign n10636 = pi8  & n10635;
  assign n10637 = ~pi8  & ~n10635;
  assign n10638 = ~n10636 & ~n10637;
  assign n10639 = n10628 & ~n10638;
  assign n10640 = n10147 & n10413;
  assign n10641 = ~n10414 & ~n10640;
  assign n10642 = ~n2098 & n9040;
  assign n10643 = n5359 & n8251;
  assign n10644 = ~n2146 & n9016;
  assign n10645 = ~n2249 & n8250;
  assign n10646 = ~n10642 & ~n10644;
  assign n10647 = ~n10645 & n10646;
  assign n10648 = ~n10643 & n10647;
  assign n10649 = pi8  & n10648;
  assign n10650 = ~pi8  & ~n10648;
  assign n10651 = ~n10649 & ~n10650;
  assign n10652 = n10641 & ~n10651;
  assign n10653 = ~n2146 & n9040;
  assign n10654 = n5343 & n8251;
  assign n10655 = ~n2347 & n8250;
  assign n10656 = ~n2249 & n9016;
  assign n10657 = ~n10653 & ~n10655;
  assign n10658 = ~n10656 & n10657;
  assign n10659 = ~n10654 & n10658;
  assign n10660 = ~pi8  & ~n10659;
  assign n10661 = pi8  & n10659;
  assign n10662 = ~n10660 & ~n10661;
  assign n10663 = n10409 & ~n10411;
  assign n10664 = ~n10412 & ~n10663;
  assign n10665 = ~n10662 & n10664;
  assign n10666 = ~n10662 & ~n10664;
  assign n10667 = n10662 & n10664;
  assign n10668 = ~n10666 & ~n10667;
  assign n10669 = ~n2412 & n8250;
  assign n10670 = n5579 & n8251;
  assign n10671 = ~n2347 & n9016;
  assign n10672 = ~n2249 & n9040;
  assign n10673 = ~n10669 & ~n10671;
  assign n10674 = ~n10672 & n10673;
  assign n10675 = ~n10670 & n10674;
  assign n10676 = ~pi8  & ~n10675;
  assign n10677 = pi8  & n10675;
  assign n10678 = ~n10676 & ~n10677;
  assign n10679 = ~n10404 & n10407;
  assign n10680 = n10404 & ~n10407;
  assign n10681 = ~n10679 & ~n10680;
  assign n10682 = ~n10678 & ~n10681;
  assign n10683 = ~n2347 & n9040;
  assign n10684 = n5596 & n8251;
  assign n10685 = ~n2496 & n8250;
  assign n10686 = ~n2412 & n9016;
  assign n10687 = ~n10683 & ~n10685;
  assign n10688 = ~n10686 & n10687;
  assign n10689 = ~n10684 & n10688;
  assign n10690 = ~pi8  & ~n10689;
  assign n10691 = pi8  & n10689;
  assign n10692 = ~n10690 & ~n10691;
  assign n10693 = n10399 & n10402;
  assign n10694 = ~n10403 & ~n10693;
  assign n10695 = ~n10692 & n10694;
  assign n10696 = ~n10692 & ~n10694;
  assign n10697 = n10692 & n10694;
  assign n10698 = ~n10696 & ~n10697;
  assign n10699 = n10202 & n10397;
  assign n10700 = ~n10398 & ~n10699;
  assign n10701 = ~n2589 & n8250;
  assign n10702 = n6016 & n8251;
  assign n10703 = ~n2496 & n9016;
  assign n10704 = ~n2412 & n9040;
  assign n10705 = ~n10701 & ~n10703;
  assign n10706 = ~n10704 & n10705;
  assign n10707 = ~n10702 & n10706;
  assign n10708 = pi8  & n10707;
  assign n10709 = ~pi8  & ~n10707;
  assign n10710 = ~n10708 & ~n10709;
  assign n10711 = n10700 & ~n10710;
  assign n10712 = n10218 & n10395;
  assign n10713 = ~n10396 & ~n10712;
  assign n10714 = ~n2496 & n9040;
  assign n10715 = n5776 & n8251;
  assign n10716 = ~n2674 & n8250;
  assign n10717 = ~n2589 & n9016;
  assign n10718 = ~n10714 & ~n10716;
  assign n10719 = ~n10717 & n10718;
  assign n10720 = ~n10715 & n10719;
  assign n10721 = pi8  & n10720;
  assign n10722 = ~pi8  & ~n10720;
  assign n10723 = ~n10721 & ~n10722;
  assign n10724 = n10713 & ~n10723;
  assign n10725 = n10391 & ~n10393;
  assign n10726 = ~n10394 & ~n10725;
  assign n10727 = ~n2674 & n9016;
  assign n10728 = n6240 & n8251;
  assign n10729 = ~n2708 & n8250;
  assign n10730 = ~n2589 & n9040;
  assign n10731 = ~n10727 & ~n10729;
  assign n10732 = ~n10730 & n10731;
  assign n10733 = ~n10728 & n10732;
  assign n10734 = pi8  & n10733;
  assign n10735 = ~pi8  & ~n10733;
  assign n10736 = ~n10734 & ~n10735;
  assign n10737 = n10726 & ~n10736;
  assign n10738 = ~n2778 & n8250;
  assign n10739 = n6393 & n8251;
  assign n10740 = ~n2708 & n9016;
  assign n10741 = ~n2674 & n9040;
  assign n10742 = ~n10738 & ~n10740;
  assign n10743 = ~n10741 & n10742;
  assign n10744 = ~n10739 & n10743;
  assign n10745 = ~pi8  & ~n10744;
  assign n10746 = pi8  & n10744;
  assign n10747 = ~n10745 & ~n10746;
  assign n10748 = n10387 & ~n10389;
  assign n10749 = ~n10390 & ~n10748;
  assign n10750 = ~n10747 & n10749;
  assign n10751 = ~n10747 & ~n10749;
  assign n10752 = n10747 & n10749;
  assign n10753 = ~n10751 & ~n10752;
  assign n10754 = ~n2708 & n9040;
  assign n10755 = n6222 & n8251;
  assign n10756 = ~n2835 & n8250;
  assign n10757 = ~n2778 & n9016;
  assign n10758 = ~n10754 & ~n10756;
  assign n10759 = ~n10757 & n10758;
  assign n10760 = ~n10755 & n10759;
  assign n10761 = ~pi8  & ~n10760;
  assign n10762 = pi8  & n10760;
  assign n10763 = ~n10761 & ~n10762;
  assign n10764 = n10382 & n10385;
  assign n10765 = ~n10386 & ~n10764;
  assign n10766 = ~n10763 & n10765;
  assign n10767 = ~n10763 & ~n10765;
  assign n10768 = n10763 & n10765;
  assign n10769 = ~n10767 & ~n10768;
  assign n10770 = ~n2919 & n8250;
  assign n10771 = n6509 & n8251;
  assign n10772 = ~n2835 & n9016;
  assign n10773 = ~n2778 & n9040;
  assign n10774 = ~n10770 & ~n10772;
  assign n10775 = ~n10773 & n10774;
  assign n10776 = ~n10771 & n10775;
  assign n10777 = ~pi8  & ~n10776;
  assign n10778 = pi8  & n10776;
  assign n10779 = ~n10777 & ~n10778;
  assign n10780 = ~n10377 & n10380;
  assign n10781 = n10377 & ~n10380;
  assign n10782 = ~n10780 & ~n10781;
  assign n10783 = ~n10779 & ~n10782;
  assign n10784 = n10287 & n10375;
  assign n10785 = ~n10376 & ~n10784;
  assign n10786 = ~n2919 & n9016;
  assign n10787 = n6809 & n8251;
  assign n10788 = ~n2951 & n8250;
  assign n10789 = ~n2835 & n9040;
  assign n10790 = ~n10786 & ~n10788;
  assign n10791 = ~n10789 & n10790;
  assign n10792 = ~n10787 & n10791;
  assign n10793 = pi8  & n10792;
  assign n10794 = ~pi8  & ~n10792;
  assign n10795 = ~n10793 & ~n10794;
  assign n10796 = n10785 & ~n10795;
  assign n10797 = n10371 & ~n10373;
  assign n10798 = ~n10374 & ~n10797;
  assign n10799 = ~n2919 & n9040;
  assign n10800 = n6821 & n8251;
  assign n10801 = ~n2951 & n9016;
  assign n10802 = ~n3031 & n8250;
  assign n10803 = ~n10799 & ~n10801;
  assign n10804 = ~n10802 & n10803;
  assign n10805 = ~n10800 & n10804;
  assign n10806 = pi8  & n10805;
  assign n10807 = ~pi8  & ~n10805;
  assign n10808 = ~n10806 & ~n10807;
  assign n10809 = n10798 & ~n10808;
  assign n10810 = n10318 & n10369;
  assign n10811 = ~n10370 & ~n10810;
  assign n10812 = ~n2951 & n9040;
  assign n10813 = n6486 & n8251;
  assign n10814 = ~n3118 & n8250;
  assign n10815 = ~n3031 & n9016;
  assign n10816 = ~n10812 & ~n10814;
  assign n10817 = ~n10815 & n10816;
  assign n10818 = ~n10813 & n10817;
  assign n10819 = pi8  & n10818;
  assign n10820 = ~pi8  & ~n10818;
  assign n10821 = ~n10819 & ~n10820;
  assign n10822 = n10811 & ~n10821;
  assign n10823 = ~n3182 & n8250;
  assign n10824 = n6863 & n8251;
  assign n10825 = ~n3118 & n9016;
  assign n10826 = ~n3031 & n9040;
  assign n10827 = ~n10823 & ~n10825;
  assign n10828 = ~n10826 & n10827;
  assign n10829 = ~n10824 & n10828;
  assign n10830 = ~pi8  & ~n10829;
  assign n10831 = pi8  & n10829;
  assign n10832 = ~n10830 & ~n10831;
  assign n10833 = n10365 & ~n10367;
  assign n10834 = ~n10368 & ~n10833;
  assign n10835 = ~n10832 & n10834;
  assign n10836 = ~n10832 & ~n10834;
  assign n10837 = n10832 & n10834;
  assign n10838 = ~n10836 & ~n10837;
  assign n10839 = ~n3118 & n9040;
  assign n10840 = n6908 & n8251;
  assign n10841 = ~n3241 & n8250;
  assign n10842 = ~n3182 & n9016;
  assign n10843 = ~n10839 & ~n10841;
  assign n10844 = ~n10842 & n10843;
  assign n10845 = ~n10840 & n10844;
  assign n10846 = pi8  & n10845;
  assign n10847 = ~pi8  & ~n10845;
  assign n10848 = ~n10846 & ~n10847;
  assign n10849 = n10353 & n10363;
  assign n10850 = ~n10364 & ~n10849;
  assign n10851 = ~n10848 & n10850;
  assign n10852 = ~n3275 & n8250;
  assign n10853 = n6959 & n8251;
  assign n10854 = ~n3241 & n9016;
  assign n10855 = ~n3182 & n9040;
  assign n10856 = ~n10852 & ~n10854;
  assign n10857 = ~n10855 & n10856;
  assign n10858 = ~n10853 & n10857;
  assign n10859 = ~pi8  & ~n10858;
  assign n10860 = pi8  & n10858;
  assign n10861 = ~n10859 & ~n10860;
  assign n10862 = pi11  & ~n10341;
  assign n10863 = n10348 & ~n10862;
  assign n10864 = ~n10348 & n10862;
  assign n10865 = ~n10863 & ~n10864;
  assign n10866 = ~n10861 & n10865;
  assign n10867 = ~n10861 & ~n10865;
  assign n10868 = n10861 & n10865;
  assign n10869 = ~n10867 & ~n10868;
  assign n10870 = ~n3241 & n9040;
  assign n10871 = n7004 & n8251;
  assign n10872 = ~n3275 & n9016;
  assign n10873 = ~n3370 & n8250;
  assign n10874 = ~n10870 & ~n10872;
  assign n10875 = ~n10873 & n10874;
  assign n10876 = ~n10871 & n10875;
  assign n10877 = pi8  & n10876;
  assign n10878 = ~pi8  & ~n10876;
  assign n10879 = ~n10877 & ~n10878;
  assign n10880 = pi11  & n10334;
  assign n10881 = ~n10339 & n10880;
  assign n10882 = n10339 & ~n10880;
  assign n10883 = ~n10881 & ~n10882;
  assign n10884 = ~n10879 & n10883;
  assign n10885 = ~n3427 & ~n8245;
  assign n10886 = ~n3427 & n9016;
  assign n10887 = ~n3485 & n9040;
  assign n10888 = ~n7720 & n8251;
  assign n10889 = ~n10886 & ~n10887;
  assign n10890 = ~n10888 & n10889;
  assign n10891 = pi8  & ~n10885;
  assign n10892 = n10890 & n10891;
  assign n10893 = ~n3427 & n8250;
  assign n10894 = n7045 & n8251;
  assign n10895 = ~n3485 & n9016;
  assign n10896 = ~n3370 & n9040;
  assign n10897 = ~n10893 & ~n10895;
  assign n10898 = ~n10896 & n10897;
  assign n10899 = ~n10894 & n10898;
  assign n10900 = n10892 & n10899;
  assign n10901 = n10334 & n10900;
  assign n10902 = ~n10334 & n10900;
  assign n10903 = n10334 & ~n10900;
  assign n10904 = ~n10902 & ~n10903;
  assign n10905 = ~n3275 & n9040;
  assign n10906 = n7102 & n8251;
  assign n10907 = ~n3485 & n8250;
  assign n10908 = ~n3370 & n9016;
  assign n10909 = ~n10905 & ~n10907;
  assign n10910 = ~n10908 & n10909;
  assign n10911 = ~n10906 & n10910;
  assign n10912 = pi8  & n10911;
  assign n10913 = ~pi8  & ~n10911;
  assign n10914 = ~n10912 & ~n10913;
  assign n10915 = ~n10904 & ~n10914;
  assign n10916 = ~n10901 & ~n10915;
  assign n10917 = n10879 & ~n10883;
  assign n10918 = ~n10884 & ~n10917;
  assign n10919 = ~n10916 & n10918;
  assign n10920 = ~n10884 & ~n10919;
  assign n10921 = ~n10869 & ~n10920;
  assign n10922 = ~n10866 & ~n10921;
  assign n10923 = n10848 & ~n10850;
  assign n10924 = ~n10851 & ~n10923;
  assign n10925 = ~n10922 & n10924;
  assign n10926 = ~n10851 & ~n10925;
  assign n10927 = ~n10838 & ~n10926;
  assign n10928 = ~n10835 & ~n10927;
  assign n10929 = n10811 & n10821;
  assign n10930 = ~n10811 & ~n10821;
  assign n10931 = ~n10929 & ~n10930;
  assign n10932 = ~n10928 & ~n10931;
  assign n10933 = ~n10822 & ~n10932;
  assign n10934 = n10798 & n10808;
  assign n10935 = ~n10798 & ~n10808;
  assign n10936 = ~n10934 & ~n10935;
  assign n10937 = ~n10933 & ~n10936;
  assign n10938 = ~n10809 & ~n10937;
  assign n10939 = ~n10785 & n10795;
  assign n10940 = ~n10796 & ~n10939;
  assign n10941 = ~n10938 & n10940;
  assign n10942 = ~n10796 & ~n10941;
  assign n10943 = n10779 & n10782;
  assign n10944 = ~n10783 & ~n10943;
  assign n10945 = ~n10942 & n10944;
  assign n10946 = ~n10783 & ~n10945;
  assign n10947 = ~n10769 & ~n10946;
  assign n10948 = ~n10766 & ~n10947;
  assign n10949 = ~n10753 & ~n10948;
  assign n10950 = ~n10750 & ~n10949;
  assign n10951 = n10726 & n10736;
  assign n10952 = ~n10726 & ~n10736;
  assign n10953 = ~n10951 & ~n10952;
  assign n10954 = ~n10950 & ~n10953;
  assign n10955 = ~n10737 & ~n10954;
  assign n10956 = n10713 & n10723;
  assign n10957 = ~n10713 & ~n10723;
  assign n10958 = ~n10956 & ~n10957;
  assign n10959 = ~n10955 & ~n10958;
  assign n10960 = ~n10724 & ~n10959;
  assign n10961 = ~n10700 & n10710;
  assign n10962 = ~n10711 & ~n10961;
  assign n10963 = ~n10960 & n10962;
  assign n10964 = ~n10711 & ~n10963;
  assign n10965 = ~n10698 & ~n10964;
  assign n10966 = ~n10695 & ~n10965;
  assign n10967 = n10678 & n10681;
  assign n10968 = ~n10682 & ~n10967;
  assign n10969 = ~n10966 & n10968;
  assign n10970 = ~n10682 & ~n10969;
  assign n10971 = ~n10668 & ~n10970;
  assign n10972 = ~n10665 & ~n10971;
  assign n10973 = n10641 & n10651;
  assign n10974 = ~n10641 & ~n10651;
  assign n10975 = ~n10973 & ~n10974;
  assign n10976 = ~n10972 & ~n10975;
  assign n10977 = ~n10652 & ~n10976;
  assign n10978 = n10628 & n10638;
  assign n10979 = ~n10628 & ~n10638;
  assign n10980 = ~n10978 & ~n10979;
  assign n10981 = ~n10977 & ~n10980;
  assign n10982 = ~n10639 & ~n10981;
  assign n10983 = ~n10615 & n10625;
  assign n10984 = ~n10626 & ~n10983;
  assign n10985 = ~n10982 & n10984;
  assign n10986 = ~n10626 & ~n10985;
  assign n10987 = n10609 & n10612;
  assign n10988 = ~n10613 & ~n10987;
  assign n10989 = ~n10986 & n10988;
  assign n10990 = ~n10613 & ~n10989;
  assign n10991 = ~n10599 & ~n10990;
  assign n10992 = ~n10596 & ~n10991;
  assign n10993 = n10572 & n10582;
  assign n10994 = ~n10572 & ~n10582;
  assign n10995 = ~n10993 & ~n10994;
  assign n10996 = ~n10992 & ~n10995;
  assign n10997 = ~n10583 & ~n10996;
  assign n10998 = n10559 & n10569;
  assign n10999 = ~n10559 & ~n10569;
  assign n11000 = ~n10998 & ~n10999;
  assign n11001 = ~n10997 & ~n11000;
  assign n11002 = ~n10570 & ~n11001;
  assign n11003 = n10546 & n10556;
  assign n11004 = ~n10546 & ~n10556;
  assign n11005 = ~n11003 & ~n11004;
  assign n11006 = ~n11002 & ~n11005;
  assign n11007 = ~n10557 & ~n11006;
  assign n11008 = n10533 & n10543;
  assign n11009 = ~n10533 & ~n10543;
  assign n11010 = ~n11008 & ~n11009;
  assign n11011 = ~n11007 & ~n11010;
  assign n11012 = ~n10544 & ~n11011;
  assign n11013 = n10520 & n10530;
  assign n11014 = ~n10520 & ~n10530;
  assign n11015 = ~n11013 & ~n11014;
  assign n11016 = ~n11012 & ~n11015;
  assign n11017 = ~n10531 & ~n11016;
  assign n11018 = n10507 & n10517;
  assign n11019 = ~n10507 & ~n10517;
  assign n11020 = ~n11018 & ~n11019;
  assign n11021 = ~n11017 & ~n11020;
  assign n11022 = ~n10518 & ~n11021;
  assign n11023 = n10494 & n10504;
  assign n11024 = ~n10494 & ~n10504;
  assign n11025 = ~n11023 & ~n11024;
  assign n11026 = ~n11022 & ~n11025;
  assign n11027 = ~n10505 & ~n11026;
  assign n11028 = n10463 & ~n10465;
  assign n11029 = ~n10466 & ~n11028;
  assign n11030 = ~n11027 & n11029;
  assign n11031 = ~n70 & n73;
  assign n11032 = ~n3883 & n11031;
  assign n11033 = n4399 & n9491;
  assign n11034 = ~n3855 & n10469;
  assign n11035 = n75 & ~n3681;
  assign n11036 = ~n11032 & ~n11034;
  assign n11037 = ~n11035 & n11036;
  assign n11038 = ~n11033 & n11037;
  assign n11039 = ~pi5  & ~n11038;
  assign n11040 = pi5  & n11038;
  assign n11041 = ~n11039 & ~n11040;
  assign n11042 = n11027 & ~n11029;
  assign n11043 = ~n11030 & ~n11042;
  assign n11044 = ~n11041 & n11043;
  assign n11045 = ~n11030 & ~n11044;
  assign n11046 = ~n10479 & ~n10483;
  assign n11047 = ~n10484 & ~n11046;
  assign n11048 = ~n11045 & n11047;
  assign n11049 = n11041 & ~n11043;
  assign n11050 = ~n11044 & ~n11049;
  assign n11051 = pi1  & ~pi2 ;
  assign n11052 = ~pi1  & pi2 ;
  assign n11053 = ~n11051 & ~n11052;
  assign n11054 = ~pi0  & ~pi1 ;
  assign n11055 = ~n11053 & n11054;
  assign n11056 = pi0  & ~n11053;
  assign n11057 = ~n3897 & n11056;
  assign n11058 = ~n11055 & ~n11057;
  assign n11059 = ~n3883 & ~n11058;
  assign n11060 = ~pi2  & n11059;
  assign n11061 = pi2  & ~n11059;
  assign n11062 = ~n11060 & ~n11061;
  assign n11063 = ~n3855 & n11031;
  assign n11064 = n3972 & n9491;
  assign n11065 = n75 & ~n987;
  assign n11066 = ~n3681 & n10469;
  assign n11067 = ~n11063 & ~n11065;
  assign n11068 = ~n11066 & n11067;
  assign n11069 = ~n11064 & n11068;
  assign n11070 = pi5  & n11069;
  assign n11071 = ~pi5  & ~n11069;
  assign n11072 = ~n11070 & ~n11071;
  assign n11073 = ~n11062 & ~n11072;
  assign n11074 = ~n11022 & n11025;
  assign n11075 = n11022 & ~n11025;
  assign n11076 = ~n11074 & ~n11075;
  assign n11077 = n11062 & n11072;
  assign n11078 = ~n11076 & ~n11077;
  assign n11079 = ~n11073 & ~n11078;
  assign n11080 = n11050 & ~n11079;
  assign n11081 = n75 & ~n878;
  assign n11082 = n3687 & n9491;
  assign n11083 = ~n987 & n10469;
  assign n11084 = ~n3681 & n11031;
  assign n11085 = ~n11081 & ~n11083;
  assign n11086 = ~n11084 & n11085;
  assign n11087 = ~n11082 & n11086;
  assign n11088 = ~pi5  & ~n11087;
  assign n11089 = pi5  & n11087;
  assign n11090 = ~n11088 & ~n11089;
  assign n11091 = ~n11017 & n11020;
  assign n11092 = n11017 & ~n11020;
  assign n11093 = ~n11091 & ~n11092;
  assign n11094 = ~n11090 & ~n11093;
  assign n11095 = ~n987 & n11031;
  assign n11096 = n3791 & n9491;
  assign n11097 = n75 & ~n1104;
  assign n11098 = ~n878 & n10469;
  assign n11099 = ~n11095 & ~n11097;
  assign n11100 = ~n11098 & n11099;
  assign n11101 = ~n11096 & n11100;
  assign n11102 = ~pi5  & ~n11101;
  assign n11103 = pi5  & n11101;
  assign n11104 = ~n11102 & ~n11103;
  assign n11105 = n11012 & n11015;
  assign n11106 = ~n11016 & ~n11105;
  assign n11107 = ~n11104 & n11106;
  assign n11108 = ~n11104 & ~n11106;
  assign n11109 = n11104 & n11106;
  assign n11110 = ~n11108 & ~n11109;
  assign n11111 = ~n1104 & n10469;
  assign n11112 = n3775 & n9491;
  assign n11113 = n75 & ~n1225;
  assign n11114 = ~n878 & n11031;
  assign n11115 = ~n11111 & ~n11113;
  assign n11116 = ~n11114 & n11115;
  assign n11117 = ~n11112 & n11116;
  assign n11118 = ~pi5  & ~n11117;
  assign n11119 = pi5  & n11117;
  assign n11120 = ~n11118 & ~n11119;
  assign n11121 = n11007 & n11010;
  assign n11122 = ~n11011 & ~n11121;
  assign n11123 = ~n11120 & n11122;
  assign n11124 = ~n11120 & ~n11122;
  assign n11125 = n11120 & n11122;
  assign n11126 = ~n11124 & ~n11125;
  assign n11127 = ~n1225 & n10469;
  assign n11128 = n4135 & n9491;
  assign n11129 = n75 & ~n1345;
  assign n11130 = ~n1104 & n11031;
  assign n11131 = ~n11127 & ~n11129;
  assign n11132 = ~n11130 & n11131;
  assign n11133 = ~n11128 & n11132;
  assign n11134 = ~pi5  & ~n11133;
  assign n11135 = pi5  & n11133;
  assign n11136 = ~n11134 & ~n11135;
  assign n11137 = ~n11002 & n11005;
  assign n11138 = n11002 & ~n11005;
  assign n11139 = ~n11137 & ~n11138;
  assign n11140 = ~n11136 & ~n11139;
  assign n11141 = ~n1345 & n10469;
  assign n11142 = n4152 & n9491;
  assign n11143 = n75 & ~n1448;
  assign n11144 = ~n1225 & n11031;
  assign n11145 = ~n11141 & ~n11143;
  assign n11146 = ~n11144 & n11145;
  assign n11147 = ~n11142 & n11146;
  assign n11148 = ~pi5  & ~n11147;
  assign n11149 = pi5  & n11147;
  assign n11150 = ~n11148 & ~n11149;
  assign n11151 = ~n10997 & n11000;
  assign n11152 = n10997 & ~n11000;
  assign n11153 = ~n11151 & ~n11152;
  assign n11154 = ~n11150 & ~n11153;
  assign n11155 = ~n1448 & n10469;
  assign n11156 = n4453 & n9491;
  assign n11157 = n75 & ~n1533;
  assign n11158 = ~n1345 & n11031;
  assign n11159 = ~n11155 & ~n11157;
  assign n11160 = ~n11158 & n11159;
  assign n11161 = ~n11156 & n11160;
  assign n11162 = ~pi5  & ~n11161;
  assign n11163 = pi5  & n11161;
  assign n11164 = ~n11162 & ~n11163;
  assign n11165 = n10992 & n10995;
  assign n11166 = ~n10996 & ~n11165;
  assign n11167 = ~n11164 & n11166;
  assign n11168 = ~n11164 & ~n11166;
  assign n11169 = n11164 & n11166;
  assign n11170 = ~n11168 & ~n11169;
  assign n11171 = n10599 & n10990;
  assign n11172 = ~n10991 & ~n11171;
  assign n11173 = ~n1533 & n10469;
  assign n11174 = n4355 & n9491;
  assign n11175 = n75 & ~n1637;
  assign n11176 = ~n1448 & n11031;
  assign n11177 = ~n11173 & ~n11175;
  assign n11178 = ~n11176 & n11177;
  assign n11179 = ~n11174 & n11178;
  assign n11180 = pi5  & n11179;
  assign n11181 = ~pi5  & ~n11179;
  assign n11182 = ~n11180 & ~n11181;
  assign n11183 = n11172 & ~n11182;
  assign n11184 = n10986 & ~n10988;
  assign n11185 = ~n10989 & ~n11184;
  assign n11186 = ~n1637 & n10469;
  assign n11187 = n4553 & n9491;
  assign n11188 = n75 & ~n1717;
  assign n11189 = ~n1533 & n11031;
  assign n11190 = ~n11186 & ~n11188;
  assign n11191 = ~n11189 & n11190;
  assign n11192 = ~n11187 & n11191;
  assign n11193 = pi5  & n11192;
  assign n11194 = ~pi5  & ~n11192;
  assign n11195 = ~n11193 & ~n11194;
  assign n11196 = n11185 & ~n11195;
  assign n11197 = ~n1717 & n10469;
  assign n11198 = n4537 & n9491;
  assign n11199 = n75 & ~n1841;
  assign n11200 = ~n1637 & n11031;
  assign n11201 = ~n11197 & ~n11199;
  assign n11202 = ~n11200 & n11201;
  assign n11203 = ~n11198 & n11202;
  assign n11204 = ~pi5  & ~n11203;
  assign n11205 = pi5  & n11203;
  assign n11206 = ~n11204 & ~n11205;
  assign n11207 = n10982 & ~n10984;
  assign n11208 = ~n10985 & ~n11207;
  assign n11209 = ~n11206 & n11208;
  assign n11210 = ~n11206 & ~n11208;
  assign n11211 = n11206 & n11208;
  assign n11212 = ~n11210 & ~n11211;
  assign n11213 = ~n1841 & n10469;
  assign n11214 = n4762 & n9491;
  assign n11215 = n75 & ~n1908;
  assign n11216 = ~n1717 & n11031;
  assign n11217 = ~n11213 & ~n11215;
  assign n11218 = ~n11216 & n11217;
  assign n11219 = ~n11214 & n11218;
  assign n11220 = ~pi5  & ~n11219;
  assign n11221 = pi5  & n11219;
  assign n11222 = ~n11220 & ~n11221;
  assign n11223 = n10977 & n10980;
  assign n11224 = ~n10981 & ~n11223;
  assign n11225 = ~n11222 & n11224;
  assign n11226 = ~n11222 & ~n11224;
  assign n11227 = n11222 & n11224;
  assign n11228 = ~n11226 & ~n11227;
  assign n11229 = ~n1908 & n10469;
  assign n11230 = n4779 & n9491;
  assign n11231 = n75 & ~n1998;
  assign n11232 = ~n1841 & n11031;
  assign n11233 = ~n11229 & ~n11231;
  assign n11234 = ~n11232 & n11233;
  assign n11235 = ~n11230 & n11234;
  assign n11236 = ~pi5  & ~n11235;
  assign n11237 = pi5  & n11235;
  assign n11238 = ~n11236 & ~n11237;
  assign n11239 = ~n10972 & n10975;
  assign n11240 = n10972 & ~n10975;
  assign n11241 = ~n11239 & ~n11240;
  assign n11242 = ~n11238 & ~n11241;
  assign n11243 = n10668 & n10970;
  assign n11244 = ~n10971 & ~n11243;
  assign n11245 = ~n1998 & n10469;
  assign n11246 = n5151 & n9491;
  assign n11247 = n75 & ~n2098;
  assign n11248 = ~n1908 & n11031;
  assign n11249 = ~n11245 & ~n11247;
  assign n11250 = ~n11248 & n11249;
  assign n11251 = ~n11246 & n11250;
  assign n11252 = pi5  & n11251;
  assign n11253 = ~pi5  & ~n11251;
  assign n11254 = ~n11252 & ~n11253;
  assign n11255 = n11244 & ~n11254;
  assign n11256 = n10966 & ~n10968;
  assign n11257 = ~n10969 & ~n11256;
  assign n11258 = ~n2098 & n10469;
  assign n11259 = n4979 & n9491;
  assign n11260 = n75 & ~n2146;
  assign n11261 = ~n1998 & n11031;
  assign n11262 = ~n11258 & ~n11260;
  assign n11263 = ~n11261 & n11262;
  assign n11264 = ~n11259 & n11263;
  assign n11265 = pi5  & n11264;
  assign n11266 = ~pi5  & ~n11264;
  assign n11267 = ~n11265 & ~n11266;
  assign n11268 = n11257 & ~n11267;
  assign n11269 = n10698 & n10964;
  assign n11270 = ~n10965 & ~n11269;
  assign n11271 = ~n2098 & n11031;
  assign n11272 = n5359 & n9491;
  assign n11273 = ~n2146 & n10469;
  assign n11274 = n75 & ~n2249;
  assign n11275 = ~n11271 & ~n11273;
  assign n11276 = ~n11274 & n11275;
  assign n11277 = ~n11272 & n11276;
  assign n11278 = pi5  & n11277;
  assign n11279 = ~pi5  & ~n11277;
  assign n11280 = ~n11278 & ~n11279;
  assign n11281 = n11270 & ~n11280;
  assign n11282 = ~n2146 & n11031;
  assign n11283 = n5343 & n9491;
  assign n11284 = n75 & ~n2347;
  assign n11285 = ~n2249 & n10469;
  assign n11286 = ~n11282 & ~n11284;
  assign n11287 = ~n11285 & n11286;
  assign n11288 = ~n11283 & n11287;
  assign n11289 = ~pi5  & ~n11288;
  assign n11290 = pi5  & n11288;
  assign n11291 = ~n11289 & ~n11290;
  assign n11292 = n10960 & ~n10962;
  assign n11293 = ~n10963 & ~n11292;
  assign n11294 = ~n11291 & n11293;
  assign n11295 = ~n11291 & ~n11293;
  assign n11296 = n11291 & n11293;
  assign n11297 = ~n11295 & ~n11296;
  assign n11298 = n75 & ~n2412;
  assign n11299 = n5579 & n9491;
  assign n11300 = ~n2347 & n10469;
  assign n11301 = ~n2249 & n11031;
  assign n11302 = ~n11298 & ~n11300;
  assign n11303 = ~n11301 & n11302;
  assign n11304 = ~n11299 & n11303;
  assign n11305 = ~pi5  & ~n11304;
  assign n11306 = pi5  & n11304;
  assign n11307 = ~n11305 & ~n11306;
  assign n11308 = ~n10955 & n10958;
  assign n11309 = n10955 & ~n10958;
  assign n11310 = ~n11308 & ~n11309;
  assign n11311 = ~n11307 & ~n11310;
  assign n11312 = ~n2347 & n11031;
  assign n11313 = n5596 & n9491;
  assign n11314 = n75 & ~n2496;
  assign n11315 = ~n2412 & n10469;
  assign n11316 = ~n11312 & ~n11314;
  assign n11317 = ~n11315 & n11316;
  assign n11318 = ~n11313 & n11317;
  assign n11319 = ~pi5  & ~n11318;
  assign n11320 = pi5  & n11318;
  assign n11321 = ~n11319 & ~n11320;
  assign n11322 = n10950 & n10953;
  assign n11323 = ~n10954 & ~n11322;
  assign n11324 = ~n11321 & n11323;
  assign n11325 = ~n11321 & ~n11323;
  assign n11326 = n11321 & n11323;
  assign n11327 = ~n11325 & ~n11326;
  assign n11328 = n10753 & n10948;
  assign n11329 = ~n10949 & ~n11328;
  assign n11330 = n75 & ~n2589;
  assign n11331 = n6016 & n9491;
  assign n11332 = ~n2496 & n10469;
  assign n11333 = ~n2412 & n11031;
  assign n11334 = ~n11330 & ~n11332;
  assign n11335 = ~n11333 & n11334;
  assign n11336 = ~n11331 & n11335;
  assign n11337 = pi5  & n11336;
  assign n11338 = ~pi5  & ~n11336;
  assign n11339 = ~n11337 & ~n11338;
  assign n11340 = n11329 & ~n11339;
  assign n11341 = n10769 & n10946;
  assign n11342 = ~n10947 & ~n11341;
  assign n11343 = ~n2496 & n11031;
  assign n11344 = n5776 & n9491;
  assign n11345 = n75 & ~n2674;
  assign n11346 = ~n2589 & n10469;
  assign n11347 = ~n11343 & ~n11345;
  assign n11348 = ~n11346 & n11347;
  assign n11349 = ~n11344 & n11348;
  assign n11350 = pi5  & n11349;
  assign n11351 = ~pi5  & ~n11349;
  assign n11352 = ~n11350 & ~n11351;
  assign n11353 = n11342 & ~n11352;
  assign n11354 = n10942 & ~n10944;
  assign n11355 = ~n10945 & ~n11354;
  assign n11356 = ~n2674 & n10469;
  assign n11357 = n6240 & n9491;
  assign n11358 = n75 & ~n2708;
  assign n11359 = ~n2589 & n11031;
  assign n11360 = ~n11356 & ~n11358;
  assign n11361 = ~n11359 & n11360;
  assign n11362 = ~n11357 & n11361;
  assign n11363 = pi5  & n11362;
  assign n11364 = ~pi5  & ~n11362;
  assign n11365 = ~n11363 & ~n11364;
  assign n11366 = n11355 & ~n11365;
  assign n11367 = n75 & ~n2778;
  assign n11368 = n6393 & n9491;
  assign n11369 = ~n2708 & n10469;
  assign n11370 = ~n2674 & n11031;
  assign n11371 = ~n11367 & ~n11369;
  assign n11372 = ~n11370 & n11371;
  assign n11373 = ~n11368 & n11372;
  assign n11374 = ~pi5  & ~n11373;
  assign n11375 = pi5  & n11373;
  assign n11376 = ~n11374 & ~n11375;
  assign n11377 = n10938 & ~n10940;
  assign n11378 = ~n10941 & ~n11377;
  assign n11379 = ~n11376 & n11378;
  assign n11380 = ~n11376 & ~n11378;
  assign n11381 = n11376 & n11378;
  assign n11382 = ~n11380 & ~n11381;
  assign n11383 = ~n2708 & n11031;
  assign n11384 = n6222 & n9491;
  assign n11385 = n75 & ~n2835;
  assign n11386 = ~n2778 & n10469;
  assign n11387 = ~n11383 & ~n11385;
  assign n11388 = ~n11386 & n11387;
  assign n11389 = ~n11384 & n11388;
  assign n11390 = ~pi5  & ~n11389;
  assign n11391 = pi5  & n11389;
  assign n11392 = ~n11390 & ~n11391;
  assign n11393 = n10933 & n10936;
  assign n11394 = ~n10937 & ~n11393;
  assign n11395 = ~n11392 & n11394;
  assign n11396 = ~n11392 & ~n11394;
  assign n11397 = n11392 & n11394;
  assign n11398 = ~n11396 & ~n11397;
  assign n11399 = n75 & ~n2919;
  assign n11400 = n6509 & n9491;
  assign n11401 = ~n2835 & n10469;
  assign n11402 = ~n2778 & n11031;
  assign n11403 = ~n11399 & ~n11401;
  assign n11404 = ~n11402 & n11403;
  assign n11405 = ~n11400 & n11404;
  assign n11406 = ~pi5  & ~n11405;
  assign n11407 = pi5  & n11405;
  assign n11408 = ~n11406 & ~n11407;
  assign n11409 = ~n10928 & n10931;
  assign n11410 = n10928 & ~n10931;
  assign n11411 = ~n11409 & ~n11410;
  assign n11412 = ~n11408 & ~n11411;
  assign n11413 = n10838 & n10926;
  assign n11414 = ~n10927 & ~n11413;
  assign n11415 = ~n2919 & n10469;
  assign n11416 = n6809 & n9491;
  assign n11417 = n75 & ~n2951;
  assign n11418 = ~n2835 & n11031;
  assign n11419 = ~n11415 & ~n11417;
  assign n11420 = ~n11418 & n11419;
  assign n11421 = ~n11416 & n11420;
  assign n11422 = pi5  & n11421;
  assign n11423 = ~pi5  & ~n11421;
  assign n11424 = ~n11422 & ~n11423;
  assign n11425 = n11414 & ~n11424;
  assign n11426 = n10922 & ~n10924;
  assign n11427 = ~n10925 & ~n11426;
  assign n11428 = ~n2919 & n11031;
  assign n11429 = n6821 & n9491;
  assign n11430 = ~n2951 & n10469;
  assign n11431 = n75 & ~n3031;
  assign n11432 = ~n11428 & ~n11430;
  assign n11433 = ~n11431 & n11432;
  assign n11434 = ~n11429 & n11433;
  assign n11435 = pi5  & n11434;
  assign n11436 = ~pi5  & ~n11434;
  assign n11437 = ~n11435 & ~n11436;
  assign n11438 = n11427 & ~n11437;
  assign n11439 = n10869 & n10920;
  assign n11440 = ~n10921 & ~n11439;
  assign n11441 = ~n2951 & n11031;
  assign n11442 = n6486 & n9491;
  assign n11443 = n75 & ~n3118;
  assign n11444 = ~n3031 & n10469;
  assign n11445 = ~n11441 & ~n11443;
  assign n11446 = ~n11444 & n11445;
  assign n11447 = ~n11442 & n11446;
  assign n11448 = pi5  & n11447;
  assign n11449 = ~pi5  & ~n11447;
  assign n11450 = ~n11448 & ~n11449;
  assign n11451 = n11440 & ~n11450;
  assign n11452 = n75 & ~n3182;
  assign n11453 = n6863 & n9491;
  assign n11454 = ~n3118 & n10469;
  assign n11455 = ~n3031 & n11031;
  assign n11456 = ~n11452 & ~n11454;
  assign n11457 = ~n11455 & n11456;
  assign n11458 = ~n11453 & n11457;
  assign n11459 = ~pi5  & ~n11458;
  assign n11460 = pi5  & n11458;
  assign n11461 = ~n11459 & ~n11460;
  assign n11462 = n10916 & ~n10918;
  assign n11463 = ~n10919 & ~n11462;
  assign n11464 = ~n11461 & n11463;
  assign n11465 = ~n11461 & ~n11463;
  assign n11466 = n11461 & n11463;
  assign n11467 = ~n11465 & ~n11466;
  assign n11468 = ~n3118 & n11031;
  assign n11469 = n6908 & n9491;
  assign n11470 = n75 & ~n3241;
  assign n11471 = ~n3182 & n10469;
  assign n11472 = ~n11468 & ~n11470;
  assign n11473 = ~n11471 & n11472;
  assign n11474 = ~n11469 & n11473;
  assign n11475 = pi5  & n11474;
  assign n11476 = ~pi5  & ~n11474;
  assign n11477 = ~n11475 & ~n11476;
  assign n11478 = n10904 & n10914;
  assign n11479 = ~n10915 & ~n11478;
  assign n11480 = ~n11477 & n11479;
  assign n11481 = n75 & ~n3275;
  assign n11482 = n6959 & n9491;
  assign n11483 = ~n3241 & n10469;
  assign n11484 = ~n3182 & n11031;
  assign n11485 = ~n11481 & ~n11483;
  assign n11486 = ~n11484 & n11485;
  assign n11487 = ~n11482 & n11486;
  assign n11488 = ~pi5  & ~n11487;
  assign n11489 = pi5  & n11487;
  assign n11490 = ~n11488 & ~n11489;
  assign n11491 = pi8  & ~n10892;
  assign n11492 = n10899 & ~n11491;
  assign n11493 = ~n10899 & n11491;
  assign n11494 = ~n11492 & ~n11493;
  assign n11495 = ~n11490 & n11494;
  assign n11496 = ~n11490 & ~n11494;
  assign n11497 = n11490 & n11494;
  assign n11498 = ~n11496 & ~n11497;
  assign n11499 = ~n3241 & n11031;
  assign n11500 = n7004 & n9491;
  assign n11501 = ~n3275 & n10469;
  assign n11502 = n75 & ~n3370;
  assign n11503 = ~n11499 & ~n11501;
  assign n11504 = ~n11502 & n11503;
  assign n11505 = ~n11500 & n11504;
  assign n11506 = pi5  & n11505;
  assign n11507 = ~pi5  & ~n11505;
  assign n11508 = ~n11506 & ~n11507;
  assign n11509 = pi8  & n10885;
  assign n11510 = ~n10890 & n11509;
  assign n11511 = n10890 & ~n11509;
  assign n11512 = ~n11510 & ~n11511;
  assign n11513 = ~n11508 & n11512;
  assign n11514 = ~n70 & ~n3427;
  assign n11515 = ~n3427 & n10469;
  assign n11516 = ~n3485 & n11031;
  assign n11517 = ~n7720 & n9491;
  assign n11518 = ~n11515 & ~n11516;
  assign n11519 = ~n11517 & n11518;
  assign n11520 = pi5  & ~n11514;
  assign n11521 = n11519 & n11520;
  assign n11522 = n75 & ~n3427;
  assign n11523 = n7045 & n9491;
  assign n11524 = ~n3485 & n10469;
  assign n11525 = ~n3370 & n11031;
  assign n11526 = ~n11522 & ~n11524;
  assign n11527 = ~n11525 & n11526;
  assign n11528 = ~n11523 & n11527;
  assign n11529 = n11521 & n11528;
  assign n11530 = n10885 & n11529;
  assign n11531 = ~n10885 & n11529;
  assign n11532 = n10885 & ~n11529;
  assign n11533 = ~n11531 & ~n11532;
  assign n11534 = ~n3275 & n11031;
  assign n11535 = n7102 & n9491;
  assign n11536 = n75 & ~n3485;
  assign n11537 = ~n3370 & n10469;
  assign n11538 = ~n11534 & ~n11536;
  assign n11539 = ~n11537 & n11538;
  assign n11540 = ~n11535 & n11539;
  assign n11541 = pi5  & n11540;
  assign n11542 = ~pi5  & ~n11540;
  assign n11543 = ~n11541 & ~n11542;
  assign n11544 = ~n11533 & ~n11543;
  assign n11545 = ~n11530 & ~n11544;
  assign n11546 = n11508 & ~n11512;
  assign n11547 = ~n11513 & ~n11546;
  assign n11548 = ~n11545 & n11547;
  assign n11549 = ~n11513 & ~n11548;
  assign n11550 = ~n11498 & ~n11549;
  assign n11551 = ~n11495 & ~n11550;
  assign n11552 = n11477 & ~n11479;
  assign n11553 = ~n11480 & ~n11552;
  assign n11554 = ~n11551 & n11553;
  assign n11555 = ~n11480 & ~n11554;
  assign n11556 = ~n11467 & ~n11555;
  assign n11557 = ~n11464 & ~n11556;
  assign n11558 = n11440 & n11450;
  assign n11559 = ~n11440 & ~n11450;
  assign n11560 = ~n11558 & ~n11559;
  assign n11561 = ~n11557 & ~n11560;
  assign n11562 = ~n11451 & ~n11561;
  assign n11563 = n11427 & n11437;
  assign n11564 = ~n11427 & ~n11437;
  assign n11565 = ~n11563 & ~n11564;
  assign n11566 = ~n11562 & ~n11565;
  assign n11567 = ~n11438 & ~n11566;
  assign n11568 = ~n11414 & n11424;
  assign n11569 = ~n11425 & ~n11568;
  assign n11570 = ~n11567 & n11569;
  assign n11571 = ~n11425 & ~n11570;
  assign n11572 = n11408 & n11411;
  assign n11573 = ~n11412 & ~n11572;
  assign n11574 = ~n11571 & n11573;
  assign n11575 = ~n11412 & ~n11574;
  assign n11576 = ~n11398 & ~n11575;
  assign n11577 = ~n11395 & ~n11576;
  assign n11578 = ~n11382 & ~n11577;
  assign n11579 = ~n11379 & ~n11578;
  assign n11580 = n11355 & n11365;
  assign n11581 = ~n11355 & ~n11365;
  assign n11582 = ~n11580 & ~n11581;
  assign n11583 = ~n11579 & ~n11582;
  assign n11584 = ~n11366 & ~n11583;
  assign n11585 = n11342 & n11352;
  assign n11586 = ~n11342 & ~n11352;
  assign n11587 = ~n11585 & ~n11586;
  assign n11588 = ~n11584 & ~n11587;
  assign n11589 = ~n11353 & ~n11588;
  assign n11590 = ~n11329 & n11339;
  assign n11591 = ~n11340 & ~n11590;
  assign n11592 = ~n11589 & n11591;
  assign n11593 = ~n11340 & ~n11592;
  assign n11594 = ~n11327 & ~n11593;
  assign n11595 = ~n11324 & ~n11594;
  assign n11596 = n11307 & n11310;
  assign n11597 = ~n11311 & ~n11596;
  assign n11598 = ~n11595 & n11597;
  assign n11599 = ~n11311 & ~n11598;
  assign n11600 = ~n11297 & ~n11599;
  assign n11601 = ~n11294 & ~n11600;
  assign n11602 = n11270 & n11280;
  assign n11603 = ~n11270 & ~n11280;
  assign n11604 = ~n11602 & ~n11603;
  assign n11605 = ~n11601 & ~n11604;
  assign n11606 = ~n11281 & ~n11605;
  assign n11607 = n11257 & n11267;
  assign n11608 = ~n11257 & ~n11267;
  assign n11609 = ~n11607 & ~n11608;
  assign n11610 = ~n11606 & ~n11609;
  assign n11611 = ~n11268 & ~n11610;
  assign n11612 = ~n11244 & n11254;
  assign n11613 = ~n11255 & ~n11612;
  assign n11614 = ~n11611 & n11613;
  assign n11615 = ~n11255 & ~n11614;
  assign n11616 = n11238 & n11241;
  assign n11617 = ~n11242 & ~n11616;
  assign n11618 = ~n11615 & n11617;
  assign n11619 = ~n11242 & ~n11618;
  assign n11620 = ~n11228 & ~n11619;
  assign n11621 = ~n11225 & ~n11620;
  assign n11622 = ~n11212 & ~n11621;
  assign n11623 = ~n11209 & ~n11622;
  assign n11624 = n11185 & n11195;
  assign n11625 = ~n11185 & ~n11195;
  assign n11626 = ~n11624 & ~n11625;
  assign n11627 = ~n11623 & ~n11626;
  assign n11628 = ~n11196 & ~n11627;
  assign n11629 = ~n11172 & n11182;
  assign n11630 = ~n11183 & ~n11629;
  assign n11631 = ~n11628 & n11630;
  assign n11632 = ~n11183 & ~n11631;
  assign n11633 = ~n11170 & ~n11632;
  assign n11634 = ~n11167 & ~n11633;
  assign n11635 = n11150 & n11153;
  assign n11636 = ~n11154 & ~n11635;
  assign n11637 = ~n11634 & n11636;
  assign n11638 = ~n11154 & ~n11637;
  assign n11639 = n11136 & n11139;
  assign n11640 = ~n11140 & ~n11639;
  assign n11641 = ~n11638 & n11640;
  assign n11642 = ~n11140 & ~n11641;
  assign n11643 = ~n11126 & ~n11642;
  assign n11644 = ~n11123 & ~n11643;
  assign n11645 = ~n11110 & ~n11644;
  assign n11646 = ~n11107 & ~n11645;
  assign n11647 = n11090 & n11093;
  assign n11648 = ~n11094 & ~n11647;
  assign n11649 = ~n11646 & n11648;
  assign n11650 = ~n11094 & ~n11649;
  assign n11651 = ~n11073 & ~n11077;
  assign n11652 = n11076 & ~n11651;
  assign n11653 = ~n11076 & n11651;
  assign n11654 = ~n11652 & ~n11653;
  assign n11655 = ~n11650 & n11654;
  assign n11656 = n11650 & ~n11654;
  assign n11657 = ~n11655 & ~n11656;
  assign n11658 = n11646 & ~n11648;
  assign n11659 = ~n11649 & ~n11658;
  assign n11660 = ~n3855 & n11055;
  assign n11661 = ~pi0  & pi1 ;
  assign n11662 = ~n3883 & n11661;
  assign n11663 = ~n3900 & n11056;
  assign n11664 = ~n11660 & ~n11662;
  assign n11665 = ~n11663 & n11664;
  assign n11666 = pi2  & n11665;
  assign n11667 = ~pi2  & ~n11665;
  assign n11668 = ~n11666 & ~n11667;
  assign n11669 = n11659 & ~n11668;
  assign n11670 = n11110 & n11644;
  assign n11671 = ~n11645 & ~n11670;
  assign n11672 = pi0  & n11053;
  assign n11673 = ~n3883 & n11672;
  assign n11674 = n4399 & n11056;
  assign n11675 = ~n3855 & n11661;
  assign n11676 = ~n3681 & n11055;
  assign n11677 = ~n11673 & ~n11675;
  assign n11678 = ~n11676 & n11677;
  assign n11679 = ~n11674 & n11678;
  assign n11680 = pi2  & n11679;
  assign n11681 = ~pi2  & ~n11679;
  assign n11682 = ~n11680 & ~n11681;
  assign n11683 = n11671 & ~n11682;
  assign n11684 = n11126 & n11642;
  assign n11685 = ~n11643 & ~n11684;
  assign n11686 = ~n3855 & n11672;
  assign n11687 = n3972 & n11056;
  assign n11688 = ~n987 & n11055;
  assign n11689 = ~n3681 & n11661;
  assign n11690 = ~n11686 & ~n11688;
  assign n11691 = ~n11689 & n11690;
  assign n11692 = ~n11687 & n11691;
  assign n11693 = pi2  & n11692;
  assign n11694 = ~pi2  & ~n11692;
  assign n11695 = ~n11693 & ~n11694;
  assign n11696 = n11685 & ~n11695;
  assign n11697 = n11638 & ~n11640;
  assign n11698 = ~n11641 & ~n11697;
  assign n11699 = ~n878 & n11055;
  assign n11700 = n3687 & n11056;
  assign n11701 = ~n987 & n11661;
  assign n11702 = ~n3681 & n11672;
  assign n11703 = ~n11699 & ~n11701;
  assign n11704 = ~n11702 & n11703;
  assign n11705 = ~n11700 & n11704;
  assign n11706 = pi2  & n11705;
  assign n11707 = ~pi2  & ~n11705;
  assign n11708 = ~n11706 & ~n11707;
  assign n11709 = n11698 & ~n11708;
  assign n11710 = n11634 & ~n11636;
  assign n11711 = ~n11637 & ~n11710;
  assign n11712 = ~n987 & n11672;
  assign n11713 = n3791 & n11056;
  assign n11714 = ~n1104 & n11055;
  assign n11715 = ~n878 & n11661;
  assign n11716 = ~n11712 & ~n11714;
  assign n11717 = ~n11715 & n11716;
  assign n11718 = ~n11713 & n11717;
  assign n11719 = pi2  & n11718;
  assign n11720 = ~pi2  & ~n11718;
  assign n11721 = ~n11719 & ~n11720;
  assign n11722 = n11711 & ~n11721;
  assign n11723 = n11711 & n11721;
  assign n11724 = ~n11711 & ~n11721;
  assign n11725 = ~n11723 & ~n11724;
  assign n11726 = ~n1104 & n11661;
  assign n11727 = n3775 & n11056;
  assign n11728 = ~n1225 & n11055;
  assign n11729 = ~n878 & n11672;
  assign n11730 = ~n11726 & ~n11728;
  assign n11731 = ~n11729 & n11730;
  assign n11732 = ~n11727 & n11731;
  assign n11733 = pi2  & n11732;
  assign n11734 = ~pi2  & ~n11732;
  assign n11735 = ~n11733 & ~n11734;
  assign n11736 = n11628 & ~n11630;
  assign n11737 = ~n11631 & ~n11736;
  assign n11738 = n11623 & n11626;
  assign n11739 = ~n11627 & ~n11738;
  assign n11740 = ~n1448 & n11661;
  assign n11741 = n4453 & n11056;
  assign n11742 = ~n1533 & n11055;
  assign n11743 = ~n1345 & n11672;
  assign n11744 = ~n11740 & ~n11742;
  assign n11745 = ~n11743 & n11744;
  assign n11746 = ~n11741 & n11745;
  assign n11747 = pi2  & n11746;
  assign n11748 = ~pi2  & ~n11746;
  assign n11749 = ~n11747 & ~n11748;
  assign n11750 = ~n1533 & n11661;
  assign n11751 = n4355 & n11056;
  assign n11752 = ~n1637 & n11055;
  assign n11753 = ~n1448 & n11672;
  assign n11754 = ~n11750 & ~n11752;
  assign n11755 = ~n11753 & n11754;
  assign n11756 = ~n11751 & n11755;
  assign n11757 = pi2  & n11756;
  assign n11758 = ~pi2  & ~n11756;
  assign n11759 = ~n11757 & ~n11758;
  assign n11760 = ~n1637 & n11661;
  assign n11761 = n4553 & n11056;
  assign n11762 = ~n1717 & n11055;
  assign n11763 = ~n1533 & n11672;
  assign n11764 = ~n11760 & ~n11762;
  assign n11765 = ~n11763 & n11764;
  assign n11766 = ~n11761 & n11765;
  assign n11767 = pi2  & n11766;
  assign n11768 = ~pi2  & ~n11766;
  assign n11769 = ~n11767 & ~n11768;
  assign n11770 = n11611 & ~n11613;
  assign n11771 = ~n11614 & ~n11770;
  assign n11772 = n11606 & n11609;
  assign n11773 = ~n11610 & ~n11772;
  assign n11774 = n11601 & n11604;
  assign n11775 = ~n11605 & ~n11774;
  assign n11776 = ~n1998 & n11661;
  assign n11777 = n5151 & n11056;
  assign n11778 = ~n2098 & n11055;
  assign n11779 = ~n1908 & n11672;
  assign n11780 = ~n11776 & ~n11778;
  assign n11781 = ~n11779 & n11780;
  assign n11782 = ~n11777 & n11781;
  assign n11783 = pi2  & n11782;
  assign n11784 = ~pi2  & ~n11782;
  assign n11785 = ~n11783 & ~n11784;
  assign n11786 = ~n2098 & n11661;
  assign n11787 = n4979 & n11056;
  assign n11788 = ~n2146 & n11055;
  assign n11789 = ~n1998 & n11672;
  assign n11790 = ~n11786 & ~n11788;
  assign n11791 = ~n11789 & n11790;
  assign n11792 = ~n11787 & n11791;
  assign n11793 = pi2  & n11792;
  assign n11794 = ~pi2  & ~n11792;
  assign n11795 = ~n11793 & ~n11794;
  assign n11796 = ~n2098 & n11672;
  assign n11797 = n5359 & n11056;
  assign n11798 = ~n2146 & n11661;
  assign n11799 = ~n2249 & n11055;
  assign n11800 = ~n11796 & ~n11798;
  assign n11801 = ~n11799 & n11800;
  assign n11802 = ~n11797 & n11801;
  assign n11803 = pi2  & n11802;
  assign n11804 = ~pi2  & ~n11802;
  assign n11805 = ~n11803 & ~n11804;
  assign n11806 = n11589 & ~n11591;
  assign n11807 = ~n11592 & ~n11806;
  assign n11808 = n11584 & n11587;
  assign n11809 = ~n11588 & ~n11808;
  assign n11810 = n11579 & n11582;
  assign n11811 = ~n11583 & ~n11810;
  assign n11812 = ~n2589 & n11055;
  assign n11813 = n6016 & n11056;
  assign n11814 = ~n2496 & n11661;
  assign n11815 = ~n2412 & n11672;
  assign n11816 = ~n11812 & ~n11814;
  assign n11817 = ~n11815 & n11816;
  assign n11818 = ~n11813 & n11817;
  assign n11819 = pi2  & n11818;
  assign n11820 = ~pi2  & ~n11818;
  assign n11821 = ~n11819 & ~n11820;
  assign n11822 = ~n2496 & n11672;
  assign n11823 = n5776 & n11056;
  assign n11824 = ~n2674 & n11055;
  assign n11825 = ~n2589 & n11661;
  assign n11826 = ~n11822 & ~n11824;
  assign n11827 = ~n11825 & n11826;
  assign n11828 = ~n11823 & n11827;
  assign n11829 = pi2  & n11828;
  assign n11830 = ~pi2  & ~n11828;
  assign n11831 = ~n11829 & ~n11830;
  assign n11832 = ~n2674 & n11661;
  assign n11833 = n6240 & n11056;
  assign n11834 = ~n2708 & n11055;
  assign n11835 = ~n2589 & n11672;
  assign n11836 = ~n11832 & ~n11834;
  assign n11837 = ~n11835 & n11836;
  assign n11838 = ~n11833 & n11837;
  assign n11839 = pi2  & n11838;
  assign n11840 = ~pi2  & ~n11838;
  assign n11841 = ~n11839 & ~n11840;
  assign n11842 = n11567 & ~n11569;
  assign n11843 = ~n11570 & ~n11842;
  assign n11844 = n11562 & n11565;
  assign n11845 = ~n11566 & ~n11844;
  assign n11846 = n11557 & n11560;
  assign n11847 = ~n11561 & ~n11846;
  assign n11848 = ~n2919 & n11661;
  assign n11849 = n6809 & n11056;
  assign n11850 = ~n2951 & n11055;
  assign n11851 = ~n2835 & n11672;
  assign n11852 = ~n11848 & ~n11850;
  assign n11853 = ~n11851 & n11852;
  assign n11854 = ~n11849 & n11853;
  assign n11855 = pi2  & n11854;
  assign n11856 = ~pi2  & ~n11854;
  assign n11857 = ~n11855 & ~n11856;
  assign n11858 = ~n2919 & n11672;
  assign n11859 = n6821 & n11056;
  assign n11860 = ~n2951 & n11661;
  assign n11861 = ~n3031 & n11055;
  assign n11862 = ~n11858 & ~n11860;
  assign n11863 = ~n11861 & n11862;
  assign n11864 = ~n11859 & n11863;
  assign n11865 = pi2  & n11864;
  assign n11866 = ~pi2  & ~n11864;
  assign n11867 = ~n11865 & ~n11866;
  assign n11868 = ~n2951 & n11672;
  assign n11869 = n6486 & n11056;
  assign n11870 = ~n3118 & n11055;
  assign n11871 = ~n3031 & n11661;
  assign n11872 = ~n11868 & ~n11870;
  assign n11873 = ~n11871 & n11872;
  assign n11874 = ~n11869 & n11873;
  assign n11875 = pi2  & n11874;
  assign n11876 = ~pi2  & ~n11874;
  assign n11877 = ~n11875 & ~n11876;
  assign n11878 = n11545 & ~n11547;
  assign n11879 = ~n11548 & ~n11878;
  assign n11880 = ~n3118 & n11672;
  assign n11881 = n6908 & n11056;
  assign n11882 = ~n3241 & n11055;
  assign n11883 = ~n3182 & n11661;
  assign n11884 = ~n11880 & ~n11882;
  assign n11885 = ~n11883 & n11884;
  assign n11886 = ~n11881 & n11885;
  assign n11887 = pi2  & n11886;
  assign n11888 = ~pi2  & ~n11886;
  assign n11889 = ~n11887 & ~n11888;
  assign n11890 = pi5  & ~n11521;
  assign n11891 = n11528 & ~n11890;
  assign n11892 = ~n11528 & n11890;
  assign n11893 = ~n11891 & ~n11892;
  assign n11894 = ~n3241 & n11672;
  assign n11895 = n7004 & n11056;
  assign n11896 = ~n3275 & n11661;
  assign n11897 = ~n3370 & n11055;
  assign n11898 = ~n11894 & ~n11896;
  assign n11899 = ~n11897 & n11898;
  assign n11900 = ~n11895 & n11899;
  assign n11901 = pi2  & n11900;
  assign n11902 = ~pi2  & ~n11900;
  assign n11903 = ~n11901 & ~n11902;
  assign n11904 = ~n3485 & n11672;
  assign n11905 = ~n3427 & n11055;
  assign n11906 = ~n3485 & n11661;
  assign n11907 = ~n3370 & n11672;
  assign n11908 = ~n11905 & ~n11906;
  assign n11909 = ~n11907 & n11908;
  assign n11910 = pi2  & ~n11909;
  assign n11911 = pi2  & n11056;
  assign n11912 = n7045 & n11911;
  assign n11913 = ~n7720 & n11911;
  assign n11914 = pi2  & n11661;
  assign n11915 = ~pi0  & ~n11914;
  assign n11916 = ~n3427 & ~n11915;
  assign n11917 = pi2  & ~n11904;
  assign n11918 = ~n11916 & n11917;
  assign n11919 = ~n11913 & n11918;
  assign n11920 = ~n11910 & n11919;
  assign n11921 = ~n11912 & n11920;
  assign n11922 = ~n11514 & ~n11921;
  assign n11923 = n11514 & n11921;
  assign n11924 = ~n3275 & n11672;
  assign n11925 = n7102 & n11056;
  assign n11926 = ~n3485 & n11055;
  assign n11927 = ~n3370 & n11661;
  assign n11928 = ~n11924 & ~n11926;
  assign n11929 = ~n11927 & n11928;
  assign n11930 = ~n11925 & n11929;
  assign n11931 = pi2  & ~n11930;
  assign n11932 = ~pi2  & n11930;
  assign n11933 = ~n11931 & ~n11932;
  assign n11934 = ~n11923 & ~n11933;
  assign n11935 = ~n11922 & ~n11934;
  assign n11936 = ~n11903 & n11935;
  assign n11937 = n11903 & ~n11935;
  assign n11938 = pi5  & n11514;
  assign n11939 = ~n11519 & n11938;
  assign n11940 = n11519 & ~n11938;
  assign n11941 = ~n11939 & ~n11940;
  assign n11942 = ~n11937 & n11941;
  assign n11943 = ~n11936 & ~n11942;
  assign n11944 = n11893 & ~n11943;
  assign n11945 = ~n11893 & n11943;
  assign n11946 = ~n3275 & n11055;
  assign n11947 = n6959 & n11056;
  assign n11948 = ~n3241 & n11661;
  assign n11949 = ~n3182 & n11672;
  assign n11950 = ~n11946 & ~n11948;
  assign n11951 = ~n11949 & n11950;
  assign n11952 = ~n11947 & n11951;
  assign n11953 = pi2  & ~n11952;
  assign n11954 = ~pi2  & n11952;
  assign n11955 = ~n11953 & ~n11954;
  assign n11956 = ~n11945 & n11955;
  assign n11957 = ~n11944 & ~n11956;
  assign n11958 = ~n11889 & ~n11957;
  assign n11959 = n11889 & n11957;
  assign n11960 = n11533 & n11543;
  assign n11961 = ~n11544 & ~n11960;
  assign n11962 = ~n11959 & n11961;
  assign n11963 = ~n11958 & ~n11962;
  assign n11964 = n11879 & ~n11963;
  assign n11965 = ~n11879 & n11963;
  assign n11966 = ~n3182 & n11055;
  assign n11967 = n6863 & n11056;
  assign n11968 = ~n3118 & n11661;
  assign n11969 = ~n3031 & n11672;
  assign n11970 = ~n11966 & ~n11968;
  assign n11971 = ~n11969 & n11970;
  assign n11972 = ~n11967 & n11971;
  assign n11973 = pi2  & ~n11972;
  assign n11974 = ~pi2  & n11972;
  assign n11975 = ~n11973 & ~n11974;
  assign n11976 = ~n11965 & n11975;
  assign n11977 = ~n11964 & ~n11976;
  assign n11978 = ~n11877 & ~n11977;
  assign n11979 = n11877 & n11977;
  assign n11980 = n11498 & n11549;
  assign n11981 = ~n11550 & ~n11980;
  assign n11982 = ~n11979 & n11981;
  assign n11983 = ~n11978 & ~n11982;
  assign n11984 = ~n11867 & ~n11983;
  assign n11985 = n11867 & n11983;
  assign n11986 = n11551 & ~n11553;
  assign n11987 = ~n11554 & ~n11986;
  assign n11988 = ~n11985 & n11987;
  assign n11989 = ~n11984 & ~n11988;
  assign n11990 = ~n11857 & ~n11989;
  assign n11991 = n11857 & n11989;
  assign n11992 = n11467 & n11555;
  assign n11993 = ~n11556 & ~n11992;
  assign n11994 = ~n11991 & n11993;
  assign n11995 = ~n11990 & ~n11994;
  assign n11996 = n11847 & ~n11995;
  assign n11997 = ~n11847 & n11995;
  assign n11998 = ~n2919 & n11055;
  assign n11999 = n6509 & n11056;
  assign n12000 = ~n2835 & n11661;
  assign n12001 = ~n2778 & n11672;
  assign n12002 = ~n11998 & ~n12000;
  assign n12003 = ~n12001 & n12002;
  assign n12004 = ~n11999 & n12003;
  assign n12005 = pi2  & ~n12004;
  assign n12006 = ~pi2  & n12004;
  assign n12007 = ~n12005 & ~n12006;
  assign n12008 = ~n11997 & n12007;
  assign n12009 = ~n11996 & ~n12008;
  assign n12010 = n11845 & ~n12009;
  assign n12011 = ~n11845 & n12009;
  assign n12012 = ~n2708 & n11672;
  assign n12013 = n6222 & n11056;
  assign n12014 = ~n2835 & n11055;
  assign n12015 = ~n2778 & n11661;
  assign n12016 = ~n12012 & ~n12014;
  assign n12017 = ~n12015 & n12016;
  assign n12018 = ~n12013 & n12017;
  assign n12019 = pi2  & ~n12018;
  assign n12020 = ~pi2  & n12018;
  assign n12021 = ~n12019 & ~n12020;
  assign n12022 = ~n12011 & n12021;
  assign n12023 = ~n12010 & ~n12022;
  assign n12024 = n11843 & ~n12023;
  assign n12025 = ~n11843 & n12023;
  assign n12026 = ~n2778 & n11055;
  assign n12027 = n6393 & n11056;
  assign n12028 = ~n2708 & n11661;
  assign n12029 = ~n2674 & n11672;
  assign n12030 = ~n12026 & ~n12028;
  assign n12031 = ~n12029 & n12030;
  assign n12032 = ~n12027 & n12031;
  assign n12033 = pi2  & ~n12032;
  assign n12034 = ~pi2  & n12032;
  assign n12035 = ~n12033 & ~n12034;
  assign n12036 = ~n12025 & n12035;
  assign n12037 = ~n12024 & ~n12036;
  assign n12038 = ~n11841 & ~n12037;
  assign n12039 = n11841 & n12037;
  assign n12040 = n11571 & ~n11573;
  assign n12041 = ~n11574 & ~n12040;
  assign n12042 = ~n12039 & n12041;
  assign n12043 = ~n12038 & ~n12042;
  assign n12044 = ~n11831 & ~n12043;
  assign n12045 = n11831 & n12043;
  assign n12046 = n11398 & n11575;
  assign n12047 = ~n11576 & ~n12046;
  assign n12048 = ~n12045 & n12047;
  assign n12049 = ~n12044 & ~n12048;
  assign n12050 = ~n11821 & ~n12049;
  assign n12051 = n11821 & n12049;
  assign n12052 = n11382 & n11577;
  assign n12053 = ~n11578 & ~n12052;
  assign n12054 = ~n12051 & n12053;
  assign n12055 = ~n12050 & ~n12054;
  assign n12056 = n11811 & ~n12055;
  assign n12057 = ~n11811 & n12055;
  assign n12058 = ~n2347 & n11672;
  assign n12059 = n5596 & n11056;
  assign n12060 = ~n2496 & n11055;
  assign n12061 = ~n2412 & n11661;
  assign n12062 = ~n12058 & ~n12060;
  assign n12063 = ~n12061 & n12062;
  assign n12064 = ~n12059 & n12063;
  assign n12065 = pi2  & ~n12064;
  assign n12066 = ~pi2  & n12064;
  assign n12067 = ~n12065 & ~n12066;
  assign n12068 = ~n12057 & n12067;
  assign n12069 = ~n12056 & ~n12068;
  assign n12070 = n11809 & ~n12069;
  assign n12071 = ~n11809 & n12069;
  assign n12072 = ~n2412 & n11055;
  assign n12073 = n5579 & n11056;
  assign n12074 = ~n2347 & n11661;
  assign n12075 = ~n2249 & n11672;
  assign n12076 = ~n12072 & ~n12074;
  assign n12077 = ~n12075 & n12076;
  assign n12078 = ~n12073 & n12077;
  assign n12079 = pi2  & ~n12078;
  assign n12080 = ~pi2  & n12078;
  assign n12081 = ~n12079 & ~n12080;
  assign n12082 = ~n12071 & n12081;
  assign n12083 = ~n12070 & ~n12082;
  assign n12084 = n11807 & ~n12083;
  assign n12085 = ~n11807 & n12083;
  assign n12086 = ~n2146 & n11672;
  assign n12087 = n5343 & n11056;
  assign n12088 = ~n2347 & n11055;
  assign n12089 = ~n2249 & n11661;
  assign n12090 = ~n12086 & ~n12088;
  assign n12091 = ~n12089 & n12090;
  assign n12092 = ~n12087 & n12091;
  assign n12093 = pi2  & ~n12092;
  assign n12094 = ~pi2  & n12092;
  assign n12095 = ~n12093 & ~n12094;
  assign n12096 = ~n12085 & n12095;
  assign n12097 = ~n12084 & ~n12096;
  assign n12098 = ~n11805 & ~n12097;
  assign n12099 = n11805 & n12097;
  assign n12100 = n11327 & n11593;
  assign n12101 = ~n11594 & ~n12100;
  assign n12102 = ~n12099 & n12101;
  assign n12103 = ~n12098 & ~n12102;
  assign n12104 = ~n11795 & ~n12103;
  assign n12105 = n11795 & n12103;
  assign n12106 = n11595 & ~n11597;
  assign n12107 = ~n11598 & ~n12106;
  assign n12108 = ~n12105 & n12107;
  assign n12109 = ~n12104 & ~n12108;
  assign n12110 = ~n11785 & ~n12109;
  assign n12111 = n11785 & n12109;
  assign n12112 = n11297 & n11599;
  assign n12113 = ~n11600 & ~n12112;
  assign n12114 = ~n12111 & n12113;
  assign n12115 = ~n12110 & ~n12114;
  assign n12116 = n11775 & ~n12115;
  assign n12117 = ~n11775 & n12115;
  assign n12118 = ~n1908 & n11661;
  assign n12119 = n4779 & n11056;
  assign n12120 = ~n1998 & n11055;
  assign n12121 = ~n1841 & n11672;
  assign n12122 = ~n12118 & ~n12120;
  assign n12123 = ~n12121 & n12122;
  assign n12124 = ~n12119 & n12123;
  assign n12125 = pi2  & ~n12124;
  assign n12126 = ~pi2  & n12124;
  assign n12127 = ~n12125 & ~n12126;
  assign n12128 = ~n12117 & n12127;
  assign n12129 = ~n12116 & ~n12128;
  assign n12130 = n11773 & ~n12129;
  assign n12131 = ~n11773 & n12129;
  assign n12132 = ~n1841 & n11661;
  assign n12133 = n4762 & n11056;
  assign n12134 = ~n1908 & n11055;
  assign n12135 = ~n1717 & n11672;
  assign n12136 = ~n12132 & ~n12134;
  assign n12137 = ~n12135 & n12136;
  assign n12138 = ~n12133 & n12137;
  assign n12139 = pi2  & ~n12138;
  assign n12140 = ~pi2  & n12138;
  assign n12141 = ~n12139 & ~n12140;
  assign n12142 = ~n12131 & n12141;
  assign n12143 = ~n12130 & ~n12142;
  assign n12144 = n11771 & ~n12143;
  assign n12145 = ~n11771 & n12143;
  assign n12146 = ~n1717 & n11661;
  assign n12147 = n4537 & n11056;
  assign n12148 = ~n1841 & n11055;
  assign n12149 = ~n1637 & n11672;
  assign n12150 = ~n12146 & ~n12148;
  assign n12151 = ~n12149 & n12150;
  assign n12152 = ~n12147 & n12151;
  assign n12153 = pi2  & ~n12152;
  assign n12154 = ~pi2  & n12152;
  assign n12155 = ~n12153 & ~n12154;
  assign n12156 = ~n12145 & n12155;
  assign n12157 = ~n12144 & ~n12156;
  assign n12158 = ~n11769 & ~n12157;
  assign n12159 = n11769 & n12157;
  assign n12160 = n11615 & ~n11617;
  assign n12161 = ~n11618 & ~n12160;
  assign n12162 = ~n12159 & n12161;
  assign n12163 = ~n12158 & ~n12162;
  assign n12164 = ~n11759 & ~n12163;
  assign n12165 = n11759 & n12163;
  assign n12166 = n11228 & n11619;
  assign n12167 = ~n11620 & ~n12166;
  assign n12168 = ~n12165 & n12167;
  assign n12169 = ~n12164 & ~n12168;
  assign n12170 = ~n11749 & ~n12169;
  assign n12171 = n11749 & n12169;
  assign n12172 = n11212 & n11621;
  assign n12173 = ~n11622 & ~n12172;
  assign n12174 = ~n12171 & n12173;
  assign n12175 = ~n12170 & ~n12174;
  assign n12176 = n11739 & ~n12175;
  assign n12177 = ~n11739 & n12175;
  assign n12178 = ~n1345 & n11661;
  assign n12179 = n4152 & n11056;
  assign n12180 = ~n1448 & n11055;
  assign n12181 = ~n1225 & n11672;
  assign n12182 = ~n12178 & ~n12180;
  assign n12183 = ~n12181 & n12182;
  assign n12184 = ~n12179 & n12183;
  assign n12185 = pi2  & ~n12184;
  assign n12186 = ~pi2  & n12184;
  assign n12187 = ~n12185 & ~n12186;
  assign n12188 = ~n12177 & n12187;
  assign n12189 = ~n12176 & ~n12188;
  assign n12190 = n11737 & ~n12189;
  assign n12191 = ~n11737 & n12189;
  assign n12192 = ~n1225 & n11661;
  assign n12193 = n4135 & n11056;
  assign n12194 = ~n1345 & n11055;
  assign n12195 = ~n1104 & n11672;
  assign n12196 = ~n12192 & ~n12194;
  assign n12197 = ~n12195 & n12196;
  assign n12198 = ~n12193 & n12197;
  assign n12199 = pi2  & ~n12198;
  assign n12200 = ~pi2  & n12198;
  assign n12201 = ~n12199 & ~n12200;
  assign n12202 = ~n12191 & n12201;
  assign n12203 = ~n12190 & ~n12202;
  assign n12204 = ~n11735 & ~n12203;
  assign n12205 = n11735 & n12203;
  assign n12206 = n11170 & n11632;
  assign n12207 = ~n11633 & ~n12206;
  assign n12208 = ~n12205 & n12207;
  assign n12209 = ~n12204 & ~n12208;
  assign n12210 = ~n11725 & ~n12209;
  assign n12211 = ~n11722 & ~n12210;
  assign n12212 = ~n11698 & n11708;
  assign n12213 = ~n11709 & ~n12212;
  assign n12214 = ~n12211 & n12213;
  assign n12215 = ~n11709 & ~n12214;
  assign n12216 = ~n11685 & n11695;
  assign n12217 = ~n11696 & ~n12216;
  assign n12218 = ~n12215 & n12217;
  assign n12219 = ~n11696 & ~n12218;
  assign n12220 = ~n11671 & n11682;
  assign n12221 = ~n11683 & ~n12220;
  assign n12222 = ~n12219 & n12221;
  assign n12223 = ~n11683 & ~n12222;
  assign n12224 = ~n11659 & n11668;
  assign n12225 = ~n11669 & ~n12224;
  assign n12226 = ~n12223 & n12225;
  assign n12227 = ~n11669 & ~n12226;
  assign n12228 = n11657 & ~n12227;
  assign n12229 = ~n11655 & ~n12228;
  assign n12230 = ~n11050 & n11079;
  assign n12231 = ~n11080 & ~n12230;
  assign n12232 = ~n12229 & n12231;
  assign n12233 = ~n11080 & ~n12232;
  assign n12234 = n11045 & ~n11047;
  assign n12235 = ~n11048 & ~n12234;
  assign n12236 = ~n12233 & n12235;
  assign n12237 = ~n11048 & ~n12236;
  assign n12238 = n10492 & ~n12237;
  assign n12239 = ~n10490 & ~n12238;
  assign n12240 = ~n9490 & n9968;
  assign n12241 = ~n9969 & ~n12240;
  assign n12242 = ~n12239 & n12241;
  assign n12243 = ~n9969 & ~n12242;
  assign n12244 = n9485 & ~n9487;
  assign n12245 = ~n9488 & ~n12244;
  assign n12246 = ~n12243 & n12245;
  assign n12247 = ~n9488 & ~n12246;
  assign n12248 = n9039 & ~n12247;
  assign n12249 = ~n9037 & ~n12248;
  assign n12250 = n8623 & ~n12249;
  assign n12251 = ~n8621 & ~n12250;
  assign n12252 = ~n7894 & n8234;
  assign n12253 = ~n8235 & ~n12252;
  assign n12254 = ~n12251 & n12253;
  assign n12255 = ~n8235 & ~n12254;
  assign n12256 = n7892 & ~n12255;
  assign n12257 = ~n7890 & ~n12256;
  assign n12258 = ~n7419 & n7579;
  assign n12259 = ~n7580 & ~n12258;
  assign n12260 = ~n12257 & n12259;
  assign n12261 = ~n7580 & ~n12260;
  assign n12262 = n7414 & ~n7416;
  assign n12263 = ~n7417 & ~n12262;
  assign n12264 = ~n12261 & n12263;
  assign n12265 = ~n7417 & ~n12264;
  assign n12266 = n7261 & ~n12265;
  assign n12267 = ~n7259 & ~n12266;
  assign n12268 = n6762 & ~n12267;
  assign n12269 = ~n6760 & ~n12268;
  assign n12270 = n6617 & ~n12269;
  assign n12271 = ~n6615 & ~n12270;
  assign n12272 = n6335 & ~n12271;
  assign n12273 = ~n6333 & ~n12272;
  assign n12274 = ~n5971 & n6110;
  assign n12275 = ~n6111 & ~n12274;
  assign n12276 = ~n12273 & n12275;
  assign n12277 = ~n6111 & ~n12276;
  assign n12278 = n5969 & ~n12277;
  assign n12279 = ~n5967 & ~n12278;
  assign n12280 = n5865 & ~n12279;
  assign n12281 = ~n5863 & ~n12280;
  assign n12282 = n5429 & ~n12281;
  assign n12283 = ~n5427 & ~n12282;
  assign n12284 = ~n5129 & n5224;
  assign n12285 = ~n5225 & ~n12284;
  assign n12286 = ~n12283 & n12285;
  assign n12287 = ~n5225 & ~n12286;
  assign n12288 = n5127 & ~n12287;
  assign n12289 = ~n5125 & ~n12288;
  assign n12290 = ~n4666 & ~n5059;
  assign n12291 = ~n5060 & ~n12290;
  assign n12292 = ~n12289 & n12291;
  assign n12293 = ~n5060 & ~n12292;
  assign n12294 = n4661 & ~n4663;
  assign n12295 = ~n4664 & ~n12294;
  assign n12296 = ~n12293 & n12295;
  assign n12297 = ~n4664 & ~n12296;
  assign n12298 = n4611 & ~n4613;
  assign n12299 = ~n4614 & ~n12298;
  assign n12300 = ~n12297 & n12299;
  assign n12301 = ~n4614 & ~n12300;
  assign n12302 = n4443 & ~n4445;
  assign n12303 = ~n4446 & ~n12302;
  assign n12304 = ~n12301 & n12303;
  assign n12305 = ~n4446 & ~n12304;
  assign n12306 = n4419 & ~n12305;
  assign n12307 = ~n4417 & ~n12306;
  assign n12308 = n3908 & n3984;
  assign n12309 = ~n3985 & ~n12308;
  assign n12310 = ~n12307 & n12309;
  assign n12311 = ~n3985 & ~n12310;
  assign n12312 = ~n3956 & ~n3961;
  assign n12313 = ~n212 & ~n1699;
  assign n12314 = n1308 & n12313;
  assign n12315 = n2658 & n12314;
  assign n12316 = n3629 & n12315;
  assign n12317 = ~n163 & ~n432;
  assign n12318 = n719 & ~n724;
  assign n12319 = n3619 & n12318;
  assign n12320 = n1170 & n1535;
  assign n12321 = n12319 & n12320;
  assign n12322 = n5523 & n7083;
  assign n12323 = n973 & n12322;
  assign n12324 = ~n168 & n900;
  assign n12325 = n2197 & n2284;
  assign n12326 = n2502 & n12317;
  assign n12327 = n12325 & n12326;
  assign n12328 = n12324 & n12327;
  assign n12329 = n12321 & n12328;
  assign n12330 = n891 & n12329;
  assign n12331 = n3638 & n12316;
  assign n12332 = n12330 & n12331;
  assign n12333 = n12323 & n12332;
  assign n12334 = ~n3955 & ~n12333;
  assign n12335 = n3955 & n12333;
  assign n12336 = ~pi29  & ~n12334;
  assign n12337 = ~n12335 & n12336;
  assign n12338 = ~pi29  & ~n12337;
  assign n12339 = ~n12334 & ~n12337;
  assign n12340 = ~n12335 & n12339;
  assign n12341 = ~n12338 & ~n12340;
  assign n12342 = ~n12312 & ~n12341;
  assign n12343 = n12312 & n12341;
  assign n12344 = ~n12342 & ~n12343;
  assign n12345 = n3694 & ~n3883;
  assign n12346 = n880 & n4399;
  assign n12347 = n3692 & ~n3855;
  assign n12348 = n748 & ~n3681;
  assign n12349 = ~n12345 & ~n12347;
  assign n12350 = ~n12348 & n12349;
  assign n12351 = ~n12346 & n12350;
  assign n12352 = n12344 & ~n12351;
  assign n12353 = ~n12344 & n12351;
  assign n12354 = ~n12352 & ~n12353;
  assign n12355 = ~n3963 & ~n3979;
  assign n12356 = ~n3980 & ~n12355;
  assign n12357 = n12354 & n12356;
  assign n12358 = ~n12354 & ~n12356;
  assign n12359 = ~n12357 & ~n12358;
  assign n12360 = ~n12311 & n12359;
  assign n12361 = n12311 & ~n12359;
  assign n12362 = ~n12360 & ~n12361;
  assign n12363 = n86 & n12362;
  assign n12364 = ~n12342 & ~n12352;
  assign n12365 = ~n427 & n3325;
  assign n12366 = n903 & n12365;
  assign n12367 = n934 & n2954;
  assign n12368 = n12366 & n12367;
  assign n12369 = n3830 & n12368;
  assign n12370 = n3867 & n5686;
  assign n12371 = n12369 & n12370;
  assign n12372 = n1185 & n12316;
  assign n12373 = n12371 & n12372;
  assign n12374 = n3660 & n12373;
  assign n12375 = ~n12339 & n12374;
  assign n12376 = n12339 & ~n12374;
  assign n12377 = ~n12375 & ~n12376;
  assign n12378 = n748 & ~n3855;
  assign n12379 = n3692 & ~n3883;
  assign n12380 = n880 & ~n3900;
  assign n12381 = ~n12378 & ~n12379;
  assign n12382 = ~n12380 & n12381;
  assign n12383 = n12377 & ~n12382;
  assign n12384 = ~n12377 & n12382;
  assign n12385 = ~n12383 & ~n12384;
  assign n12386 = ~n12364 & n12385;
  assign n12387 = n12364 & ~n12385;
  assign n12388 = ~n12386 & ~n12387;
  assign n12389 = ~n12357 & ~n12360;
  assign n12390 = n12388 & ~n12389;
  assign n12391 = ~n12388 & n12389;
  assign n12392 = ~n12390 & ~n12391;
  assign n12393 = n12362 & n12392;
  assign n12394 = n12307 & ~n12309;
  assign n12395 = ~n12310 & ~n12394;
  assign n12396 = n12362 & n12395;
  assign n12397 = ~n4419 & n12305;
  assign n12398 = ~n12306 & ~n12397;
  assign n12399 = n12395 & n12398;
  assign n12400 = n12301 & ~n12303;
  assign n12401 = ~n12304 & ~n12400;
  assign n12402 = n12398 & n12401;
  assign n12403 = n12297 & ~n12299;
  assign n12404 = ~n12300 & ~n12403;
  assign n12405 = n12401 & n12404;
  assign n12406 = n12293 & ~n12295;
  assign n12407 = ~n12296 & ~n12406;
  assign n12408 = n12404 & n12407;
  assign n12409 = n12289 & ~n12291;
  assign n12410 = ~n12292 & ~n12409;
  assign n12411 = n12407 & n12410;
  assign n12412 = ~n5127 & n12287;
  assign n12413 = ~n12288 & ~n12412;
  assign n12414 = n12410 & n12413;
  assign n12415 = n12283 & ~n12285;
  assign n12416 = ~n12286 & ~n12415;
  assign n12417 = n12413 & n12416;
  assign n12418 = ~n5429 & n12281;
  assign n12419 = ~n12282 & ~n12418;
  assign n12420 = n12416 & n12419;
  assign n12421 = ~n5865 & n12279;
  assign n12422 = ~n12280 & ~n12421;
  assign n12423 = n12419 & n12422;
  assign n12424 = ~n5969 & n12277;
  assign n12425 = ~n12278 & ~n12424;
  assign n12426 = n12422 & n12425;
  assign n12427 = n12273 & ~n12275;
  assign n12428 = ~n12276 & ~n12427;
  assign n12429 = n12425 & n12428;
  assign n12430 = ~n6335 & n12271;
  assign n12431 = ~n12272 & ~n12430;
  assign n12432 = n12428 & n12431;
  assign n12433 = ~n6617 & n12269;
  assign n12434 = ~n12270 & ~n12433;
  assign n12435 = n12431 & n12434;
  assign n12436 = ~n6762 & n12267;
  assign n12437 = ~n12268 & ~n12436;
  assign n12438 = n12434 & n12437;
  assign n12439 = ~n7261 & n12265;
  assign n12440 = ~n12266 & ~n12439;
  assign n12441 = n12437 & n12440;
  assign n12442 = n12261 & ~n12263;
  assign n12443 = ~n12264 & ~n12442;
  assign n12444 = n12440 & n12443;
  assign n12445 = n12257 & ~n12259;
  assign n12446 = ~n12260 & ~n12445;
  assign n12447 = n12443 & n12446;
  assign n12448 = ~n7892 & n12255;
  assign n12449 = ~n12256 & ~n12448;
  assign n12450 = n12446 & n12449;
  assign n12451 = n12251 & ~n12253;
  assign n12452 = ~n12254 & ~n12451;
  assign n12453 = n12449 & n12452;
  assign n12454 = ~n8623 & n12249;
  assign n12455 = ~n12250 & ~n12454;
  assign n12456 = n12452 & n12455;
  assign n12457 = ~n9039 & n12247;
  assign n12458 = ~n12248 & ~n12457;
  assign n12459 = n12455 & n12458;
  assign n12460 = n12243 & ~n12245;
  assign n12461 = ~n12246 & ~n12460;
  assign n12462 = n12458 & n12461;
  assign n12463 = n12239 & ~n12241;
  assign n12464 = ~n12242 & ~n12463;
  assign n12465 = n12461 & n12464;
  assign n12466 = ~n10492 & n12237;
  assign n12467 = ~n12238 & ~n12466;
  assign n12468 = n12464 & n12467;
  assign n12469 = n12233 & ~n12235;
  assign n12470 = ~n12236 & ~n12469;
  assign n12471 = n12467 & n12470;
  assign n12472 = n12229 & ~n12231;
  assign n12473 = ~n12232 & ~n12472;
  assign n12474 = n12470 & n12473;
  assign n12475 = ~n11657 & n12227;
  assign n12476 = ~n12228 & ~n12475;
  assign n12477 = n12473 & n12476;
  assign n12478 = n12223 & ~n12225;
  assign n12479 = ~n12226 & ~n12478;
  assign n12480 = n12476 & n12479;
  assign n12481 = n12219 & ~n12221;
  assign n12482 = ~n12222 & ~n12481;
  assign n12483 = n12479 & n12482;
  assign n12484 = n12215 & ~n12217;
  assign n12485 = ~n12218 & ~n12484;
  assign n12486 = n12482 & n12485;
  assign n12487 = ~n12482 & ~n12485;
  assign n12488 = ~n12486 & ~n12487;
  assign n12489 = n12211 & ~n12213;
  assign n12490 = ~n12214 & ~n12489;
  assign n12491 = n11725 & n12209;
  assign n12492 = ~n12210 & ~n12491;
  assign n12493 = ~n12485 & ~n12492;
  assign n12494 = n12490 & ~n12493;
  assign n12495 = n12488 & n12494;
  assign n12496 = ~n12486 & ~n12495;
  assign n12497 = ~n12479 & ~n12482;
  assign n12498 = ~n12483 & ~n12497;
  assign n12499 = ~n12496 & n12498;
  assign n12500 = ~n12483 & ~n12499;
  assign n12501 = ~n12476 & ~n12479;
  assign n12502 = ~n12480 & ~n12501;
  assign n12503 = ~n12500 & n12502;
  assign n12504 = ~n12480 & ~n12503;
  assign n12505 = ~n12473 & ~n12476;
  assign n12506 = ~n12477 & ~n12505;
  assign n12507 = ~n12504 & n12506;
  assign n12508 = ~n12477 & ~n12507;
  assign n12509 = ~n12470 & ~n12473;
  assign n12510 = ~n12474 & ~n12509;
  assign n12511 = ~n12508 & n12510;
  assign n12512 = ~n12474 & ~n12511;
  assign n12513 = ~n12467 & ~n12470;
  assign n12514 = ~n12471 & ~n12513;
  assign n12515 = ~n12512 & n12514;
  assign n12516 = ~n12471 & ~n12515;
  assign n12517 = ~n12464 & ~n12467;
  assign n12518 = ~n12468 & ~n12517;
  assign n12519 = ~n12516 & n12518;
  assign n12520 = ~n12468 & ~n12519;
  assign n12521 = ~n12461 & ~n12464;
  assign n12522 = ~n12465 & ~n12521;
  assign n12523 = ~n12520 & n12522;
  assign n12524 = ~n12465 & ~n12523;
  assign n12525 = ~n12458 & ~n12461;
  assign n12526 = ~n12462 & ~n12525;
  assign n12527 = ~n12524 & n12526;
  assign n12528 = ~n12462 & ~n12527;
  assign n12529 = ~n12455 & ~n12458;
  assign n12530 = ~n12459 & ~n12529;
  assign n12531 = ~n12528 & n12530;
  assign n12532 = ~n12459 & ~n12531;
  assign n12533 = ~n12452 & ~n12455;
  assign n12534 = ~n12456 & ~n12533;
  assign n12535 = ~n12532 & n12534;
  assign n12536 = ~n12456 & ~n12535;
  assign n12537 = ~n12449 & ~n12452;
  assign n12538 = ~n12453 & ~n12537;
  assign n12539 = ~n12536 & n12538;
  assign n12540 = ~n12453 & ~n12539;
  assign n12541 = ~n12446 & ~n12449;
  assign n12542 = ~n12450 & ~n12541;
  assign n12543 = ~n12540 & n12542;
  assign n12544 = ~n12450 & ~n12543;
  assign n12545 = ~n12443 & ~n12446;
  assign n12546 = ~n12447 & ~n12545;
  assign n12547 = ~n12544 & n12546;
  assign n12548 = ~n12447 & ~n12547;
  assign n12549 = ~n12440 & ~n12443;
  assign n12550 = ~n12444 & ~n12549;
  assign n12551 = ~n12548 & n12550;
  assign n12552 = ~n12444 & ~n12551;
  assign n12553 = ~n12437 & ~n12440;
  assign n12554 = ~n12441 & ~n12553;
  assign n12555 = ~n12552 & n12554;
  assign n12556 = ~n12441 & ~n12555;
  assign n12557 = ~n12434 & ~n12437;
  assign n12558 = ~n12438 & ~n12557;
  assign n12559 = ~n12556 & n12558;
  assign n12560 = ~n12438 & ~n12559;
  assign n12561 = ~n12431 & ~n12434;
  assign n12562 = ~n12435 & ~n12561;
  assign n12563 = ~n12560 & n12562;
  assign n12564 = ~n12435 & ~n12563;
  assign n12565 = ~n12428 & ~n12431;
  assign n12566 = ~n12432 & ~n12565;
  assign n12567 = ~n12564 & n12566;
  assign n12568 = ~n12432 & ~n12567;
  assign n12569 = ~n12425 & ~n12428;
  assign n12570 = ~n12429 & ~n12569;
  assign n12571 = ~n12568 & n12570;
  assign n12572 = ~n12429 & ~n12571;
  assign n12573 = ~n12422 & ~n12425;
  assign n12574 = ~n12426 & ~n12573;
  assign n12575 = ~n12572 & n12574;
  assign n12576 = ~n12426 & ~n12575;
  assign n12577 = ~n12419 & ~n12422;
  assign n12578 = ~n12423 & ~n12577;
  assign n12579 = ~n12576 & n12578;
  assign n12580 = ~n12423 & ~n12579;
  assign n12581 = ~n12416 & ~n12419;
  assign n12582 = ~n12420 & ~n12581;
  assign n12583 = ~n12580 & n12582;
  assign n12584 = ~n12420 & ~n12583;
  assign n12585 = ~n12413 & ~n12416;
  assign n12586 = ~n12417 & ~n12585;
  assign n12587 = ~n12584 & n12586;
  assign n12588 = ~n12417 & ~n12587;
  assign n12589 = ~n12410 & ~n12413;
  assign n12590 = ~n12414 & ~n12589;
  assign n12591 = ~n12588 & n12590;
  assign n12592 = ~n12414 & ~n12591;
  assign n12593 = ~n12407 & ~n12410;
  assign n12594 = ~n12411 & ~n12593;
  assign n12595 = ~n12592 & n12594;
  assign n12596 = ~n12411 & ~n12595;
  assign n12597 = ~n12404 & ~n12407;
  assign n12598 = ~n12408 & ~n12597;
  assign n12599 = ~n12596 & n12598;
  assign n12600 = ~n12408 & ~n12599;
  assign n12601 = ~n12401 & ~n12404;
  assign n12602 = ~n12405 & ~n12601;
  assign n12603 = ~n12600 & n12602;
  assign n12604 = ~n12405 & ~n12603;
  assign n12605 = ~n12398 & ~n12401;
  assign n12606 = ~n12402 & ~n12605;
  assign n12607 = ~n12604 & n12606;
  assign n12608 = ~n12402 & ~n12607;
  assign n12609 = ~n12395 & ~n12398;
  assign n12610 = ~n12399 & ~n12609;
  assign n12611 = ~n12608 & n12610;
  assign n12612 = ~n12399 & ~n12611;
  assign n12613 = ~n12362 & ~n12395;
  assign n12614 = ~n12396 & ~n12613;
  assign n12615 = ~n12612 & n12614;
  assign n12616 = ~n12396 & ~n12615;
  assign n12617 = ~n12362 & ~n12392;
  assign n12618 = ~n12393 & ~n12617;
  assign n12619 = ~n12616 & n12618;
  assign n12620 = ~n12393 & ~n12619;
  assign n12621 = ~n183 & ~n291;
  assign n12622 = ~n486 & n12621;
  assign n12623 = n755 & n1684;
  assign n12624 = n12622 & n12623;
  assign n12625 = n897 & n12624;
  assign n12626 = n3872 & n12625;
  assign n12627 = n12321 & n12626;
  assign n12628 = n3834 & n12627;
  assign n12629 = n12374 & ~n12628;
  assign n12630 = ~n12374 & n12628;
  assign n12631 = ~n12629 & ~n12630;
  assign n12632 = n880 & ~n3897;
  assign n12633 = ~n748 & ~n12632;
  assign n12634 = ~n3883 & ~n12633;
  assign n12635 = n12631 & n12634;
  assign n12636 = ~n12631 & ~n12634;
  assign n12637 = ~n12635 & ~n12636;
  assign n12638 = ~n12376 & ~n12382;
  assign n12639 = ~n12375 & ~n12638;
  assign n12640 = n12637 & ~n12639;
  assign n12641 = ~n12637 & n12639;
  assign n12642 = ~n12640 & ~n12641;
  assign n12643 = ~n12386 & ~n12390;
  assign n12644 = n12642 & ~n12643;
  assign n12645 = ~n12642 & n12643;
  assign n12646 = ~n12644 & ~n12645;
  assign n12647 = n12392 & n12646;
  assign n12648 = ~n12392 & ~n12646;
  assign n12649 = ~n12647 & ~n12648;
  assign n12650 = ~n12620 & n12649;
  assign n12651 = n12620 & ~n12649;
  assign n12652 = ~n12650 & ~n12651;
  assign n12653 = n4420 & n12652;
  assign n12654 = n4600 & n12392;
  assign n12655 = n4615 & n12646;
  assign n12656 = ~n12363 & ~n12654;
  assign n12657 = ~n12655 & n12656;
  assign n12658 = ~n12653 & n12657;
  assign n12659 = pi26  & n12658;
  assign n12660 = ~pi26  & ~n12658;
  assign n12661 = ~n12659 & ~n12660;
  assign n12662 = ~n247 & ~n481;
  assign n12663 = ~n601 & ~n656;
  assign n12664 = n12662 & n12663;
  assign n12665 = n3302 & n3407;
  assign n12666 = n12664 & n12665;
  assign n12667 = ~n480 & ~n902;
  assign n12668 = ~n178 & ~n237;
  assign n12669 = ~n243 & ~n317;
  assign n12670 = ~n332 & ~n599;
  assign n12671 = n12669 & n12670;
  assign n12672 = n360 & n12668;
  assign n12673 = n941 & n1305;
  assign n12674 = n1356 & n1767;
  assign n12675 = n3325 & n12667;
  assign n12676 = n12674 & n12675;
  assign n12677 = n12672 & n12673;
  assign n12678 = n2293 & n12671;
  assign n12679 = n3186 & n12678;
  assign n12680 = n12676 & n12677;
  assign n12681 = n12666 & n12680;
  assign n12682 = n5729 & n12679;
  assign n12683 = n12681 & n12682;
  assign n12684 = n3100 & n12683;
  assign n12685 = n4246 & n12684;
  assign n12686 = ~n171 & ~n188;
  assign n12687 = n1198 & n12686;
  assign n12688 = ~n126 & ~n178;
  assign n12689 = ~n438 & ~n508;
  assign n12690 = n12688 & n12689;
  assign n12691 = n1452 & n4034;
  assign n12692 = ~n135 & ~n174;
  assign n12693 = ~n270 & ~n499;
  assign n12694 = ~n604 & ~n718;
  assign n12695 = n12693 & n12694;
  assign n12696 = n244 & n12692;
  assign n12697 = n12695 & n12696;
  assign n12698 = n4881 & n12691;
  assign n12699 = n12697 & n12698;
  assign n12700 = ~n235 & ~n239;
  assign n12701 = ~n277 & ~n509;
  assign n12702 = n12700 & n12701;
  assign n12703 = n501 & n1151;
  assign n12704 = n2253 & n2473;
  assign n12705 = n12703 & n12704;
  assign n12706 = n429 & n12702;
  assign n12707 = n6984 & n12687;
  assign n12708 = n12690 & n12707;
  assign n12709 = n12705 & n12706;
  assign n12710 = n12708 & n12709;
  assign n12711 = n12699 & n12710;
  assign n12712 = n3322 & n12711;
  assign n12713 = n3933 & n5322;
  assign n12714 = n12712 & n12713;
  assign n12715 = ~n12685 & ~n12714;
  assign n12716 = ~n213 & n1764;
  assign n12717 = ~n329 & ~n379;
  assign n12718 = ~n753 & n12717;
  assign n12719 = ~n367 & ~n381;
  assign n12720 = ~n627 & n12719;
  assign n12721 = n1457 & n12720;
  assign n12722 = ~n199 & ~n352;
  assign n12723 = ~n415 & ~n430;
  assign n12724 = ~n476 & ~n566;
  assign n12725 = n12723 & n12724;
  assign n12726 = n372 & n12722;
  assign n12727 = n2206 & n2548;
  assign n12728 = n2625 & n12727;
  assign n12729 = n12725 & n12726;
  assign n12730 = n12716 & n12718;
  assign n12731 = n12729 & n12730;
  assign n12732 = n12721 & n12728;
  assign n12733 = n12731 & n12732;
  assign n12734 = n3383 & n12733;
  assign n12735 = n2380 & n12734;
  assign n12736 = n3716 & n12735;
  assign n12737 = ~n163 & ~n339;
  assign n12738 = ~n362 & ~n409;
  assign n12739 = ~n944 & n12738;
  assign n12740 = n1272 & n12737;
  assign n12741 = n1384 & n1863;
  assign n12742 = n4264 & n12741;
  assign n12743 = n12739 & n12740;
  assign n12744 = n4736 & n12743;
  assign n12745 = n12742 & n12744;
  assign n12746 = ~n337 & ~n511;
  assign n12747 = n705 & n12746;
  assign n12748 = n1035 & n1246;
  assign n12749 = n1428 & n1476;
  assign n12750 = n2007 & n12749;
  assign n12751 = n12747 & n12748;
  assign n12752 = n1279 & n2794;
  assign n12753 = n6969 & n12752;
  assign n12754 = n12750 & n12751;
  assign n12755 = n6928 & n12754;
  assign n12756 = n2389 & n12753;
  assign n12757 = n12755 & n12756;
  assign n12758 = n12745 & n12757;
  assign n12759 = n3757 & n12758;
  assign n12760 = n12736 & n12759;
  assign n12761 = ~n361 & n1136;
  assign n12762 = n3814 & n12761;
  assign n12763 = n12760 & n12762;
  assign n12764 = ~n12629 & ~n12635;
  assign n12765 = n934 & n1169;
  assign n12766 = ~n177 & ~n304;
  assign n12767 = ~n432 & n12766;
  assign n12768 = n3619 & n12767;
  assign n12769 = n12765 & n12768;
  assign n12770 = n3848 & n12769;
  assign n12771 = n3676 & n12770;
  assign n12772 = n12374 & n12771;
  assign n12773 = ~n12374 & ~n12771;
  assign n12774 = ~n12772 & ~n12773;
  assign n12775 = ~n12764 & ~n12774;
  assign n12776 = ~n12764 & n12774;
  assign n12777 = n12764 & ~n12774;
  assign n12778 = ~n12776 & ~n12777;
  assign n12779 = ~n12640 & ~n12644;
  assign n12780 = ~n12778 & ~n12779;
  assign n12781 = ~n12775 & ~n12780;
  assign n12782 = ~n12763 & n12772;
  assign n12783 = n12763 & ~n12772;
  assign n12784 = ~n12782 & ~n12783;
  assign n12785 = ~n12781 & n12784;
  assign n12786 = ~n12763 & n12785;
  assign n12787 = n5974 & n5981;
  assign n12788 = ~n12786 & ~n12787;
  assign n12789 = pi17  & ~n12788;
  assign n12790 = ~pi17  & n12788;
  assign n12791 = ~n12789 & ~n12790;
  assign n12792 = n12685 & n12714;
  assign n12793 = ~n12715 & ~n12792;
  assign n12794 = n12791 & n12793;
  assign n12795 = ~n12715 & ~n12794;
  assign n12796 = ~n183 & ~n536;
  assign n12797 = ~n1404 & n12796;
  assign n12798 = n2889 & n12317;
  assign n12799 = n12797 & n12798;
  assign n12800 = ~n307 & ~n509;
  assign n12801 = n2320 & n12800;
  assign n12802 = n2608 & n2783;
  assign n12803 = n4709 & n12802;
  assign n12804 = n6844 & n12801;
  assign n12805 = n12803 & n12804;
  assign n12806 = ~n277 & n807;
  assign n12807 = n2962 & n12806;
  assign n12808 = n418 & n12807;
  assign n12809 = n5486 & n12799;
  assign n12810 = n12808 & n12809;
  assign n12811 = n12805 & n12810;
  assign n12812 = ~n170 & ~n194;
  assign n12813 = ~n216 & ~n376;
  assign n12814 = ~n561 & ~n625;
  assign n12815 = ~n724 & ~n838;
  assign n12816 = n12814 & n12815;
  assign n12817 = n12812 & n12813;
  assign n12818 = n12816 & n12817;
  assign n12819 = ~n374 & ~n446;
  assign n12820 = ~n894 & n12819;
  assign n12821 = n298 & ~n646;
  assign n12822 = n1471 & n12821;
  assign n12823 = n12820 & n12822;
  assign n12824 = ~n430 & ~n458;
  assign n12825 = ~n689 & ~n902;
  assign n12826 = n12824 & n12825;
  assign n12827 = n160 & n1350;
  assign n12828 = n1651 & n2197;
  assign n12829 = n3204 & n12828;
  assign n12830 = n12826 & n12827;
  assign n12831 = n4829 & n12830;
  assign n12832 = n12818 & n12829;
  assign n12833 = n12831 & n12832;
  assign n12834 = n12699 & n12823;
  assign n12835 = n12833 & n12834;
  assign n12836 = n12811 & n12835;
  assign n12837 = n3341 & n12836;
  assign n12838 = ~n12795 & n12837;
  assign n12839 = n12795 & ~n12837;
  assign n12840 = ~n12838 & ~n12839;
  assign n12841 = n3692 & n12413;
  assign n12842 = n12588 & ~n12590;
  assign n12843 = ~n12591 & ~n12842;
  assign n12844 = n880 & n12843;
  assign n12845 = n748 & n12416;
  assign n12846 = n3694 & n12410;
  assign n12847 = ~n12841 & ~n12845;
  assign n12848 = ~n12846 & n12847;
  assign n12849 = ~n12844 & n12848;
  assign n12850 = n12840 & ~n12849;
  assign n12851 = ~n12838 & ~n12850;
  assign n12852 = ~n120 & ~n190;
  assign n12853 = ~n302 & ~n332;
  assign n12854 = ~n477 & n12853;
  assign n12855 = n2711 & n12854;
  assign n12856 = ~n111 & ~n299;
  assign n12857 = ~n377 & ~n499;
  assign n12858 = ~n535 & ~n603;
  assign n12859 = ~n703 & ~n893;
  assign n12860 = n12858 & n12859;
  assign n12861 = n12856 & n12857;
  assign n12862 = n1087 & n1812;
  assign n12863 = n2037 & n2625;
  assign n12864 = n12862 & n12863;
  assign n12865 = n12860 & n12861;
  assign n12866 = n1269 & n3445;
  assign n12867 = n12865 & n12866;
  assign n12868 = n12864 & n12867;
  assign n12869 = n2746 & n12868;
  assign n12870 = ~n307 & ~n523;
  assign n12871 = ~n646 & n12870;
  assign n12872 = n146 & n530;
  assign n12873 = n716 & n940;
  assign n12874 = n1284 & n2208;
  assign n12875 = n3644 & n12852;
  assign n12876 = n12874 & n12875;
  assign n12877 = n12872 & n12873;
  assign n12878 = n4889 & n12871;
  assign n12879 = n12877 & n12878;
  assign n12880 = n2102 & n12876;
  assign n12881 = n12855 & n12880;
  assign n12882 = n12879 & n12881;
  assign n12883 = n2756 & n12882;
  assign n12884 = n5677 & n12869;
  assign n12885 = n12883 & n12884;
  assign n12886 = n12837 & ~n12885;
  assign n12887 = ~n12837 & n12885;
  assign n12888 = ~n12886 & ~n12887;
  assign n12889 = n748 & n12413;
  assign n12890 = n12592 & ~n12594;
  assign n12891 = ~n12595 & ~n12890;
  assign n12892 = n880 & n12891;
  assign n12893 = n3692 & n12410;
  assign n12894 = n3694 & n12407;
  assign n12895 = ~n12889 & ~n12893;
  assign n12896 = ~n12894 & n12895;
  assign n12897 = ~n12892 & n12896;
  assign n12898 = n12888 & ~n12897;
  assign n12899 = ~n12888 & n12897;
  assign n12900 = ~n12898 & ~n12899;
  assign n12901 = ~n12851 & n12900;
  assign n12902 = n12851 & ~n12900;
  assign n12903 = ~n12901 & ~n12902;
  assign n12904 = ~n12791 & ~n12793;
  assign n12905 = ~n12794 & ~n12904;
  assign n12906 = n748 & n12419;
  assign n12907 = n12584 & ~n12586;
  assign n12908 = ~n12587 & ~n12907;
  assign n12909 = n880 & n12908;
  assign n12910 = n3692 & n12416;
  assign n12911 = n3694 & n12413;
  assign n12912 = ~n12906 & ~n12910;
  assign n12913 = ~n12911 & n12912;
  assign n12914 = ~n12909 & n12913;
  assign n12915 = n12905 & ~n12914;
  assign n12916 = ~n317 & ~n359;
  assign n12917 = ~n536 & ~n594;
  assign n12918 = ~n792 & n12917;
  assign n12919 = n413 & n12916;
  assign n12920 = n444 & n504;
  assign n12921 = n1457 & n3219;
  assign n12922 = n12920 & n12921;
  assign n12923 = n12918 & n12919;
  assign n12924 = n12922 & n12923;
  assign n12925 = ~n416 & ~n435;
  assign n12926 = ~n333 & ~n510;
  assign n12927 = ~n592 & ~n596;
  assign n12928 = n12926 & n12927;
  assign n12929 = n960 & n12928;
  assign n12930 = ~n338 & ~n534;
  assign n12931 = ~n238 & ~n356;
  assign n12932 = ~n846 & ~n989;
  assign n12933 = n12931 & n12932;
  assign n12934 = n528 & n3458;
  assign n12935 = n4269 & n5300;
  assign n12936 = n12930 & n12935;
  assign n12937 = n12933 & n12934;
  assign n12938 = n12936 & n12937;
  assign n12939 = n6414 & n12929;
  assign n12940 = n12938 & n12939;
  assign n12941 = n4856 & n12940;
  assign n12942 = ~n136 & n311;
  assign n12943 = n12941 & n12942;
  assign n12944 = n2473 & n3224;
  assign n12945 = ~n188 & ~n211;
  assign n12946 = ~n215 & ~n432;
  assign n12947 = ~n518 & n12946;
  assign n12948 = n1133 & n12945;
  assign n12949 = n2037 & n12925;
  assign n12950 = n12948 & n12949;
  assign n12951 = n2161 & n12947;
  assign n12952 = n2724 & n12944;
  assign n12953 = n12951 & n12952;
  assign n12954 = n289 & n12950;
  assign n12955 = n12953 & n12954;
  assign n12956 = n12924 & n12955;
  assign n12957 = n3396 & n12956;
  assign n12958 = n12943 & n12957;
  assign n12959 = n12685 & ~n12958;
  assign n12960 = ~n277 & ~n318;
  assign n12961 = n5550 & n12960;
  assign n12962 = ~n195 & ~n333;
  assign n12963 = ~n427 & ~n486;
  assign n12964 = ~n123 & ~n646;
  assign n12965 = n505 & n12964;
  assign n12966 = n811 & n935;
  assign n12967 = n12962 & n12963;
  assign n12968 = n12966 & n12967;
  assign n12969 = n5719 & n12965;
  assign n12970 = n12968 & n12969;
  assign n12971 = n2051 & n12970;
  assign n12972 = n3470 & n12971;
  assign n12973 = n1263 & n12972;
  assign n12974 = n12961 & n12973;
  assign n12975 = ~n136 & ~n190;
  assign n12976 = ~n334 & ~n751;
  assign n12977 = n12975 & n12976;
  assign n12978 = n528 & n1575;
  assign n12979 = n12977 & n12978;
  assign n12980 = n217 & n1754;
  assign n12981 = ~n145 & ~n238;
  assign n12982 = ~n278 & ~n365;
  assign n12983 = ~n535 & n12982;
  assign n12984 = n2350 & n12981;
  assign n12985 = n12983 & n12984;
  assign n12986 = n4831 & n4955;
  assign n12987 = n12980 & n12986;
  assign n12988 = n1586 & n12985;
  assign n12989 = n4162 & n12979;
  assign n12990 = n12988 & n12989;
  assign n12991 = n2635 & n12987;
  assign n12992 = n12990 & n12991;
  assign n12993 = n2607 & n12992;
  assign n12994 = n6842 & n12993;
  assign n12995 = ~n12974 & ~n12994;
  assign n12996 = n6622 & n6629;
  assign n12997 = ~n12786 & ~n12996;
  assign n12998 = pi14  & ~n12997;
  assign n12999 = ~pi14  & n12997;
  assign n13000 = ~n12998 & ~n12999;
  assign n13001 = n12974 & n12994;
  assign n13002 = ~n12995 & ~n13001;
  assign n13003 = n13000 & n13002;
  assign n13004 = ~n12995 & ~n13003;
  assign n13005 = n12958 & ~n13004;
  assign n13006 = ~n12958 & n13004;
  assign n13007 = ~n13005 & ~n13006;
  assign n13008 = n3692 & n12422;
  assign n13009 = n12576 & ~n12578;
  assign n13010 = ~n12579 & ~n13009;
  assign n13011 = n880 & n13010;
  assign n13012 = n748 & n12425;
  assign n13013 = n3694 & n12419;
  assign n13014 = ~n13008 & ~n13012;
  assign n13015 = ~n13013 & n13014;
  assign n13016 = ~n13011 & n13015;
  assign n13017 = n13007 & ~n13016;
  assign n13018 = ~n13005 & ~n13017;
  assign n13019 = ~n12685 & n12958;
  assign n13020 = ~n12959 & ~n13019;
  assign n13021 = ~n13018 & n13020;
  assign n13022 = ~n12959 & ~n13021;
  assign n13023 = n12905 & n12914;
  assign n13024 = ~n12905 & ~n12914;
  assign n13025 = ~n13023 & ~n13024;
  assign n13026 = ~n13022 & ~n13025;
  assign n13027 = ~n12915 & ~n13026;
  assign n13028 = ~n12840 & n12849;
  assign n13029 = ~n12850 & ~n13028;
  assign n13030 = ~n13027 & n13029;
  assign n13031 = n13027 & ~n13029;
  assign n13032 = ~n13030 & ~n13031;
  assign n13033 = n3810 & n12407;
  assign n13034 = n12600 & ~n12602;
  assign n13035 = ~n12603 & ~n13034;
  assign n13036 = n3886 & n13035;
  assign n13037 = n3884 & n12404;
  assign n13038 = n4380 & n12401;
  assign n13039 = ~n13033 & ~n13037;
  assign n13040 = ~n13038 & n13039;
  assign n13041 = ~n13036 & n13040;
  assign n13042 = pi29  & n13041;
  assign n13043 = ~pi29  & ~n13041;
  assign n13044 = ~n13042 & ~n13043;
  assign n13045 = n13032 & ~n13044;
  assign n13046 = ~n13030 & ~n13045;
  assign n13047 = n12903 & ~n13046;
  assign n13048 = ~n12901 & ~n13047;
  assign n13049 = ~n12886 & ~n12898;
  assign n13050 = n5232 & n5239;
  assign n13051 = ~n12786 & ~n13050;
  assign n13052 = pi20  & ~n13051;
  assign n13053 = ~pi20  & n13051;
  assign n13054 = ~n13052 & ~n13053;
  assign n13055 = n1453 & n2208;
  assign n13056 = ~n139 & ~n238;
  assign n13057 = ~n531 & n13056;
  assign n13058 = n1474 & n1489;
  assign n13059 = n2682 & n5474;
  assign n13060 = n12925 & n13059;
  assign n13061 = n13057 & n13058;
  assign n13062 = n13055 & n13061;
  assign n13063 = n1083 & n13060;
  assign n13064 = n3312 & n13063;
  assign n13065 = n2191 & n13062;
  assign n13066 = n13064 & n13065;
  assign n13067 = ~n270 & ~n411;
  assign n13068 = ~n439 & ~n445;
  assign n13069 = ~n721 & n13068;
  assign n13070 = n628 & n13067;
  assign n13071 = n704 & n1578;
  assign n13072 = n1697 & n1858;
  assign n13073 = n3997 & n13072;
  assign n13074 = n13070 & n13071;
  assign n13075 = n4313 & n13069;
  assign n13076 = n13074 & n13075;
  assign n13077 = n13073 & n13076;
  assign n13078 = n1922 & n3406;
  assign n13079 = n13077 & n13078;
  assign n13080 = n13066 & n13079;
  assign n13081 = n2560 & n13080;
  assign n13082 = ~n12837 & ~n13081;
  assign n13083 = n12837 & n13081;
  assign n13084 = ~n13082 & ~n13083;
  assign n13085 = n13054 & n13084;
  assign n13086 = ~n13054 & ~n13084;
  assign n13087 = ~n13085 & ~n13086;
  assign n13088 = ~n13049 & n13087;
  assign n13089 = n13049 & ~n13087;
  assign n13090 = ~n13088 & ~n13089;
  assign n13091 = n748 & n12410;
  assign n13092 = n12596 & ~n12598;
  assign n13093 = ~n12599 & ~n13092;
  assign n13094 = n880 & n13093;
  assign n13095 = n3692 & n12407;
  assign n13096 = n3694 & n12404;
  assign n13097 = ~n13091 & ~n13095;
  assign n13098 = ~n13096 & n13097;
  assign n13099 = ~n13094 & n13098;
  assign n13100 = n13090 & ~n13099;
  assign n13101 = ~n13090 & n13099;
  assign n13102 = ~n13100 & ~n13101;
  assign n13103 = ~n13048 & n13102;
  assign n13104 = n13048 & ~n13102;
  assign n13105 = ~n13103 & ~n13104;
  assign n13106 = n3810 & n12401;
  assign n13107 = n12608 & ~n12610;
  assign n13108 = ~n12611 & ~n13107;
  assign n13109 = n3886 & n13108;
  assign n13110 = n3884 & n12398;
  assign n13111 = n4380 & n12395;
  assign n13112 = ~n13106 & ~n13110;
  assign n13113 = ~n13111 & n13112;
  assign n13114 = ~n13109 & n13113;
  assign n13115 = pi29  & n13114;
  assign n13116 = ~pi29  & ~n13114;
  assign n13117 = ~n13115 & ~n13116;
  assign n13118 = n13105 & ~n13117;
  assign n13119 = ~n13105 & n13117;
  assign n13120 = ~n13118 & ~n13119;
  assign n13121 = n12661 & n13120;
  assign n13122 = ~n12661 & ~n13120;
  assign n13123 = ~n13121 & ~n13122;
  assign n13124 = ~n12903 & n13046;
  assign n13125 = ~n13047 & ~n13124;
  assign n13126 = n3810 & n12404;
  assign n13127 = n12604 & ~n12606;
  assign n13128 = ~n12607 & ~n13127;
  assign n13129 = n3886 & n13128;
  assign n13130 = n3884 & n12401;
  assign n13131 = n4380 & n12398;
  assign n13132 = ~n13126 & ~n13130;
  assign n13133 = ~n13131 & n13132;
  assign n13134 = ~n13129 & n13133;
  assign n13135 = pi29  & n13134;
  assign n13136 = ~pi29  & ~n13134;
  assign n13137 = ~n13135 & ~n13136;
  assign n13138 = n13125 & ~n13137;
  assign n13139 = n13125 & n13137;
  assign n13140 = ~n13125 & ~n13137;
  assign n13141 = ~n13139 & ~n13140;
  assign n13142 = n86 & n12395;
  assign n13143 = n12616 & ~n12618;
  assign n13144 = ~n12619 & ~n13143;
  assign n13145 = n4420 & n13144;
  assign n13146 = n4600 & n12362;
  assign n13147 = n4615 & n12392;
  assign n13148 = ~n13142 & ~n13146;
  assign n13149 = ~n13147 & n13148;
  assign n13150 = ~n13145 & n13149;
  assign n13151 = pi26  & n13150;
  assign n13152 = ~pi26  & ~n13150;
  assign n13153 = ~n13151 & ~n13152;
  assign n13154 = ~n13141 & ~n13153;
  assign n13155 = ~n13138 & ~n13154;
  assign n13156 = ~n13123 & ~n13155;
  assign n13157 = n13123 & n13155;
  assign n13158 = ~n13156 & ~n13157;
  assign n13159 = n12763 & n12772;
  assign n13160 = ~n12785 & n13159;
  assign n13161 = ~n12786 & ~n13160;
  assign n13162 = n5130 & n13161;
  assign n13163 = n12778 & n12779;
  assign n13164 = ~n12780 & ~n13163;
  assign n13165 = n12781 & ~n12784;
  assign n13166 = ~n12785 & ~n13165;
  assign n13167 = n13164 & n13166;
  assign n13168 = n12646 & n13164;
  assign n13169 = ~n12647 & ~n12650;
  assign n13170 = ~n12646 & ~n13164;
  assign n13171 = ~n13168 & ~n13170;
  assign n13172 = ~n13169 & n13171;
  assign n13173 = ~n13168 & ~n13172;
  assign n13174 = ~n13164 & ~n13166;
  assign n13175 = ~n13167 & ~n13174;
  assign n13176 = ~n13173 & n13175;
  assign n13177 = ~n13167 & ~n13176;
  assign n13178 = ~n13161 & ~n13166;
  assign n13179 = ~n13160 & n13166;
  assign n13180 = ~n13178 & ~n13179;
  assign n13181 = ~n13177 & n13180;
  assign n13182 = n13177 & ~n13180;
  assign n13183 = ~n13181 & ~n13182;
  assign n13184 = n5045 & n13183;
  assign n13185 = n5109 & n13166;
  assign n13186 = n5044 & n13164;
  assign n13187 = ~n13185 & ~n13186;
  assign n13188 = ~n13162 & n13187;
  assign n13189 = ~n13184 & n13188;
  assign n13190 = pi23  & n13189;
  assign n13191 = ~pi23  & ~n13189;
  assign n13192 = ~n13190 & ~n13191;
  assign n13193 = n13141 & n13153;
  assign n13194 = ~n13154 & ~n13193;
  assign n13195 = ~n13032 & n13044;
  assign n13196 = ~n13045 & ~n13195;
  assign n13197 = n13018 & ~n13020;
  assign n13198 = ~n13021 & ~n13197;
  assign n13199 = n748 & n12422;
  assign n13200 = n12580 & ~n12582;
  assign n13201 = ~n12583 & ~n13200;
  assign n13202 = n880 & n13201;
  assign n13203 = n3692 & n12419;
  assign n13204 = n3694 & n12416;
  assign n13205 = ~n13199 & ~n13203;
  assign n13206 = ~n13204 & n13205;
  assign n13207 = ~n13202 & n13206;
  assign n13208 = n13198 & ~n13207;
  assign n13209 = n13198 & n13207;
  assign n13210 = ~n13198 & ~n13207;
  assign n13211 = ~n13209 & ~n13210;
  assign n13212 = n3810 & n12413;
  assign n13213 = n3886 & n12891;
  assign n13214 = n3884 & n12410;
  assign n13215 = n4380 & n12407;
  assign n13216 = ~n13212 & ~n13214;
  assign n13217 = ~n13215 & n13216;
  assign n13218 = ~n13213 & n13217;
  assign n13219 = pi29  & n13218;
  assign n13220 = ~pi29  & ~n13218;
  assign n13221 = ~n13219 & ~n13220;
  assign n13222 = ~n13211 & ~n13221;
  assign n13223 = ~n13208 & ~n13222;
  assign n13224 = n13022 & ~n13025;
  assign n13225 = ~n13022 & n13025;
  assign n13226 = ~n13224 & ~n13225;
  assign n13227 = ~n13223 & ~n13226;
  assign n13228 = n3810 & n12410;
  assign n13229 = n3886 & n13093;
  assign n13230 = n3884 & n12407;
  assign n13231 = n4380 & n12404;
  assign n13232 = ~n13228 & ~n13230;
  assign n13233 = ~n13231 & n13232;
  assign n13234 = ~n13229 & n13233;
  assign n13235 = pi29  & n13234;
  assign n13236 = ~pi29  & ~n13234;
  assign n13237 = ~n13235 & ~n13236;
  assign n13238 = n13223 & n13226;
  assign n13239 = ~n13237 & ~n13238;
  assign n13240 = ~n13227 & ~n13239;
  assign n13241 = n13196 & ~n13240;
  assign n13242 = ~n13196 & n13240;
  assign n13243 = n86 & n12398;
  assign n13244 = n12612 & ~n12614;
  assign n13245 = ~n12615 & ~n13244;
  assign n13246 = n4420 & n13245;
  assign n13247 = n4600 & n12395;
  assign n13248 = n4615 & n12362;
  assign n13249 = ~n13243 & ~n13247;
  assign n13250 = ~n13248 & n13249;
  assign n13251 = ~n13246 & n13250;
  assign n13252 = pi26  & n13251;
  assign n13253 = ~pi26  & ~n13251;
  assign n13254 = ~n13252 & ~n13253;
  assign n13255 = ~n13242 & ~n13254;
  assign n13256 = ~n13241 & ~n13255;
  assign n13257 = n13194 & ~n13256;
  assign n13258 = ~n13194 & n13256;
  assign n13259 = n5044 & n12646;
  assign n13260 = n13173 & ~n13175;
  assign n13261 = ~n13176 & ~n13260;
  assign n13262 = n5045 & n13261;
  assign n13263 = n5109 & n13164;
  assign n13264 = n5130 & n13166;
  assign n13265 = ~n13259 & ~n13263;
  assign n13266 = ~n13264 & n13265;
  assign n13267 = ~n13262 & n13266;
  assign n13268 = pi23  & n13267;
  assign n13269 = ~pi23  & ~n13267;
  assign n13270 = ~n13268 & ~n13269;
  assign n13271 = ~n13258 & ~n13270;
  assign n13272 = ~n13257 & ~n13271;
  assign n13273 = n13192 & ~n13272;
  assign n13274 = ~n13192 & n13272;
  assign n13275 = ~n13273 & ~n13274;
  assign n13276 = n13158 & ~n13275;
  assign n13277 = ~n13158 & n13275;
  assign n13278 = ~n13276 & ~n13277;
  assign n13279 = n13160 & n13181;
  assign n13280 = ~n13161 & ~n13279;
  assign n13281 = n5241 & ~n13280;
  assign n13282 = n5240 & ~n13160;
  assign n13283 = ~n5853 & ~n5866;
  assign n13284 = ~n13282 & n13283;
  assign n13285 = ~n12786 & ~n13284;
  assign n13286 = ~n13281 & ~n13285;
  assign n13287 = pi20  & n13286;
  assign n13288 = ~pi20  & ~n13286;
  assign n13289 = ~n13287 & ~n13288;
  assign n13290 = n86 & n12401;
  assign n13291 = n4420 & n13108;
  assign n13292 = n4600 & n12398;
  assign n13293 = n4615 & n12395;
  assign n13294 = ~n13290 & ~n13292;
  assign n13295 = ~n13293 & n13294;
  assign n13296 = ~n13291 & n13295;
  assign n13297 = pi26  & n13296;
  assign n13298 = ~pi26  & ~n13296;
  assign n13299 = ~n13297 & ~n13298;
  assign n13300 = ~n13227 & ~n13238;
  assign n13301 = n13237 & ~n13300;
  assign n13302 = ~n13237 & n13300;
  assign n13303 = ~n13301 & ~n13302;
  assign n13304 = ~n13299 & n13303;
  assign n13305 = n13299 & n13303;
  assign n13306 = ~n13299 & ~n13303;
  assign n13307 = ~n13305 & ~n13306;
  assign n13308 = ~n13007 & n13016;
  assign n13309 = ~n13017 & ~n13308;
  assign n13310 = ~n561 & ~n894;
  assign n13311 = n848 & n13310;
  assign n13312 = n939 & n1914;
  assign n13313 = n2608 & n6196;
  assign n13314 = n13312 & n13313;
  assign n13315 = n4268 & n13311;
  assign n13316 = n13314 & n13315;
  assign n13317 = n142 & n4687;
  assign n13318 = n375 & n1642;
  assign n13319 = ~n130 & ~n328;
  assign n13320 = ~n503 & ~n534;
  assign n13321 = ~n603 & ~n838;
  assign n13322 = n13320 & n13321;
  assign n13323 = n13319 & n13322;
  assign n13324 = ~n529 & ~n698;
  assign n13325 = n1321 & n13324;
  assign n13326 = n1752 & n1890;
  assign n13327 = n3726 & n13326;
  assign n13328 = n306 & n13325;
  assign n13329 = n854 & n1265;
  assign n13330 = n2021 & n13318;
  assign n13331 = n13329 & n13330;
  assign n13332 = n13327 & n13328;
  assign n13333 = n13323 & n13332;
  assign n13334 = n13331 & n13333;
  assign n13335 = ~n237 & ~n250;
  assign n13336 = ~n253 & ~n277;
  assign n13337 = ~n314 & ~n319;
  assign n13338 = ~n365 & ~n378;
  assign n13339 = n13337 & n13338;
  assign n13340 = n13335 & n13336;
  assign n13341 = n749 & n1578;
  assign n13342 = n13340 & n13341;
  assign n13343 = n1541 & n13339;
  assign n13344 = n13317 & n13343;
  assign n13345 = n3059 & n13342;
  assign n13346 = n13344 & n13345;
  assign n13347 = n3994 & n13316;
  assign n13348 = n13346 & n13347;
  assign n13349 = n2867 & n13348;
  assign n13350 = n13334 & n13349;
  assign n13351 = n12974 & ~n13350;
  assign n13352 = ~n12974 & n13350;
  assign n13353 = ~n13351 & ~n13352;
  assign n13354 = n748 & n12431;
  assign n13355 = n12568 & ~n12570;
  assign n13356 = ~n12571 & ~n13355;
  assign n13357 = n880 & n13356;
  assign n13358 = n3692 & n12428;
  assign n13359 = n3694 & n12425;
  assign n13360 = ~n13354 & ~n13358;
  assign n13361 = ~n13359 & n13360;
  assign n13362 = ~n13357 & n13361;
  assign n13363 = n13353 & ~n13362;
  assign n13364 = ~n13351 & ~n13363;
  assign n13365 = ~n13000 & ~n13002;
  assign n13366 = ~n13003 & ~n13365;
  assign n13367 = ~n13364 & n13366;
  assign n13368 = n13364 & ~n13366;
  assign n13369 = n748 & n12428;
  assign n13370 = n12572 & ~n12574;
  assign n13371 = ~n12575 & ~n13370;
  assign n13372 = n880 & n13371;
  assign n13373 = n3692 & n12425;
  assign n13374 = n3694 & n12422;
  assign n13375 = ~n13369 & ~n13373;
  assign n13376 = ~n13374 & n13375;
  assign n13377 = ~n13372 & n13376;
  assign n13378 = ~n13368 & ~n13377;
  assign n13379 = ~n13367 & ~n13378;
  assign n13380 = n13309 & ~n13379;
  assign n13381 = ~n13309 & n13379;
  assign n13382 = ~n13380 & ~n13381;
  assign n13383 = n3810 & n12416;
  assign n13384 = n3886 & n12843;
  assign n13385 = n3884 & n12413;
  assign n13386 = n4380 & n12410;
  assign n13387 = ~n13383 & ~n13385;
  assign n13388 = ~n13386 & n13387;
  assign n13389 = ~n13384 & n13388;
  assign n13390 = pi29  & n13389;
  assign n13391 = ~pi29  & ~n13389;
  assign n13392 = ~n13390 & ~n13391;
  assign n13393 = n13382 & ~n13392;
  assign n13394 = ~n13380 & ~n13393;
  assign n13395 = n13211 & n13221;
  assign n13396 = ~n13222 & ~n13395;
  assign n13397 = ~n13394 & n13396;
  assign n13398 = n13394 & ~n13396;
  assign n13399 = n86 & n12404;
  assign n13400 = n4420 & n13128;
  assign n13401 = n4600 & n12401;
  assign n13402 = n4615 & n12398;
  assign n13403 = ~n13399 & ~n13401;
  assign n13404 = ~n13402 & n13403;
  assign n13405 = ~n13400 & n13404;
  assign n13406 = pi26  & n13405;
  assign n13407 = ~pi26  & ~n13405;
  assign n13408 = ~n13406 & ~n13407;
  assign n13409 = ~n13398 & ~n13408;
  assign n13410 = ~n13397 & ~n13409;
  assign n13411 = ~n13307 & ~n13410;
  assign n13412 = ~n13304 & ~n13411;
  assign n13413 = ~n13241 & ~n13242;
  assign n13414 = ~n13254 & n13413;
  assign n13415 = n13254 & ~n13413;
  assign n13416 = ~n13414 & ~n13415;
  assign n13417 = ~n13412 & n13416;
  assign n13418 = n13412 & ~n13416;
  assign n13419 = n5044 & n12392;
  assign n13420 = n13169 & ~n13171;
  assign n13421 = ~n13172 & ~n13420;
  assign n13422 = n5045 & n13421;
  assign n13423 = n5109 & n12646;
  assign n13424 = n5130 & n13164;
  assign n13425 = ~n13419 & ~n13423;
  assign n13426 = ~n13424 & n13425;
  assign n13427 = ~n13422 & n13426;
  assign n13428 = pi23  & n13427;
  assign n13429 = ~pi23  & ~n13427;
  assign n13430 = ~n13428 & ~n13429;
  assign n13431 = ~n13418 & ~n13430;
  assign n13432 = ~n13417 & ~n13431;
  assign n13433 = ~n13289 & ~n13432;
  assign n13434 = n13289 & n13432;
  assign n13435 = ~n13257 & ~n13258;
  assign n13436 = ~n13270 & n13435;
  assign n13437 = n13270 & ~n13435;
  assign n13438 = ~n13436 & ~n13437;
  assign n13439 = ~n13434 & n13438;
  assign n13440 = ~n13433 & ~n13439;
  assign n13441 = n13278 & ~n13440;
  assign n13442 = ~n13433 & ~n13434;
  assign n13443 = n13438 & n13442;
  assign n13444 = ~n13438 & ~n13442;
  assign n13445 = ~n13443 & ~n13444;
  assign n13446 = n13307 & n13410;
  assign n13447 = ~n13411 & ~n13446;
  assign n13448 = n5044 & n12362;
  assign n13449 = n5045 & n12652;
  assign n13450 = n5109 & n12392;
  assign n13451 = n5130 & n12646;
  assign n13452 = ~n13448 & ~n13450;
  assign n13453 = ~n13451 & n13452;
  assign n13454 = ~n13449 & n13453;
  assign n13455 = pi23  & n13454;
  assign n13456 = ~pi23  & ~n13454;
  assign n13457 = ~n13455 & ~n13456;
  assign n13458 = n13447 & ~n13457;
  assign n13459 = n13447 & n13457;
  assign n13460 = ~n13447 & ~n13457;
  assign n13461 = ~n13459 & ~n13460;
  assign n13462 = ~n13397 & ~n13398;
  assign n13463 = ~n13408 & n13462;
  assign n13464 = n13408 & ~n13462;
  assign n13465 = ~n13463 & ~n13464;
  assign n13466 = n3810 & n12419;
  assign n13467 = n3886 & n12908;
  assign n13468 = n3884 & n12416;
  assign n13469 = n4380 & n12413;
  assign n13470 = ~n13466 & ~n13468;
  assign n13471 = ~n13469 & n13470;
  assign n13472 = ~n13467 & n13471;
  assign n13473 = pi29  & n13472;
  assign n13474 = ~pi29  & ~n13472;
  assign n13475 = ~n13473 & ~n13474;
  assign n13476 = ~n13367 & ~n13368;
  assign n13477 = ~n13377 & n13476;
  assign n13478 = n13377 & ~n13476;
  assign n13479 = ~n13477 & ~n13478;
  assign n13480 = ~n13475 & n13479;
  assign n13481 = ~n200 & ~n365;
  assign n13482 = ~n520 & ~n601;
  assign n13483 = ~n685 & ~n808;
  assign n13484 = ~n1002 & ~n1051;
  assign n13485 = n13483 & n13484;
  assign n13486 = n13481 & n13482;
  assign n13487 = n901 & n2460;
  assign n13488 = n13486 & n13487;
  assign n13489 = n2194 & n13485;
  assign n13490 = n13488 & n13489;
  assign n13491 = ~n529 & ~n566;
  assign n13492 = ~n568 & n13491;
  assign n13493 = n1644 & n5523;
  assign n13494 = n13492 & n13493;
  assign n13495 = ~n148 & ~n239;
  assign n13496 = ~n245 & ~n302;
  assign n13497 = ~n356 & ~n944;
  assign n13498 = n13496 & n13497;
  assign n13499 = n797 & n13495;
  assign n13500 = n1321 & n1428;
  assign n13501 = n3325 & n4828;
  assign n13502 = n13500 & n13501;
  assign n13503 = n13498 & n13499;
  assign n13504 = n2781 & n3910;
  assign n13505 = n13503 & n13504;
  assign n13506 = n4717 & n13502;
  assign n13507 = n13494 & n13506;
  assign n13508 = n13490 & n13505;
  assign n13509 = n13507 & n13508;
  assign n13510 = n475 & n13509;
  assign n13511 = n6462 & n13510;
  assign n13512 = ~n252 & ~n839;
  assign n13513 = ~n663 & ~n703;
  assign n13514 = ~n195 & n3008;
  assign n13515 = n13513 & n13514;
  assign n13516 = n2008 & n13515;
  assign n13517 = ~n309 & ~n508;
  assign n13518 = n410 & n13517;
  assign n13519 = n1859 & n2052;
  assign n13520 = n13512 & n13519;
  assign n13521 = n812 & n13518;
  assign n13522 = n1239 & n3047;
  assign n13523 = n4829 & n13522;
  assign n13524 = n13520 & n13521;
  assign n13525 = n13523 & n13524;
  assign n13526 = n13516 & n13525;
  assign n13527 = n1469 & n2034;
  assign n13528 = n6168 & n13527;
  assign n13529 = n1045 & n13526;
  assign n13530 = n13528 & n13529;
  assign n13531 = ~n13511 & ~n13530;
  assign n13532 = n7422 & n7429;
  assign n13533 = ~n12786 & ~n13532;
  assign n13534 = pi11  & ~n13533;
  assign n13535 = ~pi11  & n13533;
  assign n13536 = ~n13534 & ~n13535;
  assign n13537 = n13511 & n13530;
  assign n13538 = ~n13531 & ~n13537;
  assign n13539 = n13536 & n13538;
  assign n13540 = ~n13531 & ~n13539;
  assign n13541 = n12974 & ~n13540;
  assign n13542 = ~n12974 & n13540;
  assign n13543 = ~n13541 & ~n13542;
  assign n13544 = n3692 & n12431;
  assign n13545 = n12564 & ~n12566;
  assign n13546 = ~n12567 & ~n13545;
  assign n13547 = n880 & n13546;
  assign n13548 = n748 & n12434;
  assign n13549 = n3694 & n12428;
  assign n13550 = ~n13544 & ~n13548;
  assign n13551 = ~n13549 & n13550;
  assign n13552 = ~n13547 & n13551;
  assign n13553 = n13543 & ~n13552;
  assign n13554 = ~n13541 & ~n13553;
  assign n13555 = ~n13353 & n13362;
  assign n13556 = ~n13363 & ~n13555;
  assign n13557 = ~n13554 & n13556;
  assign n13558 = n13554 & ~n13556;
  assign n13559 = ~n13557 & ~n13558;
  assign n13560 = ~n13536 & ~n13538;
  assign n13561 = ~n13539 & ~n13560;
  assign n13562 = n748 & n12437;
  assign n13563 = n12560 & ~n12562;
  assign n13564 = ~n12563 & ~n13563;
  assign n13565 = n880 & n13564;
  assign n13566 = n3692 & n12434;
  assign n13567 = n3694 & n12431;
  assign n13568 = ~n13562 & ~n13566;
  assign n13569 = ~n13567 & n13568;
  assign n13570 = ~n13565 & n13569;
  assign n13571 = n13561 & ~n13570;
  assign n13572 = n13561 & n13570;
  assign n13573 = ~n13561 & ~n13570;
  assign n13574 = ~n13572 & ~n13573;
  assign n13575 = ~n293 & ~n381;
  assign n13576 = ~n520 & ~n561;
  assign n13577 = ~n625 & n13576;
  assign n13578 = n1684 & n13575;
  assign n13579 = n2126 & n3723;
  assign n13580 = n5489 & n13579;
  assign n13581 = n13577 & n13578;
  assign n13582 = n13580 & n13581;
  assign n13583 = ~n183 & ~n235;
  assign n13584 = ~n376 & ~n798;
  assign n13585 = n13583 & n13584;
  assign n13586 = ~n438 & ~n460;
  assign n13587 = ~n754 & n13586;
  assign n13588 = n1538 & n13587;
  assign n13589 = ~n195 & ~n290;
  assign n13590 = ~n297 & ~n370;
  assign n13591 = ~n566 & n13590;
  assign n13592 = n513 & n13589;
  assign n13593 = n1187 & n1306;
  assign n13594 = n2253 & n2284;
  assign n13595 = n13593 & n13594;
  assign n13596 = n13591 & n13592;
  assign n13597 = n4906 & n13585;
  assign n13598 = n13596 & n13597;
  assign n13599 = n1140 & n13595;
  assign n13600 = n3300 & n13588;
  assign n13601 = n13599 & n13600;
  assign n13602 = n13598 & n13601;
  assign n13603 = n2720 & n13602;
  assign n13604 = ~n106 & ~n327;
  assign n13605 = ~n367 & ~n989;
  assign n13606 = n13604 & n13605;
  assign n13607 = n444 & n1074;
  assign n13608 = n3644 & n3988;
  assign n13609 = n13607 & n13608;
  assign n13610 = n1135 & n13606;
  assign n13611 = n2440 & n13318;
  assign n13612 = n13610 & n13611;
  assign n13613 = n13609 & n13612;
  assign n13614 = n13582 & n13613;
  assign n13615 = n4801 & n13614;
  assign n13616 = n13603 & n13615;
  assign n13617 = n13511 & ~n13616;
  assign n13618 = ~n98 & ~n106;
  assign n13619 = ~n193 & ~n382;
  assign n13620 = ~n846 & n13619;
  assign n13621 = n301 & n13618;
  assign n13622 = n660 & n1563;
  assign n13623 = n1578 & n13622;
  assign n13624 = n13620 & n13621;
  assign n13625 = n2149 & n4708;
  assign n13626 = n13624 & n13625;
  assign n13627 = n13623 & n13626;
  assign n13628 = ~n362 & ~n368;
  assign n13629 = n1424 & n13628;
  assign n13630 = ~n235 & ~n409;
  assign n13631 = ~n1002 & n13630;
  assign n13632 = n1176 & n1244;
  assign n13633 = n2360 & n13632;
  assign n13634 = n13629 & n13631;
  assign n13635 = n13633 & n13634;
  assign n13636 = ~n250 & ~n438;
  assign n13637 = ~n486 & ~n768;
  assign n13638 = n13636 & n13637;
  assign n13639 = n883 & n2043;
  assign n13640 = n2609 & n13639;
  assign n13641 = n1477 & n13638;
  assign n13642 = n12687 & n13641;
  assign n13643 = n13640 & n13642;
  assign n13644 = ~n195 & ~n383;
  assign n13645 = ~n443 & n13644;
  assign n13646 = n375 & n799;
  assign n13647 = n940 & n1403;
  assign n13648 = n2801 & n13647;
  assign n13649 = n13645 & n13646;
  assign n13650 = n418 & n1282;
  assign n13651 = n1382 & n13650;
  assign n13652 = n13648 & n13649;
  assign n13653 = n4213 & n13652;
  assign n13654 = n13635 & n13651;
  assign n13655 = n13653 & n13654;
  assign n13656 = n13627 & n13643;
  assign n13657 = n13655 & n13656;
  assign n13658 = n3073 & n13657;
  assign n13659 = ~n356 & ~n810;
  assign n13660 = n1004 & n13659;
  assign n13661 = n2460 & n2472;
  assign n13662 = n13660 & n13661;
  assign n13663 = n2550 & n13662;
  assign n13664 = n2796 & n13663;
  assign n13665 = ~n155 & ~n409;
  assign n13666 = ~n687 & n13665;
  assign n13667 = ~n237 & ~n339;
  assign n13668 = ~n370 & ~n1034;
  assign n13669 = n13667 & n13668;
  assign n13670 = n13666 & n13669;
  assign n13671 = ~n167 & ~n297;
  assign n13672 = ~n329 & ~n594;
  assign n13673 = ~n723 & ~n839;
  assign n13674 = n13672 & n13673;
  assign n13675 = n187 & n13671;
  assign n13676 = n369 & n767;
  assign n13677 = n2528 & n13676;
  assign n13678 = n13674 & n13675;
  assign n13679 = n1702 & n5488;
  assign n13680 = n13678 & n13679;
  assign n13681 = n2684 & n13677;
  assign n13682 = n13670 & n13681;
  assign n13683 = n13680 & n13682;
  assign n13684 = n13664 & n13683;
  assign n13685 = n560 & n2075;
  assign n13686 = n13684 & n13685;
  assign n13687 = ~n13658 & ~n13686;
  assign n13688 = n8242 & n8249;
  assign n13689 = ~n12786 & ~n13688;
  assign n13690 = pi8  & ~n13689;
  assign n13691 = ~pi8  & n13689;
  assign n13692 = ~n13690 & ~n13691;
  assign n13693 = n13658 & n13686;
  assign n13694 = ~n13687 & ~n13693;
  assign n13695 = n13692 & n13694;
  assign n13696 = ~n13687 & ~n13695;
  assign n13697 = n13511 & ~n13696;
  assign n13698 = ~n13511 & n13696;
  assign n13699 = ~n13697 & ~n13698;
  assign n13700 = n3692 & n12440;
  assign n13701 = n12552 & ~n12554;
  assign n13702 = ~n12555 & ~n13701;
  assign n13703 = n880 & n13702;
  assign n13704 = n748 & n12443;
  assign n13705 = n3694 & n12437;
  assign n13706 = ~n13700 & ~n13704;
  assign n13707 = ~n13705 & n13706;
  assign n13708 = ~n13703 & n13707;
  assign n13709 = n13699 & ~n13708;
  assign n13710 = ~n13697 & ~n13709;
  assign n13711 = ~n13511 & n13616;
  assign n13712 = ~n13617 & ~n13711;
  assign n13713 = ~n13710 & n13712;
  assign n13714 = ~n13617 & ~n13713;
  assign n13715 = ~n13574 & ~n13714;
  assign n13716 = ~n13571 & ~n13715;
  assign n13717 = ~n13543 & n13552;
  assign n13718 = ~n13553 & ~n13717;
  assign n13719 = ~n13716 & n13718;
  assign n13720 = n13716 & ~n13718;
  assign n13721 = ~n13719 & ~n13720;
  assign n13722 = n3810 & n12425;
  assign n13723 = n3886 & n13010;
  assign n13724 = n3884 & n12422;
  assign n13725 = n4380 & n12419;
  assign n13726 = ~n13722 & ~n13724;
  assign n13727 = ~n13725 & n13726;
  assign n13728 = ~n13723 & n13727;
  assign n13729 = pi29  & n13728;
  assign n13730 = ~pi29  & ~n13728;
  assign n13731 = ~n13729 & ~n13730;
  assign n13732 = n13721 & ~n13731;
  assign n13733 = ~n13719 & ~n13732;
  assign n13734 = n13559 & ~n13733;
  assign n13735 = ~n13557 & ~n13734;
  assign n13736 = n13475 & ~n13479;
  assign n13737 = ~n13480 & ~n13736;
  assign n13738 = ~n13735 & n13737;
  assign n13739 = ~n13480 & ~n13738;
  assign n13740 = ~n13382 & n13392;
  assign n13741 = ~n13393 & ~n13740;
  assign n13742 = ~n13739 & n13741;
  assign n13743 = n13739 & ~n13741;
  assign n13744 = n86 & n12407;
  assign n13745 = n4420 & n13035;
  assign n13746 = n4600 & n12404;
  assign n13747 = n4615 & n12401;
  assign n13748 = ~n13744 & ~n13746;
  assign n13749 = ~n13747 & n13748;
  assign n13750 = ~n13745 & n13749;
  assign n13751 = pi26  & n13750;
  assign n13752 = ~pi26  & ~n13750;
  assign n13753 = ~n13751 & ~n13752;
  assign n13754 = ~n13743 & ~n13753;
  assign n13755 = ~n13742 & ~n13754;
  assign n13756 = n13465 & ~n13755;
  assign n13757 = ~n13465 & n13755;
  assign n13758 = n5044 & n12395;
  assign n13759 = n5045 & n13144;
  assign n13760 = n5109 & n12362;
  assign n13761 = n5130 & n12392;
  assign n13762 = ~n13758 & ~n13760;
  assign n13763 = ~n13761 & n13762;
  assign n13764 = ~n13759 & n13763;
  assign n13765 = pi23  & n13764;
  assign n13766 = ~pi23  & ~n13764;
  assign n13767 = ~n13765 & ~n13766;
  assign n13768 = ~n13757 & ~n13767;
  assign n13769 = ~n13756 & ~n13768;
  assign n13770 = ~n13461 & ~n13769;
  assign n13771 = ~n13458 & ~n13770;
  assign n13772 = ~n13417 & ~n13418;
  assign n13773 = ~n13430 & n13772;
  assign n13774 = n13430 & ~n13772;
  assign n13775 = ~n13773 & ~n13774;
  assign n13776 = ~n13771 & n13775;
  assign n13777 = n13771 & ~n13775;
  assign n13778 = n5866 & ~n12786;
  assign n13779 = ~n13160 & ~n13181;
  assign n13780 = ~n13279 & ~n13779;
  assign n13781 = ~n13179 & ~n13780;
  assign n13782 = n5241 & ~n13781;
  assign n13783 = n5240 & n13166;
  assign n13784 = n5853 & n13161;
  assign n13785 = ~n13778 & ~n13783;
  assign n13786 = ~n13784 & n13785;
  assign n13787 = ~n13782 & n13786;
  assign n13788 = pi20  & n13787;
  assign n13789 = ~pi20  & ~n13787;
  assign n13790 = ~n13788 & ~n13789;
  assign n13791 = ~n13777 & ~n13790;
  assign n13792 = ~n13776 & ~n13791;
  assign n13793 = n13445 & ~n13792;
  assign n13794 = ~n13445 & n13792;
  assign n13795 = ~n13793 & ~n13794;
  assign n13796 = n5866 & n13161;
  assign n13797 = n5241 & n13183;
  assign n13798 = n5853 & n13166;
  assign n13799 = n5240 & n13164;
  assign n13800 = ~n13798 & ~n13799;
  assign n13801 = ~n13796 & n13800;
  assign n13802 = ~n13797 & n13801;
  assign n13803 = pi20  & n13802;
  assign n13804 = ~pi20  & ~n13802;
  assign n13805 = ~n13803 & ~n13804;
  assign n13806 = ~n13756 & ~n13757;
  assign n13807 = ~n13767 & n13806;
  assign n13808 = n13767 & ~n13806;
  assign n13809 = ~n13807 & ~n13808;
  assign n13810 = n13735 & ~n13737;
  assign n13811 = ~n13738 & ~n13810;
  assign n13812 = n86 & n12410;
  assign n13813 = n4420 & n13093;
  assign n13814 = n4600 & n12407;
  assign n13815 = n4615 & n12404;
  assign n13816 = ~n13812 & ~n13814;
  assign n13817 = ~n13815 & n13816;
  assign n13818 = ~n13813 & n13817;
  assign n13819 = pi26  & n13818;
  assign n13820 = ~pi26  & ~n13818;
  assign n13821 = ~n13819 & ~n13820;
  assign n13822 = n13811 & ~n13821;
  assign n13823 = n13811 & n13821;
  assign n13824 = ~n13811 & ~n13821;
  assign n13825 = ~n13823 & ~n13824;
  assign n13826 = ~n13559 & n13733;
  assign n13827 = ~n13734 & ~n13826;
  assign n13828 = n3810 & n12422;
  assign n13829 = n3886 & n13201;
  assign n13830 = n3884 & n12419;
  assign n13831 = n4380 & n12416;
  assign n13832 = ~n13828 & ~n13830;
  assign n13833 = ~n13831 & n13832;
  assign n13834 = ~n13829 & n13833;
  assign n13835 = pi29  & n13834;
  assign n13836 = ~pi29  & ~n13834;
  assign n13837 = ~n13835 & ~n13836;
  assign n13838 = n13827 & ~n13837;
  assign n13839 = n13827 & n13837;
  assign n13840 = ~n13827 & ~n13837;
  assign n13841 = ~n13839 & ~n13840;
  assign n13842 = n86 & n12413;
  assign n13843 = n4420 & n12891;
  assign n13844 = n4600 & n12410;
  assign n13845 = n4615 & n12407;
  assign n13846 = ~n13842 & ~n13844;
  assign n13847 = ~n13845 & n13846;
  assign n13848 = ~n13843 & n13847;
  assign n13849 = pi26  & n13848;
  assign n13850 = ~pi26  & ~n13848;
  assign n13851 = ~n13849 & ~n13850;
  assign n13852 = ~n13841 & ~n13851;
  assign n13853 = ~n13838 & ~n13852;
  assign n13854 = ~n13825 & ~n13853;
  assign n13855 = ~n13822 & ~n13854;
  assign n13856 = ~n13742 & ~n13743;
  assign n13857 = ~n13753 & n13856;
  assign n13858 = n13753 & ~n13856;
  assign n13859 = ~n13857 & ~n13858;
  assign n13860 = ~n13855 & n13859;
  assign n13861 = n13855 & ~n13859;
  assign n13862 = n5044 & n12398;
  assign n13863 = n5045 & n13245;
  assign n13864 = n5109 & n12395;
  assign n13865 = n5130 & n12362;
  assign n13866 = ~n13862 & ~n13864;
  assign n13867 = ~n13865 & n13866;
  assign n13868 = ~n13863 & n13867;
  assign n13869 = pi23  & n13868;
  assign n13870 = ~pi23  & ~n13868;
  assign n13871 = ~n13869 & ~n13870;
  assign n13872 = ~n13861 & ~n13871;
  assign n13873 = ~n13860 & ~n13872;
  assign n13874 = n13809 & ~n13873;
  assign n13875 = ~n13809 & n13873;
  assign n13876 = n5240 & n12646;
  assign n13877 = n5241 & n13261;
  assign n13878 = n5853 & n13164;
  assign n13879 = n5866 & n13166;
  assign n13880 = ~n13876 & ~n13878;
  assign n13881 = ~n13879 & n13880;
  assign n13882 = ~n13877 & n13881;
  assign n13883 = pi20  & n13882;
  assign n13884 = ~pi20  & ~n13882;
  assign n13885 = ~n13883 & ~n13884;
  assign n13886 = ~n13875 & ~n13885;
  assign n13887 = ~n13874 & ~n13886;
  assign n13888 = ~n13805 & ~n13887;
  assign n13889 = n13461 & n13769;
  assign n13890 = ~n13770 & ~n13889;
  assign n13891 = n13805 & ~n13887;
  assign n13892 = ~n13805 & n13887;
  assign n13893 = ~n13891 & ~n13892;
  assign n13894 = n13890 & ~n13893;
  assign n13895 = ~n13888 & ~n13894;
  assign n13896 = ~n13776 & ~n13777;
  assign n13897 = ~n13790 & n13896;
  assign n13898 = n13790 & ~n13896;
  assign n13899 = ~n13897 & ~n13898;
  assign n13900 = ~n13895 & n13899;
  assign n13901 = n13895 & n13899;
  assign n13902 = ~n13895 & ~n13899;
  assign n13903 = ~n13901 & ~n13902;
  assign n13904 = ~n13890 & n13893;
  assign n13905 = ~n13894 & ~n13904;
  assign n13906 = n5983 & ~n13280;
  assign n13907 = n5982 & ~n13160;
  assign n13908 = ~n6323 & ~n6336;
  assign n13909 = ~n13907 & n13908;
  assign n13910 = ~n12786 & ~n13909;
  assign n13911 = ~n13906 & ~n13910;
  assign n13912 = pi17  & n13911;
  assign n13913 = ~pi17  & ~n13911;
  assign n13914 = ~n13912 & ~n13913;
  assign n13915 = n13825 & n13853;
  assign n13916 = ~n13854 & ~n13915;
  assign n13917 = n5044 & n12401;
  assign n13918 = n5045 & n13108;
  assign n13919 = n5109 & n12398;
  assign n13920 = n5130 & n12395;
  assign n13921 = ~n13917 & ~n13919;
  assign n13922 = ~n13920 & n13921;
  assign n13923 = ~n13918 & n13922;
  assign n13924 = pi23  & n13923;
  assign n13925 = ~pi23  & ~n13923;
  assign n13926 = ~n13924 & ~n13925;
  assign n13927 = n13916 & ~n13926;
  assign n13928 = n13916 & n13926;
  assign n13929 = ~n13916 & ~n13926;
  assign n13930 = ~n13928 & ~n13929;
  assign n13931 = n13841 & n13851;
  assign n13932 = ~n13852 & ~n13931;
  assign n13933 = ~n13721 & n13731;
  assign n13934 = ~n13732 & ~n13933;
  assign n13935 = n13710 & ~n13712;
  assign n13936 = ~n13713 & ~n13935;
  assign n13937 = n748 & n12440;
  assign n13938 = n12556 & ~n12558;
  assign n13939 = ~n12559 & ~n13938;
  assign n13940 = n880 & n13939;
  assign n13941 = n3692 & n12437;
  assign n13942 = n3694 & n12434;
  assign n13943 = ~n13937 & ~n13941;
  assign n13944 = ~n13942 & n13943;
  assign n13945 = ~n13940 & n13944;
  assign n13946 = n13936 & ~n13945;
  assign n13947 = n13936 & n13945;
  assign n13948 = ~n13936 & ~n13945;
  assign n13949 = ~n13947 & ~n13948;
  assign n13950 = n3810 & n12431;
  assign n13951 = n3886 & n13356;
  assign n13952 = n3884 & n12428;
  assign n13953 = n4380 & n12425;
  assign n13954 = ~n13950 & ~n13952;
  assign n13955 = ~n13953 & n13954;
  assign n13956 = ~n13951 & n13955;
  assign n13957 = pi29  & n13956;
  assign n13958 = ~pi29  & ~n13956;
  assign n13959 = ~n13957 & ~n13958;
  assign n13960 = ~n13949 & ~n13959;
  assign n13961 = ~n13946 & ~n13960;
  assign n13962 = ~n13574 & n13714;
  assign n13963 = n13574 & ~n13714;
  assign n13964 = ~n13962 & ~n13963;
  assign n13965 = ~n13961 & ~n13964;
  assign n13966 = n3810 & n12428;
  assign n13967 = n3886 & n13371;
  assign n13968 = n3884 & n12425;
  assign n13969 = n4380 & n12422;
  assign n13970 = ~n13966 & ~n13968;
  assign n13971 = ~n13969 & n13970;
  assign n13972 = ~n13967 & n13971;
  assign n13973 = pi29  & n13972;
  assign n13974 = ~pi29  & ~n13972;
  assign n13975 = ~n13973 & ~n13974;
  assign n13976 = n13961 & n13964;
  assign n13977 = ~n13975 & ~n13976;
  assign n13978 = ~n13965 & ~n13977;
  assign n13979 = n13934 & ~n13978;
  assign n13980 = ~n13934 & n13978;
  assign n13981 = n86 & n12416;
  assign n13982 = n4420 & n12843;
  assign n13983 = n4600 & n12413;
  assign n13984 = n4615 & n12410;
  assign n13985 = ~n13981 & ~n13983;
  assign n13986 = ~n13984 & n13985;
  assign n13987 = ~n13982 & n13986;
  assign n13988 = pi26  & n13987;
  assign n13989 = ~pi26  & ~n13987;
  assign n13990 = ~n13988 & ~n13989;
  assign n13991 = ~n13980 & ~n13990;
  assign n13992 = ~n13979 & ~n13991;
  assign n13993 = n13932 & ~n13992;
  assign n13994 = ~n13932 & n13992;
  assign n13995 = n5044 & n12404;
  assign n13996 = n5045 & n13128;
  assign n13997 = n5109 & n12401;
  assign n13998 = n5130 & n12398;
  assign n13999 = ~n13995 & ~n13997;
  assign n14000 = ~n13998 & n13999;
  assign n14001 = ~n13996 & n14000;
  assign n14002 = pi23  & n14001;
  assign n14003 = ~pi23  & ~n14001;
  assign n14004 = ~n14002 & ~n14003;
  assign n14005 = ~n13994 & ~n14004;
  assign n14006 = ~n13993 & ~n14005;
  assign n14007 = ~n13930 & ~n14006;
  assign n14008 = ~n13927 & ~n14007;
  assign n14009 = ~n13860 & ~n13861;
  assign n14010 = ~n13871 & n14009;
  assign n14011 = n13871 & ~n14009;
  assign n14012 = ~n14010 & ~n14011;
  assign n14013 = ~n14008 & n14012;
  assign n14014 = n14008 & ~n14012;
  assign n14015 = n5240 & n12392;
  assign n14016 = n5241 & n13421;
  assign n14017 = n5853 & n12646;
  assign n14018 = n5866 & n13164;
  assign n14019 = ~n14015 & ~n14017;
  assign n14020 = ~n14018 & n14019;
  assign n14021 = ~n14016 & n14020;
  assign n14022 = pi20  & n14021;
  assign n14023 = ~pi20  & ~n14021;
  assign n14024 = ~n14022 & ~n14023;
  assign n14025 = ~n14014 & ~n14024;
  assign n14026 = ~n14013 & ~n14025;
  assign n14027 = ~n13914 & ~n14026;
  assign n14028 = n13914 & n14026;
  assign n14029 = ~n13874 & ~n13875;
  assign n14030 = ~n13885 & n14029;
  assign n14031 = n13885 & ~n14029;
  assign n14032 = ~n14030 & ~n14031;
  assign n14033 = ~n14028 & n14032;
  assign n14034 = ~n14027 & ~n14033;
  assign n14035 = n13905 & ~n14034;
  assign n14036 = ~n14027 & ~n14028;
  assign n14037 = n14032 & n14036;
  assign n14038 = ~n14032 & ~n14036;
  assign n14039 = ~n14037 & ~n14038;
  assign n14040 = n13930 & n14006;
  assign n14041 = ~n14007 & ~n14040;
  assign n14042 = n5240 & n12362;
  assign n14043 = n5241 & n12652;
  assign n14044 = n5853 & n12392;
  assign n14045 = n5866 & n12646;
  assign n14046 = ~n14042 & ~n14044;
  assign n14047 = ~n14045 & n14046;
  assign n14048 = ~n14043 & n14047;
  assign n14049 = pi20  & n14048;
  assign n14050 = ~pi20  & ~n14048;
  assign n14051 = ~n14049 & ~n14050;
  assign n14052 = n14041 & ~n14051;
  assign n14053 = n14041 & n14051;
  assign n14054 = ~n14041 & ~n14051;
  assign n14055 = ~n14053 & ~n14054;
  assign n14056 = ~n13993 & ~n13994;
  assign n14057 = ~n14004 & n14056;
  assign n14058 = n14004 & ~n14056;
  assign n14059 = ~n14057 & ~n14058;
  assign n14060 = n86 & n12419;
  assign n14061 = n4420 & n12908;
  assign n14062 = n4600 & n12416;
  assign n14063 = n4615 & n12413;
  assign n14064 = ~n14060 & ~n14062;
  assign n14065 = ~n14063 & n14064;
  assign n14066 = ~n14061 & n14065;
  assign n14067 = pi26  & n14066;
  assign n14068 = ~pi26  & ~n14066;
  assign n14069 = ~n14067 & ~n14068;
  assign n14070 = ~n13965 & ~n13976;
  assign n14071 = n13975 & ~n14070;
  assign n14072 = ~n13975 & n14070;
  assign n14073 = ~n14071 & ~n14072;
  assign n14074 = ~n14069 & n14073;
  assign n14075 = n14069 & n14073;
  assign n14076 = ~n14069 & ~n14073;
  assign n14077 = ~n14075 & ~n14076;
  assign n14078 = ~n13699 & n13708;
  assign n14079 = ~n13709 & ~n14078;
  assign n14080 = ~n116 & ~n625;
  assign n14081 = n2007 & n14080;
  assign n14082 = ~n106 & ~n237;
  assign n14083 = ~n594 & ~n1034;
  assign n14084 = n3010 & n14083;
  assign n14085 = n436 & n14082;
  assign n14086 = n600 & n1451;
  assign n14087 = n2891 & n2934;
  assign n14088 = n14086 & n14087;
  assign n14089 = n14084 & n14085;
  assign n14090 = n5632 & n14081;
  assign n14091 = n14089 & n14090;
  assign n14092 = n1111 & n14088;
  assign n14093 = n14091 & n14092;
  assign n14094 = n1150 & n14093;
  assign n14095 = n2648 & n14094;
  assign n14096 = n2738 & n14095;
  assign n14097 = n13658 & ~n14096;
  assign n14098 = n11053 & n11054;
  assign n14099 = ~pi2  & ~n14098;
  assign n14100 = ~n12786 & n14099;
  assign n14101 = pi2  & n12786;
  assign n14102 = ~n14100 & ~n14101;
  assign n14103 = ~n126 & ~n242;
  assign n14104 = ~n308 & ~n309;
  assign n14105 = ~n411 & ~n604;
  assign n14106 = ~n723 & n14105;
  assign n14107 = n14103 & n14104;
  assign n14108 = n150 & n562;
  assign n14109 = n1423 & n2043;
  assign n14110 = n2501 & n14109;
  assign n14111 = n14107 & n14108;
  assign n14112 = n14106 & n14111;
  assign n14113 = n1195 & n14110;
  assign n14114 = n14112 & n14113;
  assign n14115 = ~n415 & ~n435;
  assign n14116 = n431 & n14115;
  assign n14117 = n13585 & n14116;
  assign n14118 = n1473 & n2658;
  assign n14119 = n1910 & n2979;
  assign n14120 = n4302 & n12980;
  assign n14121 = n14119 & n14120;
  assign n14122 = n3720 & n14118;
  assign n14123 = n14117 & n14122;
  assign n14124 = n3308 & n14121;
  assign n14125 = n14123 & n14124;
  assign n14126 = n14114 & n14125;
  assign n14127 = ~n327 & ~n364;
  assign n14128 = n146 & n14127;
  assign n14129 = n1005 & n1510;
  assign n14130 = n3327 & n4004;
  assign n14131 = n14129 & n14130;
  assign n14132 = n4313 & n14128;
  assign n14133 = n14131 & n14132;
  assign n14134 = n6467 & n6971;
  assign n14135 = n14133 & n14134;
  assign n14136 = n4107 & n13490;
  assign n14137 = n14135 & n14136;
  assign n14138 = n14126 & n14137;
  assign n14139 = n14102 & ~n14138;
  assign n14140 = n14102 & n14138;
  assign n14141 = ~n14102 & ~n14138;
  assign n14142 = ~n14140 & ~n14141;
  assign n14143 = ~n10469 & ~n11031;
  assign n14144 = n73 & n14143;
  assign n14145 = ~n12786 & ~n14144;
  assign n14146 = ~pi5  & n14145;
  assign n14147 = pi5  & ~n14145;
  assign n14148 = ~n14146 & ~n14147;
  assign n14149 = ~n14142 & n14148;
  assign n14150 = ~n14139 & ~n14149;
  assign n14151 = n13658 & ~n14150;
  assign n14152 = ~n13658 & n14150;
  assign n14153 = ~n14151 & ~n14152;
  assign n14154 = n3692 & n12449;
  assign n14155 = n12540 & ~n12542;
  assign n14156 = ~n12543 & ~n14155;
  assign n14157 = n880 & n14156;
  assign n14158 = n748 & n12452;
  assign n14159 = n3694 & n12446;
  assign n14160 = ~n14154 & ~n14158;
  assign n14161 = ~n14159 & n14160;
  assign n14162 = ~n14157 & n14161;
  assign n14163 = n14153 & ~n14162;
  assign n14164 = ~n14151 & ~n14163;
  assign n14165 = ~n13658 & n14096;
  assign n14166 = ~n14097 & ~n14165;
  assign n14167 = ~n14164 & n14166;
  assign n14168 = ~n14097 & ~n14167;
  assign n14169 = ~n13692 & ~n13694;
  assign n14170 = ~n13695 & ~n14169;
  assign n14171 = ~n14168 & n14170;
  assign n14172 = n14168 & ~n14170;
  assign n14173 = n748 & n12446;
  assign n14174 = n12548 & ~n12550;
  assign n14175 = ~n12551 & ~n14174;
  assign n14176 = n880 & n14175;
  assign n14177 = n3692 & n12443;
  assign n14178 = n3694 & n12440;
  assign n14179 = ~n14173 & ~n14177;
  assign n14180 = ~n14178 & n14179;
  assign n14181 = ~n14176 & n14180;
  assign n14182 = ~n14172 & ~n14181;
  assign n14183 = ~n14171 & ~n14182;
  assign n14184 = n14079 & ~n14183;
  assign n14185 = ~n14079 & n14183;
  assign n14186 = ~n14184 & ~n14185;
  assign n14187 = n3810 & n12434;
  assign n14188 = n3886 & n13546;
  assign n14189 = n3884 & n12431;
  assign n14190 = n4380 & n12428;
  assign n14191 = ~n14187 & ~n14189;
  assign n14192 = ~n14190 & n14191;
  assign n14193 = ~n14188 & n14192;
  assign n14194 = pi29  & n14193;
  assign n14195 = ~pi29  & ~n14193;
  assign n14196 = ~n14194 & ~n14195;
  assign n14197 = n14186 & ~n14196;
  assign n14198 = ~n14184 & ~n14197;
  assign n14199 = n13949 & n13959;
  assign n14200 = ~n13960 & ~n14199;
  assign n14201 = ~n14198 & n14200;
  assign n14202 = n14198 & ~n14200;
  assign n14203 = n86 & n12422;
  assign n14204 = n4420 & n13201;
  assign n14205 = n4600 & n12419;
  assign n14206 = n4615 & n12416;
  assign n14207 = ~n14203 & ~n14205;
  assign n14208 = ~n14206 & n14207;
  assign n14209 = ~n14204 & n14208;
  assign n14210 = pi26  & n14209;
  assign n14211 = ~pi26  & ~n14209;
  assign n14212 = ~n14210 & ~n14211;
  assign n14213 = ~n14202 & ~n14212;
  assign n14214 = ~n14201 & ~n14213;
  assign n14215 = ~n14077 & ~n14214;
  assign n14216 = ~n14074 & ~n14215;
  assign n14217 = ~n13979 & ~n13980;
  assign n14218 = ~n13990 & n14217;
  assign n14219 = n13990 & ~n14217;
  assign n14220 = ~n14218 & ~n14219;
  assign n14221 = ~n14216 & n14220;
  assign n14222 = n14216 & ~n14220;
  assign n14223 = n5044 & n12407;
  assign n14224 = n5045 & n13035;
  assign n14225 = n5109 & n12404;
  assign n14226 = n5130 & n12401;
  assign n14227 = ~n14223 & ~n14225;
  assign n14228 = ~n14226 & n14227;
  assign n14229 = ~n14224 & n14228;
  assign n14230 = pi23  & n14229;
  assign n14231 = ~pi23  & ~n14229;
  assign n14232 = ~n14230 & ~n14231;
  assign n14233 = ~n14222 & ~n14232;
  assign n14234 = ~n14221 & ~n14233;
  assign n14235 = n14059 & ~n14234;
  assign n14236 = ~n14059 & n14234;
  assign n14237 = n5240 & n12395;
  assign n14238 = n5241 & n13144;
  assign n14239 = n5853 & n12362;
  assign n14240 = n5866 & n12392;
  assign n14241 = ~n14237 & ~n14239;
  assign n14242 = ~n14240 & n14241;
  assign n14243 = ~n14238 & n14242;
  assign n14244 = pi20  & n14243;
  assign n14245 = ~pi20  & ~n14243;
  assign n14246 = ~n14244 & ~n14245;
  assign n14247 = ~n14236 & ~n14246;
  assign n14248 = ~n14235 & ~n14247;
  assign n14249 = ~n14055 & ~n14248;
  assign n14250 = ~n14052 & ~n14249;
  assign n14251 = ~n14013 & ~n14014;
  assign n14252 = ~n14024 & n14251;
  assign n14253 = n14024 & ~n14251;
  assign n14254 = ~n14252 & ~n14253;
  assign n14255 = ~n14250 & n14254;
  assign n14256 = n14250 & ~n14254;
  assign n14257 = n6336 & ~n12786;
  assign n14258 = n5983 & ~n13781;
  assign n14259 = n5982 & n13166;
  assign n14260 = n6323 & n13161;
  assign n14261 = ~n14257 & ~n14259;
  assign n14262 = ~n14260 & n14261;
  assign n14263 = ~n14258 & n14262;
  assign n14264 = pi17  & n14263;
  assign n14265 = ~pi17  & ~n14263;
  assign n14266 = ~n14264 & ~n14265;
  assign n14267 = ~n14256 & ~n14266;
  assign n14268 = ~n14255 & ~n14267;
  assign n14269 = n14039 & ~n14268;
  assign n14270 = ~n14039 & n14268;
  assign n14271 = ~n14269 & ~n14270;
  assign n14272 = n6336 & n13161;
  assign n14273 = n5983 & n13183;
  assign n14274 = n6323 & n13166;
  assign n14275 = n5982 & n13164;
  assign n14276 = ~n14274 & ~n14275;
  assign n14277 = ~n14272 & n14276;
  assign n14278 = ~n14273 & n14277;
  assign n14279 = pi17  & n14278;
  assign n14280 = ~pi17  & ~n14278;
  assign n14281 = ~n14279 & ~n14280;
  assign n14282 = ~n14235 & ~n14236;
  assign n14283 = ~n14246 & n14282;
  assign n14284 = n14246 & ~n14282;
  assign n14285 = ~n14283 & ~n14284;
  assign n14286 = n14077 & n14214;
  assign n14287 = ~n14215 & ~n14286;
  assign n14288 = n5044 & n12410;
  assign n14289 = n5045 & n13093;
  assign n14290 = n5109 & n12407;
  assign n14291 = n5130 & n12404;
  assign n14292 = ~n14288 & ~n14290;
  assign n14293 = ~n14291 & n14292;
  assign n14294 = ~n14289 & n14293;
  assign n14295 = pi23  & n14294;
  assign n14296 = ~pi23  & ~n14294;
  assign n14297 = ~n14295 & ~n14296;
  assign n14298 = n14287 & ~n14297;
  assign n14299 = n14287 & n14297;
  assign n14300 = ~n14287 & ~n14297;
  assign n14301 = ~n14299 & ~n14300;
  assign n14302 = ~n14201 & ~n14202;
  assign n14303 = ~n14212 & n14302;
  assign n14304 = n14212 & ~n14302;
  assign n14305 = ~n14303 & ~n14304;
  assign n14306 = n3810 & n12437;
  assign n14307 = n3886 & n13564;
  assign n14308 = n3884 & n12434;
  assign n14309 = n4380 & n12431;
  assign n14310 = ~n14306 & ~n14308;
  assign n14311 = ~n14309 & n14310;
  assign n14312 = ~n14307 & n14311;
  assign n14313 = pi29  & n14312;
  assign n14314 = ~pi29  & ~n14312;
  assign n14315 = ~n14313 & ~n14314;
  assign n14316 = ~n14171 & ~n14172;
  assign n14317 = ~n14181 & n14316;
  assign n14318 = n14181 & ~n14316;
  assign n14319 = ~n14317 & ~n14318;
  assign n14320 = ~n14315 & n14319;
  assign n14321 = n14164 & ~n14166;
  assign n14322 = ~n14167 & ~n14321;
  assign n14323 = n748 & n12449;
  assign n14324 = n12544 & ~n12546;
  assign n14325 = ~n12547 & ~n14324;
  assign n14326 = n880 & n14325;
  assign n14327 = n3692 & n12446;
  assign n14328 = n3694 & n12443;
  assign n14329 = ~n14323 & ~n14327;
  assign n14330 = ~n14328 & n14329;
  assign n14331 = ~n14326 & n14330;
  assign n14332 = n14322 & ~n14331;
  assign n14333 = n14322 & n14331;
  assign n14334 = ~n14322 & ~n14331;
  assign n14335 = ~n14333 & ~n14334;
  assign n14336 = ~n145 & ~n159;
  assign n14337 = ~n171 & ~n174;
  assign n14338 = ~n376 & ~n525;
  assign n14339 = ~n663 & ~n1051;
  assign n14340 = n14338 & n14339;
  assign n14341 = n14336 & n14337;
  assign n14342 = n1403 & n2682;
  assign n14343 = n2892 & n3033;
  assign n14344 = n14342 & n14343;
  assign n14345 = n14340 & n14341;
  assign n14346 = n14344 & n14345;
  assign n14347 = n2110 & n3379;
  assign n14348 = n14346 & n14347;
  assign n14349 = n326 & n14348;
  assign n14350 = n823 & n14349;
  assign n14351 = n4033 & n14350;
  assign n14352 = ~n14102 & ~n14351;
  assign n14353 = ~n304 & n1429;
  assign n14354 = n12930 & n14353;
  assign n14355 = ~n116 & ~n253;
  assign n14356 = ~n270 & ~n718;
  assign n14357 = n533 & n14355;
  assign n14358 = n1151 & n14356;
  assign n14359 = n2157 & n2561;
  assign n14360 = n2757 & n4687;
  assign n14361 = n14359 & n14360;
  assign n14362 = n14357 & n14358;
  assign n14363 = n2748 & n3655;
  assign n14364 = n14362 & n14363;
  assign n14365 = n12721 & n14361;
  assign n14366 = n14354 & n14365;
  assign n14367 = n1569 & n14364;
  assign n14368 = n1778 & n14367;
  assign n14369 = n14366 & n14368;
  assign n14370 = n14126 & n14369;
  assign n14371 = ~n14102 & ~n14370;
  assign n14372 = n14102 & n14370;
  assign n14373 = ~n14371 & ~n14372;
  assign n14374 = ~n510 & ~n639;
  assign n14375 = ~n937 & n14374;
  assign n14376 = n4925 & n6929;
  assign n14377 = n14375 & n14376;
  assign n14378 = n1021 & n14377;
  assign n14379 = ~n592 & ~n648;
  assign n14380 = ~n1032 & n14379;
  assign n14381 = ~n245 & ~n566;
  assign n14382 = ~n1699 & n14381;
  assign n14383 = n565 & n2837;
  assign n14384 = n3007 & n14383;
  assign n14385 = n14382 & n14384;
  assign n14386 = ~n149 & ~n276;
  assign n14387 = ~n334 & ~n355;
  assign n14388 = ~n638 & n14387;
  assign n14389 = n487 & n14386;
  assign n14390 = n1486 & n2167;
  assign n14391 = n3204 & n14390;
  assign n14392 = n14388 & n14389;
  assign n14393 = n3936 & n4110;
  assign n14394 = n14392 & n14393;
  assign n14395 = n14391 & n14394;
  assign n14396 = n2525 & n14385;
  assign n14397 = n14395 & n14396;
  assign n14398 = ~n174 & ~n309;
  assign n14399 = ~n364 & n14398;
  assign n14400 = n2254 & n2528;
  assign n14401 = n14399 & n14400;
  assign n14402 = n14397 & n14401;
  assign n14403 = ~n171 & ~n353;
  assign n14404 = ~n368 & ~n1002;
  assign n14405 = n14403 & n14404;
  assign n14406 = n298 & n1576;
  assign n14407 = n3407 & n14406;
  assign n14408 = n219 & n14405;
  assign n14409 = n13585 & n14380;
  assign n14410 = n14408 & n14409;
  assign n14411 = n2575 & n14407;
  assign n14412 = n14410 & n14411;
  assign n14413 = n14378 & n14412;
  assign n14414 = n12869 & n14413;
  assign n14415 = n14402 & n14414;
  assign n14416 = ~n14102 & ~n14415;
  assign n14417 = n14102 & n14415;
  assign n14418 = n748 & n12464;
  assign n14419 = n12524 & ~n12526;
  assign n14420 = ~n12527 & ~n14419;
  assign n14421 = n880 & n14420;
  assign n14422 = n3692 & n12461;
  assign n14423 = n3694 & n12458;
  assign n14424 = ~n14418 & ~n14422;
  assign n14425 = ~n14423 & n14424;
  assign n14426 = ~n14421 & n14425;
  assign n14427 = ~n14417 & ~n14426;
  assign n14428 = ~n14416 & ~n14427;
  assign n14429 = n14373 & ~n14428;
  assign n14430 = ~n14371 & ~n14429;
  assign n14431 = n14102 & n14351;
  assign n14432 = ~n14352 & ~n14431;
  assign n14433 = ~n14430 & n14432;
  assign n14434 = ~n14352 & ~n14433;
  assign n14435 = n14142 & ~n14148;
  assign n14436 = ~n14149 & ~n14435;
  assign n14437 = ~n14434 & n14436;
  assign n14438 = n14434 & ~n14436;
  assign n14439 = ~n14437 & ~n14438;
  assign n14440 = n748 & n12455;
  assign n14441 = n12536 & ~n12538;
  assign n14442 = ~n12539 & ~n14441;
  assign n14443 = n880 & n14442;
  assign n14444 = n3692 & n12452;
  assign n14445 = n3694 & n12449;
  assign n14446 = ~n14440 & ~n14444;
  assign n14447 = ~n14445 & n14446;
  assign n14448 = ~n14443 & n14447;
  assign n14449 = n14439 & ~n14448;
  assign n14450 = ~n14437 & ~n14449;
  assign n14451 = ~n14153 & n14162;
  assign n14452 = ~n14163 & ~n14451;
  assign n14453 = ~n14450 & n14452;
  assign n14454 = n14450 & ~n14452;
  assign n14455 = ~n14453 & ~n14454;
  assign n14456 = n3810 & n12443;
  assign n14457 = n3886 & n13702;
  assign n14458 = n3884 & n12440;
  assign n14459 = n4380 & n12437;
  assign n14460 = ~n14456 & ~n14458;
  assign n14461 = ~n14459 & n14460;
  assign n14462 = ~n14457 & n14461;
  assign n14463 = pi29  & n14462;
  assign n14464 = ~pi29  & ~n14462;
  assign n14465 = ~n14463 & ~n14464;
  assign n14466 = n14455 & ~n14465;
  assign n14467 = ~n14453 & ~n14466;
  assign n14468 = ~n14335 & ~n14467;
  assign n14469 = ~n14332 & ~n14468;
  assign n14470 = n14315 & ~n14319;
  assign n14471 = ~n14320 & ~n14470;
  assign n14472 = ~n14469 & n14471;
  assign n14473 = ~n14320 & ~n14472;
  assign n14474 = ~n14186 & n14196;
  assign n14475 = ~n14197 & ~n14474;
  assign n14476 = ~n14473 & n14475;
  assign n14477 = n14473 & ~n14475;
  assign n14478 = n86 & n12425;
  assign n14479 = n4420 & n13010;
  assign n14480 = n4600 & n12422;
  assign n14481 = n4615 & n12419;
  assign n14482 = ~n14478 & ~n14480;
  assign n14483 = ~n14481 & n14482;
  assign n14484 = ~n14479 & n14483;
  assign n14485 = pi26  & n14484;
  assign n14486 = ~pi26  & ~n14484;
  assign n14487 = ~n14485 & ~n14486;
  assign n14488 = ~n14477 & ~n14487;
  assign n14489 = ~n14476 & ~n14488;
  assign n14490 = n14305 & ~n14489;
  assign n14491 = ~n14305 & n14489;
  assign n14492 = n5044 & n12413;
  assign n14493 = n5045 & n12891;
  assign n14494 = n5109 & n12410;
  assign n14495 = n5130 & n12407;
  assign n14496 = ~n14492 & ~n14494;
  assign n14497 = ~n14495 & n14496;
  assign n14498 = ~n14493 & n14497;
  assign n14499 = pi23  & n14498;
  assign n14500 = ~pi23  & ~n14498;
  assign n14501 = ~n14499 & ~n14500;
  assign n14502 = ~n14491 & ~n14501;
  assign n14503 = ~n14490 & ~n14502;
  assign n14504 = ~n14301 & ~n14503;
  assign n14505 = ~n14298 & ~n14504;
  assign n14506 = ~n14221 & ~n14222;
  assign n14507 = ~n14232 & n14506;
  assign n14508 = n14232 & ~n14506;
  assign n14509 = ~n14507 & ~n14508;
  assign n14510 = ~n14505 & n14509;
  assign n14511 = n14505 & ~n14509;
  assign n14512 = n5240 & n12398;
  assign n14513 = n5241 & n13245;
  assign n14514 = n5853 & n12395;
  assign n14515 = n5866 & n12362;
  assign n14516 = ~n14512 & ~n14514;
  assign n14517 = ~n14515 & n14516;
  assign n14518 = ~n14513 & n14517;
  assign n14519 = pi20  & n14518;
  assign n14520 = ~pi20  & ~n14518;
  assign n14521 = ~n14519 & ~n14520;
  assign n14522 = ~n14511 & ~n14521;
  assign n14523 = ~n14510 & ~n14522;
  assign n14524 = n14285 & ~n14523;
  assign n14525 = ~n14285 & n14523;
  assign n14526 = n5982 & n12646;
  assign n14527 = n5983 & n13261;
  assign n14528 = n6323 & n13164;
  assign n14529 = n6336 & n13166;
  assign n14530 = ~n14526 & ~n14528;
  assign n14531 = ~n14529 & n14530;
  assign n14532 = ~n14527 & n14531;
  assign n14533 = pi17  & n14532;
  assign n14534 = ~pi17  & ~n14532;
  assign n14535 = ~n14533 & ~n14534;
  assign n14536 = ~n14525 & ~n14535;
  assign n14537 = ~n14524 & ~n14536;
  assign n14538 = ~n14281 & ~n14537;
  assign n14539 = n14055 & n14248;
  assign n14540 = ~n14249 & ~n14539;
  assign n14541 = n14281 & ~n14537;
  assign n14542 = ~n14281 & n14537;
  assign n14543 = ~n14541 & ~n14542;
  assign n14544 = n14540 & ~n14543;
  assign n14545 = ~n14538 & ~n14544;
  assign n14546 = ~n14255 & ~n14256;
  assign n14547 = ~n14266 & n14546;
  assign n14548 = n14266 & ~n14546;
  assign n14549 = ~n14547 & ~n14548;
  assign n14550 = ~n14545 & n14549;
  assign n14551 = n14545 & n14549;
  assign n14552 = ~n14545 & ~n14549;
  assign n14553 = ~n14551 & ~n14552;
  assign n14554 = ~n14540 & n14543;
  assign n14555 = ~n14544 & ~n14554;
  assign n14556 = n6631 & ~n13280;
  assign n14557 = n6630 & ~n13160;
  assign n14558 = ~n7238 & ~n7262;
  assign n14559 = ~n14557 & n14558;
  assign n14560 = ~n12786 & ~n14559;
  assign n14561 = ~n14556 & ~n14560;
  assign n14562 = pi14  & n14561;
  assign n14563 = ~pi14  & ~n14561;
  assign n14564 = ~n14562 & ~n14563;
  assign n14565 = n14301 & n14503;
  assign n14566 = ~n14504 & ~n14565;
  assign n14567 = n5240 & n12401;
  assign n14568 = n5241 & n13108;
  assign n14569 = n5853 & n12398;
  assign n14570 = n5866 & n12395;
  assign n14571 = ~n14567 & ~n14569;
  assign n14572 = ~n14570 & n14571;
  assign n14573 = ~n14568 & n14572;
  assign n14574 = pi20  & n14573;
  assign n14575 = ~pi20  & ~n14573;
  assign n14576 = ~n14574 & ~n14575;
  assign n14577 = n14566 & ~n14576;
  assign n14578 = n14566 & n14576;
  assign n14579 = ~n14566 & ~n14576;
  assign n14580 = ~n14578 & ~n14579;
  assign n14581 = ~n14490 & ~n14491;
  assign n14582 = ~n14501 & n14581;
  assign n14583 = n14501 & ~n14581;
  assign n14584 = ~n14582 & ~n14583;
  assign n14585 = n14469 & ~n14471;
  assign n14586 = ~n14472 & ~n14585;
  assign n14587 = n86 & n12428;
  assign n14588 = n4420 & n13371;
  assign n14589 = n4600 & n12425;
  assign n14590 = n4615 & n12422;
  assign n14591 = ~n14587 & ~n14589;
  assign n14592 = ~n14590 & n14591;
  assign n14593 = ~n14588 & n14592;
  assign n14594 = pi26  & n14593;
  assign n14595 = ~pi26  & ~n14593;
  assign n14596 = ~n14594 & ~n14595;
  assign n14597 = n14586 & ~n14596;
  assign n14598 = n14586 & n14596;
  assign n14599 = ~n14586 & ~n14596;
  assign n14600 = ~n14598 & ~n14599;
  assign n14601 = n14335 & n14467;
  assign n14602 = ~n14468 & ~n14601;
  assign n14603 = n3810 & n12440;
  assign n14604 = n3886 & n13939;
  assign n14605 = n3884 & n12437;
  assign n14606 = n4380 & n12434;
  assign n14607 = ~n14603 & ~n14605;
  assign n14608 = ~n14606 & n14607;
  assign n14609 = ~n14604 & n14608;
  assign n14610 = pi29  & n14609;
  assign n14611 = ~pi29  & ~n14609;
  assign n14612 = ~n14610 & ~n14611;
  assign n14613 = n14602 & ~n14612;
  assign n14614 = n14602 & n14612;
  assign n14615 = ~n14602 & ~n14612;
  assign n14616 = ~n14614 & ~n14615;
  assign n14617 = n86 & n12431;
  assign n14618 = n4420 & n13356;
  assign n14619 = n4600 & n12428;
  assign n14620 = n4615 & n12425;
  assign n14621 = ~n14617 & ~n14619;
  assign n14622 = ~n14620 & n14621;
  assign n14623 = ~n14618 & n14622;
  assign n14624 = pi26  & n14623;
  assign n14625 = ~pi26  & ~n14623;
  assign n14626 = ~n14624 & ~n14625;
  assign n14627 = ~n14616 & ~n14626;
  assign n14628 = ~n14613 & ~n14627;
  assign n14629 = ~n14600 & ~n14628;
  assign n14630 = ~n14597 & ~n14629;
  assign n14631 = ~n14476 & ~n14477;
  assign n14632 = ~n14487 & n14631;
  assign n14633 = n14487 & ~n14631;
  assign n14634 = ~n14632 & ~n14633;
  assign n14635 = ~n14630 & n14634;
  assign n14636 = n14630 & ~n14634;
  assign n14637 = n5044 & n12416;
  assign n14638 = n5045 & n12843;
  assign n14639 = n5109 & n12413;
  assign n14640 = n5130 & n12410;
  assign n14641 = ~n14637 & ~n14639;
  assign n14642 = ~n14640 & n14641;
  assign n14643 = ~n14638 & n14642;
  assign n14644 = pi23  & n14643;
  assign n14645 = ~pi23  & ~n14643;
  assign n14646 = ~n14644 & ~n14645;
  assign n14647 = ~n14636 & ~n14646;
  assign n14648 = ~n14635 & ~n14647;
  assign n14649 = n14584 & ~n14648;
  assign n14650 = ~n14584 & n14648;
  assign n14651 = n5240 & n12404;
  assign n14652 = n5241 & n13128;
  assign n14653 = n5853 & n12401;
  assign n14654 = n5866 & n12398;
  assign n14655 = ~n14651 & ~n14653;
  assign n14656 = ~n14654 & n14655;
  assign n14657 = ~n14652 & n14656;
  assign n14658 = pi20  & n14657;
  assign n14659 = ~pi20  & ~n14657;
  assign n14660 = ~n14658 & ~n14659;
  assign n14661 = ~n14650 & ~n14660;
  assign n14662 = ~n14649 & ~n14661;
  assign n14663 = ~n14580 & ~n14662;
  assign n14664 = ~n14577 & ~n14663;
  assign n14665 = ~n14510 & ~n14511;
  assign n14666 = ~n14521 & n14665;
  assign n14667 = n14521 & ~n14665;
  assign n14668 = ~n14666 & ~n14667;
  assign n14669 = ~n14664 & n14668;
  assign n14670 = n14664 & ~n14668;
  assign n14671 = n5982 & n12392;
  assign n14672 = n5983 & n13421;
  assign n14673 = n6323 & n12646;
  assign n14674 = n6336 & n13164;
  assign n14675 = ~n14671 & ~n14673;
  assign n14676 = ~n14674 & n14675;
  assign n14677 = ~n14672 & n14676;
  assign n14678 = pi17  & n14677;
  assign n14679 = ~pi17  & ~n14677;
  assign n14680 = ~n14678 & ~n14679;
  assign n14681 = ~n14670 & ~n14680;
  assign n14682 = ~n14669 & ~n14681;
  assign n14683 = ~n14564 & ~n14682;
  assign n14684 = n14564 & n14682;
  assign n14685 = ~n14524 & ~n14525;
  assign n14686 = ~n14535 & n14685;
  assign n14687 = n14535 & ~n14685;
  assign n14688 = ~n14686 & ~n14687;
  assign n14689 = ~n14684 & n14688;
  assign n14690 = ~n14683 & ~n14689;
  assign n14691 = n14555 & ~n14690;
  assign n14692 = ~n14683 & ~n14684;
  assign n14693 = n14688 & n14692;
  assign n14694 = ~n14688 & ~n14692;
  assign n14695 = ~n14693 & ~n14694;
  assign n14696 = n14580 & n14662;
  assign n14697 = ~n14663 & ~n14696;
  assign n14698 = n5982 & n12362;
  assign n14699 = n5983 & n12652;
  assign n14700 = n6323 & n12392;
  assign n14701 = n6336 & n12646;
  assign n14702 = ~n14698 & ~n14700;
  assign n14703 = ~n14701 & n14702;
  assign n14704 = ~n14699 & n14703;
  assign n14705 = pi17  & n14704;
  assign n14706 = ~pi17  & ~n14704;
  assign n14707 = ~n14705 & ~n14706;
  assign n14708 = n14697 & ~n14707;
  assign n14709 = n14697 & n14707;
  assign n14710 = ~n14697 & ~n14707;
  assign n14711 = ~n14709 & ~n14710;
  assign n14712 = ~n14649 & ~n14650;
  assign n14713 = ~n14660 & n14712;
  assign n14714 = n14660 & ~n14712;
  assign n14715 = ~n14713 & ~n14714;
  assign n14716 = n14600 & n14628;
  assign n14717 = ~n14629 & ~n14716;
  assign n14718 = n5044 & n12419;
  assign n14719 = n5045 & n12908;
  assign n14720 = n5109 & n12416;
  assign n14721 = n5130 & n12413;
  assign n14722 = ~n14718 & ~n14720;
  assign n14723 = ~n14721 & n14722;
  assign n14724 = ~n14719 & n14723;
  assign n14725 = pi23  & n14724;
  assign n14726 = ~pi23  & ~n14724;
  assign n14727 = ~n14725 & ~n14726;
  assign n14728 = n14717 & ~n14727;
  assign n14729 = n14717 & n14727;
  assign n14730 = ~n14717 & ~n14727;
  assign n14731 = ~n14729 & ~n14730;
  assign n14732 = ~n14616 & n14626;
  assign n14733 = n14616 & ~n14626;
  assign n14734 = ~n14732 & ~n14733;
  assign n14735 = ~n14455 & n14465;
  assign n14736 = ~n14466 & ~n14735;
  assign n14737 = n14430 & ~n14432;
  assign n14738 = ~n14433 & ~n14737;
  assign n14739 = n748 & n12458;
  assign n14740 = n12532 & ~n12534;
  assign n14741 = ~n12535 & ~n14740;
  assign n14742 = n880 & n14741;
  assign n14743 = n3692 & n12455;
  assign n14744 = n3694 & n12452;
  assign n14745 = ~n14739 & ~n14743;
  assign n14746 = ~n14744 & n14745;
  assign n14747 = ~n14742 & n14746;
  assign n14748 = n14738 & ~n14747;
  assign n14749 = n14738 & n14747;
  assign n14750 = ~n14738 & ~n14747;
  assign n14751 = ~n14749 & ~n14750;
  assign n14752 = ~n14373 & n14428;
  assign n14753 = ~n14429 & ~n14752;
  assign n14754 = n748 & n12461;
  assign n14755 = n12528 & ~n12530;
  assign n14756 = ~n12531 & ~n14755;
  assign n14757 = n880 & n14756;
  assign n14758 = n3692 & n12458;
  assign n14759 = n3694 & n12455;
  assign n14760 = ~n14754 & ~n14758;
  assign n14761 = ~n14759 & n14760;
  assign n14762 = ~n14757 & n14761;
  assign n14763 = n14753 & ~n14762;
  assign n14764 = n14753 & n14762;
  assign n14765 = ~n14753 & ~n14762;
  assign n14766 = ~n14764 & ~n14765;
  assign n14767 = ~n98 & ~n235;
  assign n14768 = ~n526 & ~n661;
  assign n14769 = ~n1034 & n14768;
  assign n14770 = n14767 & n14769;
  assign n14771 = n3704 & n14770;
  assign n14772 = ~n106 & ~n129;
  assign n14773 = ~n216 & n14772;
  assign n14774 = n354 & n375;
  assign n14775 = n593 & n1230;
  assign n14776 = n1383 & n3409;
  assign n14777 = n14775 & n14776;
  assign n14778 = n14773 & n14774;
  assign n14779 = n3385 & n4266;
  assign n14780 = n14778 & n14779;
  assign n14781 = n2971 & n14777;
  assign n14782 = n13494 & n14781;
  assign n14783 = n14771 & n14780;
  assign n14784 = n14782 & n14783;
  assign n14785 = n1696 & n14784;
  assign n14786 = n5322 & n14785;
  assign n14787 = n3692 & n12464;
  assign n14788 = n12520 & ~n12522;
  assign n14789 = ~n12523 & ~n14788;
  assign n14790 = n880 & n14789;
  assign n14791 = n748 & n12467;
  assign n14792 = n3694 & n12461;
  assign n14793 = ~n14787 & ~n14791;
  assign n14794 = ~n14792 & n14793;
  assign n14795 = ~n14790 & n14794;
  assign n14796 = ~n14786 & ~n14795;
  assign n14797 = ~n155 & ~n291;
  assign n14798 = ~n317 & ~n376;
  assign n14799 = ~n415 & ~n814;
  assign n14800 = n14798 & n14799;
  assign n14801 = n1424 & n14797;
  assign n14802 = n1452 & n2042;
  assign n14803 = n3408 & n3459;
  assign n14804 = n4164 & n14803;
  assign n14805 = n14801 & n14802;
  assign n14806 = n14800 & n14805;
  assign n14807 = n3127 & n14804;
  assign n14808 = n14806 & n14807;
  assign n14809 = n714 & n6410;
  assign n14810 = n14808 & n14809;
  assign n14811 = n1562 & n14810;
  assign n14812 = n1984 & n14811;
  assign n14813 = n3692 & n12467;
  assign n14814 = n12516 & ~n12518;
  assign n14815 = ~n12519 & ~n14814;
  assign n14816 = n880 & n14815;
  assign n14817 = n748 & n12470;
  assign n14818 = n3694 & n12464;
  assign n14819 = ~n14813 & ~n14817;
  assign n14820 = ~n14818 & n14819;
  assign n14821 = ~n14816 & n14820;
  assign n14822 = ~n14812 & ~n14821;
  assign n14823 = ~n302 & ~n378;
  assign n14824 = ~n411 & ~n502;
  assign n14825 = ~n723 & n14824;
  assign n14826 = n602 & n14823;
  assign n14827 = n1890 & n2451;
  assign n14828 = n14826 & n14827;
  assign n14829 = n2396 & n14825;
  assign n14830 = n3324 & n3646;
  assign n14831 = n4829 & n14830;
  assign n14832 = n14828 & n14829;
  assign n14833 = n14831 & n14832;
  assign n14834 = n3253 & n14833;
  assign n14835 = n2519 & n14834;
  assign n14836 = n14402 & n14835;
  assign n14837 = n3692 & n12470;
  assign n14838 = n12512 & ~n12514;
  assign n14839 = ~n12515 & ~n14838;
  assign n14840 = n880 & n14839;
  assign n14841 = n748 & n12473;
  assign n14842 = n3694 & n12467;
  assign n14843 = ~n14837 & ~n14841;
  assign n14844 = ~n14842 & n14843;
  assign n14845 = ~n14840 & n14844;
  assign n14846 = ~n14836 & ~n14845;
  assign n14847 = n3692 & n12473;
  assign n14848 = n12508 & ~n12510;
  assign n14849 = ~n12511 & ~n14848;
  assign n14850 = n880 & n14849;
  assign n14851 = n748 & n12476;
  assign n14852 = n3694 & n12470;
  assign n14853 = ~n14847 & ~n14851;
  assign n14854 = ~n14852 & n14853;
  assign n14855 = ~n14850 & n14854;
  assign n14856 = ~n93 & ~n299;
  assign n14857 = ~n312 & ~n329;
  assign n14858 = n14856 & n14857;
  assign n14859 = n1151 & n1884;
  assign n14860 = n14858 & n14859;
  assign n14861 = ~n193 & ~n197;
  assign n14862 = ~n291 & ~n480;
  assign n14863 = n14861 & n14862;
  assign n14864 = n164 & n1270;
  assign n14865 = n1351 & n2201;
  assign n14866 = n4887 & n14865;
  assign n14867 = n14863 & n14864;
  assign n14868 = n717 & n2396;
  assign n14869 = n14867 & n14868;
  assign n14870 = n14860 & n14866;
  assign n14871 = n14869 & n14870;
  assign n14872 = n1059 & n4300;
  assign n14873 = n14871 & n14872;
  assign n14874 = n4101 & n14873;
  assign n14875 = ~n14855 & ~n14874;
  assign n14876 = ~n167 & ~n355;
  assign n14877 = ~n1487 & n14876;
  assign n14878 = ~n129 & ~n273;
  assign n14879 = ~n333 & ~n482;
  assign n14880 = ~n525 & ~n536;
  assign n14881 = ~n636 & n14880;
  assign n14882 = n14878 & n14879;
  assign n14883 = n1669 & n14882;
  assign n14884 = n2264 & n14881;
  assign n14885 = n13317 & n14877;
  assign n14886 = n14884 & n14885;
  assign n14887 = n4273 & n14883;
  assign n14888 = n14886 & n14887;
  assign n14889 = n6923 & n14888;
  assign n14890 = n749 & n1136;
  assign n14891 = ~n184 & ~n313;
  assign n14892 = n272 & n14891;
  assign n14893 = n1243 & n3007;
  assign n14894 = n12963 & n14893;
  assign n14895 = n717 & n14892;
  assign n14896 = n3632 & n5646;
  assign n14897 = n13629 & n14890;
  assign n14898 = n14896 & n14897;
  assign n14899 = n14894 & n14895;
  assign n14900 = n3649 & n14899;
  assign n14901 = n14898 & n14900;
  assign n14902 = ~n196 & ~n539;
  assign n14903 = n240 & n14902;
  assign n14904 = ~n148 & ~n174;
  assign n14905 = ~n215 & ~n334;
  assign n14906 = n14904 & n14905;
  assign n14907 = n160 & n1151;
  assign n14908 = n2757 & n3325;
  assign n14909 = n12852 & n14908;
  assign n14910 = n14906 & n14907;
  assign n14911 = n442 & n2196;
  assign n14912 = n14903 & n14911;
  assign n14913 = n14909 & n14910;
  assign n14914 = n3439 & n6846;
  assign n14915 = n14913 & n14914;
  assign n14916 = n13316 & n14912;
  assign n14917 = n14915 & n14916;
  assign n14918 = n14889 & n14917;
  assign n14919 = n14901 & n14918;
  assign n14920 = n3692 & n12476;
  assign n14921 = n12504 & ~n12506;
  assign n14922 = ~n12507 & ~n14921;
  assign n14923 = n880 & n14922;
  assign n14924 = n748 & n12479;
  assign n14925 = n3694 & n12473;
  assign n14926 = ~n14920 & ~n14924;
  assign n14927 = ~n14925 & n14926;
  assign n14928 = ~n14923 & n14927;
  assign n14929 = ~n14919 & ~n14928;
  assign n14930 = ~n374 & ~n377;
  assign n14931 = ~n414 & ~n753;
  assign n14932 = n14930 & n14931;
  assign n14933 = n1005 & n1429;
  assign n14934 = n1642 & n2040;
  assign n14935 = n2108 & n2658;
  assign n14936 = n3205 & n14935;
  assign n14937 = n14933 & n14934;
  assign n14938 = n517 & n14932;
  assign n14939 = n3722 & n14938;
  assign n14940 = n14936 & n14937;
  assign n14941 = n14939 & n14940;
  assign n14942 = n2217 & n14941;
  assign n14943 = n13664 & n14942;
  assign n14944 = ~n370 & ~n522;
  assign n14945 = ~n751 & n14944;
  assign n14946 = n254 & n417;
  assign n14947 = n933 & n1321;
  assign n14948 = n1779 & n2868;
  assign n14949 = n14947 & n14948;
  assign n14950 = n14945 & n14946;
  assign n14951 = n14949 & n14950;
  assign n14952 = n2594 & n14951;
  assign n14953 = n3743 & n14952;
  assign n14954 = n12745 & n14953;
  assign n14955 = n14943 & n14954;
  assign n14956 = n3692 & n12479;
  assign n14957 = n12500 & ~n12502;
  assign n14958 = ~n12503 & ~n14957;
  assign n14959 = n880 & n14958;
  assign n14960 = n748 & n12482;
  assign n14961 = n3694 & n12476;
  assign n14962 = ~n14956 & ~n14960;
  assign n14963 = ~n14961 & n14962;
  assign n14964 = ~n14959 & n14963;
  assign n14965 = ~n14955 & ~n14964;
  assign n14966 = ~n661 & n1722;
  assign n14967 = n12667 & n14966;
  assign n14968 = ~n243 & ~n309;
  assign n14969 = ~n894 & n14968;
  assign n14970 = n4269 & n14969;
  assign n14971 = n1030 & n14970;
  assign n14972 = ~n236 & ~n255;
  assign n14973 = ~n283 & ~n365;
  assign n14974 = ~n535 & ~n638;
  assign n14975 = ~n653 & ~n937;
  assign n14976 = n14974 & n14975;
  assign n14977 = n14972 & n14973;
  assign n14978 = n1430 & n14977;
  assign n14979 = n418 & n14976;
  assign n14980 = n3822 & n14979;
  assign n14981 = n14967 & n14978;
  assign n14982 = n14980 & n14981;
  assign n14983 = n13582 & n14971;
  assign n14984 = n14982 & n14983;
  assign n14985 = ~n247 & ~n259;
  assign n14986 = ~n437 & ~n502;
  assign n14987 = ~n810 & n14986;
  assign n14988 = n413 & n14985;
  assign n14989 = n660 & n759;
  assign n14990 = n2548 & n14989;
  assign n14991 = n14987 & n14988;
  assign n14992 = n2001 & n14991;
  assign n14993 = n1583 & n14990;
  assign n14994 = n5290 & n14993;
  assign n14995 = n14992 & n14994;
  assign n14996 = n3045 & n14995;
  assign n14997 = n14984 & n14996;
  assign n14998 = n234 & n14997;
  assign n14999 = n3692 & n12482;
  assign n15000 = n12496 & ~n12498;
  assign n15001 = ~n12499 & ~n15000;
  assign n15002 = n880 & n15001;
  assign n15003 = n748 & n12485;
  assign n15004 = n3694 & n12479;
  assign n15005 = ~n14999 & ~n15003;
  assign n15006 = ~n15004 & n15005;
  assign n15007 = ~n15002 & n15006;
  assign n15008 = ~n14998 & ~n15007;
  assign n15009 = ~n155 & ~n246;
  assign n15010 = ~n564 & ~n648;
  assign n15011 = ~n922 & n15010;
  assign n15012 = n657 & n15009;
  assign n15013 = n1351 & n1663;
  assign n15014 = n4326 & n15013;
  assign n15015 = n15011 & n15012;
  assign n15016 = n15014 & n15015;
  assign n15017 = n930 & n3346;
  assign n15018 = n6888 & n15017;
  assign n15019 = n5751 & n15016;
  assign n15020 = n15018 & n15019;
  assign n15021 = n624 & n3930;
  assign n15022 = n15020 & n15021;
  assign n15023 = n4324 & n15022;
  assign n15024 = n3692 & n12485;
  assign n15025 = ~n12488 & ~n12494;
  assign n15026 = ~n12495 & ~n15025;
  assign n15027 = n880 & n15026;
  assign n15028 = n748 & n12490;
  assign n15029 = n3694 & n12482;
  assign n15030 = ~n15024 & ~n15028;
  assign n15031 = ~n15029 & n15030;
  assign n15032 = ~n15027 & n15031;
  assign n15033 = ~n15023 & ~n15032;
  assign n15034 = ~n15023 & n15032;
  assign n15035 = n15023 & ~n15032;
  assign n15036 = ~n15034 & ~n15035;
  assign n15037 = ~n123 & ~n380;
  assign n15038 = ~n361 & ~n536;
  assign n15039 = ~n596 & n15038;
  assign n15040 = n664 & n15037;
  assign n15041 = n15039 & n15040;
  assign n15042 = n2036 & n15041;
  assign n15043 = ~n196 & ~n213;
  assign n15044 = ~n477 & ~n1032;
  assign n15045 = n15043 & n15044;
  assign n15046 = n647 & n1049;
  assign n15047 = n1122 & n1188;
  assign n15048 = n15046 & n15047;
  assign n15049 = n3661 & n15045;
  assign n15050 = n15048 & n15049;
  assign n15051 = n571 & n916;
  assign n15052 = n14860 & n15051;
  assign n15053 = n15042 & n15050;
  assign n15054 = n15052 & n15053;
  assign n15055 = ~n199 & ~n689;
  assign n15056 = ~n937 & n15055;
  assign n15057 = n487 & n540;
  assign n15058 = n1915 & n2309;
  assign n15059 = n15057 & n15058;
  assign n15060 = n15056 & n15059;
  assign n15061 = n844 & n2854;
  assign n15062 = n2874 & n2936;
  assign n15063 = n15061 & n15062;
  assign n15064 = n15060 & n15063;
  assign n15065 = n6982 & n15064;
  assign n15066 = n15054 & n15065;
  assign n15067 = n3148 & n15066;
  assign n15068 = n3694 & n12490;
  assign n15069 = n3692 & n12492;
  assign n15070 = n12490 & ~n12492;
  assign n15071 = ~n12490 & n12492;
  assign n15072 = ~n15070 & ~n15071;
  assign n15073 = n880 & ~n15072;
  assign n15074 = ~n15068 & ~n15069;
  assign n15075 = ~n15073 & n15074;
  assign n15076 = ~n15067 & ~n15075;
  assign n15077 = n1779 & n1884;
  assign n15078 = ~n515 & ~n648;
  assign n15079 = ~n1699 & n15078;
  assign n15080 = ~n163 & ~n314;
  assign n15081 = ~n353 & ~n509;
  assign n15082 = ~n814 & n15081;
  assign n15083 = n895 & n15080;
  assign n15084 = n2024 & n2309;
  assign n15085 = n15083 & n15084;
  assign n15086 = n1721 & n15082;
  assign n15087 = n15077 & n15079;
  assign n15088 = n15086 & n15087;
  assign n15089 = n15085 & n15088;
  assign n15090 = ~n136 & ~n153;
  assign n15091 = ~n155 & ~n199;
  assign n15092 = ~n281 & ~n304;
  assign n15093 = ~n526 & ~n689;
  assign n15094 = ~n1051 & n15093;
  assign n15095 = n15091 & n15092;
  assign n15096 = n479 & n15090;
  assign n15097 = n883 & n1673;
  assign n15098 = n2207 & n15097;
  assign n15099 = n15095 & n15096;
  assign n15100 = n1379 & n15094;
  assign n15101 = n3707 & n3936;
  assign n15102 = n15100 & n15101;
  assign n15103 = n15098 & n15099;
  assign n15104 = n15102 & n15103;
  assign n15105 = n14378 & n15104;
  assign n15106 = n15089 & n15105;
  assign n15107 = n13603 & n15106;
  assign n15108 = n15076 & ~n15107;
  assign n15109 = ~n15076 & n15107;
  assign n15110 = n748 & n12492;
  assign n15111 = n12485 & ~n15070;
  assign n15112 = ~n12485 & n15070;
  assign n15113 = ~n15111 & ~n15112;
  assign n15114 = n880 & ~n15113;
  assign n15115 = n3692 & n12490;
  assign n15116 = n3694 & n12485;
  assign n15117 = ~n15110 & ~n15115;
  assign n15118 = ~n15116 & n15117;
  assign n15119 = ~n15114 & n15118;
  assign n15120 = ~n15109 & ~n15119;
  assign n15121 = ~n15108 & ~n15120;
  assign n15122 = ~n15036 & ~n15121;
  assign n15123 = ~n15033 & ~n15122;
  assign n15124 = ~n14998 & n15007;
  assign n15125 = n14998 & ~n15007;
  assign n15126 = ~n15124 & ~n15125;
  assign n15127 = ~n15123 & ~n15126;
  assign n15128 = ~n15008 & ~n15127;
  assign n15129 = ~n14955 & n14964;
  assign n15130 = n14955 & ~n14964;
  assign n15131 = ~n15129 & ~n15130;
  assign n15132 = ~n15128 & ~n15131;
  assign n15133 = ~n14965 & ~n15132;
  assign n15134 = ~n14919 & n14928;
  assign n15135 = n14919 & ~n14928;
  assign n15136 = ~n15134 & ~n15135;
  assign n15137 = ~n15133 & ~n15136;
  assign n15138 = ~n14929 & ~n15137;
  assign n15139 = n14855 & ~n14874;
  assign n15140 = ~n14855 & n14874;
  assign n15141 = ~n15139 & ~n15140;
  assign n15142 = ~n15138 & ~n15141;
  assign n15143 = ~n14875 & ~n15142;
  assign n15144 = ~n14836 & n14845;
  assign n15145 = n14836 & ~n14845;
  assign n15146 = ~n15144 & ~n15145;
  assign n15147 = ~n15143 & ~n15146;
  assign n15148 = ~n14846 & ~n15147;
  assign n15149 = ~n14812 & n14821;
  assign n15150 = n14812 & ~n14821;
  assign n15151 = ~n15149 & ~n15150;
  assign n15152 = ~n15148 & ~n15151;
  assign n15153 = ~n14822 & ~n15152;
  assign n15154 = ~n14786 & n14795;
  assign n15155 = n14786 & ~n14795;
  assign n15156 = ~n15154 & ~n15155;
  assign n15157 = ~n15153 & ~n15156;
  assign n15158 = ~n14796 & ~n15157;
  assign n15159 = ~n14416 & ~n14417;
  assign n15160 = ~n14426 & n15159;
  assign n15161 = n14426 & ~n15159;
  assign n15162 = ~n15160 & ~n15161;
  assign n15163 = ~n15158 & n15162;
  assign n15164 = n15158 & ~n15162;
  assign n15165 = ~n15163 & ~n15164;
  assign n15166 = n3810 & n12455;
  assign n15167 = n3886 & n14442;
  assign n15168 = n3884 & n12452;
  assign n15169 = n4380 & n12449;
  assign n15170 = ~n15166 & ~n15168;
  assign n15171 = ~n15169 & n15170;
  assign n15172 = ~n15167 & n15171;
  assign n15173 = pi29  & n15172;
  assign n15174 = ~pi29  & ~n15172;
  assign n15175 = ~n15173 & ~n15174;
  assign n15176 = n15165 & ~n15175;
  assign n15177 = ~n15163 & ~n15176;
  assign n15178 = ~n14766 & ~n15177;
  assign n15179 = ~n14763 & ~n15178;
  assign n15180 = ~n14751 & ~n15179;
  assign n15181 = ~n14748 & ~n15180;
  assign n15182 = ~n14439 & n14448;
  assign n15183 = ~n14449 & ~n15182;
  assign n15184 = ~n15181 & n15183;
  assign n15185 = n15181 & ~n15183;
  assign n15186 = n3810 & n12446;
  assign n15187 = n3886 & n14175;
  assign n15188 = n3884 & n12443;
  assign n15189 = n4380 & n12440;
  assign n15190 = ~n15186 & ~n15188;
  assign n15191 = ~n15189 & n15190;
  assign n15192 = ~n15187 & n15191;
  assign n15193 = pi29  & n15192;
  assign n15194 = ~pi29  & ~n15192;
  assign n15195 = ~n15193 & ~n15194;
  assign n15196 = ~n15185 & ~n15195;
  assign n15197 = ~n15184 & ~n15196;
  assign n15198 = n14736 & ~n15197;
  assign n15199 = ~n14736 & n15197;
  assign n15200 = n86 & n12434;
  assign n15201 = n4420 & n13546;
  assign n15202 = n4600 & n12431;
  assign n15203 = n4615 & n12428;
  assign n15204 = ~n15200 & ~n15202;
  assign n15205 = ~n15203 & n15204;
  assign n15206 = ~n15201 & n15205;
  assign n15207 = pi26  & n15206;
  assign n15208 = ~pi26  & ~n15206;
  assign n15209 = ~n15207 & ~n15208;
  assign n15210 = ~n15199 & ~n15209;
  assign n15211 = ~n15198 & ~n15210;
  assign n15212 = ~n14734 & ~n15211;
  assign n15213 = n14734 & n15211;
  assign n15214 = n5044 & n12422;
  assign n15215 = n5045 & n13201;
  assign n15216 = n5109 & n12419;
  assign n15217 = n5130 & n12416;
  assign n15218 = ~n15214 & ~n15216;
  assign n15219 = ~n15217 & n15218;
  assign n15220 = ~n15215 & n15219;
  assign n15221 = pi23  & n15220;
  assign n15222 = ~pi23  & ~n15220;
  assign n15223 = ~n15221 & ~n15222;
  assign n15224 = ~n15213 & ~n15223;
  assign n15225 = ~n15212 & ~n15224;
  assign n15226 = ~n14731 & ~n15225;
  assign n15227 = ~n14728 & ~n15226;
  assign n15228 = ~n14635 & ~n14636;
  assign n15229 = ~n14646 & n15228;
  assign n15230 = n14646 & ~n15228;
  assign n15231 = ~n15229 & ~n15230;
  assign n15232 = ~n15227 & n15231;
  assign n15233 = n15227 & ~n15231;
  assign n15234 = n5240 & n12407;
  assign n15235 = n5241 & n13035;
  assign n15236 = n5853 & n12404;
  assign n15237 = n5866 & n12401;
  assign n15238 = ~n15234 & ~n15236;
  assign n15239 = ~n15237 & n15238;
  assign n15240 = ~n15235 & n15239;
  assign n15241 = pi20  & n15240;
  assign n15242 = ~pi20  & ~n15240;
  assign n15243 = ~n15241 & ~n15242;
  assign n15244 = ~n15233 & ~n15243;
  assign n15245 = ~n15232 & ~n15244;
  assign n15246 = n14715 & ~n15245;
  assign n15247 = ~n14715 & n15245;
  assign n15248 = n5982 & n12395;
  assign n15249 = n5983 & n13144;
  assign n15250 = n6323 & n12362;
  assign n15251 = n6336 & n12392;
  assign n15252 = ~n15248 & ~n15250;
  assign n15253 = ~n15251 & n15252;
  assign n15254 = ~n15249 & n15253;
  assign n15255 = pi17  & n15254;
  assign n15256 = ~pi17  & ~n15254;
  assign n15257 = ~n15255 & ~n15256;
  assign n15258 = ~n15247 & ~n15257;
  assign n15259 = ~n15246 & ~n15258;
  assign n15260 = ~n14711 & ~n15259;
  assign n15261 = ~n14708 & ~n15260;
  assign n15262 = ~n14669 & ~n14670;
  assign n15263 = ~n14680 & n15262;
  assign n15264 = n14680 & ~n15262;
  assign n15265 = ~n15263 & ~n15264;
  assign n15266 = ~n15261 & n15265;
  assign n15267 = n15261 & ~n15265;
  assign n15268 = n7262 & ~n12786;
  assign n15269 = n6631 & ~n13781;
  assign n15270 = n6630 & n13166;
  assign n15271 = n7238 & n13161;
  assign n15272 = ~n15268 & ~n15270;
  assign n15273 = ~n15271 & n15272;
  assign n15274 = ~n15269 & n15273;
  assign n15275 = pi14  & n15274;
  assign n15276 = ~pi14  & ~n15274;
  assign n15277 = ~n15275 & ~n15276;
  assign n15278 = ~n15267 & ~n15277;
  assign n15279 = ~n15266 & ~n15278;
  assign n15280 = n14695 & ~n15279;
  assign n15281 = ~n14695 & n15279;
  assign n15282 = ~n15280 & ~n15281;
  assign n15283 = n7262 & n13161;
  assign n15284 = n6631 & n13183;
  assign n15285 = n7238 & n13166;
  assign n15286 = n6630 & n13164;
  assign n15287 = ~n15285 & ~n15286;
  assign n15288 = ~n15283 & n15287;
  assign n15289 = ~n15284 & n15288;
  assign n15290 = pi14  & n15289;
  assign n15291 = ~pi14  & ~n15289;
  assign n15292 = ~n15290 & ~n15291;
  assign n15293 = ~n15246 & ~n15247;
  assign n15294 = ~n15257 & n15293;
  assign n15295 = n15257 & ~n15293;
  assign n15296 = ~n15294 & ~n15295;
  assign n15297 = n14731 & n15225;
  assign n15298 = ~n15226 & ~n15297;
  assign n15299 = n5240 & n12410;
  assign n15300 = n5241 & n13093;
  assign n15301 = n5853 & n12407;
  assign n15302 = n5866 & n12404;
  assign n15303 = ~n15299 & ~n15301;
  assign n15304 = ~n15302 & n15303;
  assign n15305 = ~n15300 & n15304;
  assign n15306 = pi20  & n15305;
  assign n15307 = ~pi20  & ~n15305;
  assign n15308 = ~n15306 & ~n15307;
  assign n15309 = n15298 & ~n15308;
  assign n15310 = n15298 & n15308;
  assign n15311 = ~n15298 & ~n15308;
  assign n15312 = ~n15310 & ~n15311;
  assign n15313 = ~n15212 & ~n15213;
  assign n15314 = ~n15223 & n15313;
  assign n15315 = n15223 & ~n15313;
  assign n15316 = ~n15314 & ~n15315;
  assign n15317 = n86 & n12437;
  assign n15318 = n4420 & n13564;
  assign n15319 = n4600 & n12434;
  assign n15320 = n4615 & n12431;
  assign n15321 = ~n15317 & ~n15319;
  assign n15322 = ~n15320 & n15321;
  assign n15323 = ~n15318 & n15322;
  assign n15324 = pi26  & n15323;
  assign n15325 = ~pi26  & ~n15323;
  assign n15326 = ~n15324 & ~n15325;
  assign n15327 = ~n15184 & ~n15185;
  assign n15328 = ~n15195 & n15327;
  assign n15329 = n15195 & ~n15327;
  assign n15330 = ~n15328 & ~n15329;
  assign n15331 = ~n15326 & n15330;
  assign n15332 = n14751 & n15179;
  assign n15333 = ~n15180 & ~n15332;
  assign n15334 = n3810 & n12449;
  assign n15335 = n3886 & n14325;
  assign n15336 = n3884 & n12446;
  assign n15337 = n4380 & n12443;
  assign n15338 = ~n15334 & ~n15336;
  assign n15339 = ~n15337 & n15338;
  assign n15340 = ~n15335 & n15339;
  assign n15341 = pi29  & n15340;
  assign n15342 = ~pi29  & ~n15340;
  assign n15343 = ~n15341 & ~n15342;
  assign n15344 = n15333 & ~n15343;
  assign n15345 = n15333 & n15343;
  assign n15346 = ~n15333 & ~n15343;
  assign n15347 = ~n15345 & ~n15346;
  assign n15348 = n86 & n12440;
  assign n15349 = n4420 & n13939;
  assign n15350 = n4600 & n12437;
  assign n15351 = n4615 & n12434;
  assign n15352 = ~n15348 & ~n15350;
  assign n15353 = ~n15351 & n15352;
  assign n15354 = ~n15349 & n15353;
  assign n15355 = pi26  & n15354;
  assign n15356 = ~pi26  & ~n15354;
  assign n15357 = ~n15355 & ~n15356;
  assign n15358 = ~n15347 & ~n15357;
  assign n15359 = ~n15344 & ~n15358;
  assign n15360 = n15326 & ~n15330;
  assign n15361 = ~n15331 & ~n15360;
  assign n15362 = ~n15359 & n15361;
  assign n15363 = ~n15331 & ~n15362;
  assign n15364 = ~n15198 & ~n15199;
  assign n15365 = ~n15209 & n15364;
  assign n15366 = n15209 & ~n15364;
  assign n15367 = ~n15365 & ~n15366;
  assign n15368 = ~n15363 & n15367;
  assign n15369 = n15363 & ~n15367;
  assign n15370 = n5044 & n12425;
  assign n15371 = n5045 & n13010;
  assign n15372 = n5109 & n12422;
  assign n15373 = n5130 & n12419;
  assign n15374 = ~n15370 & ~n15372;
  assign n15375 = ~n15373 & n15374;
  assign n15376 = ~n15371 & n15375;
  assign n15377 = pi23  & n15376;
  assign n15378 = ~pi23  & ~n15376;
  assign n15379 = ~n15377 & ~n15378;
  assign n15380 = ~n15369 & ~n15379;
  assign n15381 = ~n15368 & ~n15380;
  assign n15382 = n15316 & ~n15381;
  assign n15383 = ~n15316 & n15381;
  assign n15384 = n5240 & n12413;
  assign n15385 = n5241 & n12891;
  assign n15386 = n5853 & n12410;
  assign n15387 = n5866 & n12407;
  assign n15388 = ~n15384 & ~n15386;
  assign n15389 = ~n15387 & n15388;
  assign n15390 = ~n15385 & n15389;
  assign n15391 = pi20  & n15390;
  assign n15392 = ~pi20  & ~n15390;
  assign n15393 = ~n15391 & ~n15392;
  assign n15394 = ~n15383 & ~n15393;
  assign n15395 = ~n15382 & ~n15394;
  assign n15396 = ~n15312 & ~n15395;
  assign n15397 = ~n15309 & ~n15396;
  assign n15398 = ~n15232 & ~n15233;
  assign n15399 = ~n15243 & n15398;
  assign n15400 = n15243 & ~n15398;
  assign n15401 = ~n15399 & ~n15400;
  assign n15402 = ~n15397 & n15401;
  assign n15403 = n15397 & ~n15401;
  assign n15404 = n5982 & n12398;
  assign n15405 = n5983 & n13245;
  assign n15406 = n6323 & n12395;
  assign n15407 = n6336 & n12362;
  assign n15408 = ~n15404 & ~n15406;
  assign n15409 = ~n15407 & n15408;
  assign n15410 = ~n15405 & n15409;
  assign n15411 = pi17  & n15410;
  assign n15412 = ~pi17  & ~n15410;
  assign n15413 = ~n15411 & ~n15412;
  assign n15414 = ~n15403 & ~n15413;
  assign n15415 = ~n15402 & ~n15414;
  assign n15416 = n15296 & ~n15415;
  assign n15417 = ~n15296 & n15415;
  assign n15418 = n6630 & n12646;
  assign n15419 = n6631 & n13261;
  assign n15420 = n7238 & n13164;
  assign n15421 = n7262 & n13166;
  assign n15422 = ~n15418 & ~n15420;
  assign n15423 = ~n15421 & n15422;
  assign n15424 = ~n15419 & n15423;
  assign n15425 = pi14  & n15424;
  assign n15426 = ~pi14  & ~n15424;
  assign n15427 = ~n15425 & ~n15426;
  assign n15428 = ~n15417 & ~n15427;
  assign n15429 = ~n15416 & ~n15428;
  assign n15430 = ~n15292 & ~n15429;
  assign n15431 = n14711 & n15259;
  assign n15432 = ~n15260 & ~n15431;
  assign n15433 = n15292 & ~n15429;
  assign n15434 = ~n15292 & n15429;
  assign n15435 = ~n15433 & ~n15434;
  assign n15436 = n15432 & ~n15435;
  assign n15437 = ~n15430 & ~n15436;
  assign n15438 = ~n15266 & ~n15267;
  assign n15439 = ~n15277 & n15438;
  assign n15440 = n15277 & ~n15438;
  assign n15441 = ~n15439 & ~n15440;
  assign n15442 = ~n15437 & n15441;
  assign n15443 = n15437 & n15441;
  assign n15444 = ~n15437 & ~n15441;
  assign n15445 = ~n15443 & ~n15444;
  assign n15446 = ~n15432 & n15435;
  assign n15447 = ~n15436 & ~n15446;
  assign n15448 = n7431 & ~n13280;
  assign n15449 = n7430 & ~n13160;
  assign n15450 = ~n7869 & ~n7895;
  assign n15451 = ~n15449 & n15450;
  assign n15452 = ~n12786 & ~n15451;
  assign n15453 = ~n15448 & ~n15452;
  assign n15454 = pi11  & n15453;
  assign n15455 = ~pi11  & ~n15453;
  assign n15456 = ~n15454 & ~n15455;
  assign n15457 = n15312 & n15395;
  assign n15458 = ~n15396 & ~n15457;
  assign n15459 = n5982 & n12401;
  assign n15460 = n5983 & n13108;
  assign n15461 = n6323 & n12398;
  assign n15462 = n6336 & n12395;
  assign n15463 = ~n15459 & ~n15461;
  assign n15464 = ~n15462 & n15463;
  assign n15465 = ~n15460 & n15464;
  assign n15466 = pi17  & n15465;
  assign n15467 = ~pi17  & ~n15465;
  assign n15468 = ~n15466 & ~n15467;
  assign n15469 = n15458 & ~n15468;
  assign n15470 = n15458 & n15468;
  assign n15471 = ~n15458 & ~n15468;
  assign n15472 = ~n15470 & ~n15471;
  assign n15473 = ~n15382 & ~n15383;
  assign n15474 = ~n15393 & n15473;
  assign n15475 = n15393 & ~n15473;
  assign n15476 = ~n15474 & ~n15475;
  assign n15477 = n15359 & ~n15361;
  assign n15478 = ~n15362 & ~n15477;
  assign n15479 = n5044 & n12428;
  assign n15480 = n5045 & n13371;
  assign n15481 = n5109 & n12425;
  assign n15482 = n5130 & n12422;
  assign n15483 = ~n15479 & ~n15481;
  assign n15484 = ~n15482 & n15483;
  assign n15485 = ~n15480 & n15484;
  assign n15486 = pi23  & n15485;
  assign n15487 = ~pi23  & ~n15485;
  assign n15488 = ~n15486 & ~n15487;
  assign n15489 = n15478 & ~n15488;
  assign n15490 = n15478 & n15488;
  assign n15491 = ~n15478 & ~n15488;
  assign n15492 = ~n15490 & ~n15491;
  assign n15493 = ~n15347 & n15357;
  assign n15494 = n15347 & ~n15357;
  assign n15495 = ~n15493 & ~n15494;
  assign n15496 = n14766 & n15177;
  assign n15497 = ~n15178 & ~n15496;
  assign n15498 = n3810 & n12452;
  assign n15499 = n3886 & n14156;
  assign n15500 = n3884 & n12449;
  assign n15501 = n4380 & n12446;
  assign n15502 = ~n15498 & ~n15500;
  assign n15503 = ~n15501 & n15502;
  assign n15504 = ~n15499 & n15503;
  assign n15505 = pi29  & n15504;
  assign n15506 = ~pi29  & ~n15504;
  assign n15507 = ~n15505 & ~n15506;
  assign n15508 = n15497 & ~n15507;
  assign n15509 = n15497 & n15507;
  assign n15510 = ~n15497 & ~n15507;
  assign n15511 = ~n15509 & ~n15510;
  assign n15512 = n4600 & n12440;
  assign n15513 = n4420 & n13702;
  assign n15514 = n86 & n12443;
  assign n15515 = n4615 & n12437;
  assign n15516 = ~n15512 & ~n15514;
  assign n15517 = ~n15515 & n15516;
  assign n15518 = ~n15513 & n15517;
  assign n15519 = pi26  & n15518;
  assign n15520 = ~pi26  & ~n15518;
  assign n15521 = ~n15519 & ~n15520;
  assign n15522 = ~n15511 & ~n15521;
  assign n15523 = ~n15508 & ~n15522;
  assign n15524 = ~n15495 & ~n15523;
  assign n15525 = n15495 & n15523;
  assign n15526 = n5044 & n12431;
  assign n15527 = n5045 & n13356;
  assign n15528 = n5109 & n12428;
  assign n15529 = n5130 & n12425;
  assign n15530 = ~n15526 & ~n15528;
  assign n15531 = ~n15529 & n15530;
  assign n15532 = ~n15527 & n15531;
  assign n15533 = pi23  & n15532;
  assign n15534 = ~pi23  & ~n15532;
  assign n15535 = ~n15533 & ~n15534;
  assign n15536 = ~n15525 & ~n15535;
  assign n15537 = ~n15524 & ~n15536;
  assign n15538 = ~n15492 & ~n15537;
  assign n15539 = ~n15489 & ~n15538;
  assign n15540 = ~n15368 & ~n15369;
  assign n15541 = ~n15379 & n15540;
  assign n15542 = n15379 & ~n15540;
  assign n15543 = ~n15541 & ~n15542;
  assign n15544 = ~n15539 & n15543;
  assign n15545 = n15539 & ~n15543;
  assign n15546 = n5240 & n12416;
  assign n15547 = n5241 & n12843;
  assign n15548 = n5853 & n12413;
  assign n15549 = n5866 & n12410;
  assign n15550 = ~n15546 & ~n15548;
  assign n15551 = ~n15549 & n15550;
  assign n15552 = ~n15547 & n15551;
  assign n15553 = pi20  & n15552;
  assign n15554 = ~pi20  & ~n15552;
  assign n15555 = ~n15553 & ~n15554;
  assign n15556 = ~n15545 & ~n15555;
  assign n15557 = ~n15544 & ~n15556;
  assign n15558 = n15476 & ~n15557;
  assign n15559 = ~n15476 & n15557;
  assign n15560 = n5982 & n12404;
  assign n15561 = n5983 & n13128;
  assign n15562 = n6323 & n12401;
  assign n15563 = n6336 & n12398;
  assign n15564 = ~n15560 & ~n15562;
  assign n15565 = ~n15563 & n15564;
  assign n15566 = ~n15561 & n15565;
  assign n15567 = pi17  & n15566;
  assign n15568 = ~pi17  & ~n15566;
  assign n15569 = ~n15567 & ~n15568;
  assign n15570 = ~n15559 & ~n15569;
  assign n15571 = ~n15558 & ~n15570;
  assign n15572 = ~n15472 & ~n15571;
  assign n15573 = ~n15469 & ~n15572;
  assign n15574 = ~n15402 & ~n15403;
  assign n15575 = ~n15413 & n15574;
  assign n15576 = n15413 & ~n15574;
  assign n15577 = ~n15575 & ~n15576;
  assign n15578 = ~n15573 & n15577;
  assign n15579 = n15573 & ~n15577;
  assign n15580 = n6630 & n12392;
  assign n15581 = n6631 & n13421;
  assign n15582 = n7238 & n12646;
  assign n15583 = n7262 & n13164;
  assign n15584 = ~n15580 & ~n15582;
  assign n15585 = ~n15583 & n15584;
  assign n15586 = ~n15581 & n15585;
  assign n15587 = pi14  & n15586;
  assign n15588 = ~pi14  & ~n15586;
  assign n15589 = ~n15587 & ~n15588;
  assign n15590 = ~n15579 & ~n15589;
  assign n15591 = ~n15578 & ~n15590;
  assign n15592 = ~n15456 & ~n15591;
  assign n15593 = n15456 & n15591;
  assign n15594 = ~n15416 & ~n15417;
  assign n15595 = ~n15427 & n15594;
  assign n15596 = n15427 & ~n15594;
  assign n15597 = ~n15595 & ~n15596;
  assign n15598 = ~n15593 & n15597;
  assign n15599 = ~n15592 & ~n15598;
  assign n15600 = n15447 & ~n15599;
  assign n15601 = ~n15592 & ~n15593;
  assign n15602 = n15597 & n15601;
  assign n15603 = ~n15597 & ~n15601;
  assign n15604 = ~n15602 & ~n15603;
  assign n15605 = n15472 & n15571;
  assign n15606 = ~n15572 & ~n15605;
  assign n15607 = n6630 & n12362;
  assign n15608 = n6631 & n12652;
  assign n15609 = n7238 & n12392;
  assign n15610 = n7262 & n12646;
  assign n15611 = ~n15607 & ~n15609;
  assign n15612 = ~n15610 & n15611;
  assign n15613 = ~n15608 & n15612;
  assign n15614 = pi14  & n15613;
  assign n15615 = ~pi14  & ~n15613;
  assign n15616 = ~n15614 & ~n15615;
  assign n15617 = n15606 & ~n15616;
  assign n15618 = n15606 & n15616;
  assign n15619 = ~n15606 & ~n15616;
  assign n15620 = ~n15618 & ~n15619;
  assign n15621 = ~n15558 & ~n15559;
  assign n15622 = ~n15569 & n15621;
  assign n15623 = n15569 & ~n15621;
  assign n15624 = ~n15622 & ~n15623;
  assign n15625 = n15492 & n15537;
  assign n15626 = ~n15538 & ~n15625;
  assign n15627 = n5240 & n12419;
  assign n15628 = n5241 & n12908;
  assign n15629 = n5853 & n12416;
  assign n15630 = n5866 & n12413;
  assign n15631 = ~n15627 & ~n15629;
  assign n15632 = ~n15630 & n15631;
  assign n15633 = ~n15628 & n15632;
  assign n15634 = pi20  & n15633;
  assign n15635 = ~pi20  & ~n15633;
  assign n15636 = ~n15634 & ~n15635;
  assign n15637 = n15626 & ~n15636;
  assign n15638 = n15626 & n15636;
  assign n15639 = ~n15626 & ~n15636;
  assign n15640 = ~n15638 & ~n15639;
  assign n15641 = ~n15524 & ~n15525;
  assign n15642 = ~n15535 & n15641;
  assign n15643 = n15535 & ~n15641;
  assign n15644 = ~n15642 & ~n15643;
  assign n15645 = ~n15511 & n15521;
  assign n15646 = n15511 & ~n15521;
  assign n15647 = ~n15645 & ~n15646;
  assign n15648 = n3810 & n12458;
  assign n15649 = n3886 & n14741;
  assign n15650 = n3884 & n12455;
  assign n15651 = n4380 & n12452;
  assign n15652 = ~n15648 & ~n15650;
  assign n15653 = ~n15651 & n15652;
  assign n15654 = ~n15649 & n15653;
  assign n15655 = pi29  & n15654;
  assign n15656 = ~pi29  & ~n15654;
  assign n15657 = ~n15655 & ~n15656;
  assign n15658 = n15153 & n15156;
  assign n15659 = ~n15157 & ~n15658;
  assign n15660 = ~n15657 & n15659;
  assign n15661 = n3810 & n12461;
  assign n15662 = n3886 & n14756;
  assign n15663 = n3884 & n12458;
  assign n15664 = n4380 & n12455;
  assign n15665 = ~n15661 & ~n15663;
  assign n15666 = ~n15664 & n15665;
  assign n15667 = ~n15662 & n15666;
  assign n15668 = pi29  & n15667;
  assign n15669 = ~pi29  & ~n15667;
  assign n15670 = ~n15668 & ~n15669;
  assign n15671 = n15148 & n15151;
  assign n15672 = ~n15152 & ~n15671;
  assign n15673 = ~n15670 & n15672;
  assign n15674 = n3810 & n12464;
  assign n15675 = n3886 & n14420;
  assign n15676 = n3884 & n12461;
  assign n15677 = n4380 & n12458;
  assign n15678 = ~n15674 & ~n15676;
  assign n15679 = ~n15677 & n15678;
  assign n15680 = ~n15675 & n15679;
  assign n15681 = pi29  & n15680;
  assign n15682 = ~pi29  & ~n15680;
  assign n15683 = ~n15681 & ~n15682;
  assign n15684 = n15143 & n15146;
  assign n15685 = ~n15147 & ~n15684;
  assign n15686 = ~n15683 & n15685;
  assign n15687 = n3810 & n12467;
  assign n15688 = n3886 & n14789;
  assign n15689 = n3884 & n12464;
  assign n15690 = n4380 & n12461;
  assign n15691 = ~n15687 & ~n15689;
  assign n15692 = ~n15690 & n15691;
  assign n15693 = ~n15688 & n15692;
  assign n15694 = pi29  & n15693;
  assign n15695 = ~pi29  & ~n15693;
  assign n15696 = ~n15694 & ~n15695;
  assign n15697 = n15138 & n15141;
  assign n15698 = ~n15142 & ~n15697;
  assign n15699 = ~n15696 & n15698;
  assign n15700 = n3810 & n12470;
  assign n15701 = n3886 & n14815;
  assign n15702 = n3884 & n12467;
  assign n15703 = n4380 & n12464;
  assign n15704 = ~n15700 & ~n15702;
  assign n15705 = ~n15703 & n15704;
  assign n15706 = ~n15701 & n15705;
  assign n15707 = pi29  & n15706;
  assign n15708 = ~pi29  & ~n15706;
  assign n15709 = ~n15707 & ~n15708;
  assign n15710 = n15133 & n15136;
  assign n15711 = ~n15137 & ~n15710;
  assign n15712 = ~n15709 & n15711;
  assign n15713 = n3810 & n12473;
  assign n15714 = n3886 & n14839;
  assign n15715 = n3884 & n12470;
  assign n15716 = n4380 & n12467;
  assign n15717 = ~n15713 & ~n15715;
  assign n15718 = ~n15716 & n15717;
  assign n15719 = ~n15714 & n15718;
  assign n15720 = ~pi29  & ~n15719;
  assign n15721 = pi29  & n15719;
  assign n15722 = ~n15720 & ~n15721;
  assign n15723 = n15128 & n15131;
  assign n15724 = ~n15132 & ~n15723;
  assign n15725 = ~n15722 & n15724;
  assign n15726 = ~n15722 & ~n15724;
  assign n15727 = n15722 & n15724;
  assign n15728 = ~n15726 & ~n15727;
  assign n15729 = n3810 & n12476;
  assign n15730 = n3886 & n14849;
  assign n15731 = n3884 & n12473;
  assign n15732 = n4380 & n12470;
  assign n15733 = ~n15729 & ~n15731;
  assign n15734 = ~n15732 & n15733;
  assign n15735 = ~n15730 & n15734;
  assign n15736 = ~pi29  & ~n15735;
  assign n15737 = pi29  & n15735;
  assign n15738 = ~n15736 & ~n15737;
  assign n15739 = n15123 & n15126;
  assign n15740 = ~n15127 & ~n15739;
  assign n15741 = ~n15738 & n15740;
  assign n15742 = ~n15738 & ~n15740;
  assign n15743 = n15738 & n15740;
  assign n15744 = ~n15742 & ~n15743;
  assign n15745 = n3810 & n12479;
  assign n15746 = n3886 & n14922;
  assign n15747 = n3884 & n12476;
  assign n15748 = n4380 & n12473;
  assign n15749 = ~n15745 & ~n15747;
  assign n15750 = ~n15748 & n15749;
  assign n15751 = ~n15746 & n15750;
  assign n15752 = ~pi29  & ~n15751;
  assign n15753 = pi29  & n15751;
  assign n15754 = ~n15752 & ~n15753;
  assign n15755 = n15036 & n15121;
  assign n15756 = ~n15122 & ~n15755;
  assign n15757 = ~n15754 & n15756;
  assign n15758 = ~n15754 & ~n15756;
  assign n15759 = n15754 & n15756;
  assign n15760 = ~n15758 & ~n15759;
  assign n15761 = n3810 & n12482;
  assign n15762 = n3886 & n14958;
  assign n15763 = n3884 & n12479;
  assign n15764 = n4380 & n12476;
  assign n15765 = ~n15761 & ~n15763;
  assign n15766 = ~n15764 & n15765;
  assign n15767 = ~n15762 & n15766;
  assign n15768 = ~pi29  & ~n15767;
  assign n15769 = pi29  & n15767;
  assign n15770 = ~n15768 & ~n15769;
  assign n15771 = ~n15108 & ~n15109;
  assign n15772 = ~n15119 & n15771;
  assign n15773 = n15119 & ~n15771;
  assign n15774 = ~n15772 & ~n15773;
  assign n15775 = ~n15770 & n15774;
  assign n15776 = n3810 & n12485;
  assign n15777 = n3886 & n15001;
  assign n15778 = n3884 & n12482;
  assign n15779 = n4380 & n12479;
  assign n15780 = ~n15776 & ~n15778;
  assign n15781 = ~n15779 & n15780;
  assign n15782 = ~n15777 & n15781;
  assign n15783 = ~pi29  & ~n15782;
  assign n15784 = pi29  & n15782;
  assign n15785 = ~n15783 & ~n15784;
  assign n15786 = ~n15067 & n15075;
  assign n15787 = n15067 & ~n15075;
  assign n15788 = ~n15786 & ~n15787;
  assign n15789 = ~n15785 & ~n15788;
  assign n15790 = ~n746 & n12492;
  assign n15791 = ~n3807 & n12492;
  assign n15792 = n3884 & n12492;
  assign n15793 = n4380 & n12490;
  assign n15794 = n3886 & ~n15072;
  assign n15795 = ~n15792 & ~n15793;
  assign n15796 = ~n15794 & n15795;
  assign n15797 = pi29  & ~n15791;
  assign n15798 = n15796 & n15797;
  assign n15799 = n3810 & n12492;
  assign n15800 = n3886 & ~n15113;
  assign n15801 = n3884 & n12490;
  assign n15802 = n4380 & n12485;
  assign n15803 = ~n15799 & ~n15801;
  assign n15804 = ~n15802 & n15803;
  assign n15805 = ~n15800 & n15804;
  assign n15806 = n15798 & n15805;
  assign n15807 = n15790 & n15806;
  assign n15808 = n3810 & n12490;
  assign n15809 = n3886 & n15026;
  assign n15810 = n3884 & n12485;
  assign n15811 = n4380 & n12482;
  assign n15812 = ~n15808 & ~n15810;
  assign n15813 = ~n15811 & n15812;
  assign n15814 = ~n15809 & n15813;
  assign n15815 = ~pi29  & ~n15814;
  assign n15816 = pi29  & n15814;
  assign n15817 = ~n15815 & ~n15816;
  assign n15818 = ~n15790 & n15806;
  assign n15819 = n15790 & ~n15806;
  assign n15820 = ~n15818 & ~n15819;
  assign n15821 = ~n15817 & ~n15820;
  assign n15822 = ~n15807 & ~n15821;
  assign n15823 = n15785 & n15788;
  assign n15824 = ~n15789 & ~n15823;
  assign n15825 = ~n15822 & n15824;
  assign n15826 = ~n15789 & ~n15825;
  assign n15827 = n15770 & ~n15774;
  assign n15828 = ~n15775 & ~n15827;
  assign n15829 = ~n15826 & n15828;
  assign n15830 = ~n15775 & ~n15829;
  assign n15831 = ~n15760 & ~n15830;
  assign n15832 = ~n15757 & ~n15831;
  assign n15833 = ~n15744 & ~n15832;
  assign n15834 = ~n15741 & ~n15833;
  assign n15835 = ~n15728 & ~n15834;
  assign n15836 = ~n15725 & ~n15835;
  assign n15837 = n15709 & ~n15711;
  assign n15838 = ~n15712 & ~n15837;
  assign n15839 = ~n15836 & n15838;
  assign n15840 = ~n15712 & ~n15839;
  assign n15841 = n15696 & ~n15698;
  assign n15842 = ~n15699 & ~n15841;
  assign n15843 = ~n15840 & n15842;
  assign n15844 = ~n15699 & ~n15843;
  assign n15845 = n15683 & ~n15685;
  assign n15846 = ~n15686 & ~n15845;
  assign n15847 = ~n15844 & n15846;
  assign n15848 = ~n15686 & ~n15847;
  assign n15849 = n15670 & ~n15672;
  assign n15850 = ~n15673 & ~n15849;
  assign n15851 = ~n15848 & n15850;
  assign n15852 = ~n15673 & ~n15851;
  assign n15853 = n15657 & ~n15659;
  assign n15854 = ~n15660 & ~n15853;
  assign n15855 = ~n15852 & n15854;
  assign n15856 = ~n15660 & ~n15855;
  assign n15857 = ~n15165 & n15175;
  assign n15858 = ~n15176 & ~n15857;
  assign n15859 = ~n15856 & n15858;
  assign n15860 = n15856 & ~n15858;
  assign n15861 = n86 & n12446;
  assign n15862 = n4420 & n14175;
  assign n15863 = n4600 & n12443;
  assign n15864 = n4615 & n12440;
  assign n15865 = ~n15861 & ~n15863;
  assign n15866 = ~n15864 & n15865;
  assign n15867 = ~n15862 & n15866;
  assign n15868 = pi26  & n15867;
  assign n15869 = ~pi26  & ~n15867;
  assign n15870 = ~n15868 & ~n15869;
  assign n15871 = ~n15860 & ~n15870;
  assign n15872 = ~n15859 & ~n15871;
  assign n15873 = ~n15647 & ~n15872;
  assign n15874 = n15647 & n15872;
  assign n15875 = n5044 & n12434;
  assign n15876 = n5045 & n13546;
  assign n15877 = n5109 & n12431;
  assign n15878 = n5130 & n12428;
  assign n15879 = ~n15875 & ~n15877;
  assign n15880 = ~n15878 & n15879;
  assign n15881 = ~n15876 & n15880;
  assign n15882 = pi23  & n15881;
  assign n15883 = ~pi23  & ~n15881;
  assign n15884 = ~n15882 & ~n15883;
  assign n15885 = ~n15874 & ~n15884;
  assign n15886 = ~n15873 & ~n15885;
  assign n15887 = n15644 & ~n15886;
  assign n15888 = ~n15644 & n15886;
  assign n15889 = n5240 & n12422;
  assign n15890 = n5241 & n13201;
  assign n15891 = n5853 & n12419;
  assign n15892 = n5866 & n12416;
  assign n15893 = ~n15889 & ~n15891;
  assign n15894 = ~n15892 & n15893;
  assign n15895 = ~n15890 & n15894;
  assign n15896 = pi20  & n15895;
  assign n15897 = ~pi20  & ~n15895;
  assign n15898 = ~n15896 & ~n15897;
  assign n15899 = ~n15888 & ~n15898;
  assign n15900 = ~n15887 & ~n15899;
  assign n15901 = ~n15640 & ~n15900;
  assign n15902 = ~n15637 & ~n15901;
  assign n15903 = ~n15544 & ~n15545;
  assign n15904 = ~n15555 & n15903;
  assign n15905 = n15555 & ~n15903;
  assign n15906 = ~n15904 & ~n15905;
  assign n15907 = ~n15902 & n15906;
  assign n15908 = n15902 & ~n15906;
  assign n15909 = n5982 & n12407;
  assign n15910 = n5983 & n13035;
  assign n15911 = n6323 & n12404;
  assign n15912 = n6336 & n12401;
  assign n15913 = ~n15909 & ~n15911;
  assign n15914 = ~n15912 & n15913;
  assign n15915 = ~n15910 & n15914;
  assign n15916 = pi17  & n15915;
  assign n15917 = ~pi17  & ~n15915;
  assign n15918 = ~n15916 & ~n15917;
  assign n15919 = ~n15908 & ~n15918;
  assign n15920 = ~n15907 & ~n15919;
  assign n15921 = n15624 & ~n15920;
  assign n15922 = ~n15624 & n15920;
  assign n15923 = n6630 & n12395;
  assign n15924 = n6631 & n13144;
  assign n15925 = n7238 & n12362;
  assign n15926 = n7262 & n12392;
  assign n15927 = ~n15923 & ~n15925;
  assign n15928 = ~n15926 & n15927;
  assign n15929 = ~n15924 & n15928;
  assign n15930 = pi14  & n15929;
  assign n15931 = ~pi14  & ~n15929;
  assign n15932 = ~n15930 & ~n15931;
  assign n15933 = ~n15922 & ~n15932;
  assign n15934 = ~n15921 & ~n15933;
  assign n15935 = ~n15620 & ~n15934;
  assign n15936 = ~n15617 & ~n15935;
  assign n15937 = ~n15578 & ~n15579;
  assign n15938 = ~n15589 & n15937;
  assign n15939 = n15589 & ~n15937;
  assign n15940 = ~n15938 & ~n15939;
  assign n15941 = ~n15936 & n15940;
  assign n15942 = n15936 & ~n15940;
  assign n15943 = n7895 & ~n12786;
  assign n15944 = n7431 & ~n13781;
  assign n15945 = n7430 & n13166;
  assign n15946 = n7869 & n13161;
  assign n15947 = ~n15943 & ~n15945;
  assign n15948 = ~n15946 & n15947;
  assign n15949 = ~n15944 & n15948;
  assign n15950 = pi11  & n15949;
  assign n15951 = ~pi11  & ~n15949;
  assign n15952 = ~n15950 & ~n15951;
  assign n15953 = ~n15942 & ~n15952;
  assign n15954 = ~n15941 & ~n15953;
  assign n15955 = n15604 & ~n15954;
  assign n15956 = ~n15604 & n15954;
  assign n15957 = ~n15955 & ~n15956;
  assign n15958 = n7895 & n13161;
  assign n15959 = n7431 & n13183;
  assign n15960 = n7869 & n13166;
  assign n15961 = n7430 & n13164;
  assign n15962 = ~n15960 & ~n15961;
  assign n15963 = ~n15958 & n15962;
  assign n15964 = ~n15959 & n15963;
  assign n15965 = pi11  & n15964;
  assign n15966 = ~pi11  & ~n15964;
  assign n15967 = ~n15965 & ~n15966;
  assign n15968 = ~n15921 & ~n15922;
  assign n15969 = ~n15932 & n15968;
  assign n15970 = n15932 & ~n15968;
  assign n15971 = ~n15969 & ~n15970;
  assign n15972 = n15640 & n15900;
  assign n15973 = ~n15901 & ~n15972;
  assign n15974 = n5982 & n12410;
  assign n15975 = n5983 & n13093;
  assign n15976 = n6323 & n12407;
  assign n15977 = n6336 & n12404;
  assign n15978 = ~n15974 & ~n15976;
  assign n15979 = ~n15977 & n15978;
  assign n15980 = ~n15975 & n15979;
  assign n15981 = pi17  & n15980;
  assign n15982 = ~pi17  & ~n15980;
  assign n15983 = ~n15981 & ~n15982;
  assign n15984 = n15973 & ~n15983;
  assign n15985 = n15973 & n15983;
  assign n15986 = ~n15973 & ~n15983;
  assign n15987 = ~n15985 & ~n15986;
  assign n15988 = ~n15887 & ~n15888;
  assign n15989 = ~n15898 & n15988;
  assign n15990 = n15898 & ~n15988;
  assign n15991 = ~n15989 & ~n15990;
  assign n15992 = ~n15873 & ~n15874;
  assign n15993 = ~n15884 & n15992;
  assign n15994 = n15884 & ~n15992;
  assign n15995 = ~n15993 & ~n15994;
  assign n15996 = n15852 & ~n15854;
  assign n15997 = ~n15855 & ~n15996;
  assign n15998 = n86 & n12449;
  assign n15999 = n4420 & n14325;
  assign n16000 = n4600 & n12446;
  assign n16001 = n4615 & n12443;
  assign n16002 = ~n15998 & ~n16000;
  assign n16003 = ~n16001 & n16002;
  assign n16004 = ~n15999 & n16003;
  assign n16005 = pi26  & n16004;
  assign n16006 = ~pi26  & ~n16004;
  assign n16007 = ~n16005 & ~n16006;
  assign n16008 = n15997 & ~n16007;
  assign n16009 = n15848 & ~n15850;
  assign n16010 = ~n15851 & ~n16009;
  assign n16011 = n86 & n12452;
  assign n16012 = n4420 & n14156;
  assign n16013 = n4600 & n12449;
  assign n16014 = n4615 & n12446;
  assign n16015 = ~n16011 & ~n16013;
  assign n16016 = ~n16014 & n16015;
  assign n16017 = ~n16012 & n16016;
  assign n16018 = pi26  & n16017;
  assign n16019 = ~pi26  & ~n16017;
  assign n16020 = ~n16018 & ~n16019;
  assign n16021 = n16010 & ~n16020;
  assign n16022 = n15844 & ~n15846;
  assign n16023 = ~n15847 & ~n16022;
  assign n16024 = n86 & n12455;
  assign n16025 = n4420 & n14442;
  assign n16026 = n4600 & n12452;
  assign n16027 = n4615 & n12449;
  assign n16028 = ~n16024 & ~n16026;
  assign n16029 = ~n16027 & n16028;
  assign n16030 = ~n16025 & n16029;
  assign n16031 = pi26  & n16030;
  assign n16032 = ~pi26  & ~n16030;
  assign n16033 = ~n16031 & ~n16032;
  assign n16034 = n16023 & ~n16033;
  assign n16035 = n15840 & ~n15842;
  assign n16036 = ~n15843 & ~n16035;
  assign n16037 = n86 & n12458;
  assign n16038 = n4420 & n14741;
  assign n16039 = n4600 & n12455;
  assign n16040 = n4615 & n12452;
  assign n16041 = ~n16037 & ~n16039;
  assign n16042 = ~n16040 & n16041;
  assign n16043 = ~n16038 & n16042;
  assign n16044 = pi26  & n16043;
  assign n16045 = ~pi26  & ~n16043;
  assign n16046 = ~n16044 & ~n16045;
  assign n16047 = n16036 & ~n16046;
  assign n16048 = n15836 & ~n15838;
  assign n16049 = ~n15839 & ~n16048;
  assign n16050 = n86 & n12461;
  assign n16051 = n4420 & n14756;
  assign n16052 = n4600 & n12458;
  assign n16053 = n4615 & n12455;
  assign n16054 = ~n16050 & ~n16052;
  assign n16055 = ~n16053 & n16054;
  assign n16056 = ~n16051 & n16055;
  assign n16057 = pi26  & n16056;
  assign n16058 = ~pi26  & ~n16056;
  assign n16059 = ~n16057 & ~n16058;
  assign n16060 = n16049 & ~n16059;
  assign n16061 = n15728 & n15834;
  assign n16062 = ~n15835 & ~n16061;
  assign n16063 = n86 & n12464;
  assign n16064 = n4420 & n14420;
  assign n16065 = n4600 & n12461;
  assign n16066 = n4615 & n12458;
  assign n16067 = ~n16063 & ~n16065;
  assign n16068 = ~n16066 & n16067;
  assign n16069 = ~n16064 & n16068;
  assign n16070 = pi26  & n16069;
  assign n16071 = ~pi26  & ~n16069;
  assign n16072 = ~n16070 & ~n16071;
  assign n16073 = n16062 & ~n16072;
  assign n16074 = n15744 & n15832;
  assign n16075 = ~n15833 & ~n16074;
  assign n16076 = n86 & n12467;
  assign n16077 = n4420 & n14789;
  assign n16078 = n4600 & n12464;
  assign n16079 = n4615 & n12461;
  assign n16080 = ~n16076 & ~n16078;
  assign n16081 = ~n16079 & n16080;
  assign n16082 = ~n16077 & n16081;
  assign n16083 = pi26  & n16082;
  assign n16084 = ~pi26  & ~n16082;
  assign n16085 = ~n16083 & ~n16084;
  assign n16086 = n16075 & ~n16085;
  assign n16087 = n15760 & n15830;
  assign n16088 = ~n15831 & ~n16087;
  assign n16089 = n86 & n12470;
  assign n16090 = n4420 & n14815;
  assign n16091 = n4600 & n12467;
  assign n16092 = n4615 & n12464;
  assign n16093 = ~n16089 & ~n16091;
  assign n16094 = ~n16092 & n16093;
  assign n16095 = ~n16090 & n16094;
  assign n16096 = pi26  & n16095;
  assign n16097 = ~pi26  & ~n16095;
  assign n16098 = ~n16096 & ~n16097;
  assign n16099 = n16088 & ~n16098;
  assign n16100 = n15826 & ~n15828;
  assign n16101 = ~n15829 & ~n16100;
  assign n16102 = n4600 & n12470;
  assign n16103 = n4420 & n14839;
  assign n16104 = n86 & n12473;
  assign n16105 = n4615 & n12467;
  assign n16106 = ~n16102 & ~n16104;
  assign n16107 = ~n16105 & n16106;
  assign n16108 = ~n16103 & n16107;
  assign n16109 = pi26  & n16108;
  assign n16110 = ~pi26  & ~n16108;
  assign n16111 = ~n16109 & ~n16110;
  assign n16112 = n16101 & ~n16111;
  assign n16113 = n86 & n12476;
  assign n16114 = n4420 & n14849;
  assign n16115 = n4600 & n12473;
  assign n16116 = n4615 & n12470;
  assign n16117 = ~n16113 & ~n16115;
  assign n16118 = ~n16116 & n16117;
  assign n16119 = ~n16114 & n16118;
  assign n16120 = pi26  & n16119;
  assign n16121 = ~pi26  & ~n16119;
  assign n16122 = ~n16120 & ~n16121;
  assign n16123 = n15822 & ~n15824;
  assign n16124 = ~n15825 & ~n16123;
  assign n16125 = ~n16122 & n16124;
  assign n16126 = n4600 & n12476;
  assign n16127 = n4420 & n14922;
  assign n16128 = n86 & n12479;
  assign n16129 = n4615 & n12473;
  assign n16130 = ~n16126 & ~n16128;
  assign n16131 = ~n16129 & n16130;
  assign n16132 = ~n16127 & n16131;
  assign n16133 = ~pi26  & ~n16132;
  assign n16134 = pi26  & n16132;
  assign n16135 = ~n16133 & ~n16134;
  assign n16136 = n15817 & n15820;
  assign n16137 = ~n15821 & ~n16136;
  assign n16138 = ~n16135 & n16137;
  assign n16139 = ~n16135 & ~n16137;
  assign n16140 = n16135 & n16137;
  assign n16141 = ~n16139 & ~n16140;
  assign n16142 = n86 & n12482;
  assign n16143 = n4420 & n14958;
  assign n16144 = n4600 & n12479;
  assign n16145 = n4615 & n12476;
  assign n16146 = ~n16142 & ~n16144;
  assign n16147 = ~n16145 & n16146;
  assign n16148 = ~n16143 & n16147;
  assign n16149 = ~pi26  & ~n16148;
  assign n16150 = pi26  & n16148;
  assign n16151 = ~n16149 & ~n16150;
  assign n16152 = pi29  & ~n15798;
  assign n16153 = n15805 & ~n16152;
  assign n16154 = ~n15805 & n16152;
  assign n16155 = ~n16153 & ~n16154;
  assign n16156 = ~n16151 & n16155;
  assign n16157 = ~n16151 & ~n16155;
  assign n16158 = n16151 & n16155;
  assign n16159 = ~n16157 & ~n16158;
  assign n16160 = n86 & n12485;
  assign n16161 = n4420 & n15001;
  assign n16162 = n4600 & n12482;
  assign n16163 = n4615 & n12479;
  assign n16164 = ~n16160 & ~n16162;
  assign n16165 = ~n16163 & n16164;
  assign n16166 = ~n16161 & n16165;
  assign n16167 = pi26  & n16166;
  assign n16168 = ~pi26  & ~n16166;
  assign n16169 = ~n16167 & ~n16168;
  assign n16170 = pi29  & n15791;
  assign n16171 = ~n15796 & n16170;
  assign n16172 = n15796 & ~n16170;
  assign n16173 = ~n16171 & ~n16172;
  assign n16174 = ~n16169 & n16173;
  assign n16175 = ~n81 & n12492;
  assign n16176 = n4615 & n12490;
  assign n16177 = n4600 & n12492;
  assign n16178 = n4420 & ~n15072;
  assign n16179 = ~n16176 & ~n16177;
  assign n16180 = ~n16178 & n16179;
  assign n16181 = pi26  & ~n16175;
  assign n16182 = n16180 & n16181;
  assign n16183 = n86 & n12492;
  assign n16184 = n4420 & ~n15113;
  assign n16185 = n4600 & n12490;
  assign n16186 = n4615 & n12485;
  assign n16187 = ~n16183 & ~n16185;
  assign n16188 = ~n16186 & n16187;
  assign n16189 = ~n16184 & n16188;
  assign n16190 = n16182 & n16189;
  assign n16191 = n15791 & n16190;
  assign n16192 = ~n15791 & n16190;
  assign n16193 = n15791 & ~n16190;
  assign n16194 = ~n16192 & ~n16193;
  assign n16195 = n86 & n12490;
  assign n16196 = n4420 & n15026;
  assign n16197 = n4600 & n12485;
  assign n16198 = n4615 & n12482;
  assign n16199 = ~n16195 & ~n16197;
  assign n16200 = ~n16198 & n16199;
  assign n16201 = ~n16196 & n16200;
  assign n16202 = pi26  & n16201;
  assign n16203 = ~pi26  & ~n16201;
  assign n16204 = ~n16202 & ~n16203;
  assign n16205 = ~n16194 & ~n16204;
  assign n16206 = ~n16191 & ~n16205;
  assign n16207 = n16169 & ~n16173;
  assign n16208 = ~n16174 & ~n16207;
  assign n16209 = ~n16206 & n16208;
  assign n16210 = ~n16174 & ~n16209;
  assign n16211 = ~n16159 & ~n16210;
  assign n16212 = ~n16156 & ~n16211;
  assign n16213 = ~n16141 & ~n16212;
  assign n16214 = ~n16138 & ~n16213;
  assign n16215 = n16122 & n16124;
  assign n16216 = ~n16122 & ~n16124;
  assign n16217 = ~n16215 & ~n16216;
  assign n16218 = ~n16214 & ~n16217;
  assign n16219 = ~n16125 & ~n16218;
  assign n16220 = n16101 & n16111;
  assign n16221 = ~n16101 & ~n16111;
  assign n16222 = ~n16220 & ~n16221;
  assign n16223 = ~n16219 & ~n16222;
  assign n16224 = ~n16112 & ~n16223;
  assign n16225 = n16088 & n16098;
  assign n16226 = ~n16088 & ~n16098;
  assign n16227 = ~n16225 & ~n16226;
  assign n16228 = ~n16224 & ~n16227;
  assign n16229 = ~n16099 & ~n16228;
  assign n16230 = n16075 & n16085;
  assign n16231 = ~n16075 & ~n16085;
  assign n16232 = ~n16230 & ~n16231;
  assign n16233 = ~n16229 & ~n16232;
  assign n16234 = ~n16086 & ~n16233;
  assign n16235 = n16062 & n16072;
  assign n16236 = ~n16062 & ~n16072;
  assign n16237 = ~n16235 & ~n16236;
  assign n16238 = ~n16234 & ~n16237;
  assign n16239 = ~n16073 & ~n16238;
  assign n16240 = n16049 & n16059;
  assign n16241 = ~n16049 & ~n16059;
  assign n16242 = ~n16240 & ~n16241;
  assign n16243 = ~n16239 & ~n16242;
  assign n16244 = ~n16060 & ~n16243;
  assign n16245 = n16036 & n16046;
  assign n16246 = ~n16036 & ~n16046;
  assign n16247 = ~n16245 & ~n16246;
  assign n16248 = ~n16244 & ~n16247;
  assign n16249 = ~n16047 & ~n16248;
  assign n16250 = n16023 & n16033;
  assign n16251 = ~n16023 & ~n16033;
  assign n16252 = ~n16250 & ~n16251;
  assign n16253 = ~n16249 & ~n16252;
  assign n16254 = ~n16034 & ~n16253;
  assign n16255 = n16010 & n16020;
  assign n16256 = ~n16010 & ~n16020;
  assign n16257 = ~n16255 & ~n16256;
  assign n16258 = ~n16254 & ~n16257;
  assign n16259 = ~n16021 & ~n16258;
  assign n16260 = ~n15997 & n16007;
  assign n16261 = ~n16008 & ~n16260;
  assign n16262 = ~n16259 & n16261;
  assign n16263 = ~n16008 & ~n16262;
  assign n16264 = ~n15859 & ~n15860;
  assign n16265 = ~n15870 & n16264;
  assign n16266 = n15870 & ~n16264;
  assign n16267 = ~n16265 & ~n16266;
  assign n16268 = ~n16263 & n16267;
  assign n16269 = n16263 & ~n16267;
  assign n16270 = n5044 & n12437;
  assign n16271 = n5045 & n13564;
  assign n16272 = n5109 & n12434;
  assign n16273 = n5130 & n12431;
  assign n16274 = ~n16270 & ~n16272;
  assign n16275 = ~n16273 & n16274;
  assign n16276 = ~n16271 & n16275;
  assign n16277 = pi23  & n16276;
  assign n16278 = ~pi23  & ~n16276;
  assign n16279 = ~n16277 & ~n16278;
  assign n16280 = ~n16269 & ~n16279;
  assign n16281 = ~n16268 & ~n16280;
  assign n16282 = n15995 & ~n16281;
  assign n16283 = ~n15995 & n16281;
  assign n16284 = n5240 & n12425;
  assign n16285 = n5241 & n13010;
  assign n16286 = n5853 & n12422;
  assign n16287 = n5866 & n12419;
  assign n16288 = ~n16284 & ~n16286;
  assign n16289 = ~n16287 & n16288;
  assign n16290 = ~n16285 & n16289;
  assign n16291 = pi20  & n16290;
  assign n16292 = ~pi20  & ~n16290;
  assign n16293 = ~n16291 & ~n16292;
  assign n16294 = ~n16283 & ~n16293;
  assign n16295 = ~n16282 & ~n16294;
  assign n16296 = n15991 & ~n16295;
  assign n16297 = ~n15991 & n16295;
  assign n16298 = n5982 & n12413;
  assign n16299 = n5983 & n12891;
  assign n16300 = n6323 & n12410;
  assign n16301 = n6336 & n12407;
  assign n16302 = ~n16298 & ~n16300;
  assign n16303 = ~n16301 & n16302;
  assign n16304 = ~n16299 & n16303;
  assign n16305 = pi17  & n16304;
  assign n16306 = ~pi17  & ~n16304;
  assign n16307 = ~n16305 & ~n16306;
  assign n16308 = ~n16297 & ~n16307;
  assign n16309 = ~n16296 & ~n16308;
  assign n16310 = ~n15987 & ~n16309;
  assign n16311 = ~n15984 & ~n16310;
  assign n16312 = ~n15907 & ~n15908;
  assign n16313 = ~n15918 & n16312;
  assign n16314 = n15918 & ~n16312;
  assign n16315 = ~n16313 & ~n16314;
  assign n16316 = ~n16311 & n16315;
  assign n16317 = n16311 & ~n16315;
  assign n16318 = n6630 & n12398;
  assign n16319 = n6631 & n13245;
  assign n16320 = n7238 & n12395;
  assign n16321 = n7262 & n12362;
  assign n16322 = ~n16318 & ~n16320;
  assign n16323 = ~n16321 & n16322;
  assign n16324 = ~n16319 & n16323;
  assign n16325 = pi14  & n16324;
  assign n16326 = ~pi14  & ~n16324;
  assign n16327 = ~n16325 & ~n16326;
  assign n16328 = ~n16317 & ~n16327;
  assign n16329 = ~n16316 & ~n16328;
  assign n16330 = n15971 & ~n16329;
  assign n16331 = ~n15971 & n16329;
  assign n16332 = n7430 & n12646;
  assign n16333 = n7431 & n13261;
  assign n16334 = n7869 & n13164;
  assign n16335 = n7895 & n13166;
  assign n16336 = ~n16332 & ~n16334;
  assign n16337 = ~n16335 & n16336;
  assign n16338 = ~n16333 & n16337;
  assign n16339 = pi11  & n16338;
  assign n16340 = ~pi11  & ~n16338;
  assign n16341 = ~n16339 & ~n16340;
  assign n16342 = ~n16331 & ~n16341;
  assign n16343 = ~n16330 & ~n16342;
  assign n16344 = ~n15967 & ~n16343;
  assign n16345 = n15620 & n15934;
  assign n16346 = ~n15935 & ~n16345;
  assign n16347 = n15967 & ~n16343;
  assign n16348 = ~n15967 & n16343;
  assign n16349 = ~n16347 & ~n16348;
  assign n16350 = n16346 & ~n16349;
  assign n16351 = ~n16344 & ~n16350;
  assign n16352 = ~n15941 & ~n15942;
  assign n16353 = ~n15952 & n16352;
  assign n16354 = n15952 & ~n16352;
  assign n16355 = ~n16353 & ~n16354;
  assign n16356 = ~n16351 & n16355;
  assign n16357 = n16351 & n16355;
  assign n16358 = ~n16351 & ~n16355;
  assign n16359 = ~n16357 & ~n16358;
  assign n16360 = ~n16346 & n16349;
  assign n16361 = ~n16350 & ~n16360;
  assign n16362 = n8251 & ~n13280;
  assign n16363 = n8250 & ~n13160;
  assign n16364 = ~n9016 & ~n9040;
  assign n16365 = ~n16363 & n16364;
  assign n16366 = ~n12786 & ~n16365;
  assign n16367 = ~n16362 & ~n16366;
  assign n16368 = pi8  & n16367;
  assign n16369 = ~pi8  & ~n16367;
  assign n16370 = ~n16368 & ~n16369;
  assign n16371 = n15987 & n16309;
  assign n16372 = ~n16310 & ~n16371;
  assign n16373 = n6630 & n12401;
  assign n16374 = n6631 & n13108;
  assign n16375 = n7238 & n12398;
  assign n16376 = n7262 & n12395;
  assign n16377 = ~n16373 & ~n16375;
  assign n16378 = ~n16376 & n16377;
  assign n16379 = ~n16374 & n16378;
  assign n16380 = pi14  & n16379;
  assign n16381 = ~pi14  & ~n16379;
  assign n16382 = ~n16380 & ~n16381;
  assign n16383 = n16372 & ~n16382;
  assign n16384 = n16372 & n16382;
  assign n16385 = ~n16372 & ~n16382;
  assign n16386 = ~n16384 & ~n16385;
  assign n16387 = ~n16296 & ~n16297;
  assign n16388 = ~n16307 & n16387;
  assign n16389 = n16307 & ~n16387;
  assign n16390 = ~n16388 & ~n16389;
  assign n16391 = ~n16282 & ~n16283;
  assign n16392 = ~n16293 & n16391;
  assign n16393 = n16293 & ~n16391;
  assign n16394 = ~n16392 & ~n16393;
  assign n16395 = n5044 & n12440;
  assign n16396 = n5045 & n13939;
  assign n16397 = n5109 & n12437;
  assign n16398 = n5130 & n12434;
  assign n16399 = ~n16395 & ~n16397;
  assign n16400 = ~n16398 & n16399;
  assign n16401 = ~n16396 & n16400;
  assign n16402 = ~pi23  & ~n16401;
  assign n16403 = pi23  & n16401;
  assign n16404 = ~n16402 & ~n16403;
  assign n16405 = n16259 & ~n16261;
  assign n16406 = ~n16262 & ~n16405;
  assign n16407 = ~n16404 & n16406;
  assign n16408 = ~n16404 & ~n16406;
  assign n16409 = n16404 & n16406;
  assign n16410 = ~n16408 & ~n16409;
  assign n16411 = n5044 & n12443;
  assign n16412 = n5045 & n13702;
  assign n16413 = n5109 & n12440;
  assign n16414 = n5130 & n12437;
  assign n16415 = ~n16411 & ~n16413;
  assign n16416 = ~n16414 & n16415;
  assign n16417 = ~n16412 & n16416;
  assign n16418 = ~pi23  & ~n16417;
  assign n16419 = pi23  & n16417;
  assign n16420 = ~n16418 & ~n16419;
  assign n16421 = n16254 & n16257;
  assign n16422 = ~n16258 & ~n16421;
  assign n16423 = ~n16420 & n16422;
  assign n16424 = ~n16420 & ~n16422;
  assign n16425 = n16420 & n16422;
  assign n16426 = ~n16424 & ~n16425;
  assign n16427 = n5044 & n12446;
  assign n16428 = n5045 & n14175;
  assign n16429 = n5109 & n12443;
  assign n16430 = n5130 & n12440;
  assign n16431 = ~n16427 & ~n16429;
  assign n16432 = ~n16430 & n16431;
  assign n16433 = ~n16428 & n16432;
  assign n16434 = ~pi23  & ~n16433;
  assign n16435 = pi23  & n16433;
  assign n16436 = ~n16434 & ~n16435;
  assign n16437 = n16249 & n16252;
  assign n16438 = ~n16253 & ~n16437;
  assign n16439 = ~n16436 & n16438;
  assign n16440 = ~n16436 & ~n16438;
  assign n16441 = n16436 & n16438;
  assign n16442 = ~n16440 & ~n16441;
  assign n16443 = n5044 & n12449;
  assign n16444 = n5045 & n14325;
  assign n16445 = n5109 & n12446;
  assign n16446 = n5130 & n12443;
  assign n16447 = ~n16443 & ~n16445;
  assign n16448 = ~n16446 & n16447;
  assign n16449 = ~n16444 & n16448;
  assign n16450 = ~pi23  & ~n16449;
  assign n16451 = pi23  & n16449;
  assign n16452 = ~n16450 & ~n16451;
  assign n16453 = n16244 & n16247;
  assign n16454 = ~n16248 & ~n16453;
  assign n16455 = ~n16452 & n16454;
  assign n16456 = ~n16452 & ~n16454;
  assign n16457 = n16452 & n16454;
  assign n16458 = ~n16456 & ~n16457;
  assign n16459 = n5044 & n12452;
  assign n16460 = n5045 & n14156;
  assign n16461 = n5109 & n12449;
  assign n16462 = n5130 & n12446;
  assign n16463 = ~n16459 & ~n16461;
  assign n16464 = ~n16462 & n16463;
  assign n16465 = ~n16460 & n16464;
  assign n16466 = ~pi23  & ~n16465;
  assign n16467 = pi23  & n16465;
  assign n16468 = ~n16466 & ~n16467;
  assign n16469 = n16239 & n16242;
  assign n16470 = ~n16243 & ~n16469;
  assign n16471 = ~n16468 & n16470;
  assign n16472 = ~n16468 & ~n16470;
  assign n16473 = n16468 & n16470;
  assign n16474 = ~n16472 & ~n16473;
  assign n16475 = n5044 & n12455;
  assign n16476 = n5045 & n14442;
  assign n16477 = n5109 & n12452;
  assign n16478 = n5130 & n12449;
  assign n16479 = ~n16475 & ~n16477;
  assign n16480 = ~n16478 & n16479;
  assign n16481 = ~n16476 & n16480;
  assign n16482 = ~pi23  & ~n16481;
  assign n16483 = pi23  & n16481;
  assign n16484 = ~n16482 & ~n16483;
  assign n16485 = ~n16234 & n16237;
  assign n16486 = n16234 & ~n16237;
  assign n16487 = ~n16485 & ~n16486;
  assign n16488 = ~n16484 & ~n16487;
  assign n16489 = n5044 & n12458;
  assign n16490 = n5045 & n14741;
  assign n16491 = n5109 & n12455;
  assign n16492 = n5130 & n12452;
  assign n16493 = ~n16489 & ~n16491;
  assign n16494 = ~n16492 & n16493;
  assign n16495 = ~n16490 & n16494;
  assign n16496 = ~pi23  & ~n16495;
  assign n16497 = pi23  & n16495;
  assign n16498 = ~n16496 & ~n16497;
  assign n16499 = ~n16229 & n16232;
  assign n16500 = n16229 & ~n16232;
  assign n16501 = ~n16499 & ~n16500;
  assign n16502 = ~n16498 & ~n16501;
  assign n16503 = n5044 & n12461;
  assign n16504 = n5045 & n14756;
  assign n16505 = n5109 & n12458;
  assign n16506 = n5130 & n12455;
  assign n16507 = ~n16503 & ~n16505;
  assign n16508 = ~n16506 & n16507;
  assign n16509 = ~n16504 & n16508;
  assign n16510 = ~pi23  & ~n16509;
  assign n16511 = pi23  & n16509;
  assign n16512 = ~n16510 & ~n16511;
  assign n16513 = ~n16224 & n16227;
  assign n16514 = n16224 & ~n16227;
  assign n16515 = ~n16513 & ~n16514;
  assign n16516 = ~n16512 & ~n16515;
  assign n16517 = n5044 & n12464;
  assign n16518 = n5045 & n14420;
  assign n16519 = n5109 & n12461;
  assign n16520 = n5130 & n12458;
  assign n16521 = ~n16517 & ~n16519;
  assign n16522 = ~n16520 & n16521;
  assign n16523 = ~n16518 & n16522;
  assign n16524 = ~pi23  & ~n16523;
  assign n16525 = pi23  & n16523;
  assign n16526 = ~n16524 & ~n16525;
  assign n16527 = n16219 & n16222;
  assign n16528 = ~n16223 & ~n16527;
  assign n16529 = ~n16526 & n16528;
  assign n16530 = ~n16526 & ~n16528;
  assign n16531 = n16526 & n16528;
  assign n16532 = ~n16530 & ~n16531;
  assign n16533 = n5044 & n12467;
  assign n16534 = n5045 & n14789;
  assign n16535 = n5109 & n12464;
  assign n16536 = n5130 & n12461;
  assign n16537 = ~n16533 & ~n16535;
  assign n16538 = ~n16536 & n16537;
  assign n16539 = ~n16534 & n16538;
  assign n16540 = ~pi23  & ~n16539;
  assign n16541 = pi23  & n16539;
  assign n16542 = ~n16540 & ~n16541;
  assign n16543 = n16214 & n16217;
  assign n16544 = ~n16218 & ~n16543;
  assign n16545 = ~n16542 & n16544;
  assign n16546 = ~n16542 & ~n16544;
  assign n16547 = n16542 & n16544;
  assign n16548 = ~n16546 & ~n16547;
  assign n16549 = n16141 & n16212;
  assign n16550 = ~n16213 & ~n16549;
  assign n16551 = n5044 & n12470;
  assign n16552 = n5045 & n14815;
  assign n16553 = n5109 & n12467;
  assign n16554 = n5130 & n12464;
  assign n16555 = ~n16551 & ~n16553;
  assign n16556 = ~n16554 & n16555;
  assign n16557 = ~n16552 & n16556;
  assign n16558 = pi23  & n16557;
  assign n16559 = ~pi23  & ~n16557;
  assign n16560 = ~n16558 & ~n16559;
  assign n16561 = n16550 & ~n16560;
  assign n16562 = n16159 & n16210;
  assign n16563 = ~n16211 & ~n16562;
  assign n16564 = n5044 & n12473;
  assign n16565 = n5045 & n14839;
  assign n16566 = n5109 & n12470;
  assign n16567 = n5130 & n12467;
  assign n16568 = ~n16564 & ~n16566;
  assign n16569 = ~n16567 & n16568;
  assign n16570 = ~n16565 & n16569;
  assign n16571 = pi23  & n16570;
  assign n16572 = ~pi23  & ~n16570;
  assign n16573 = ~n16571 & ~n16572;
  assign n16574 = n16563 & ~n16573;
  assign n16575 = n5044 & n12476;
  assign n16576 = n5045 & n14849;
  assign n16577 = n5109 & n12473;
  assign n16578 = n5130 & n12470;
  assign n16579 = ~n16575 & ~n16577;
  assign n16580 = ~n16578 & n16579;
  assign n16581 = ~n16576 & n16580;
  assign n16582 = ~pi23  & ~n16581;
  assign n16583 = pi23  & n16581;
  assign n16584 = ~n16582 & ~n16583;
  assign n16585 = n16206 & ~n16208;
  assign n16586 = ~n16209 & ~n16585;
  assign n16587 = ~n16584 & n16586;
  assign n16588 = ~n16584 & ~n16586;
  assign n16589 = n16584 & n16586;
  assign n16590 = ~n16588 & ~n16589;
  assign n16591 = n5044 & n12479;
  assign n16592 = n5045 & n14922;
  assign n16593 = n5109 & n12476;
  assign n16594 = n5130 & n12473;
  assign n16595 = ~n16591 & ~n16593;
  assign n16596 = ~n16594 & n16595;
  assign n16597 = ~n16592 & n16596;
  assign n16598 = pi23  & n16597;
  assign n16599 = ~pi23  & ~n16597;
  assign n16600 = ~n16598 & ~n16599;
  assign n16601 = n16194 & n16204;
  assign n16602 = ~n16205 & ~n16601;
  assign n16603 = ~n16600 & n16602;
  assign n16604 = n5044 & n12482;
  assign n16605 = n5045 & n14958;
  assign n16606 = n5109 & n12479;
  assign n16607 = n5130 & n12476;
  assign n16608 = ~n16604 & ~n16606;
  assign n16609 = ~n16607 & n16608;
  assign n16610 = ~n16605 & n16609;
  assign n16611 = ~pi23  & ~n16610;
  assign n16612 = pi23  & n16610;
  assign n16613 = ~n16611 & ~n16612;
  assign n16614 = pi26  & ~n16182;
  assign n16615 = n16189 & ~n16614;
  assign n16616 = ~n16189 & n16614;
  assign n16617 = ~n16615 & ~n16616;
  assign n16618 = ~n16613 & n16617;
  assign n16619 = ~n16613 & ~n16617;
  assign n16620 = n16613 & n16617;
  assign n16621 = ~n16619 & ~n16620;
  assign n16622 = n5044 & n12485;
  assign n16623 = n5045 & n15001;
  assign n16624 = n5109 & n12482;
  assign n16625 = n5130 & n12479;
  assign n16626 = ~n16622 & ~n16624;
  assign n16627 = ~n16625 & n16626;
  assign n16628 = ~n16623 & n16627;
  assign n16629 = pi23  & n16628;
  assign n16630 = ~pi23  & ~n16628;
  assign n16631 = ~n16629 & ~n16630;
  assign n16632 = pi26  & n16175;
  assign n16633 = ~n16180 & n16632;
  assign n16634 = n16180 & ~n16632;
  assign n16635 = ~n16633 & ~n16634;
  assign n16636 = ~n16631 & n16635;
  assign n16637 = ~n5042 & n12492;
  assign n16638 = n5109 & n12492;
  assign n16639 = n5130 & n12490;
  assign n16640 = n5045 & ~n15072;
  assign n16641 = ~n16638 & ~n16639;
  assign n16642 = ~n16640 & n16641;
  assign n16643 = pi23  & ~n16637;
  assign n16644 = n16642 & n16643;
  assign n16645 = n5044 & n12492;
  assign n16646 = n5045 & ~n15113;
  assign n16647 = n5109 & n12490;
  assign n16648 = n5130 & n12485;
  assign n16649 = ~n16645 & ~n16647;
  assign n16650 = ~n16648 & n16649;
  assign n16651 = ~n16646 & n16650;
  assign n16652 = n16644 & n16651;
  assign n16653 = n16175 & n16652;
  assign n16654 = ~n16175 & n16652;
  assign n16655 = n16175 & ~n16652;
  assign n16656 = ~n16654 & ~n16655;
  assign n16657 = n5044 & n12490;
  assign n16658 = n5045 & n15026;
  assign n16659 = n5109 & n12485;
  assign n16660 = n5130 & n12482;
  assign n16661 = ~n16657 & ~n16659;
  assign n16662 = ~n16660 & n16661;
  assign n16663 = ~n16658 & n16662;
  assign n16664 = pi23  & n16663;
  assign n16665 = ~pi23  & ~n16663;
  assign n16666 = ~n16664 & ~n16665;
  assign n16667 = ~n16656 & ~n16666;
  assign n16668 = ~n16653 & ~n16667;
  assign n16669 = n16631 & ~n16635;
  assign n16670 = ~n16636 & ~n16669;
  assign n16671 = ~n16668 & n16670;
  assign n16672 = ~n16636 & ~n16671;
  assign n16673 = ~n16621 & ~n16672;
  assign n16674 = ~n16618 & ~n16673;
  assign n16675 = n16600 & ~n16602;
  assign n16676 = ~n16603 & ~n16675;
  assign n16677 = ~n16674 & n16676;
  assign n16678 = ~n16603 & ~n16677;
  assign n16679 = ~n16590 & ~n16678;
  assign n16680 = ~n16587 & ~n16679;
  assign n16681 = n16563 & n16573;
  assign n16682 = ~n16563 & ~n16573;
  assign n16683 = ~n16681 & ~n16682;
  assign n16684 = ~n16680 & ~n16683;
  assign n16685 = ~n16574 & ~n16684;
  assign n16686 = ~n16550 & n16560;
  assign n16687 = ~n16561 & ~n16686;
  assign n16688 = ~n16685 & n16687;
  assign n16689 = ~n16561 & ~n16688;
  assign n16690 = ~n16548 & ~n16689;
  assign n16691 = ~n16545 & ~n16690;
  assign n16692 = ~n16532 & ~n16691;
  assign n16693 = ~n16529 & ~n16692;
  assign n16694 = n16512 & n16515;
  assign n16695 = ~n16516 & ~n16694;
  assign n16696 = ~n16693 & n16695;
  assign n16697 = ~n16516 & ~n16696;
  assign n16698 = n16498 & n16501;
  assign n16699 = ~n16502 & ~n16698;
  assign n16700 = ~n16697 & n16699;
  assign n16701 = ~n16502 & ~n16700;
  assign n16702 = n16484 & n16487;
  assign n16703 = ~n16488 & ~n16702;
  assign n16704 = ~n16701 & n16703;
  assign n16705 = ~n16488 & ~n16704;
  assign n16706 = ~n16474 & ~n16705;
  assign n16707 = ~n16471 & ~n16706;
  assign n16708 = ~n16458 & ~n16707;
  assign n16709 = ~n16455 & ~n16708;
  assign n16710 = ~n16442 & ~n16709;
  assign n16711 = ~n16439 & ~n16710;
  assign n16712 = ~n16426 & ~n16711;
  assign n16713 = ~n16423 & ~n16712;
  assign n16714 = ~n16410 & ~n16713;
  assign n16715 = ~n16407 & ~n16714;
  assign n16716 = ~n16268 & ~n16269;
  assign n16717 = ~n16279 & n16716;
  assign n16718 = n16279 & ~n16716;
  assign n16719 = ~n16717 & ~n16718;
  assign n16720 = ~n16715 & n16719;
  assign n16721 = n16715 & ~n16719;
  assign n16722 = n5240 & n12428;
  assign n16723 = n5241 & n13371;
  assign n16724 = n5853 & n12425;
  assign n16725 = n5866 & n12422;
  assign n16726 = ~n16722 & ~n16724;
  assign n16727 = ~n16725 & n16726;
  assign n16728 = ~n16723 & n16727;
  assign n16729 = pi20  & n16728;
  assign n16730 = ~pi20  & ~n16728;
  assign n16731 = ~n16729 & ~n16730;
  assign n16732 = ~n16721 & ~n16731;
  assign n16733 = ~n16720 & ~n16732;
  assign n16734 = n16394 & ~n16733;
  assign n16735 = ~n16394 & n16733;
  assign n16736 = n5982 & n12416;
  assign n16737 = n5983 & n12843;
  assign n16738 = n6323 & n12413;
  assign n16739 = n6336 & n12410;
  assign n16740 = ~n16736 & ~n16738;
  assign n16741 = ~n16739 & n16740;
  assign n16742 = ~n16737 & n16741;
  assign n16743 = pi17  & n16742;
  assign n16744 = ~pi17  & ~n16742;
  assign n16745 = ~n16743 & ~n16744;
  assign n16746 = ~n16735 & ~n16745;
  assign n16747 = ~n16734 & ~n16746;
  assign n16748 = n16390 & ~n16747;
  assign n16749 = ~n16390 & n16747;
  assign n16750 = n6630 & n12404;
  assign n16751 = n6631 & n13128;
  assign n16752 = n7238 & n12401;
  assign n16753 = n7262 & n12398;
  assign n16754 = ~n16750 & ~n16752;
  assign n16755 = ~n16753 & n16754;
  assign n16756 = ~n16751 & n16755;
  assign n16757 = pi14  & n16756;
  assign n16758 = ~pi14  & ~n16756;
  assign n16759 = ~n16757 & ~n16758;
  assign n16760 = ~n16749 & ~n16759;
  assign n16761 = ~n16748 & ~n16760;
  assign n16762 = ~n16386 & ~n16761;
  assign n16763 = ~n16383 & ~n16762;
  assign n16764 = ~n16316 & ~n16317;
  assign n16765 = ~n16327 & n16764;
  assign n16766 = n16327 & ~n16764;
  assign n16767 = ~n16765 & ~n16766;
  assign n16768 = ~n16763 & n16767;
  assign n16769 = n16763 & ~n16767;
  assign n16770 = n7430 & n12392;
  assign n16771 = n7431 & n13421;
  assign n16772 = n7869 & n12646;
  assign n16773 = n7895 & n13164;
  assign n16774 = ~n16770 & ~n16772;
  assign n16775 = ~n16773 & n16774;
  assign n16776 = ~n16771 & n16775;
  assign n16777 = pi11  & n16776;
  assign n16778 = ~pi11  & ~n16776;
  assign n16779 = ~n16777 & ~n16778;
  assign n16780 = ~n16769 & ~n16779;
  assign n16781 = ~n16768 & ~n16780;
  assign n16782 = ~n16370 & ~n16781;
  assign n16783 = n16370 & n16781;
  assign n16784 = ~n16330 & ~n16331;
  assign n16785 = ~n16341 & n16784;
  assign n16786 = n16341 & ~n16784;
  assign n16787 = ~n16785 & ~n16786;
  assign n16788 = ~n16783 & n16787;
  assign n16789 = ~n16782 & ~n16788;
  assign n16790 = n16361 & ~n16789;
  assign n16791 = ~n16782 & ~n16783;
  assign n16792 = n16787 & n16791;
  assign n16793 = ~n16787 & ~n16791;
  assign n16794 = ~n16792 & ~n16793;
  assign n16795 = n16386 & n16761;
  assign n16796 = ~n16762 & ~n16795;
  assign n16797 = n7430 & n12362;
  assign n16798 = n7431 & n12652;
  assign n16799 = n7869 & n12392;
  assign n16800 = n7895 & n12646;
  assign n16801 = ~n16797 & ~n16799;
  assign n16802 = ~n16800 & n16801;
  assign n16803 = ~n16798 & n16802;
  assign n16804 = pi11  & n16803;
  assign n16805 = ~pi11  & ~n16803;
  assign n16806 = ~n16804 & ~n16805;
  assign n16807 = n16796 & ~n16806;
  assign n16808 = n16796 & n16806;
  assign n16809 = ~n16796 & ~n16806;
  assign n16810 = ~n16808 & ~n16809;
  assign n16811 = ~n16748 & ~n16749;
  assign n16812 = ~n16759 & n16811;
  assign n16813 = n16759 & ~n16811;
  assign n16814 = ~n16812 & ~n16813;
  assign n16815 = ~n16734 & ~n16735;
  assign n16816 = ~n16745 & n16815;
  assign n16817 = n16745 & ~n16815;
  assign n16818 = ~n16816 & ~n16817;
  assign n16819 = n16410 & n16713;
  assign n16820 = ~n16714 & ~n16819;
  assign n16821 = n5240 & n12431;
  assign n16822 = n5241 & n13356;
  assign n16823 = n5853 & n12428;
  assign n16824 = n5866 & n12425;
  assign n16825 = ~n16821 & ~n16823;
  assign n16826 = ~n16824 & n16825;
  assign n16827 = ~n16822 & n16826;
  assign n16828 = pi20  & n16827;
  assign n16829 = ~pi20  & ~n16827;
  assign n16830 = ~n16828 & ~n16829;
  assign n16831 = n16820 & ~n16830;
  assign n16832 = n16426 & n16711;
  assign n16833 = ~n16712 & ~n16832;
  assign n16834 = n5240 & n12434;
  assign n16835 = n5241 & n13546;
  assign n16836 = n5853 & n12431;
  assign n16837 = n5866 & n12428;
  assign n16838 = ~n16834 & ~n16836;
  assign n16839 = ~n16837 & n16838;
  assign n16840 = ~n16835 & n16839;
  assign n16841 = pi20  & n16840;
  assign n16842 = ~pi20  & ~n16840;
  assign n16843 = ~n16841 & ~n16842;
  assign n16844 = n16833 & ~n16843;
  assign n16845 = n16442 & n16709;
  assign n16846 = ~n16710 & ~n16845;
  assign n16847 = n5240 & n12437;
  assign n16848 = n5241 & n13564;
  assign n16849 = n5853 & n12434;
  assign n16850 = n5866 & n12431;
  assign n16851 = ~n16847 & ~n16849;
  assign n16852 = ~n16850 & n16851;
  assign n16853 = ~n16848 & n16852;
  assign n16854 = pi20  & n16853;
  assign n16855 = ~pi20  & ~n16853;
  assign n16856 = ~n16854 & ~n16855;
  assign n16857 = n16846 & ~n16856;
  assign n16858 = n16458 & n16707;
  assign n16859 = ~n16708 & ~n16858;
  assign n16860 = n5240 & n12440;
  assign n16861 = n5241 & n13939;
  assign n16862 = n5853 & n12437;
  assign n16863 = n5866 & n12434;
  assign n16864 = ~n16860 & ~n16862;
  assign n16865 = ~n16863 & n16864;
  assign n16866 = ~n16861 & n16865;
  assign n16867 = pi20  & n16866;
  assign n16868 = ~pi20  & ~n16866;
  assign n16869 = ~n16867 & ~n16868;
  assign n16870 = n16859 & ~n16869;
  assign n16871 = n16474 & n16705;
  assign n16872 = ~n16706 & ~n16871;
  assign n16873 = n5240 & n12443;
  assign n16874 = n5241 & n13702;
  assign n16875 = n5853 & n12440;
  assign n16876 = n5866 & n12437;
  assign n16877 = ~n16873 & ~n16875;
  assign n16878 = ~n16876 & n16877;
  assign n16879 = ~n16874 & n16878;
  assign n16880 = pi20  & n16879;
  assign n16881 = ~pi20  & ~n16879;
  assign n16882 = ~n16880 & ~n16881;
  assign n16883 = n16872 & ~n16882;
  assign n16884 = n16701 & ~n16703;
  assign n16885 = ~n16704 & ~n16884;
  assign n16886 = n5240 & n12446;
  assign n16887 = n5241 & n14175;
  assign n16888 = n5853 & n12443;
  assign n16889 = n5866 & n12440;
  assign n16890 = ~n16886 & ~n16888;
  assign n16891 = ~n16889 & n16890;
  assign n16892 = ~n16887 & n16891;
  assign n16893 = pi20  & n16892;
  assign n16894 = ~pi20  & ~n16892;
  assign n16895 = ~n16893 & ~n16894;
  assign n16896 = n16885 & ~n16895;
  assign n16897 = n16697 & ~n16699;
  assign n16898 = ~n16700 & ~n16897;
  assign n16899 = n5240 & n12449;
  assign n16900 = n5241 & n14325;
  assign n16901 = n5853 & n12446;
  assign n16902 = n5866 & n12443;
  assign n16903 = ~n16899 & ~n16901;
  assign n16904 = ~n16902 & n16903;
  assign n16905 = ~n16900 & n16904;
  assign n16906 = pi20  & n16905;
  assign n16907 = ~pi20  & ~n16905;
  assign n16908 = ~n16906 & ~n16907;
  assign n16909 = n16898 & ~n16908;
  assign n16910 = n16693 & ~n16695;
  assign n16911 = ~n16696 & ~n16910;
  assign n16912 = n5240 & n12452;
  assign n16913 = n5241 & n14156;
  assign n16914 = n5853 & n12449;
  assign n16915 = n5866 & n12446;
  assign n16916 = ~n16912 & ~n16914;
  assign n16917 = ~n16915 & n16916;
  assign n16918 = ~n16913 & n16917;
  assign n16919 = pi20  & n16918;
  assign n16920 = ~pi20  & ~n16918;
  assign n16921 = ~n16919 & ~n16920;
  assign n16922 = n16911 & ~n16921;
  assign n16923 = n16532 & n16691;
  assign n16924 = ~n16692 & ~n16923;
  assign n16925 = n5240 & n12455;
  assign n16926 = n5241 & n14442;
  assign n16927 = n5853 & n12452;
  assign n16928 = n5866 & n12449;
  assign n16929 = ~n16925 & ~n16927;
  assign n16930 = ~n16928 & n16929;
  assign n16931 = ~n16926 & n16930;
  assign n16932 = pi20  & n16931;
  assign n16933 = ~pi20  & ~n16931;
  assign n16934 = ~n16932 & ~n16933;
  assign n16935 = n16924 & ~n16934;
  assign n16936 = n16548 & n16689;
  assign n16937 = ~n16690 & ~n16936;
  assign n16938 = n5240 & n12458;
  assign n16939 = n5241 & n14741;
  assign n16940 = n5853 & n12455;
  assign n16941 = n5866 & n12452;
  assign n16942 = ~n16938 & ~n16940;
  assign n16943 = ~n16941 & n16942;
  assign n16944 = ~n16939 & n16943;
  assign n16945 = pi20  & n16944;
  assign n16946 = ~pi20  & ~n16944;
  assign n16947 = ~n16945 & ~n16946;
  assign n16948 = n16937 & ~n16947;
  assign n16949 = n5240 & n12461;
  assign n16950 = n5241 & n14756;
  assign n16951 = n5853 & n12458;
  assign n16952 = n5866 & n12455;
  assign n16953 = ~n16949 & ~n16951;
  assign n16954 = ~n16952 & n16953;
  assign n16955 = ~n16950 & n16954;
  assign n16956 = ~pi20  & ~n16955;
  assign n16957 = pi20  & n16955;
  assign n16958 = ~n16956 & ~n16957;
  assign n16959 = n16685 & ~n16687;
  assign n16960 = ~n16688 & ~n16959;
  assign n16961 = ~n16958 & n16960;
  assign n16962 = ~n16958 & ~n16960;
  assign n16963 = n16958 & n16960;
  assign n16964 = ~n16962 & ~n16963;
  assign n16965 = n5240 & n12464;
  assign n16966 = n5241 & n14420;
  assign n16967 = n5853 & n12461;
  assign n16968 = n5866 & n12458;
  assign n16969 = ~n16965 & ~n16967;
  assign n16970 = ~n16968 & n16969;
  assign n16971 = ~n16966 & n16970;
  assign n16972 = ~pi20  & ~n16971;
  assign n16973 = pi20  & n16971;
  assign n16974 = ~n16972 & ~n16973;
  assign n16975 = ~n16680 & n16683;
  assign n16976 = n16680 & ~n16683;
  assign n16977 = ~n16975 & ~n16976;
  assign n16978 = ~n16974 & ~n16977;
  assign n16979 = n16590 & n16678;
  assign n16980 = ~n16679 & ~n16979;
  assign n16981 = n5240 & n12467;
  assign n16982 = n5241 & n14789;
  assign n16983 = n5853 & n12464;
  assign n16984 = n5866 & n12461;
  assign n16985 = ~n16981 & ~n16983;
  assign n16986 = ~n16984 & n16985;
  assign n16987 = ~n16982 & n16986;
  assign n16988 = pi20  & n16987;
  assign n16989 = ~pi20  & ~n16987;
  assign n16990 = ~n16988 & ~n16989;
  assign n16991 = n16980 & ~n16990;
  assign n16992 = n16674 & ~n16676;
  assign n16993 = ~n16677 & ~n16992;
  assign n16994 = n5240 & n12470;
  assign n16995 = n5241 & n14815;
  assign n16996 = n5853 & n12467;
  assign n16997 = n5866 & n12464;
  assign n16998 = ~n16994 & ~n16996;
  assign n16999 = ~n16997 & n16998;
  assign n17000 = ~n16995 & n16999;
  assign n17001 = pi20  & n17000;
  assign n17002 = ~pi20  & ~n17000;
  assign n17003 = ~n17001 & ~n17002;
  assign n17004 = n16993 & ~n17003;
  assign n17005 = n16621 & n16672;
  assign n17006 = ~n16673 & ~n17005;
  assign n17007 = n5240 & n12473;
  assign n17008 = n5241 & n14839;
  assign n17009 = n5853 & n12470;
  assign n17010 = n5866 & n12467;
  assign n17011 = ~n17007 & ~n17009;
  assign n17012 = ~n17010 & n17011;
  assign n17013 = ~n17008 & n17012;
  assign n17014 = pi20  & n17013;
  assign n17015 = ~pi20  & ~n17013;
  assign n17016 = ~n17014 & ~n17015;
  assign n17017 = n17006 & ~n17016;
  assign n17018 = n5240 & n12476;
  assign n17019 = n5241 & n14849;
  assign n17020 = n5853 & n12473;
  assign n17021 = n5866 & n12470;
  assign n17022 = ~n17018 & ~n17020;
  assign n17023 = ~n17021 & n17022;
  assign n17024 = ~n17019 & n17023;
  assign n17025 = ~pi20  & ~n17024;
  assign n17026 = pi20  & n17024;
  assign n17027 = ~n17025 & ~n17026;
  assign n17028 = n16668 & ~n16670;
  assign n17029 = ~n16671 & ~n17028;
  assign n17030 = ~n17027 & n17029;
  assign n17031 = ~n17027 & ~n17029;
  assign n17032 = n17027 & n17029;
  assign n17033 = ~n17031 & ~n17032;
  assign n17034 = n5240 & n12479;
  assign n17035 = n5241 & n14922;
  assign n17036 = n5853 & n12476;
  assign n17037 = n5866 & n12473;
  assign n17038 = ~n17034 & ~n17036;
  assign n17039 = ~n17037 & n17038;
  assign n17040 = ~n17035 & n17039;
  assign n17041 = pi20  & n17040;
  assign n17042 = ~pi20  & ~n17040;
  assign n17043 = ~n17041 & ~n17042;
  assign n17044 = n16656 & n16666;
  assign n17045 = ~n16667 & ~n17044;
  assign n17046 = ~n17043 & n17045;
  assign n17047 = n5240 & n12482;
  assign n17048 = n5241 & n14958;
  assign n17049 = n5853 & n12479;
  assign n17050 = n5866 & n12476;
  assign n17051 = ~n17047 & ~n17049;
  assign n17052 = ~n17050 & n17051;
  assign n17053 = ~n17048 & n17052;
  assign n17054 = ~pi20  & ~n17053;
  assign n17055 = pi20  & n17053;
  assign n17056 = ~n17054 & ~n17055;
  assign n17057 = pi23  & ~n16644;
  assign n17058 = n16651 & ~n17057;
  assign n17059 = ~n16651 & n17057;
  assign n17060 = ~n17058 & ~n17059;
  assign n17061 = ~n17056 & n17060;
  assign n17062 = ~n17056 & ~n17060;
  assign n17063 = n17056 & n17060;
  assign n17064 = ~n17062 & ~n17063;
  assign n17065 = n5240 & n12485;
  assign n17066 = n5241 & n15001;
  assign n17067 = n5853 & n12482;
  assign n17068 = n5866 & n12479;
  assign n17069 = ~n17065 & ~n17067;
  assign n17070 = ~n17068 & n17069;
  assign n17071 = ~n17066 & n17070;
  assign n17072 = pi20  & n17071;
  assign n17073 = ~pi20  & ~n17071;
  assign n17074 = ~n17072 & ~n17073;
  assign n17075 = pi23  & n16637;
  assign n17076 = ~n16642 & n17075;
  assign n17077 = n16642 & ~n17075;
  assign n17078 = ~n17076 & ~n17077;
  assign n17079 = ~n17074 & n17078;
  assign n17080 = ~n5235 & n12492;
  assign n17081 = n5853 & n12492;
  assign n17082 = n5866 & n12490;
  assign n17083 = n5241 & ~n15072;
  assign n17084 = ~n17081 & ~n17082;
  assign n17085 = ~n17083 & n17084;
  assign n17086 = pi20  & ~n17080;
  assign n17087 = n17085 & n17086;
  assign n17088 = n5240 & n12492;
  assign n17089 = n5241 & ~n15113;
  assign n17090 = n5853 & n12490;
  assign n17091 = n5866 & n12485;
  assign n17092 = ~n17088 & ~n17090;
  assign n17093 = ~n17091 & n17092;
  assign n17094 = ~n17089 & n17093;
  assign n17095 = n17087 & n17094;
  assign n17096 = n16637 & n17095;
  assign n17097 = ~n16637 & n17095;
  assign n17098 = n16637 & ~n17095;
  assign n17099 = ~n17097 & ~n17098;
  assign n17100 = n5240 & n12490;
  assign n17101 = n5241 & n15026;
  assign n17102 = n5853 & n12485;
  assign n17103 = n5866 & n12482;
  assign n17104 = ~n17100 & ~n17102;
  assign n17105 = ~n17103 & n17104;
  assign n17106 = ~n17101 & n17105;
  assign n17107 = pi20  & n17106;
  assign n17108 = ~pi20  & ~n17106;
  assign n17109 = ~n17107 & ~n17108;
  assign n17110 = ~n17099 & ~n17109;
  assign n17111 = ~n17096 & ~n17110;
  assign n17112 = n17074 & ~n17078;
  assign n17113 = ~n17079 & ~n17112;
  assign n17114 = ~n17111 & n17113;
  assign n17115 = ~n17079 & ~n17114;
  assign n17116 = ~n17064 & ~n17115;
  assign n17117 = ~n17061 & ~n17116;
  assign n17118 = n17043 & ~n17045;
  assign n17119 = ~n17046 & ~n17118;
  assign n17120 = ~n17117 & n17119;
  assign n17121 = ~n17046 & ~n17120;
  assign n17122 = ~n17033 & ~n17121;
  assign n17123 = ~n17030 & ~n17122;
  assign n17124 = n17006 & n17016;
  assign n17125 = ~n17006 & ~n17016;
  assign n17126 = ~n17124 & ~n17125;
  assign n17127 = ~n17123 & ~n17126;
  assign n17128 = ~n17017 & ~n17127;
  assign n17129 = n16993 & n17003;
  assign n17130 = ~n16993 & ~n17003;
  assign n17131 = ~n17129 & ~n17130;
  assign n17132 = ~n17128 & ~n17131;
  assign n17133 = ~n17004 & ~n17132;
  assign n17134 = ~n16980 & n16990;
  assign n17135 = ~n16991 & ~n17134;
  assign n17136 = ~n17133 & n17135;
  assign n17137 = ~n16991 & ~n17136;
  assign n17138 = n16974 & n16977;
  assign n17139 = ~n16978 & ~n17138;
  assign n17140 = ~n17137 & n17139;
  assign n17141 = ~n16978 & ~n17140;
  assign n17142 = ~n16964 & ~n17141;
  assign n17143 = ~n16961 & ~n17142;
  assign n17144 = n16937 & n16947;
  assign n17145 = ~n16937 & ~n16947;
  assign n17146 = ~n17144 & ~n17145;
  assign n17147 = ~n17143 & ~n17146;
  assign n17148 = ~n16948 & ~n17147;
  assign n17149 = n16924 & n16934;
  assign n17150 = ~n16924 & ~n16934;
  assign n17151 = ~n17149 & ~n17150;
  assign n17152 = ~n17148 & ~n17151;
  assign n17153 = ~n16935 & ~n17152;
  assign n17154 = n16911 & n16921;
  assign n17155 = ~n16911 & ~n16921;
  assign n17156 = ~n17154 & ~n17155;
  assign n17157 = ~n17153 & ~n17156;
  assign n17158 = ~n16922 & ~n17157;
  assign n17159 = n16898 & n16908;
  assign n17160 = ~n16898 & ~n16908;
  assign n17161 = ~n17159 & ~n17160;
  assign n17162 = ~n17158 & ~n17161;
  assign n17163 = ~n16909 & ~n17162;
  assign n17164 = n16885 & n16895;
  assign n17165 = ~n16885 & ~n16895;
  assign n17166 = ~n17164 & ~n17165;
  assign n17167 = ~n17163 & ~n17166;
  assign n17168 = ~n16896 & ~n17167;
  assign n17169 = n16872 & n16882;
  assign n17170 = ~n16872 & ~n16882;
  assign n17171 = ~n17169 & ~n17170;
  assign n17172 = ~n17168 & ~n17171;
  assign n17173 = ~n16883 & ~n17172;
  assign n17174 = n16859 & n16869;
  assign n17175 = ~n16859 & ~n16869;
  assign n17176 = ~n17174 & ~n17175;
  assign n17177 = ~n17173 & ~n17176;
  assign n17178 = ~n16870 & ~n17177;
  assign n17179 = n16846 & n16856;
  assign n17180 = ~n16846 & ~n16856;
  assign n17181 = ~n17179 & ~n17180;
  assign n17182 = ~n17178 & ~n17181;
  assign n17183 = ~n16857 & ~n17182;
  assign n17184 = n16833 & n16843;
  assign n17185 = ~n16833 & ~n16843;
  assign n17186 = ~n17184 & ~n17185;
  assign n17187 = ~n17183 & ~n17186;
  assign n17188 = ~n16844 & ~n17187;
  assign n17189 = ~n16820 & n16830;
  assign n17190 = ~n16831 & ~n17189;
  assign n17191 = ~n17188 & n17190;
  assign n17192 = ~n16831 & ~n17191;
  assign n17193 = ~n16720 & ~n16721;
  assign n17194 = ~n16731 & n17193;
  assign n17195 = n16731 & ~n17193;
  assign n17196 = ~n17194 & ~n17195;
  assign n17197 = ~n17192 & n17196;
  assign n17198 = n17192 & ~n17196;
  assign n17199 = n5982 & n12419;
  assign n17200 = n5983 & n12908;
  assign n17201 = n6323 & n12416;
  assign n17202 = n6336 & n12413;
  assign n17203 = ~n17199 & ~n17201;
  assign n17204 = ~n17202 & n17203;
  assign n17205 = ~n17200 & n17204;
  assign n17206 = pi17  & n17205;
  assign n17207 = ~pi17  & ~n17205;
  assign n17208 = ~n17206 & ~n17207;
  assign n17209 = ~n17198 & ~n17208;
  assign n17210 = ~n17197 & ~n17209;
  assign n17211 = n16818 & ~n17210;
  assign n17212 = ~n16818 & n17210;
  assign n17213 = n6630 & n12407;
  assign n17214 = n6631 & n13035;
  assign n17215 = n7238 & n12404;
  assign n17216 = n7262 & n12401;
  assign n17217 = ~n17213 & ~n17215;
  assign n17218 = ~n17216 & n17217;
  assign n17219 = ~n17214 & n17218;
  assign n17220 = pi14  & n17219;
  assign n17221 = ~pi14  & ~n17219;
  assign n17222 = ~n17220 & ~n17221;
  assign n17223 = ~n17212 & ~n17222;
  assign n17224 = ~n17211 & ~n17223;
  assign n17225 = n16814 & ~n17224;
  assign n17226 = ~n16814 & n17224;
  assign n17227 = n7430 & n12395;
  assign n17228 = n7431 & n13144;
  assign n17229 = n7869 & n12362;
  assign n17230 = n7895 & n12392;
  assign n17231 = ~n17227 & ~n17229;
  assign n17232 = ~n17230 & n17231;
  assign n17233 = ~n17228 & n17232;
  assign n17234 = pi11  & n17233;
  assign n17235 = ~pi11  & ~n17233;
  assign n17236 = ~n17234 & ~n17235;
  assign n17237 = ~n17226 & ~n17236;
  assign n17238 = ~n17225 & ~n17237;
  assign n17239 = ~n16810 & ~n17238;
  assign n17240 = ~n16807 & ~n17239;
  assign n17241 = ~n16768 & ~n16769;
  assign n17242 = ~n16779 & n17241;
  assign n17243 = n16779 & ~n17241;
  assign n17244 = ~n17242 & ~n17243;
  assign n17245 = ~n17240 & n17244;
  assign n17246 = n17240 & ~n17244;
  assign n17247 = n9040 & ~n12786;
  assign n17248 = n8251 & ~n13781;
  assign n17249 = n8250 & n13166;
  assign n17250 = n9016 & n13161;
  assign n17251 = ~n17247 & ~n17249;
  assign n17252 = ~n17250 & n17251;
  assign n17253 = ~n17248 & n17252;
  assign n17254 = pi8  & n17253;
  assign n17255 = ~pi8  & ~n17253;
  assign n17256 = ~n17254 & ~n17255;
  assign n17257 = ~n17246 & ~n17256;
  assign n17258 = ~n17245 & ~n17257;
  assign n17259 = n16794 & ~n17258;
  assign n17260 = ~n16794 & n17258;
  assign n17261 = ~n17259 & ~n17260;
  assign n17262 = n9040 & n13161;
  assign n17263 = n8251 & n13183;
  assign n17264 = n9016 & n13166;
  assign n17265 = n8250 & n13164;
  assign n17266 = ~n17264 & ~n17265;
  assign n17267 = ~n17262 & n17266;
  assign n17268 = ~n17263 & n17267;
  assign n17269 = pi8  & n17268;
  assign n17270 = ~pi8  & ~n17268;
  assign n17271 = ~n17269 & ~n17270;
  assign n17272 = ~n17225 & ~n17226;
  assign n17273 = ~n17236 & n17272;
  assign n17274 = n17236 & ~n17272;
  assign n17275 = ~n17273 & ~n17274;
  assign n17276 = ~n17211 & ~n17212;
  assign n17277 = ~n17222 & n17276;
  assign n17278 = n17222 & ~n17276;
  assign n17279 = ~n17277 & ~n17278;
  assign n17280 = n5982 & n12422;
  assign n17281 = n5983 & n13201;
  assign n17282 = n6323 & n12419;
  assign n17283 = n6336 & n12416;
  assign n17284 = ~n17280 & ~n17282;
  assign n17285 = ~n17283 & n17284;
  assign n17286 = ~n17281 & n17285;
  assign n17287 = ~pi17  & ~n17286;
  assign n17288 = pi17  & n17286;
  assign n17289 = ~n17287 & ~n17288;
  assign n17290 = n17188 & ~n17190;
  assign n17291 = ~n17191 & ~n17290;
  assign n17292 = ~n17289 & n17291;
  assign n17293 = ~n17289 & ~n17291;
  assign n17294 = n17289 & n17291;
  assign n17295 = ~n17293 & ~n17294;
  assign n17296 = n5982 & n12425;
  assign n17297 = n5983 & n13010;
  assign n17298 = n6323 & n12422;
  assign n17299 = n6336 & n12419;
  assign n17300 = ~n17296 & ~n17298;
  assign n17301 = ~n17299 & n17300;
  assign n17302 = ~n17297 & n17301;
  assign n17303 = ~pi17  & ~n17302;
  assign n17304 = pi17  & n17302;
  assign n17305 = ~n17303 & ~n17304;
  assign n17306 = ~n17183 & n17186;
  assign n17307 = n17183 & ~n17186;
  assign n17308 = ~n17306 & ~n17307;
  assign n17309 = ~n17305 & ~n17308;
  assign n17310 = n5982 & n12428;
  assign n17311 = n5983 & n13371;
  assign n17312 = n6323 & n12425;
  assign n17313 = n6336 & n12422;
  assign n17314 = ~n17310 & ~n17312;
  assign n17315 = ~n17313 & n17314;
  assign n17316 = ~n17311 & n17315;
  assign n17317 = ~pi17  & ~n17316;
  assign n17318 = pi17  & n17316;
  assign n17319 = ~n17317 & ~n17318;
  assign n17320 = ~n17178 & n17181;
  assign n17321 = n17178 & ~n17181;
  assign n17322 = ~n17320 & ~n17321;
  assign n17323 = ~n17319 & ~n17322;
  assign n17324 = n5982 & n12431;
  assign n17325 = n5983 & n13356;
  assign n17326 = n6323 & n12428;
  assign n17327 = n6336 & n12425;
  assign n17328 = ~n17324 & ~n17326;
  assign n17329 = ~n17327 & n17328;
  assign n17330 = ~n17325 & n17329;
  assign n17331 = ~pi17  & ~n17330;
  assign n17332 = pi17  & n17330;
  assign n17333 = ~n17331 & ~n17332;
  assign n17334 = ~n17173 & n17176;
  assign n17335 = n17173 & ~n17176;
  assign n17336 = ~n17334 & ~n17335;
  assign n17337 = ~n17333 & ~n17336;
  assign n17338 = n5982 & n12434;
  assign n17339 = n5983 & n13546;
  assign n17340 = n6323 & n12431;
  assign n17341 = n6336 & n12428;
  assign n17342 = ~n17338 & ~n17340;
  assign n17343 = ~n17341 & n17342;
  assign n17344 = ~n17339 & n17343;
  assign n17345 = ~pi17  & ~n17344;
  assign n17346 = pi17  & n17344;
  assign n17347 = ~n17345 & ~n17346;
  assign n17348 = ~n17168 & n17171;
  assign n17349 = n17168 & ~n17171;
  assign n17350 = ~n17348 & ~n17349;
  assign n17351 = ~n17347 & ~n17350;
  assign n17352 = n5982 & n12437;
  assign n17353 = n5983 & n13564;
  assign n17354 = n6323 & n12434;
  assign n17355 = n6336 & n12431;
  assign n17356 = ~n17352 & ~n17354;
  assign n17357 = ~n17355 & n17356;
  assign n17358 = ~n17353 & n17357;
  assign n17359 = ~pi17  & ~n17358;
  assign n17360 = pi17  & n17358;
  assign n17361 = ~n17359 & ~n17360;
  assign n17362 = n17163 & n17166;
  assign n17363 = ~n17167 & ~n17362;
  assign n17364 = ~n17361 & n17363;
  assign n17365 = ~n17361 & ~n17363;
  assign n17366 = n17361 & n17363;
  assign n17367 = ~n17365 & ~n17366;
  assign n17368 = n5982 & n12440;
  assign n17369 = n5983 & n13939;
  assign n17370 = n6323 & n12437;
  assign n17371 = n6336 & n12434;
  assign n17372 = ~n17368 & ~n17370;
  assign n17373 = ~n17371 & n17372;
  assign n17374 = ~n17369 & n17373;
  assign n17375 = ~pi17  & ~n17374;
  assign n17376 = pi17  & n17374;
  assign n17377 = ~n17375 & ~n17376;
  assign n17378 = n17158 & n17161;
  assign n17379 = ~n17162 & ~n17378;
  assign n17380 = ~n17377 & n17379;
  assign n17381 = ~n17377 & ~n17379;
  assign n17382 = n17377 & n17379;
  assign n17383 = ~n17381 & ~n17382;
  assign n17384 = n5982 & n12443;
  assign n17385 = n5983 & n13702;
  assign n17386 = n6323 & n12440;
  assign n17387 = n6336 & n12437;
  assign n17388 = ~n17384 & ~n17386;
  assign n17389 = ~n17387 & n17388;
  assign n17390 = ~n17385 & n17389;
  assign n17391 = ~pi17  & ~n17390;
  assign n17392 = pi17  & n17390;
  assign n17393 = ~n17391 & ~n17392;
  assign n17394 = n17153 & n17156;
  assign n17395 = ~n17157 & ~n17394;
  assign n17396 = ~n17393 & n17395;
  assign n17397 = ~n17393 & ~n17395;
  assign n17398 = n17393 & n17395;
  assign n17399 = ~n17397 & ~n17398;
  assign n17400 = n5982 & n12446;
  assign n17401 = n5983 & n14175;
  assign n17402 = n6323 & n12443;
  assign n17403 = n6336 & n12440;
  assign n17404 = ~n17400 & ~n17402;
  assign n17405 = ~n17403 & n17404;
  assign n17406 = ~n17401 & n17405;
  assign n17407 = ~pi17  & ~n17406;
  assign n17408 = pi17  & n17406;
  assign n17409 = ~n17407 & ~n17408;
  assign n17410 = ~n17148 & n17151;
  assign n17411 = n17148 & ~n17151;
  assign n17412 = ~n17410 & ~n17411;
  assign n17413 = ~n17409 & ~n17412;
  assign n17414 = n5982 & n12449;
  assign n17415 = n5983 & n14325;
  assign n17416 = n6323 & n12446;
  assign n17417 = n6336 & n12443;
  assign n17418 = ~n17414 & ~n17416;
  assign n17419 = ~n17417 & n17418;
  assign n17420 = ~n17415 & n17419;
  assign n17421 = ~pi17  & ~n17420;
  assign n17422 = pi17  & n17420;
  assign n17423 = ~n17421 & ~n17422;
  assign n17424 = ~n17143 & n17146;
  assign n17425 = n17143 & ~n17146;
  assign n17426 = ~n17424 & ~n17425;
  assign n17427 = ~n17423 & ~n17426;
  assign n17428 = n16964 & n17141;
  assign n17429 = ~n17142 & ~n17428;
  assign n17430 = n5982 & n12452;
  assign n17431 = n5983 & n14156;
  assign n17432 = n6323 & n12449;
  assign n17433 = n6336 & n12446;
  assign n17434 = ~n17430 & ~n17432;
  assign n17435 = ~n17433 & n17434;
  assign n17436 = ~n17431 & n17435;
  assign n17437 = pi17  & n17436;
  assign n17438 = ~pi17  & ~n17436;
  assign n17439 = ~n17437 & ~n17438;
  assign n17440 = n17429 & ~n17439;
  assign n17441 = n17137 & ~n17139;
  assign n17442 = ~n17140 & ~n17441;
  assign n17443 = n5982 & n12455;
  assign n17444 = n5983 & n14442;
  assign n17445 = n6323 & n12452;
  assign n17446 = n6336 & n12449;
  assign n17447 = ~n17443 & ~n17445;
  assign n17448 = ~n17446 & n17447;
  assign n17449 = ~n17444 & n17448;
  assign n17450 = pi17  & n17449;
  assign n17451 = ~pi17  & ~n17449;
  assign n17452 = ~n17450 & ~n17451;
  assign n17453 = n17442 & ~n17452;
  assign n17454 = n5982 & n12458;
  assign n17455 = n5983 & n14741;
  assign n17456 = n6323 & n12455;
  assign n17457 = n6336 & n12452;
  assign n17458 = ~n17454 & ~n17456;
  assign n17459 = ~n17457 & n17458;
  assign n17460 = ~n17455 & n17459;
  assign n17461 = ~pi17  & ~n17460;
  assign n17462 = pi17  & n17460;
  assign n17463 = ~n17461 & ~n17462;
  assign n17464 = n17133 & ~n17135;
  assign n17465 = ~n17136 & ~n17464;
  assign n17466 = ~n17463 & n17465;
  assign n17467 = ~n17463 & ~n17465;
  assign n17468 = n17463 & n17465;
  assign n17469 = ~n17467 & ~n17468;
  assign n17470 = n5982 & n12461;
  assign n17471 = n5983 & n14756;
  assign n17472 = n6323 & n12458;
  assign n17473 = n6336 & n12455;
  assign n17474 = ~n17470 & ~n17472;
  assign n17475 = ~n17473 & n17474;
  assign n17476 = ~n17471 & n17475;
  assign n17477 = ~pi17  & ~n17476;
  assign n17478 = pi17  & n17476;
  assign n17479 = ~n17477 & ~n17478;
  assign n17480 = n17128 & n17131;
  assign n17481 = ~n17132 & ~n17480;
  assign n17482 = ~n17479 & n17481;
  assign n17483 = ~n17479 & ~n17481;
  assign n17484 = n17479 & n17481;
  assign n17485 = ~n17483 & ~n17484;
  assign n17486 = n5982 & n12464;
  assign n17487 = n5983 & n14420;
  assign n17488 = n6323 & n12461;
  assign n17489 = n6336 & n12458;
  assign n17490 = ~n17486 & ~n17488;
  assign n17491 = ~n17489 & n17490;
  assign n17492 = ~n17487 & n17491;
  assign n17493 = ~pi17  & ~n17492;
  assign n17494 = pi17  & n17492;
  assign n17495 = ~n17493 & ~n17494;
  assign n17496 = ~n17123 & n17126;
  assign n17497 = n17123 & ~n17126;
  assign n17498 = ~n17496 & ~n17497;
  assign n17499 = ~n17495 & ~n17498;
  assign n17500 = n17033 & n17121;
  assign n17501 = ~n17122 & ~n17500;
  assign n17502 = n5982 & n12467;
  assign n17503 = n5983 & n14789;
  assign n17504 = n6323 & n12464;
  assign n17505 = n6336 & n12461;
  assign n17506 = ~n17502 & ~n17504;
  assign n17507 = ~n17505 & n17506;
  assign n17508 = ~n17503 & n17507;
  assign n17509 = pi17  & n17508;
  assign n17510 = ~pi17  & ~n17508;
  assign n17511 = ~n17509 & ~n17510;
  assign n17512 = n17501 & ~n17511;
  assign n17513 = n17117 & ~n17119;
  assign n17514 = ~n17120 & ~n17513;
  assign n17515 = n5982 & n12470;
  assign n17516 = n5983 & n14815;
  assign n17517 = n6323 & n12467;
  assign n17518 = n6336 & n12464;
  assign n17519 = ~n17515 & ~n17517;
  assign n17520 = ~n17518 & n17519;
  assign n17521 = ~n17516 & n17520;
  assign n17522 = pi17  & n17521;
  assign n17523 = ~pi17  & ~n17521;
  assign n17524 = ~n17522 & ~n17523;
  assign n17525 = n17514 & ~n17524;
  assign n17526 = n17064 & n17115;
  assign n17527 = ~n17116 & ~n17526;
  assign n17528 = n5982 & n12473;
  assign n17529 = n5983 & n14839;
  assign n17530 = n6323 & n12470;
  assign n17531 = n6336 & n12467;
  assign n17532 = ~n17528 & ~n17530;
  assign n17533 = ~n17531 & n17532;
  assign n17534 = ~n17529 & n17533;
  assign n17535 = pi17  & n17534;
  assign n17536 = ~pi17  & ~n17534;
  assign n17537 = ~n17535 & ~n17536;
  assign n17538 = n17527 & ~n17537;
  assign n17539 = n5982 & n12476;
  assign n17540 = n5983 & n14849;
  assign n17541 = n6323 & n12473;
  assign n17542 = n6336 & n12470;
  assign n17543 = ~n17539 & ~n17541;
  assign n17544 = ~n17542 & n17543;
  assign n17545 = ~n17540 & n17544;
  assign n17546 = ~pi17  & ~n17545;
  assign n17547 = pi17  & n17545;
  assign n17548 = ~n17546 & ~n17547;
  assign n17549 = n17111 & ~n17113;
  assign n17550 = ~n17114 & ~n17549;
  assign n17551 = ~n17548 & n17550;
  assign n17552 = ~n17548 & ~n17550;
  assign n17553 = n17548 & n17550;
  assign n17554 = ~n17552 & ~n17553;
  assign n17555 = n5982 & n12479;
  assign n17556 = n5983 & n14922;
  assign n17557 = n6323 & n12476;
  assign n17558 = n6336 & n12473;
  assign n17559 = ~n17555 & ~n17557;
  assign n17560 = ~n17558 & n17559;
  assign n17561 = ~n17556 & n17560;
  assign n17562 = pi17  & n17561;
  assign n17563 = ~pi17  & ~n17561;
  assign n17564 = ~n17562 & ~n17563;
  assign n17565 = n17099 & n17109;
  assign n17566 = ~n17110 & ~n17565;
  assign n17567 = ~n17564 & n17566;
  assign n17568 = n5982 & n12482;
  assign n17569 = n5983 & n14958;
  assign n17570 = n6323 & n12479;
  assign n17571 = n6336 & n12476;
  assign n17572 = ~n17568 & ~n17570;
  assign n17573 = ~n17571 & n17572;
  assign n17574 = ~n17569 & n17573;
  assign n17575 = ~pi17  & ~n17574;
  assign n17576 = pi17  & n17574;
  assign n17577 = ~n17575 & ~n17576;
  assign n17578 = pi20  & ~n17087;
  assign n17579 = n17094 & ~n17578;
  assign n17580 = ~n17094 & n17578;
  assign n17581 = ~n17579 & ~n17580;
  assign n17582 = ~n17577 & n17581;
  assign n17583 = ~n17577 & ~n17581;
  assign n17584 = n17577 & n17581;
  assign n17585 = ~n17583 & ~n17584;
  assign n17586 = n5982 & n12485;
  assign n17587 = n5983 & n15001;
  assign n17588 = n6323 & n12482;
  assign n17589 = n6336 & n12479;
  assign n17590 = ~n17586 & ~n17588;
  assign n17591 = ~n17589 & n17590;
  assign n17592 = ~n17587 & n17591;
  assign n17593 = pi17  & n17592;
  assign n17594 = ~pi17  & ~n17592;
  assign n17595 = ~n17593 & ~n17594;
  assign n17596 = pi20  & n17080;
  assign n17597 = ~n17085 & n17596;
  assign n17598 = n17085 & ~n17596;
  assign n17599 = ~n17597 & ~n17598;
  assign n17600 = ~n17595 & n17599;
  assign n17601 = ~n5980 & n12492;
  assign n17602 = n6323 & n12492;
  assign n17603 = n6336 & n12490;
  assign n17604 = n5983 & ~n15072;
  assign n17605 = ~n17602 & ~n17603;
  assign n17606 = ~n17604 & n17605;
  assign n17607 = pi17  & ~n17601;
  assign n17608 = n17606 & n17607;
  assign n17609 = n5982 & n12492;
  assign n17610 = n5983 & ~n15113;
  assign n17611 = n6323 & n12490;
  assign n17612 = n6336 & n12485;
  assign n17613 = ~n17609 & ~n17611;
  assign n17614 = ~n17612 & n17613;
  assign n17615 = ~n17610 & n17614;
  assign n17616 = n17608 & n17615;
  assign n17617 = n17080 & n17616;
  assign n17618 = ~n17080 & n17616;
  assign n17619 = n17080 & ~n17616;
  assign n17620 = ~n17618 & ~n17619;
  assign n17621 = n5982 & n12490;
  assign n17622 = n5983 & n15026;
  assign n17623 = n6323 & n12485;
  assign n17624 = n6336 & n12482;
  assign n17625 = ~n17621 & ~n17623;
  assign n17626 = ~n17624 & n17625;
  assign n17627 = ~n17622 & n17626;
  assign n17628 = pi17  & n17627;
  assign n17629 = ~pi17  & ~n17627;
  assign n17630 = ~n17628 & ~n17629;
  assign n17631 = ~n17620 & ~n17630;
  assign n17632 = ~n17617 & ~n17631;
  assign n17633 = n17595 & ~n17599;
  assign n17634 = ~n17600 & ~n17633;
  assign n17635 = ~n17632 & n17634;
  assign n17636 = ~n17600 & ~n17635;
  assign n17637 = ~n17585 & ~n17636;
  assign n17638 = ~n17582 & ~n17637;
  assign n17639 = n17564 & ~n17566;
  assign n17640 = ~n17567 & ~n17639;
  assign n17641 = ~n17638 & n17640;
  assign n17642 = ~n17567 & ~n17641;
  assign n17643 = ~n17554 & ~n17642;
  assign n17644 = ~n17551 & ~n17643;
  assign n17645 = n17527 & n17537;
  assign n17646 = ~n17527 & ~n17537;
  assign n17647 = ~n17645 & ~n17646;
  assign n17648 = ~n17644 & ~n17647;
  assign n17649 = ~n17538 & ~n17648;
  assign n17650 = n17514 & n17524;
  assign n17651 = ~n17514 & ~n17524;
  assign n17652 = ~n17650 & ~n17651;
  assign n17653 = ~n17649 & ~n17652;
  assign n17654 = ~n17525 & ~n17653;
  assign n17655 = ~n17501 & n17511;
  assign n17656 = ~n17512 & ~n17655;
  assign n17657 = ~n17654 & n17656;
  assign n17658 = ~n17512 & ~n17657;
  assign n17659 = n17495 & n17498;
  assign n17660 = ~n17499 & ~n17659;
  assign n17661 = ~n17658 & n17660;
  assign n17662 = ~n17499 & ~n17661;
  assign n17663 = ~n17485 & ~n17662;
  assign n17664 = ~n17482 & ~n17663;
  assign n17665 = ~n17469 & ~n17664;
  assign n17666 = ~n17466 & ~n17665;
  assign n17667 = n17442 & n17452;
  assign n17668 = ~n17442 & ~n17452;
  assign n17669 = ~n17667 & ~n17668;
  assign n17670 = ~n17666 & ~n17669;
  assign n17671 = ~n17453 & ~n17670;
  assign n17672 = ~n17429 & n17439;
  assign n17673 = ~n17440 & ~n17672;
  assign n17674 = ~n17671 & n17673;
  assign n17675 = ~n17440 & ~n17674;
  assign n17676 = n17423 & n17426;
  assign n17677 = ~n17427 & ~n17676;
  assign n17678 = ~n17675 & n17677;
  assign n17679 = ~n17427 & ~n17678;
  assign n17680 = n17409 & n17412;
  assign n17681 = ~n17413 & ~n17680;
  assign n17682 = ~n17679 & n17681;
  assign n17683 = ~n17413 & ~n17682;
  assign n17684 = ~n17399 & ~n17683;
  assign n17685 = ~n17396 & ~n17684;
  assign n17686 = ~n17383 & ~n17685;
  assign n17687 = ~n17380 & ~n17686;
  assign n17688 = ~n17367 & ~n17687;
  assign n17689 = ~n17364 & ~n17688;
  assign n17690 = n17347 & n17350;
  assign n17691 = ~n17351 & ~n17690;
  assign n17692 = ~n17689 & n17691;
  assign n17693 = ~n17351 & ~n17692;
  assign n17694 = n17333 & n17336;
  assign n17695 = ~n17337 & ~n17694;
  assign n17696 = ~n17693 & n17695;
  assign n17697 = ~n17337 & ~n17696;
  assign n17698 = n17319 & n17322;
  assign n17699 = ~n17323 & ~n17698;
  assign n17700 = ~n17697 & n17699;
  assign n17701 = ~n17323 & ~n17700;
  assign n17702 = n17305 & n17308;
  assign n17703 = ~n17309 & ~n17702;
  assign n17704 = ~n17701 & n17703;
  assign n17705 = ~n17309 & ~n17704;
  assign n17706 = ~n17295 & ~n17705;
  assign n17707 = ~n17292 & ~n17706;
  assign n17708 = ~n17197 & ~n17198;
  assign n17709 = ~n17208 & n17708;
  assign n17710 = n17208 & ~n17708;
  assign n17711 = ~n17709 & ~n17710;
  assign n17712 = ~n17707 & n17711;
  assign n17713 = n17707 & ~n17711;
  assign n17714 = n6630 & n12410;
  assign n17715 = n6631 & n13093;
  assign n17716 = n7238 & n12407;
  assign n17717 = n7262 & n12404;
  assign n17718 = ~n17714 & ~n17716;
  assign n17719 = ~n17717 & n17718;
  assign n17720 = ~n17715 & n17719;
  assign n17721 = pi14  & n17720;
  assign n17722 = ~pi14  & ~n17720;
  assign n17723 = ~n17721 & ~n17722;
  assign n17724 = ~n17713 & ~n17723;
  assign n17725 = ~n17712 & ~n17724;
  assign n17726 = n17279 & ~n17725;
  assign n17727 = ~n17279 & n17725;
  assign n17728 = n7430 & n12398;
  assign n17729 = n7431 & n13245;
  assign n17730 = n7869 & n12395;
  assign n17731 = n7895 & n12362;
  assign n17732 = ~n17728 & ~n17730;
  assign n17733 = ~n17731 & n17732;
  assign n17734 = ~n17729 & n17733;
  assign n17735 = pi11  & n17734;
  assign n17736 = ~pi11  & ~n17734;
  assign n17737 = ~n17735 & ~n17736;
  assign n17738 = ~n17727 & ~n17737;
  assign n17739 = ~n17726 & ~n17738;
  assign n17740 = n17275 & ~n17739;
  assign n17741 = ~n17275 & n17739;
  assign n17742 = n8250 & n12646;
  assign n17743 = n8251 & n13261;
  assign n17744 = n9016 & n13164;
  assign n17745 = n9040 & n13166;
  assign n17746 = ~n17742 & ~n17744;
  assign n17747 = ~n17745 & n17746;
  assign n17748 = ~n17743 & n17747;
  assign n17749 = pi8  & n17748;
  assign n17750 = ~pi8  & ~n17748;
  assign n17751 = ~n17749 & ~n17750;
  assign n17752 = ~n17741 & ~n17751;
  assign n17753 = ~n17740 & ~n17752;
  assign n17754 = ~n17271 & ~n17753;
  assign n17755 = n17271 & ~n17753;
  assign n17756 = ~n17271 & n17753;
  assign n17757 = ~n17755 & ~n17756;
  assign n17758 = n16810 & n17238;
  assign n17759 = ~n17239 & ~n17758;
  assign n17760 = ~n17757 & n17759;
  assign n17761 = ~n17754 & ~n17760;
  assign n17762 = ~n17245 & ~n17246;
  assign n17763 = ~n17256 & n17762;
  assign n17764 = n17256 & ~n17762;
  assign n17765 = ~n17763 & ~n17764;
  assign n17766 = ~n17761 & n17765;
  assign n17767 = n17761 & n17765;
  assign n17768 = ~n17761 & ~n17765;
  assign n17769 = ~n17767 & ~n17768;
  assign n17770 = n17757 & ~n17759;
  assign n17771 = ~n17760 & ~n17770;
  assign n17772 = n9491 & ~n13280;
  assign n17773 = n74 & ~n13160;
  assign n17774 = n14143 & ~n17773;
  assign n17775 = ~n12786 & ~n17774;
  assign n17776 = ~n17772 & ~n17775;
  assign n17777 = pi5  & n17776;
  assign n17778 = ~pi5  & ~n17776;
  assign n17779 = ~n17777 & ~n17778;
  assign n17780 = ~n17726 & ~n17727;
  assign n17781 = ~n17737 & n17780;
  assign n17782 = n17737 & ~n17780;
  assign n17783 = ~n17781 & ~n17782;
  assign n17784 = n17295 & n17705;
  assign n17785 = ~n17706 & ~n17784;
  assign n17786 = n6630 & n12413;
  assign n17787 = n6631 & n12891;
  assign n17788 = n7238 & n12410;
  assign n17789 = n7262 & n12407;
  assign n17790 = ~n17786 & ~n17788;
  assign n17791 = ~n17789 & n17790;
  assign n17792 = ~n17787 & n17791;
  assign n17793 = pi14  & n17792;
  assign n17794 = ~pi14  & ~n17792;
  assign n17795 = ~n17793 & ~n17794;
  assign n17796 = n17785 & ~n17795;
  assign n17797 = n17701 & ~n17703;
  assign n17798 = ~n17704 & ~n17797;
  assign n17799 = n6630 & n12416;
  assign n17800 = n6631 & n12843;
  assign n17801 = n7238 & n12413;
  assign n17802 = n7262 & n12410;
  assign n17803 = ~n17799 & ~n17801;
  assign n17804 = ~n17802 & n17803;
  assign n17805 = ~n17800 & n17804;
  assign n17806 = pi14  & n17805;
  assign n17807 = ~pi14  & ~n17805;
  assign n17808 = ~n17806 & ~n17807;
  assign n17809 = n17798 & ~n17808;
  assign n17810 = n17697 & ~n17699;
  assign n17811 = ~n17700 & ~n17810;
  assign n17812 = n6630 & n12419;
  assign n17813 = n6631 & n12908;
  assign n17814 = n7238 & n12416;
  assign n17815 = n7262 & n12413;
  assign n17816 = ~n17812 & ~n17814;
  assign n17817 = ~n17815 & n17816;
  assign n17818 = ~n17813 & n17817;
  assign n17819 = pi14  & n17818;
  assign n17820 = ~pi14  & ~n17818;
  assign n17821 = ~n17819 & ~n17820;
  assign n17822 = n17811 & ~n17821;
  assign n17823 = n17693 & ~n17695;
  assign n17824 = ~n17696 & ~n17823;
  assign n17825 = n6630 & n12422;
  assign n17826 = n6631 & n13201;
  assign n17827 = n7238 & n12419;
  assign n17828 = n7262 & n12416;
  assign n17829 = ~n17825 & ~n17827;
  assign n17830 = ~n17828 & n17829;
  assign n17831 = ~n17826 & n17830;
  assign n17832 = pi14  & n17831;
  assign n17833 = ~pi14  & ~n17831;
  assign n17834 = ~n17832 & ~n17833;
  assign n17835 = n17824 & ~n17834;
  assign n17836 = n17689 & ~n17691;
  assign n17837 = ~n17692 & ~n17836;
  assign n17838 = n6630 & n12425;
  assign n17839 = n6631 & n13010;
  assign n17840 = n7238 & n12422;
  assign n17841 = n7262 & n12419;
  assign n17842 = ~n17838 & ~n17840;
  assign n17843 = ~n17841 & n17842;
  assign n17844 = ~n17839 & n17843;
  assign n17845 = pi14  & n17844;
  assign n17846 = ~pi14  & ~n17844;
  assign n17847 = ~n17845 & ~n17846;
  assign n17848 = n17837 & ~n17847;
  assign n17849 = n17367 & n17687;
  assign n17850 = ~n17688 & ~n17849;
  assign n17851 = n6630 & n12428;
  assign n17852 = n6631 & n13371;
  assign n17853 = n7238 & n12425;
  assign n17854 = n7262 & n12422;
  assign n17855 = ~n17851 & ~n17853;
  assign n17856 = ~n17854 & n17855;
  assign n17857 = ~n17852 & n17856;
  assign n17858 = pi14  & n17857;
  assign n17859 = ~pi14  & ~n17857;
  assign n17860 = ~n17858 & ~n17859;
  assign n17861 = n17850 & ~n17860;
  assign n17862 = n17383 & n17685;
  assign n17863 = ~n17686 & ~n17862;
  assign n17864 = n6630 & n12431;
  assign n17865 = n6631 & n13356;
  assign n17866 = n7238 & n12428;
  assign n17867 = n7262 & n12425;
  assign n17868 = ~n17864 & ~n17866;
  assign n17869 = ~n17867 & n17868;
  assign n17870 = ~n17865 & n17869;
  assign n17871 = pi14  & n17870;
  assign n17872 = ~pi14  & ~n17870;
  assign n17873 = ~n17871 & ~n17872;
  assign n17874 = n17863 & ~n17873;
  assign n17875 = n17399 & n17683;
  assign n17876 = ~n17684 & ~n17875;
  assign n17877 = n6630 & n12434;
  assign n17878 = n6631 & n13546;
  assign n17879 = n7238 & n12431;
  assign n17880 = n7262 & n12428;
  assign n17881 = ~n17877 & ~n17879;
  assign n17882 = ~n17880 & n17881;
  assign n17883 = ~n17878 & n17882;
  assign n17884 = pi14  & n17883;
  assign n17885 = ~pi14  & ~n17883;
  assign n17886 = ~n17884 & ~n17885;
  assign n17887 = n17876 & ~n17886;
  assign n17888 = n17679 & ~n17681;
  assign n17889 = ~n17682 & ~n17888;
  assign n17890 = n6630 & n12437;
  assign n17891 = n6631 & n13564;
  assign n17892 = n7238 & n12434;
  assign n17893 = n7262 & n12431;
  assign n17894 = ~n17890 & ~n17892;
  assign n17895 = ~n17893 & n17894;
  assign n17896 = ~n17891 & n17895;
  assign n17897 = pi14  & n17896;
  assign n17898 = ~pi14  & ~n17896;
  assign n17899 = ~n17897 & ~n17898;
  assign n17900 = n17889 & ~n17899;
  assign n17901 = n17675 & ~n17677;
  assign n17902 = ~n17678 & ~n17901;
  assign n17903 = n6630 & n12440;
  assign n17904 = n6631 & n13939;
  assign n17905 = n7238 & n12437;
  assign n17906 = n7262 & n12434;
  assign n17907 = ~n17903 & ~n17905;
  assign n17908 = ~n17906 & n17907;
  assign n17909 = ~n17904 & n17908;
  assign n17910 = pi14  & n17909;
  assign n17911 = ~pi14  & ~n17909;
  assign n17912 = ~n17910 & ~n17911;
  assign n17913 = n17902 & ~n17912;
  assign n17914 = n6630 & n12443;
  assign n17915 = n6631 & n13702;
  assign n17916 = n7238 & n12440;
  assign n17917 = n7262 & n12437;
  assign n17918 = ~n17914 & ~n17916;
  assign n17919 = ~n17917 & n17918;
  assign n17920 = ~n17915 & n17919;
  assign n17921 = ~pi14  & ~n17920;
  assign n17922 = pi14  & n17920;
  assign n17923 = ~n17921 & ~n17922;
  assign n17924 = n17671 & ~n17673;
  assign n17925 = ~n17674 & ~n17924;
  assign n17926 = ~n17923 & n17925;
  assign n17927 = ~n17923 & ~n17925;
  assign n17928 = n17923 & n17925;
  assign n17929 = ~n17927 & ~n17928;
  assign n17930 = n6630 & n12446;
  assign n17931 = n6631 & n14175;
  assign n17932 = n7238 & n12443;
  assign n17933 = n7262 & n12440;
  assign n17934 = ~n17930 & ~n17932;
  assign n17935 = ~n17933 & n17934;
  assign n17936 = ~n17931 & n17935;
  assign n17937 = ~pi14  & ~n17936;
  assign n17938 = pi14  & n17936;
  assign n17939 = ~n17937 & ~n17938;
  assign n17940 = n17666 & n17669;
  assign n17941 = ~n17670 & ~n17940;
  assign n17942 = ~n17939 & n17941;
  assign n17943 = ~n17939 & ~n17941;
  assign n17944 = n17939 & n17941;
  assign n17945 = ~n17943 & ~n17944;
  assign n17946 = n17469 & n17664;
  assign n17947 = ~n17665 & ~n17946;
  assign n17948 = n6630 & n12449;
  assign n17949 = n6631 & n14325;
  assign n17950 = n7238 & n12446;
  assign n17951 = n7262 & n12443;
  assign n17952 = ~n17948 & ~n17950;
  assign n17953 = ~n17951 & n17952;
  assign n17954 = ~n17949 & n17953;
  assign n17955 = pi14  & n17954;
  assign n17956 = ~pi14  & ~n17954;
  assign n17957 = ~n17955 & ~n17956;
  assign n17958 = n17947 & ~n17957;
  assign n17959 = n17485 & n17662;
  assign n17960 = ~n17663 & ~n17959;
  assign n17961 = n6630 & n12452;
  assign n17962 = n6631 & n14156;
  assign n17963 = n7238 & n12449;
  assign n17964 = n7262 & n12446;
  assign n17965 = ~n17961 & ~n17963;
  assign n17966 = ~n17964 & n17965;
  assign n17967 = ~n17962 & n17966;
  assign n17968 = pi14  & n17967;
  assign n17969 = ~pi14  & ~n17967;
  assign n17970 = ~n17968 & ~n17969;
  assign n17971 = n17960 & ~n17970;
  assign n17972 = n17658 & ~n17660;
  assign n17973 = ~n17661 & ~n17972;
  assign n17974 = n6630 & n12455;
  assign n17975 = n6631 & n14442;
  assign n17976 = n7238 & n12452;
  assign n17977 = n7262 & n12449;
  assign n17978 = ~n17974 & ~n17976;
  assign n17979 = ~n17977 & n17978;
  assign n17980 = ~n17975 & n17979;
  assign n17981 = pi14  & n17980;
  assign n17982 = ~pi14  & ~n17980;
  assign n17983 = ~n17981 & ~n17982;
  assign n17984 = n17973 & ~n17983;
  assign n17985 = n6630 & n12458;
  assign n17986 = n6631 & n14741;
  assign n17987 = n7238 & n12455;
  assign n17988 = n7262 & n12452;
  assign n17989 = ~n17985 & ~n17987;
  assign n17990 = ~n17988 & n17989;
  assign n17991 = ~n17986 & n17990;
  assign n17992 = ~pi14  & ~n17991;
  assign n17993 = pi14  & n17991;
  assign n17994 = ~n17992 & ~n17993;
  assign n17995 = n17654 & ~n17656;
  assign n17996 = ~n17657 & ~n17995;
  assign n17997 = ~n17994 & n17996;
  assign n17998 = ~n17994 & ~n17996;
  assign n17999 = n17994 & n17996;
  assign n18000 = ~n17998 & ~n17999;
  assign n18001 = n6630 & n12461;
  assign n18002 = n6631 & n14756;
  assign n18003 = n7238 & n12458;
  assign n18004 = n7262 & n12455;
  assign n18005 = ~n18001 & ~n18003;
  assign n18006 = ~n18004 & n18005;
  assign n18007 = ~n18002 & n18006;
  assign n18008 = ~pi14  & ~n18007;
  assign n18009 = pi14  & n18007;
  assign n18010 = ~n18008 & ~n18009;
  assign n18011 = n17649 & n17652;
  assign n18012 = ~n17653 & ~n18011;
  assign n18013 = ~n18010 & n18012;
  assign n18014 = ~n18010 & ~n18012;
  assign n18015 = n18010 & n18012;
  assign n18016 = ~n18014 & ~n18015;
  assign n18017 = n6630 & n12464;
  assign n18018 = n6631 & n14420;
  assign n18019 = n7238 & n12461;
  assign n18020 = n7262 & n12458;
  assign n18021 = ~n18017 & ~n18019;
  assign n18022 = ~n18020 & n18021;
  assign n18023 = ~n18018 & n18022;
  assign n18024 = ~pi14  & ~n18023;
  assign n18025 = pi14  & n18023;
  assign n18026 = ~n18024 & ~n18025;
  assign n18027 = ~n17644 & n17647;
  assign n18028 = n17644 & ~n17647;
  assign n18029 = ~n18027 & ~n18028;
  assign n18030 = ~n18026 & ~n18029;
  assign n18031 = n17554 & n17642;
  assign n18032 = ~n17643 & ~n18031;
  assign n18033 = n6630 & n12467;
  assign n18034 = n6631 & n14789;
  assign n18035 = n7238 & n12464;
  assign n18036 = n7262 & n12461;
  assign n18037 = ~n18033 & ~n18035;
  assign n18038 = ~n18036 & n18037;
  assign n18039 = ~n18034 & n18038;
  assign n18040 = pi14  & n18039;
  assign n18041 = ~pi14  & ~n18039;
  assign n18042 = ~n18040 & ~n18041;
  assign n18043 = n18032 & ~n18042;
  assign n18044 = n17638 & ~n17640;
  assign n18045 = ~n17641 & ~n18044;
  assign n18046 = n6630 & n12470;
  assign n18047 = n6631 & n14815;
  assign n18048 = n7238 & n12467;
  assign n18049 = n7262 & n12464;
  assign n18050 = ~n18046 & ~n18048;
  assign n18051 = ~n18049 & n18050;
  assign n18052 = ~n18047 & n18051;
  assign n18053 = pi14  & n18052;
  assign n18054 = ~pi14  & ~n18052;
  assign n18055 = ~n18053 & ~n18054;
  assign n18056 = n18045 & ~n18055;
  assign n18057 = n17585 & n17636;
  assign n18058 = ~n17637 & ~n18057;
  assign n18059 = n6630 & n12473;
  assign n18060 = n6631 & n14839;
  assign n18061 = n7238 & n12470;
  assign n18062 = n7262 & n12467;
  assign n18063 = ~n18059 & ~n18061;
  assign n18064 = ~n18062 & n18063;
  assign n18065 = ~n18060 & n18064;
  assign n18066 = pi14  & n18065;
  assign n18067 = ~pi14  & ~n18065;
  assign n18068 = ~n18066 & ~n18067;
  assign n18069 = n18058 & ~n18068;
  assign n18070 = n6630 & n12476;
  assign n18071 = n6631 & n14849;
  assign n18072 = n7238 & n12473;
  assign n18073 = n7262 & n12470;
  assign n18074 = ~n18070 & ~n18072;
  assign n18075 = ~n18073 & n18074;
  assign n18076 = ~n18071 & n18075;
  assign n18077 = ~pi14  & ~n18076;
  assign n18078 = pi14  & n18076;
  assign n18079 = ~n18077 & ~n18078;
  assign n18080 = n17632 & ~n17634;
  assign n18081 = ~n17635 & ~n18080;
  assign n18082 = ~n18079 & n18081;
  assign n18083 = ~n18079 & ~n18081;
  assign n18084 = n18079 & n18081;
  assign n18085 = ~n18083 & ~n18084;
  assign n18086 = n6630 & n12479;
  assign n18087 = n6631 & n14922;
  assign n18088 = n7238 & n12476;
  assign n18089 = n7262 & n12473;
  assign n18090 = ~n18086 & ~n18088;
  assign n18091 = ~n18089 & n18090;
  assign n18092 = ~n18087 & n18091;
  assign n18093 = pi14  & n18092;
  assign n18094 = ~pi14  & ~n18092;
  assign n18095 = ~n18093 & ~n18094;
  assign n18096 = n17620 & n17630;
  assign n18097 = ~n17631 & ~n18096;
  assign n18098 = ~n18095 & n18097;
  assign n18099 = n6630 & n12482;
  assign n18100 = n6631 & n14958;
  assign n18101 = n7238 & n12479;
  assign n18102 = n7262 & n12476;
  assign n18103 = ~n18099 & ~n18101;
  assign n18104 = ~n18102 & n18103;
  assign n18105 = ~n18100 & n18104;
  assign n18106 = ~pi14  & ~n18105;
  assign n18107 = pi14  & n18105;
  assign n18108 = ~n18106 & ~n18107;
  assign n18109 = pi17  & ~n17608;
  assign n18110 = n17615 & ~n18109;
  assign n18111 = ~n17615 & n18109;
  assign n18112 = ~n18110 & ~n18111;
  assign n18113 = ~n18108 & n18112;
  assign n18114 = ~n18108 & ~n18112;
  assign n18115 = n18108 & n18112;
  assign n18116 = ~n18114 & ~n18115;
  assign n18117 = n6630 & n12485;
  assign n18118 = n6631 & n15001;
  assign n18119 = n7238 & n12482;
  assign n18120 = n7262 & n12479;
  assign n18121 = ~n18117 & ~n18119;
  assign n18122 = ~n18120 & n18121;
  assign n18123 = ~n18118 & n18122;
  assign n18124 = pi14  & n18123;
  assign n18125 = ~pi14  & ~n18123;
  assign n18126 = ~n18124 & ~n18125;
  assign n18127 = pi17  & n17601;
  assign n18128 = ~n17606 & n18127;
  assign n18129 = n17606 & ~n18127;
  assign n18130 = ~n18128 & ~n18129;
  assign n18131 = ~n18126 & n18130;
  assign n18132 = ~n6628 & n12492;
  assign n18133 = n7238 & n12492;
  assign n18134 = n7262 & n12490;
  assign n18135 = n6631 & ~n15072;
  assign n18136 = ~n18133 & ~n18134;
  assign n18137 = ~n18135 & n18136;
  assign n18138 = pi14  & ~n18132;
  assign n18139 = n18137 & n18138;
  assign n18140 = n6630 & n12492;
  assign n18141 = n6631 & ~n15113;
  assign n18142 = n7238 & n12490;
  assign n18143 = n7262 & n12485;
  assign n18144 = ~n18140 & ~n18142;
  assign n18145 = ~n18143 & n18144;
  assign n18146 = ~n18141 & n18145;
  assign n18147 = n18139 & n18146;
  assign n18148 = n17601 & n18147;
  assign n18149 = ~n17601 & n18147;
  assign n18150 = n17601 & ~n18147;
  assign n18151 = ~n18149 & ~n18150;
  assign n18152 = n6630 & n12490;
  assign n18153 = n6631 & n15026;
  assign n18154 = n7238 & n12485;
  assign n18155 = n7262 & n12482;
  assign n18156 = ~n18152 & ~n18154;
  assign n18157 = ~n18155 & n18156;
  assign n18158 = ~n18153 & n18157;
  assign n18159 = pi14  & n18158;
  assign n18160 = ~pi14  & ~n18158;
  assign n18161 = ~n18159 & ~n18160;
  assign n18162 = ~n18151 & ~n18161;
  assign n18163 = ~n18148 & ~n18162;
  assign n18164 = n18126 & ~n18130;
  assign n18165 = ~n18131 & ~n18164;
  assign n18166 = ~n18163 & n18165;
  assign n18167 = ~n18131 & ~n18166;
  assign n18168 = ~n18116 & ~n18167;
  assign n18169 = ~n18113 & ~n18168;
  assign n18170 = n18095 & ~n18097;
  assign n18171 = ~n18098 & ~n18170;
  assign n18172 = ~n18169 & n18171;
  assign n18173 = ~n18098 & ~n18172;
  assign n18174 = ~n18085 & ~n18173;
  assign n18175 = ~n18082 & ~n18174;
  assign n18176 = n18058 & n18068;
  assign n18177 = ~n18058 & ~n18068;
  assign n18178 = ~n18176 & ~n18177;
  assign n18179 = ~n18175 & ~n18178;
  assign n18180 = ~n18069 & ~n18179;
  assign n18181 = n18045 & n18055;
  assign n18182 = ~n18045 & ~n18055;
  assign n18183 = ~n18181 & ~n18182;
  assign n18184 = ~n18180 & ~n18183;
  assign n18185 = ~n18056 & ~n18184;
  assign n18186 = ~n18032 & n18042;
  assign n18187 = ~n18043 & ~n18186;
  assign n18188 = ~n18185 & n18187;
  assign n18189 = ~n18043 & ~n18188;
  assign n18190 = n18026 & n18029;
  assign n18191 = ~n18030 & ~n18190;
  assign n18192 = ~n18189 & n18191;
  assign n18193 = ~n18030 & ~n18192;
  assign n18194 = ~n18016 & ~n18193;
  assign n18195 = ~n18013 & ~n18194;
  assign n18196 = ~n18000 & ~n18195;
  assign n18197 = ~n17997 & ~n18196;
  assign n18198 = n17973 & n17983;
  assign n18199 = ~n17973 & ~n17983;
  assign n18200 = ~n18198 & ~n18199;
  assign n18201 = ~n18197 & ~n18200;
  assign n18202 = ~n17984 & ~n18201;
  assign n18203 = n17960 & n17970;
  assign n18204 = ~n17960 & ~n17970;
  assign n18205 = ~n18203 & ~n18204;
  assign n18206 = ~n18202 & ~n18205;
  assign n18207 = ~n17971 & ~n18206;
  assign n18208 = ~n17947 & n17957;
  assign n18209 = ~n17958 & ~n18208;
  assign n18210 = ~n18207 & n18209;
  assign n18211 = ~n17958 & ~n18210;
  assign n18212 = ~n17945 & ~n18211;
  assign n18213 = ~n17942 & ~n18212;
  assign n18214 = ~n17929 & ~n18213;
  assign n18215 = ~n17926 & ~n18214;
  assign n18216 = n17902 & n17912;
  assign n18217 = ~n17902 & ~n17912;
  assign n18218 = ~n18216 & ~n18217;
  assign n18219 = ~n18215 & ~n18218;
  assign n18220 = ~n17913 & ~n18219;
  assign n18221 = n17889 & n17899;
  assign n18222 = ~n17889 & ~n17899;
  assign n18223 = ~n18221 & ~n18222;
  assign n18224 = ~n18220 & ~n18223;
  assign n18225 = ~n17900 & ~n18224;
  assign n18226 = n17876 & n17886;
  assign n18227 = ~n17876 & ~n17886;
  assign n18228 = ~n18226 & ~n18227;
  assign n18229 = ~n18225 & ~n18228;
  assign n18230 = ~n17887 & ~n18229;
  assign n18231 = n17863 & n17873;
  assign n18232 = ~n17863 & ~n17873;
  assign n18233 = ~n18231 & ~n18232;
  assign n18234 = ~n18230 & ~n18233;
  assign n18235 = ~n17874 & ~n18234;
  assign n18236 = n17850 & n17860;
  assign n18237 = ~n17850 & ~n17860;
  assign n18238 = ~n18236 & ~n18237;
  assign n18239 = ~n18235 & ~n18238;
  assign n18240 = ~n17861 & ~n18239;
  assign n18241 = n17837 & n17847;
  assign n18242 = ~n17837 & ~n17847;
  assign n18243 = ~n18241 & ~n18242;
  assign n18244 = ~n18240 & ~n18243;
  assign n18245 = ~n17848 & ~n18244;
  assign n18246 = n17824 & n17834;
  assign n18247 = ~n17824 & ~n17834;
  assign n18248 = ~n18246 & ~n18247;
  assign n18249 = ~n18245 & ~n18248;
  assign n18250 = ~n17835 & ~n18249;
  assign n18251 = n17811 & n17821;
  assign n18252 = ~n17811 & ~n17821;
  assign n18253 = ~n18251 & ~n18252;
  assign n18254 = ~n18250 & ~n18253;
  assign n18255 = ~n17822 & ~n18254;
  assign n18256 = n17798 & n17808;
  assign n18257 = ~n17798 & ~n17808;
  assign n18258 = ~n18256 & ~n18257;
  assign n18259 = ~n18255 & ~n18258;
  assign n18260 = ~n17809 & ~n18259;
  assign n18261 = ~n17785 & n17795;
  assign n18262 = ~n17796 & ~n18261;
  assign n18263 = ~n18260 & n18262;
  assign n18264 = ~n17796 & ~n18263;
  assign n18265 = ~n17712 & ~n17713;
  assign n18266 = ~n17723 & n18265;
  assign n18267 = n17723 & ~n18265;
  assign n18268 = ~n18266 & ~n18267;
  assign n18269 = ~n18264 & n18268;
  assign n18270 = n18264 & ~n18268;
  assign n18271 = n7430 & n12401;
  assign n18272 = n7431 & n13108;
  assign n18273 = n7869 & n12398;
  assign n18274 = n7895 & n12395;
  assign n18275 = ~n18271 & ~n18273;
  assign n18276 = ~n18274 & n18275;
  assign n18277 = ~n18272 & n18276;
  assign n18278 = pi11  & n18277;
  assign n18279 = ~pi11  & ~n18277;
  assign n18280 = ~n18278 & ~n18279;
  assign n18281 = ~n18270 & ~n18280;
  assign n18282 = ~n18269 & ~n18281;
  assign n18283 = n17783 & ~n18282;
  assign n18284 = ~n17783 & n18282;
  assign n18285 = n8250 & n12392;
  assign n18286 = n8251 & n13421;
  assign n18287 = n9016 & n12646;
  assign n18288 = n9040 & n13164;
  assign n18289 = ~n18285 & ~n18287;
  assign n18290 = ~n18288 & n18289;
  assign n18291 = ~n18286 & n18290;
  assign n18292 = pi8  & n18291;
  assign n18293 = ~pi8  & ~n18291;
  assign n18294 = ~n18292 & ~n18293;
  assign n18295 = ~n18284 & ~n18294;
  assign n18296 = ~n18283 & ~n18295;
  assign n18297 = ~n17779 & ~n18296;
  assign n18298 = n17779 & n18296;
  assign n18299 = ~n17740 & ~n17741;
  assign n18300 = ~n17751 & n18299;
  assign n18301 = n17751 & ~n18299;
  assign n18302 = ~n18300 & ~n18301;
  assign n18303 = ~n18298 & n18302;
  assign n18304 = ~n18297 & ~n18303;
  assign n18305 = n17771 & ~n18304;
  assign n18306 = ~n18297 & ~n18298;
  assign n18307 = n18302 & n18306;
  assign n18308 = ~n18302 & ~n18306;
  assign n18309 = ~n18307 & ~n18308;
  assign n18310 = ~n18283 & ~n18284;
  assign n18311 = ~n18294 & n18310;
  assign n18312 = n18294 & ~n18310;
  assign n18313 = ~n18311 & ~n18312;
  assign n18314 = n7430 & n12404;
  assign n18315 = n7431 & n13128;
  assign n18316 = n7869 & n12401;
  assign n18317 = n7895 & n12398;
  assign n18318 = ~n18314 & ~n18316;
  assign n18319 = ~n18317 & n18318;
  assign n18320 = ~n18315 & n18319;
  assign n18321 = ~pi11  & ~n18320;
  assign n18322 = pi11  & n18320;
  assign n18323 = ~n18321 & ~n18322;
  assign n18324 = n18260 & ~n18262;
  assign n18325 = ~n18263 & ~n18324;
  assign n18326 = ~n18323 & n18325;
  assign n18327 = ~n18323 & ~n18325;
  assign n18328 = n18323 & n18325;
  assign n18329 = ~n18327 & ~n18328;
  assign n18330 = n7430 & n12407;
  assign n18331 = n7431 & n13035;
  assign n18332 = n7869 & n12404;
  assign n18333 = n7895 & n12401;
  assign n18334 = ~n18330 & ~n18332;
  assign n18335 = ~n18333 & n18334;
  assign n18336 = ~n18331 & n18335;
  assign n18337 = ~pi11  & ~n18336;
  assign n18338 = pi11  & n18336;
  assign n18339 = ~n18337 & ~n18338;
  assign n18340 = n18255 & n18258;
  assign n18341 = ~n18259 & ~n18340;
  assign n18342 = ~n18339 & n18341;
  assign n18343 = ~n18339 & ~n18341;
  assign n18344 = n18339 & n18341;
  assign n18345 = ~n18343 & ~n18344;
  assign n18346 = n7430 & n12410;
  assign n18347 = n7431 & n13093;
  assign n18348 = n7869 & n12407;
  assign n18349 = n7895 & n12404;
  assign n18350 = ~n18346 & ~n18348;
  assign n18351 = ~n18349 & n18350;
  assign n18352 = ~n18347 & n18351;
  assign n18353 = ~pi11  & ~n18352;
  assign n18354 = pi11  & n18352;
  assign n18355 = ~n18353 & ~n18354;
  assign n18356 = n18250 & n18253;
  assign n18357 = ~n18254 & ~n18356;
  assign n18358 = ~n18355 & n18357;
  assign n18359 = ~n18355 & ~n18357;
  assign n18360 = n18355 & n18357;
  assign n18361 = ~n18359 & ~n18360;
  assign n18362 = n7430 & n12413;
  assign n18363 = n7431 & n12891;
  assign n18364 = n7869 & n12410;
  assign n18365 = n7895 & n12407;
  assign n18366 = ~n18362 & ~n18364;
  assign n18367 = ~n18365 & n18366;
  assign n18368 = ~n18363 & n18367;
  assign n18369 = ~pi11  & ~n18368;
  assign n18370 = pi11  & n18368;
  assign n18371 = ~n18369 & ~n18370;
  assign n18372 = n18245 & n18248;
  assign n18373 = ~n18249 & ~n18372;
  assign n18374 = ~n18371 & n18373;
  assign n18375 = ~n18371 & ~n18373;
  assign n18376 = n18371 & n18373;
  assign n18377 = ~n18375 & ~n18376;
  assign n18378 = n7430 & n12416;
  assign n18379 = n7431 & n12843;
  assign n18380 = n7869 & n12413;
  assign n18381 = n7895 & n12410;
  assign n18382 = ~n18378 & ~n18380;
  assign n18383 = ~n18381 & n18382;
  assign n18384 = ~n18379 & n18383;
  assign n18385 = ~pi11  & ~n18384;
  assign n18386 = pi11  & n18384;
  assign n18387 = ~n18385 & ~n18386;
  assign n18388 = n18240 & n18243;
  assign n18389 = ~n18244 & ~n18388;
  assign n18390 = ~n18387 & n18389;
  assign n18391 = ~n18387 & ~n18389;
  assign n18392 = n18387 & n18389;
  assign n18393 = ~n18391 & ~n18392;
  assign n18394 = n7430 & n12419;
  assign n18395 = n7431 & n12908;
  assign n18396 = n7869 & n12416;
  assign n18397 = n7895 & n12413;
  assign n18398 = ~n18394 & ~n18396;
  assign n18399 = ~n18397 & n18398;
  assign n18400 = ~n18395 & n18399;
  assign n18401 = ~pi11  & ~n18400;
  assign n18402 = pi11  & n18400;
  assign n18403 = ~n18401 & ~n18402;
  assign n18404 = ~n18235 & n18238;
  assign n18405 = n18235 & ~n18238;
  assign n18406 = ~n18404 & ~n18405;
  assign n18407 = ~n18403 & ~n18406;
  assign n18408 = n7430 & n12422;
  assign n18409 = n7431 & n13201;
  assign n18410 = n7869 & n12419;
  assign n18411 = n7895 & n12416;
  assign n18412 = ~n18408 & ~n18410;
  assign n18413 = ~n18411 & n18412;
  assign n18414 = ~n18409 & n18413;
  assign n18415 = ~pi11  & ~n18414;
  assign n18416 = pi11  & n18414;
  assign n18417 = ~n18415 & ~n18416;
  assign n18418 = ~n18230 & n18233;
  assign n18419 = n18230 & ~n18233;
  assign n18420 = ~n18418 & ~n18419;
  assign n18421 = ~n18417 & ~n18420;
  assign n18422 = n7430 & n12425;
  assign n18423 = n7431 & n13010;
  assign n18424 = n7869 & n12422;
  assign n18425 = n7895 & n12419;
  assign n18426 = ~n18422 & ~n18424;
  assign n18427 = ~n18425 & n18426;
  assign n18428 = ~n18423 & n18427;
  assign n18429 = ~pi11  & ~n18428;
  assign n18430 = pi11  & n18428;
  assign n18431 = ~n18429 & ~n18430;
  assign n18432 = ~n18225 & n18228;
  assign n18433 = n18225 & ~n18228;
  assign n18434 = ~n18432 & ~n18433;
  assign n18435 = ~n18431 & ~n18434;
  assign n18436 = n7430 & n12428;
  assign n18437 = n7431 & n13371;
  assign n18438 = n7869 & n12425;
  assign n18439 = n7895 & n12422;
  assign n18440 = ~n18436 & ~n18438;
  assign n18441 = ~n18439 & n18440;
  assign n18442 = ~n18437 & n18441;
  assign n18443 = ~pi11  & ~n18442;
  assign n18444 = pi11  & n18442;
  assign n18445 = ~n18443 & ~n18444;
  assign n18446 = n18220 & n18223;
  assign n18447 = ~n18224 & ~n18446;
  assign n18448 = ~n18445 & n18447;
  assign n18449 = ~n18445 & ~n18447;
  assign n18450 = n18445 & n18447;
  assign n18451 = ~n18449 & ~n18450;
  assign n18452 = n7430 & n12431;
  assign n18453 = n7431 & n13356;
  assign n18454 = n7869 & n12428;
  assign n18455 = n7895 & n12425;
  assign n18456 = ~n18452 & ~n18454;
  assign n18457 = ~n18455 & n18456;
  assign n18458 = ~n18453 & n18457;
  assign n18459 = ~pi11  & ~n18458;
  assign n18460 = pi11  & n18458;
  assign n18461 = ~n18459 & ~n18460;
  assign n18462 = n18215 & n18218;
  assign n18463 = ~n18219 & ~n18462;
  assign n18464 = ~n18461 & n18463;
  assign n18465 = ~n18461 & ~n18463;
  assign n18466 = n18461 & n18463;
  assign n18467 = ~n18465 & ~n18466;
  assign n18468 = n17929 & n18213;
  assign n18469 = ~n18214 & ~n18468;
  assign n18470 = n7430 & n12434;
  assign n18471 = n7431 & n13546;
  assign n18472 = n7869 & n12431;
  assign n18473 = n7895 & n12428;
  assign n18474 = ~n18470 & ~n18472;
  assign n18475 = ~n18473 & n18474;
  assign n18476 = ~n18471 & n18475;
  assign n18477 = pi11  & n18476;
  assign n18478 = ~pi11  & ~n18476;
  assign n18479 = ~n18477 & ~n18478;
  assign n18480 = n18469 & ~n18479;
  assign n18481 = n17945 & n18211;
  assign n18482 = ~n18212 & ~n18481;
  assign n18483 = n7430 & n12437;
  assign n18484 = n7431 & n13564;
  assign n18485 = n7869 & n12434;
  assign n18486 = n7895 & n12431;
  assign n18487 = ~n18483 & ~n18485;
  assign n18488 = ~n18486 & n18487;
  assign n18489 = ~n18484 & n18488;
  assign n18490 = pi11  & n18489;
  assign n18491 = ~pi11  & ~n18489;
  assign n18492 = ~n18490 & ~n18491;
  assign n18493 = n18482 & ~n18492;
  assign n18494 = n7430 & n12440;
  assign n18495 = n7431 & n13939;
  assign n18496 = n7869 & n12437;
  assign n18497 = n7895 & n12434;
  assign n18498 = ~n18494 & ~n18496;
  assign n18499 = ~n18497 & n18498;
  assign n18500 = ~n18495 & n18499;
  assign n18501 = ~pi11  & ~n18500;
  assign n18502 = pi11  & n18500;
  assign n18503 = ~n18501 & ~n18502;
  assign n18504 = n18207 & ~n18209;
  assign n18505 = ~n18210 & ~n18504;
  assign n18506 = ~n18503 & n18505;
  assign n18507 = ~n18503 & ~n18505;
  assign n18508 = n18503 & n18505;
  assign n18509 = ~n18507 & ~n18508;
  assign n18510 = n7430 & n12443;
  assign n18511 = n7431 & n13702;
  assign n18512 = n7869 & n12440;
  assign n18513 = n7895 & n12437;
  assign n18514 = ~n18510 & ~n18512;
  assign n18515 = ~n18513 & n18514;
  assign n18516 = ~n18511 & n18515;
  assign n18517 = ~pi11  & ~n18516;
  assign n18518 = pi11  & n18516;
  assign n18519 = ~n18517 & ~n18518;
  assign n18520 = ~n18202 & n18205;
  assign n18521 = n18202 & ~n18205;
  assign n18522 = ~n18520 & ~n18521;
  assign n18523 = ~n18519 & ~n18522;
  assign n18524 = n7430 & n12446;
  assign n18525 = n7431 & n14175;
  assign n18526 = n7869 & n12443;
  assign n18527 = n7895 & n12440;
  assign n18528 = ~n18524 & ~n18526;
  assign n18529 = ~n18527 & n18528;
  assign n18530 = ~n18525 & n18529;
  assign n18531 = ~pi11  & ~n18530;
  assign n18532 = pi11  & n18530;
  assign n18533 = ~n18531 & ~n18532;
  assign n18534 = n18197 & n18200;
  assign n18535 = ~n18201 & ~n18534;
  assign n18536 = ~n18533 & n18535;
  assign n18537 = ~n18533 & ~n18535;
  assign n18538 = n18533 & n18535;
  assign n18539 = ~n18537 & ~n18538;
  assign n18540 = n18000 & n18195;
  assign n18541 = ~n18196 & ~n18540;
  assign n18542 = n7430 & n12449;
  assign n18543 = n7431 & n14325;
  assign n18544 = n7869 & n12446;
  assign n18545 = n7895 & n12443;
  assign n18546 = ~n18542 & ~n18544;
  assign n18547 = ~n18545 & n18546;
  assign n18548 = ~n18543 & n18547;
  assign n18549 = pi11  & n18548;
  assign n18550 = ~pi11  & ~n18548;
  assign n18551 = ~n18549 & ~n18550;
  assign n18552 = n18541 & ~n18551;
  assign n18553 = n18016 & n18193;
  assign n18554 = ~n18194 & ~n18553;
  assign n18555 = n7430 & n12452;
  assign n18556 = n7431 & n14156;
  assign n18557 = n7869 & n12449;
  assign n18558 = n7895 & n12446;
  assign n18559 = ~n18555 & ~n18557;
  assign n18560 = ~n18558 & n18559;
  assign n18561 = ~n18556 & n18560;
  assign n18562 = pi11  & n18561;
  assign n18563 = ~pi11  & ~n18561;
  assign n18564 = ~n18562 & ~n18563;
  assign n18565 = n18554 & ~n18564;
  assign n18566 = n18189 & ~n18191;
  assign n18567 = ~n18192 & ~n18566;
  assign n18568 = n7430 & n12455;
  assign n18569 = n7431 & n14442;
  assign n18570 = n7869 & n12452;
  assign n18571 = n7895 & n12449;
  assign n18572 = ~n18568 & ~n18570;
  assign n18573 = ~n18571 & n18572;
  assign n18574 = ~n18569 & n18573;
  assign n18575 = pi11  & n18574;
  assign n18576 = ~pi11  & ~n18574;
  assign n18577 = ~n18575 & ~n18576;
  assign n18578 = n18567 & ~n18577;
  assign n18579 = n7430 & n12458;
  assign n18580 = n7431 & n14741;
  assign n18581 = n7869 & n12455;
  assign n18582 = n7895 & n12452;
  assign n18583 = ~n18579 & ~n18581;
  assign n18584 = ~n18582 & n18583;
  assign n18585 = ~n18580 & n18584;
  assign n18586 = ~pi11  & ~n18585;
  assign n18587 = pi11  & n18585;
  assign n18588 = ~n18586 & ~n18587;
  assign n18589 = n18185 & ~n18187;
  assign n18590 = ~n18188 & ~n18589;
  assign n18591 = ~n18588 & n18590;
  assign n18592 = ~n18588 & ~n18590;
  assign n18593 = n18588 & n18590;
  assign n18594 = ~n18592 & ~n18593;
  assign n18595 = n7430 & n12461;
  assign n18596 = n7431 & n14756;
  assign n18597 = n7869 & n12458;
  assign n18598 = n7895 & n12455;
  assign n18599 = ~n18595 & ~n18597;
  assign n18600 = ~n18598 & n18599;
  assign n18601 = ~n18596 & n18600;
  assign n18602 = ~pi11  & ~n18601;
  assign n18603 = pi11  & n18601;
  assign n18604 = ~n18602 & ~n18603;
  assign n18605 = n18180 & n18183;
  assign n18606 = ~n18184 & ~n18605;
  assign n18607 = ~n18604 & n18606;
  assign n18608 = ~n18604 & ~n18606;
  assign n18609 = n18604 & n18606;
  assign n18610 = ~n18608 & ~n18609;
  assign n18611 = n7430 & n12464;
  assign n18612 = n7431 & n14420;
  assign n18613 = n7869 & n12461;
  assign n18614 = n7895 & n12458;
  assign n18615 = ~n18611 & ~n18613;
  assign n18616 = ~n18614 & n18615;
  assign n18617 = ~n18612 & n18616;
  assign n18618 = ~pi11  & ~n18617;
  assign n18619 = pi11  & n18617;
  assign n18620 = ~n18618 & ~n18619;
  assign n18621 = ~n18175 & n18178;
  assign n18622 = n18175 & ~n18178;
  assign n18623 = ~n18621 & ~n18622;
  assign n18624 = ~n18620 & ~n18623;
  assign n18625 = n18085 & n18173;
  assign n18626 = ~n18174 & ~n18625;
  assign n18627 = n7430 & n12467;
  assign n18628 = n7431 & n14789;
  assign n18629 = n7869 & n12464;
  assign n18630 = n7895 & n12461;
  assign n18631 = ~n18627 & ~n18629;
  assign n18632 = ~n18630 & n18631;
  assign n18633 = ~n18628 & n18632;
  assign n18634 = pi11  & n18633;
  assign n18635 = ~pi11  & ~n18633;
  assign n18636 = ~n18634 & ~n18635;
  assign n18637 = n18626 & ~n18636;
  assign n18638 = n18169 & ~n18171;
  assign n18639 = ~n18172 & ~n18638;
  assign n18640 = n7430 & n12470;
  assign n18641 = n7431 & n14815;
  assign n18642 = n7869 & n12467;
  assign n18643 = n7895 & n12464;
  assign n18644 = ~n18640 & ~n18642;
  assign n18645 = ~n18643 & n18644;
  assign n18646 = ~n18641 & n18645;
  assign n18647 = pi11  & n18646;
  assign n18648 = ~pi11  & ~n18646;
  assign n18649 = ~n18647 & ~n18648;
  assign n18650 = n18639 & ~n18649;
  assign n18651 = n18116 & n18167;
  assign n18652 = ~n18168 & ~n18651;
  assign n18653 = n7430 & n12473;
  assign n18654 = n7431 & n14839;
  assign n18655 = n7869 & n12470;
  assign n18656 = n7895 & n12467;
  assign n18657 = ~n18653 & ~n18655;
  assign n18658 = ~n18656 & n18657;
  assign n18659 = ~n18654 & n18658;
  assign n18660 = pi11  & n18659;
  assign n18661 = ~pi11  & ~n18659;
  assign n18662 = ~n18660 & ~n18661;
  assign n18663 = n18652 & ~n18662;
  assign n18664 = n7430 & n12476;
  assign n18665 = n7431 & n14849;
  assign n18666 = n7869 & n12473;
  assign n18667 = n7895 & n12470;
  assign n18668 = ~n18664 & ~n18666;
  assign n18669 = ~n18667 & n18668;
  assign n18670 = ~n18665 & n18669;
  assign n18671 = ~pi11  & ~n18670;
  assign n18672 = pi11  & n18670;
  assign n18673 = ~n18671 & ~n18672;
  assign n18674 = n18163 & ~n18165;
  assign n18675 = ~n18166 & ~n18674;
  assign n18676 = ~n18673 & n18675;
  assign n18677 = ~n18673 & ~n18675;
  assign n18678 = n18673 & n18675;
  assign n18679 = ~n18677 & ~n18678;
  assign n18680 = n7430 & n12479;
  assign n18681 = n7431 & n14922;
  assign n18682 = n7869 & n12476;
  assign n18683 = n7895 & n12473;
  assign n18684 = ~n18680 & ~n18682;
  assign n18685 = ~n18683 & n18684;
  assign n18686 = ~n18681 & n18685;
  assign n18687 = pi11  & n18686;
  assign n18688 = ~pi11  & ~n18686;
  assign n18689 = ~n18687 & ~n18688;
  assign n18690 = n18151 & n18161;
  assign n18691 = ~n18162 & ~n18690;
  assign n18692 = ~n18689 & n18691;
  assign n18693 = n7430 & n12482;
  assign n18694 = n7431 & n14958;
  assign n18695 = n7869 & n12479;
  assign n18696 = n7895 & n12476;
  assign n18697 = ~n18693 & ~n18695;
  assign n18698 = ~n18696 & n18697;
  assign n18699 = ~n18694 & n18698;
  assign n18700 = ~pi11  & ~n18699;
  assign n18701 = pi11  & n18699;
  assign n18702 = ~n18700 & ~n18701;
  assign n18703 = pi14  & ~n18139;
  assign n18704 = n18146 & ~n18703;
  assign n18705 = ~n18146 & n18703;
  assign n18706 = ~n18704 & ~n18705;
  assign n18707 = ~n18702 & n18706;
  assign n18708 = ~n18702 & ~n18706;
  assign n18709 = n18702 & n18706;
  assign n18710 = ~n18708 & ~n18709;
  assign n18711 = n7430 & n12485;
  assign n18712 = n7431 & n15001;
  assign n18713 = n7869 & n12482;
  assign n18714 = n7895 & n12479;
  assign n18715 = ~n18711 & ~n18713;
  assign n18716 = ~n18714 & n18715;
  assign n18717 = ~n18712 & n18716;
  assign n18718 = pi11  & n18717;
  assign n18719 = ~pi11  & ~n18717;
  assign n18720 = ~n18718 & ~n18719;
  assign n18721 = pi14  & n18132;
  assign n18722 = ~n18137 & n18721;
  assign n18723 = n18137 & ~n18721;
  assign n18724 = ~n18722 & ~n18723;
  assign n18725 = ~n18720 & n18724;
  assign n18726 = ~n7425 & n12492;
  assign n18727 = n7869 & n12492;
  assign n18728 = n7895 & n12490;
  assign n18729 = n7431 & ~n15072;
  assign n18730 = ~n18727 & ~n18728;
  assign n18731 = ~n18729 & n18730;
  assign n18732 = pi11  & ~n18726;
  assign n18733 = n18731 & n18732;
  assign n18734 = n7430 & n12492;
  assign n18735 = n7431 & ~n15113;
  assign n18736 = n7869 & n12490;
  assign n18737 = n7895 & n12485;
  assign n18738 = ~n18734 & ~n18736;
  assign n18739 = ~n18737 & n18738;
  assign n18740 = ~n18735 & n18739;
  assign n18741 = n18733 & n18740;
  assign n18742 = n18132 & n18741;
  assign n18743 = ~n18132 & n18741;
  assign n18744 = n18132 & ~n18741;
  assign n18745 = ~n18743 & ~n18744;
  assign n18746 = n7430 & n12490;
  assign n18747 = n7431 & n15026;
  assign n18748 = n7869 & n12485;
  assign n18749 = n7895 & n12482;
  assign n18750 = ~n18746 & ~n18748;
  assign n18751 = ~n18749 & n18750;
  assign n18752 = ~n18747 & n18751;
  assign n18753 = pi11  & n18752;
  assign n18754 = ~pi11  & ~n18752;
  assign n18755 = ~n18753 & ~n18754;
  assign n18756 = ~n18745 & ~n18755;
  assign n18757 = ~n18742 & ~n18756;
  assign n18758 = n18720 & ~n18724;
  assign n18759 = ~n18725 & ~n18758;
  assign n18760 = ~n18757 & n18759;
  assign n18761 = ~n18725 & ~n18760;
  assign n18762 = ~n18710 & ~n18761;
  assign n18763 = ~n18707 & ~n18762;
  assign n18764 = n18689 & ~n18691;
  assign n18765 = ~n18692 & ~n18764;
  assign n18766 = ~n18763 & n18765;
  assign n18767 = ~n18692 & ~n18766;
  assign n18768 = ~n18679 & ~n18767;
  assign n18769 = ~n18676 & ~n18768;
  assign n18770 = n18652 & n18662;
  assign n18771 = ~n18652 & ~n18662;
  assign n18772 = ~n18770 & ~n18771;
  assign n18773 = ~n18769 & ~n18772;
  assign n18774 = ~n18663 & ~n18773;
  assign n18775 = n18639 & n18649;
  assign n18776 = ~n18639 & ~n18649;
  assign n18777 = ~n18775 & ~n18776;
  assign n18778 = ~n18774 & ~n18777;
  assign n18779 = ~n18650 & ~n18778;
  assign n18780 = ~n18626 & n18636;
  assign n18781 = ~n18637 & ~n18780;
  assign n18782 = ~n18779 & n18781;
  assign n18783 = ~n18637 & ~n18782;
  assign n18784 = n18620 & n18623;
  assign n18785 = ~n18624 & ~n18784;
  assign n18786 = ~n18783 & n18785;
  assign n18787 = ~n18624 & ~n18786;
  assign n18788 = ~n18610 & ~n18787;
  assign n18789 = ~n18607 & ~n18788;
  assign n18790 = ~n18594 & ~n18789;
  assign n18791 = ~n18591 & ~n18790;
  assign n18792 = n18567 & n18577;
  assign n18793 = ~n18567 & ~n18577;
  assign n18794 = ~n18792 & ~n18793;
  assign n18795 = ~n18791 & ~n18794;
  assign n18796 = ~n18578 & ~n18795;
  assign n18797 = n18554 & n18564;
  assign n18798 = ~n18554 & ~n18564;
  assign n18799 = ~n18797 & ~n18798;
  assign n18800 = ~n18796 & ~n18799;
  assign n18801 = ~n18565 & ~n18800;
  assign n18802 = ~n18541 & n18551;
  assign n18803 = ~n18552 & ~n18802;
  assign n18804 = ~n18801 & n18803;
  assign n18805 = ~n18552 & ~n18804;
  assign n18806 = ~n18539 & ~n18805;
  assign n18807 = ~n18536 & ~n18806;
  assign n18808 = n18519 & n18522;
  assign n18809 = ~n18523 & ~n18808;
  assign n18810 = ~n18807 & n18809;
  assign n18811 = ~n18523 & ~n18810;
  assign n18812 = ~n18509 & ~n18811;
  assign n18813 = ~n18506 & ~n18812;
  assign n18814 = n18482 & n18492;
  assign n18815 = ~n18482 & ~n18492;
  assign n18816 = ~n18814 & ~n18815;
  assign n18817 = ~n18813 & ~n18816;
  assign n18818 = ~n18493 & ~n18817;
  assign n18819 = ~n18469 & n18479;
  assign n18820 = ~n18480 & ~n18819;
  assign n18821 = ~n18818 & n18820;
  assign n18822 = ~n18480 & ~n18821;
  assign n18823 = ~n18467 & ~n18822;
  assign n18824 = ~n18464 & ~n18823;
  assign n18825 = ~n18451 & ~n18824;
  assign n18826 = ~n18448 & ~n18825;
  assign n18827 = n18431 & n18434;
  assign n18828 = ~n18435 & ~n18827;
  assign n18829 = ~n18826 & n18828;
  assign n18830 = ~n18435 & ~n18829;
  assign n18831 = n18417 & n18420;
  assign n18832 = ~n18421 & ~n18831;
  assign n18833 = ~n18830 & n18832;
  assign n18834 = ~n18421 & ~n18833;
  assign n18835 = n18403 & n18406;
  assign n18836 = ~n18407 & ~n18835;
  assign n18837 = ~n18834 & n18836;
  assign n18838 = ~n18407 & ~n18837;
  assign n18839 = ~n18393 & ~n18838;
  assign n18840 = ~n18390 & ~n18839;
  assign n18841 = ~n18377 & ~n18840;
  assign n18842 = ~n18374 & ~n18841;
  assign n18843 = ~n18361 & ~n18842;
  assign n18844 = ~n18358 & ~n18843;
  assign n18845 = ~n18345 & ~n18844;
  assign n18846 = ~n18342 & ~n18845;
  assign n18847 = ~n18329 & ~n18846;
  assign n18848 = ~n18326 & ~n18847;
  assign n18849 = ~n18269 & ~n18270;
  assign n18850 = ~n18280 & n18849;
  assign n18851 = n18280 & ~n18849;
  assign n18852 = ~n18850 & ~n18851;
  assign n18853 = ~n18848 & n18852;
  assign n18854 = n18848 & ~n18852;
  assign n18855 = n8250 & n12362;
  assign n18856 = n8251 & n12652;
  assign n18857 = n9016 & n12392;
  assign n18858 = n9040 & n12646;
  assign n18859 = ~n18855 & ~n18857;
  assign n18860 = ~n18858 & n18859;
  assign n18861 = ~n18856 & n18860;
  assign n18862 = pi8  & n18861;
  assign n18863 = ~pi8  & ~n18861;
  assign n18864 = ~n18862 & ~n18863;
  assign n18865 = ~n18854 & ~n18864;
  assign n18866 = ~n18853 & ~n18865;
  assign n18867 = n18313 & ~n18866;
  assign n18868 = ~n18313 & n18866;
  assign n18869 = n11031 & ~n12786;
  assign n18870 = n9491 & ~n13781;
  assign n18871 = n75 & n13166;
  assign n18872 = n10469 & n13161;
  assign n18873 = ~n18869 & ~n18871;
  assign n18874 = ~n18872 & n18873;
  assign n18875 = ~n18870 & n18874;
  assign n18876 = pi5  & n18875;
  assign n18877 = ~pi5  & ~n18875;
  assign n18878 = ~n18876 & ~n18877;
  assign n18879 = ~n18868 & ~n18878;
  assign n18880 = ~n18867 & ~n18879;
  assign n18881 = n18309 & ~n18880;
  assign n18882 = ~n18309 & n18880;
  assign n18883 = ~n18881 & ~n18882;
  assign n18884 = ~n18867 & ~n18868;
  assign n18885 = ~n18878 & n18884;
  assign n18886 = n18878 & ~n18884;
  assign n18887 = ~n18885 & ~n18886;
  assign n18888 = n18329 & n18846;
  assign n18889 = ~n18847 & ~n18888;
  assign n18890 = n8250 & n12395;
  assign n18891 = n8251 & n13144;
  assign n18892 = n9016 & n12362;
  assign n18893 = n9040 & n12392;
  assign n18894 = ~n18890 & ~n18892;
  assign n18895 = ~n18893 & n18894;
  assign n18896 = ~n18891 & n18895;
  assign n18897 = pi8  & n18896;
  assign n18898 = ~pi8  & ~n18896;
  assign n18899 = ~n18897 & ~n18898;
  assign n18900 = n18889 & ~n18899;
  assign n18901 = n18345 & n18844;
  assign n18902 = ~n18845 & ~n18901;
  assign n18903 = n8250 & n12398;
  assign n18904 = n8251 & n13245;
  assign n18905 = n9016 & n12395;
  assign n18906 = n9040 & n12362;
  assign n18907 = ~n18903 & ~n18905;
  assign n18908 = ~n18906 & n18907;
  assign n18909 = ~n18904 & n18908;
  assign n18910 = pi8  & n18909;
  assign n18911 = ~pi8  & ~n18909;
  assign n18912 = ~n18910 & ~n18911;
  assign n18913 = n18902 & ~n18912;
  assign n18914 = n18361 & n18842;
  assign n18915 = ~n18843 & ~n18914;
  assign n18916 = n8250 & n12401;
  assign n18917 = n8251 & n13108;
  assign n18918 = n9016 & n12398;
  assign n18919 = n9040 & n12395;
  assign n18920 = ~n18916 & ~n18918;
  assign n18921 = ~n18919 & n18920;
  assign n18922 = ~n18917 & n18921;
  assign n18923 = pi8  & n18922;
  assign n18924 = ~pi8  & ~n18922;
  assign n18925 = ~n18923 & ~n18924;
  assign n18926 = n18915 & ~n18925;
  assign n18927 = n18377 & n18840;
  assign n18928 = ~n18841 & ~n18927;
  assign n18929 = n8250 & n12404;
  assign n18930 = n8251 & n13128;
  assign n18931 = n9016 & n12401;
  assign n18932 = n9040 & n12398;
  assign n18933 = ~n18929 & ~n18931;
  assign n18934 = ~n18932 & n18933;
  assign n18935 = ~n18930 & n18934;
  assign n18936 = pi8  & n18935;
  assign n18937 = ~pi8  & ~n18935;
  assign n18938 = ~n18936 & ~n18937;
  assign n18939 = n18928 & ~n18938;
  assign n18940 = n18393 & n18838;
  assign n18941 = ~n18839 & ~n18940;
  assign n18942 = n8250 & n12407;
  assign n18943 = n8251 & n13035;
  assign n18944 = n9016 & n12404;
  assign n18945 = n9040 & n12401;
  assign n18946 = ~n18942 & ~n18944;
  assign n18947 = ~n18945 & n18946;
  assign n18948 = ~n18943 & n18947;
  assign n18949 = pi8  & n18948;
  assign n18950 = ~pi8  & ~n18948;
  assign n18951 = ~n18949 & ~n18950;
  assign n18952 = n18941 & ~n18951;
  assign n18953 = n18834 & ~n18836;
  assign n18954 = ~n18837 & ~n18953;
  assign n18955 = n8250 & n12410;
  assign n18956 = n8251 & n13093;
  assign n18957 = n9016 & n12407;
  assign n18958 = n9040 & n12404;
  assign n18959 = ~n18955 & ~n18957;
  assign n18960 = ~n18958 & n18959;
  assign n18961 = ~n18956 & n18960;
  assign n18962 = pi8  & n18961;
  assign n18963 = ~pi8  & ~n18961;
  assign n18964 = ~n18962 & ~n18963;
  assign n18965 = n18954 & ~n18964;
  assign n18966 = n18830 & ~n18832;
  assign n18967 = ~n18833 & ~n18966;
  assign n18968 = n8250 & n12413;
  assign n18969 = n8251 & n12891;
  assign n18970 = n9016 & n12410;
  assign n18971 = n9040 & n12407;
  assign n18972 = ~n18968 & ~n18970;
  assign n18973 = ~n18971 & n18972;
  assign n18974 = ~n18969 & n18973;
  assign n18975 = pi8  & n18974;
  assign n18976 = ~pi8  & ~n18974;
  assign n18977 = ~n18975 & ~n18976;
  assign n18978 = n18967 & ~n18977;
  assign n18979 = n18826 & ~n18828;
  assign n18980 = ~n18829 & ~n18979;
  assign n18981 = n8250 & n12416;
  assign n18982 = n8251 & n12843;
  assign n18983 = n9016 & n12413;
  assign n18984 = n9040 & n12410;
  assign n18985 = ~n18981 & ~n18983;
  assign n18986 = ~n18984 & n18985;
  assign n18987 = ~n18982 & n18986;
  assign n18988 = pi8  & n18987;
  assign n18989 = ~pi8  & ~n18987;
  assign n18990 = ~n18988 & ~n18989;
  assign n18991 = n18980 & ~n18990;
  assign n18992 = n18451 & n18824;
  assign n18993 = ~n18825 & ~n18992;
  assign n18994 = n8250 & n12419;
  assign n18995 = n8251 & n12908;
  assign n18996 = n9016 & n12416;
  assign n18997 = n9040 & n12413;
  assign n18998 = ~n18994 & ~n18996;
  assign n18999 = ~n18997 & n18998;
  assign n19000 = ~n18995 & n18999;
  assign n19001 = pi8  & n19000;
  assign n19002 = ~pi8  & ~n19000;
  assign n19003 = ~n19001 & ~n19002;
  assign n19004 = n18993 & ~n19003;
  assign n19005 = n18467 & n18822;
  assign n19006 = ~n18823 & ~n19005;
  assign n19007 = n8250 & n12422;
  assign n19008 = n8251 & n13201;
  assign n19009 = n9016 & n12419;
  assign n19010 = n9040 & n12416;
  assign n19011 = ~n19007 & ~n19009;
  assign n19012 = ~n19010 & n19011;
  assign n19013 = ~n19008 & n19012;
  assign n19014 = pi8  & n19013;
  assign n19015 = ~pi8  & ~n19013;
  assign n19016 = ~n19014 & ~n19015;
  assign n19017 = n19006 & ~n19016;
  assign n19018 = n8250 & n12425;
  assign n19019 = n8251 & n13010;
  assign n19020 = n9016 & n12422;
  assign n19021 = n9040 & n12419;
  assign n19022 = ~n19018 & ~n19020;
  assign n19023 = ~n19021 & n19022;
  assign n19024 = ~n19019 & n19023;
  assign n19025 = ~pi8  & ~n19024;
  assign n19026 = pi8  & n19024;
  assign n19027 = ~n19025 & ~n19026;
  assign n19028 = n18818 & ~n18820;
  assign n19029 = ~n18821 & ~n19028;
  assign n19030 = ~n19027 & n19029;
  assign n19031 = ~n19027 & ~n19029;
  assign n19032 = n19027 & n19029;
  assign n19033 = ~n19031 & ~n19032;
  assign n19034 = n8250 & n12428;
  assign n19035 = n8251 & n13371;
  assign n19036 = n9016 & n12425;
  assign n19037 = n9040 & n12422;
  assign n19038 = ~n19034 & ~n19036;
  assign n19039 = ~n19037 & n19038;
  assign n19040 = ~n19035 & n19039;
  assign n19041 = ~pi8  & ~n19040;
  assign n19042 = pi8  & n19040;
  assign n19043 = ~n19041 & ~n19042;
  assign n19044 = ~n18813 & n18816;
  assign n19045 = n18813 & ~n18816;
  assign n19046 = ~n19044 & ~n19045;
  assign n19047 = ~n19043 & ~n19046;
  assign n19048 = n18509 & n18811;
  assign n19049 = ~n18812 & ~n19048;
  assign n19050 = n8250 & n12431;
  assign n19051 = n8251 & n13356;
  assign n19052 = n9016 & n12428;
  assign n19053 = n9040 & n12425;
  assign n19054 = ~n19050 & ~n19052;
  assign n19055 = ~n19053 & n19054;
  assign n19056 = ~n19051 & n19055;
  assign n19057 = pi8  & n19056;
  assign n19058 = ~pi8  & ~n19056;
  assign n19059 = ~n19057 & ~n19058;
  assign n19060 = n19049 & ~n19059;
  assign n19061 = n18807 & ~n18809;
  assign n19062 = ~n18810 & ~n19061;
  assign n19063 = n8250 & n12434;
  assign n19064 = n8251 & n13546;
  assign n19065 = n9016 & n12431;
  assign n19066 = n9040 & n12428;
  assign n19067 = ~n19063 & ~n19065;
  assign n19068 = ~n19066 & n19067;
  assign n19069 = ~n19064 & n19068;
  assign n19070 = pi8  & n19069;
  assign n19071 = ~pi8  & ~n19069;
  assign n19072 = ~n19070 & ~n19071;
  assign n19073 = n19062 & ~n19072;
  assign n19074 = n18539 & n18805;
  assign n19075 = ~n18806 & ~n19074;
  assign n19076 = n8250 & n12437;
  assign n19077 = n8251 & n13564;
  assign n19078 = n9016 & n12434;
  assign n19079 = n9040 & n12431;
  assign n19080 = ~n19076 & ~n19078;
  assign n19081 = ~n19079 & n19080;
  assign n19082 = ~n19077 & n19081;
  assign n19083 = pi8  & n19082;
  assign n19084 = ~pi8  & ~n19082;
  assign n19085 = ~n19083 & ~n19084;
  assign n19086 = n19075 & ~n19085;
  assign n19087 = n8250 & n12440;
  assign n19088 = n8251 & n13939;
  assign n19089 = n9016 & n12437;
  assign n19090 = n9040 & n12434;
  assign n19091 = ~n19087 & ~n19089;
  assign n19092 = ~n19090 & n19091;
  assign n19093 = ~n19088 & n19092;
  assign n19094 = ~pi8  & ~n19093;
  assign n19095 = pi8  & n19093;
  assign n19096 = ~n19094 & ~n19095;
  assign n19097 = n18801 & ~n18803;
  assign n19098 = ~n18804 & ~n19097;
  assign n19099 = ~n19096 & n19098;
  assign n19100 = ~n19096 & ~n19098;
  assign n19101 = n19096 & n19098;
  assign n19102 = ~n19100 & ~n19101;
  assign n19103 = n8250 & n12443;
  assign n19104 = n8251 & n13702;
  assign n19105 = n9016 & n12440;
  assign n19106 = n9040 & n12437;
  assign n19107 = ~n19103 & ~n19105;
  assign n19108 = ~n19106 & n19107;
  assign n19109 = ~n19104 & n19108;
  assign n19110 = ~pi8  & ~n19109;
  assign n19111 = pi8  & n19109;
  assign n19112 = ~n19110 & ~n19111;
  assign n19113 = ~n18796 & n18799;
  assign n19114 = n18796 & ~n18799;
  assign n19115 = ~n19113 & ~n19114;
  assign n19116 = ~n19112 & ~n19115;
  assign n19117 = n8250 & n12446;
  assign n19118 = n8251 & n14175;
  assign n19119 = n9016 & n12443;
  assign n19120 = n9040 & n12440;
  assign n19121 = ~n19117 & ~n19119;
  assign n19122 = ~n19120 & n19121;
  assign n19123 = ~n19118 & n19122;
  assign n19124 = ~pi8  & ~n19123;
  assign n19125 = pi8  & n19123;
  assign n19126 = ~n19124 & ~n19125;
  assign n19127 = n18791 & n18794;
  assign n19128 = ~n18795 & ~n19127;
  assign n19129 = ~n19126 & n19128;
  assign n19130 = ~n19126 & ~n19128;
  assign n19131 = n19126 & n19128;
  assign n19132 = ~n19130 & ~n19131;
  assign n19133 = n18594 & n18789;
  assign n19134 = ~n18790 & ~n19133;
  assign n19135 = n8250 & n12449;
  assign n19136 = n8251 & n14325;
  assign n19137 = n9016 & n12446;
  assign n19138 = n9040 & n12443;
  assign n19139 = ~n19135 & ~n19137;
  assign n19140 = ~n19138 & n19139;
  assign n19141 = ~n19136 & n19140;
  assign n19142 = pi8  & n19141;
  assign n19143 = ~pi8  & ~n19141;
  assign n19144 = ~n19142 & ~n19143;
  assign n19145 = n19134 & ~n19144;
  assign n19146 = n18610 & n18787;
  assign n19147 = ~n18788 & ~n19146;
  assign n19148 = n8250 & n12452;
  assign n19149 = n8251 & n14156;
  assign n19150 = n9016 & n12449;
  assign n19151 = n9040 & n12446;
  assign n19152 = ~n19148 & ~n19150;
  assign n19153 = ~n19151 & n19152;
  assign n19154 = ~n19149 & n19153;
  assign n19155 = pi8  & n19154;
  assign n19156 = ~pi8  & ~n19154;
  assign n19157 = ~n19155 & ~n19156;
  assign n19158 = n19147 & ~n19157;
  assign n19159 = n18783 & ~n18785;
  assign n19160 = ~n18786 & ~n19159;
  assign n19161 = n8250 & n12455;
  assign n19162 = n8251 & n14442;
  assign n19163 = n9016 & n12452;
  assign n19164 = n9040 & n12449;
  assign n19165 = ~n19161 & ~n19163;
  assign n19166 = ~n19164 & n19165;
  assign n19167 = ~n19162 & n19166;
  assign n19168 = pi8  & n19167;
  assign n19169 = ~pi8  & ~n19167;
  assign n19170 = ~n19168 & ~n19169;
  assign n19171 = n19160 & ~n19170;
  assign n19172 = n8250 & n12458;
  assign n19173 = n8251 & n14741;
  assign n19174 = n9016 & n12455;
  assign n19175 = n9040 & n12452;
  assign n19176 = ~n19172 & ~n19174;
  assign n19177 = ~n19175 & n19176;
  assign n19178 = ~n19173 & n19177;
  assign n19179 = ~pi8  & ~n19178;
  assign n19180 = pi8  & n19178;
  assign n19181 = ~n19179 & ~n19180;
  assign n19182 = n18779 & ~n18781;
  assign n19183 = ~n18782 & ~n19182;
  assign n19184 = ~n19181 & n19183;
  assign n19185 = ~n19181 & ~n19183;
  assign n19186 = n19181 & n19183;
  assign n19187 = ~n19185 & ~n19186;
  assign n19188 = n8250 & n12461;
  assign n19189 = n8251 & n14756;
  assign n19190 = n9016 & n12458;
  assign n19191 = n9040 & n12455;
  assign n19192 = ~n19188 & ~n19190;
  assign n19193 = ~n19191 & n19192;
  assign n19194 = ~n19189 & n19193;
  assign n19195 = ~pi8  & ~n19194;
  assign n19196 = pi8  & n19194;
  assign n19197 = ~n19195 & ~n19196;
  assign n19198 = n18774 & n18777;
  assign n19199 = ~n18778 & ~n19198;
  assign n19200 = ~n19197 & n19199;
  assign n19201 = ~n19197 & ~n19199;
  assign n19202 = n19197 & n19199;
  assign n19203 = ~n19201 & ~n19202;
  assign n19204 = n8250 & n12464;
  assign n19205 = n8251 & n14420;
  assign n19206 = n9016 & n12461;
  assign n19207 = n9040 & n12458;
  assign n19208 = ~n19204 & ~n19206;
  assign n19209 = ~n19207 & n19208;
  assign n19210 = ~n19205 & n19209;
  assign n19211 = ~pi8  & ~n19210;
  assign n19212 = pi8  & n19210;
  assign n19213 = ~n19211 & ~n19212;
  assign n19214 = ~n18769 & n18772;
  assign n19215 = n18769 & ~n18772;
  assign n19216 = ~n19214 & ~n19215;
  assign n19217 = ~n19213 & ~n19216;
  assign n19218 = n18679 & n18767;
  assign n19219 = ~n18768 & ~n19218;
  assign n19220 = n8250 & n12467;
  assign n19221 = n8251 & n14789;
  assign n19222 = n9016 & n12464;
  assign n19223 = n9040 & n12461;
  assign n19224 = ~n19220 & ~n19222;
  assign n19225 = ~n19223 & n19224;
  assign n19226 = ~n19221 & n19225;
  assign n19227 = pi8  & n19226;
  assign n19228 = ~pi8  & ~n19226;
  assign n19229 = ~n19227 & ~n19228;
  assign n19230 = n19219 & ~n19229;
  assign n19231 = n18763 & ~n18765;
  assign n19232 = ~n18766 & ~n19231;
  assign n19233 = n8250 & n12470;
  assign n19234 = n8251 & n14815;
  assign n19235 = n9016 & n12467;
  assign n19236 = n9040 & n12464;
  assign n19237 = ~n19233 & ~n19235;
  assign n19238 = ~n19236 & n19237;
  assign n19239 = ~n19234 & n19238;
  assign n19240 = pi8  & n19239;
  assign n19241 = ~pi8  & ~n19239;
  assign n19242 = ~n19240 & ~n19241;
  assign n19243 = n19232 & ~n19242;
  assign n19244 = n18710 & n18761;
  assign n19245 = ~n18762 & ~n19244;
  assign n19246 = n8250 & n12473;
  assign n19247 = n8251 & n14839;
  assign n19248 = n9016 & n12470;
  assign n19249 = n9040 & n12467;
  assign n19250 = ~n19246 & ~n19248;
  assign n19251 = ~n19249 & n19250;
  assign n19252 = ~n19247 & n19251;
  assign n19253 = pi8  & n19252;
  assign n19254 = ~pi8  & ~n19252;
  assign n19255 = ~n19253 & ~n19254;
  assign n19256 = n19245 & ~n19255;
  assign n19257 = n8250 & n12476;
  assign n19258 = n8251 & n14849;
  assign n19259 = n9016 & n12473;
  assign n19260 = n9040 & n12470;
  assign n19261 = ~n19257 & ~n19259;
  assign n19262 = ~n19260 & n19261;
  assign n19263 = ~n19258 & n19262;
  assign n19264 = ~pi8  & ~n19263;
  assign n19265 = pi8  & n19263;
  assign n19266 = ~n19264 & ~n19265;
  assign n19267 = n18757 & ~n18759;
  assign n19268 = ~n18760 & ~n19267;
  assign n19269 = ~n19266 & n19268;
  assign n19270 = ~n19266 & ~n19268;
  assign n19271 = n19266 & n19268;
  assign n19272 = ~n19270 & ~n19271;
  assign n19273 = n8250 & n12479;
  assign n19274 = n8251 & n14922;
  assign n19275 = n9016 & n12476;
  assign n19276 = n9040 & n12473;
  assign n19277 = ~n19273 & ~n19275;
  assign n19278 = ~n19276 & n19277;
  assign n19279 = ~n19274 & n19278;
  assign n19280 = pi8  & n19279;
  assign n19281 = ~pi8  & ~n19279;
  assign n19282 = ~n19280 & ~n19281;
  assign n19283 = n18745 & n18755;
  assign n19284 = ~n18756 & ~n19283;
  assign n19285 = ~n19282 & n19284;
  assign n19286 = n8250 & n12482;
  assign n19287 = n8251 & n14958;
  assign n19288 = n9016 & n12479;
  assign n19289 = n9040 & n12476;
  assign n19290 = ~n19286 & ~n19288;
  assign n19291 = ~n19289 & n19290;
  assign n19292 = ~n19287 & n19291;
  assign n19293 = ~pi8  & ~n19292;
  assign n19294 = pi8  & n19292;
  assign n19295 = ~n19293 & ~n19294;
  assign n19296 = pi11  & ~n18733;
  assign n19297 = n18740 & ~n19296;
  assign n19298 = ~n18740 & n19296;
  assign n19299 = ~n19297 & ~n19298;
  assign n19300 = ~n19295 & n19299;
  assign n19301 = ~n19295 & ~n19299;
  assign n19302 = n19295 & n19299;
  assign n19303 = ~n19301 & ~n19302;
  assign n19304 = n8250 & n12485;
  assign n19305 = n8251 & n15001;
  assign n19306 = n9016 & n12482;
  assign n19307 = n9040 & n12479;
  assign n19308 = ~n19304 & ~n19306;
  assign n19309 = ~n19307 & n19308;
  assign n19310 = ~n19305 & n19309;
  assign n19311 = pi8  & n19310;
  assign n19312 = ~pi8  & ~n19310;
  assign n19313 = ~n19311 & ~n19312;
  assign n19314 = pi11  & n18726;
  assign n19315 = ~n18731 & n19314;
  assign n19316 = n18731 & ~n19314;
  assign n19317 = ~n19315 & ~n19316;
  assign n19318 = ~n19313 & n19317;
  assign n19319 = ~n8245 & n12492;
  assign n19320 = n9016 & n12492;
  assign n19321 = n9040 & n12490;
  assign n19322 = n8251 & ~n15072;
  assign n19323 = ~n19320 & ~n19321;
  assign n19324 = ~n19322 & n19323;
  assign n19325 = pi8  & ~n19319;
  assign n19326 = n19324 & n19325;
  assign n19327 = n8250 & n12492;
  assign n19328 = n8251 & ~n15113;
  assign n19329 = n9016 & n12490;
  assign n19330 = n9040 & n12485;
  assign n19331 = ~n19327 & ~n19329;
  assign n19332 = ~n19330 & n19331;
  assign n19333 = ~n19328 & n19332;
  assign n19334 = n19326 & n19333;
  assign n19335 = n18726 & n19334;
  assign n19336 = ~n18726 & n19334;
  assign n19337 = n18726 & ~n19334;
  assign n19338 = ~n19336 & ~n19337;
  assign n19339 = n8250 & n12490;
  assign n19340 = n8251 & n15026;
  assign n19341 = n9016 & n12485;
  assign n19342 = n9040 & n12482;
  assign n19343 = ~n19339 & ~n19341;
  assign n19344 = ~n19342 & n19343;
  assign n19345 = ~n19340 & n19344;
  assign n19346 = pi8  & n19345;
  assign n19347 = ~pi8  & ~n19345;
  assign n19348 = ~n19346 & ~n19347;
  assign n19349 = ~n19338 & ~n19348;
  assign n19350 = ~n19335 & ~n19349;
  assign n19351 = n19313 & ~n19317;
  assign n19352 = ~n19318 & ~n19351;
  assign n19353 = ~n19350 & n19352;
  assign n19354 = ~n19318 & ~n19353;
  assign n19355 = ~n19303 & ~n19354;
  assign n19356 = ~n19300 & ~n19355;
  assign n19357 = n19282 & ~n19284;
  assign n19358 = ~n19285 & ~n19357;
  assign n19359 = ~n19356 & n19358;
  assign n19360 = ~n19285 & ~n19359;
  assign n19361 = ~n19272 & ~n19360;
  assign n19362 = ~n19269 & ~n19361;
  assign n19363 = n19245 & n19255;
  assign n19364 = ~n19245 & ~n19255;
  assign n19365 = ~n19363 & ~n19364;
  assign n19366 = ~n19362 & ~n19365;
  assign n19367 = ~n19256 & ~n19366;
  assign n19368 = n19232 & n19242;
  assign n19369 = ~n19232 & ~n19242;
  assign n19370 = ~n19368 & ~n19369;
  assign n19371 = ~n19367 & ~n19370;
  assign n19372 = ~n19243 & ~n19371;
  assign n19373 = ~n19219 & n19229;
  assign n19374 = ~n19230 & ~n19373;
  assign n19375 = ~n19372 & n19374;
  assign n19376 = ~n19230 & ~n19375;
  assign n19377 = n19213 & n19216;
  assign n19378 = ~n19217 & ~n19377;
  assign n19379 = ~n19376 & n19378;
  assign n19380 = ~n19217 & ~n19379;
  assign n19381 = ~n19203 & ~n19380;
  assign n19382 = ~n19200 & ~n19381;
  assign n19383 = ~n19187 & ~n19382;
  assign n19384 = ~n19184 & ~n19383;
  assign n19385 = n19160 & n19170;
  assign n19386 = ~n19160 & ~n19170;
  assign n19387 = ~n19385 & ~n19386;
  assign n19388 = ~n19384 & ~n19387;
  assign n19389 = ~n19171 & ~n19388;
  assign n19390 = n19147 & n19157;
  assign n19391 = ~n19147 & ~n19157;
  assign n19392 = ~n19390 & ~n19391;
  assign n19393 = ~n19389 & ~n19392;
  assign n19394 = ~n19158 & ~n19393;
  assign n19395 = ~n19134 & n19144;
  assign n19396 = ~n19145 & ~n19395;
  assign n19397 = ~n19394 & n19396;
  assign n19398 = ~n19145 & ~n19397;
  assign n19399 = ~n19132 & ~n19398;
  assign n19400 = ~n19129 & ~n19399;
  assign n19401 = n19112 & n19115;
  assign n19402 = ~n19116 & ~n19401;
  assign n19403 = ~n19400 & n19402;
  assign n19404 = ~n19116 & ~n19403;
  assign n19405 = ~n19102 & ~n19404;
  assign n19406 = ~n19099 & ~n19405;
  assign n19407 = n19075 & n19085;
  assign n19408 = ~n19075 & ~n19085;
  assign n19409 = ~n19407 & ~n19408;
  assign n19410 = ~n19406 & ~n19409;
  assign n19411 = ~n19086 & ~n19410;
  assign n19412 = n19062 & n19072;
  assign n19413 = ~n19062 & ~n19072;
  assign n19414 = ~n19412 & ~n19413;
  assign n19415 = ~n19411 & ~n19414;
  assign n19416 = ~n19073 & ~n19415;
  assign n19417 = ~n19049 & n19059;
  assign n19418 = ~n19060 & ~n19417;
  assign n19419 = ~n19416 & n19418;
  assign n19420 = ~n19060 & ~n19419;
  assign n19421 = n19043 & n19046;
  assign n19422 = ~n19047 & ~n19421;
  assign n19423 = ~n19420 & n19422;
  assign n19424 = ~n19047 & ~n19423;
  assign n19425 = ~n19033 & ~n19424;
  assign n19426 = ~n19030 & ~n19425;
  assign n19427 = n19006 & n19016;
  assign n19428 = ~n19006 & ~n19016;
  assign n19429 = ~n19427 & ~n19428;
  assign n19430 = ~n19426 & ~n19429;
  assign n19431 = ~n19017 & ~n19430;
  assign n19432 = n18993 & n19003;
  assign n19433 = ~n18993 & ~n19003;
  assign n19434 = ~n19432 & ~n19433;
  assign n19435 = ~n19431 & ~n19434;
  assign n19436 = ~n19004 & ~n19435;
  assign n19437 = n18980 & n18990;
  assign n19438 = ~n18980 & ~n18990;
  assign n19439 = ~n19437 & ~n19438;
  assign n19440 = ~n19436 & ~n19439;
  assign n19441 = ~n18991 & ~n19440;
  assign n19442 = n18967 & n18977;
  assign n19443 = ~n18967 & ~n18977;
  assign n19444 = ~n19442 & ~n19443;
  assign n19445 = ~n19441 & ~n19444;
  assign n19446 = ~n18978 & ~n19445;
  assign n19447 = n18954 & n18964;
  assign n19448 = ~n18954 & ~n18964;
  assign n19449 = ~n19447 & ~n19448;
  assign n19450 = ~n19446 & ~n19449;
  assign n19451 = ~n18965 & ~n19450;
  assign n19452 = n18941 & n18951;
  assign n19453 = ~n18941 & ~n18951;
  assign n19454 = ~n19452 & ~n19453;
  assign n19455 = ~n19451 & ~n19454;
  assign n19456 = ~n18952 & ~n19455;
  assign n19457 = n18928 & n18938;
  assign n19458 = ~n18928 & ~n18938;
  assign n19459 = ~n19457 & ~n19458;
  assign n19460 = ~n19456 & ~n19459;
  assign n19461 = ~n18939 & ~n19460;
  assign n19462 = n18915 & n18925;
  assign n19463 = ~n18915 & ~n18925;
  assign n19464 = ~n19462 & ~n19463;
  assign n19465 = ~n19461 & ~n19464;
  assign n19466 = ~n18926 & ~n19465;
  assign n19467 = n18902 & n18912;
  assign n19468 = ~n18902 & ~n18912;
  assign n19469 = ~n19467 & ~n19468;
  assign n19470 = ~n19466 & ~n19469;
  assign n19471 = ~n18913 & ~n19470;
  assign n19472 = ~n18889 & n18899;
  assign n19473 = ~n18900 & ~n19472;
  assign n19474 = ~n19471 & n19473;
  assign n19475 = ~n18900 & ~n19474;
  assign n19476 = ~n18853 & ~n18854;
  assign n19477 = ~n18864 & n19476;
  assign n19478 = n18864 & ~n19476;
  assign n19479 = ~n19477 & ~n19478;
  assign n19480 = ~n19475 & n19479;
  assign n19481 = n19475 & ~n19479;
  assign n19482 = n11031 & n13161;
  assign n19483 = n9491 & n13183;
  assign n19484 = n10469 & n13166;
  assign n19485 = n75 & n13164;
  assign n19486 = ~n19484 & ~n19485;
  assign n19487 = ~n19482 & n19486;
  assign n19488 = ~n19483 & n19487;
  assign n19489 = pi5  & n19488;
  assign n19490 = ~pi5  & ~n19488;
  assign n19491 = ~n19489 & ~n19490;
  assign n19492 = ~n19481 & ~n19491;
  assign n19493 = ~n19480 & ~n19492;
  assign n19494 = n18887 & ~n19493;
  assign n19495 = ~n18887 & n19493;
  assign n19496 = ~n19494 & ~n19495;
  assign n19497 = n75 & n12646;
  assign n19498 = n9491 & n13261;
  assign n19499 = n10469 & n13164;
  assign n19500 = n11031 & n13166;
  assign n19501 = ~n19497 & ~n19499;
  assign n19502 = ~n19500 & n19501;
  assign n19503 = ~n19498 & n19502;
  assign n19504 = ~pi5  & ~n19503;
  assign n19505 = pi5  & n19503;
  assign n19506 = ~n19504 & ~n19505;
  assign n19507 = n19471 & ~n19473;
  assign n19508 = ~n19474 & ~n19507;
  assign n19509 = ~n19506 & n19508;
  assign n19510 = ~n19506 & ~n19508;
  assign n19511 = n19506 & n19508;
  assign n19512 = ~n19510 & ~n19511;
  assign n19513 = n11056 & ~n13280;
  assign n19514 = ~n11054 & ~n11056;
  assign n19515 = n11055 & ~n13160;
  assign n19516 = ~n19514 & ~n19515;
  assign n19517 = ~n12786 & ~n19516;
  assign n19518 = ~n19513 & ~n19517;
  assign n19519 = pi2  & n19518;
  assign n19520 = ~pi2  & ~n19518;
  assign n19521 = ~n19519 & ~n19520;
  assign n19522 = ~n19512 & ~n19521;
  assign n19523 = ~n19509 & ~n19522;
  assign n19524 = ~n19480 & ~n19481;
  assign n19525 = ~n19491 & n19524;
  assign n19526 = n19491 & ~n19524;
  assign n19527 = ~n19525 & ~n19526;
  assign n19528 = ~n19523 & n19527;
  assign n19529 = n19523 & ~n19527;
  assign n19530 = ~n19528 & ~n19529;
  assign n19531 = n75 & n12392;
  assign n19532 = n9491 & n13421;
  assign n19533 = n10469 & n12646;
  assign n19534 = n11031 & n13164;
  assign n19535 = ~n19531 & ~n19533;
  assign n19536 = ~n19534 & n19535;
  assign n19537 = ~n19532 & n19536;
  assign n19538 = ~pi5  & ~n19537;
  assign n19539 = pi5  & n19537;
  assign n19540 = ~n19538 & ~n19539;
  assign n19541 = ~n19466 & n19469;
  assign n19542 = n19466 & ~n19469;
  assign n19543 = ~n19541 & ~n19542;
  assign n19544 = ~n19540 & ~n19543;
  assign n19545 = n75 & n12362;
  assign n19546 = n9491 & n12652;
  assign n19547 = n10469 & n12392;
  assign n19548 = n11031 & n12646;
  assign n19549 = ~n19545 & ~n19547;
  assign n19550 = ~n19548 & n19549;
  assign n19551 = ~n19546 & n19550;
  assign n19552 = ~pi5  & ~n19551;
  assign n19553 = pi5  & n19551;
  assign n19554 = ~n19552 & ~n19553;
  assign n19555 = ~n19461 & n19464;
  assign n19556 = n19461 & ~n19464;
  assign n19557 = ~n19555 & ~n19556;
  assign n19558 = ~n19554 & ~n19557;
  assign n19559 = n75 & n12395;
  assign n19560 = n9491 & n13144;
  assign n19561 = n10469 & n12362;
  assign n19562 = n11031 & n12392;
  assign n19563 = ~n19559 & ~n19561;
  assign n19564 = ~n19562 & n19563;
  assign n19565 = ~n19560 & n19564;
  assign n19566 = ~pi5  & ~n19565;
  assign n19567 = pi5  & n19565;
  assign n19568 = ~n19566 & ~n19567;
  assign n19569 = ~n19456 & n19459;
  assign n19570 = n19456 & ~n19459;
  assign n19571 = ~n19569 & ~n19570;
  assign n19572 = ~n19568 & ~n19571;
  assign n19573 = n75 & n12398;
  assign n19574 = n9491 & n13245;
  assign n19575 = n10469 & n12395;
  assign n19576 = n11031 & n12362;
  assign n19577 = ~n19573 & ~n19575;
  assign n19578 = ~n19576 & n19577;
  assign n19579 = ~n19574 & n19578;
  assign n19580 = ~pi5  & ~n19579;
  assign n19581 = pi5  & n19579;
  assign n19582 = ~n19580 & ~n19581;
  assign n19583 = ~n19451 & n19454;
  assign n19584 = n19451 & ~n19454;
  assign n19585 = ~n19583 & ~n19584;
  assign n19586 = ~n19582 & ~n19585;
  assign n19587 = n75 & n12401;
  assign n19588 = n9491 & n13108;
  assign n19589 = n10469 & n12398;
  assign n19590 = n11031 & n12395;
  assign n19591 = ~n19587 & ~n19589;
  assign n19592 = ~n19590 & n19591;
  assign n19593 = ~n19588 & n19592;
  assign n19594 = ~pi5  & ~n19593;
  assign n19595 = pi5  & n19593;
  assign n19596 = ~n19594 & ~n19595;
  assign n19597 = n19446 & n19449;
  assign n19598 = ~n19450 & ~n19597;
  assign n19599 = ~n19596 & n19598;
  assign n19600 = ~n19596 & ~n19598;
  assign n19601 = n19596 & n19598;
  assign n19602 = ~n19600 & ~n19601;
  assign n19603 = n75 & n12404;
  assign n19604 = n9491 & n13128;
  assign n19605 = n10469 & n12401;
  assign n19606 = n11031 & n12398;
  assign n19607 = ~n19603 & ~n19605;
  assign n19608 = ~n19606 & n19607;
  assign n19609 = ~n19604 & n19608;
  assign n19610 = ~pi5  & ~n19609;
  assign n19611 = pi5  & n19609;
  assign n19612 = ~n19610 & ~n19611;
  assign n19613 = n19441 & n19444;
  assign n19614 = ~n19445 & ~n19613;
  assign n19615 = ~n19612 & n19614;
  assign n19616 = ~n19612 & ~n19614;
  assign n19617 = n19612 & n19614;
  assign n19618 = ~n19616 & ~n19617;
  assign n19619 = n75 & n12407;
  assign n19620 = n9491 & n13035;
  assign n19621 = n10469 & n12404;
  assign n19622 = n11031 & n12401;
  assign n19623 = ~n19619 & ~n19621;
  assign n19624 = ~n19622 & n19623;
  assign n19625 = ~n19620 & n19624;
  assign n19626 = ~pi5  & ~n19625;
  assign n19627 = pi5  & n19625;
  assign n19628 = ~n19626 & ~n19627;
  assign n19629 = n19436 & n19439;
  assign n19630 = ~n19440 & ~n19629;
  assign n19631 = ~n19628 & n19630;
  assign n19632 = ~n19628 & ~n19630;
  assign n19633 = n19628 & n19630;
  assign n19634 = ~n19632 & ~n19633;
  assign n19635 = n75 & n12410;
  assign n19636 = n9491 & n13093;
  assign n19637 = n10469 & n12407;
  assign n19638 = n11031 & n12404;
  assign n19639 = ~n19635 & ~n19637;
  assign n19640 = ~n19638 & n19639;
  assign n19641 = ~n19636 & n19640;
  assign n19642 = ~pi5  & ~n19641;
  assign n19643 = pi5  & n19641;
  assign n19644 = ~n19642 & ~n19643;
  assign n19645 = ~n19431 & n19434;
  assign n19646 = n19431 & ~n19434;
  assign n19647 = ~n19645 & ~n19646;
  assign n19648 = ~n19644 & ~n19647;
  assign n19649 = n75 & n12413;
  assign n19650 = n9491 & n12891;
  assign n19651 = n10469 & n12410;
  assign n19652 = n11031 & n12407;
  assign n19653 = ~n19649 & ~n19651;
  assign n19654 = ~n19652 & n19653;
  assign n19655 = ~n19650 & n19654;
  assign n19656 = ~pi5  & ~n19655;
  assign n19657 = pi5  & n19655;
  assign n19658 = ~n19656 & ~n19657;
  assign n19659 = ~n19426 & n19429;
  assign n19660 = n19426 & ~n19429;
  assign n19661 = ~n19659 & ~n19660;
  assign n19662 = ~n19658 & ~n19661;
  assign n19663 = n19033 & n19424;
  assign n19664 = ~n19425 & ~n19663;
  assign n19665 = n75 & n12416;
  assign n19666 = n9491 & n12843;
  assign n19667 = n10469 & n12413;
  assign n19668 = n11031 & n12410;
  assign n19669 = ~n19665 & ~n19667;
  assign n19670 = ~n19668 & n19669;
  assign n19671 = ~n19666 & n19670;
  assign n19672 = pi5  & n19671;
  assign n19673 = ~pi5  & ~n19671;
  assign n19674 = ~n19672 & ~n19673;
  assign n19675 = n19664 & ~n19674;
  assign n19676 = n19420 & ~n19422;
  assign n19677 = ~n19423 & ~n19676;
  assign n19678 = n75 & n12419;
  assign n19679 = n9491 & n12908;
  assign n19680 = n10469 & n12416;
  assign n19681 = n11031 & n12413;
  assign n19682 = ~n19678 & ~n19680;
  assign n19683 = ~n19681 & n19682;
  assign n19684 = ~n19679 & n19683;
  assign n19685 = pi5  & n19684;
  assign n19686 = ~pi5  & ~n19684;
  assign n19687 = ~n19685 & ~n19686;
  assign n19688 = n19677 & ~n19687;
  assign n19689 = n75 & n12422;
  assign n19690 = n9491 & n13201;
  assign n19691 = n10469 & n12419;
  assign n19692 = n11031 & n12416;
  assign n19693 = ~n19689 & ~n19691;
  assign n19694 = ~n19692 & n19693;
  assign n19695 = ~n19690 & n19694;
  assign n19696 = ~pi5  & ~n19695;
  assign n19697 = pi5  & n19695;
  assign n19698 = ~n19696 & ~n19697;
  assign n19699 = n19416 & ~n19418;
  assign n19700 = ~n19419 & ~n19699;
  assign n19701 = ~n19698 & n19700;
  assign n19702 = ~n19698 & ~n19700;
  assign n19703 = n19698 & n19700;
  assign n19704 = ~n19702 & ~n19703;
  assign n19705 = n75 & n12425;
  assign n19706 = n9491 & n13010;
  assign n19707 = n10469 & n12422;
  assign n19708 = n11031 & n12419;
  assign n19709 = ~n19705 & ~n19707;
  assign n19710 = ~n19708 & n19709;
  assign n19711 = ~n19706 & n19710;
  assign n19712 = ~pi5  & ~n19711;
  assign n19713 = pi5  & n19711;
  assign n19714 = ~n19712 & ~n19713;
  assign n19715 = n19411 & n19414;
  assign n19716 = ~n19415 & ~n19715;
  assign n19717 = ~n19714 & n19716;
  assign n19718 = ~n19714 & ~n19716;
  assign n19719 = n19714 & n19716;
  assign n19720 = ~n19718 & ~n19719;
  assign n19721 = n75 & n12428;
  assign n19722 = n9491 & n13371;
  assign n19723 = n10469 & n12425;
  assign n19724 = n11031 & n12422;
  assign n19725 = ~n19721 & ~n19723;
  assign n19726 = ~n19724 & n19725;
  assign n19727 = ~n19722 & n19726;
  assign n19728 = ~pi5  & ~n19727;
  assign n19729 = pi5  & n19727;
  assign n19730 = ~n19728 & ~n19729;
  assign n19731 = ~n19406 & n19409;
  assign n19732 = n19406 & ~n19409;
  assign n19733 = ~n19731 & ~n19732;
  assign n19734 = ~n19730 & ~n19733;
  assign n19735 = n19102 & n19404;
  assign n19736 = ~n19405 & ~n19735;
  assign n19737 = n75 & n12431;
  assign n19738 = n9491 & n13356;
  assign n19739 = n10469 & n12428;
  assign n19740 = n11031 & n12425;
  assign n19741 = ~n19737 & ~n19739;
  assign n19742 = ~n19740 & n19741;
  assign n19743 = ~n19738 & n19742;
  assign n19744 = pi5  & n19743;
  assign n19745 = ~pi5  & ~n19743;
  assign n19746 = ~n19744 & ~n19745;
  assign n19747 = n19736 & ~n19746;
  assign n19748 = n19400 & ~n19402;
  assign n19749 = ~n19403 & ~n19748;
  assign n19750 = n75 & n12434;
  assign n19751 = n9491 & n13546;
  assign n19752 = n10469 & n12431;
  assign n19753 = n11031 & n12428;
  assign n19754 = ~n19750 & ~n19752;
  assign n19755 = ~n19753 & n19754;
  assign n19756 = ~n19751 & n19755;
  assign n19757 = pi5  & n19756;
  assign n19758 = ~pi5  & ~n19756;
  assign n19759 = ~n19757 & ~n19758;
  assign n19760 = n19749 & ~n19759;
  assign n19761 = n19132 & n19398;
  assign n19762 = ~n19399 & ~n19761;
  assign n19763 = n75 & n12437;
  assign n19764 = n9491 & n13564;
  assign n19765 = n10469 & n12434;
  assign n19766 = n11031 & n12431;
  assign n19767 = ~n19763 & ~n19765;
  assign n19768 = ~n19766 & n19767;
  assign n19769 = ~n19764 & n19768;
  assign n19770 = pi5  & n19769;
  assign n19771 = ~pi5  & ~n19769;
  assign n19772 = ~n19770 & ~n19771;
  assign n19773 = n19762 & ~n19772;
  assign n19774 = n75 & n12440;
  assign n19775 = n9491 & n13939;
  assign n19776 = n10469 & n12437;
  assign n19777 = n11031 & n12434;
  assign n19778 = ~n19774 & ~n19776;
  assign n19779 = ~n19777 & n19778;
  assign n19780 = ~n19775 & n19779;
  assign n19781 = ~pi5  & ~n19780;
  assign n19782 = pi5  & n19780;
  assign n19783 = ~n19781 & ~n19782;
  assign n19784 = n19394 & ~n19396;
  assign n19785 = ~n19397 & ~n19784;
  assign n19786 = ~n19783 & n19785;
  assign n19787 = ~n19783 & ~n19785;
  assign n19788 = n19783 & n19785;
  assign n19789 = ~n19787 & ~n19788;
  assign n19790 = n75 & n12443;
  assign n19791 = n9491 & n13702;
  assign n19792 = n10469 & n12440;
  assign n19793 = n11031 & n12437;
  assign n19794 = ~n19790 & ~n19792;
  assign n19795 = ~n19793 & n19794;
  assign n19796 = ~n19791 & n19795;
  assign n19797 = ~pi5  & ~n19796;
  assign n19798 = pi5  & n19796;
  assign n19799 = ~n19797 & ~n19798;
  assign n19800 = ~n19389 & n19392;
  assign n19801 = n19389 & ~n19392;
  assign n19802 = ~n19800 & ~n19801;
  assign n19803 = ~n19799 & ~n19802;
  assign n19804 = n75 & n12446;
  assign n19805 = n9491 & n14175;
  assign n19806 = n10469 & n12443;
  assign n19807 = n11031 & n12440;
  assign n19808 = ~n19804 & ~n19806;
  assign n19809 = ~n19807 & n19808;
  assign n19810 = ~n19805 & n19809;
  assign n19811 = ~pi5  & ~n19810;
  assign n19812 = pi5  & n19810;
  assign n19813 = ~n19811 & ~n19812;
  assign n19814 = n19384 & n19387;
  assign n19815 = ~n19388 & ~n19814;
  assign n19816 = ~n19813 & n19815;
  assign n19817 = ~n19813 & ~n19815;
  assign n19818 = n19813 & n19815;
  assign n19819 = ~n19817 & ~n19818;
  assign n19820 = n19187 & n19382;
  assign n19821 = ~n19383 & ~n19820;
  assign n19822 = n75 & n12449;
  assign n19823 = n9491 & n14325;
  assign n19824 = n10469 & n12446;
  assign n19825 = n11031 & n12443;
  assign n19826 = ~n19822 & ~n19824;
  assign n19827 = ~n19825 & n19826;
  assign n19828 = ~n19823 & n19827;
  assign n19829 = pi5  & n19828;
  assign n19830 = ~pi5  & ~n19828;
  assign n19831 = ~n19829 & ~n19830;
  assign n19832 = n19821 & ~n19831;
  assign n19833 = n19203 & n19380;
  assign n19834 = ~n19381 & ~n19833;
  assign n19835 = n75 & n12452;
  assign n19836 = n9491 & n14156;
  assign n19837 = n10469 & n12449;
  assign n19838 = n11031 & n12446;
  assign n19839 = ~n19835 & ~n19837;
  assign n19840 = ~n19838 & n19839;
  assign n19841 = ~n19836 & n19840;
  assign n19842 = pi5  & n19841;
  assign n19843 = ~pi5  & ~n19841;
  assign n19844 = ~n19842 & ~n19843;
  assign n19845 = n19834 & ~n19844;
  assign n19846 = n19376 & ~n19378;
  assign n19847 = ~n19379 & ~n19846;
  assign n19848 = n75 & n12455;
  assign n19849 = n9491 & n14442;
  assign n19850 = n10469 & n12452;
  assign n19851 = n11031 & n12449;
  assign n19852 = ~n19848 & ~n19850;
  assign n19853 = ~n19851 & n19852;
  assign n19854 = ~n19849 & n19853;
  assign n19855 = pi5  & n19854;
  assign n19856 = ~pi5  & ~n19854;
  assign n19857 = ~n19855 & ~n19856;
  assign n19858 = n19847 & ~n19857;
  assign n19859 = n75 & n12458;
  assign n19860 = n9491 & n14741;
  assign n19861 = n10469 & n12455;
  assign n19862 = n11031 & n12452;
  assign n19863 = ~n19859 & ~n19861;
  assign n19864 = ~n19862 & n19863;
  assign n19865 = ~n19860 & n19864;
  assign n19866 = ~pi5  & ~n19865;
  assign n19867 = pi5  & n19865;
  assign n19868 = ~n19866 & ~n19867;
  assign n19869 = n19372 & ~n19374;
  assign n19870 = ~n19375 & ~n19869;
  assign n19871 = ~n19868 & n19870;
  assign n19872 = ~n19868 & ~n19870;
  assign n19873 = n19868 & n19870;
  assign n19874 = ~n19872 & ~n19873;
  assign n19875 = n75 & n12461;
  assign n19876 = n9491 & n14756;
  assign n19877 = n10469 & n12458;
  assign n19878 = n11031 & n12455;
  assign n19879 = ~n19875 & ~n19877;
  assign n19880 = ~n19878 & n19879;
  assign n19881 = ~n19876 & n19880;
  assign n19882 = ~pi5  & ~n19881;
  assign n19883 = pi5  & n19881;
  assign n19884 = ~n19882 & ~n19883;
  assign n19885 = n19367 & n19370;
  assign n19886 = ~n19371 & ~n19885;
  assign n19887 = ~n19884 & n19886;
  assign n19888 = ~n19884 & ~n19886;
  assign n19889 = n19884 & n19886;
  assign n19890 = ~n19888 & ~n19889;
  assign n19891 = n75 & n12464;
  assign n19892 = n9491 & n14420;
  assign n19893 = n10469 & n12461;
  assign n19894 = n11031 & n12458;
  assign n19895 = ~n19891 & ~n19893;
  assign n19896 = ~n19894 & n19895;
  assign n19897 = ~n19892 & n19896;
  assign n19898 = ~pi5  & ~n19897;
  assign n19899 = pi5  & n19897;
  assign n19900 = ~n19898 & ~n19899;
  assign n19901 = ~n19362 & n19365;
  assign n19902 = n19362 & ~n19365;
  assign n19903 = ~n19901 & ~n19902;
  assign n19904 = ~n19900 & ~n19903;
  assign n19905 = n19272 & n19360;
  assign n19906 = ~n19361 & ~n19905;
  assign n19907 = n75 & n12467;
  assign n19908 = n9491 & n14789;
  assign n19909 = n10469 & n12464;
  assign n19910 = n11031 & n12461;
  assign n19911 = ~n19907 & ~n19909;
  assign n19912 = ~n19910 & n19911;
  assign n19913 = ~n19908 & n19912;
  assign n19914 = pi5  & n19913;
  assign n19915 = ~pi5  & ~n19913;
  assign n19916 = ~n19914 & ~n19915;
  assign n19917 = n19906 & ~n19916;
  assign n19918 = n19356 & ~n19358;
  assign n19919 = ~n19359 & ~n19918;
  assign n19920 = n75 & n12470;
  assign n19921 = n9491 & n14815;
  assign n19922 = n10469 & n12467;
  assign n19923 = n11031 & n12464;
  assign n19924 = ~n19920 & ~n19922;
  assign n19925 = ~n19923 & n19924;
  assign n19926 = ~n19921 & n19925;
  assign n19927 = pi5  & n19926;
  assign n19928 = ~pi5  & ~n19926;
  assign n19929 = ~n19927 & ~n19928;
  assign n19930 = n19919 & ~n19929;
  assign n19931 = n19303 & n19354;
  assign n19932 = ~n19355 & ~n19931;
  assign n19933 = n75 & n12473;
  assign n19934 = n9491 & n14839;
  assign n19935 = n10469 & n12470;
  assign n19936 = n11031 & n12467;
  assign n19937 = ~n19933 & ~n19935;
  assign n19938 = ~n19936 & n19937;
  assign n19939 = ~n19934 & n19938;
  assign n19940 = pi5  & n19939;
  assign n19941 = ~pi5  & ~n19939;
  assign n19942 = ~n19940 & ~n19941;
  assign n19943 = n19932 & ~n19942;
  assign n19944 = n75 & n12476;
  assign n19945 = n9491 & n14849;
  assign n19946 = n10469 & n12473;
  assign n19947 = n11031 & n12470;
  assign n19948 = ~n19944 & ~n19946;
  assign n19949 = ~n19947 & n19948;
  assign n19950 = ~n19945 & n19949;
  assign n19951 = ~pi5  & ~n19950;
  assign n19952 = pi5  & n19950;
  assign n19953 = ~n19951 & ~n19952;
  assign n19954 = n19350 & ~n19352;
  assign n19955 = ~n19353 & ~n19954;
  assign n19956 = ~n19953 & n19955;
  assign n19957 = ~n19953 & ~n19955;
  assign n19958 = n19953 & n19955;
  assign n19959 = ~n19957 & ~n19958;
  assign n19960 = n75 & n12479;
  assign n19961 = n9491 & n14922;
  assign n19962 = n10469 & n12476;
  assign n19963 = n11031 & n12473;
  assign n19964 = ~n19960 & ~n19962;
  assign n19965 = ~n19963 & n19964;
  assign n19966 = ~n19961 & n19965;
  assign n19967 = pi5  & n19966;
  assign n19968 = ~pi5  & ~n19966;
  assign n19969 = ~n19967 & ~n19968;
  assign n19970 = n19338 & n19348;
  assign n19971 = ~n19349 & ~n19970;
  assign n19972 = ~n19969 & n19971;
  assign n19973 = n75 & n12482;
  assign n19974 = n9491 & n14958;
  assign n19975 = n10469 & n12479;
  assign n19976 = n11031 & n12476;
  assign n19977 = ~n19973 & ~n19975;
  assign n19978 = ~n19976 & n19977;
  assign n19979 = ~n19974 & n19978;
  assign n19980 = ~pi5  & ~n19979;
  assign n19981 = pi5  & n19979;
  assign n19982 = ~n19980 & ~n19981;
  assign n19983 = pi8  & ~n19326;
  assign n19984 = n19333 & ~n19983;
  assign n19985 = ~n19333 & n19983;
  assign n19986 = ~n19984 & ~n19985;
  assign n19987 = ~n19982 & n19986;
  assign n19988 = ~n19982 & ~n19986;
  assign n19989 = n19982 & n19986;
  assign n19990 = ~n19988 & ~n19989;
  assign n19991 = n75 & n12485;
  assign n19992 = n9491 & n15001;
  assign n19993 = n10469 & n12482;
  assign n19994 = n11031 & n12479;
  assign n19995 = ~n19991 & ~n19993;
  assign n19996 = ~n19994 & n19995;
  assign n19997 = ~n19992 & n19996;
  assign n19998 = pi5  & n19997;
  assign n19999 = ~pi5  & ~n19997;
  assign n20000 = ~n19998 & ~n19999;
  assign n20001 = pi8  & n19319;
  assign n20002 = ~n19324 & n20001;
  assign n20003 = n19324 & ~n20001;
  assign n20004 = ~n20002 & ~n20003;
  assign n20005 = ~n20000 & n20004;
  assign n20006 = ~n70 & n12492;
  assign n20007 = n10469 & n12492;
  assign n20008 = n11031 & n12490;
  assign n20009 = n9491 & ~n15072;
  assign n20010 = ~n20007 & ~n20008;
  assign n20011 = ~n20009 & n20010;
  assign n20012 = pi5  & ~n20006;
  assign n20013 = n20011 & n20012;
  assign n20014 = n75 & n12492;
  assign n20015 = n9491 & ~n15113;
  assign n20016 = n10469 & n12490;
  assign n20017 = n11031 & n12485;
  assign n20018 = ~n20014 & ~n20016;
  assign n20019 = ~n20017 & n20018;
  assign n20020 = ~n20015 & n20019;
  assign n20021 = n20013 & n20020;
  assign n20022 = n19319 & n20021;
  assign n20023 = ~n19319 & n20021;
  assign n20024 = n19319 & ~n20021;
  assign n20025 = ~n20023 & ~n20024;
  assign n20026 = n75 & n12490;
  assign n20027 = n9491 & n15026;
  assign n20028 = n10469 & n12485;
  assign n20029 = n11031 & n12482;
  assign n20030 = ~n20026 & ~n20028;
  assign n20031 = ~n20029 & n20030;
  assign n20032 = ~n20027 & n20031;
  assign n20033 = pi5  & n20032;
  assign n20034 = ~pi5  & ~n20032;
  assign n20035 = ~n20033 & ~n20034;
  assign n20036 = ~n20025 & ~n20035;
  assign n20037 = ~n20022 & ~n20036;
  assign n20038 = n20000 & ~n20004;
  assign n20039 = ~n20005 & ~n20038;
  assign n20040 = ~n20037 & n20039;
  assign n20041 = ~n20005 & ~n20040;
  assign n20042 = ~n19990 & ~n20041;
  assign n20043 = ~n19987 & ~n20042;
  assign n20044 = n19969 & ~n19971;
  assign n20045 = ~n19972 & ~n20044;
  assign n20046 = ~n20043 & n20045;
  assign n20047 = ~n19972 & ~n20046;
  assign n20048 = ~n19959 & ~n20047;
  assign n20049 = ~n19956 & ~n20048;
  assign n20050 = n19932 & n19942;
  assign n20051 = ~n19932 & ~n19942;
  assign n20052 = ~n20050 & ~n20051;
  assign n20053 = ~n20049 & ~n20052;
  assign n20054 = ~n19943 & ~n20053;
  assign n20055 = n19919 & n19929;
  assign n20056 = ~n19919 & ~n19929;
  assign n20057 = ~n20055 & ~n20056;
  assign n20058 = ~n20054 & ~n20057;
  assign n20059 = ~n19930 & ~n20058;
  assign n20060 = ~n19906 & n19916;
  assign n20061 = ~n19917 & ~n20060;
  assign n20062 = ~n20059 & n20061;
  assign n20063 = ~n19917 & ~n20062;
  assign n20064 = n19900 & n19903;
  assign n20065 = ~n19904 & ~n20064;
  assign n20066 = ~n20063 & n20065;
  assign n20067 = ~n19904 & ~n20066;
  assign n20068 = ~n19890 & ~n20067;
  assign n20069 = ~n19887 & ~n20068;
  assign n20070 = ~n19874 & ~n20069;
  assign n20071 = ~n19871 & ~n20070;
  assign n20072 = n19847 & n19857;
  assign n20073 = ~n19847 & ~n19857;
  assign n20074 = ~n20072 & ~n20073;
  assign n20075 = ~n20071 & ~n20074;
  assign n20076 = ~n19858 & ~n20075;
  assign n20077 = n19834 & n19844;
  assign n20078 = ~n19834 & ~n19844;
  assign n20079 = ~n20077 & ~n20078;
  assign n20080 = ~n20076 & ~n20079;
  assign n20081 = ~n19845 & ~n20080;
  assign n20082 = ~n19821 & n19831;
  assign n20083 = ~n19832 & ~n20082;
  assign n20084 = ~n20081 & n20083;
  assign n20085 = ~n19832 & ~n20084;
  assign n20086 = ~n19819 & ~n20085;
  assign n20087 = ~n19816 & ~n20086;
  assign n20088 = n19799 & n19802;
  assign n20089 = ~n19803 & ~n20088;
  assign n20090 = ~n20087 & n20089;
  assign n20091 = ~n19803 & ~n20090;
  assign n20092 = ~n19789 & ~n20091;
  assign n20093 = ~n19786 & ~n20092;
  assign n20094 = n19762 & n19772;
  assign n20095 = ~n19762 & ~n19772;
  assign n20096 = ~n20094 & ~n20095;
  assign n20097 = ~n20093 & ~n20096;
  assign n20098 = ~n19773 & ~n20097;
  assign n20099 = n19749 & n19759;
  assign n20100 = ~n19749 & ~n19759;
  assign n20101 = ~n20099 & ~n20100;
  assign n20102 = ~n20098 & ~n20101;
  assign n20103 = ~n19760 & ~n20102;
  assign n20104 = ~n19736 & n19746;
  assign n20105 = ~n19747 & ~n20104;
  assign n20106 = ~n20103 & n20105;
  assign n20107 = ~n19747 & ~n20106;
  assign n20108 = n19730 & n19733;
  assign n20109 = ~n19734 & ~n20108;
  assign n20110 = ~n20107 & n20109;
  assign n20111 = ~n19734 & ~n20110;
  assign n20112 = ~n19720 & ~n20111;
  assign n20113 = ~n19717 & ~n20112;
  assign n20114 = ~n19704 & ~n20113;
  assign n20115 = ~n19701 & ~n20114;
  assign n20116 = n19677 & n19687;
  assign n20117 = ~n19677 & ~n19687;
  assign n20118 = ~n20116 & ~n20117;
  assign n20119 = ~n20115 & ~n20118;
  assign n20120 = ~n19688 & ~n20119;
  assign n20121 = ~n19664 & n19674;
  assign n20122 = ~n19675 & ~n20121;
  assign n20123 = ~n20120 & n20122;
  assign n20124 = ~n19675 & ~n20123;
  assign n20125 = n19658 & n19661;
  assign n20126 = ~n19662 & ~n20125;
  assign n20127 = ~n20124 & n20126;
  assign n20128 = ~n19662 & ~n20127;
  assign n20129 = n19644 & n19647;
  assign n20130 = ~n19648 & ~n20129;
  assign n20131 = ~n20128 & n20130;
  assign n20132 = ~n19648 & ~n20131;
  assign n20133 = ~n19634 & ~n20132;
  assign n20134 = ~n19631 & ~n20133;
  assign n20135 = ~n19618 & ~n20134;
  assign n20136 = ~n19615 & ~n20135;
  assign n20137 = ~n19602 & ~n20136;
  assign n20138 = ~n19599 & ~n20137;
  assign n20139 = n19582 & n19585;
  assign n20140 = ~n19586 & ~n20139;
  assign n20141 = ~n20138 & n20140;
  assign n20142 = ~n19586 & ~n20141;
  assign n20143 = n19568 & n19571;
  assign n20144 = ~n19572 & ~n20143;
  assign n20145 = ~n20142 & n20144;
  assign n20146 = ~n19572 & ~n20145;
  assign n20147 = n19554 & n19557;
  assign n20148 = ~n19558 & ~n20147;
  assign n20149 = ~n20146 & n20148;
  assign n20150 = ~n19558 & ~n20149;
  assign n20151 = n19540 & n19543;
  assign n20152 = ~n19544 & ~n20151;
  assign n20153 = ~n20150 & n20152;
  assign n20154 = ~n19544 & ~n20153;
  assign n20155 = n19512 & n19521;
  assign n20156 = ~n19522 & ~n20155;
  assign n20157 = ~n20154 & n20156;
  assign n20158 = n20154 & ~n20156;
  assign n20159 = ~n20157 & ~n20158;
  assign n20160 = n20150 & ~n20152;
  assign n20161 = ~n20153 & ~n20160;
  assign n20162 = n11672 & ~n12786;
  assign n20163 = n11056 & ~n13781;
  assign n20164 = n11055 & n13166;
  assign n20165 = n11661 & n13161;
  assign n20166 = ~n20162 & ~n20164;
  assign n20167 = ~n20165 & n20166;
  assign n20168 = ~n20163 & n20167;
  assign n20169 = pi2  & n20168;
  assign n20170 = ~pi2  & ~n20168;
  assign n20171 = ~n20169 & ~n20170;
  assign n20172 = n20161 & ~n20171;
  assign n20173 = n20146 & ~n20148;
  assign n20174 = ~n20149 & ~n20173;
  assign n20175 = n11672 & n13161;
  assign n20176 = n11056 & n13183;
  assign n20177 = n11661 & n13166;
  assign n20178 = n11055 & n13164;
  assign n20179 = ~n20177 & ~n20178;
  assign n20180 = ~n20175 & n20179;
  assign n20181 = ~n20176 & n20180;
  assign n20182 = pi2  & n20181;
  assign n20183 = ~pi2  & ~n20181;
  assign n20184 = ~n20182 & ~n20183;
  assign n20185 = n20174 & ~n20184;
  assign n20186 = n20142 & ~n20144;
  assign n20187 = ~n20145 & ~n20186;
  assign n20188 = n11055 & n12646;
  assign n20189 = n11056 & n13261;
  assign n20190 = n11661 & n13164;
  assign n20191 = n11672 & n13166;
  assign n20192 = ~n20188 & ~n20190;
  assign n20193 = ~n20191 & n20192;
  assign n20194 = ~n20189 & n20193;
  assign n20195 = pi2  & n20194;
  assign n20196 = ~pi2  & ~n20194;
  assign n20197 = ~n20195 & ~n20196;
  assign n20198 = n20187 & ~n20197;
  assign n20199 = n20138 & ~n20140;
  assign n20200 = ~n20141 & ~n20199;
  assign n20201 = n11055 & n12392;
  assign n20202 = n11056 & n13421;
  assign n20203 = n11661 & n12646;
  assign n20204 = n11672 & n13164;
  assign n20205 = ~n20201 & ~n20203;
  assign n20206 = ~n20204 & n20205;
  assign n20207 = ~n20202 & n20206;
  assign n20208 = pi2  & n20207;
  assign n20209 = ~pi2  & ~n20207;
  assign n20210 = ~n20208 & ~n20209;
  assign n20211 = n20200 & ~n20210;
  assign n20212 = n19602 & n20136;
  assign n20213 = ~n20137 & ~n20212;
  assign n20214 = n11055 & n12362;
  assign n20215 = n11056 & n12652;
  assign n20216 = n11661 & n12392;
  assign n20217 = n11672 & n12646;
  assign n20218 = ~n20214 & ~n20216;
  assign n20219 = ~n20217 & n20218;
  assign n20220 = ~n20215 & n20219;
  assign n20221 = pi2  & n20220;
  assign n20222 = ~pi2  & ~n20220;
  assign n20223 = ~n20221 & ~n20222;
  assign n20224 = n20213 & ~n20223;
  assign n20225 = n19618 & n20134;
  assign n20226 = ~n20135 & ~n20225;
  assign n20227 = n11055 & n12395;
  assign n20228 = n11056 & n13144;
  assign n20229 = n11661 & n12362;
  assign n20230 = n11672 & n12392;
  assign n20231 = ~n20227 & ~n20229;
  assign n20232 = ~n20230 & n20231;
  assign n20233 = ~n20228 & n20232;
  assign n20234 = pi2  & n20233;
  assign n20235 = ~pi2  & ~n20233;
  assign n20236 = ~n20234 & ~n20235;
  assign n20237 = n20226 & ~n20236;
  assign n20238 = n19634 & n20132;
  assign n20239 = ~n20133 & ~n20238;
  assign n20240 = n11055 & n12398;
  assign n20241 = n11056 & n13245;
  assign n20242 = n11661 & n12395;
  assign n20243 = n11672 & n12362;
  assign n20244 = ~n20240 & ~n20242;
  assign n20245 = ~n20243 & n20244;
  assign n20246 = ~n20241 & n20245;
  assign n20247 = pi2  & n20246;
  assign n20248 = ~pi2  & ~n20246;
  assign n20249 = ~n20247 & ~n20248;
  assign n20250 = n20239 & ~n20249;
  assign n20251 = n20128 & ~n20130;
  assign n20252 = ~n20131 & ~n20251;
  assign n20253 = n11055 & n12401;
  assign n20254 = n11056 & n13108;
  assign n20255 = n11661 & n12398;
  assign n20256 = n11672 & n12395;
  assign n20257 = ~n20253 & ~n20255;
  assign n20258 = ~n20256 & n20257;
  assign n20259 = ~n20254 & n20258;
  assign n20260 = pi2  & n20259;
  assign n20261 = ~pi2  & ~n20259;
  assign n20262 = ~n20260 & ~n20261;
  assign n20263 = n20252 & ~n20262;
  assign n20264 = n20124 & ~n20126;
  assign n20265 = ~n20127 & ~n20264;
  assign n20266 = n11055 & n12404;
  assign n20267 = n11056 & n13128;
  assign n20268 = n11661 & n12401;
  assign n20269 = n11672 & n12398;
  assign n20270 = ~n20266 & ~n20268;
  assign n20271 = ~n20269 & n20270;
  assign n20272 = ~n20267 & n20271;
  assign n20273 = pi2  & n20272;
  assign n20274 = ~pi2  & ~n20272;
  assign n20275 = ~n20273 & ~n20274;
  assign n20276 = n20265 & ~n20275;
  assign n20277 = n20265 & n20275;
  assign n20278 = ~n20265 & ~n20275;
  assign n20279 = ~n20277 & ~n20278;
  assign n20280 = n20120 & ~n20122;
  assign n20281 = ~n20123 & ~n20280;
  assign n20282 = n20115 & n20118;
  assign n20283 = ~n20119 & ~n20282;
  assign n20284 = n11055 & n12413;
  assign n20285 = n11056 & n12891;
  assign n20286 = n11661 & n12410;
  assign n20287 = n11672 & n12407;
  assign n20288 = ~n20284 & ~n20286;
  assign n20289 = ~n20287 & n20288;
  assign n20290 = ~n20285 & n20289;
  assign n20291 = pi2  & n20290;
  assign n20292 = ~pi2  & ~n20290;
  assign n20293 = ~n20291 & ~n20292;
  assign n20294 = n11055 & n12416;
  assign n20295 = n11056 & n12843;
  assign n20296 = n11661 & n12413;
  assign n20297 = n11672 & n12410;
  assign n20298 = ~n20294 & ~n20296;
  assign n20299 = ~n20297 & n20298;
  assign n20300 = ~n20295 & n20299;
  assign n20301 = pi2  & n20300;
  assign n20302 = ~pi2  & ~n20300;
  assign n20303 = ~n20301 & ~n20302;
  assign n20304 = n11055 & n12419;
  assign n20305 = n11056 & n12908;
  assign n20306 = n11661 & n12416;
  assign n20307 = n11672 & n12413;
  assign n20308 = ~n20304 & ~n20306;
  assign n20309 = ~n20307 & n20308;
  assign n20310 = ~n20305 & n20309;
  assign n20311 = pi2  & n20310;
  assign n20312 = ~pi2  & ~n20310;
  assign n20313 = ~n20311 & ~n20312;
  assign n20314 = n20103 & ~n20105;
  assign n20315 = ~n20106 & ~n20314;
  assign n20316 = n20098 & n20101;
  assign n20317 = ~n20102 & ~n20316;
  assign n20318 = n20093 & n20096;
  assign n20319 = ~n20097 & ~n20318;
  assign n20320 = n11055 & n12431;
  assign n20321 = n11056 & n13356;
  assign n20322 = n11661 & n12428;
  assign n20323 = n11672 & n12425;
  assign n20324 = ~n20320 & ~n20322;
  assign n20325 = ~n20323 & n20324;
  assign n20326 = ~n20321 & n20325;
  assign n20327 = pi2  & n20326;
  assign n20328 = ~pi2  & ~n20326;
  assign n20329 = ~n20327 & ~n20328;
  assign n20330 = n11055 & n12434;
  assign n20331 = n11056 & n13546;
  assign n20332 = n11661 & n12431;
  assign n20333 = n11672 & n12428;
  assign n20334 = ~n20330 & ~n20332;
  assign n20335 = ~n20333 & n20334;
  assign n20336 = ~n20331 & n20335;
  assign n20337 = pi2  & n20336;
  assign n20338 = ~pi2  & ~n20336;
  assign n20339 = ~n20337 & ~n20338;
  assign n20340 = n11055 & n12437;
  assign n20341 = n11056 & n13564;
  assign n20342 = n11661 & n12434;
  assign n20343 = n11672 & n12431;
  assign n20344 = ~n20340 & ~n20342;
  assign n20345 = ~n20343 & n20344;
  assign n20346 = ~n20341 & n20345;
  assign n20347 = pi2  & n20346;
  assign n20348 = ~pi2  & ~n20346;
  assign n20349 = ~n20347 & ~n20348;
  assign n20350 = n20081 & ~n20083;
  assign n20351 = ~n20084 & ~n20350;
  assign n20352 = n20076 & n20079;
  assign n20353 = ~n20080 & ~n20352;
  assign n20354 = n20071 & n20074;
  assign n20355 = ~n20075 & ~n20354;
  assign n20356 = n11055 & n12449;
  assign n20357 = n11056 & n14325;
  assign n20358 = n11661 & n12446;
  assign n20359 = n11672 & n12443;
  assign n20360 = ~n20356 & ~n20358;
  assign n20361 = ~n20359 & n20360;
  assign n20362 = ~n20357 & n20361;
  assign n20363 = pi2  & n20362;
  assign n20364 = ~pi2  & ~n20362;
  assign n20365 = ~n20363 & ~n20364;
  assign n20366 = n11055 & n12452;
  assign n20367 = n11056 & n14156;
  assign n20368 = n11661 & n12449;
  assign n20369 = n11672 & n12446;
  assign n20370 = ~n20366 & ~n20368;
  assign n20371 = ~n20369 & n20370;
  assign n20372 = ~n20367 & n20371;
  assign n20373 = pi2  & n20372;
  assign n20374 = ~pi2  & ~n20372;
  assign n20375 = ~n20373 & ~n20374;
  assign n20376 = n11055 & n12455;
  assign n20377 = n11056 & n14442;
  assign n20378 = n11661 & n12452;
  assign n20379 = n11672 & n12449;
  assign n20380 = ~n20376 & ~n20378;
  assign n20381 = ~n20379 & n20380;
  assign n20382 = ~n20377 & n20381;
  assign n20383 = pi2  & n20382;
  assign n20384 = ~pi2  & ~n20382;
  assign n20385 = ~n20383 & ~n20384;
  assign n20386 = n20059 & ~n20061;
  assign n20387 = ~n20062 & ~n20386;
  assign n20388 = n20054 & n20057;
  assign n20389 = ~n20058 & ~n20388;
  assign n20390 = n20049 & n20052;
  assign n20391 = ~n20053 & ~n20390;
  assign n20392 = n11055 & n12467;
  assign n20393 = n11056 & n14789;
  assign n20394 = n11661 & n12464;
  assign n20395 = n11672 & n12461;
  assign n20396 = ~n20392 & ~n20394;
  assign n20397 = ~n20395 & n20396;
  assign n20398 = ~n20393 & n20397;
  assign n20399 = pi2  & n20398;
  assign n20400 = ~pi2  & ~n20398;
  assign n20401 = ~n20399 & ~n20400;
  assign n20402 = n11055 & n12470;
  assign n20403 = n11056 & n14815;
  assign n20404 = n11661 & n12467;
  assign n20405 = n11672 & n12464;
  assign n20406 = ~n20402 & ~n20404;
  assign n20407 = ~n20405 & n20406;
  assign n20408 = ~n20403 & n20407;
  assign n20409 = pi2  & n20408;
  assign n20410 = ~pi2  & ~n20408;
  assign n20411 = ~n20409 & ~n20410;
  assign n20412 = n11055 & n12473;
  assign n20413 = n11056 & n14839;
  assign n20414 = n11661 & n12470;
  assign n20415 = n11672 & n12467;
  assign n20416 = ~n20412 & ~n20414;
  assign n20417 = ~n20415 & n20416;
  assign n20418 = ~n20413 & n20417;
  assign n20419 = pi2  & n20418;
  assign n20420 = ~pi2  & ~n20418;
  assign n20421 = ~n20419 & ~n20420;
  assign n20422 = n20037 & ~n20039;
  assign n20423 = ~n20040 & ~n20422;
  assign n20424 = n11055 & n12479;
  assign n20425 = n11056 & n14922;
  assign n20426 = n11661 & n12476;
  assign n20427 = n11672 & n12473;
  assign n20428 = ~n20424 & ~n20426;
  assign n20429 = ~n20427 & n20428;
  assign n20430 = ~n20425 & n20429;
  assign n20431 = pi2  & n20430;
  assign n20432 = ~pi2  & ~n20430;
  assign n20433 = ~n20431 & ~n20432;
  assign n20434 = pi5  & ~n20013;
  assign n20435 = n20020 & ~n20434;
  assign n20436 = ~n20020 & n20434;
  assign n20437 = ~n20435 & ~n20436;
  assign n20438 = n11055 & n12485;
  assign n20439 = n11056 & n15001;
  assign n20440 = n11661 & n12482;
  assign n20441 = n11672 & n12479;
  assign n20442 = ~n20438 & ~n20440;
  assign n20443 = ~n20441 & n20442;
  assign n20444 = ~n20439 & n20443;
  assign n20445 = pi2  & n20444;
  assign n20446 = ~pi2  & ~n20444;
  assign n20447 = ~n20445 & ~n20446;
  assign n20448 = ~n11054 & n12492;
  assign n20449 = n11055 & n12492;
  assign n20450 = n11661 & n12490;
  assign n20451 = n11672 & n12485;
  assign n20452 = ~n20449 & ~n20450;
  assign n20453 = ~n20451 & n20452;
  assign n20454 = pi2  & ~n20453;
  assign n20455 = ~n12485 & n15072;
  assign n20456 = n11911 & ~n20455;
  assign n20457 = pi2  & n11672;
  assign n20458 = n12490 & n20457;
  assign n20459 = pi2  & ~n20448;
  assign n20460 = ~n20458 & n20459;
  assign n20461 = ~n20456 & n20460;
  assign n20462 = ~n20454 & n20461;
  assign n20463 = ~n20006 & ~n20462;
  assign n20464 = n20006 & n20462;
  assign n20465 = n11055 & n12490;
  assign n20466 = n11056 & n15026;
  assign n20467 = n11661 & n12485;
  assign n20468 = n11672 & n12482;
  assign n20469 = ~n20465 & ~n20467;
  assign n20470 = ~n20468 & n20469;
  assign n20471 = ~n20466 & n20470;
  assign n20472 = pi2  & ~n20471;
  assign n20473 = ~pi2  & n20471;
  assign n20474 = ~n20472 & ~n20473;
  assign n20475 = ~n20464 & ~n20474;
  assign n20476 = ~n20463 & ~n20475;
  assign n20477 = ~n20447 & n20476;
  assign n20478 = n20447 & ~n20476;
  assign n20479 = pi5  & n20006;
  assign n20480 = ~n20011 & n20479;
  assign n20481 = n20011 & ~n20479;
  assign n20482 = ~n20480 & ~n20481;
  assign n20483 = ~n20478 & n20482;
  assign n20484 = ~n20477 & ~n20483;
  assign n20485 = n20437 & ~n20484;
  assign n20486 = ~n20437 & n20484;
  assign n20487 = n11055 & n12482;
  assign n20488 = n11056 & n14958;
  assign n20489 = n11661 & n12479;
  assign n20490 = n11672 & n12476;
  assign n20491 = ~n20487 & ~n20489;
  assign n20492 = ~n20490 & n20491;
  assign n20493 = ~n20488 & n20492;
  assign n20494 = pi2  & ~n20493;
  assign n20495 = ~pi2  & n20493;
  assign n20496 = ~n20494 & ~n20495;
  assign n20497 = ~n20486 & n20496;
  assign n20498 = ~n20485 & ~n20497;
  assign n20499 = ~n20433 & ~n20498;
  assign n20500 = n20433 & n20498;
  assign n20501 = n20025 & n20035;
  assign n20502 = ~n20036 & ~n20501;
  assign n20503 = ~n20500 & n20502;
  assign n20504 = ~n20499 & ~n20503;
  assign n20505 = n20423 & ~n20504;
  assign n20506 = ~n20423 & n20504;
  assign n20507 = n11055 & n12476;
  assign n20508 = n11056 & n14849;
  assign n20509 = n11661 & n12473;
  assign n20510 = n11672 & n12470;
  assign n20511 = ~n20507 & ~n20509;
  assign n20512 = ~n20510 & n20511;
  assign n20513 = ~n20508 & n20512;
  assign n20514 = pi2  & ~n20513;
  assign n20515 = ~pi2  & n20513;
  assign n20516 = ~n20514 & ~n20515;
  assign n20517 = ~n20506 & n20516;
  assign n20518 = ~n20505 & ~n20517;
  assign n20519 = ~n20421 & ~n20518;
  assign n20520 = n20421 & n20518;
  assign n20521 = n19990 & n20041;
  assign n20522 = ~n20042 & ~n20521;
  assign n20523 = ~n20520 & n20522;
  assign n20524 = ~n20519 & ~n20523;
  assign n20525 = ~n20411 & ~n20524;
  assign n20526 = n20411 & n20524;
  assign n20527 = n20043 & ~n20045;
  assign n20528 = ~n20046 & ~n20527;
  assign n20529 = ~n20526 & n20528;
  assign n20530 = ~n20525 & ~n20529;
  assign n20531 = ~n20401 & ~n20530;
  assign n20532 = n20401 & n20530;
  assign n20533 = n19959 & n20047;
  assign n20534 = ~n20048 & ~n20533;
  assign n20535 = ~n20532 & n20534;
  assign n20536 = ~n20531 & ~n20535;
  assign n20537 = n20391 & ~n20536;
  assign n20538 = ~n20391 & n20536;
  assign n20539 = n11055 & n12464;
  assign n20540 = n11056 & n14420;
  assign n20541 = n11661 & n12461;
  assign n20542 = n11672 & n12458;
  assign n20543 = ~n20539 & ~n20541;
  assign n20544 = ~n20542 & n20543;
  assign n20545 = ~n20540 & n20544;
  assign n20546 = pi2  & ~n20545;
  assign n20547 = ~pi2  & n20545;
  assign n20548 = ~n20546 & ~n20547;
  assign n20549 = ~n20538 & n20548;
  assign n20550 = ~n20537 & ~n20549;
  assign n20551 = n20389 & ~n20550;
  assign n20552 = ~n20389 & n20550;
  assign n20553 = n11055 & n12461;
  assign n20554 = n11056 & n14756;
  assign n20555 = n11661 & n12458;
  assign n20556 = n11672 & n12455;
  assign n20557 = ~n20553 & ~n20555;
  assign n20558 = ~n20556 & n20557;
  assign n20559 = ~n20554 & n20558;
  assign n20560 = pi2  & ~n20559;
  assign n20561 = ~pi2  & n20559;
  assign n20562 = ~n20560 & ~n20561;
  assign n20563 = ~n20552 & n20562;
  assign n20564 = ~n20551 & ~n20563;
  assign n20565 = n20387 & ~n20564;
  assign n20566 = ~n20387 & n20564;
  assign n20567 = n11055 & n12458;
  assign n20568 = n11056 & n14741;
  assign n20569 = n11661 & n12455;
  assign n20570 = n11672 & n12452;
  assign n20571 = ~n20567 & ~n20569;
  assign n20572 = ~n20570 & n20571;
  assign n20573 = ~n20568 & n20572;
  assign n20574 = pi2  & ~n20573;
  assign n20575 = ~pi2  & n20573;
  assign n20576 = ~n20574 & ~n20575;
  assign n20577 = ~n20566 & n20576;
  assign n20578 = ~n20565 & ~n20577;
  assign n20579 = ~n20385 & ~n20578;
  assign n20580 = n20385 & n20578;
  assign n20581 = n20063 & ~n20065;
  assign n20582 = ~n20066 & ~n20581;
  assign n20583 = ~n20580 & n20582;
  assign n20584 = ~n20579 & ~n20583;
  assign n20585 = ~n20375 & ~n20584;
  assign n20586 = n20375 & n20584;
  assign n20587 = n19890 & n20067;
  assign n20588 = ~n20068 & ~n20587;
  assign n20589 = ~n20586 & n20588;
  assign n20590 = ~n20585 & ~n20589;
  assign n20591 = ~n20365 & ~n20590;
  assign n20592 = n20365 & n20590;
  assign n20593 = n19874 & n20069;
  assign n20594 = ~n20070 & ~n20593;
  assign n20595 = ~n20592 & n20594;
  assign n20596 = ~n20591 & ~n20595;
  assign n20597 = n20355 & ~n20596;
  assign n20598 = ~n20355 & n20596;
  assign n20599 = n11055 & n12446;
  assign n20600 = n11056 & n14175;
  assign n20601 = n11661 & n12443;
  assign n20602 = n11672 & n12440;
  assign n20603 = ~n20599 & ~n20601;
  assign n20604 = ~n20602 & n20603;
  assign n20605 = ~n20600 & n20604;
  assign n20606 = pi2  & ~n20605;
  assign n20607 = ~pi2  & n20605;
  assign n20608 = ~n20606 & ~n20607;
  assign n20609 = ~n20598 & n20608;
  assign n20610 = ~n20597 & ~n20609;
  assign n20611 = n20353 & ~n20610;
  assign n20612 = ~n20353 & n20610;
  assign n20613 = n11055 & n12443;
  assign n20614 = n11056 & n13702;
  assign n20615 = n11661 & n12440;
  assign n20616 = n11672 & n12437;
  assign n20617 = ~n20613 & ~n20615;
  assign n20618 = ~n20616 & n20617;
  assign n20619 = ~n20614 & n20618;
  assign n20620 = pi2  & ~n20619;
  assign n20621 = ~pi2  & n20619;
  assign n20622 = ~n20620 & ~n20621;
  assign n20623 = ~n20612 & n20622;
  assign n20624 = ~n20611 & ~n20623;
  assign n20625 = n20351 & ~n20624;
  assign n20626 = ~n20351 & n20624;
  assign n20627 = n11055 & n12440;
  assign n20628 = n11056 & n13939;
  assign n20629 = n11661 & n12437;
  assign n20630 = n11672 & n12434;
  assign n20631 = ~n20627 & ~n20629;
  assign n20632 = ~n20630 & n20631;
  assign n20633 = ~n20628 & n20632;
  assign n20634 = pi2  & ~n20633;
  assign n20635 = ~pi2  & n20633;
  assign n20636 = ~n20634 & ~n20635;
  assign n20637 = ~n20626 & n20636;
  assign n20638 = ~n20625 & ~n20637;
  assign n20639 = ~n20349 & ~n20638;
  assign n20640 = n20349 & n20638;
  assign n20641 = n19819 & n20085;
  assign n20642 = ~n20086 & ~n20641;
  assign n20643 = ~n20640 & n20642;
  assign n20644 = ~n20639 & ~n20643;
  assign n20645 = ~n20339 & ~n20644;
  assign n20646 = n20339 & n20644;
  assign n20647 = n20087 & ~n20089;
  assign n20648 = ~n20090 & ~n20647;
  assign n20649 = ~n20646 & n20648;
  assign n20650 = ~n20645 & ~n20649;
  assign n20651 = ~n20329 & ~n20650;
  assign n20652 = n20329 & n20650;
  assign n20653 = n19789 & n20091;
  assign n20654 = ~n20092 & ~n20653;
  assign n20655 = ~n20652 & n20654;
  assign n20656 = ~n20651 & ~n20655;
  assign n20657 = n20319 & ~n20656;
  assign n20658 = ~n20319 & n20656;
  assign n20659 = n11055 & n12428;
  assign n20660 = n11056 & n13371;
  assign n20661 = n11661 & n12425;
  assign n20662 = n11672 & n12422;
  assign n20663 = ~n20659 & ~n20661;
  assign n20664 = ~n20662 & n20663;
  assign n20665 = ~n20660 & n20664;
  assign n20666 = pi2  & ~n20665;
  assign n20667 = ~pi2  & n20665;
  assign n20668 = ~n20666 & ~n20667;
  assign n20669 = ~n20658 & n20668;
  assign n20670 = ~n20657 & ~n20669;
  assign n20671 = n20317 & ~n20670;
  assign n20672 = ~n20317 & n20670;
  assign n20673 = n11055 & n12425;
  assign n20674 = n11056 & n13010;
  assign n20675 = n11661 & n12422;
  assign n20676 = n11672 & n12419;
  assign n20677 = ~n20673 & ~n20675;
  assign n20678 = ~n20676 & n20677;
  assign n20679 = ~n20674 & n20678;
  assign n20680 = pi2  & ~n20679;
  assign n20681 = ~pi2  & n20679;
  assign n20682 = ~n20680 & ~n20681;
  assign n20683 = ~n20672 & n20682;
  assign n20684 = ~n20671 & ~n20683;
  assign n20685 = n20315 & ~n20684;
  assign n20686 = ~n20315 & n20684;
  assign n20687 = n11055 & n12422;
  assign n20688 = n11056 & n13201;
  assign n20689 = n11661 & n12419;
  assign n20690 = n11672 & n12416;
  assign n20691 = ~n20687 & ~n20689;
  assign n20692 = ~n20690 & n20691;
  assign n20693 = ~n20688 & n20692;
  assign n20694 = pi2  & ~n20693;
  assign n20695 = ~pi2  & n20693;
  assign n20696 = ~n20694 & ~n20695;
  assign n20697 = ~n20686 & n20696;
  assign n20698 = ~n20685 & ~n20697;
  assign n20699 = ~n20313 & ~n20698;
  assign n20700 = n20313 & n20698;
  assign n20701 = n20107 & ~n20109;
  assign n20702 = ~n20110 & ~n20701;
  assign n20703 = ~n20700 & n20702;
  assign n20704 = ~n20699 & ~n20703;
  assign n20705 = ~n20303 & ~n20704;
  assign n20706 = n20303 & n20704;
  assign n20707 = n19720 & n20111;
  assign n20708 = ~n20112 & ~n20707;
  assign n20709 = ~n20706 & n20708;
  assign n20710 = ~n20705 & ~n20709;
  assign n20711 = ~n20293 & ~n20710;
  assign n20712 = n20293 & n20710;
  assign n20713 = n19704 & n20113;
  assign n20714 = ~n20114 & ~n20713;
  assign n20715 = ~n20712 & n20714;
  assign n20716 = ~n20711 & ~n20715;
  assign n20717 = n20283 & ~n20716;
  assign n20718 = ~n20283 & n20716;
  assign n20719 = n11055 & n12410;
  assign n20720 = n11056 & n13093;
  assign n20721 = n11661 & n12407;
  assign n20722 = n11672 & n12404;
  assign n20723 = ~n20719 & ~n20721;
  assign n20724 = ~n20722 & n20723;
  assign n20725 = ~n20720 & n20724;
  assign n20726 = pi2  & ~n20725;
  assign n20727 = ~pi2  & n20725;
  assign n20728 = ~n20726 & ~n20727;
  assign n20729 = ~n20718 & n20728;
  assign n20730 = ~n20717 & ~n20729;
  assign n20731 = n20281 & ~n20730;
  assign n20732 = ~n20281 & n20730;
  assign n20733 = n11055 & n12407;
  assign n20734 = n11056 & n13035;
  assign n20735 = n11661 & n12404;
  assign n20736 = n11672 & n12401;
  assign n20737 = ~n20733 & ~n20735;
  assign n20738 = ~n20736 & n20737;
  assign n20739 = ~n20734 & n20738;
  assign n20740 = pi2  & ~n20739;
  assign n20741 = ~pi2  & n20739;
  assign n20742 = ~n20740 & ~n20741;
  assign n20743 = ~n20732 & n20742;
  assign n20744 = ~n20731 & ~n20743;
  assign n20745 = ~n20279 & ~n20744;
  assign n20746 = ~n20276 & ~n20745;
  assign n20747 = ~n20252 & n20262;
  assign n20748 = ~n20263 & ~n20747;
  assign n20749 = ~n20746 & n20748;
  assign n20750 = ~n20263 & ~n20749;
  assign n20751 = ~n20239 & n20249;
  assign n20752 = ~n20250 & ~n20751;
  assign n20753 = ~n20750 & n20752;
  assign n20754 = ~n20250 & ~n20753;
  assign n20755 = ~n20226 & n20236;
  assign n20756 = ~n20237 & ~n20755;
  assign n20757 = ~n20754 & n20756;
  assign n20758 = ~n20237 & ~n20757;
  assign n20759 = ~n20213 & n20223;
  assign n20760 = ~n20224 & ~n20759;
  assign n20761 = ~n20758 & n20760;
  assign n20762 = ~n20224 & ~n20761;
  assign n20763 = ~n20200 & n20210;
  assign n20764 = ~n20211 & ~n20763;
  assign n20765 = ~n20762 & n20764;
  assign n20766 = ~n20211 & ~n20765;
  assign n20767 = ~n20187 & n20197;
  assign n20768 = ~n20198 & ~n20767;
  assign n20769 = ~n20766 & n20768;
  assign n20770 = ~n20198 & ~n20769;
  assign n20771 = ~n20174 & n20184;
  assign n20772 = ~n20185 & ~n20771;
  assign n20773 = ~n20770 & n20772;
  assign n20774 = ~n20185 & ~n20773;
  assign n20775 = ~n20161 & n20171;
  assign n20776 = ~n20172 & ~n20775;
  assign n20777 = ~n20774 & n20776;
  assign n20778 = ~n20172 & ~n20777;
  assign n20779 = n20159 & ~n20778;
  assign n20780 = ~n20157 & ~n20779;
  assign n20781 = n19530 & ~n20780;
  assign n20782 = ~n19528 & ~n20781;
  assign n20783 = n19496 & ~n20782;
  assign n20784 = ~n19494 & ~n20783;
  assign n20785 = n18883 & ~n20784;
  assign n20786 = ~n18881 & ~n20785;
  assign n20787 = ~n17771 & n18304;
  assign n20788 = ~n18305 & ~n20787;
  assign n20789 = ~n20786 & n20788;
  assign n20790 = ~n18305 & ~n20789;
  assign n20791 = ~n17769 & ~n20790;
  assign n20792 = ~n17766 & ~n20791;
  assign n20793 = n17261 & ~n20792;
  assign n20794 = ~n17259 & ~n20793;
  assign n20795 = ~n16361 & n16789;
  assign n20796 = ~n16790 & ~n20795;
  assign n20797 = ~n20794 & n20796;
  assign n20798 = ~n16790 & ~n20797;
  assign n20799 = ~n16359 & ~n20798;
  assign n20800 = ~n16356 & ~n20799;
  assign n20801 = n15957 & ~n20800;
  assign n20802 = ~n15955 & ~n20801;
  assign n20803 = ~n15447 & n15599;
  assign n20804 = ~n15600 & ~n20803;
  assign n20805 = ~n20802 & n20804;
  assign n20806 = ~n15600 & ~n20805;
  assign n20807 = ~n15445 & ~n20806;
  assign n20808 = ~n15442 & ~n20807;
  assign n20809 = n15282 & ~n20808;
  assign n20810 = ~n15280 & ~n20809;
  assign n20811 = ~n14555 & n14690;
  assign n20812 = ~n14691 & ~n20811;
  assign n20813 = ~n20810 & n20812;
  assign n20814 = ~n14691 & ~n20813;
  assign n20815 = ~n14553 & ~n20814;
  assign n20816 = ~n14550 & ~n20815;
  assign n20817 = n14271 & ~n20816;
  assign n20818 = ~n14269 & ~n20817;
  assign n20819 = ~n13905 & n14034;
  assign n20820 = ~n14035 & ~n20819;
  assign n20821 = ~n20818 & n20820;
  assign n20822 = ~n14035 & ~n20821;
  assign n20823 = ~n13903 & ~n20822;
  assign n20824 = ~n13900 & ~n20823;
  assign n20825 = n13795 & ~n20824;
  assign n20826 = ~n13793 & ~n20825;
  assign n20827 = ~n13278 & n13440;
  assign n20828 = ~n13441 & ~n20827;
  assign n20829 = ~n20826 & n20828;
  assign n20830 = ~n13441 & ~n20829;
  assign n20831 = ~n13192 & ~n13272;
  assign n20832 = ~n13276 & ~n20831;
  assign n20833 = n5130 & ~n12786;
  assign n20834 = n5045 & ~n13781;
  assign n20835 = n5044 & n13166;
  assign n20836 = n5109 & n13161;
  assign n20837 = ~n20833 & ~n20835;
  assign n20838 = ~n20836 & n20837;
  assign n20839 = ~n20834 & n20838;
  assign n20840 = pi23  & n20839;
  assign n20841 = ~pi23  & ~n20839;
  assign n20842 = ~n20840 & ~n20841;
  assign n20843 = ~n12661 & n13120;
  assign n20844 = ~n13156 & ~n20843;
  assign n20845 = n86 & n12392;
  assign n20846 = n4420 & n13421;
  assign n20847 = n4600 & n12646;
  assign n20848 = n4615 & n13164;
  assign n20849 = ~n20845 & ~n20847;
  assign n20850 = ~n20848 & n20849;
  assign n20851 = ~n20846 & n20850;
  assign n20852 = pi26  & n20851;
  assign n20853 = ~pi26  & ~n20851;
  assign n20854 = ~n20852 & ~n20853;
  assign n20855 = ~n13082 & ~n13085;
  assign n20856 = n12736 & ~n20855;
  assign n20857 = ~n12736 & n20855;
  assign n20858 = ~n20856 & ~n20857;
  assign n20859 = n3692 & n12404;
  assign n20860 = n880 & n13035;
  assign n20861 = n748 & n12407;
  assign n20862 = n3694 & n12401;
  assign n20863 = ~n20859 & ~n20861;
  assign n20864 = ~n20862 & n20863;
  assign n20865 = ~n20860 & n20864;
  assign n20866 = n20858 & ~n20865;
  assign n20867 = ~n20858 & n20865;
  assign n20868 = ~n20866 & ~n20867;
  assign n20869 = ~n13088 & n13099;
  assign n20870 = ~n13089 & ~n20869;
  assign n20871 = n20868 & n20870;
  assign n20872 = ~n20868 & ~n20870;
  assign n20873 = ~n20871 & ~n20872;
  assign n20874 = n3810 & n12398;
  assign n20875 = n3886 & n13245;
  assign n20876 = n3884 & n12395;
  assign n20877 = n4380 & n12362;
  assign n20878 = ~n20874 & ~n20876;
  assign n20879 = ~n20877 & n20878;
  assign n20880 = ~n20875 & n20879;
  assign n20881 = pi29  & n20880;
  assign n20882 = ~pi29  & ~n20880;
  assign n20883 = ~n20881 & ~n20882;
  assign n20884 = n20873 & ~n20883;
  assign n20885 = ~n20873 & n20883;
  assign n20886 = ~n20884 & ~n20885;
  assign n20887 = ~n13104 & ~n13117;
  assign n20888 = ~n13103 & ~n20887;
  assign n20889 = n20886 & ~n20888;
  assign n20890 = ~n20886 & n20888;
  assign n20891 = ~n20889 & ~n20890;
  assign n20892 = ~n20854 & n20891;
  assign n20893 = n20854 & ~n20891;
  assign n20894 = ~n20892 & ~n20893;
  assign n20895 = ~n20844 & n20894;
  assign n20896 = n20844 & ~n20894;
  assign n20897 = ~n20895 & ~n20896;
  assign n20898 = ~n20842 & ~n20897;
  assign n20899 = n20842 & n20897;
  assign n20900 = ~n20898 & ~n20899;
  assign n20901 = ~n20832 & ~n20900;
  assign n20902 = n20832 & n20900;
  assign n20903 = ~n20901 & ~n20902;
  assign n20904 = ~n20830 & n20903;
  assign n20905 = n20830 & ~n20903;
  assign n20906 = ~n20904 & ~n20905;
  assign n20907 = n75 & n20906;
  assign n20908 = n5045 & ~n13280;
  assign n20909 = n5044 & ~n13160;
  assign n20910 = ~n5109 & ~n5130;
  assign n20911 = ~n20909 & n20910;
  assign n20912 = ~n12786 & ~n20911;
  assign n20913 = ~n20908 & ~n20912;
  assign n20914 = pi23  & n20913;
  assign n20915 = ~pi23  & ~n20913;
  assign n20916 = ~n20914 & ~n20915;
  assign n20917 = ~n20854 & ~n20890;
  assign n20918 = ~n20889 & ~n20917;
  assign n20919 = ~n20916 & ~n20918;
  assign n20920 = n20916 & n20918;
  assign n20921 = ~n20919 & ~n20920;
  assign n20922 = ~n20871 & ~n20884;
  assign n20923 = ~n20856 & ~n20866;
  assign n20924 = ~n408 & ~n703;
  assign n20925 = n514 & n20924;
  assign n20926 = n533 & n1914;
  assign n20927 = n3101 & n3717;
  assign n20928 = n4102 & n20927;
  assign n20929 = n20925 & n20926;
  assign n20930 = n757 & n3725;
  assign n20931 = n20929 & n20930;
  assign n20932 = n20928 & n20931;
  assign n20933 = ~n111 & ~n246;
  assign n20934 = ~n412 & ~n592;
  assign n20935 = ~n597 & n20934;
  assign n20936 = n942 & n20933;
  assign n20937 = n1187 & n1291;
  assign n20938 = n1864 & n20937;
  assign n20939 = n20935 & n20936;
  assign n20940 = n20938 & n20939;
  assign n20941 = n1028 & n4056;
  assign n20942 = n6157 & n20941;
  assign n20943 = n20940 & n20942;
  assign n20944 = n20932 & n20943;
  assign n20945 = n12811 & n20944;
  assign n20946 = n4879 & n20945;
  assign n20947 = ~n12736 & n20946;
  assign n20948 = n12736 & ~n20946;
  assign n20949 = ~n20947 & ~n20948;
  assign n20950 = ~n20923 & n20949;
  assign n20951 = n20923 & ~n20949;
  assign n20952 = ~n20950 & ~n20951;
  assign n20953 = n748 & n12404;
  assign n20954 = n880 & n13128;
  assign n20955 = n3692 & n12401;
  assign n20956 = n3694 & n12398;
  assign n20957 = ~n20953 & ~n20955;
  assign n20958 = ~n20956 & n20957;
  assign n20959 = ~n20954 & n20958;
  assign n20960 = n20952 & n20959;
  assign n20961 = ~n20952 & ~n20959;
  assign n20962 = ~n20960 & ~n20961;
  assign n20963 = n3810 & n12395;
  assign n20964 = n3886 & n13144;
  assign n20965 = n3884 & n12362;
  assign n20966 = n4380 & n12392;
  assign n20967 = ~n20963 & ~n20965;
  assign n20968 = ~n20966 & n20967;
  assign n20969 = ~n20964 & n20968;
  assign n20970 = pi29  & n20969;
  assign n20971 = ~pi29  & ~n20969;
  assign n20972 = ~n20970 & ~n20971;
  assign n20973 = ~n20962 & ~n20972;
  assign n20974 = n20962 & n20972;
  assign n20975 = ~n20973 & ~n20974;
  assign n20976 = ~n20922 & n20975;
  assign n20977 = n20922 & ~n20975;
  assign n20978 = ~n20976 & ~n20977;
  assign n20979 = n86 & n12646;
  assign n20980 = n4420 & n13261;
  assign n20981 = n4600 & n13164;
  assign n20982 = n4615 & n13166;
  assign n20983 = ~n20979 & ~n20981;
  assign n20984 = ~n20982 & n20983;
  assign n20985 = ~n20980 & n20984;
  assign n20986 = pi26  & n20985;
  assign n20987 = ~pi26  & ~n20985;
  assign n20988 = ~n20986 & ~n20987;
  assign n20989 = n20978 & ~n20988;
  assign n20990 = ~n20978 & n20988;
  assign n20991 = ~n20989 & ~n20990;
  assign n20992 = n20921 & n20991;
  assign n20993 = ~n20921 & ~n20991;
  assign n20994 = ~n20992 & ~n20993;
  assign n20995 = n20842 & ~n20895;
  assign n20996 = ~n20896 & ~n20995;
  assign n20997 = n20994 & n20996;
  assign n20998 = ~n20994 & ~n20996;
  assign n20999 = ~n20997 & ~n20998;
  assign n21000 = ~n20901 & ~n20904;
  assign n21001 = n20999 & ~n21000;
  assign n21002 = ~n20999 & n21000;
  assign n21003 = ~n21001 & ~n21002;
  assign n21004 = n20906 & n21003;
  assign n21005 = n20826 & ~n20828;
  assign n21006 = ~n20829 & ~n21005;
  assign n21007 = n20906 & n21006;
  assign n21008 = ~n13795 & n20824;
  assign n21009 = ~n20825 & ~n21008;
  assign n21010 = n21006 & n21009;
  assign n21011 = n13903 & n20822;
  assign n21012 = ~n20823 & ~n21011;
  assign n21013 = n21009 & n21012;
  assign n21014 = n20818 & ~n20820;
  assign n21015 = ~n20821 & ~n21014;
  assign n21016 = n21012 & n21015;
  assign n21017 = ~n14271 & n20816;
  assign n21018 = ~n20817 & ~n21017;
  assign n21019 = n21015 & n21018;
  assign n21020 = n14553 & n20814;
  assign n21021 = ~n20815 & ~n21020;
  assign n21022 = n21018 & n21021;
  assign n21023 = n20810 & ~n20812;
  assign n21024 = ~n20813 & ~n21023;
  assign n21025 = n21021 & n21024;
  assign n21026 = ~n15282 & n20808;
  assign n21027 = ~n20809 & ~n21026;
  assign n21028 = n21024 & n21027;
  assign n21029 = n15445 & n20806;
  assign n21030 = ~n20807 & ~n21029;
  assign n21031 = n21027 & n21030;
  assign n21032 = n20802 & ~n20804;
  assign n21033 = ~n20805 & ~n21032;
  assign n21034 = n21030 & n21033;
  assign n21035 = ~n15957 & n20800;
  assign n21036 = ~n20801 & ~n21035;
  assign n21037 = n21033 & n21036;
  assign n21038 = n16359 & n20798;
  assign n21039 = ~n20799 & ~n21038;
  assign n21040 = n21036 & n21039;
  assign n21041 = n20794 & ~n20796;
  assign n21042 = ~n20797 & ~n21041;
  assign n21043 = n21039 & n21042;
  assign n21044 = ~n17261 & n20792;
  assign n21045 = ~n20793 & ~n21044;
  assign n21046 = n21042 & n21045;
  assign n21047 = n17769 & n20790;
  assign n21048 = ~n20791 & ~n21047;
  assign n21049 = n21045 & n21048;
  assign n21050 = n20786 & ~n20788;
  assign n21051 = ~n20789 & ~n21050;
  assign n21052 = n21048 & n21051;
  assign n21053 = ~n18883 & n20784;
  assign n21054 = ~n20785 & ~n21053;
  assign n21055 = n21051 & n21054;
  assign n21056 = ~n19496 & n20782;
  assign n21057 = ~n20783 & ~n21056;
  assign n21058 = n21054 & n21057;
  assign n21059 = ~n19530 & n20780;
  assign n21060 = ~n20781 & ~n21059;
  assign n21061 = n21057 & n21060;
  assign n21062 = ~n20159 & n20778;
  assign n21063 = ~n20779 & ~n21062;
  assign n21064 = n21060 & n21063;
  assign n21065 = n20774 & ~n20776;
  assign n21066 = ~n20777 & ~n21065;
  assign n21067 = n21063 & n21066;
  assign n21068 = n20770 & ~n20772;
  assign n21069 = ~n20773 & ~n21068;
  assign n21070 = n21066 & n21069;
  assign n21071 = n20766 & ~n20768;
  assign n21072 = ~n20769 & ~n21071;
  assign n21073 = n21069 & n21072;
  assign n21074 = n20762 & ~n20764;
  assign n21075 = ~n20765 & ~n21074;
  assign n21076 = n21072 & n21075;
  assign n21077 = n20758 & ~n20760;
  assign n21078 = ~n20761 & ~n21077;
  assign n21079 = n21075 & n21078;
  assign n21080 = n20754 & ~n20756;
  assign n21081 = ~n20757 & ~n21080;
  assign n21082 = n21078 & n21081;
  assign n21083 = n20750 & ~n20752;
  assign n21084 = ~n20753 & ~n21083;
  assign n21085 = n21081 & n21084;
  assign n21086 = ~n21081 & ~n21084;
  assign n21087 = ~n21085 & ~n21086;
  assign n21088 = n20746 & ~n20748;
  assign n21089 = ~n20749 & ~n21088;
  assign n21090 = n20279 & n20744;
  assign n21091 = ~n20745 & ~n21090;
  assign n21092 = ~n21084 & ~n21091;
  assign n21093 = n21089 & ~n21092;
  assign n21094 = n21087 & n21093;
  assign n21095 = ~n21085 & ~n21094;
  assign n21096 = ~n21078 & ~n21081;
  assign n21097 = ~n21082 & ~n21096;
  assign n21098 = ~n21095 & n21097;
  assign n21099 = ~n21082 & ~n21098;
  assign n21100 = ~n21075 & ~n21078;
  assign n21101 = ~n21079 & ~n21100;
  assign n21102 = ~n21099 & n21101;
  assign n21103 = ~n21079 & ~n21102;
  assign n21104 = ~n21072 & ~n21075;
  assign n21105 = ~n21076 & ~n21104;
  assign n21106 = ~n21103 & n21105;
  assign n21107 = ~n21076 & ~n21106;
  assign n21108 = ~n21069 & ~n21072;
  assign n21109 = ~n21073 & ~n21108;
  assign n21110 = ~n21107 & n21109;
  assign n21111 = ~n21073 & ~n21110;
  assign n21112 = ~n21066 & ~n21069;
  assign n21113 = ~n21070 & ~n21112;
  assign n21114 = ~n21111 & n21113;
  assign n21115 = ~n21070 & ~n21114;
  assign n21116 = ~n21063 & ~n21066;
  assign n21117 = ~n21067 & ~n21116;
  assign n21118 = ~n21115 & n21117;
  assign n21119 = ~n21067 & ~n21118;
  assign n21120 = ~n21060 & ~n21063;
  assign n21121 = ~n21064 & ~n21120;
  assign n21122 = ~n21119 & n21121;
  assign n21123 = ~n21064 & ~n21122;
  assign n21124 = ~n21057 & ~n21060;
  assign n21125 = ~n21061 & ~n21124;
  assign n21126 = ~n21123 & n21125;
  assign n21127 = ~n21061 & ~n21126;
  assign n21128 = ~n21054 & ~n21057;
  assign n21129 = ~n21058 & ~n21128;
  assign n21130 = ~n21127 & n21129;
  assign n21131 = ~n21058 & ~n21130;
  assign n21132 = ~n21051 & ~n21054;
  assign n21133 = ~n21055 & ~n21132;
  assign n21134 = ~n21131 & n21133;
  assign n21135 = ~n21055 & ~n21134;
  assign n21136 = ~n21048 & ~n21051;
  assign n21137 = ~n21052 & ~n21136;
  assign n21138 = ~n21135 & n21137;
  assign n21139 = ~n21052 & ~n21138;
  assign n21140 = ~n21045 & ~n21048;
  assign n21141 = ~n21049 & ~n21140;
  assign n21142 = ~n21139 & n21141;
  assign n21143 = ~n21049 & ~n21142;
  assign n21144 = ~n21042 & ~n21045;
  assign n21145 = ~n21046 & ~n21144;
  assign n21146 = ~n21143 & n21145;
  assign n21147 = ~n21046 & ~n21146;
  assign n21148 = ~n21039 & ~n21042;
  assign n21149 = ~n21043 & ~n21148;
  assign n21150 = ~n21147 & n21149;
  assign n21151 = ~n21043 & ~n21150;
  assign n21152 = ~n21036 & ~n21039;
  assign n21153 = ~n21040 & ~n21152;
  assign n21154 = ~n21151 & n21153;
  assign n21155 = ~n21040 & ~n21154;
  assign n21156 = ~n21033 & ~n21036;
  assign n21157 = ~n21037 & ~n21156;
  assign n21158 = ~n21155 & n21157;
  assign n21159 = ~n21037 & ~n21158;
  assign n21160 = ~n21030 & ~n21033;
  assign n21161 = ~n21034 & ~n21160;
  assign n21162 = ~n21159 & n21161;
  assign n21163 = ~n21034 & ~n21162;
  assign n21164 = ~n21027 & ~n21030;
  assign n21165 = ~n21031 & ~n21164;
  assign n21166 = ~n21163 & n21165;
  assign n21167 = ~n21031 & ~n21166;
  assign n21168 = ~n21024 & ~n21027;
  assign n21169 = ~n21028 & ~n21168;
  assign n21170 = ~n21167 & n21169;
  assign n21171 = ~n21028 & ~n21170;
  assign n21172 = ~n21021 & ~n21024;
  assign n21173 = ~n21025 & ~n21172;
  assign n21174 = ~n21171 & n21173;
  assign n21175 = ~n21025 & ~n21174;
  assign n21176 = ~n21018 & ~n21021;
  assign n21177 = ~n21022 & ~n21176;
  assign n21178 = ~n21175 & n21177;
  assign n21179 = ~n21022 & ~n21178;
  assign n21180 = ~n21015 & ~n21018;
  assign n21181 = ~n21019 & ~n21180;
  assign n21182 = ~n21179 & n21181;
  assign n21183 = ~n21019 & ~n21182;
  assign n21184 = ~n21012 & ~n21015;
  assign n21185 = ~n21016 & ~n21184;
  assign n21186 = ~n21183 & n21185;
  assign n21187 = ~n21016 & ~n21186;
  assign n21188 = ~n21009 & ~n21012;
  assign n21189 = ~n21013 & ~n21188;
  assign n21190 = ~n21187 & n21189;
  assign n21191 = ~n21013 & ~n21190;
  assign n21192 = ~n21006 & ~n21009;
  assign n21193 = ~n21010 & ~n21192;
  assign n21194 = ~n21191 & n21193;
  assign n21195 = ~n21010 & ~n21194;
  assign n21196 = ~n20906 & ~n21006;
  assign n21197 = ~n21007 & ~n21196;
  assign n21198 = ~n21195 & n21197;
  assign n21199 = ~n21007 & ~n21198;
  assign n21200 = ~n20906 & ~n21003;
  assign n21201 = ~n21004 & ~n21200;
  assign n21202 = ~n21199 & n21201;
  assign n21203 = ~n21004 & ~n21202;
  assign n21204 = ~n20997 & ~n21001;
  assign n21205 = n4615 & n13161;
  assign n21206 = n4420 & n13183;
  assign n21207 = n4600 & n13166;
  assign n21208 = n86 & n13164;
  assign n21209 = ~n21207 & ~n21208;
  assign n21210 = ~n21205 & n21209;
  assign n21211 = ~n21206 & n21210;
  assign n21212 = pi26  & n21211;
  assign n21213 = ~pi26  & ~n21211;
  assign n21214 = ~n21212 & ~n21213;
  assign n21215 = ~n20976 & n20988;
  assign n21216 = ~n20977 & ~n21215;
  assign n21217 = n21214 & n21216;
  assign n21218 = ~n21214 & ~n21216;
  assign n21219 = ~n21217 & ~n21218;
  assign n21220 = n20952 & ~n20959;
  assign n21221 = ~n20973 & ~n21220;
  assign n21222 = ~n20947 & ~n20950;
  assign n21223 = n5036 & n5043;
  assign n21224 = ~n12786 & ~n21223;
  assign n21225 = pi23  & ~n21224;
  assign n21226 = ~pi23  & n21224;
  assign n21227 = ~n21225 & ~n21226;
  assign n21228 = ~n111 & ~n235;
  assign n21229 = ~n300 & ~n358;
  assign n21230 = n21228 & n21229;
  assign n21231 = n600 & n1123;
  assign n21232 = n1306 & n1752;
  assign n21233 = n4164 & n6967;
  assign n21234 = n21232 & n21233;
  assign n21235 = n21230 & n21231;
  assign n21236 = n6872 & n21235;
  assign n21237 = n796 & n21234;
  assign n21238 = n21236 & n21237;
  assign n21239 = n5298 & n21238;
  assign n21240 = n13643 & n15089;
  assign n21241 = n21239 & n21240;
  assign n21242 = n12941 & n21241;
  assign n21243 = n20946 & n21242;
  assign n21244 = ~n20946 & ~n21242;
  assign n21245 = ~n21243 & ~n21244;
  assign n21246 = n21227 & n21245;
  assign n21247 = ~n21227 & ~n21245;
  assign n21248 = ~n21246 & ~n21247;
  assign n21249 = ~n21222 & n21248;
  assign n21250 = n21222 & ~n21248;
  assign n21251 = ~n21249 & ~n21250;
  assign n21252 = n748 & n12401;
  assign n21253 = n880 & n13108;
  assign n21254 = n3692 & n12398;
  assign n21255 = n3694 & n12395;
  assign n21256 = ~n21252 & ~n21254;
  assign n21257 = ~n21255 & n21256;
  assign n21258 = ~n21253 & n21257;
  assign n21259 = n21251 & ~n21258;
  assign n21260 = ~n21251 & n21258;
  assign n21261 = ~n21259 & ~n21260;
  assign n21262 = n21221 & ~n21261;
  assign n21263 = ~n21221 & n21261;
  assign n21264 = ~n21262 & ~n21263;
  assign n21265 = n3810 & n12362;
  assign n21266 = n3886 & n12652;
  assign n21267 = n3884 & n12392;
  assign n21268 = n4380 & n12646;
  assign n21269 = ~n21265 & ~n21267;
  assign n21270 = ~n21268 & n21269;
  assign n21271 = ~n21266 & n21270;
  assign n21272 = pi29  & n21271;
  assign n21273 = ~pi29  & ~n21271;
  assign n21274 = ~n21272 & ~n21273;
  assign n21275 = n21264 & ~n21274;
  assign n21276 = ~n21264 & n21274;
  assign n21277 = ~n21275 & ~n21276;
  assign n21278 = ~n21219 & n21277;
  assign n21279 = n21219 & ~n21277;
  assign n21280 = ~n21278 & ~n21279;
  assign n21281 = ~n20919 & ~n20991;
  assign n21282 = ~n20920 & ~n21281;
  assign n21283 = n21280 & n21282;
  assign n21284 = ~n21280 & ~n21282;
  assign n21285 = ~n21283 & ~n21284;
  assign n21286 = ~n21204 & n21285;
  assign n21287 = n21204 & ~n21285;
  assign n21288 = ~n21286 & ~n21287;
  assign n21289 = n21003 & n21288;
  assign n21290 = ~n21003 & ~n21288;
  assign n21291 = ~n21289 & ~n21290;
  assign n21292 = ~n21203 & n21291;
  assign n21293 = n21203 & ~n21291;
  assign n21294 = ~n21292 & ~n21293;
  assign n21295 = n9491 & n21294;
  assign n21296 = n10469 & n21003;
  assign n21297 = n11031 & n21288;
  assign n21298 = ~n20907 & ~n21296;
  assign n21299 = ~n21297 & n21298;
  assign n21300 = ~n21295 & n21299;
  assign n21301 = ~pi5  & ~n21300;
  assign n21302 = pi5  & n21300;
  assign n21303 = ~n21301 & ~n21302;
  assign n21304 = n7430 & n21027;
  assign n21305 = n21171 & ~n21173;
  assign n21306 = ~n21174 & ~n21305;
  assign n21307 = n7431 & n21306;
  assign n21308 = n7869 & n21024;
  assign n21309 = n7895 & n21021;
  assign n21310 = ~n21304 & ~n21308;
  assign n21311 = ~n21309 & n21310;
  assign n21312 = ~n21307 & n21311;
  assign n21313 = ~pi11  & ~n21312;
  assign n21314 = pi11  & n21312;
  assign n21315 = ~n21313 & ~n21314;
  assign n21316 = n5240 & n21060;
  assign n21317 = n21127 & ~n21129;
  assign n21318 = ~n21130 & ~n21317;
  assign n21319 = n5241 & n21318;
  assign n21320 = n5853 & n21057;
  assign n21321 = n5866 & n21054;
  assign n21322 = ~n21316 & ~n21320;
  assign n21323 = ~n21321 & n21322;
  assign n21324 = ~n21319 & n21323;
  assign n21325 = ~pi20  & ~n21324;
  assign n21326 = pi20  & n21324;
  assign n21327 = ~n21325 & ~n21326;
  assign n21328 = n86 & n21081;
  assign n21329 = n21099 & ~n21101;
  assign n21330 = ~n21102 & ~n21329;
  assign n21331 = n4420 & n21330;
  assign n21332 = n4600 & n21078;
  assign n21333 = n4615 & n21075;
  assign n21334 = ~n21328 & ~n21332;
  assign n21335 = ~n21333 & n21334;
  assign n21336 = ~n21331 & n21335;
  assign n21337 = ~pi26  & ~n21336;
  assign n21338 = pi26  & n21336;
  assign n21339 = ~n21337 & ~n21338;
  assign n21340 = ~n3807 & n21091;
  assign n21341 = n3884 & n21091;
  assign n21342 = n4380 & n21089;
  assign n21343 = n21089 & ~n21091;
  assign n21344 = ~n21089 & n21091;
  assign n21345 = ~n21343 & ~n21344;
  assign n21346 = n3886 & ~n21345;
  assign n21347 = ~n21341 & ~n21342;
  assign n21348 = ~n21346 & n21347;
  assign n21349 = pi29  & ~n21340;
  assign n21350 = n21348 & n21349;
  assign n21351 = pi29  & ~n21350;
  assign n21352 = n3810 & n21091;
  assign n21353 = n21084 & ~n21343;
  assign n21354 = ~n21084 & n21343;
  assign n21355 = ~n21353 & ~n21354;
  assign n21356 = n3886 & ~n21355;
  assign n21357 = n3884 & n21089;
  assign n21358 = n4380 & n21084;
  assign n21359 = ~n21352 & ~n21357;
  assign n21360 = ~n21358 & n21359;
  assign n21361 = ~n21356 & n21360;
  assign n21362 = ~n21351 & n21361;
  assign n21363 = n21351 & ~n21361;
  assign n21364 = ~n21362 & ~n21363;
  assign n21365 = ~n21339 & ~n21364;
  assign n21366 = n21339 & n21364;
  assign n21367 = ~n21365 & ~n21366;
  assign n21368 = n86 & n21084;
  assign n21369 = n21095 & ~n21097;
  assign n21370 = ~n21098 & ~n21369;
  assign n21371 = n4420 & n21370;
  assign n21372 = n4600 & n21081;
  assign n21373 = n4615 & n21078;
  assign n21374 = ~n21368 & ~n21372;
  assign n21375 = ~n21373 & n21374;
  assign n21376 = ~n21371 & n21375;
  assign n21377 = pi26  & n21376;
  assign n21378 = ~pi26  & ~n21376;
  assign n21379 = ~n21377 & ~n21378;
  assign n21380 = pi29  & n21340;
  assign n21381 = ~n21348 & n21380;
  assign n21382 = n21348 & ~n21380;
  assign n21383 = ~n21381 & ~n21382;
  assign n21384 = ~n21379 & n21383;
  assign n21385 = ~n81 & n21091;
  assign n21386 = n4600 & n21091;
  assign n21387 = n4615 & n21089;
  assign n21388 = n4420 & ~n21345;
  assign n21389 = ~n21386 & ~n21387;
  assign n21390 = ~n21388 & n21389;
  assign n21391 = pi26  & ~n21385;
  assign n21392 = n21390 & n21391;
  assign n21393 = n86 & n21091;
  assign n21394 = n4420 & ~n21355;
  assign n21395 = n4600 & n21089;
  assign n21396 = n4615 & n21084;
  assign n21397 = ~n21393 & ~n21395;
  assign n21398 = ~n21396 & n21397;
  assign n21399 = ~n21394 & n21398;
  assign n21400 = n21392 & n21399;
  assign n21401 = n21340 & n21400;
  assign n21402 = ~n21340 & n21400;
  assign n21403 = n21340 & ~n21400;
  assign n21404 = ~n21402 & ~n21403;
  assign n21405 = n86 & n21089;
  assign n21406 = ~n21087 & ~n21093;
  assign n21407 = ~n21094 & ~n21406;
  assign n21408 = n4420 & n21407;
  assign n21409 = n4600 & n21084;
  assign n21410 = n4615 & n21081;
  assign n21411 = ~n21405 & ~n21409;
  assign n21412 = ~n21410 & n21411;
  assign n21413 = ~n21408 & n21412;
  assign n21414 = pi26  & n21413;
  assign n21415 = ~pi26  & ~n21413;
  assign n21416 = ~n21414 & ~n21415;
  assign n21417 = ~n21404 & ~n21416;
  assign n21418 = ~n21401 & ~n21417;
  assign n21419 = n21379 & ~n21383;
  assign n21420 = ~n21384 & ~n21419;
  assign n21421 = ~n21418 & n21420;
  assign n21422 = ~n21384 & ~n21421;
  assign n21423 = ~n21367 & ~n21422;
  assign n21424 = n21367 & n21422;
  assign n21425 = ~n21423 & ~n21424;
  assign n21426 = n5044 & n21072;
  assign n21427 = n21111 & ~n21113;
  assign n21428 = ~n21114 & ~n21427;
  assign n21429 = n5045 & n21428;
  assign n21430 = n5109 & n21069;
  assign n21431 = n5130 & n21066;
  assign n21432 = ~n21426 & ~n21430;
  assign n21433 = ~n21431 & n21432;
  assign n21434 = ~n21429 & n21433;
  assign n21435 = pi23  & n21434;
  assign n21436 = ~pi23  & ~n21434;
  assign n21437 = ~n21435 & ~n21436;
  assign n21438 = n21425 & ~n21437;
  assign n21439 = n5044 & n21075;
  assign n21440 = n21107 & ~n21109;
  assign n21441 = ~n21110 & ~n21440;
  assign n21442 = n5045 & n21441;
  assign n21443 = n5109 & n21072;
  assign n21444 = n5130 & n21069;
  assign n21445 = ~n21439 & ~n21443;
  assign n21446 = ~n21444 & n21445;
  assign n21447 = ~n21442 & n21446;
  assign n21448 = ~pi23  & ~n21447;
  assign n21449 = pi23  & n21447;
  assign n21450 = ~n21448 & ~n21449;
  assign n21451 = n21418 & ~n21420;
  assign n21452 = ~n21421 & ~n21451;
  assign n21453 = ~n21450 & n21452;
  assign n21454 = ~n21450 & ~n21452;
  assign n21455 = n21450 & n21452;
  assign n21456 = ~n21454 & ~n21455;
  assign n21457 = n5044 & n21078;
  assign n21458 = n21103 & ~n21105;
  assign n21459 = ~n21106 & ~n21458;
  assign n21460 = n5045 & n21459;
  assign n21461 = n5109 & n21075;
  assign n21462 = n5130 & n21072;
  assign n21463 = ~n21457 & ~n21461;
  assign n21464 = ~n21462 & n21463;
  assign n21465 = ~n21460 & n21464;
  assign n21466 = pi23  & n21465;
  assign n21467 = ~pi23  & ~n21465;
  assign n21468 = ~n21466 & ~n21467;
  assign n21469 = n21404 & n21416;
  assign n21470 = ~n21417 & ~n21469;
  assign n21471 = ~n21468 & n21470;
  assign n21472 = n5044 & n21081;
  assign n21473 = n5045 & n21330;
  assign n21474 = n5109 & n21078;
  assign n21475 = n5130 & n21075;
  assign n21476 = ~n21472 & ~n21474;
  assign n21477 = ~n21475 & n21476;
  assign n21478 = ~n21473 & n21477;
  assign n21479 = ~pi23  & ~n21478;
  assign n21480 = pi23  & n21478;
  assign n21481 = ~n21479 & ~n21480;
  assign n21482 = pi26  & ~n21392;
  assign n21483 = n21399 & ~n21482;
  assign n21484 = ~n21399 & n21482;
  assign n21485 = ~n21483 & ~n21484;
  assign n21486 = ~n21481 & n21485;
  assign n21487 = ~n21481 & ~n21485;
  assign n21488 = n21481 & n21485;
  assign n21489 = ~n21487 & ~n21488;
  assign n21490 = n5044 & n21084;
  assign n21491 = n5045 & n21370;
  assign n21492 = n5109 & n21081;
  assign n21493 = n5130 & n21078;
  assign n21494 = ~n21490 & ~n21492;
  assign n21495 = ~n21493 & n21494;
  assign n21496 = ~n21491 & n21495;
  assign n21497 = pi23  & n21496;
  assign n21498 = ~pi23  & ~n21496;
  assign n21499 = ~n21497 & ~n21498;
  assign n21500 = pi26  & n21385;
  assign n21501 = ~n21390 & n21500;
  assign n21502 = n21390 & ~n21500;
  assign n21503 = ~n21501 & ~n21502;
  assign n21504 = ~n21499 & n21503;
  assign n21505 = ~n5042 & n21091;
  assign n21506 = n5109 & n21091;
  assign n21507 = n5130 & n21089;
  assign n21508 = n5045 & ~n21345;
  assign n21509 = ~n21506 & ~n21507;
  assign n21510 = ~n21508 & n21509;
  assign n21511 = pi23  & ~n21505;
  assign n21512 = n21510 & n21511;
  assign n21513 = n5044 & n21091;
  assign n21514 = n5045 & ~n21355;
  assign n21515 = n5109 & n21089;
  assign n21516 = n5130 & n21084;
  assign n21517 = ~n21513 & ~n21515;
  assign n21518 = ~n21516 & n21517;
  assign n21519 = ~n21514 & n21518;
  assign n21520 = n21512 & n21519;
  assign n21521 = n21385 & n21520;
  assign n21522 = ~n21385 & n21520;
  assign n21523 = n21385 & ~n21520;
  assign n21524 = ~n21522 & ~n21523;
  assign n21525 = n5044 & n21089;
  assign n21526 = n5045 & n21407;
  assign n21527 = n5109 & n21084;
  assign n21528 = n5130 & n21081;
  assign n21529 = ~n21525 & ~n21527;
  assign n21530 = ~n21528 & n21529;
  assign n21531 = ~n21526 & n21530;
  assign n21532 = pi23  & n21531;
  assign n21533 = ~pi23  & ~n21531;
  assign n21534 = ~n21532 & ~n21533;
  assign n21535 = ~n21524 & ~n21534;
  assign n21536 = ~n21521 & ~n21535;
  assign n21537 = n21499 & ~n21503;
  assign n21538 = ~n21504 & ~n21537;
  assign n21539 = ~n21536 & n21538;
  assign n21540 = ~n21504 & ~n21539;
  assign n21541 = ~n21489 & ~n21540;
  assign n21542 = ~n21486 & ~n21541;
  assign n21543 = n21468 & ~n21470;
  assign n21544 = ~n21471 & ~n21543;
  assign n21545 = ~n21542 & n21544;
  assign n21546 = ~n21471 & ~n21545;
  assign n21547 = ~n21456 & ~n21546;
  assign n21548 = ~n21453 & ~n21547;
  assign n21549 = n21425 & n21437;
  assign n21550 = ~n21425 & ~n21437;
  assign n21551 = ~n21549 & ~n21550;
  assign n21552 = ~n21548 & ~n21551;
  assign n21553 = ~n21438 & ~n21552;
  assign n21554 = n86 & n21078;
  assign n21555 = n4420 & n21459;
  assign n21556 = n4600 & n21075;
  assign n21557 = n4615 & n21072;
  assign n21558 = ~n21554 & ~n21556;
  assign n21559 = ~n21557 & n21558;
  assign n21560 = ~n21555 & n21559;
  assign n21561 = ~pi26  & ~n21560;
  assign n21562 = pi26  & n21560;
  assign n21563 = ~n21561 & ~n21562;
  assign n21564 = n3810 & n21089;
  assign n21565 = n3886 & n21407;
  assign n21566 = n3884 & n21084;
  assign n21567 = n4380 & n21081;
  assign n21568 = ~n21564 & ~n21566;
  assign n21569 = ~n21567 & n21568;
  assign n21570 = ~n21565 & n21569;
  assign n21571 = ~pi29  & ~n21570;
  assign n21572 = pi29  & n21570;
  assign n21573 = ~n21571 & ~n21572;
  assign n21574 = n21350 & n21361;
  assign n21575 = ~n746 & n21091;
  assign n21576 = n21574 & ~n21575;
  assign n21577 = ~n21574 & n21575;
  assign n21578 = ~n21576 & ~n21577;
  assign n21579 = ~n21573 & ~n21578;
  assign n21580 = n21573 & n21578;
  assign n21581 = ~n21579 & ~n21580;
  assign n21582 = ~n21563 & ~n21581;
  assign n21583 = n21563 & n21581;
  assign n21584 = ~n21582 & ~n21583;
  assign n21585 = ~n21339 & n21364;
  assign n21586 = ~n21423 & ~n21585;
  assign n21587 = ~n21584 & ~n21586;
  assign n21588 = n21584 & n21586;
  assign n21589 = ~n21587 & ~n21588;
  assign n21590 = n5044 & n21069;
  assign n21591 = n21115 & ~n21117;
  assign n21592 = ~n21118 & ~n21591;
  assign n21593 = n5045 & n21592;
  assign n21594 = n5109 & n21066;
  assign n21595 = n5130 & n21063;
  assign n21596 = ~n21590 & ~n21594;
  assign n21597 = ~n21595 & n21596;
  assign n21598 = ~n21593 & n21597;
  assign n21599 = pi23  & n21598;
  assign n21600 = ~pi23  & ~n21598;
  assign n21601 = ~n21599 & ~n21600;
  assign n21602 = n21589 & ~n21601;
  assign n21603 = ~n21589 & n21601;
  assign n21604 = ~n21602 & ~n21603;
  assign n21605 = ~n21553 & n21604;
  assign n21606 = n21553 & ~n21604;
  assign n21607 = ~n21605 & ~n21606;
  assign n21608 = ~n21327 & ~n21607;
  assign n21609 = n21327 & n21607;
  assign n21610 = ~n21608 & ~n21609;
  assign n21611 = n5240 & n21063;
  assign n21612 = n21123 & ~n21125;
  assign n21613 = ~n21126 & ~n21612;
  assign n21614 = n5241 & n21613;
  assign n21615 = n5853 & n21060;
  assign n21616 = n5866 & n21057;
  assign n21617 = ~n21611 & ~n21615;
  assign n21618 = ~n21616 & n21617;
  assign n21619 = ~n21614 & n21618;
  assign n21620 = ~pi20  & ~n21619;
  assign n21621 = pi20  & n21619;
  assign n21622 = ~n21620 & ~n21621;
  assign n21623 = ~n21548 & n21551;
  assign n21624 = n21548 & ~n21551;
  assign n21625 = ~n21623 & ~n21624;
  assign n21626 = ~n21622 & ~n21625;
  assign n21627 = n21456 & n21546;
  assign n21628 = ~n21547 & ~n21627;
  assign n21629 = n5240 & n21066;
  assign n21630 = n21119 & ~n21121;
  assign n21631 = ~n21122 & ~n21630;
  assign n21632 = n5241 & n21631;
  assign n21633 = n5853 & n21063;
  assign n21634 = n5866 & n21060;
  assign n21635 = ~n21629 & ~n21633;
  assign n21636 = ~n21634 & n21635;
  assign n21637 = ~n21632 & n21636;
  assign n21638 = pi20  & n21637;
  assign n21639 = ~pi20  & ~n21637;
  assign n21640 = ~n21638 & ~n21639;
  assign n21641 = n21628 & ~n21640;
  assign n21642 = n21542 & ~n21544;
  assign n21643 = ~n21545 & ~n21642;
  assign n21644 = n5240 & n21069;
  assign n21645 = n5241 & n21592;
  assign n21646 = n5853 & n21066;
  assign n21647 = n5866 & n21063;
  assign n21648 = ~n21644 & ~n21646;
  assign n21649 = ~n21647 & n21648;
  assign n21650 = ~n21645 & n21649;
  assign n21651 = pi20  & n21650;
  assign n21652 = ~pi20  & ~n21650;
  assign n21653 = ~n21651 & ~n21652;
  assign n21654 = n21643 & ~n21653;
  assign n21655 = n21489 & n21540;
  assign n21656 = ~n21541 & ~n21655;
  assign n21657 = n5240 & n21072;
  assign n21658 = n5241 & n21428;
  assign n21659 = n5853 & n21069;
  assign n21660 = n5866 & n21066;
  assign n21661 = ~n21657 & ~n21659;
  assign n21662 = ~n21660 & n21661;
  assign n21663 = ~n21658 & n21662;
  assign n21664 = pi20  & n21663;
  assign n21665 = ~pi20  & ~n21663;
  assign n21666 = ~n21664 & ~n21665;
  assign n21667 = n21656 & ~n21666;
  assign n21668 = n5240 & n21075;
  assign n21669 = n5241 & n21441;
  assign n21670 = n5853 & n21072;
  assign n21671 = n5866 & n21069;
  assign n21672 = ~n21668 & ~n21670;
  assign n21673 = ~n21671 & n21672;
  assign n21674 = ~n21669 & n21673;
  assign n21675 = ~pi20  & ~n21674;
  assign n21676 = pi20  & n21674;
  assign n21677 = ~n21675 & ~n21676;
  assign n21678 = n21536 & ~n21538;
  assign n21679 = ~n21539 & ~n21678;
  assign n21680 = ~n21677 & n21679;
  assign n21681 = ~n21677 & ~n21679;
  assign n21682 = n21677 & n21679;
  assign n21683 = ~n21681 & ~n21682;
  assign n21684 = n5240 & n21078;
  assign n21685 = n5241 & n21459;
  assign n21686 = n5853 & n21075;
  assign n21687 = n5866 & n21072;
  assign n21688 = ~n21684 & ~n21686;
  assign n21689 = ~n21687 & n21688;
  assign n21690 = ~n21685 & n21689;
  assign n21691 = pi20  & n21690;
  assign n21692 = ~pi20  & ~n21690;
  assign n21693 = ~n21691 & ~n21692;
  assign n21694 = n21524 & n21534;
  assign n21695 = ~n21535 & ~n21694;
  assign n21696 = ~n21693 & n21695;
  assign n21697 = n5240 & n21081;
  assign n21698 = n5241 & n21330;
  assign n21699 = n5853 & n21078;
  assign n21700 = n5866 & n21075;
  assign n21701 = ~n21697 & ~n21699;
  assign n21702 = ~n21700 & n21701;
  assign n21703 = ~n21698 & n21702;
  assign n21704 = ~pi20  & ~n21703;
  assign n21705 = pi20  & n21703;
  assign n21706 = ~n21704 & ~n21705;
  assign n21707 = pi23  & ~n21512;
  assign n21708 = n21519 & ~n21707;
  assign n21709 = ~n21519 & n21707;
  assign n21710 = ~n21708 & ~n21709;
  assign n21711 = ~n21706 & n21710;
  assign n21712 = ~n21706 & ~n21710;
  assign n21713 = n21706 & n21710;
  assign n21714 = ~n21712 & ~n21713;
  assign n21715 = n5240 & n21084;
  assign n21716 = n5241 & n21370;
  assign n21717 = n5853 & n21081;
  assign n21718 = n5866 & n21078;
  assign n21719 = ~n21715 & ~n21717;
  assign n21720 = ~n21718 & n21719;
  assign n21721 = ~n21716 & n21720;
  assign n21722 = pi20  & n21721;
  assign n21723 = ~pi20  & ~n21721;
  assign n21724 = ~n21722 & ~n21723;
  assign n21725 = pi23  & n21505;
  assign n21726 = ~n21510 & n21725;
  assign n21727 = n21510 & ~n21725;
  assign n21728 = ~n21726 & ~n21727;
  assign n21729 = ~n21724 & n21728;
  assign n21730 = ~n5235 & n21091;
  assign n21731 = n5853 & n21091;
  assign n21732 = n5866 & n21089;
  assign n21733 = n5241 & ~n21345;
  assign n21734 = ~n21731 & ~n21732;
  assign n21735 = ~n21733 & n21734;
  assign n21736 = pi20  & ~n21730;
  assign n21737 = n21735 & n21736;
  assign n21738 = n5240 & n21091;
  assign n21739 = n5241 & ~n21355;
  assign n21740 = n5853 & n21089;
  assign n21741 = n5866 & n21084;
  assign n21742 = ~n21738 & ~n21740;
  assign n21743 = ~n21741 & n21742;
  assign n21744 = ~n21739 & n21743;
  assign n21745 = n21737 & n21744;
  assign n21746 = n21505 & n21745;
  assign n21747 = ~n21505 & n21745;
  assign n21748 = n21505 & ~n21745;
  assign n21749 = ~n21747 & ~n21748;
  assign n21750 = n5240 & n21089;
  assign n21751 = n5241 & n21407;
  assign n21752 = n5853 & n21084;
  assign n21753 = n5866 & n21081;
  assign n21754 = ~n21750 & ~n21752;
  assign n21755 = ~n21753 & n21754;
  assign n21756 = ~n21751 & n21755;
  assign n21757 = pi20  & n21756;
  assign n21758 = ~pi20  & ~n21756;
  assign n21759 = ~n21757 & ~n21758;
  assign n21760 = ~n21749 & ~n21759;
  assign n21761 = ~n21746 & ~n21760;
  assign n21762 = n21724 & ~n21728;
  assign n21763 = ~n21729 & ~n21762;
  assign n21764 = ~n21761 & n21763;
  assign n21765 = ~n21729 & ~n21764;
  assign n21766 = ~n21714 & ~n21765;
  assign n21767 = ~n21711 & ~n21766;
  assign n21768 = n21693 & ~n21695;
  assign n21769 = ~n21696 & ~n21768;
  assign n21770 = ~n21767 & n21769;
  assign n21771 = ~n21696 & ~n21770;
  assign n21772 = ~n21683 & ~n21771;
  assign n21773 = ~n21680 & ~n21772;
  assign n21774 = n21656 & n21666;
  assign n21775 = ~n21656 & ~n21666;
  assign n21776 = ~n21774 & ~n21775;
  assign n21777 = ~n21773 & ~n21776;
  assign n21778 = ~n21667 & ~n21777;
  assign n21779 = n21643 & n21653;
  assign n21780 = ~n21643 & ~n21653;
  assign n21781 = ~n21779 & ~n21780;
  assign n21782 = ~n21778 & ~n21781;
  assign n21783 = ~n21654 & ~n21782;
  assign n21784 = ~n21628 & n21640;
  assign n21785 = ~n21641 & ~n21784;
  assign n21786 = ~n21783 & n21785;
  assign n21787 = ~n21641 & ~n21786;
  assign n21788 = n21622 & n21625;
  assign n21789 = ~n21626 & ~n21788;
  assign n21790 = ~n21787 & n21789;
  assign n21791 = ~n21626 & ~n21790;
  assign n21792 = ~n21610 & ~n21791;
  assign n21793 = n21610 & n21791;
  assign n21794 = ~n21792 & ~n21793;
  assign n21795 = n5982 & n21051;
  assign n21796 = n21139 & ~n21141;
  assign n21797 = ~n21142 & ~n21796;
  assign n21798 = n5983 & n21797;
  assign n21799 = n6323 & n21048;
  assign n21800 = n6336 & n21045;
  assign n21801 = ~n21795 & ~n21799;
  assign n21802 = ~n21800 & n21801;
  assign n21803 = ~n21798 & n21802;
  assign n21804 = pi17  & n21803;
  assign n21805 = ~pi17  & ~n21803;
  assign n21806 = ~n21804 & ~n21805;
  assign n21807 = n21794 & ~n21806;
  assign n21808 = n21787 & ~n21789;
  assign n21809 = ~n21790 & ~n21808;
  assign n21810 = n5982 & n21054;
  assign n21811 = n21135 & ~n21137;
  assign n21812 = ~n21138 & ~n21811;
  assign n21813 = n5983 & n21812;
  assign n21814 = n6323 & n21051;
  assign n21815 = n6336 & n21048;
  assign n21816 = ~n21810 & ~n21814;
  assign n21817 = ~n21815 & n21816;
  assign n21818 = ~n21813 & n21817;
  assign n21819 = pi17  & n21818;
  assign n21820 = ~pi17  & ~n21818;
  assign n21821 = ~n21819 & ~n21820;
  assign n21822 = n21809 & ~n21821;
  assign n21823 = n5982 & n21057;
  assign n21824 = n21131 & ~n21133;
  assign n21825 = ~n21134 & ~n21824;
  assign n21826 = n5983 & n21825;
  assign n21827 = n6323 & n21054;
  assign n21828 = n6336 & n21051;
  assign n21829 = ~n21823 & ~n21827;
  assign n21830 = ~n21828 & n21829;
  assign n21831 = ~n21826 & n21830;
  assign n21832 = ~pi17  & ~n21831;
  assign n21833 = pi17  & n21831;
  assign n21834 = ~n21832 & ~n21833;
  assign n21835 = n21783 & ~n21785;
  assign n21836 = ~n21786 & ~n21835;
  assign n21837 = ~n21834 & n21836;
  assign n21838 = ~n21834 & ~n21836;
  assign n21839 = n21834 & n21836;
  assign n21840 = ~n21838 & ~n21839;
  assign n21841 = n5982 & n21060;
  assign n21842 = n5983 & n21318;
  assign n21843 = n6323 & n21057;
  assign n21844 = n6336 & n21054;
  assign n21845 = ~n21841 & ~n21843;
  assign n21846 = ~n21844 & n21845;
  assign n21847 = ~n21842 & n21846;
  assign n21848 = ~pi17  & ~n21847;
  assign n21849 = pi17  & n21847;
  assign n21850 = ~n21848 & ~n21849;
  assign n21851 = n21778 & n21781;
  assign n21852 = ~n21782 & ~n21851;
  assign n21853 = ~n21850 & n21852;
  assign n21854 = ~n21850 & ~n21852;
  assign n21855 = n21850 & n21852;
  assign n21856 = ~n21854 & ~n21855;
  assign n21857 = n5982 & n21063;
  assign n21858 = n5983 & n21613;
  assign n21859 = n6323 & n21060;
  assign n21860 = n6336 & n21057;
  assign n21861 = ~n21857 & ~n21859;
  assign n21862 = ~n21860 & n21861;
  assign n21863 = ~n21858 & n21862;
  assign n21864 = ~pi17  & ~n21863;
  assign n21865 = pi17  & n21863;
  assign n21866 = ~n21864 & ~n21865;
  assign n21867 = ~n21773 & n21776;
  assign n21868 = n21773 & ~n21776;
  assign n21869 = ~n21867 & ~n21868;
  assign n21870 = ~n21866 & ~n21869;
  assign n21871 = n21683 & n21771;
  assign n21872 = ~n21772 & ~n21871;
  assign n21873 = n5982 & n21066;
  assign n21874 = n5983 & n21631;
  assign n21875 = n6323 & n21063;
  assign n21876 = n6336 & n21060;
  assign n21877 = ~n21873 & ~n21875;
  assign n21878 = ~n21876 & n21877;
  assign n21879 = ~n21874 & n21878;
  assign n21880 = pi17  & n21879;
  assign n21881 = ~pi17  & ~n21879;
  assign n21882 = ~n21880 & ~n21881;
  assign n21883 = n21872 & ~n21882;
  assign n21884 = n21767 & ~n21769;
  assign n21885 = ~n21770 & ~n21884;
  assign n21886 = n5982 & n21069;
  assign n21887 = n5983 & n21592;
  assign n21888 = n6323 & n21066;
  assign n21889 = n6336 & n21063;
  assign n21890 = ~n21886 & ~n21888;
  assign n21891 = ~n21889 & n21890;
  assign n21892 = ~n21887 & n21891;
  assign n21893 = pi17  & n21892;
  assign n21894 = ~pi17  & ~n21892;
  assign n21895 = ~n21893 & ~n21894;
  assign n21896 = n21885 & ~n21895;
  assign n21897 = n21714 & n21765;
  assign n21898 = ~n21766 & ~n21897;
  assign n21899 = n5982 & n21072;
  assign n21900 = n5983 & n21428;
  assign n21901 = n6323 & n21069;
  assign n21902 = n6336 & n21066;
  assign n21903 = ~n21899 & ~n21901;
  assign n21904 = ~n21902 & n21903;
  assign n21905 = ~n21900 & n21904;
  assign n21906 = pi17  & n21905;
  assign n21907 = ~pi17  & ~n21905;
  assign n21908 = ~n21906 & ~n21907;
  assign n21909 = n21898 & ~n21908;
  assign n21910 = n5982 & n21075;
  assign n21911 = n5983 & n21441;
  assign n21912 = n6323 & n21072;
  assign n21913 = n6336 & n21069;
  assign n21914 = ~n21910 & ~n21912;
  assign n21915 = ~n21913 & n21914;
  assign n21916 = ~n21911 & n21915;
  assign n21917 = ~pi17  & ~n21916;
  assign n21918 = pi17  & n21916;
  assign n21919 = ~n21917 & ~n21918;
  assign n21920 = n21761 & ~n21763;
  assign n21921 = ~n21764 & ~n21920;
  assign n21922 = ~n21919 & n21921;
  assign n21923 = ~n21919 & ~n21921;
  assign n21924 = n21919 & n21921;
  assign n21925 = ~n21923 & ~n21924;
  assign n21926 = n5982 & n21078;
  assign n21927 = n5983 & n21459;
  assign n21928 = n6323 & n21075;
  assign n21929 = n6336 & n21072;
  assign n21930 = ~n21926 & ~n21928;
  assign n21931 = ~n21929 & n21930;
  assign n21932 = ~n21927 & n21931;
  assign n21933 = pi17  & n21932;
  assign n21934 = ~pi17  & ~n21932;
  assign n21935 = ~n21933 & ~n21934;
  assign n21936 = n21749 & n21759;
  assign n21937 = ~n21760 & ~n21936;
  assign n21938 = ~n21935 & n21937;
  assign n21939 = n5982 & n21081;
  assign n21940 = n5983 & n21330;
  assign n21941 = n6323 & n21078;
  assign n21942 = n6336 & n21075;
  assign n21943 = ~n21939 & ~n21941;
  assign n21944 = ~n21942 & n21943;
  assign n21945 = ~n21940 & n21944;
  assign n21946 = ~pi17  & ~n21945;
  assign n21947 = pi17  & n21945;
  assign n21948 = ~n21946 & ~n21947;
  assign n21949 = pi20  & ~n21737;
  assign n21950 = n21744 & ~n21949;
  assign n21951 = ~n21744 & n21949;
  assign n21952 = ~n21950 & ~n21951;
  assign n21953 = ~n21948 & n21952;
  assign n21954 = ~n21948 & ~n21952;
  assign n21955 = n21948 & n21952;
  assign n21956 = ~n21954 & ~n21955;
  assign n21957 = n5982 & n21084;
  assign n21958 = n5983 & n21370;
  assign n21959 = n6323 & n21081;
  assign n21960 = n6336 & n21078;
  assign n21961 = ~n21957 & ~n21959;
  assign n21962 = ~n21960 & n21961;
  assign n21963 = ~n21958 & n21962;
  assign n21964 = pi17  & n21963;
  assign n21965 = ~pi17  & ~n21963;
  assign n21966 = ~n21964 & ~n21965;
  assign n21967 = pi20  & n21730;
  assign n21968 = ~n21735 & n21967;
  assign n21969 = n21735 & ~n21967;
  assign n21970 = ~n21968 & ~n21969;
  assign n21971 = ~n21966 & n21970;
  assign n21972 = ~n5980 & n21091;
  assign n21973 = n6323 & n21091;
  assign n21974 = n6336 & n21089;
  assign n21975 = n5983 & ~n21345;
  assign n21976 = ~n21973 & ~n21974;
  assign n21977 = ~n21975 & n21976;
  assign n21978 = pi17  & ~n21972;
  assign n21979 = n21977 & n21978;
  assign n21980 = n5982 & n21091;
  assign n21981 = n5983 & ~n21355;
  assign n21982 = n6323 & n21089;
  assign n21983 = n6336 & n21084;
  assign n21984 = ~n21980 & ~n21982;
  assign n21985 = ~n21983 & n21984;
  assign n21986 = ~n21981 & n21985;
  assign n21987 = n21979 & n21986;
  assign n21988 = n21730 & n21987;
  assign n21989 = ~n21730 & n21987;
  assign n21990 = n21730 & ~n21987;
  assign n21991 = ~n21989 & ~n21990;
  assign n21992 = n5982 & n21089;
  assign n21993 = n5983 & n21407;
  assign n21994 = n6323 & n21084;
  assign n21995 = n6336 & n21081;
  assign n21996 = ~n21992 & ~n21994;
  assign n21997 = ~n21995 & n21996;
  assign n21998 = ~n21993 & n21997;
  assign n21999 = pi17  & n21998;
  assign n22000 = ~pi17  & ~n21998;
  assign n22001 = ~n21999 & ~n22000;
  assign n22002 = ~n21991 & ~n22001;
  assign n22003 = ~n21988 & ~n22002;
  assign n22004 = n21966 & ~n21970;
  assign n22005 = ~n21971 & ~n22004;
  assign n22006 = ~n22003 & n22005;
  assign n22007 = ~n21971 & ~n22006;
  assign n22008 = ~n21956 & ~n22007;
  assign n22009 = ~n21953 & ~n22008;
  assign n22010 = n21935 & ~n21937;
  assign n22011 = ~n21938 & ~n22010;
  assign n22012 = ~n22009 & n22011;
  assign n22013 = ~n21938 & ~n22012;
  assign n22014 = ~n21925 & ~n22013;
  assign n22015 = ~n21922 & ~n22014;
  assign n22016 = n21898 & n21908;
  assign n22017 = ~n21898 & ~n21908;
  assign n22018 = ~n22016 & ~n22017;
  assign n22019 = ~n22015 & ~n22018;
  assign n22020 = ~n21909 & ~n22019;
  assign n22021 = n21885 & n21895;
  assign n22022 = ~n21885 & ~n21895;
  assign n22023 = ~n22021 & ~n22022;
  assign n22024 = ~n22020 & ~n22023;
  assign n22025 = ~n21896 & ~n22024;
  assign n22026 = ~n21872 & n21882;
  assign n22027 = ~n21883 & ~n22026;
  assign n22028 = ~n22025 & n22027;
  assign n22029 = ~n21883 & ~n22028;
  assign n22030 = n21866 & n21869;
  assign n22031 = ~n21870 & ~n22030;
  assign n22032 = ~n22029 & n22031;
  assign n22033 = ~n21870 & ~n22032;
  assign n22034 = ~n21856 & ~n22033;
  assign n22035 = ~n21853 & ~n22034;
  assign n22036 = ~n21840 & ~n22035;
  assign n22037 = ~n21837 & ~n22036;
  assign n22038 = n21809 & n21821;
  assign n22039 = ~n21809 & ~n21821;
  assign n22040 = ~n22038 & ~n22039;
  assign n22041 = ~n22037 & ~n22040;
  assign n22042 = ~n21822 & ~n22041;
  assign n22043 = ~n21794 & n21806;
  assign n22044 = ~n21807 & ~n22043;
  assign n22045 = ~n22042 & n22044;
  assign n22046 = ~n21807 & ~n22045;
  assign n22047 = n5982 & n21048;
  assign n22048 = n21143 & ~n21145;
  assign n22049 = ~n21146 & ~n22048;
  assign n22050 = n5983 & n22049;
  assign n22051 = n6323 & n21045;
  assign n22052 = n6336 & n21042;
  assign n22053 = ~n22047 & ~n22051;
  assign n22054 = ~n22052 & n22053;
  assign n22055 = ~n22050 & n22054;
  assign n22056 = ~pi17  & ~n22055;
  assign n22057 = pi17  & n22055;
  assign n22058 = ~n22056 & ~n22057;
  assign n22059 = ~n21327 & n21607;
  assign n22060 = ~n21792 & ~n22059;
  assign n22061 = n5044 & n21066;
  assign n22062 = n5045 & n21631;
  assign n22063 = n5109 & n21063;
  assign n22064 = n5130 & n21060;
  assign n22065 = ~n22061 & ~n22063;
  assign n22066 = ~n22064 & n22065;
  assign n22067 = ~n22062 & n22066;
  assign n22068 = ~pi23  & ~n22067;
  assign n22069 = pi23  & n22067;
  assign n22070 = ~n22068 & ~n22069;
  assign n22071 = ~n21563 & n21581;
  assign n22072 = ~n21587 & ~n22071;
  assign n22073 = n86 & n21075;
  assign n22074 = n4420 & n21441;
  assign n22075 = n4600 & n21072;
  assign n22076 = n4615 & n21069;
  assign n22077 = ~n22073 & ~n22075;
  assign n22078 = ~n22076 & n22077;
  assign n22079 = ~n22074 & n22078;
  assign n22080 = pi26  & n22079;
  assign n22081 = ~pi26  & ~n22079;
  assign n22082 = ~n22080 & ~n22081;
  assign n22083 = n21574 & n21575;
  assign n22084 = ~n21579 & ~n22083;
  assign n22085 = n3810 & n21084;
  assign n22086 = n3886 & n21370;
  assign n22087 = n3884 & n21081;
  assign n22088 = n4380 & n21078;
  assign n22089 = ~n22085 & ~n22087;
  assign n22090 = ~n22088 & n22089;
  assign n22091 = ~n22086 & n22090;
  assign n22092 = ~pi29  & ~n22091;
  assign n22093 = pi29  & n22091;
  assign n22094 = ~n22092 & ~n22093;
  assign n22095 = ~n143 & ~n258;
  assign n22096 = ~n278 & ~n414;
  assign n22097 = ~n416 & n22096;
  assign n22098 = n635 & n22095;
  assign n22099 = n797 & n1230;
  assign n22100 = n1247 & n1358;
  assign n22101 = n1470 & n22100;
  assign n22102 = n22098 & n22099;
  assign n22103 = n22097 & n22102;
  assign n22104 = n22101 & n22103;
  assign n22105 = ~n284 & ~n371;
  assign n22106 = ~n520 & ~n1699;
  assign n22107 = n22105 & n22106;
  assign n22108 = n440 & n479;
  assign n22109 = n752 & n1429;
  assign n22110 = n3016 & n3407;
  assign n22111 = n3837 & n4063;
  assign n22112 = n22110 & n22111;
  assign n22113 = n22108 & n22109;
  assign n22114 = n3836 & n22107;
  assign n22115 = n4689 & n22114;
  assign n22116 = n22112 & n22113;
  assign n22117 = n13323 & n22116;
  assign n22118 = n22115 & n22117;
  assign n22119 = ~n297 & ~n332;
  assign n22120 = ~n338 & ~n568;
  assign n22121 = ~n687 & n22120;
  assign n22122 = n448 & n22119;
  assign n22123 = n1306 & n1403;
  assign n22124 = n1476 & n2037;
  assign n22125 = n22123 & n22124;
  assign n22126 = n22121 & n22122;
  assign n22127 = n2850 & n7017;
  assign n22128 = n22126 & n22127;
  assign n22129 = n1957 & n22125;
  assign n22130 = n14967 & n22129;
  assign n22131 = n22128 & n22130;
  assign n22132 = n22104 & n22131;
  assign n22133 = n14889 & n22118;
  assign n22134 = n22132 & n22133;
  assign n22135 = n3694 & n21089;
  assign n22136 = n3692 & n21091;
  assign n22137 = n880 & ~n21345;
  assign n22138 = ~n22135 & ~n22136;
  assign n22139 = ~n22137 & n22138;
  assign n22140 = ~n22134 & n22139;
  assign n22141 = n22134 & ~n22139;
  assign n22142 = ~n22140 & ~n22141;
  assign n22143 = ~n22094 & ~n22142;
  assign n22144 = n22094 & n22142;
  assign n22145 = ~n22143 & ~n22144;
  assign n22146 = ~n22084 & n22145;
  assign n22147 = n22084 & ~n22145;
  assign n22148 = ~n22146 & ~n22147;
  assign n22149 = n22082 & n22148;
  assign n22150 = ~n22082 & ~n22148;
  assign n22151 = ~n22149 & ~n22150;
  assign n22152 = ~n22072 & ~n22151;
  assign n22153 = n22072 & n22151;
  assign n22154 = ~n22152 & ~n22153;
  assign n22155 = ~n22070 & ~n22154;
  assign n22156 = n22070 & n22154;
  assign n22157 = ~n22155 & ~n22156;
  assign n22158 = ~n21602 & ~n21605;
  assign n22159 = n22157 & n22158;
  assign n22160 = ~n22157 & ~n22158;
  assign n22161 = ~n22159 & ~n22160;
  assign n22162 = n5240 & n21057;
  assign n22163 = n5241 & n21825;
  assign n22164 = n5853 & n21054;
  assign n22165 = n5866 & n21051;
  assign n22166 = ~n22162 & ~n22164;
  assign n22167 = ~n22165 & n22166;
  assign n22168 = ~n22163 & n22167;
  assign n22169 = pi20  & n22168;
  assign n22170 = ~pi20  & ~n22168;
  assign n22171 = ~n22169 & ~n22170;
  assign n22172 = n22161 & n22171;
  assign n22173 = ~n22161 & ~n22171;
  assign n22174 = ~n22172 & ~n22173;
  assign n22175 = ~n22060 & n22174;
  assign n22176 = n22060 & ~n22174;
  assign n22177 = ~n22175 & ~n22176;
  assign n22178 = ~n22058 & ~n22177;
  assign n22179 = n22058 & n22177;
  assign n22180 = ~n22178 & ~n22179;
  assign n22181 = ~n22046 & n22180;
  assign n22182 = n22046 & ~n22180;
  assign n22183 = ~n22181 & ~n22182;
  assign n22184 = n6630 & n21039;
  assign n22185 = n21155 & ~n21157;
  assign n22186 = ~n21158 & ~n22185;
  assign n22187 = n6631 & n22186;
  assign n22188 = n7238 & n21036;
  assign n22189 = n7262 & n21033;
  assign n22190 = ~n22184 & ~n22188;
  assign n22191 = ~n22189 & n22190;
  assign n22192 = ~n22187 & n22191;
  assign n22193 = pi14  & n22192;
  assign n22194 = ~pi14  & ~n22192;
  assign n22195 = ~n22193 & ~n22194;
  assign n22196 = n22183 & ~n22195;
  assign n22197 = n6630 & n21042;
  assign n22198 = n21151 & ~n21153;
  assign n22199 = ~n21154 & ~n22198;
  assign n22200 = n6631 & n22199;
  assign n22201 = n7238 & n21039;
  assign n22202 = n7262 & n21036;
  assign n22203 = ~n22197 & ~n22201;
  assign n22204 = ~n22202 & n22203;
  assign n22205 = ~n22200 & n22204;
  assign n22206 = ~pi14  & ~n22205;
  assign n22207 = pi14  & n22205;
  assign n22208 = ~n22206 & ~n22207;
  assign n22209 = n22042 & ~n22044;
  assign n22210 = ~n22045 & ~n22209;
  assign n22211 = ~n22208 & n22210;
  assign n22212 = ~n22208 & ~n22210;
  assign n22213 = n22208 & n22210;
  assign n22214 = ~n22212 & ~n22213;
  assign n22215 = n6630 & n21045;
  assign n22216 = n21147 & ~n21149;
  assign n22217 = ~n21150 & ~n22216;
  assign n22218 = n6631 & n22217;
  assign n22219 = n7238 & n21042;
  assign n22220 = n7262 & n21039;
  assign n22221 = ~n22215 & ~n22219;
  assign n22222 = ~n22220 & n22221;
  assign n22223 = ~n22218 & n22222;
  assign n22224 = ~pi14  & ~n22223;
  assign n22225 = pi14  & n22223;
  assign n22226 = ~n22224 & ~n22225;
  assign n22227 = n22037 & n22040;
  assign n22228 = ~n22041 & ~n22227;
  assign n22229 = ~n22226 & n22228;
  assign n22230 = ~n22226 & ~n22228;
  assign n22231 = n22226 & n22228;
  assign n22232 = ~n22230 & ~n22231;
  assign n22233 = n21840 & n22035;
  assign n22234 = ~n22036 & ~n22233;
  assign n22235 = n6630 & n21048;
  assign n22236 = n6631 & n22049;
  assign n22237 = n7238 & n21045;
  assign n22238 = n7262 & n21042;
  assign n22239 = ~n22235 & ~n22237;
  assign n22240 = ~n22238 & n22239;
  assign n22241 = ~n22236 & n22240;
  assign n22242 = pi14  & n22241;
  assign n22243 = ~pi14  & ~n22241;
  assign n22244 = ~n22242 & ~n22243;
  assign n22245 = n22234 & ~n22244;
  assign n22246 = n21856 & n22033;
  assign n22247 = ~n22034 & ~n22246;
  assign n22248 = n6630 & n21051;
  assign n22249 = n6631 & n21797;
  assign n22250 = n7238 & n21048;
  assign n22251 = n7262 & n21045;
  assign n22252 = ~n22248 & ~n22250;
  assign n22253 = ~n22251 & n22252;
  assign n22254 = ~n22249 & n22253;
  assign n22255 = pi14  & n22254;
  assign n22256 = ~pi14  & ~n22254;
  assign n22257 = ~n22255 & ~n22256;
  assign n22258 = n22247 & ~n22257;
  assign n22259 = n22029 & ~n22031;
  assign n22260 = ~n22032 & ~n22259;
  assign n22261 = n6630 & n21054;
  assign n22262 = n6631 & n21812;
  assign n22263 = n7238 & n21051;
  assign n22264 = n7262 & n21048;
  assign n22265 = ~n22261 & ~n22263;
  assign n22266 = ~n22264 & n22265;
  assign n22267 = ~n22262 & n22266;
  assign n22268 = pi14  & n22267;
  assign n22269 = ~pi14  & ~n22267;
  assign n22270 = ~n22268 & ~n22269;
  assign n22271 = n22260 & ~n22270;
  assign n22272 = n6630 & n21057;
  assign n22273 = n6631 & n21825;
  assign n22274 = n7238 & n21054;
  assign n22275 = n7262 & n21051;
  assign n22276 = ~n22272 & ~n22274;
  assign n22277 = ~n22275 & n22276;
  assign n22278 = ~n22273 & n22277;
  assign n22279 = ~pi14  & ~n22278;
  assign n22280 = pi14  & n22278;
  assign n22281 = ~n22279 & ~n22280;
  assign n22282 = n22025 & ~n22027;
  assign n22283 = ~n22028 & ~n22282;
  assign n22284 = ~n22281 & n22283;
  assign n22285 = ~n22281 & ~n22283;
  assign n22286 = n22281 & n22283;
  assign n22287 = ~n22285 & ~n22286;
  assign n22288 = n6630 & n21060;
  assign n22289 = n6631 & n21318;
  assign n22290 = n7238 & n21057;
  assign n22291 = n7262 & n21054;
  assign n22292 = ~n22288 & ~n22290;
  assign n22293 = ~n22291 & n22292;
  assign n22294 = ~n22289 & n22293;
  assign n22295 = ~pi14  & ~n22294;
  assign n22296 = pi14  & n22294;
  assign n22297 = ~n22295 & ~n22296;
  assign n22298 = n22020 & n22023;
  assign n22299 = ~n22024 & ~n22298;
  assign n22300 = ~n22297 & n22299;
  assign n22301 = ~n22297 & ~n22299;
  assign n22302 = n22297 & n22299;
  assign n22303 = ~n22301 & ~n22302;
  assign n22304 = n6630 & n21063;
  assign n22305 = n6631 & n21613;
  assign n22306 = n7238 & n21060;
  assign n22307 = n7262 & n21057;
  assign n22308 = ~n22304 & ~n22306;
  assign n22309 = ~n22307 & n22308;
  assign n22310 = ~n22305 & n22309;
  assign n22311 = ~pi14  & ~n22310;
  assign n22312 = pi14  & n22310;
  assign n22313 = ~n22311 & ~n22312;
  assign n22314 = ~n22015 & n22018;
  assign n22315 = n22015 & ~n22018;
  assign n22316 = ~n22314 & ~n22315;
  assign n22317 = ~n22313 & ~n22316;
  assign n22318 = n21925 & n22013;
  assign n22319 = ~n22014 & ~n22318;
  assign n22320 = n6630 & n21066;
  assign n22321 = n6631 & n21631;
  assign n22322 = n7238 & n21063;
  assign n22323 = n7262 & n21060;
  assign n22324 = ~n22320 & ~n22322;
  assign n22325 = ~n22323 & n22324;
  assign n22326 = ~n22321 & n22325;
  assign n22327 = pi14  & n22326;
  assign n22328 = ~pi14  & ~n22326;
  assign n22329 = ~n22327 & ~n22328;
  assign n22330 = n22319 & ~n22329;
  assign n22331 = n22009 & ~n22011;
  assign n22332 = ~n22012 & ~n22331;
  assign n22333 = n6630 & n21069;
  assign n22334 = n6631 & n21592;
  assign n22335 = n7238 & n21066;
  assign n22336 = n7262 & n21063;
  assign n22337 = ~n22333 & ~n22335;
  assign n22338 = ~n22336 & n22337;
  assign n22339 = ~n22334 & n22338;
  assign n22340 = pi14  & n22339;
  assign n22341 = ~pi14  & ~n22339;
  assign n22342 = ~n22340 & ~n22341;
  assign n22343 = n22332 & ~n22342;
  assign n22344 = n21956 & n22007;
  assign n22345 = ~n22008 & ~n22344;
  assign n22346 = n6630 & n21072;
  assign n22347 = n6631 & n21428;
  assign n22348 = n7238 & n21069;
  assign n22349 = n7262 & n21066;
  assign n22350 = ~n22346 & ~n22348;
  assign n22351 = ~n22349 & n22350;
  assign n22352 = ~n22347 & n22351;
  assign n22353 = pi14  & n22352;
  assign n22354 = ~pi14  & ~n22352;
  assign n22355 = ~n22353 & ~n22354;
  assign n22356 = n22345 & ~n22355;
  assign n22357 = n6630 & n21075;
  assign n22358 = n6631 & n21441;
  assign n22359 = n7238 & n21072;
  assign n22360 = n7262 & n21069;
  assign n22361 = ~n22357 & ~n22359;
  assign n22362 = ~n22360 & n22361;
  assign n22363 = ~n22358 & n22362;
  assign n22364 = ~pi14  & ~n22363;
  assign n22365 = pi14  & n22363;
  assign n22366 = ~n22364 & ~n22365;
  assign n22367 = n22003 & ~n22005;
  assign n22368 = ~n22006 & ~n22367;
  assign n22369 = ~n22366 & n22368;
  assign n22370 = ~n22366 & ~n22368;
  assign n22371 = n22366 & n22368;
  assign n22372 = ~n22370 & ~n22371;
  assign n22373 = n6630 & n21078;
  assign n22374 = n6631 & n21459;
  assign n22375 = n7238 & n21075;
  assign n22376 = n7262 & n21072;
  assign n22377 = ~n22373 & ~n22375;
  assign n22378 = ~n22376 & n22377;
  assign n22379 = ~n22374 & n22378;
  assign n22380 = pi14  & n22379;
  assign n22381 = ~pi14  & ~n22379;
  assign n22382 = ~n22380 & ~n22381;
  assign n22383 = n21991 & n22001;
  assign n22384 = ~n22002 & ~n22383;
  assign n22385 = ~n22382 & n22384;
  assign n22386 = n6630 & n21081;
  assign n22387 = n6631 & n21330;
  assign n22388 = n7238 & n21078;
  assign n22389 = n7262 & n21075;
  assign n22390 = ~n22386 & ~n22388;
  assign n22391 = ~n22389 & n22390;
  assign n22392 = ~n22387 & n22391;
  assign n22393 = ~pi14  & ~n22392;
  assign n22394 = pi14  & n22392;
  assign n22395 = ~n22393 & ~n22394;
  assign n22396 = pi17  & ~n21979;
  assign n22397 = n21986 & ~n22396;
  assign n22398 = ~n21986 & n22396;
  assign n22399 = ~n22397 & ~n22398;
  assign n22400 = ~n22395 & n22399;
  assign n22401 = ~n22395 & ~n22399;
  assign n22402 = n22395 & n22399;
  assign n22403 = ~n22401 & ~n22402;
  assign n22404 = n6630 & n21084;
  assign n22405 = n6631 & n21370;
  assign n22406 = n7238 & n21081;
  assign n22407 = n7262 & n21078;
  assign n22408 = ~n22404 & ~n22406;
  assign n22409 = ~n22407 & n22408;
  assign n22410 = ~n22405 & n22409;
  assign n22411 = pi14  & n22410;
  assign n22412 = ~pi14  & ~n22410;
  assign n22413 = ~n22411 & ~n22412;
  assign n22414 = pi17  & n21972;
  assign n22415 = ~n21977 & n22414;
  assign n22416 = n21977 & ~n22414;
  assign n22417 = ~n22415 & ~n22416;
  assign n22418 = ~n22413 & n22417;
  assign n22419 = ~n6628 & n21091;
  assign n22420 = n7238 & n21091;
  assign n22421 = n7262 & n21089;
  assign n22422 = n6631 & ~n21345;
  assign n22423 = ~n22420 & ~n22421;
  assign n22424 = ~n22422 & n22423;
  assign n22425 = pi14  & ~n22419;
  assign n22426 = n22424 & n22425;
  assign n22427 = n6630 & n21091;
  assign n22428 = n6631 & ~n21355;
  assign n22429 = n7238 & n21089;
  assign n22430 = n7262 & n21084;
  assign n22431 = ~n22427 & ~n22429;
  assign n22432 = ~n22430 & n22431;
  assign n22433 = ~n22428 & n22432;
  assign n22434 = n22426 & n22433;
  assign n22435 = n21972 & n22434;
  assign n22436 = ~n21972 & n22434;
  assign n22437 = n21972 & ~n22434;
  assign n22438 = ~n22436 & ~n22437;
  assign n22439 = n6630 & n21089;
  assign n22440 = n6631 & n21407;
  assign n22441 = n7238 & n21084;
  assign n22442 = n7262 & n21081;
  assign n22443 = ~n22439 & ~n22441;
  assign n22444 = ~n22442 & n22443;
  assign n22445 = ~n22440 & n22444;
  assign n22446 = pi14  & n22445;
  assign n22447 = ~pi14  & ~n22445;
  assign n22448 = ~n22446 & ~n22447;
  assign n22449 = ~n22438 & ~n22448;
  assign n22450 = ~n22435 & ~n22449;
  assign n22451 = n22413 & ~n22417;
  assign n22452 = ~n22418 & ~n22451;
  assign n22453 = ~n22450 & n22452;
  assign n22454 = ~n22418 & ~n22453;
  assign n22455 = ~n22403 & ~n22454;
  assign n22456 = ~n22400 & ~n22455;
  assign n22457 = n22382 & ~n22384;
  assign n22458 = ~n22385 & ~n22457;
  assign n22459 = ~n22456 & n22458;
  assign n22460 = ~n22385 & ~n22459;
  assign n22461 = ~n22372 & ~n22460;
  assign n22462 = ~n22369 & ~n22461;
  assign n22463 = n22345 & n22355;
  assign n22464 = ~n22345 & ~n22355;
  assign n22465 = ~n22463 & ~n22464;
  assign n22466 = ~n22462 & ~n22465;
  assign n22467 = ~n22356 & ~n22466;
  assign n22468 = n22332 & n22342;
  assign n22469 = ~n22332 & ~n22342;
  assign n22470 = ~n22468 & ~n22469;
  assign n22471 = ~n22467 & ~n22470;
  assign n22472 = ~n22343 & ~n22471;
  assign n22473 = ~n22319 & n22329;
  assign n22474 = ~n22330 & ~n22473;
  assign n22475 = ~n22472 & n22474;
  assign n22476 = ~n22330 & ~n22475;
  assign n22477 = n22313 & n22316;
  assign n22478 = ~n22317 & ~n22477;
  assign n22479 = ~n22476 & n22478;
  assign n22480 = ~n22317 & ~n22479;
  assign n22481 = ~n22303 & ~n22480;
  assign n22482 = ~n22300 & ~n22481;
  assign n22483 = ~n22287 & ~n22482;
  assign n22484 = ~n22284 & ~n22483;
  assign n22485 = n22260 & n22270;
  assign n22486 = ~n22260 & ~n22270;
  assign n22487 = ~n22485 & ~n22486;
  assign n22488 = ~n22484 & ~n22487;
  assign n22489 = ~n22271 & ~n22488;
  assign n22490 = n22247 & n22257;
  assign n22491 = ~n22247 & ~n22257;
  assign n22492 = ~n22490 & ~n22491;
  assign n22493 = ~n22489 & ~n22492;
  assign n22494 = ~n22258 & ~n22493;
  assign n22495 = ~n22234 & n22244;
  assign n22496 = ~n22245 & ~n22495;
  assign n22497 = ~n22494 & n22496;
  assign n22498 = ~n22245 & ~n22497;
  assign n22499 = ~n22232 & ~n22498;
  assign n22500 = ~n22229 & ~n22499;
  assign n22501 = ~n22214 & ~n22500;
  assign n22502 = ~n22211 & ~n22501;
  assign n22503 = n22183 & n22195;
  assign n22504 = ~n22183 & ~n22195;
  assign n22505 = ~n22503 & ~n22504;
  assign n22506 = ~n22502 & ~n22505;
  assign n22507 = ~n22196 & ~n22506;
  assign n22508 = ~n22178 & ~n22181;
  assign n22509 = n5982 & n21045;
  assign n22510 = n5983 & n22217;
  assign n22511 = n6323 & n21042;
  assign n22512 = n6336 & n21039;
  assign n22513 = ~n22509 & ~n22511;
  assign n22514 = ~n22512 & n22513;
  assign n22515 = ~n22510 & n22514;
  assign n22516 = ~pi17  & ~n22515;
  assign n22517 = pi17  & n22515;
  assign n22518 = ~n22516 & ~n22517;
  assign n22519 = n22161 & ~n22171;
  assign n22520 = ~n22060 & ~n22174;
  assign n22521 = ~n22519 & ~n22520;
  assign n22522 = n5044 & n21063;
  assign n22523 = n5045 & n21613;
  assign n22524 = n5109 & n21060;
  assign n22525 = n5130 & n21057;
  assign n22526 = ~n22522 & ~n22524;
  assign n22527 = ~n22525 & n22526;
  assign n22528 = ~n22523 & n22527;
  assign n22529 = ~pi23  & ~n22528;
  assign n22530 = pi23  & n22528;
  assign n22531 = ~n22529 & ~n22530;
  assign n22532 = ~n22082 & n22148;
  assign n22533 = ~n22152 & ~n22532;
  assign n22534 = ~n22143 & ~n22146;
  assign n22535 = n3810 & n21081;
  assign n22536 = n3886 & n21330;
  assign n22537 = n3884 & n21078;
  assign n22538 = n4380 & n21075;
  assign n22539 = ~n22535 & ~n22537;
  assign n22540 = ~n22538 & n22539;
  assign n22541 = ~n22536 & n22540;
  assign n22542 = ~pi29  & ~n22541;
  assign n22543 = pi29  & n22541;
  assign n22544 = ~n22542 & ~n22543;
  assign n22545 = ~n22134 & ~n22139;
  assign n22546 = ~n256 & ~n317;
  assign n22547 = ~n603 & n22546;
  assign n22548 = ~n278 & ~n432;
  assign n22549 = ~n486 & ~n792;
  assign n22550 = n22548 & n22549;
  assign n22551 = n160 & n935;
  assign n22552 = n958 & n1489;
  assign n22553 = n1779 & n4934;
  assign n22554 = n12930 & n22553;
  assign n22555 = n22551 & n22552;
  assign n22556 = n22547 & n22550;
  assign n22557 = n22555 & n22556;
  assign n22558 = n1953 & n22554;
  assign n22559 = n4053 & n4473;
  assign n22560 = n22558 & n22559;
  assign n22561 = n5658 & n22557;
  assign n22562 = n22560 & n22561;
  assign n22563 = n6941 & n22562;
  assign n22564 = n14889 & n22563;
  assign n22565 = n22545 & ~n22564;
  assign n22566 = ~n22545 & n22564;
  assign n22567 = ~n22565 & ~n22566;
  assign n22568 = n748 & n21091;
  assign n22569 = n880 & ~n21355;
  assign n22570 = n3692 & n21089;
  assign n22571 = n3694 & n21084;
  assign n22572 = ~n22568 & ~n22570;
  assign n22573 = ~n22571 & n22572;
  assign n22574 = ~n22569 & n22573;
  assign n22575 = n22567 & ~n22574;
  assign n22576 = ~n22567 & n22574;
  assign n22577 = ~n22575 & ~n22576;
  assign n22578 = ~n22544 & n22577;
  assign n22579 = n22544 & ~n22577;
  assign n22580 = ~n22578 & ~n22579;
  assign n22581 = n22534 & ~n22580;
  assign n22582 = ~n22534 & n22580;
  assign n22583 = ~n22581 & ~n22582;
  assign n22584 = n86 & n21072;
  assign n22585 = n4420 & n21428;
  assign n22586 = n4600 & n21069;
  assign n22587 = n4615 & n21066;
  assign n22588 = ~n22584 & ~n22586;
  assign n22589 = ~n22587 & n22588;
  assign n22590 = ~n22585 & n22589;
  assign n22591 = pi26  & n22590;
  assign n22592 = ~pi26  & ~n22590;
  assign n22593 = ~n22591 & ~n22592;
  assign n22594 = n22583 & n22593;
  assign n22595 = ~n22583 & ~n22593;
  assign n22596 = ~n22594 & ~n22595;
  assign n22597 = ~n22533 & ~n22596;
  assign n22598 = n22533 & n22596;
  assign n22599 = ~n22597 & ~n22598;
  assign n22600 = ~n22531 & ~n22599;
  assign n22601 = n22531 & n22599;
  assign n22602 = ~n22600 & ~n22601;
  assign n22603 = ~n22070 & n22154;
  assign n22604 = ~n22160 & ~n22603;
  assign n22605 = n22602 & n22604;
  assign n22606 = ~n22602 & ~n22604;
  assign n22607 = ~n22605 & ~n22606;
  assign n22608 = n5240 & n21054;
  assign n22609 = n5241 & n21812;
  assign n22610 = n5853 & n21051;
  assign n22611 = n5866 & n21048;
  assign n22612 = ~n22608 & ~n22610;
  assign n22613 = ~n22611 & n22612;
  assign n22614 = ~n22609 & n22613;
  assign n22615 = pi20  & n22614;
  assign n22616 = ~pi20  & ~n22614;
  assign n22617 = ~n22615 & ~n22616;
  assign n22618 = n22607 & n22617;
  assign n22619 = ~n22607 & ~n22617;
  assign n22620 = ~n22618 & ~n22619;
  assign n22621 = ~n22521 & n22620;
  assign n22622 = n22521 & ~n22620;
  assign n22623 = ~n22621 & ~n22622;
  assign n22624 = ~n22518 & ~n22623;
  assign n22625 = n22518 & n22623;
  assign n22626 = ~n22624 & ~n22625;
  assign n22627 = n22508 & ~n22626;
  assign n22628 = ~n22508 & n22626;
  assign n22629 = ~n22627 & ~n22628;
  assign n22630 = n6630 & n21036;
  assign n22631 = n21159 & ~n21161;
  assign n22632 = ~n21162 & ~n22631;
  assign n22633 = n6631 & n22632;
  assign n22634 = n7238 & n21033;
  assign n22635 = n7262 & n21030;
  assign n22636 = ~n22630 & ~n22634;
  assign n22637 = ~n22635 & n22636;
  assign n22638 = ~n22633 & n22637;
  assign n22639 = pi14  & n22638;
  assign n22640 = ~pi14  & ~n22638;
  assign n22641 = ~n22639 & ~n22640;
  assign n22642 = n22629 & n22641;
  assign n22643 = ~n22629 & ~n22641;
  assign n22644 = ~n22642 & ~n22643;
  assign n22645 = ~n22507 & ~n22644;
  assign n22646 = n22507 & n22644;
  assign n22647 = ~n22645 & ~n22646;
  assign n22648 = ~n21315 & n22647;
  assign n22649 = ~n21315 & ~n22647;
  assign n22650 = n21315 & n22647;
  assign n22651 = ~n22649 & ~n22650;
  assign n22652 = n7430 & n21030;
  assign n22653 = n21167 & ~n21169;
  assign n22654 = ~n21170 & ~n22653;
  assign n22655 = n7431 & n22654;
  assign n22656 = n7869 & n21027;
  assign n22657 = n7895 & n21024;
  assign n22658 = ~n22652 & ~n22656;
  assign n22659 = ~n22657 & n22658;
  assign n22660 = ~n22655 & n22659;
  assign n22661 = ~pi11  & ~n22660;
  assign n22662 = pi11  & n22660;
  assign n22663 = ~n22661 & ~n22662;
  assign n22664 = n22502 & n22505;
  assign n22665 = ~n22506 & ~n22664;
  assign n22666 = ~n22663 & n22665;
  assign n22667 = ~n22663 & ~n22665;
  assign n22668 = n22663 & n22665;
  assign n22669 = ~n22667 & ~n22668;
  assign n22670 = n22214 & n22500;
  assign n22671 = ~n22501 & ~n22670;
  assign n22672 = n7430 & n21033;
  assign n22673 = n21163 & ~n21165;
  assign n22674 = ~n21166 & ~n22673;
  assign n22675 = n7431 & n22674;
  assign n22676 = n7869 & n21030;
  assign n22677 = n7895 & n21027;
  assign n22678 = ~n22672 & ~n22676;
  assign n22679 = ~n22677 & n22678;
  assign n22680 = ~n22675 & n22679;
  assign n22681 = pi11  & n22680;
  assign n22682 = ~pi11  & ~n22680;
  assign n22683 = ~n22681 & ~n22682;
  assign n22684 = n22671 & ~n22683;
  assign n22685 = n22232 & n22498;
  assign n22686 = ~n22499 & ~n22685;
  assign n22687 = n7430 & n21036;
  assign n22688 = n7431 & n22632;
  assign n22689 = n7869 & n21033;
  assign n22690 = n7895 & n21030;
  assign n22691 = ~n22687 & ~n22689;
  assign n22692 = ~n22690 & n22691;
  assign n22693 = ~n22688 & n22692;
  assign n22694 = pi11  & n22693;
  assign n22695 = ~pi11  & ~n22693;
  assign n22696 = ~n22694 & ~n22695;
  assign n22697 = n22686 & ~n22696;
  assign n22698 = n7430 & n21039;
  assign n22699 = n7431 & n22186;
  assign n22700 = n7869 & n21036;
  assign n22701 = n7895 & n21033;
  assign n22702 = ~n22698 & ~n22700;
  assign n22703 = ~n22701 & n22702;
  assign n22704 = ~n22699 & n22703;
  assign n22705 = ~pi11  & ~n22704;
  assign n22706 = pi11  & n22704;
  assign n22707 = ~n22705 & ~n22706;
  assign n22708 = n22494 & ~n22496;
  assign n22709 = ~n22497 & ~n22708;
  assign n22710 = ~n22707 & n22709;
  assign n22711 = ~n22707 & ~n22709;
  assign n22712 = n22707 & n22709;
  assign n22713 = ~n22711 & ~n22712;
  assign n22714 = n7430 & n21042;
  assign n22715 = n7431 & n22199;
  assign n22716 = n7869 & n21039;
  assign n22717 = n7895 & n21036;
  assign n22718 = ~n22714 & ~n22716;
  assign n22719 = ~n22717 & n22718;
  assign n22720 = ~n22715 & n22719;
  assign n22721 = ~pi11  & ~n22720;
  assign n22722 = pi11  & n22720;
  assign n22723 = ~n22721 & ~n22722;
  assign n22724 = ~n22489 & n22492;
  assign n22725 = n22489 & ~n22492;
  assign n22726 = ~n22724 & ~n22725;
  assign n22727 = ~n22723 & ~n22726;
  assign n22728 = n7430 & n21045;
  assign n22729 = n7431 & n22217;
  assign n22730 = n7869 & n21042;
  assign n22731 = n7895 & n21039;
  assign n22732 = ~n22728 & ~n22730;
  assign n22733 = ~n22731 & n22732;
  assign n22734 = ~n22729 & n22733;
  assign n22735 = ~pi11  & ~n22734;
  assign n22736 = pi11  & n22734;
  assign n22737 = ~n22735 & ~n22736;
  assign n22738 = n22484 & n22487;
  assign n22739 = ~n22488 & ~n22738;
  assign n22740 = ~n22737 & n22739;
  assign n22741 = ~n22737 & ~n22739;
  assign n22742 = n22737 & n22739;
  assign n22743 = ~n22741 & ~n22742;
  assign n22744 = n22287 & n22482;
  assign n22745 = ~n22483 & ~n22744;
  assign n22746 = n7430 & n21048;
  assign n22747 = n7431 & n22049;
  assign n22748 = n7869 & n21045;
  assign n22749 = n7895 & n21042;
  assign n22750 = ~n22746 & ~n22748;
  assign n22751 = ~n22749 & n22750;
  assign n22752 = ~n22747 & n22751;
  assign n22753 = pi11  & n22752;
  assign n22754 = ~pi11  & ~n22752;
  assign n22755 = ~n22753 & ~n22754;
  assign n22756 = n22745 & ~n22755;
  assign n22757 = n22303 & n22480;
  assign n22758 = ~n22481 & ~n22757;
  assign n22759 = n7430 & n21051;
  assign n22760 = n7431 & n21797;
  assign n22761 = n7869 & n21048;
  assign n22762 = n7895 & n21045;
  assign n22763 = ~n22759 & ~n22761;
  assign n22764 = ~n22762 & n22763;
  assign n22765 = ~n22760 & n22764;
  assign n22766 = pi11  & n22765;
  assign n22767 = ~pi11  & ~n22765;
  assign n22768 = ~n22766 & ~n22767;
  assign n22769 = n22758 & ~n22768;
  assign n22770 = n22476 & ~n22478;
  assign n22771 = ~n22479 & ~n22770;
  assign n22772 = n7430 & n21054;
  assign n22773 = n7431 & n21812;
  assign n22774 = n7869 & n21051;
  assign n22775 = n7895 & n21048;
  assign n22776 = ~n22772 & ~n22774;
  assign n22777 = ~n22775 & n22776;
  assign n22778 = ~n22773 & n22777;
  assign n22779 = pi11  & n22778;
  assign n22780 = ~pi11  & ~n22778;
  assign n22781 = ~n22779 & ~n22780;
  assign n22782 = n22771 & ~n22781;
  assign n22783 = n7430 & n21057;
  assign n22784 = n7431 & n21825;
  assign n22785 = n7869 & n21054;
  assign n22786 = n7895 & n21051;
  assign n22787 = ~n22783 & ~n22785;
  assign n22788 = ~n22786 & n22787;
  assign n22789 = ~n22784 & n22788;
  assign n22790 = ~pi11  & ~n22789;
  assign n22791 = pi11  & n22789;
  assign n22792 = ~n22790 & ~n22791;
  assign n22793 = n22472 & ~n22474;
  assign n22794 = ~n22475 & ~n22793;
  assign n22795 = ~n22792 & n22794;
  assign n22796 = ~n22792 & ~n22794;
  assign n22797 = n22792 & n22794;
  assign n22798 = ~n22796 & ~n22797;
  assign n22799 = n7430 & n21060;
  assign n22800 = n7431 & n21318;
  assign n22801 = n7869 & n21057;
  assign n22802 = n7895 & n21054;
  assign n22803 = ~n22799 & ~n22801;
  assign n22804 = ~n22802 & n22803;
  assign n22805 = ~n22800 & n22804;
  assign n22806 = ~pi11  & ~n22805;
  assign n22807 = pi11  & n22805;
  assign n22808 = ~n22806 & ~n22807;
  assign n22809 = n22467 & n22470;
  assign n22810 = ~n22471 & ~n22809;
  assign n22811 = ~n22808 & n22810;
  assign n22812 = ~n22808 & ~n22810;
  assign n22813 = n22808 & n22810;
  assign n22814 = ~n22812 & ~n22813;
  assign n22815 = n7430 & n21063;
  assign n22816 = n7431 & n21613;
  assign n22817 = n7869 & n21060;
  assign n22818 = n7895 & n21057;
  assign n22819 = ~n22815 & ~n22817;
  assign n22820 = ~n22818 & n22819;
  assign n22821 = ~n22816 & n22820;
  assign n22822 = ~pi11  & ~n22821;
  assign n22823 = pi11  & n22821;
  assign n22824 = ~n22822 & ~n22823;
  assign n22825 = ~n22462 & n22465;
  assign n22826 = n22462 & ~n22465;
  assign n22827 = ~n22825 & ~n22826;
  assign n22828 = ~n22824 & ~n22827;
  assign n22829 = n22372 & n22460;
  assign n22830 = ~n22461 & ~n22829;
  assign n22831 = n7430 & n21066;
  assign n22832 = n7431 & n21631;
  assign n22833 = n7869 & n21063;
  assign n22834 = n7895 & n21060;
  assign n22835 = ~n22831 & ~n22833;
  assign n22836 = ~n22834 & n22835;
  assign n22837 = ~n22832 & n22836;
  assign n22838 = pi11  & n22837;
  assign n22839 = ~pi11  & ~n22837;
  assign n22840 = ~n22838 & ~n22839;
  assign n22841 = n22830 & ~n22840;
  assign n22842 = n22456 & ~n22458;
  assign n22843 = ~n22459 & ~n22842;
  assign n22844 = n7430 & n21069;
  assign n22845 = n7431 & n21592;
  assign n22846 = n7869 & n21066;
  assign n22847 = n7895 & n21063;
  assign n22848 = ~n22844 & ~n22846;
  assign n22849 = ~n22847 & n22848;
  assign n22850 = ~n22845 & n22849;
  assign n22851 = pi11  & n22850;
  assign n22852 = ~pi11  & ~n22850;
  assign n22853 = ~n22851 & ~n22852;
  assign n22854 = n22843 & ~n22853;
  assign n22855 = n22403 & n22454;
  assign n22856 = ~n22455 & ~n22855;
  assign n22857 = n7430 & n21072;
  assign n22858 = n7431 & n21428;
  assign n22859 = n7869 & n21069;
  assign n22860 = n7895 & n21066;
  assign n22861 = ~n22857 & ~n22859;
  assign n22862 = ~n22860 & n22861;
  assign n22863 = ~n22858 & n22862;
  assign n22864 = pi11  & n22863;
  assign n22865 = ~pi11  & ~n22863;
  assign n22866 = ~n22864 & ~n22865;
  assign n22867 = n22856 & ~n22866;
  assign n22868 = n7430 & n21075;
  assign n22869 = n7431 & n21441;
  assign n22870 = n7869 & n21072;
  assign n22871 = n7895 & n21069;
  assign n22872 = ~n22868 & ~n22870;
  assign n22873 = ~n22871 & n22872;
  assign n22874 = ~n22869 & n22873;
  assign n22875 = ~pi11  & ~n22874;
  assign n22876 = pi11  & n22874;
  assign n22877 = ~n22875 & ~n22876;
  assign n22878 = n22450 & ~n22452;
  assign n22879 = ~n22453 & ~n22878;
  assign n22880 = ~n22877 & n22879;
  assign n22881 = ~n22877 & ~n22879;
  assign n22882 = n22877 & n22879;
  assign n22883 = ~n22881 & ~n22882;
  assign n22884 = n7430 & n21078;
  assign n22885 = n7431 & n21459;
  assign n22886 = n7869 & n21075;
  assign n22887 = n7895 & n21072;
  assign n22888 = ~n22884 & ~n22886;
  assign n22889 = ~n22887 & n22888;
  assign n22890 = ~n22885 & n22889;
  assign n22891 = pi11  & n22890;
  assign n22892 = ~pi11  & ~n22890;
  assign n22893 = ~n22891 & ~n22892;
  assign n22894 = n22438 & n22448;
  assign n22895 = ~n22449 & ~n22894;
  assign n22896 = ~n22893 & n22895;
  assign n22897 = n7430 & n21081;
  assign n22898 = n7431 & n21330;
  assign n22899 = n7869 & n21078;
  assign n22900 = n7895 & n21075;
  assign n22901 = ~n22897 & ~n22899;
  assign n22902 = ~n22900 & n22901;
  assign n22903 = ~n22898 & n22902;
  assign n22904 = ~pi11  & ~n22903;
  assign n22905 = pi11  & n22903;
  assign n22906 = ~n22904 & ~n22905;
  assign n22907 = pi14  & ~n22426;
  assign n22908 = n22433 & ~n22907;
  assign n22909 = ~n22433 & n22907;
  assign n22910 = ~n22908 & ~n22909;
  assign n22911 = ~n22906 & n22910;
  assign n22912 = ~n22906 & ~n22910;
  assign n22913 = n22906 & n22910;
  assign n22914 = ~n22912 & ~n22913;
  assign n22915 = n7430 & n21084;
  assign n22916 = n7431 & n21370;
  assign n22917 = n7869 & n21081;
  assign n22918 = n7895 & n21078;
  assign n22919 = ~n22915 & ~n22917;
  assign n22920 = ~n22918 & n22919;
  assign n22921 = ~n22916 & n22920;
  assign n22922 = pi11  & n22921;
  assign n22923 = ~pi11  & ~n22921;
  assign n22924 = ~n22922 & ~n22923;
  assign n22925 = pi14  & n22419;
  assign n22926 = ~n22424 & n22925;
  assign n22927 = n22424 & ~n22925;
  assign n22928 = ~n22926 & ~n22927;
  assign n22929 = ~n22924 & n22928;
  assign n22930 = ~n7425 & n21091;
  assign n22931 = n7869 & n21091;
  assign n22932 = n7895 & n21089;
  assign n22933 = n7431 & ~n21345;
  assign n22934 = ~n22931 & ~n22932;
  assign n22935 = ~n22933 & n22934;
  assign n22936 = pi11  & ~n22930;
  assign n22937 = n22935 & n22936;
  assign n22938 = n7430 & n21091;
  assign n22939 = n7431 & ~n21355;
  assign n22940 = n7869 & n21089;
  assign n22941 = n7895 & n21084;
  assign n22942 = ~n22938 & ~n22940;
  assign n22943 = ~n22941 & n22942;
  assign n22944 = ~n22939 & n22943;
  assign n22945 = n22937 & n22944;
  assign n22946 = n22419 & n22945;
  assign n22947 = ~n22419 & n22945;
  assign n22948 = n22419 & ~n22945;
  assign n22949 = ~n22947 & ~n22948;
  assign n22950 = n7430 & n21089;
  assign n22951 = n7431 & n21407;
  assign n22952 = n7869 & n21084;
  assign n22953 = n7895 & n21081;
  assign n22954 = ~n22950 & ~n22952;
  assign n22955 = ~n22953 & n22954;
  assign n22956 = ~n22951 & n22955;
  assign n22957 = pi11  & n22956;
  assign n22958 = ~pi11  & ~n22956;
  assign n22959 = ~n22957 & ~n22958;
  assign n22960 = ~n22949 & ~n22959;
  assign n22961 = ~n22946 & ~n22960;
  assign n22962 = n22924 & ~n22928;
  assign n22963 = ~n22929 & ~n22962;
  assign n22964 = ~n22961 & n22963;
  assign n22965 = ~n22929 & ~n22964;
  assign n22966 = ~n22914 & ~n22965;
  assign n22967 = ~n22911 & ~n22966;
  assign n22968 = n22893 & ~n22895;
  assign n22969 = ~n22896 & ~n22968;
  assign n22970 = ~n22967 & n22969;
  assign n22971 = ~n22896 & ~n22970;
  assign n22972 = ~n22883 & ~n22971;
  assign n22973 = ~n22880 & ~n22972;
  assign n22974 = n22856 & n22866;
  assign n22975 = ~n22856 & ~n22866;
  assign n22976 = ~n22974 & ~n22975;
  assign n22977 = ~n22973 & ~n22976;
  assign n22978 = ~n22867 & ~n22977;
  assign n22979 = n22843 & n22853;
  assign n22980 = ~n22843 & ~n22853;
  assign n22981 = ~n22979 & ~n22980;
  assign n22982 = ~n22978 & ~n22981;
  assign n22983 = ~n22854 & ~n22982;
  assign n22984 = ~n22830 & n22840;
  assign n22985 = ~n22841 & ~n22984;
  assign n22986 = ~n22983 & n22985;
  assign n22987 = ~n22841 & ~n22986;
  assign n22988 = n22824 & n22827;
  assign n22989 = ~n22828 & ~n22988;
  assign n22990 = ~n22987 & n22989;
  assign n22991 = ~n22828 & ~n22990;
  assign n22992 = ~n22814 & ~n22991;
  assign n22993 = ~n22811 & ~n22992;
  assign n22994 = ~n22798 & ~n22993;
  assign n22995 = ~n22795 & ~n22994;
  assign n22996 = n22771 & n22781;
  assign n22997 = ~n22771 & ~n22781;
  assign n22998 = ~n22996 & ~n22997;
  assign n22999 = ~n22995 & ~n22998;
  assign n23000 = ~n22782 & ~n22999;
  assign n23001 = n22758 & n22768;
  assign n23002 = ~n22758 & ~n22768;
  assign n23003 = ~n23001 & ~n23002;
  assign n23004 = ~n23000 & ~n23003;
  assign n23005 = ~n22769 & ~n23004;
  assign n23006 = ~n22745 & n22755;
  assign n23007 = ~n22756 & ~n23006;
  assign n23008 = ~n23005 & n23007;
  assign n23009 = ~n22756 & ~n23008;
  assign n23010 = ~n22743 & ~n23009;
  assign n23011 = ~n22740 & ~n23010;
  assign n23012 = n22723 & n22726;
  assign n23013 = ~n22727 & ~n23012;
  assign n23014 = ~n23011 & n23013;
  assign n23015 = ~n22727 & ~n23014;
  assign n23016 = ~n22713 & ~n23015;
  assign n23017 = ~n22710 & ~n23016;
  assign n23018 = n22686 & n22696;
  assign n23019 = ~n22686 & ~n22696;
  assign n23020 = ~n23018 & ~n23019;
  assign n23021 = ~n23017 & ~n23020;
  assign n23022 = ~n22697 & ~n23021;
  assign n23023 = ~n22671 & n22683;
  assign n23024 = ~n22684 & ~n23023;
  assign n23025 = ~n23022 & n23024;
  assign n23026 = ~n22684 & ~n23025;
  assign n23027 = ~n22669 & ~n23026;
  assign n23028 = ~n22666 & ~n23027;
  assign n23029 = ~n22651 & ~n23028;
  assign n23030 = ~n22648 & ~n23029;
  assign n23031 = n7430 & n21024;
  assign n23032 = n21175 & ~n21177;
  assign n23033 = ~n21178 & ~n23032;
  assign n23034 = n7431 & n23033;
  assign n23035 = n7869 & n21021;
  assign n23036 = n7895 & n21018;
  assign n23037 = ~n23031 & ~n23035;
  assign n23038 = ~n23036 & n23037;
  assign n23039 = ~n23034 & n23038;
  assign n23040 = ~pi11  & ~n23039;
  assign n23041 = pi11  & n23039;
  assign n23042 = ~n23040 & ~n23041;
  assign n23043 = n22629 & ~n22641;
  assign n23044 = ~n22645 & ~n23043;
  assign n23045 = n5982 & n21042;
  assign n23046 = n5983 & n22199;
  assign n23047 = n6323 & n21039;
  assign n23048 = n6336 & n21036;
  assign n23049 = ~n23045 & ~n23047;
  assign n23050 = ~n23048 & n23049;
  assign n23051 = ~n23046 & n23050;
  assign n23052 = ~pi17  & ~n23051;
  assign n23053 = pi17  & n23051;
  assign n23054 = ~n23052 & ~n23053;
  assign n23055 = n22607 & ~n22617;
  assign n23056 = ~n22521 & ~n22620;
  assign n23057 = ~n23055 & ~n23056;
  assign n23058 = ~n22531 & n22599;
  assign n23059 = ~n22606 & ~n23058;
  assign n23060 = n5044 & n21060;
  assign n23061 = n5045 & n21318;
  assign n23062 = n5109 & n21057;
  assign n23063 = n5130 & n21054;
  assign n23064 = ~n23060 & ~n23062;
  assign n23065 = ~n23063 & n23064;
  assign n23066 = ~n23061 & n23065;
  assign n23067 = ~pi23  & ~n23066;
  assign n23068 = pi23  & n23066;
  assign n23069 = ~n23067 & ~n23068;
  assign n23070 = n22583 & ~n22593;
  assign n23071 = ~n22597 & ~n23070;
  assign n23072 = n3810 & n21078;
  assign n23073 = n3886 & n21459;
  assign n23074 = n3884 & n21075;
  assign n23075 = n4380 & n21072;
  assign n23076 = ~n23072 & ~n23074;
  assign n23077 = ~n23075 & n23076;
  assign n23078 = ~n23073 & n23077;
  assign n23079 = ~pi29  & ~n23078;
  assign n23080 = pi29  & n23078;
  assign n23081 = ~n23079 & ~n23080;
  assign n23082 = ~n281 & ~n627;
  assign n23083 = n354 & n23082;
  assign n23084 = ~n274 & ~n299;
  assign n23085 = n2727 & n23084;
  assign n23086 = n164 & n428;
  assign n23087 = n487 & n600;
  assign n23088 = n633 & n1035;
  assign n23089 = n5474 & n23088;
  assign n23090 = n23086 & n23087;
  assign n23091 = n23083 & n23085;
  assign n23092 = n23090 & n23091;
  assign n23093 = n2444 & n23089;
  assign n23094 = n23092 & n23093;
  assign n23095 = n4507 & n5713;
  assign n23096 = n23094 & n23095;
  assign n23097 = n1882 & n23096;
  assign n23098 = n2747 & n23097;
  assign n23099 = n3692 & n21084;
  assign n23100 = n880 & n21407;
  assign n23101 = n748 & n21089;
  assign n23102 = n3694 & n21081;
  assign n23103 = ~n23099 & ~n23101;
  assign n23104 = ~n23102 & n23103;
  assign n23105 = ~n23100 & n23104;
  assign n23106 = ~n23098 & n23105;
  assign n23107 = n23098 & ~n23105;
  assign n23108 = ~n23106 & ~n23107;
  assign n23109 = ~n22566 & ~n22574;
  assign n23110 = ~n22565 & ~n23109;
  assign n23111 = ~n23108 & ~n23110;
  assign n23112 = n23108 & n23110;
  assign n23113 = ~n23111 & ~n23112;
  assign n23114 = ~n23081 & ~n23113;
  assign n23115 = n23081 & n23113;
  assign n23116 = ~n23114 & ~n23115;
  assign n23117 = ~n22578 & ~n22582;
  assign n23118 = n23116 & n23117;
  assign n23119 = ~n23116 & ~n23117;
  assign n23120 = ~n23118 & ~n23119;
  assign n23121 = n86 & n21069;
  assign n23122 = n4420 & n21592;
  assign n23123 = n4600 & n21066;
  assign n23124 = n4615 & n21063;
  assign n23125 = ~n23121 & ~n23123;
  assign n23126 = ~n23124 & n23125;
  assign n23127 = ~n23122 & n23126;
  assign n23128 = pi26  & n23127;
  assign n23129 = ~pi26  & ~n23127;
  assign n23130 = ~n23128 & ~n23129;
  assign n23131 = n23120 & n23130;
  assign n23132 = ~n23120 & ~n23130;
  assign n23133 = ~n23131 & ~n23132;
  assign n23134 = ~n23071 & n23133;
  assign n23135 = n23071 & ~n23133;
  assign n23136 = ~n23134 & ~n23135;
  assign n23137 = ~n23069 & ~n23136;
  assign n23138 = n23069 & n23136;
  assign n23139 = ~n23137 & ~n23138;
  assign n23140 = n23059 & ~n23139;
  assign n23141 = ~n23059 & n23139;
  assign n23142 = ~n23140 & ~n23141;
  assign n23143 = n5240 & n21051;
  assign n23144 = n5241 & n21797;
  assign n23145 = n5853 & n21048;
  assign n23146 = n5866 & n21045;
  assign n23147 = ~n23143 & ~n23145;
  assign n23148 = ~n23146 & n23147;
  assign n23149 = ~n23144 & n23148;
  assign n23150 = pi20  & n23149;
  assign n23151 = ~pi20  & ~n23149;
  assign n23152 = ~n23150 & ~n23151;
  assign n23153 = n23142 & n23152;
  assign n23154 = ~n23142 & ~n23152;
  assign n23155 = ~n23153 & ~n23154;
  assign n23156 = ~n23057 & ~n23155;
  assign n23157 = n23057 & n23155;
  assign n23158 = ~n23156 & ~n23157;
  assign n23159 = ~n23054 & ~n23158;
  assign n23160 = n23054 & n23158;
  assign n23161 = ~n23159 & ~n23160;
  assign n23162 = ~n22624 & ~n22628;
  assign n23163 = n23161 & n23162;
  assign n23164 = ~n23161 & ~n23162;
  assign n23165 = ~n23163 & ~n23164;
  assign n23166 = n6630 & n21033;
  assign n23167 = n6631 & n22674;
  assign n23168 = n7238 & n21030;
  assign n23169 = n7262 & n21027;
  assign n23170 = ~n23166 & ~n23168;
  assign n23171 = ~n23169 & n23170;
  assign n23172 = ~n23167 & n23171;
  assign n23173 = pi14  & n23172;
  assign n23174 = ~pi14  & ~n23172;
  assign n23175 = ~n23173 & ~n23174;
  assign n23176 = n23165 & n23175;
  assign n23177 = ~n23165 & ~n23175;
  assign n23178 = ~n23176 & ~n23177;
  assign n23179 = ~n23044 & n23178;
  assign n23180 = n23044 & ~n23178;
  assign n23181 = ~n23179 & ~n23180;
  assign n23182 = ~n23042 & ~n23181;
  assign n23183 = n23042 & n23181;
  assign n23184 = ~n23182 & ~n23183;
  assign n23185 = n23030 & ~n23184;
  assign n23186 = ~n23030 & n23184;
  assign n23187 = ~n23185 & ~n23186;
  assign n23188 = n8250 & n21015;
  assign n23189 = n21187 & ~n21189;
  assign n23190 = ~n21190 & ~n23189;
  assign n23191 = n8251 & n23190;
  assign n23192 = n9016 & n21012;
  assign n23193 = n9040 & n21009;
  assign n23194 = ~n23188 & ~n23192;
  assign n23195 = ~n23193 & n23194;
  assign n23196 = ~n23191 & n23195;
  assign n23197 = pi8  & n23196;
  assign n23198 = ~pi8  & ~n23196;
  assign n23199 = ~n23197 & ~n23198;
  assign n23200 = n23187 & ~n23199;
  assign n23201 = n22651 & n23028;
  assign n23202 = ~n23029 & ~n23201;
  assign n23203 = n8250 & n21018;
  assign n23204 = n21183 & ~n21185;
  assign n23205 = ~n21186 & ~n23204;
  assign n23206 = n8251 & n23205;
  assign n23207 = n9016 & n21015;
  assign n23208 = n9040 & n21012;
  assign n23209 = ~n23203 & ~n23207;
  assign n23210 = ~n23208 & n23209;
  assign n23211 = ~n23206 & n23210;
  assign n23212 = pi8  & n23211;
  assign n23213 = ~pi8  & ~n23211;
  assign n23214 = ~n23212 & ~n23213;
  assign n23215 = n23202 & ~n23214;
  assign n23216 = n22669 & n23026;
  assign n23217 = ~n23027 & ~n23216;
  assign n23218 = n8250 & n21021;
  assign n23219 = n21179 & ~n21181;
  assign n23220 = ~n21182 & ~n23219;
  assign n23221 = n8251 & n23220;
  assign n23222 = n9016 & n21018;
  assign n23223 = n9040 & n21015;
  assign n23224 = ~n23218 & ~n23222;
  assign n23225 = ~n23223 & n23224;
  assign n23226 = ~n23221 & n23225;
  assign n23227 = pi8  & n23226;
  assign n23228 = ~pi8  & ~n23226;
  assign n23229 = ~n23227 & ~n23228;
  assign n23230 = n23217 & ~n23229;
  assign n23231 = n8250 & n21024;
  assign n23232 = n8251 & n23033;
  assign n23233 = n9016 & n21021;
  assign n23234 = n9040 & n21018;
  assign n23235 = ~n23231 & ~n23233;
  assign n23236 = ~n23234 & n23235;
  assign n23237 = ~n23232 & n23236;
  assign n23238 = ~pi8  & ~n23237;
  assign n23239 = pi8  & n23237;
  assign n23240 = ~n23238 & ~n23239;
  assign n23241 = n23022 & ~n23024;
  assign n23242 = ~n23025 & ~n23241;
  assign n23243 = ~n23240 & n23242;
  assign n23244 = ~n23240 & ~n23242;
  assign n23245 = n23240 & n23242;
  assign n23246 = ~n23244 & ~n23245;
  assign n23247 = n8250 & n21027;
  assign n23248 = n8251 & n21306;
  assign n23249 = n9016 & n21024;
  assign n23250 = n9040 & n21021;
  assign n23251 = ~n23247 & ~n23249;
  assign n23252 = ~n23250 & n23251;
  assign n23253 = ~n23248 & n23252;
  assign n23254 = ~pi8  & ~n23253;
  assign n23255 = pi8  & n23253;
  assign n23256 = ~n23254 & ~n23255;
  assign n23257 = ~n23017 & n23020;
  assign n23258 = n23017 & ~n23020;
  assign n23259 = ~n23257 & ~n23258;
  assign n23260 = ~n23256 & ~n23259;
  assign n23261 = n22713 & n23015;
  assign n23262 = ~n23016 & ~n23261;
  assign n23263 = n8250 & n21030;
  assign n23264 = n8251 & n22654;
  assign n23265 = n9016 & n21027;
  assign n23266 = n9040 & n21024;
  assign n23267 = ~n23263 & ~n23265;
  assign n23268 = ~n23266 & n23267;
  assign n23269 = ~n23264 & n23268;
  assign n23270 = pi8  & n23269;
  assign n23271 = ~pi8  & ~n23269;
  assign n23272 = ~n23270 & ~n23271;
  assign n23273 = n23262 & ~n23272;
  assign n23274 = n23011 & ~n23013;
  assign n23275 = ~n23014 & ~n23274;
  assign n23276 = n8250 & n21033;
  assign n23277 = n8251 & n22674;
  assign n23278 = n9016 & n21030;
  assign n23279 = n9040 & n21027;
  assign n23280 = ~n23276 & ~n23278;
  assign n23281 = ~n23279 & n23280;
  assign n23282 = ~n23277 & n23281;
  assign n23283 = pi8  & n23282;
  assign n23284 = ~pi8  & ~n23282;
  assign n23285 = ~n23283 & ~n23284;
  assign n23286 = n23275 & ~n23285;
  assign n23287 = n22743 & n23009;
  assign n23288 = ~n23010 & ~n23287;
  assign n23289 = n8250 & n21036;
  assign n23290 = n8251 & n22632;
  assign n23291 = n9016 & n21033;
  assign n23292 = n9040 & n21030;
  assign n23293 = ~n23289 & ~n23291;
  assign n23294 = ~n23292 & n23293;
  assign n23295 = ~n23290 & n23294;
  assign n23296 = pi8  & n23295;
  assign n23297 = ~pi8  & ~n23295;
  assign n23298 = ~n23296 & ~n23297;
  assign n23299 = n23288 & ~n23298;
  assign n23300 = n8250 & n21039;
  assign n23301 = n8251 & n22186;
  assign n23302 = n9016 & n21036;
  assign n23303 = n9040 & n21033;
  assign n23304 = ~n23300 & ~n23302;
  assign n23305 = ~n23303 & n23304;
  assign n23306 = ~n23301 & n23305;
  assign n23307 = ~pi8  & ~n23306;
  assign n23308 = pi8  & n23306;
  assign n23309 = ~n23307 & ~n23308;
  assign n23310 = n23005 & ~n23007;
  assign n23311 = ~n23008 & ~n23310;
  assign n23312 = ~n23309 & n23311;
  assign n23313 = ~n23309 & ~n23311;
  assign n23314 = n23309 & n23311;
  assign n23315 = ~n23313 & ~n23314;
  assign n23316 = n8250 & n21042;
  assign n23317 = n8251 & n22199;
  assign n23318 = n9016 & n21039;
  assign n23319 = n9040 & n21036;
  assign n23320 = ~n23316 & ~n23318;
  assign n23321 = ~n23319 & n23320;
  assign n23322 = ~n23317 & n23321;
  assign n23323 = ~pi8  & ~n23322;
  assign n23324 = pi8  & n23322;
  assign n23325 = ~n23323 & ~n23324;
  assign n23326 = ~n23000 & n23003;
  assign n23327 = n23000 & ~n23003;
  assign n23328 = ~n23326 & ~n23327;
  assign n23329 = ~n23325 & ~n23328;
  assign n23330 = n8250 & n21045;
  assign n23331 = n8251 & n22217;
  assign n23332 = n9016 & n21042;
  assign n23333 = n9040 & n21039;
  assign n23334 = ~n23330 & ~n23332;
  assign n23335 = ~n23333 & n23334;
  assign n23336 = ~n23331 & n23335;
  assign n23337 = ~pi8  & ~n23336;
  assign n23338 = pi8  & n23336;
  assign n23339 = ~n23337 & ~n23338;
  assign n23340 = n22995 & n22998;
  assign n23341 = ~n22999 & ~n23340;
  assign n23342 = ~n23339 & n23341;
  assign n23343 = ~n23339 & ~n23341;
  assign n23344 = n23339 & n23341;
  assign n23345 = ~n23343 & ~n23344;
  assign n23346 = n22798 & n22993;
  assign n23347 = ~n22994 & ~n23346;
  assign n23348 = n8250 & n21048;
  assign n23349 = n8251 & n22049;
  assign n23350 = n9016 & n21045;
  assign n23351 = n9040 & n21042;
  assign n23352 = ~n23348 & ~n23350;
  assign n23353 = ~n23351 & n23352;
  assign n23354 = ~n23349 & n23353;
  assign n23355 = pi8  & n23354;
  assign n23356 = ~pi8  & ~n23354;
  assign n23357 = ~n23355 & ~n23356;
  assign n23358 = n23347 & ~n23357;
  assign n23359 = n22814 & n22991;
  assign n23360 = ~n22992 & ~n23359;
  assign n23361 = n8250 & n21051;
  assign n23362 = n8251 & n21797;
  assign n23363 = n9016 & n21048;
  assign n23364 = n9040 & n21045;
  assign n23365 = ~n23361 & ~n23363;
  assign n23366 = ~n23364 & n23365;
  assign n23367 = ~n23362 & n23366;
  assign n23368 = pi8  & n23367;
  assign n23369 = ~pi8  & ~n23367;
  assign n23370 = ~n23368 & ~n23369;
  assign n23371 = n23360 & ~n23370;
  assign n23372 = n22987 & ~n22989;
  assign n23373 = ~n22990 & ~n23372;
  assign n23374 = n8250 & n21054;
  assign n23375 = n8251 & n21812;
  assign n23376 = n9016 & n21051;
  assign n23377 = n9040 & n21048;
  assign n23378 = ~n23374 & ~n23376;
  assign n23379 = ~n23377 & n23378;
  assign n23380 = ~n23375 & n23379;
  assign n23381 = pi8  & n23380;
  assign n23382 = ~pi8  & ~n23380;
  assign n23383 = ~n23381 & ~n23382;
  assign n23384 = n23373 & ~n23383;
  assign n23385 = n8250 & n21057;
  assign n23386 = n8251 & n21825;
  assign n23387 = n9016 & n21054;
  assign n23388 = n9040 & n21051;
  assign n23389 = ~n23385 & ~n23387;
  assign n23390 = ~n23388 & n23389;
  assign n23391 = ~n23386 & n23390;
  assign n23392 = ~pi8  & ~n23391;
  assign n23393 = pi8  & n23391;
  assign n23394 = ~n23392 & ~n23393;
  assign n23395 = n22983 & ~n22985;
  assign n23396 = ~n22986 & ~n23395;
  assign n23397 = ~n23394 & n23396;
  assign n23398 = ~n23394 & ~n23396;
  assign n23399 = n23394 & n23396;
  assign n23400 = ~n23398 & ~n23399;
  assign n23401 = n8250 & n21060;
  assign n23402 = n8251 & n21318;
  assign n23403 = n9016 & n21057;
  assign n23404 = n9040 & n21054;
  assign n23405 = ~n23401 & ~n23403;
  assign n23406 = ~n23404 & n23405;
  assign n23407 = ~n23402 & n23406;
  assign n23408 = ~pi8  & ~n23407;
  assign n23409 = pi8  & n23407;
  assign n23410 = ~n23408 & ~n23409;
  assign n23411 = n22978 & n22981;
  assign n23412 = ~n22982 & ~n23411;
  assign n23413 = ~n23410 & n23412;
  assign n23414 = ~n23410 & ~n23412;
  assign n23415 = n23410 & n23412;
  assign n23416 = ~n23414 & ~n23415;
  assign n23417 = n8250 & n21063;
  assign n23418 = n8251 & n21613;
  assign n23419 = n9016 & n21060;
  assign n23420 = n9040 & n21057;
  assign n23421 = ~n23417 & ~n23419;
  assign n23422 = ~n23420 & n23421;
  assign n23423 = ~n23418 & n23422;
  assign n23424 = ~pi8  & ~n23423;
  assign n23425 = pi8  & n23423;
  assign n23426 = ~n23424 & ~n23425;
  assign n23427 = ~n22973 & n22976;
  assign n23428 = n22973 & ~n22976;
  assign n23429 = ~n23427 & ~n23428;
  assign n23430 = ~n23426 & ~n23429;
  assign n23431 = n22883 & n22971;
  assign n23432 = ~n22972 & ~n23431;
  assign n23433 = n8250 & n21066;
  assign n23434 = n8251 & n21631;
  assign n23435 = n9016 & n21063;
  assign n23436 = n9040 & n21060;
  assign n23437 = ~n23433 & ~n23435;
  assign n23438 = ~n23436 & n23437;
  assign n23439 = ~n23434 & n23438;
  assign n23440 = pi8  & n23439;
  assign n23441 = ~pi8  & ~n23439;
  assign n23442 = ~n23440 & ~n23441;
  assign n23443 = n23432 & ~n23442;
  assign n23444 = n22967 & ~n22969;
  assign n23445 = ~n22970 & ~n23444;
  assign n23446 = n8250 & n21069;
  assign n23447 = n8251 & n21592;
  assign n23448 = n9016 & n21066;
  assign n23449 = n9040 & n21063;
  assign n23450 = ~n23446 & ~n23448;
  assign n23451 = ~n23449 & n23450;
  assign n23452 = ~n23447 & n23451;
  assign n23453 = pi8  & n23452;
  assign n23454 = ~pi8  & ~n23452;
  assign n23455 = ~n23453 & ~n23454;
  assign n23456 = n23445 & ~n23455;
  assign n23457 = n22914 & n22965;
  assign n23458 = ~n22966 & ~n23457;
  assign n23459 = n8250 & n21072;
  assign n23460 = n8251 & n21428;
  assign n23461 = n9016 & n21069;
  assign n23462 = n9040 & n21066;
  assign n23463 = ~n23459 & ~n23461;
  assign n23464 = ~n23462 & n23463;
  assign n23465 = ~n23460 & n23464;
  assign n23466 = pi8  & n23465;
  assign n23467 = ~pi8  & ~n23465;
  assign n23468 = ~n23466 & ~n23467;
  assign n23469 = n23458 & ~n23468;
  assign n23470 = n8250 & n21075;
  assign n23471 = n8251 & n21441;
  assign n23472 = n9016 & n21072;
  assign n23473 = n9040 & n21069;
  assign n23474 = ~n23470 & ~n23472;
  assign n23475 = ~n23473 & n23474;
  assign n23476 = ~n23471 & n23475;
  assign n23477 = ~pi8  & ~n23476;
  assign n23478 = pi8  & n23476;
  assign n23479 = ~n23477 & ~n23478;
  assign n23480 = n22961 & ~n22963;
  assign n23481 = ~n22964 & ~n23480;
  assign n23482 = ~n23479 & n23481;
  assign n23483 = ~n23479 & ~n23481;
  assign n23484 = n23479 & n23481;
  assign n23485 = ~n23483 & ~n23484;
  assign n23486 = n8250 & n21078;
  assign n23487 = n8251 & n21459;
  assign n23488 = n9016 & n21075;
  assign n23489 = n9040 & n21072;
  assign n23490 = ~n23486 & ~n23488;
  assign n23491 = ~n23489 & n23490;
  assign n23492 = ~n23487 & n23491;
  assign n23493 = pi8  & n23492;
  assign n23494 = ~pi8  & ~n23492;
  assign n23495 = ~n23493 & ~n23494;
  assign n23496 = n22949 & n22959;
  assign n23497 = ~n22960 & ~n23496;
  assign n23498 = ~n23495 & n23497;
  assign n23499 = n8250 & n21081;
  assign n23500 = n8251 & n21330;
  assign n23501 = n9016 & n21078;
  assign n23502 = n9040 & n21075;
  assign n23503 = ~n23499 & ~n23501;
  assign n23504 = ~n23502 & n23503;
  assign n23505 = ~n23500 & n23504;
  assign n23506 = ~pi8  & ~n23505;
  assign n23507 = pi8  & n23505;
  assign n23508 = ~n23506 & ~n23507;
  assign n23509 = pi11  & ~n22937;
  assign n23510 = n22944 & ~n23509;
  assign n23511 = ~n22944 & n23509;
  assign n23512 = ~n23510 & ~n23511;
  assign n23513 = ~n23508 & n23512;
  assign n23514 = ~n23508 & ~n23512;
  assign n23515 = n23508 & n23512;
  assign n23516 = ~n23514 & ~n23515;
  assign n23517 = n8250 & n21084;
  assign n23518 = n8251 & n21370;
  assign n23519 = n9016 & n21081;
  assign n23520 = n9040 & n21078;
  assign n23521 = ~n23517 & ~n23519;
  assign n23522 = ~n23520 & n23521;
  assign n23523 = ~n23518 & n23522;
  assign n23524 = pi8  & n23523;
  assign n23525 = ~pi8  & ~n23523;
  assign n23526 = ~n23524 & ~n23525;
  assign n23527 = pi11  & n22930;
  assign n23528 = ~n22935 & n23527;
  assign n23529 = n22935 & ~n23527;
  assign n23530 = ~n23528 & ~n23529;
  assign n23531 = ~n23526 & n23530;
  assign n23532 = ~n8245 & n21091;
  assign n23533 = n9016 & n21091;
  assign n23534 = n9040 & n21089;
  assign n23535 = n8251 & ~n21345;
  assign n23536 = ~n23533 & ~n23534;
  assign n23537 = ~n23535 & n23536;
  assign n23538 = pi8  & ~n23532;
  assign n23539 = n23537 & n23538;
  assign n23540 = n8250 & n21091;
  assign n23541 = n8251 & ~n21355;
  assign n23542 = n9016 & n21089;
  assign n23543 = n9040 & n21084;
  assign n23544 = ~n23540 & ~n23542;
  assign n23545 = ~n23543 & n23544;
  assign n23546 = ~n23541 & n23545;
  assign n23547 = n23539 & n23546;
  assign n23548 = n22930 & n23547;
  assign n23549 = ~n22930 & n23547;
  assign n23550 = n22930 & ~n23547;
  assign n23551 = ~n23549 & ~n23550;
  assign n23552 = n8250 & n21089;
  assign n23553 = n8251 & n21407;
  assign n23554 = n9016 & n21084;
  assign n23555 = n9040 & n21081;
  assign n23556 = ~n23552 & ~n23554;
  assign n23557 = ~n23555 & n23556;
  assign n23558 = ~n23553 & n23557;
  assign n23559 = pi8  & n23558;
  assign n23560 = ~pi8  & ~n23558;
  assign n23561 = ~n23559 & ~n23560;
  assign n23562 = ~n23551 & ~n23561;
  assign n23563 = ~n23548 & ~n23562;
  assign n23564 = n23526 & ~n23530;
  assign n23565 = ~n23531 & ~n23564;
  assign n23566 = ~n23563 & n23565;
  assign n23567 = ~n23531 & ~n23566;
  assign n23568 = ~n23516 & ~n23567;
  assign n23569 = ~n23513 & ~n23568;
  assign n23570 = n23495 & ~n23497;
  assign n23571 = ~n23498 & ~n23570;
  assign n23572 = ~n23569 & n23571;
  assign n23573 = ~n23498 & ~n23572;
  assign n23574 = ~n23485 & ~n23573;
  assign n23575 = ~n23482 & ~n23574;
  assign n23576 = n23458 & n23468;
  assign n23577 = ~n23458 & ~n23468;
  assign n23578 = ~n23576 & ~n23577;
  assign n23579 = ~n23575 & ~n23578;
  assign n23580 = ~n23469 & ~n23579;
  assign n23581 = n23445 & n23455;
  assign n23582 = ~n23445 & ~n23455;
  assign n23583 = ~n23581 & ~n23582;
  assign n23584 = ~n23580 & ~n23583;
  assign n23585 = ~n23456 & ~n23584;
  assign n23586 = ~n23432 & n23442;
  assign n23587 = ~n23443 & ~n23586;
  assign n23588 = ~n23585 & n23587;
  assign n23589 = ~n23443 & ~n23588;
  assign n23590 = n23426 & n23429;
  assign n23591 = ~n23430 & ~n23590;
  assign n23592 = ~n23589 & n23591;
  assign n23593 = ~n23430 & ~n23592;
  assign n23594 = ~n23416 & ~n23593;
  assign n23595 = ~n23413 & ~n23594;
  assign n23596 = ~n23400 & ~n23595;
  assign n23597 = ~n23397 & ~n23596;
  assign n23598 = n23373 & n23383;
  assign n23599 = ~n23373 & ~n23383;
  assign n23600 = ~n23598 & ~n23599;
  assign n23601 = ~n23597 & ~n23600;
  assign n23602 = ~n23384 & ~n23601;
  assign n23603 = n23360 & n23370;
  assign n23604 = ~n23360 & ~n23370;
  assign n23605 = ~n23603 & ~n23604;
  assign n23606 = ~n23602 & ~n23605;
  assign n23607 = ~n23371 & ~n23606;
  assign n23608 = ~n23347 & n23357;
  assign n23609 = ~n23358 & ~n23608;
  assign n23610 = ~n23607 & n23609;
  assign n23611 = ~n23358 & ~n23610;
  assign n23612 = ~n23345 & ~n23611;
  assign n23613 = ~n23342 & ~n23612;
  assign n23614 = n23325 & n23328;
  assign n23615 = ~n23329 & ~n23614;
  assign n23616 = ~n23613 & n23615;
  assign n23617 = ~n23329 & ~n23616;
  assign n23618 = ~n23315 & ~n23617;
  assign n23619 = ~n23312 & ~n23618;
  assign n23620 = n23288 & n23298;
  assign n23621 = ~n23288 & ~n23298;
  assign n23622 = ~n23620 & ~n23621;
  assign n23623 = ~n23619 & ~n23622;
  assign n23624 = ~n23299 & ~n23623;
  assign n23625 = n23275 & n23285;
  assign n23626 = ~n23275 & ~n23285;
  assign n23627 = ~n23625 & ~n23626;
  assign n23628 = ~n23624 & ~n23627;
  assign n23629 = ~n23286 & ~n23628;
  assign n23630 = ~n23262 & n23272;
  assign n23631 = ~n23273 & ~n23630;
  assign n23632 = ~n23629 & n23631;
  assign n23633 = ~n23273 & ~n23632;
  assign n23634 = n23256 & n23259;
  assign n23635 = ~n23260 & ~n23634;
  assign n23636 = ~n23633 & n23635;
  assign n23637 = ~n23260 & ~n23636;
  assign n23638 = ~n23246 & ~n23637;
  assign n23639 = ~n23243 & ~n23638;
  assign n23640 = n23217 & n23229;
  assign n23641 = ~n23217 & ~n23229;
  assign n23642 = ~n23640 & ~n23641;
  assign n23643 = ~n23639 & ~n23642;
  assign n23644 = ~n23230 & ~n23643;
  assign n23645 = n23202 & n23214;
  assign n23646 = ~n23202 & ~n23214;
  assign n23647 = ~n23645 & ~n23646;
  assign n23648 = ~n23644 & ~n23647;
  assign n23649 = ~n23215 & ~n23648;
  assign n23650 = n23187 & n23199;
  assign n23651 = ~n23187 & ~n23199;
  assign n23652 = ~n23650 & ~n23651;
  assign n23653 = ~n23649 & ~n23652;
  assign n23654 = ~n23200 & ~n23653;
  assign n23655 = ~n23182 & ~n23186;
  assign n23656 = n7430 & n21021;
  assign n23657 = n7431 & n23220;
  assign n23658 = n7869 & n21018;
  assign n23659 = n7895 & n21015;
  assign n23660 = ~n23656 & ~n23658;
  assign n23661 = ~n23659 & n23660;
  assign n23662 = ~n23657 & n23661;
  assign n23663 = ~pi11  & ~n23662;
  assign n23664 = pi11  & n23662;
  assign n23665 = ~n23663 & ~n23664;
  assign n23666 = n23165 & ~n23175;
  assign n23667 = ~n23044 & ~n23178;
  assign n23668 = ~n23666 & ~n23667;
  assign n23669 = n5982 & n21039;
  assign n23670 = n5983 & n22186;
  assign n23671 = n6323 & n21036;
  assign n23672 = n6336 & n21033;
  assign n23673 = ~n23669 & ~n23671;
  assign n23674 = ~n23672 & n23673;
  assign n23675 = ~n23670 & n23674;
  assign n23676 = ~pi17  & ~n23675;
  assign n23677 = pi17  & n23675;
  assign n23678 = ~n23676 & ~n23677;
  assign n23679 = n23142 & ~n23152;
  assign n23680 = ~n23156 & ~n23679;
  assign n23681 = ~n23137 & ~n23141;
  assign n23682 = n5044 & n21057;
  assign n23683 = n5045 & n21825;
  assign n23684 = n5109 & n21054;
  assign n23685 = n5130 & n21051;
  assign n23686 = ~n23682 & ~n23684;
  assign n23687 = ~n23685 & n23686;
  assign n23688 = ~n23683 & n23687;
  assign n23689 = ~pi23  & ~n23688;
  assign n23690 = pi23  & n23688;
  assign n23691 = ~n23689 & ~n23690;
  assign n23692 = n23120 & ~n23130;
  assign n23693 = ~n23071 & ~n23133;
  assign n23694 = ~n23692 & ~n23693;
  assign n23695 = n3810 & n21075;
  assign n23696 = n3886 & n21441;
  assign n23697 = n3884 & n21072;
  assign n23698 = n4380 & n21069;
  assign n23699 = ~n23695 & ~n23697;
  assign n23700 = ~n23698 & n23699;
  assign n23701 = ~n23696 & n23700;
  assign n23702 = ~pi29  & ~n23701;
  assign n23703 = pi29  & n23701;
  assign n23704 = ~n23702 & ~n23703;
  assign n23705 = ~n23098 & ~n23105;
  assign n23706 = ~n23111 & ~n23705;
  assign n23707 = ~n299 & ~n437;
  assign n23708 = ~n460 & ~n518;
  assign n23709 = ~n566 & ~n687;
  assign n23710 = n23708 & n23709;
  assign n23711 = n244 & n23707;
  assign n23712 = n4858 & n23711;
  assign n23713 = n1152 & n23710;
  assign n23714 = n1916 & n6170;
  assign n23715 = n23713 & n23714;
  assign n23716 = n12818 & n23712;
  assign n23717 = n23715 & n23716;
  assign n23718 = n12805 & n23717;
  assign n23719 = n20932 & n23718;
  assign n23720 = n14943 & n23719;
  assign n23721 = n3692 & n21081;
  assign n23722 = n880 & n21370;
  assign n23723 = n748 & n21084;
  assign n23724 = n3694 & n21078;
  assign n23725 = ~n23721 & ~n23723;
  assign n23726 = ~n23724 & n23725;
  assign n23727 = ~n23722 & n23726;
  assign n23728 = ~n23720 & n23727;
  assign n23729 = n23720 & ~n23727;
  assign n23730 = ~n23728 & ~n23729;
  assign n23731 = ~n23706 & ~n23730;
  assign n23732 = n23706 & n23730;
  assign n23733 = ~n23731 & ~n23732;
  assign n23734 = ~n23704 & ~n23733;
  assign n23735 = n23704 & n23733;
  assign n23736 = ~n23734 & ~n23735;
  assign n23737 = ~n23081 & n23113;
  assign n23738 = ~n23119 & ~n23737;
  assign n23739 = n23736 & n23738;
  assign n23740 = ~n23736 & ~n23738;
  assign n23741 = ~n23739 & ~n23740;
  assign n23742 = n86 & n21066;
  assign n23743 = n4420 & n21631;
  assign n23744 = n4600 & n21063;
  assign n23745 = n4615 & n21060;
  assign n23746 = ~n23742 & ~n23744;
  assign n23747 = ~n23745 & n23746;
  assign n23748 = ~n23743 & n23747;
  assign n23749 = pi26  & n23748;
  assign n23750 = ~pi26  & ~n23748;
  assign n23751 = ~n23749 & ~n23750;
  assign n23752 = n23741 & n23751;
  assign n23753 = ~n23741 & ~n23751;
  assign n23754 = ~n23752 & ~n23753;
  assign n23755 = ~n23694 & n23754;
  assign n23756 = n23694 & ~n23754;
  assign n23757 = ~n23755 & ~n23756;
  assign n23758 = ~n23691 & ~n23757;
  assign n23759 = n23691 & n23757;
  assign n23760 = ~n23758 & ~n23759;
  assign n23761 = n23681 & ~n23760;
  assign n23762 = ~n23681 & n23760;
  assign n23763 = ~n23761 & ~n23762;
  assign n23764 = n5240 & n21048;
  assign n23765 = n5241 & n22049;
  assign n23766 = n5853 & n21045;
  assign n23767 = n5866 & n21042;
  assign n23768 = ~n23764 & ~n23766;
  assign n23769 = ~n23767 & n23768;
  assign n23770 = ~n23765 & n23769;
  assign n23771 = pi20  & n23770;
  assign n23772 = ~pi20  & ~n23770;
  assign n23773 = ~n23771 & ~n23772;
  assign n23774 = n23763 & n23773;
  assign n23775 = ~n23763 & ~n23773;
  assign n23776 = ~n23774 & ~n23775;
  assign n23777 = ~n23680 & ~n23776;
  assign n23778 = n23680 & n23776;
  assign n23779 = ~n23777 & ~n23778;
  assign n23780 = ~n23678 & ~n23779;
  assign n23781 = n23678 & n23779;
  assign n23782 = ~n23780 & ~n23781;
  assign n23783 = ~n23054 & n23158;
  assign n23784 = ~n23164 & ~n23783;
  assign n23785 = n23782 & n23784;
  assign n23786 = ~n23782 & ~n23784;
  assign n23787 = ~n23785 & ~n23786;
  assign n23788 = n6630 & n21030;
  assign n23789 = n6631 & n22654;
  assign n23790 = n7238 & n21027;
  assign n23791 = n7262 & n21024;
  assign n23792 = ~n23788 & ~n23790;
  assign n23793 = ~n23791 & n23792;
  assign n23794 = ~n23789 & n23793;
  assign n23795 = pi14  & n23794;
  assign n23796 = ~pi14  & ~n23794;
  assign n23797 = ~n23795 & ~n23796;
  assign n23798 = n23787 & n23797;
  assign n23799 = ~n23787 & ~n23797;
  assign n23800 = ~n23798 & ~n23799;
  assign n23801 = ~n23668 & n23800;
  assign n23802 = n23668 & ~n23800;
  assign n23803 = ~n23801 & ~n23802;
  assign n23804 = ~n23665 & ~n23803;
  assign n23805 = n23665 & n23803;
  assign n23806 = ~n23804 & ~n23805;
  assign n23807 = n23655 & ~n23806;
  assign n23808 = ~n23655 & n23806;
  assign n23809 = ~n23807 & ~n23808;
  assign n23810 = n8250 & n21012;
  assign n23811 = n21191 & ~n21193;
  assign n23812 = ~n21194 & ~n23811;
  assign n23813 = n8251 & n23812;
  assign n23814 = n9016 & n21009;
  assign n23815 = n9040 & n21006;
  assign n23816 = ~n23810 & ~n23814;
  assign n23817 = ~n23815 & n23816;
  assign n23818 = ~n23813 & n23817;
  assign n23819 = pi8  & n23818;
  assign n23820 = ~pi8  & ~n23818;
  assign n23821 = ~n23819 & ~n23820;
  assign n23822 = n23809 & n23821;
  assign n23823 = ~n23809 & ~n23821;
  assign n23824 = ~n23822 & ~n23823;
  assign n23825 = ~n23654 & ~n23824;
  assign n23826 = n23654 & n23824;
  assign n23827 = ~n23825 & ~n23826;
  assign n23828 = ~n21303 & ~n23827;
  assign n23829 = n21303 & n23827;
  assign n23830 = ~n23828 & ~n23829;
  assign n23831 = n75 & n21006;
  assign n23832 = n21199 & ~n21201;
  assign n23833 = ~n21202 & ~n23832;
  assign n23834 = n9491 & n23833;
  assign n23835 = n10469 & n20906;
  assign n23836 = n11031 & n21003;
  assign n23837 = ~n23831 & ~n23835;
  assign n23838 = ~n23836 & n23837;
  assign n23839 = ~n23834 & n23838;
  assign n23840 = ~pi5  & ~n23839;
  assign n23841 = pi5  & n23839;
  assign n23842 = ~n23840 & ~n23841;
  assign n23843 = n23649 & n23652;
  assign n23844 = ~n23653 & ~n23843;
  assign n23845 = ~n23842 & n23844;
  assign n23846 = ~n23842 & ~n23844;
  assign n23847 = n23842 & n23844;
  assign n23848 = ~n23846 & ~n23847;
  assign n23849 = n75 & n21009;
  assign n23850 = n21195 & ~n21197;
  assign n23851 = ~n21198 & ~n23850;
  assign n23852 = n9491 & n23851;
  assign n23853 = n10469 & n21006;
  assign n23854 = n11031 & n20906;
  assign n23855 = ~n23849 & ~n23853;
  assign n23856 = ~n23854 & n23855;
  assign n23857 = ~n23852 & n23856;
  assign n23858 = ~pi5  & ~n23857;
  assign n23859 = pi5  & n23857;
  assign n23860 = ~n23858 & ~n23859;
  assign n23861 = ~n23644 & n23647;
  assign n23862 = n23644 & ~n23647;
  assign n23863 = ~n23861 & ~n23862;
  assign n23864 = ~n23860 & ~n23863;
  assign n23865 = n75 & n21012;
  assign n23866 = n9491 & n23812;
  assign n23867 = n10469 & n21009;
  assign n23868 = n11031 & n21006;
  assign n23869 = ~n23865 & ~n23867;
  assign n23870 = ~n23868 & n23869;
  assign n23871 = ~n23866 & n23870;
  assign n23872 = ~pi5  & ~n23871;
  assign n23873 = pi5  & n23871;
  assign n23874 = ~n23872 & ~n23873;
  assign n23875 = ~n23639 & n23642;
  assign n23876 = n23639 & ~n23642;
  assign n23877 = ~n23875 & ~n23876;
  assign n23878 = ~n23874 & ~n23877;
  assign n23879 = n23246 & n23637;
  assign n23880 = ~n23638 & ~n23879;
  assign n23881 = n75 & n21015;
  assign n23882 = n9491 & n23190;
  assign n23883 = n10469 & n21012;
  assign n23884 = n11031 & n21009;
  assign n23885 = ~n23881 & ~n23883;
  assign n23886 = ~n23884 & n23885;
  assign n23887 = ~n23882 & n23886;
  assign n23888 = pi5  & n23887;
  assign n23889 = ~pi5  & ~n23887;
  assign n23890 = ~n23888 & ~n23889;
  assign n23891 = n23880 & ~n23890;
  assign n23892 = n23633 & ~n23635;
  assign n23893 = ~n23636 & ~n23892;
  assign n23894 = n75 & n21018;
  assign n23895 = n9491 & n23205;
  assign n23896 = n10469 & n21015;
  assign n23897 = n11031 & n21012;
  assign n23898 = ~n23894 & ~n23896;
  assign n23899 = ~n23897 & n23898;
  assign n23900 = ~n23895 & n23899;
  assign n23901 = pi5  & n23900;
  assign n23902 = ~pi5  & ~n23900;
  assign n23903 = ~n23901 & ~n23902;
  assign n23904 = n23893 & ~n23903;
  assign n23905 = n75 & n21021;
  assign n23906 = n9491 & n23220;
  assign n23907 = n10469 & n21018;
  assign n23908 = n11031 & n21015;
  assign n23909 = ~n23905 & ~n23907;
  assign n23910 = ~n23908 & n23909;
  assign n23911 = ~n23906 & n23910;
  assign n23912 = ~pi5  & ~n23911;
  assign n23913 = pi5  & n23911;
  assign n23914 = ~n23912 & ~n23913;
  assign n23915 = n23629 & ~n23631;
  assign n23916 = ~n23632 & ~n23915;
  assign n23917 = ~n23914 & n23916;
  assign n23918 = ~n23914 & ~n23916;
  assign n23919 = n23914 & n23916;
  assign n23920 = ~n23918 & ~n23919;
  assign n23921 = n75 & n21024;
  assign n23922 = n9491 & n23033;
  assign n23923 = n10469 & n21021;
  assign n23924 = n11031 & n21018;
  assign n23925 = ~n23921 & ~n23923;
  assign n23926 = ~n23924 & n23925;
  assign n23927 = ~n23922 & n23926;
  assign n23928 = ~pi5  & ~n23927;
  assign n23929 = pi5  & n23927;
  assign n23930 = ~n23928 & ~n23929;
  assign n23931 = n23624 & n23627;
  assign n23932 = ~n23628 & ~n23931;
  assign n23933 = ~n23930 & n23932;
  assign n23934 = ~n23930 & ~n23932;
  assign n23935 = n23930 & n23932;
  assign n23936 = ~n23934 & ~n23935;
  assign n23937 = n75 & n21027;
  assign n23938 = n9491 & n21306;
  assign n23939 = n10469 & n21024;
  assign n23940 = n11031 & n21021;
  assign n23941 = ~n23937 & ~n23939;
  assign n23942 = ~n23940 & n23941;
  assign n23943 = ~n23938 & n23942;
  assign n23944 = ~pi5  & ~n23943;
  assign n23945 = pi5  & n23943;
  assign n23946 = ~n23944 & ~n23945;
  assign n23947 = ~n23619 & n23622;
  assign n23948 = n23619 & ~n23622;
  assign n23949 = ~n23947 & ~n23948;
  assign n23950 = ~n23946 & ~n23949;
  assign n23951 = n23315 & n23617;
  assign n23952 = ~n23618 & ~n23951;
  assign n23953 = n75 & n21030;
  assign n23954 = n9491 & n22654;
  assign n23955 = n10469 & n21027;
  assign n23956 = n11031 & n21024;
  assign n23957 = ~n23953 & ~n23955;
  assign n23958 = ~n23956 & n23957;
  assign n23959 = ~n23954 & n23958;
  assign n23960 = pi5  & n23959;
  assign n23961 = ~pi5  & ~n23959;
  assign n23962 = ~n23960 & ~n23961;
  assign n23963 = n23952 & ~n23962;
  assign n23964 = n23613 & ~n23615;
  assign n23965 = ~n23616 & ~n23964;
  assign n23966 = n75 & n21033;
  assign n23967 = n9491 & n22674;
  assign n23968 = n10469 & n21030;
  assign n23969 = n11031 & n21027;
  assign n23970 = ~n23966 & ~n23968;
  assign n23971 = ~n23969 & n23970;
  assign n23972 = ~n23967 & n23971;
  assign n23973 = pi5  & n23972;
  assign n23974 = ~pi5  & ~n23972;
  assign n23975 = ~n23973 & ~n23974;
  assign n23976 = n23965 & ~n23975;
  assign n23977 = n23345 & n23611;
  assign n23978 = ~n23612 & ~n23977;
  assign n23979 = n75 & n21036;
  assign n23980 = n9491 & n22632;
  assign n23981 = n10469 & n21033;
  assign n23982 = n11031 & n21030;
  assign n23983 = ~n23979 & ~n23981;
  assign n23984 = ~n23982 & n23983;
  assign n23985 = ~n23980 & n23984;
  assign n23986 = pi5  & n23985;
  assign n23987 = ~pi5  & ~n23985;
  assign n23988 = ~n23986 & ~n23987;
  assign n23989 = n23978 & ~n23988;
  assign n23990 = n75 & n21039;
  assign n23991 = n9491 & n22186;
  assign n23992 = n10469 & n21036;
  assign n23993 = n11031 & n21033;
  assign n23994 = ~n23990 & ~n23992;
  assign n23995 = ~n23993 & n23994;
  assign n23996 = ~n23991 & n23995;
  assign n23997 = ~pi5  & ~n23996;
  assign n23998 = pi5  & n23996;
  assign n23999 = ~n23997 & ~n23998;
  assign n24000 = n23607 & ~n23609;
  assign n24001 = ~n23610 & ~n24000;
  assign n24002 = ~n23999 & n24001;
  assign n24003 = ~n23999 & ~n24001;
  assign n24004 = n23999 & n24001;
  assign n24005 = ~n24003 & ~n24004;
  assign n24006 = n75 & n21042;
  assign n24007 = n9491 & n22199;
  assign n24008 = n10469 & n21039;
  assign n24009 = n11031 & n21036;
  assign n24010 = ~n24006 & ~n24008;
  assign n24011 = ~n24009 & n24010;
  assign n24012 = ~n24007 & n24011;
  assign n24013 = ~pi5  & ~n24012;
  assign n24014 = pi5  & n24012;
  assign n24015 = ~n24013 & ~n24014;
  assign n24016 = ~n23602 & n23605;
  assign n24017 = n23602 & ~n23605;
  assign n24018 = ~n24016 & ~n24017;
  assign n24019 = ~n24015 & ~n24018;
  assign n24020 = n75 & n21045;
  assign n24021 = n9491 & n22217;
  assign n24022 = n10469 & n21042;
  assign n24023 = n11031 & n21039;
  assign n24024 = ~n24020 & ~n24022;
  assign n24025 = ~n24023 & n24024;
  assign n24026 = ~n24021 & n24025;
  assign n24027 = ~pi5  & ~n24026;
  assign n24028 = pi5  & n24026;
  assign n24029 = ~n24027 & ~n24028;
  assign n24030 = n23597 & n23600;
  assign n24031 = ~n23601 & ~n24030;
  assign n24032 = ~n24029 & n24031;
  assign n24033 = ~n24029 & ~n24031;
  assign n24034 = n24029 & n24031;
  assign n24035 = ~n24033 & ~n24034;
  assign n24036 = n23400 & n23595;
  assign n24037 = ~n23596 & ~n24036;
  assign n24038 = n75 & n21048;
  assign n24039 = n9491 & n22049;
  assign n24040 = n10469 & n21045;
  assign n24041 = n11031 & n21042;
  assign n24042 = ~n24038 & ~n24040;
  assign n24043 = ~n24041 & n24042;
  assign n24044 = ~n24039 & n24043;
  assign n24045 = pi5  & n24044;
  assign n24046 = ~pi5  & ~n24044;
  assign n24047 = ~n24045 & ~n24046;
  assign n24048 = n24037 & ~n24047;
  assign n24049 = n23416 & n23593;
  assign n24050 = ~n23594 & ~n24049;
  assign n24051 = n75 & n21051;
  assign n24052 = n9491 & n21797;
  assign n24053 = n10469 & n21048;
  assign n24054 = n11031 & n21045;
  assign n24055 = ~n24051 & ~n24053;
  assign n24056 = ~n24054 & n24055;
  assign n24057 = ~n24052 & n24056;
  assign n24058 = pi5  & n24057;
  assign n24059 = ~pi5  & ~n24057;
  assign n24060 = ~n24058 & ~n24059;
  assign n24061 = n24050 & ~n24060;
  assign n24062 = n23589 & ~n23591;
  assign n24063 = ~n23592 & ~n24062;
  assign n24064 = n75 & n21054;
  assign n24065 = n9491 & n21812;
  assign n24066 = n10469 & n21051;
  assign n24067 = n11031 & n21048;
  assign n24068 = ~n24064 & ~n24066;
  assign n24069 = ~n24067 & n24068;
  assign n24070 = ~n24065 & n24069;
  assign n24071 = pi5  & n24070;
  assign n24072 = ~pi5  & ~n24070;
  assign n24073 = ~n24071 & ~n24072;
  assign n24074 = n24063 & ~n24073;
  assign n24075 = n75 & n21057;
  assign n24076 = n9491 & n21825;
  assign n24077 = n10469 & n21054;
  assign n24078 = n11031 & n21051;
  assign n24079 = ~n24075 & ~n24077;
  assign n24080 = ~n24078 & n24079;
  assign n24081 = ~n24076 & n24080;
  assign n24082 = ~pi5  & ~n24081;
  assign n24083 = pi5  & n24081;
  assign n24084 = ~n24082 & ~n24083;
  assign n24085 = n23585 & ~n23587;
  assign n24086 = ~n23588 & ~n24085;
  assign n24087 = ~n24084 & n24086;
  assign n24088 = ~n24084 & ~n24086;
  assign n24089 = n24084 & n24086;
  assign n24090 = ~n24088 & ~n24089;
  assign n24091 = n75 & n21060;
  assign n24092 = n9491 & n21318;
  assign n24093 = n10469 & n21057;
  assign n24094 = n11031 & n21054;
  assign n24095 = ~n24091 & ~n24093;
  assign n24096 = ~n24094 & n24095;
  assign n24097 = ~n24092 & n24096;
  assign n24098 = ~pi5  & ~n24097;
  assign n24099 = pi5  & n24097;
  assign n24100 = ~n24098 & ~n24099;
  assign n24101 = n23580 & n23583;
  assign n24102 = ~n23584 & ~n24101;
  assign n24103 = ~n24100 & n24102;
  assign n24104 = ~n24100 & ~n24102;
  assign n24105 = n24100 & n24102;
  assign n24106 = ~n24104 & ~n24105;
  assign n24107 = n75 & n21063;
  assign n24108 = n9491 & n21613;
  assign n24109 = n10469 & n21060;
  assign n24110 = n11031 & n21057;
  assign n24111 = ~n24107 & ~n24109;
  assign n24112 = ~n24110 & n24111;
  assign n24113 = ~n24108 & n24112;
  assign n24114 = ~pi5  & ~n24113;
  assign n24115 = pi5  & n24113;
  assign n24116 = ~n24114 & ~n24115;
  assign n24117 = ~n23575 & n23578;
  assign n24118 = n23575 & ~n23578;
  assign n24119 = ~n24117 & ~n24118;
  assign n24120 = ~n24116 & ~n24119;
  assign n24121 = n23485 & n23573;
  assign n24122 = ~n23574 & ~n24121;
  assign n24123 = n75 & n21066;
  assign n24124 = n9491 & n21631;
  assign n24125 = n10469 & n21063;
  assign n24126 = n11031 & n21060;
  assign n24127 = ~n24123 & ~n24125;
  assign n24128 = ~n24126 & n24127;
  assign n24129 = ~n24124 & n24128;
  assign n24130 = pi5  & n24129;
  assign n24131 = ~pi5  & ~n24129;
  assign n24132 = ~n24130 & ~n24131;
  assign n24133 = n24122 & ~n24132;
  assign n24134 = n23569 & ~n23571;
  assign n24135 = ~n23572 & ~n24134;
  assign n24136 = n75 & n21069;
  assign n24137 = n9491 & n21592;
  assign n24138 = n10469 & n21066;
  assign n24139 = n11031 & n21063;
  assign n24140 = ~n24136 & ~n24138;
  assign n24141 = ~n24139 & n24140;
  assign n24142 = ~n24137 & n24141;
  assign n24143 = pi5  & n24142;
  assign n24144 = ~pi5  & ~n24142;
  assign n24145 = ~n24143 & ~n24144;
  assign n24146 = n24135 & ~n24145;
  assign n24147 = n23516 & n23567;
  assign n24148 = ~n23568 & ~n24147;
  assign n24149 = n75 & n21072;
  assign n24150 = n9491 & n21428;
  assign n24151 = n10469 & n21069;
  assign n24152 = n11031 & n21066;
  assign n24153 = ~n24149 & ~n24151;
  assign n24154 = ~n24152 & n24153;
  assign n24155 = ~n24150 & n24154;
  assign n24156 = pi5  & n24155;
  assign n24157 = ~pi5  & ~n24155;
  assign n24158 = ~n24156 & ~n24157;
  assign n24159 = n24148 & ~n24158;
  assign n24160 = n75 & n21075;
  assign n24161 = n9491 & n21441;
  assign n24162 = n10469 & n21072;
  assign n24163 = n11031 & n21069;
  assign n24164 = ~n24160 & ~n24162;
  assign n24165 = ~n24163 & n24164;
  assign n24166 = ~n24161 & n24165;
  assign n24167 = ~pi5  & ~n24166;
  assign n24168 = pi5  & n24166;
  assign n24169 = ~n24167 & ~n24168;
  assign n24170 = n23563 & ~n23565;
  assign n24171 = ~n23566 & ~n24170;
  assign n24172 = ~n24169 & n24171;
  assign n24173 = ~n24169 & ~n24171;
  assign n24174 = n24169 & n24171;
  assign n24175 = ~n24173 & ~n24174;
  assign n24176 = n75 & n21078;
  assign n24177 = n9491 & n21459;
  assign n24178 = n10469 & n21075;
  assign n24179 = n11031 & n21072;
  assign n24180 = ~n24176 & ~n24178;
  assign n24181 = ~n24179 & n24180;
  assign n24182 = ~n24177 & n24181;
  assign n24183 = pi5  & n24182;
  assign n24184 = ~pi5  & ~n24182;
  assign n24185 = ~n24183 & ~n24184;
  assign n24186 = n23551 & n23561;
  assign n24187 = ~n23562 & ~n24186;
  assign n24188 = ~n24185 & n24187;
  assign n24189 = n75 & n21081;
  assign n24190 = n9491 & n21330;
  assign n24191 = n10469 & n21078;
  assign n24192 = n11031 & n21075;
  assign n24193 = ~n24189 & ~n24191;
  assign n24194 = ~n24192 & n24193;
  assign n24195 = ~n24190 & n24194;
  assign n24196 = ~pi5  & ~n24195;
  assign n24197 = pi5  & n24195;
  assign n24198 = ~n24196 & ~n24197;
  assign n24199 = pi8  & ~n23539;
  assign n24200 = n23546 & ~n24199;
  assign n24201 = ~n23546 & n24199;
  assign n24202 = ~n24200 & ~n24201;
  assign n24203 = ~n24198 & n24202;
  assign n24204 = ~n24198 & ~n24202;
  assign n24205 = n24198 & n24202;
  assign n24206 = ~n24204 & ~n24205;
  assign n24207 = n75 & n21084;
  assign n24208 = n9491 & n21370;
  assign n24209 = n10469 & n21081;
  assign n24210 = n11031 & n21078;
  assign n24211 = ~n24207 & ~n24209;
  assign n24212 = ~n24210 & n24211;
  assign n24213 = ~n24208 & n24212;
  assign n24214 = pi5  & n24213;
  assign n24215 = ~pi5  & ~n24213;
  assign n24216 = ~n24214 & ~n24215;
  assign n24217 = pi8  & n23532;
  assign n24218 = ~n23537 & n24217;
  assign n24219 = n23537 & ~n24217;
  assign n24220 = ~n24218 & ~n24219;
  assign n24221 = ~n24216 & n24220;
  assign n24222 = ~n70 & n21091;
  assign n24223 = n10469 & n21091;
  assign n24224 = n11031 & n21089;
  assign n24225 = n9491 & ~n21345;
  assign n24226 = ~n24223 & ~n24224;
  assign n24227 = ~n24225 & n24226;
  assign n24228 = pi5  & ~n24222;
  assign n24229 = n24227 & n24228;
  assign n24230 = n75 & n21091;
  assign n24231 = n9491 & ~n21355;
  assign n24232 = n10469 & n21089;
  assign n24233 = n11031 & n21084;
  assign n24234 = ~n24230 & ~n24232;
  assign n24235 = ~n24233 & n24234;
  assign n24236 = ~n24231 & n24235;
  assign n24237 = n24229 & n24236;
  assign n24238 = n23532 & n24237;
  assign n24239 = ~n23532 & n24237;
  assign n24240 = n23532 & ~n24237;
  assign n24241 = ~n24239 & ~n24240;
  assign n24242 = n75 & n21089;
  assign n24243 = n9491 & n21407;
  assign n24244 = n10469 & n21084;
  assign n24245 = n11031 & n21081;
  assign n24246 = ~n24242 & ~n24244;
  assign n24247 = ~n24245 & n24246;
  assign n24248 = ~n24243 & n24247;
  assign n24249 = pi5  & n24248;
  assign n24250 = ~pi5  & ~n24248;
  assign n24251 = ~n24249 & ~n24250;
  assign n24252 = ~n24241 & ~n24251;
  assign n24253 = ~n24238 & ~n24252;
  assign n24254 = n24216 & ~n24220;
  assign n24255 = ~n24221 & ~n24254;
  assign n24256 = ~n24253 & n24255;
  assign n24257 = ~n24221 & ~n24256;
  assign n24258 = ~n24206 & ~n24257;
  assign n24259 = ~n24203 & ~n24258;
  assign n24260 = n24185 & ~n24187;
  assign n24261 = ~n24188 & ~n24260;
  assign n24262 = ~n24259 & n24261;
  assign n24263 = ~n24188 & ~n24262;
  assign n24264 = ~n24175 & ~n24263;
  assign n24265 = ~n24172 & ~n24264;
  assign n24266 = n24148 & n24158;
  assign n24267 = ~n24148 & ~n24158;
  assign n24268 = ~n24266 & ~n24267;
  assign n24269 = ~n24265 & ~n24268;
  assign n24270 = ~n24159 & ~n24269;
  assign n24271 = n24135 & n24145;
  assign n24272 = ~n24135 & ~n24145;
  assign n24273 = ~n24271 & ~n24272;
  assign n24274 = ~n24270 & ~n24273;
  assign n24275 = ~n24146 & ~n24274;
  assign n24276 = ~n24122 & n24132;
  assign n24277 = ~n24133 & ~n24276;
  assign n24278 = ~n24275 & n24277;
  assign n24279 = ~n24133 & ~n24278;
  assign n24280 = n24116 & n24119;
  assign n24281 = ~n24120 & ~n24280;
  assign n24282 = ~n24279 & n24281;
  assign n24283 = ~n24120 & ~n24282;
  assign n24284 = ~n24106 & ~n24283;
  assign n24285 = ~n24103 & ~n24284;
  assign n24286 = ~n24090 & ~n24285;
  assign n24287 = ~n24087 & ~n24286;
  assign n24288 = n24063 & n24073;
  assign n24289 = ~n24063 & ~n24073;
  assign n24290 = ~n24288 & ~n24289;
  assign n24291 = ~n24287 & ~n24290;
  assign n24292 = ~n24074 & ~n24291;
  assign n24293 = n24050 & n24060;
  assign n24294 = ~n24050 & ~n24060;
  assign n24295 = ~n24293 & ~n24294;
  assign n24296 = ~n24292 & ~n24295;
  assign n24297 = ~n24061 & ~n24296;
  assign n24298 = ~n24037 & n24047;
  assign n24299 = ~n24048 & ~n24298;
  assign n24300 = ~n24297 & n24299;
  assign n24301 = ~n24048 & ~n24300;
  assign n24302 = ~n24035 & ~n24301;
  assign n24303 = ~n24032 & ~n24302;
  assign n24304 = n24015 & n24018;
  assign n24305 = ~n24019 & ~n24304;
  assign n24306 = ~n24303 & n24305;
  assign n24307 = ~n24019 & ~n24306;
  assign n24308 = ~n24005 & ~n24307;
  assign n24309 = ~n24002 & ~n24308;
  assign n24310 = n23978 & n23988;
  assign n24311 = ~n23978 & ~n23988;
  assign n24312 = ~n24310 & ~n24311;
  assign n24313 = ~n24309 & ~n24312;
  assign n24314 = ~n23989 & ~n24313;
  assign n24315 = n23965 & n23975;
  assign n24316 = ~n23965 & ~n23975;
  assign n24317 = ~n24315 & ~n24316;
  assign n24318 = ~n24314 & ~n24317;
  assign n24319 = ~n23976 & ~n24318;
  assign n24320 = ~n23952 & n23962;
  assign n24321 = ~n23963 & ~n24320;
  assign n24322 = ~n24319 & n24321;
  assign n24323 = ~n23963 & ~n24322;
  assign n24324 = n23946 & n23949;
  assign n24325 = ~n23950 & ~n24324;
  assign n24326 = ~n24323 & n24325;
  assign n24327 = ~n23950 & ~n24326;
  assign n24328 = ~n23936 & ~n24327;
  assign n24329 = ~n23933 & ~n24328;
  assign n24330 = ~n23920 & ~n24329;
  assign n24331 = ~n23917 & ~n24330;
  assign n24332 = n23893 & n23903;
  assign n24333 = ~n23893 & ~n23903;
  assign n24334 = ~n24332 & ~n24333;
  assign n24335 = ~n24331 & ~n24334;
  assign n24336 = ~n23904 & ~n24335;
  assign n24337 = ~n23880 & n23890;
  assign n24338 = ~n23891 & ~n24337;
  assign n24339 = ~n24336 & n24338;
  assign n24340 = ~n23891 & ~n24339;
  assign n24341 = n23874 & n23877;
  assign n24342 = ~n23878 & ~n24341;
  assign n24343 = ~n24340 & n24342;
  assign n24344 = ~n23878 & ~n24343;
  assign n24345 = n23860 & n23863;
  assign n24346 = ~n23864 & ~n24345;
  assign n24347 = ~n24344 & n24346;
  assign n24348 = ~n23864 & ~n24347;
  assign n24349 = ~n23848 & ~n24348;
  assign n24350 = ~n23845 & ~n24349;
  assign n24351 = n23830 & n24350;
  assign n24352 = ~n23830 & ~n24350;
  assign n24353 = ~n24351 & ~n24352;
  assign n24354 = ~n21283 & ~n21286;
  assign n24355 = ~n21244 & ~n21246;
  assign n24356 = ~n106 & ~n355;
  assign n24357 = ~n361 & ~n703;
  assign n24358 = n24356 & n24357;
  assign n24359 = n1752 & n24358;
  assign n24360 = n943 & n7060;
  assign n24361 = n24359 & n24360;
  assign n24362 = ~n120 & ~n312;
  assign n24363 = ~n634 & n24362;
  assign n24364 = n797 & n1229;
  assign n24365 = n1245 & n3016;
  assign n24366 = n24364 & n24365;
  assign n24367 = n24363 & n24366;
  assign n24368 = n776 & n24367;
  assign n24369 = n24361 & n24368;
  assign n24370 = n12316 & n24369;
  assign n24371 = n1073 & n24370;
  assign n24372 = ~n24355 & n24371;
  assign n24373 = n24355 & ~n24371;
  assign n24374 = ~n24372 & ~n24373;
  assign n24375 = n3692 & n12395;
  assign n24376 = n880 & n13245;
  assign n24377 = n748 & n12398;
  assign n24378 = n3694 & n12362;
  assign n24379 = ~n24375 & ~n24377;
  assign n24380 = ~n24378 & n24379;
  assign n24381 = ~n24376 & n24380;
  assign n24382 = n24374 & ~n24381;
  assign n24383 = ~n24374 & n24381;
  assign n24384 = ~n24382 & ~n24383;
  assign n24385 = ~n21249 & n21258;
  assign n24386 = ~n21250 & ~n24385;
  assign n24387 = n24384 & n24386;
  assign n24388 = ~n24384 & ~n24386;
  assign n24389 = ~n24387 & ~n24388;
  assign n24390 = n3810 & n12392;
  assign n24391 = n3886 & n13421;
  assign n24392 = n3884 & n12646;
  assign n24393 = n4380 & n13164;
  assign n24394 = ~n24390 & ~n24392;
  assign n24395 = ~n24393 & n24394;
  assign n24396 = ~n24391 & n24395;
  assign n24397 = pi29  & n24396;
  assign n24398 = ~pi29  & ~n24396;
  assign n24399 = ~n24397 & ~n24398;
  assign n24400 = n24389 & ~n24399;
  assign n24401 = ~n24389 & n24399;
  assign n24402 = ~n24400 & ~n24401;
  assign n24403 = ~n21263 & n21274;
  assign n24404 = ~n21262 & ~n24403;
  assign n24405 = n24402 & n24404;
  assign n24406 = ~n24402 & ~n24404;
  assign n24407 = ~n24405 & ~n24406;
  assign n24408 = n4615 & ~n12786;
  assign n24409 = n4420 & ~n13781;
  assign n24410 = n86 & n13166;
  assign n24411 = n4600 & n13161;
  assign n24412 = ~n24408 & ~n24410;
  assign n24413 = ~n24411 & n24412;
  assign n24414 = ~n24409 & n24413;
  assign n24415 = pi26  & n24414;
  assign n24416 = ~pi26  & ~n24414;
  assign n24417 = ~n24415 & ~n24416;
  assign n24418 = n24407 & n24417;
  assign n24419 = ~n24407 & ~n24417;
  assign n24420 = ~n24418 & ~n24419;
  assign n24421 = ~n21214 & n21216;
  assign n24422 = ~n21278 & ~n24421;
  assign n24423 = ~n24420 & ~n24422;
  assign n24424 = n24420 & n24422;
  assign n24425 = ~n24423 & ~n24424;
  assign n24426 = ~n24354 & n24425;
  assign n24427 = n24354 & ~n24425;
  assign n24428 = ~n24426 & ~n24427;
  assign n24429 = n11055 & n24428;
  assign n24430 = ~n24423 & ~n24426;
  assign n24431 = ~n24372 & ~n24382;
  assign n24432 = ~n634 & ~n937;
  assign n24433 = n905 & n24432;
  assign n24434 = n2934 & n6171;
  assign n24435 = n24433 & n24434;
  assign n24436 = n1574 & n1985;
  assign n24437 = n24435 & n24436;
  assign n24438 = n921 & n24437;
  assign n24439 = n3625 & n24438;
  assign n24440 = n12316 & n24439;
  assign n24441 = n866 & n24440;
  assign n24442 = ~n24371 & n24441;
  assign n24443 = n24371 & ~n24441;
  assign n24444 = ~n24442 & ~n24443;
  assign n24445 = n748 & n12395;
  assign n24446 = n880 & n13144;
  assign n24447 = n3692 & n12362;
  assign n24448 = n3694 & n12392;
  assign n24449 = ~n24445 & ~n24447;
  assign n24450 = ~n24448 & n24449;
  assign n24451 = ~n24446 & n24450;
  assign n24452 = n24444 & ~n24451;
  assign n24453 = ~n24444 & n24451;
  assign n24454 = ~n24452 & ~n24453;
  assign n24455 = n24431 & ~n24454;
  assign n24456 = ~n24431 & n24454;
  assign n24457 = ~n24455 & ~n24456;
  assign n24458 = ~n24387 & ~n24400;
  assign n24459 = ~n24457 & n24458;
  assign n24460 = n24457 & ~n24458;
  assign n24461 = ~n24459 & ~n24460;
  assign n24462 = n4420 & ~n13280;
  assign n24463 = n86 & ~n13160;
  assign n24464 = ~n4600 & ~n4615;
  assign n24465 = ~n24463 & n24464;
  assign n24466 = ~n12786 & ~n24465;
  assign n24467 = ~n24462 & ~n24466;
  assign n24468 = ~pi26  & ~n24467;
  assign n24469 = pi26  & n24467;
  assign n24470 = ~n24468 & ~n24469;
  assign n24471 = n3810 & n12646;
  assign n24472 = n3886 & n13261;
  assign n24473 = n3884 & n13164;
  assign n24474 = n4380 & n13166;
  assign n24475 = ~n24471 & ~n24473;
  assign n24476 = ~n24474 & n24475;
  assign n24477 = ~n24472 & n24476;
  assign n24478 = pi29  & n24477;
  assign n24479 = ~pi29  & ~n24477;
  assign n24480 = ~n24478 & ~n24479;
  assign n24481 = ~n24470 & n24480;
  assign n24482 = n24470 & ~n24480;
  assign n24483 = ~n24481 & ~n24482;
  assign n24484 = ~n24461 & n24483;
  assign n24485 = n24461 & ~n24483;
  assign n24486 = ~n24484 & ~n24485;
  assign n24487 = ~n24406 & ~n24417;
  assign n24488 = ~n24405 & ~n24487;
  assign n24489 = n24486 & ~n24488;
  assign n24490 = ~n24486 & n24488;
  assign n24491 = ~n24489 & ~n24490;
  assign n24492 = ~n24430 & n24491;
  assign n24493 = n24430 & ~n24491;
  assign n24494 = ~n24492 & ~n24493;
  assign n24495 = n24428 & n24494;
  assign n24496 = n21288 & n24428;
  assign n24497 = ~n21289 & ~n21292;
  assign n24498 = ~n21288 & ~n24428;
  assign n24499 = ~n24496 & ~n24498;
  assign n24500 = ~n24497 & n24499;
  assign n24501 = ~n24496 & ~n24500;
  assign n24502 = ~n24428 & ~n24494;
  assign n24503 = ~n24495 & ~n24502;
  assign n24504 = ~n24501 & n24503;
  assign n24505 = ~n24495 & ~n24504;
  assign n24506 = ~n24489 & ~n24492;
  assign n24507 = ~n24456 & ~n24460;
  assign n24508 = n4380 & n13161;
  assign n24509 = n3886 & n13183;
  assign n24510 = n3884 & n13166;
  assign n24511 = n3810 & n13164;
  assign n24512 = ~n24510 & ~n24511;
  assign n24513 = ~n24508 & n24512;
  assign n24514 = ~n24509 & n24513;
  assign n24515 = pi29  & n24514;
  assign n24516 = ~pi29  & ~n24514;
  assign n24517 = ~n24515 & ~n24516;
  assign n24518 = ~n24443 & ~n24452;
  assign n24519 = n78 & n85;
  assign n24520 = ~n12786 & ~n24519;
  assign n24521 = pi26  & ~n24520;
  assign n24522 = ~pi26  & n24520;
  assign n24523 = ~n24521 & ~n24522;
  assign n24524 = n3851 & n3857;
  assign n24525 = ~n183 & ~n304;
  assign n24526 = n447 & n24525;
  assign n24527 = n3614 & n24526;
  assign n24528 = n3660 & n24527;
  assign n24529 = n24524 & n24528;
  assign n24530 = n24371 & n24529;
  assign n24531 = ~n24371 & ~n24529;
  assign n24532 = ~n24530 & ~n24531;
  assign n24533 = n24523 & n24532;
  assign n24534 = ~n24523 & ~n24532;
  assign n24535 = ~n24533 & ~n24534;
  assign n24536 = ~n24518 & n24535;
  assign n24537 = n24518 & ~n24535;
  assign n24538 = ~n24536 & ~n24537;
  assign n24539 = n748 & n12362;
  assign n24540 = n880 & n12652;
  assign n24541 = n3692 & n12392;
  assign n24542 = n3694 & n12646;
  assign n24543 = ~n24539 & ~n24541;
  assign n24544 = ~n24542 & n24543;
  assign n24545 = ~n24540 & n24544;
  assign n24546 = n24538 & ~n24545;
  assign n24547 = ~n24538 & n24545;
  assign n24548 = ~n24546 & ~n24547;
  assign n24549 = ~n24517 & n24548;
  assign n24550 = n24517 & ~n24548;
  assign n24551 = ~n24549 & ~n24550;
  assign n24552 = n24507 & ~n24551;
  assign n24553 = ~n24507 & n24551;
  assign n24554 = ~n24552 & ~n24553;
  assign n24555 = ~n24470 & ~n24480;
  assign n24556 = ~n24485 & ~n24555;
  assign n24557 = n24554 & ~n24556;
  assign n24558 = ~n24554 & n24556;
  assign n24559 = ~n24557 & ~n24558;
  assign n24560 = n24506 & ~n24559;
  assign n24561 = ~n24506 & n24559;
  assign n24562 = ~n24560 & ~n24561;
  assign n24563 = n24494 & n24562;
  assign n24564 = ~n24494 & ~n24562;
  assign n24565 = ~n24563 & ~n24564;
  assign n24566 = ~n24505 & n24565;
  assign n24567 = n24505 & ~n24565;
  assign n24568 = ~n24566 & ~n24567;
  assign n24569 = n11056 & n24568;
  assign n24570 = n11661 & n24494;
  assign n24571 = n11672 & n24562;
  assign n24572 = ~n24429 & ~n24570;
  assign n24573 = ~n24571 & n24572;
  assign n24574 = ~n24569 & n24573;
  assign n24575 = pi2  & n24574;
  assign n24576 = ~pi2  & ~n24574;
  assign n24577 = ~n24575 & ~n24576;
  assign n24578 = n24353 & ~n24577;
  assign n24579 = n24353 & n24577;
  assign n24580 = ~n24353 & ~n24577;
  assign n24581 = ~n24579 & ~n24580;
  assign n24582 = n11055 & n21288;
  assign n24583 = n24501 & ~n24503;
  assign n24584 = ~n24504 & ~n24583;
  assign n24585 = n11056 & n24584;
  assign n24586 = n11661 & n24428;
  assign n24587 = n11672 & n24494;
  assign n24588 = ~n24582 & ~n24586;
  assign n24589 = ~n24587 & n24588;
  assign n24590 = ~n24585 & n24589;
  assign n24591 = pi2  & n24590;
  assign n24592 = ~pi2  & ~n24590;
  assign n24593 = ~n24591 & ~n24592;
  assign n24594 = n11055 & n21003;
  assign n24595 = n24497 & ~n24499;
  assign n24596 = ~n24500 & ~n24595;
  assign n24597 = n11056 & n24596;
  assign n24598 = n11661 & n21288;
  assign n24599 = n11672 & n24428;
  assign n24600 = ~n24594 & ~n24598;
  assign n24601 = ~n24599 & n24600;
  assign n24602 = ~n24597 & n24601;
  assign n24603 = pi2  & n24602;
  assign n24604 = ~pi2  & ~n24602;
  assign n24605 = ~n24603 & ~n24604;
  assign n24606 = n11055 & n20906;
  assign n24607 = n11056 & n21294;
  assign n24608 = n11661 & n21003;
  assign n24609 = n11672 & n21288;
  assign n24610 = ~n24606 & ~n24608;
  assign n24611 = ~n24609 & n24610;
  assign n24612 = ~n24607 & n24611;
  assign n24613 = pi2  & n24612;
  assign n24614 = ~pi2  & ~n24612;
  assign n24615 = ~n24613 & ~n24614;
  assign n24616 = n24336 & ~n24338;
  assign n24617 = ~n24339 & ~n24616;
  assign n24618 = n24331 & n24334;
  assign n24619 = ~n24335 & ~n24618;
  assign n24620 = n11055 & n21012;
  assign n24621 = n11056 & n23812;
  assign n24622 = n11661 & n21009;
  assign n24623 = n11672 & n21006;
  assign n24624 = ~n24620 & ~n24622;
  assign n24625 = ~n24623 & n24624;
  assign n24626 = ~n24621 & n24625;
  assign n24627 = pi2  & n24626;
  assign n24628 = ~pi2  & ~n24626;
  assign n24629 = ~n24627 & ~n24628;
  assign n24630 = n11055 & n21015;
  assign n24631 = n11056 & n23190;
  assign n24632 = n11661 & n21012;
  assign n24633 = n11672 & n21009;
  assign n24634 = ~n24630 & ~n24632;
  assign n24635 = ~n24633 & n24634;
  assign n24636 = ~n24631 & n24635;
  assign n24637 = pi2  & n24636;
  assign n24638 = ~pi2  & ~n24636;
  assign n24639 = ~n24637 & ~n24638;
  assign n24640 = n11055 & n21018;
  assign n24641 = n11056 & n23205;
  assign n24642 = n11661 & n21015;
  assign n24643 = n11672 & n21012;
  assign n24644 = ~n24640 & ~n24642;
  assign n24645 = ~n24643 & n24644;
  assign n24646 = ~n24641 & n24645;
  assign n24647 = pi2  & n24646;
  assign n24648 = ~pi2  & ~n24646;
  assign n24649 = ~n24647 & ~n24648;
  assign n24650 = n24319 & ~n24321;
  assign n24651 = ~n24322 & ~n24650;
  assign n24652 = n24314 & n24317;
  assign n24653 = ~n24318 & ~n24652;
  assign n24654 = n24309 & n24312;
  assign n24655 = ~n24313 & ~n24654;
  assign n24656 = n11055 & n21030;
  assign n24657 = n11056 & n22654;
  assign n24658 = n11661 & n21027;
  assign n24659 = n11672 & n21024;
  assign n24660 = ~n24656 & ~n24658;
  assign n24661 = ~n24659 & n24660;
  assign n24662 = ~n24657 & n24661;
  assign n24663 = pi2  & n24662;
  assign n24664 = ~pi2  & ~n24662;
  assign n24665 = ~n24663 & ~n24664;
  assign n24666 = n11055 & n21033;
  assign n24667 = n11056 & n22674;
  assign n24668 = n11661 & n21030;
  assign n24669 = n11672 & n21027;
  assign n24670 = ~n24666 & ~n24668;
  assign n24671 = ~n24669 & n24670;
  assign n24672 = ~n24667 & n24671;
  assign n24673 = pi2  & n24672;
  assign n24674 = ~pi2  & ~n24672;
  assign n24675 = ~n24673 & ~n24674;
  assign n24676 = n11055 & n21036;
  assign n24677 = n11056 & n22632;
  assign n24678 = n11661 & n21033;
  assign n24679 = n11672 & n21030;
  assign n24680 = ~n24676 & ~n24678;
  assign n24681 = ~n24679 & n24680;
  assign n24682 = ~n24677 & n24681;
  assign n24683 = pi2  & n24682;
  assign n24684 = ~pi2  & ~n24682;
  assign n24685 = ~n24683 & ~n24684;
  assign n24686 = n24297 & ~n24299;
  assign n24687 = ~n24300 & ~n24686;
  assign n24688 = n24292 & n24295;
  assign n24689 = ~n24296 & ~n24688;
  assign n24690 = n24287 & n24290;
  assign n24691 = ~n24291 & ~n24690;
  assign n24692 = n11055 & n21048;
  assign n24693 = n11056 & n22049;
  assign n24694 = n11661 & n21045;
  assign n24695 = n11672 & n21042;
  assign n24696 = ~n24692 & ~n24694;
  assign n24697 = ~n24695 & n24696;
  assign n24698 = ~n24693 & n24697;
  assign n24699 = pi2  & n24698;
  assign n24700 = ~pi2  & ~n24698;
  assign n24701 = ~n24699 & ~n24700;
  assign n24702 = n11055 & n21051;
  assign n24703 = n11056 & n21797;
  assign n24704 = n11661 & n21048;
  assign n24705 = n11672 & n21045;
  assign n24706 = ~n24702 & ~n24704;
  assign n24707 = ~n24705 & n24706;
  assign n24708 = ~n24703 & n24707;
  assign n24709 = pi2  & n24708;
  assign n24710 = ~pi2  & ~n24708;
  assign n24711 = ~n24709 & ~n24710;
  assign n24712 = n11055 & n21054;
  assign n24713 = n11056 & n21812;
  assign n24714 = n11661 & n21051;
  assign n24715 = n11672 & n21048;
  assign n24716 = ~n24712 & ~n24714;
  assign n24717 = ~n24715 & n24716;
  assign n24718 = ~n24713 & n24717;
  assign n24719 = pi2  & n24718;
  assign n24720 = ~pi2  & ~n24718;
  assign n24721 = ~n24719 & ~n24720;
  assign n24722 = n24275 & ~n24277;
  assign n24723 = ~n24278 & ~n24722;
  assign n24724 = n24270 & n24273;
  assign n24725 = ~n24274 & ~n24724;
  assign n24726 = n24265 & n24268;
  assign n24727 = ~n24269 & ~n24726;
  assign n24728 = n11055 & n21066;
  assign n24729 = n11056 & n21631;
  assign n24730 = n11661 & n21063;
  assign n24731 = n11672 & n21060;
  assign n24732 = ~n24728 & ~n24730;
  assign n24733 = ~n24731 & n24732;
  assign n24734 = ~n24729 & n24733;
  assign n24735 = pi2  & n24734;
  assign n24736 = ~pi2  & ~n24734;
  assign n24737 = ~n24735 & ~n24736;
  assign n24738 = n11055 & n21069;
  assign n24739 = n11056 & n21592;
  assign n24740 = n11661 & n21066;
  assign n24741 = n11672 & n21063;
  assign n24742 = ~n24738 & ~n24740;
  assign n24743 = ~n24741 & n24742;
  assign n24744 = ~n24739 & n24743;
  assign n24745 = pi2  & n24744;
  assign n24746 = ~pi2  & ~n24744;
  assign n24747 = ~n24745 & ~n24746;
  assign n24748 = n11055 & n21072;
  assign n24749 = n11056 & n21428;
  assign n24750 = n11661 & n21069;
  assign n24751 = n11672 & n21066;
  assign n24752 = ~n24748 & ~n24750;
  assign n24753 = ~n24751 & n24752;
  assign n24754 = ~n24749 & n24753;
  assign n24755 = pi2  & n24754;
  assign n24756 = ~pi2  & ~n24754;
  assign n24757 = ~n24755 & ~n24756;
  assign n24758 = n24253 & ~n24255;
  assign n24759 = ~n24256 & ~n24758;
  assign n24760 = n11055 & n21078;
  assign n24761 = n11056 & n21459;
  assign n24762 = n11661 & n21075;
  assign n24763 = n11672 & n21072;
  assign n24764 = ~n24760 & ~n24762;
  assign n24765 = ~n24763 & n24764;
  assign n24766 = ~n24761 & n24765;
  assign n24767 = pi2  & n24766;
  assign n24768 = ~pi2  & ~n24766;
  assign n24769 = ~n24767 & ~n24768;
  assign n24770 = pi5  & ~n24229;
  assign n24771 = n24236 & ~n24770;
  assign n24772 = ~n24236 & n24770;
  assign n24773 = ~n24771 & ~n24772;
  assign n24774 = n11055 & n21084;
  assign n24775 = n11056 & n21370;
  assign n24776 = n11661 & n21081;
  assign n24777 = n11672 & n21078;
  assign n24778 = ~n24774 & ~n24776;
  assign n24779 = ~n24777 & n24778;
  assign n24780 = ~n24775 & n24779;
  assign n24781 = pi2  & n24780;
  assign n24782 = ~pi2  & ~n24780;
  assign n24783 = ~n24781 & ~n24782;
  assign n24784 = ~n11054 & n21091;
  assign n24785 = n11055 & n21091;
  assign n24786 = n11661 & n21089;
  assign n24787 = n11672 & n21084;
  assign n24788 = ~n24785 & ~n24786;
  assign n24789 = ~n24787 & n24788;
  assign n24790 = pi2  & ~n24789;
  assign n24791 = ~n21084 & n21345;
  assign n24792 = n11911 & ~n24791;
  assign n24793 = n20457 & n21089;
  assign n24794 = pi2  & ~n24784;
  assign n24795 = ~n24793 & n24794;
  assign n24796 = ~n24792 & n24795;
  assign n24797 = ~n24790 & n24796;
  assign n24798 = ~n24222 & ~n24797;
  assign n24799 = n24222 & n24797;
  assign n24800 = n11055 & n21089;
  assign n24801 = n11056 & n21407;
  assign n24802 = n11661 & n21084;
  assign n24803 = n11672 & n21081;
  assign n24804 = ~n24800 & ~n24802;
  assign n24805 = ~n24803 & n24804;
  assign n24806 = ~n24801 & n24805;
  assign n24807 = pi2  & ~n24806;
  assign n24808 = ~pi2  & n24806;
  assign n24809 = ~n24807 & ~n24808;
  assign n24810 = ~n24799 & ~n24809;
  assign n24811 = ~n24798 & ~n24810;
  assign n24812 = ~n24783 & n24811;
  assign n24813 = n24783 & ~n24811;
  assign n24814 = pi5  & n24222;
  assign n24815 = ~n24227 & n24814;
  assign n24816 = n24227 & ~n24814;
  assign n24817 = ~n24815 & ~n24816;
  assign n24818 = ~n24813 & n24817;
  assign n24819 = ~n24812 & ~n24818;
  assign n24820 = n24773 & ~n24819;
  assign n24821 = ~n24773 & n24819;
  assign n24822 = n11055 & n21081;
  assign n24823 = n11056 & n21330;
  assign n24824 = n11661 & n21078;
  assign n24825 = n11672 & n21075;
  assign n24826 = ~n24822 & ~n24824;
  assign n24827 = ~n24825 & n24826;
  assign n24828 = ~n24823 & n24827;
  assign n24829 = pi2  & ~n24828;
  assign n24830 = ~pi2  & n24828;
  assign n24831 = ~n24829 & ~n24830;
  assign n24832 = ~n24821 & n24831;
  assign n24833 = ~n24820 & ~n24832;
  assign n24834 = ~n24769 & ~n24833;
  assign n24835 = n24769 & n24833;
  assign n24836 = n24241 & n24251;
  assign n24837 = ~n24252 & ~n24836;
  assign n24838 = ~n24835 & n24837;
  assign n24839 = ~n24834 & ~n24838;
  assign n24840 = n24759 & ~n24839;
  assign n24841 = ~n24759 & n24839;
  assign n24842 = n11055 & n21075;
  assign n24843 = n11056 & n21441;
  assign n24844 = n11661 & n21072;
  assign n24845 = n11672 & n21069;
  assign n24846 = ~n24842 & ~n24844;
  assign n24847 = ~n24845 & n24846;
  assign n24848 = ~n24843 & n24847;
  assign n24849 = pi2  & ~n24848;
  assign n24850 = ~pi2  & n24848;
  assign n24851 = ~n24849 & ~n24850;
  assign n24852 = ~n24841 & n24851;
  assign n24853 = ~n24840 & ~n24852;
  assign n24854 = ~n24757 & ~n24853;
  assign n24855 = n24757 & n24853;
  assign n24856 = n24206 & n24257;
  assign n24857 = ~n24258 & ~n24856;
  assign n24858 = ~n24855 & n24857;
  assign n24859 = ~n24854 & ~n24858;
  assign n24860 = ~n24747 & ~n24859;
  assign n24861 = n24747 & n24859;
  assign n24862 = n24259 & ~n24261;
  assign n24863 = ~n24262 & ~n24862;
  assign n24864 = ~n24861 & n24863;
  assign n24865 = ~n24860 & ~n24864;
  assign n24866 = ~n24737 & ~n24865;
  assign n24867 = n24737 & n24865;
  assign n24868 = n24175 & n24263;
  assign n24869 = ~n24264 & ~n24868;
  assign n24870 = ~n24867 & n24869;
  assign n24871 = ~n24866 & ~n24870;
  assign n24872 = n24727 & ~n24871;
  assign n24873 = ~n24727 & n24871;
  assign n24874 = n11055 & n21063;
  assign n24875 = n11056 & n21613;
  assign n24876 = n11661 & n21060;
  assign n24877 = n11672 & n21057;
  assign n24878 = ~n24874 & ~n24876;
  assign n24879 = ~n24877 & n24878;
  assign n24880 = ~n24875 & n24879;
  assign n24881 = pi2  & ~n24880;
  assign n24882 = ~pi2  & n24880;
  assign n24883 = ~n24881 & ~n24882;
  assign n24884 = ~n24873 & n24883;
  assign n24885 = ~n24872 & ~n24884;
  assign n24886 = n24725 & ~n24885;
  assign n24887 = ~n24725 & n24885;
  assign n24888 = n11055 & n21060;
  assign n24889 = n11056 & n21318;
  assign n24890 = n11661 & n21057;
  assign n24891 = n11672 & n21054;
  assign n24892 = ~n24888 & ~n24890;
  assign n24893 = ~n24891 & n24892;
  assign n24894 = ~n24889 & n24893;
  assign n24895 = pi2  & ~n24894;
  assign n24896 = ~pi2  & n24894;
  assign n24897 = ~n24895 & ~n24896;
  assign n24898 = ~n24887 & n24897;
  assign n24899 = ~n24886 & ~n24898;
  assign n24900 = n24723 & ~n24899;
  assign n24901 = ~n24723 & n24899;
  assign n24902 = n11055 & n21057;
  assign n24903 = n11056 & n21825;
  assign n24904 = n11661 & n21054;
  assign n24905 = n11672 & n21051;
  assign n24906 = ~n24902 & ~n24904;
  assign n24907 = ~n24905 & n24906;
  assign n24908 = ~n24903 & n24907;
  assign n24909 = pi2  & ~n24908;
  assign n24910 = ~pi2  & n24908;
  assign n24911 = ~n24909 & ~n24910;
  assign n24912 = ~n24901 & n24911;
  assign n24913 = ~n24900 & ~n24912;
  assign n24914 = ~n24721 & ~n24913;
  assign n24915 = n24721 & n24913;
  assign n24916 = n24279 & ~n24281;
  assign n24917 = ~n24282 & ~n24916;
  assign n24918 = ~n24915 & n24917;
  assign n24919 = ~n24914 & ~n24918;
  assign n24920 = ~n24711 & ~n24919;
  assign n24921 = n24711 & n24919;
  assign n24922 = n24106 & n24283;
  assign n24923 = ~n24284 & ~n24922;
  assign n24924 = ~n24921 & n24923;
  assign n24925 = ~n24920 & ~n24924;
  assign n24926 = ~n24701 & ~n24925;
  assign n24927 = n24701 & n24925;
  assign n24928 = n24090 & n24285;
  assign n24929 = ~n24286 & ~n24928;
  assign n24930 = ~n24927 & n24929;
  assign n24931 = ~n24926 & ~n24930;
  assign n24932 = n24691 & ~n24931;
  assign n24933 = ~n24691 & n24931;
  assign n24934 = n11055 & n21045;
  assign n24935 = n11056 & n22217;
  assign n24936 = n11661 & n21042;
  assign n24937 = n11672 & n21039;
  assign n24938 = ~n24934 & ~n24936;
  assign n24939 = ~n24937 & n24938;
  assign n24940 = ~n24935 & n24939;
  assign n24941 = pi2  & ~n24940;
  assign n24942 = ~pi2  & n24940;
  assign n24943 = ~n24941 & ~n24942;
  assign n24944 = ~n24933 & n24943;
  assign n24945 = ~n24932 & ~n24944;
  assign n24946 = n24689 & ~n24945;
  assign n24947 = ~n24689 & n24945;
  assign n24948 = n11055 & n21042;
  assign n24949 = n11056 & n22199;
  assign n24950 = n11661 & n21039;
  assign n24951 = n11672 & n21036;
  assign n24952 = ~n24948 & ~n24950;
  assign n24953 = ~n24951 & n24952;
  assign n24954 = ~n24949 & n24953;
  assign n24955 = pi2  & ~n24954;
  assign n24956 = ~pi2  & n24954;
  assign n24957 = ~n24955 & ~n24956;
  assign n24958 = ~n24947 & n24957;
  assign n24959 = ~n24946 & ~n24958;
  assign n24960 = n24687 & ~n24959;
  assign n24961 = ~n24687 & n24959;
  assign n24962 = n11055 & n21039;
  assign n24963 = n11056 & n22186;
  assign n24964 = n11661 & n21036;
  assign n24965 = n11672 & n21033;
  assign n24966 = ~n24962 & ~n24964;
  assign n24967 = ~n24965 & n24966;
  assign n24968 = ~n24963 & n24967;
  assign n24969 = pi2  & ~n24968;
  assign n24970 = ~pi2  & n24968;
  assign n24971 = ~n24969 & ~n24970;
  assign n24972 = ~n24961 & n24971;
  assign n24973 = ~n24960 & ~n24972;
  assign n24974 = ~n24685 & ~n24973;
  assign n24975 = n24685 & n24973;
  assign n24976 = n24035 & n24301;
  assign n24977 = ~n24302 & ~n24976;
  assign n24978 = ~n24975 & n24977;
  assign n24979 = ~n24974 & ~n24978;
  assign n24980 = ~n24675 & ~n24979;
  assign n24981 = n24675 & n24979;
  assign n24982 = n24303 & ~n24305;
  assign n24983 = ~n24306 & ~n24982;
  assign n24984 = ~n24981 & n24983;
  assign n24985 = ~n24980 & ~n24984;
  assign n24986 = ~n24665 & ~n24985;
  assign n24987 = n24665 & n24985;
  assign n24988 = n24005 & n24307;
  assign n24989 = ~n24308 & ~n24988;
  assign n24990 = ~n24987 & n24989;
  assign n24991 = ~n24986 & ~n24990;
  assign n24992 = n24655 & ~n24991;
  assign n24993 = ~n24655 & n24991;
  assign n24994 = n11055 & n21027;
  assign n24995 = n11056 & n21306;
  assign n24996 = n11661 & n21024;
  assign n24997 = n11672 & n21021;
  assign n24998 = ~n24994 & ~n24996;
  assign n24999 = ~n24997 & n24998;
  assign n25000 = ~n24995 & n24999;
  assign n25001 = pi2  & ~n25000;
  assign n25002 = ~pi2  & n25000;
  assign n25003 = ~n25001 & ~n25002;
  assign n25004 = ~n24993 & n25003;
  assign n25005 = ~n24992 & ~n25004;
  assign n25006 = n24653 & ~n25005;
  assign n25007 = ~n24653 & n25005;
  assign n25008 = n11055 & n21024;
  assign n25009 = n11056 & n23033;
  assign n25010 = n11661 & n21021;
  assign n25011 = n11672 & n21018;
  assign n25012 = ~n25008 & ~n25010;
  assign n25013 = ~n25011 & n25012;
  assign n25014 = ~n25009 & n25013;
  assign n25015 = pi2  & ~n25014;
  assign n25016 = ~pi2  & n25014;
  assign n25017 = ~n25015 & ~n25016;
  assign n25018 = ~n25007 & n25017;
  assign n25019 = ~n25006 & ~n25018;
  assign n25020 = n24651 & ~n25019;
  assign n25021 = ~n24651 & n25019;
  assign n25022 = n11055 & n21021;
  assign n25023 = n11056 & n23220;
  assign n25024 = n11661 & n21018;
  assign n25025 = n11672 & n21015;
  assign n25026 = ~n25022 & ~n25024;
  assign n25027 = ~n25025 & n25026;
  assign n25028 = ~n25023 & n25027;
  assign n25029 = pi2  & ~n25028;
  assign n25030 = ~pi2  & n25028;
  assign n25031 = ~n25029 & ~n25030;
  assign n25032 = ~n25021 & n25031;
  assign n25033 = ~n25020 & ~n25032;
  assign n25034 = ~n24649 & ~n25033;
  assign n25035 = n24649 & n25033;
  assign n25036 = n24323 & ~n24325;
  assign n25037 = ~n24326 & ~n25036;
  assign n25038 = ~n25035 & n25037;
  assign n25039 = ~n25034 & ~n25038;
  assign n25040 = ~n24639 & ~n25039;
  assign n25041 = n24639 & n25039;
  assign n25042 = n23936 & n24327;
  assign n25043 = ~n24328 & ~n25042;
  assign n25044 = ~n25041 & n25043;
  assign n25045 = ~n25040 & ~n25044;
  assign n25046 = ~n24629 & ~n25045;
  assign n25047 = n24629 & n25045;
  assign n25048 = n23920 & n24329;
  assign n25049 = ~n24330 & ~n25048;
  assign n25050 = ~n25047 & n25049;
  assign n25051 = ~n25046 & ~n25050;
  assign n25052 = n24619 & ~n25051;
  assign n25053 = ~n24619 & n25051;
  assign n25054 = n11055 & n21009;
  assign n25055 = n11056 & n23851;
  assign n25056 = n11661 & n21006;
  assign n25057 = n11672 & n20906;
  assign n25058 = ~n25054 & ~n25056;
  assign n25059 = ~n25057 & n25058;
  assign n25060 = ~n25055 & n25059;
  assign n25061 = pi2  & ~n25060;
  assign n25062 = ~pi2  & n25060;
  assign n25063 = ~n25061 & ~n25062;
  assign n25064 = ~n25053 & n25063;
  assign n25065 = ~n25052 & ~n25064;
  assign n25066 = n24617 & ~n25065;
  assign n25067 = ~n24617 & n25065;
  assign n25068 = n11055 & n21006;
  assign n25069 = n11056 & n23833;
  assign n25070 = n11661 & n20906;
  assign n25071 = n11672 & n21003;
  assign n25072 = ~n25068 & ~n25070;
  assign n25073 = ~n25071 & n25072;
  assign n25074 = ~n25069 & n25073;
  assign n25075 = pi2  & ~n25074;
  assign n25076 = ~pi2  & n25074;
  assign n25077 = ~n25075 & ~n25076;
  assign n25078 = ~n25067 & n25077;
  assign n25079 = ~n25066 & ~n25078;
  assign n25080 = ~n24615 & ~n25079;
  assign n25081 = n24615 & n25079;
  assign n25082 = n24340 & ~n24342;
  assign n25083 = ~n24343 & ~n25082;
  assign n25084 = ~n25081 & n25083;
  assign n25085 = ~n25080 & ~n25084;
  assign n25086 = ~n24605 & ~n25085;
  assign n25087 = n24605 & n25085;
  assign n25088 = n24344 & ~n24346;
  assign n25089 = ~n24347 & ~n25088;
  assign n25090 = ~n25087 & n25089;
  assign n25091 = ~n25086 & ~n25090;
  assign n25092 = ~n24593 & ~n25091;
  assign n25093 = n24593 & n25091;
  assign n25094 = n23848 & n24348;
  assign n25095 = ~n24349 & ~n25094;
  assign n25096 = ~n25093 & n25095;
  assign n25097 = ~n25092 & ~n25096;
  assign n25098 = ~n24581 & ~n25097;
  assign n25099 = ~n24578 & ~n25098;
  assign n25100 = n75 & n21003;
  assign n25101 = n9491 & n24596;
  assign n25102 = n10469 & n21288;
  assign n25103 = n11031 & n24428;
  assign n25104 = ~n25100 & ~n25102;
  assign n25105 = ~n25103 & n25104;
  assign n25106 = ~n25101 & n25105;
  assign n25107 = ~pi5  & ~n25106;
  assign n25108 = pi5  & n25106;
  assign n25109 = ~n25107 & ~n25108;
  assign n25110 = n23809 & ~n23821;
  assign n25111 = ~n23825 & ~n25110;
  assign n25112 = ~n23804 & ~n23808;
  assign n25113 = n7430 & n21018;
  assign n25114 = n7431 & n23205;
  assign n25115 = n7869 & n21015;
  assign n25116 = n7895 & n21012;
  assign n25117 = ~n25113 & ~n25115;
  assign n25118 = ~n25116 & n25117;
  assign n25119 = ~n25114 & n25118;
  assign n25120 = ~pi11  & ~n25119;
  assign n25121 = pi11  & n25119;
  assign n25122 = ~n25120 & ~n25121;
  assign n25123 = n23787 & ~n23797;
  assign n25124 = ~n23668 & ~n23800;
  assign n25125 = ~n25123 & ~n25124;
  assign n25126 = n5982 & n21036;
  assign n25127 = n5983 & n22632;
  assign n25128 = n6323 & n21033;
  assign n25129 = n6336 & n21030;
  assign n25130 = ~n25126 & ~n25128;
  assign n25131 = ~n25129 & n25130;
  assign n25132 = ~n25127 & n25131;
  assign n25133 = ~pi17  & ~n25132;
  assign n25134 = pi17  & n25132;
  assign n25135 = ~n25133 & ~n25134;
  assign n25136 = n23763 & ~n23773;
  assign n25137 = ~n23777 & ~n25136;
  assign n25138 = ~n23758 & ~n23762;
  assign n25139 = n5044 & n21054;
  assign n25140 = n5045 & n21812;
  assign n25141 = n5109 & n21051;
  assign n25142 = n5130 & n21048;
  assign n25143 = ~n25139 & ~n25141;
  assign n25144 = ~n25142 & n25143;
  assign n25145 = ~n25140 & n25144;
  assign n25146 = ~pi23  & ~n25145;
  assign n25147 = pi23  & n25145;
  assign n25148 = ~n25146 & ~n25147;
  assign n25149 = n23741 & ~n23751;
  assign n25150 = ~n23694 & ~n23754;
  assign n25151 = ~n25149 & ~n25150;
  assign n25152 = n3810 & n21072;
  assign n25153 = n3886 & n21428;
  assign n25154 = n3884 & n21069;
  assign n25155 = n4380 & n21066;
  assign n25156 = ~n25152 & ~n25154;
  assign n25157 = ~n25155 & n25156;
  assign n25158 = ~n25153 & n25157;
  assign n25159 = ~pi29  & ~n25158;
  assign n25160 = pi29  & n25158;
  assign n25161 = ~n25159 & ~n25160;
  assign n25162 = ~n23720 & ~n23727;
  assign n25163 = ~n23731 & ~n25162;
  assign n25164 = ~n156 & ~n329;
  assign n25165 = ~n376 & ~n838;
  assign n25166 = n25164 & n25165;
  assign n25167 = n298 & n354;
  assign n25168 = n1122 & n1420;
  assign n25169 = n1859 & n3911;
  assign n25170 = n25168 & n25169;
  assign n25171 = n25166 & n25167;
  assign n25172 = n2678 & n25171;
  assign n25173 = n5273 & n25170;
  assign n25174 = n12666 & n25173;
  assign n25175 = n4332 & n25172;
  assign n25176 = n25174 & n25175;
  assign n25177 = n4844 & n25176;
  assign n25178 = n12943 & n25177;
  assign n25179 = n3692 & n21078;
  assign n25180 = n880 & n21330;
  assign n25181 = n748 & n21081;
  assign n25182 = n3694 & n21075;
  assign n25183 = ~n25179 & ~n25181;
  assign n25184 = ~n25182 & n25183;
  assign n25185 = ~n25180 & n25184;
  assign n25186 = ~n25178 & n25185;
  assign n25187 = n25178 & ~n25185;
  assign n25188 = ~n25186 & ~n25187;
  assign n25189 = ~n25163 & ~n25188;
  assign n25190 = n25163 & n25188;
  assign n25191 = ~n25189 & ~n25190;
  assign n25192 = ~n25161 & ~n25191;
  assign n25193 = n25161 & n25191;
  assign n25194 = ~n25192 & ~n25193;
  assign n25195 = ~n23704 & n23733;
  assign n25196 = ~n23740 & ~n25195;
  assign n25197 = n25194 & n25196;
  assign n25198 = ~n25194 & ~n25196;
  assign n25199 = ~n25197 & ~n25198;
  assign n25200 = n86 & n21063;
  assign n25201 = n4420 & n21613;
  assign n25202 = n4600 & n21060;
  assign n25203 = n4615 & n21057;
  assign n25204 = ~n25200 & ~n25202;
  assign n25205 = ~n25203 & n25204;
  assign n25206 = ~n25201 & n25205;
  assign n25207 = pi26  & n25206;
  assign n25208 = ~pi26  & ~n25206;
  assign n25209 = ~n25207 & ~n25208;
  assign n25210 = n25199 & n25209;
  assign n25211 = ~n25199 & ~n25209;
  assign n25212 = ~n25210 & ~n25211;
  assign n25213 = ~n25151 & n25212;
  assign n25214 = n25151 & ~n25212;
  assign n25215 = ~n25213 & ~n25214;
  assign n25216 = ~n25148 & ~n25215;
  assign n25217 = n25148 & n25215;
  assign n25218 = ~n25216 & ~n25217;
  assign n25219 = n25138 & ~n25218;
  assign n25220 = ~n25138 & n25218;
  assign n25221 = ~n25219 & ~n25220;
  assign n25222 = n5240 & n21045;
  assign n25223 = n5241 & n22217;
  assign n25224 = n5853 & n21042;
  assign n25225 = n5866 & n21039;
  assign n25226 = ~n25222 & ~n25224;
  assign n25227 = ~n25225 & n25226;
  assign n25228 = ~n25223 & n25227;
  assign n25229 = pi20  & n25228;
  assign n25230 = ~pi20  & ~n25228;
  assign n25231 = ~n25229 & ~n25230;
  assign n25232 = n25221 & n25231;
  assign n25233 = ~n25221 & ~n25231;
  assign n25234 = ~n25232 & ~n25233;
  assign n25235 = ~n25137 & ~n25234;
  assign n25236 = n25137 & n25234;
  assign n25237 = ~n25235 & ~n25236;
  assign n25238 = ~n25135 & ~n25237;
  assign n25239 = n25135 & n25237;
  assign n25240 = ~n25238 & ~n25239;
  assign n25241 = ~n23678 & n23779;
  assign n25242 = ~n23786 & ~n25241;
  assign n25243 = n25240 & n25242;
  assign n25244 = ~n25240 & ~n25242;
  assign n25245 = ~n25243 & ~n25244;
  assign n25246 = n6630 & n21027;
  assign n25247 = n6631 & n21306;
  assign n25248 = n7238 & n21024;
  assign n25249 = n7262 & n21021;
  assign n25250 = ~n25246 & ~n25248;
  assign n25251 = ~n25249 & n25250;
  assign n25252 = ~n25247 & n25251;
  assign n25253 = pi14  & n25252;
  assign n25254 = ~pi14  & ~n25252;
  assign n25255 = ~n25253 & ~n25254;
  assign n25256 = n25245 & n25255;
  assign n25257 = ~n25245 & ~n25255;
  assign n25258 = ~n25256 & ~n25257;
  assign n25259 = ~n25125 & n25258;
  assign n25260 = n25125 & ~n25258;
  assign n25261 = ~n25259 & ~n25260;
  assign n25262 = ~n25122 & ~n25261;
  assign n25263 = n25122 & n25261;
  assign n25264 = ~n25262 & ~n25263;
  assign n25265 = n25112 & ~n25264;
  assign n25266 = ~n25112 & n25264;
  assign n25267 = ~n25265 & ~n25266;
  assign n25268 = n8250 & n21009;
  assign n25269 = n8251 & n23851;
  assign n25270 = n9016 & n21006;
  assign n25271 = n9040 & n20906;
  assign n25272 = ~n25268 & ~n25270;
  assign n25273 = ~n25271 & n25272;
  assign n25274 = ~n25269 & n25273;
  assign n25275 = pi8  & n25274;
  assign n25276 = ~pi8  & ~n25274;
  assign n25277 = ~n25275 & ~n25276;
  assign n25278 = n25267 & n25277;
  assign n25279 = ~n25267 & ~n25277;
  assign n25280 = ~n25278 & ~n25279;
  assign n25281 = ~n25111 & ~n25280;
  assign n25282 = n25111 & n25280;
  assign n25283 = ~n25281 & ~n25282;
  assign n25284 = ~n25109 & ~n25283;
  assign n25285 = n25109 & n25283;
  assign n25286 = ~n25284 & ~n25285;
  assign n25287 = ~n21303 & n23827;
  assign n25288 = ~n24352 & ~n25287;
  assign n25289 = n25286 & n25288;
  assign n25290 = ~n25286 & ~n25288;
  assign n25291 = ~n25289 & ~n25290;
  assign n25292 = n11055 & n24494;
  assign n25293 = ~n24563 & ~n24566;
  assign n25294 = ~n24557 & ~n24561;
  assign n25295 = ~n24549 & ~n24553;
  assign n25296 = ~n24531 & ~n24533;
  assign n25297 = ~n304 & n3880;
  assign n25298 = n3673 & n25297;
  assign n25299 = n24524 & n25298;
  assign n25300 = ~n25296 & n25299;
  assign n25301 = n25296 & ~n25299;
  assign n25302 = ~n25300 & ~n25301;
  assign n25303 = n748 & n12392;
  assign n25304 = n880 & n13421;
  assign n25305 = n3692 & n12646;
  assign n25306 = n3694 & n13164;
  assign n25307 = ~n25303 & ~n25305;
  assign n25308 = ~n25306 & n25307;
  assign n25309 = ~n25304 & n25308;
  assign n25310 = n25302 & ~n25309;
  assign n25311 = ~n25302 & n25309;
  assign n25312 = ~n25310 & ~n25311;
  assign n25313 = ~n24536 & n24545;
  assign n25314 = ~n24537 & ~n25313;
  assign n25315 = ~n25312 & ~n25314;
  assign n25316 = n25312 & n25314;
  assign n25317 = ~n25315 & ~n25316;
  assign n25318 = n4380 & ~n12786;
  assign n25319 = n3886 & ~n13781;
  assign n25320 = n3810 & n13166;
  assign n25321 = n3884 & n13161;
  assign n25322 = ~n25318 & ~n25320;
  assign n25323 = ~n25321 & n25322;
  assign n25324 = ~n25319 & n25323;
  assign n25325 = pi29  & n25324;
  assign n25326 = ~pi29  & ~n25324;
  assign n25327 = ~n25325 & ~n25326;
  assign n25328 = n25317 & ~n25327;
  assign n25329 = ~n25317 & n25327;
  assign n25330 = ~n25328 & ~n25329;
  assign n25331 = ~n25295 & n25330;
  assign n25332 = n25295 & ~n25330;
  assign n25333 = ~n25331 & ~n25332;
  assign n25334 = ~n25294 & n25333;
  assign n25335 = n25294 & ~n25333;
  assign n25336 = ~n25334 & ~n25335;
  assign n25337 = n24562 & n25336;
  assign n25338 = ~n24562 & ~n25336;
  assign n25339 = ~n25337 & ~n25338;
  assign n25340 = ~n25293 & n25339;
  assign n25341 = n25293 & ~n25339;
  assign n25342 = ~n25340 & ~n25341;
  assign n25343 = n11056 & n25342;
  assign n25344 = n11661 & n24562;
  assign n25345 = n11672 & n25336;
  assign n25346 = ~n25292 & ~n25344;
  assign n25347 = ~n25345 & n25346;
  assign n25348 = ~n25343 & n25347;
  assign n25349 = pi2  & n25348;
  assign n25350 = ~pi2  & ~n25348;
  assign n25351 = ~n25349 & ~n25350;
  assign n25352 = n25291 & ~n25351;
  assign n25353 = ~n25291 & n25351;
  assign n25354 = ~n25352 & ~n25353;
  assign n25355 = ~n25099 & n25354;
  assign n25356 = n25099 & ~n25354;
  assign n25357 = ~n25355 & ~n25356;
  assign n25358 = n24581 & ~n25097;
  assign n25359 = ~n24581 & n25097;
  assign n25360 = ~n25358 & ~n25359;
  assign n25361 = n25357 & ~n25360;
  assign n25362 = ~n25357 & n25360;
  assign po0  = ~n25361 & ~n25362;
  assign n25364 = ~n25352 & ~n25355;
  assign n25365 = ~n25109 & n25283;
  assign n25366 = ~n25290 & ~n25365;
  assign n25367 = n75 & n21288;
  assign n25368 = n9491 & n24584;
  assign n25369 = n10469 & n24428;
  assign n25370 = n11031 & n24494;
  assign n25371 = ~n25367 & ~n25369;
  assign n25372 = ~n25370 & n25371;
  assign n25373 = ~n25368 & n25372;
  assign n25374 = ~pi5  & ~n25373;
  assign n25375 = pi5  & n25373;
  assign n25376 = ~n25374 & ~n25375;
  assign n25377 = n25267 & ~n25277;
  assign n25378 = ~n25281 & ~n25377;
  assign n25379 = n7430 & n21015;
  assign n25380 = n7431 & n23190;
  assign n25381 = n7869 & n21012;
  assign n25382 = n7895 & n21009;
  assign n25383 = ~n25379 & ~n25381;
  assign n25384 = ~n25382 & n25383;
  assign n25385 = ~n25380 & n25384;
  assign n25386 = ~pi11  & ~n25385;
  assign n25387 = pi11  & n25385;
  assign n25388 = ~n25386 & ~n25387;
  assign n25389 = n25245 & ~n25255;
  assign n25390 = ~n25125 & ~n25258;
  assign n25391 = ~n25389 & ~n25390;
  assign n25392 = ~n25135 & n25237;
  assign n25393 = ~n25244 & ~n25392;
  assign n25394 = n5982 & n21033;
  assign n25395 = n5983 & n22674;
  assign n25396 = n6323 & n21030;
  assign n25397 = n6336 & n21027;
  assign n25398 = ~n25394 & ~n25396;
  assign n25399 = ~n25397 & n25398;
  assign n25400 = ~n25395 & n25399;
  assign n25401 = ~pi17  & ~n25400;
  assign n25402 = pi17  & n25400;
  assign n25403 = ~n25401 & ~n25402;
  assign n25404 = n25221 & ~n25231;
  assign n25405 = ~n25235 & ~n25404;
  assign n25406 = n5044 & n21051;
  assign n25407 = n5045 & n21797;
  assign n25408 = n5109 & n21048;
  assign n25409 = n5130 & n21045;
  assign n25410 = ~n25406 & ~n25408;
  assign n25411 = ~n25409 & n25410;
  assign n25412 = ~n25407 & n25411;
  assign n25413 = ~pi23  & ~n25412;
  assign n25414 = pi23  & n25412;
  assign n25415 = ~n25413 & ~n25414;
  assign n25416 = n25199 & ~n25209;
  assign n25417 = ~n25151 & ~n25212;
  assign n25418 = ~n25416 & ~n25417;
  assign n25419 = ~n25161 & n25191;
  assign n25420 = ~n25198 & ~n25419;
  assign n25421 = n3810 & n21069;
  assign n25422 = n3886 & n21592;
  assign n25423 = n3884 & n21066;
  assign n25424 = n4380 & n21063;
  assign n25425 = ~n25421 & ~n25423;
  assign n25426 = ~n25424 & n25425;
  assign n25427 = ~n25422 & n25426;
  assign n25428 = pi29  & n25427;
  assign n25429 = ~pi29  & ~n25427;
  assign n25430 = ~n25428 & ~n25429;
  assign n25431 = ~n25178 & ~n25185;
  assign n25432 = ~n25189 & ~n25431;
  assign n25433 = ~n282 & ~n370;
  assign n25434 = ~n411 & ~n634;
  assign n25435 = n2261 & n25434;
  assign n25436 = n142 & n25433;
  assign n25437 = n298 & n514;
  assign n25438 = n2452 & n2473;
  assign n25439 = n3325 & n25438;
  assign n25440 = n25436 & n25437;
  assign n25441 = n1280 & n25435;
  assign n25442 = n2804 & n25441;
  assign n25443 = n25439 & n25440;
  assign n25444 = n6944 & n25443;
  assign n25445 = n7024 & n25442;
  assign n25446 = n25444 & n25445;
  assign n25447 = n3163 & n13627;
  assign n25448 = n25446 & n25447;
  assign n25449 = n1376 & n25448;
  assign n25450 = n3692 & n21075;
  assign n25451 = n880 & n21459;
  assign n25452 = n748 & n21078;
  assign n25453 = n3694 & n21072;
  assign n25454 = ~n25450 & ~n25452;
  assign n25455 = ~n25453 & n25454;
  assign n25456 = ~n25451 & n25455;
  assign n25457 = ~n25449 & n25456;
  assign n25458 = n25449 & ~n25456;
  assign n25459 = ~n25457 & ~n25458;
  assign n25460 = ~n25432 & ~n25459;
  assign n25461 = n25432 & n25459;
  assign n25462 = ~n25460 & ~n25461;
  assign n25463 = ~n25430 & n25462;
  assign n25464 = n25430 & ~n25462;
  assign n25465 = ~n25463 & ~n25464;
  assign n25466 = ~n25420 & n25465;
  assign n25467 = n25420 & ~n25465;
  assign n25468 = ~n25466 & ~n25467;
  assign n25469 = n86 & n21060;
  assign n25470 = n4420 & n21318;
  assign n25471 = n4600 & n21057;
  assign n25472 = n4615 & n21054;
  assign n25473 = ~n25469 & ~n25471;
  assign n25474 = ~n25472 & n25473;
  assign n25475 = ~n25470 & n25474;
  assign n25476 = pi26  & n25475;
  assign n25477 = ~pi26  & ~n25475;
  assign n25478 = ~n25476 & ~n25477;
  assign n25479 = n25468 & n25478;
  assign n25480 = ~n25468 & ~n25478;
  assign n25481 = ~n25479 & ~n25480;
  assign n25482 = ~n25418 & ~n25481;
  assign n25483 = n25418 & n25481;
  assign n25484 = ~n25482 & ~n25483;
  assign n25485 = ~n25415 & ~n25484;
  assign n25486 = n25415 & n25484;
  assign n25487 = ~n25485 & ~n25486;
  assign n25488 = ~n25216 & ~n25220;
  assign n25489 = n25487 & n25488;
  assign n25490 = ~n25487 & ~n25488;
  assign n25491 = ~n25489 & ~n25490;
  assign n25492 = n5240 & n21042;
  assign n25493 = n5241 & n22199;
  assign n25494 = n5853 & n21039;
  assign n25495 = n5866 & n21036;
  assign n25496 = ~n25492 & ~n25494;
  assign n25497 = ~n25495 & n25496;
  assign n25498 = ~n25493 & n25497;
  assign n25499 = pi20  & n25498;
  assign n25500 = ~pi20  & ~n25498;
  assign n25501 = ~n25499 & ~n25500;
  assign n25502 = n25491 & n25501;
  assign n25503 = ~n25491 & ~n25501;
  assign n25504 = ~n25502 & ~n25503;
  assign n25505 = ~n25405 & n25504;
  assign n25506 = n25405 & ~n25504;
  assign n25507 = ~n25505 & ~n25506;
  assign n25508 = ~n25403 & ~n25507;
  assign n25509 = n25403 & n25507;
  assign n25510 = ~n25508 & ~n25509;
  assign n25511 = n25393 & ~n25510;
  assign n25512 = ~n25393 & n25510;
  assign n25513 = ~n25511 & ~n25512;
  assign n25514 = n6630 & n21024;
  assign n25515 = n6631 & n23033;
  assign n25516 = n7238 & n21021;
  assign n25517 = n7262 & n21018;
  assign n25518 = ~n25514 & ~n25516;
  assign n25519 = ~n25517 & n25518;
  assign n25520 = ~n25515 & n25519;
  assign n25521 = pi14  & n25520;
  assign n25522 = ~pi14  & ~n25520;
  assign n25523 = ~n25521 & ~n25522;
  assign n25524 = n25513 & n25523;
  assign n25525 = ~n25513 & ~n25523;
  assign n25526 = ~n25524 & ~n25525;
  assign n25527 = ~n25391 & ~n25526;
  assign n25528 = n25391 & n25526;
  assign n25529 = ~n25527 & ~n25528;
  assign n25530 = ~n25388 & ~n25529;
  assign n25531 = n25388 & n25529;
  assign n25532 = ~n25530 & ~n25531;
  assign n25533 = ~n25262 & ~n25266;
  assign n25534 = n25532 & n25533;
  assign n25535 = ~n25532 & ~n25533;
  assign n25536 = ~n25534 & ~n25535;
  assign n25537 = n8250 & n21006;
  assign n25538 = n8251 & n23833;
  assign n25539 = n9016 & n20906;
  assign n25540 = n9040 & n21003;
  assign n25541 = ~n25537 & ~n25539;
  assign n25542 = ~n25540 & n25541;
  assign n25543 = ~n25538 & n25542;
  assign n25544 = pi8  & n25543;
  assign n25545 = ~pi8  & ~n25543;
  assign n25546 = ~n25544 & ~n25545;
  assign n25547 = n25536 & n25546;
  assign n25548 = ~n25536 & ~n25546;
  assign n25549 = ~n25547 & ~n25548;
  assign n25550 = ~n25378 & n25549;
  assign n25551 = n25378 & ~n25549;
  assign n25552 = ~n25550 & ~n25551;
  assign n25553 = ~n25376 & ~n25552;
  assign n25554 = n25376 & n25552;
  assign n25555 = ~n25553 & ~n25554;
  assign n25556 = n25366 & ~n25555;
  assign n25557 = ~n25366 & n25555;
  assign n25558 = ~n25556 & ~n25557;
  assign n25559 = n11055 & n24562;
  assign n25560 = ~n25337 & ~n25340;
  assign n25561 = ~n25331 & ~n25334;
  assign n25562 = ~n25316 & ~n25328;
  assign n25563 = n3810 & n13161;
  assign n25564 = n3886 & ~n13280;
  assign n25565 = ~n3809 & ~n3886;
  assign n25566 = ~n12786 & n25565;
  assign n25567 = ~n25563 & ~n25566;
  assign n25568 = ~n25564 & n25567;
  assign n25569 = ~pi29  & ~n25568;
  assign n25570 = pi29  & n25568;
  assign n25571 = ~n25569 & ~n25570;
  assign n25572 = n748 & n12646;
  assign n25573 = n880 & n13261;
  assign n25574 = n3692 & n13164;
  assign n25575 = n3694 & n13166;
  assign n25576 = ~n25572 & ~n25574;
  assign n25577 = ~n25575 & n25576;
  assign n25578 = ~n25573 & n25577;
  assign n25579 = ~n25571 & n25578;
  assign n25580 = n25571 & ~n25578;
  assign n25581 = ~n25579 & ~n25580;
  assign n25582 = n3834 & n3882;
  assign n25583 = n25299 & ~n25582;
  assign n25584 = ~n25299 & n25582;
  assign n25585 = ~n25583 & ~n25584;
  assign n25586 = ~n25300 & n25309;
  assign n25587 = ~n25301 & ~n25586;
  assign n25588 = n25585 & n25587;
  assign n25589 = ~n25585 & ~n25587;
  assign n25590 = ~n25588 & ~n25589;
  assign n25591 = ~n25581 & n25590;
  assign n25592 = n25581 & ~n25590;
  assign n25593 = ~n25591 & ~n25592;
  assign n25594 = ~n25562 & n25593;
  assign n25595 = n25562 & ~n25593;
  assign n25596 = ~n25594 & ~n25595;
  assign n25597 = ~n25561 & n25596;
  assign n25598 = n25561 & ~n25596;
  assign n25599 = ~n25597 & ~n25598;
  assign n25600 = ~n25336 & ~n25599;
  assign n25601 = n25336 & n25599;
  assign n25602 = ~n25600 & ~n25601;
  assign n25603 = ~n25560 & n25602;
  assign n25604 = n25560 & ~n25602;
  assign n25605 = ~n25603 & ~n25604;
  assign n25606 = n11056 & n25605;
  assign n25607 = n11661 & n25336;
  assign n25608 = n11672 & n25599;
  assign n25609 = ~n25559 & ~n25607;
  assign n25610 = ~n25608 & n25609;
  assign n25611 = ~n25606 & n25610;
  assign n25612 = pi2  & n25611;
  assign n25613 = ~pi2  & ~n25611;
  assign n25614 = ~n25612 & ~n25613;
  assign n25615 = n25558 & ~n25614;
  assign n25616 = ~n25558 & n25614;
  assign n25617 = ~n25615 & ~n25616;
  assign n25618 = ~n25364 & n25617;
  assign n25619 = n25364 & ~n25617;
  assign n25620 = ~n25618 & ~n25619;
  assign n25621 = n25361 & n25620;
  assign n25622 = ~n25361 & ~n25620;
  assign po1  = ~n25621 & ~n25622;
  assign n25624 = ~n25615 & ~n25618;
  assign n25625 = ~n25553 & ~n25557;
  assign n25626 = n75 & n24428;
  assign n25627 = n9491 & n24568;
  assign n25628 = n10469 & n24494;
  assign n25629 = n11031 & n24562;
  assign n25630 = ~n25626 & ~n25628;
  assign n25631 = ~n25629 & n25630;
  assign n25632 = ~n25627 & n25631;
  assign n25633 = ~pi5  & ~n25632;
  assign n25634 = pi5  & n25632;
  assign n25635 = ~n25633 & ~n25634;
  assign n25636 = n25536 & ~n25546;
  assign n25637 = ~n25378 & ~n25549;
  assign n25638 = ~n25636 & ~n25637;
  assign n25639 = n7430 & n21012;
  assign n25640 = n7431 & n23812;
  assign n25641 = n7869 & n21009;
  assign n25642 = n7895 & n21006;
  assign n25643 = ~n25639 & ~n25641;
  assign n25644 = ~n25642 & n25643;
  assign n25645 = ~n25640 & n25644;
  assign n25646 = ~pi11  & ~n25645;
  assign n25647 = pi11  & n25645;
  assign n25648 = ~n25646 & ~n25647;
  assign n25649 = n25513 & ~n25523;
  assign n25650 = ~n25527 & ~n25649;
  assign n25651 = ~n25508 & ~n25512;
  assign n25652 = n5982 & n21030;
  assign n25653 = n5983 & n22654;
  assign n25654 = n6323 & n21027;
  assign n25655 = n6336 & n21024;
  assign n25656 = ~n25652 & ~n25654;
  assign n25657 = ~n25655 & n25656;
  assign n25658 = ~n25653 & n25657;
  assign n25659 = ~pi17  & ~n25658;
  assign n25660 = pi17  & n25658;
  assign n25661 = ~n25659 & ~n25660;
  assign n25662 = n25491 & ~n25501;
  assign n25663 = ~n25405 & ~n25504;
  assign n25664 = ~n25662 & ~n25663;
  assign n25665 = n5044 & n21048;
  assign n25666 = n5045 & n22049;
  assign n25667 = n5109 & n21045;
  assign n25668 = n5130 & n21042;
  assign n25669 = ~n25665 & ~n25667;
  assign n25670 = ~n25668 & n25669;
  assign n25671 = ~n25666 & n25670;
  assign n25672 = ~pi23  & ~n25671;
  assign n25673 = pi23  & n25671;
  assign n25674 = ~n25672 & ~n25673;
  assign n25675 = n25468 & ~n25478;
  assign n25676 = ~n25482 & ~n25675;
  assign n25677 = ~n25463 & ~n25466;
  assign n25678 = n3810 & n21066;
  assign n25679 = n3886 & n21631;
  assign n25680 = n3884 & n21063;
  assign n25681 = n4380 & n21060;
  assign n25682 = ~n25678 & ~n25680;
  assign n25683 = ~n25681 & n25682;
  assign n25684 = ~n25679 & n25683;
  assign n25685 = pi29  & n25684;
  assign n25686 = ~pi29  & ~n25684;
  assign n25687 = ~n25685 & ~n25686;
  assign n25688 = ~n25449 & ~n25456;
  assign n25689 = ~n25460 & ~n25688;
  assign n25690 = ~n520 & ~n592;
  assign n25691 = ~n599 & ~n639;
  assign n25692 = ~n1032 & n25691;
  assign n25693 = n598 & n25690;
  assign n25694 = n785 & n938;
  assign n25695 = n1306 & n3128;
  assign n25696 = n25694 & n25695;
  assign n25697 = n25692 & n25693;
  assign n25698 = n1700 & n12980;
  assign n25699 = n13666 & n25698;
  assign n25700 = n25696 & n25697;
  assign n25701 = n2623 & n7058;
  assign n25702 = n25700 & n25701;
  assign n25703 = n4312 & n25699;
  assign n25704 = n25702 & n25703;
  assign n25705 = n2435 & n25704;
  assign n25706 = n4287 & n25705;
  assign n25707 = n3692 & n21072;
  assign n25708 = n880 & n21441;
  assign n25709 = n748 & n21075;
  assign n25710 = n3694 & n21069;
  assign n25711 = ~n25707 & ~n25709;
  assign n25712 = ~n25710 & n25711;
  assign n25713 = ~n25708 & n25712;
  assign n25714 = ~n25706 & n25713;
  assign n25715 = n25706 & ~n25713;
  assign n25716 = ~n25714 & ~n25715;
  assign n25717 = ~n25689 & ~n25716;
  assign n25718 = n25689 & n25716;
  assign n25719 = ~n25717 & ~n25718;
  assign n25720 = ~n25687 & n25719;
  assign n25721 = n25687 & ~n25719;
  assign n25722 = ~n25720 & ~n25721;
  assign n25723 = ~n25677 & n25722;
  assign n25724 = n25677 & ~n25722;
  assign n25725 = ~n25723 & ~n25724;
  assign n25726 = n86 & n21057;
  assign n25727 = n4420 & n21825;
  assign n25728 = n4600 & n21054;
  assign n25729 = n4615 & n21051;
  assign n25730 = ~n25726 & ~n25728;
  assign n25731 = ~n25729 & n25730;
  assign n25732 = ~n25727 & n25731;
  assign n25733 = pi26  & n25732;
  assign n25734 = ~pi26  & ~n25732;
  assign n25735 = ~n25733 & ~n25734;
  assign n25736 = n25725 & n25735;
  assign n25737 = ~n25725 & ~n25735;
  assign n25738 = ~n25736 & ~n25737;
  assign n25739 = ~n25676 & ~n25738;
  assign n25740 = n25676 & n25738;
  assign n25741 = ~n25739 & ~n25740;
  assign n25742 = ~n25674 & ~n25741;
  assign n25743 = n25674 & n25741;
  assign n25744 = ~n25742 & ~n25743;
  assign n25745 = ~n25415 & n25484;
  assign n25746 = ~n25490 & ~n25745;
  assign n25747 = n25744 & n25746;
  assign n25748 = ~n25744 & ~n25746;
  assign n25749 = ~n25747 & ~n25748;
  assign n25750 = n5240 & n21039;
  assign n25751 = n5241 & n22186;
  assign n25752 = n5853 & n21036;
  assign n25753 = n5866 & n21033;
  assign n25754 = ~n25750 & ~n25752;
  assign n25755 = ~n25753 & n25754;
  assign n25756 = ~n25751 & n25755;
  assign n25757 = pi20  & n25756;
  assign n25758 = ~pi20  & ~n25756;
  assign n25759 = ~n25757 & ~n25758;
  assign n25760 = n25749 & n25759;
  assign n25761 = ~n25749 & ~n25759;
  assign n25762 = ~n25760 & ~n25761;
  assign n25763 = ~n25664 & n25762;
  assign n25764 = n25664 & ~n25762;
  assign n25765 = ~n25763 & ~n25764;
  assign n25766 = ~n25661 & ~n25765;
  assign n25767 = n25661 & n25765;
  assign n25768 = ~n25766 & ~n25767;
  assign n25769 = n25651 & ~n25768;
  assign n25770 = ~n25651 & n25768;
  assign n25771 = ~n25769 & ~n25770;
  assign n25772 = n6630 & n21021;
  assign n25773 = n6631 & n23220;
  assign n25774 = n7238 & n21018;
  assign n25775 = n7262 & n21015;
  assign n25776 = ~n25772 & ~n25774;
  assign n25777 = ~n25775 & n25776;
  assign n25778 = ~n25773 & n25777;
  assign n25779 = pi14  & n25778;
  assign n25780 = ~pi14  & ~n25778;
  assign n25781 = ~n25779 & ~n25780;
  assign n25782 = n25771 & n25781;
  assign n25783 = ~n25771 & ~n25781;
  assign n25784 = ~n25782 & ~n25783;
  assign n25785 = ~n25650 & ~n25784;
  assign n25786 = n25650 & n25784;
  assign n25787 = ~n25785 & ~n25786;
  assign n25788 = ~n25648 & ~n25787;
  assign n25789 = n25648 & n25787;
  assign n25790 = ~n25788 & ~n25789;
  assign n25791 = ~n25388 & n25529;
  assign n25792 = ~n25535 & ~n25791;
  assign n25793 = n25790 & n25792;
  assign n25794 = ~n25790 & ~n25792;
  assign n25795 = ~n25793 & ~n25794;
  assign n25796 = n8250 & n20906;
  assign n25797 = n8251 & n21294;
  assign n25798 = n9016 & n21003;
  assign n25799 = n9040 & n21288;
  assign n25800 = ~n25796 & ~n25798;
  assign n25801 = ~n25799 & n25800;
  assign n25802 = ~n25797 & n25801;
  assign n25803 = pi8  & n25802;
  assign n25804 = ~pi8  & ~n25802;
  assign n25805 = ~n25803 & ~n25804;
  assign n25806 = n25795 & n25805;
  assign n25807 = ~n25795 & ~n25805;
  assign n25808 = ~n25806 & ~n25807;
  assign n25809 = ~n25638 & n25808;
  assign n25810 = n25638 & ~n25808;
  assign n25811 = ~n25809 & ~n25810;
  assign n25812 = ~n25635 & ~n25811;
  assign n25813 = n25635 & n25811;
  assign n25814 = ~n25812 & ~n25813;
  assign n25815 = n25625 & ~n25814;
  assign n25816 = ~n25625 & n25814;
  assign n25817 = ~n25815 & ~n25816;
  assign n25818 = n11055 & n25336;
  assign n25819 = ~n25601 & ~n25603;
  assign n25820 = ~n25594 & ~n25597;
  assign n25821 = ~n25571 & ~n25578;
  assign n25822 = ~n25591 & ~n25821;
  assign n25823 = ~n25584 & ~n25588;
  assign n25824 = n3804 & n3809;
  assign n25825 = ~n12786 & ~n25824;
  assign n25826 = pi29  & ~n25825;
  assign n25827 = ~pi29  & n25825;
  assign n25828 = ~n25826 & ~n25827;
  assign n25829 = n12760 & n25582;
  assign n25830 = ~n12760 & ~n25582;
  assign n25831 = ~n25829 & ~n25830;
  assign n25832 = n25828 & n25831;
  assign n25833 = ~n25828 & ~n25831;
  assign n25834 = ~n25832 & ~n25833;
  assign n25835 = n3694 & n13161;
  assign n25836 = n880 & n13183;
  assign n25837 = n3692 & n13166;
  assign n25838 = n748 & n13164;
  assign n25839 = ~n25837 & ~n25838;
  assign n25840 = ~n25835 & n25839;
  assign n25841 = ~n25836 & n25840;
  assign n25842 = n25834 & n25841;
  assign n25843 = ~n25834 & ~n25841;
  assign n25844 = ~n25842 & ~n25843;
  assign n25845 = ~n25823 & ~n25844;
  assign n25846 = n25823 & n25844;
  assign n25847 = ~n25845 & ~n25846;
  assign n25848 = ~n25822 & n25847;
  assign n25849 = n25822 & ~n25847;
  assign n25850 = ~n25848 & ~n25849;
  assign n25851 = ~n25820 & n25850;
  assign n25852 = n25820 & ~n25850;
  assign n25853 = ~n25851 & ~n25852;
  assign n25854 = ~n25599 & ~n25853;
  assign n25855 = n25599 & n25853;
  assign n25856 = ~n25854 & ~n25855;
  assign n25857 = ~n25819 & n25856;
  assign n25858 = n25819 & ~n25856;
  assign n25859 = ~n25857 & ~n25858;
  assign n25860 = n11056 & n25859;
  assign n25861 = n11661 & n25599;
  assign n25862 = n11672 & n25853;
  assign n25863 = ~n25818 & ~n25861;
  assign n25864 = ~n25862 & n25863;
  assign n25865 = ~n25860 & n25864;
  assign n25866 = pi2  & n25865;
  assign n25867 = ~pi2  & ~n25865;
  assign n25868 = ~n25866 & ~n25867;
  assign n25869 = n25817 & ~n25868;
  assign n25870 = ~n25817 & n25868;
  assign n25871 = ~n25869 & ~n25870;
  assign n25872 = ~n25624 & n25871;
  assign n25873 = n25624 & ~n25871;
  assign n25874 = ~n25872 & ~n25873;
  assign n25875 = n25621 & n25874;
  assign n25876 = ~n25621 & ~n25874;
  assign po2  = ~n25875 & ~n25876;
  assign n25878 = ~n25869 & ~n25872;
  assign n25879 = ~n25812 & ~n25816;
  assign n25880 = n75 & n24494;
  assign n25881 = n9491 & n25342;
  assign n25882 = n10469 & n24562;
  assign n25883 = n11031 & n25336;
  assign n25884 = ~n25880 & ~n25882;
  assign n25885 = ~n25883 & n25884;
  assign n25886 = ~n25881 & n25885;
  assign n25887 = ~pi5  & ~n25886;
  assign n25888 = pi5  & n25886;
  assign n25889 = ~n25887 & ~n25888;
  assign n25890 = n25795 & ~n25805;
  assign n25891 = ~n25638 & ~n25808;
  assign n25892 = ~n25890 & ~n25891;
  assign n25893 = n7430 & n21009;
  assign n25894 = n7431 & n23851;
  assign n25895 = n7869 & n21006;
  assign n25896 = n7895 & n20906;
  assign n25897 = ~n25893 & ~n25895;
  assign n25898 = ~n25896 & n25897;
  assign n25899 = ~n25894 & n25898;
  assign n25900 = ~pi11  & ~n25899;
  assign n25901 = pi11  & n25899;
  assign n25902 = ~n25900 & ~n25901;
  assign n25903 = n25771 & ~n25781;
  assign n25904 = ~n25785 & ~n25903;
  assign n25905 = ~n25766 & ~n25770;
  assign n25906 = n5982 & n21027;
  assign n25907 = n5983 & n21306;
  assign n25908 = n6323 & n21024;
  assign n25909 = n6336 & n21021;
  assign n25910 = ~n25906 & ~n25908;
  assign n25911 = ~n25909 & n25910;
  assign n25912 = ~n25907 & n25911;
  assign n25913 = ~pi17  & ~n25912;
  assign n25914 = pi17  & n25912;
  assign n25915 = ~n25913 & ~n25914;
  assign n25916 = n25749 & ~n25759;
  assign n25917 = ~n25664 & ~n25762;
  assign n25918 = ~n25916 & ~n25917;
  assign n25919 = n5044 & n21045;
  assign n25920 = n5045 & n22217;
  assign n25921 = n5109 & n21042;
  assign n25922 = n5130 & n21039;
  assign n25923 = ~n25919 & ~n25921;
  assign n25924 = ~n25922 & n25923;
  assign n25925 = ~n25920 & n25924;
  assign n25926 = ~pi23  & ~n25925;
  assign n25927 = pi23  & n25925;
  assign n25928 = ~n25926 & ~n25927;
  assign n25929 = n25725 & ~n25735;
  assign n25930 = ~n25739 & ~n25929;
  assign n25931 = ~n25720 & ~n25723;
  assign n25932 = n3810 & n21063;
  assign n25933 = n3886 & n21613;
  assign n25934 = n3884 & n21060;
  assign n25935 = n4380 & n21057;
  assign n25936 = ~n25932 & ~n25934;
  assign n25937 = ~n25935 & n25936;
  assign n25938 = ~n25933 & n25937;
  assign n25939 = pi29  & n25938;
  assign n25940 = ~pi29  & ~n25938;
  assign n25941 = ~n25939 & ~n25940;
  assign n25942 = ~n25706 & ~n25713;
  assign n25943 = ~n25717 & ~n25942;
  assign n25944 = n500 & n1356;
  assign n25945 = n1380 & n25944;
  assign n25946 = ~n200 & ~n770;
  assign n25947 = n478 & n25946;
  assign n25948 = n1012 & n1538;
  assign n25949 = n3128 & n25948;
  assign n25950 = n2499 & n25947;
  assign n25951 = n2521 & n5270;
  assign n25952 = n25950 & n25951;
  assign n25953 = n25945 & n25949;
  assign n25954 = n25952 & n25953;
  assign n25955 = n14771 & n25954;
  assign n25956 = n2990 & n25955;
  assign n25957 = n4081 & n7082;
  assign n25958 = n25956 & n25957;
  assign n25959 = n3692 & n21069;
  assign n25960 = n880 & n21428;
  assign n25961 = n748 & n21072;
  assign n25962 = n3694 & n21066;
  assign n25963 = ~n25959 & ~n25961;
  assign n25964 = ~n25962 & n25963;
  assign n25965 = ~n25960 & n25964;
  assign n25966 = ~n25958 & n25965;
  assign n25967 = n25958 & ~n25965;
  assign n25968 = ~n25966 & ~n25967;
  assign n25969 = ~n25943 & ~n25968;
  assign n25970 = n25943 & n25968;
  assign n25971 = ~n25969 & ~n25970;
  assign n25972 = ~n25941 & n25971;
  assign n25973 = n25941 & ~n25971;
  assign n25974 = ~n25972 & ~n25973;
  assign n25975 = ~n25931 & n25974;
  assign n25976 = n25931 & ~n25974;
  assign n25977 = ~n25975 & ~n25976;
  assign n25978 = n86 & n21054;
  assign n25979 = n4420 & n21812;
  assign n25980 = n4600 & n21051;
  assign n25981 = n4615 & n21048;
  assign n25982 = ~n25978 & ~n25980;
  assign n25983 = ~n25981 & n25982;
  assign n25984 = ~n25979 & n25983;
  assign n25985 = pi26  & n25984;
  assign n25986 = ~pi26  & ~n25984;
  assign n25987 = ~n25985 & ~n25986;
  assign n25988 = n25977 & n25987;
  assign n25989 = ~n25977 & ~n25987;
  assign n25990 = ~n25988 & ~n25989;
  assign n25991 = ~n25930 & ~n25990;
  assign n25992 = n25930 & n25990;
  assign n25993 = ~n25991 & ~n25992;
  assign n25994 = ~n25928 & ~n25993;
  assign n25995 = n25928 & n25993;
  assign n25996 = ~n25994 & ~n25995;
  assign n25997 = ~n25674 & n25741;
  assign n25998 = ~n25748 & ~n25997;
  assign n25999 = n25996 & n25998;
  assign n26000 = ~n25996 & ~n25998;
  assign n26001 = ~n25999 & ~n26000;
  assign n26002 = n5240 & n21036;
  assign n26003 = n5241 & n22632;
  assign n26004 = n5853 & n21033;
  assign n26005 = n5866 & n21030;
  assign n26006 = ~n26002 & ~n26004;
  assign n26007 = ~n26005 & n26006;
  assign n26008 = ~n26003 & n26007;
  assign n26009 = pi20  & n26008;
  assign n26010 = ~pi20  & ~n26008;
  assign n26011 = ~n26009 & ~n26010;
  assign n26012 = n26001 & n26011;
  assign n26013 = ~n26001 & ~n26011;
  assign n26014 = ~n26012 & ~n26013;
  assign n26015 = ~n25918 & n26014;
  assign n26016 = n25918 & ~n26014;
  assign n26017 = ~n26015 & ~n26016;
  assign n26018 = ~n25915 & ~n26017;
  assign n26019 = n25915 & n26017;
  assign n26020 = ~n26018 & ~n26019;
  assign n26021 = n25905 & ~n26020;
  assign n26022 = ~n25905 & n26020;
  assign n26023 = ~n26021 & ~n26022;
  assign n26024 = n6630 & n21018;
  assign n26025 = n6631 & n23205;
  assign n26026 = n7238 & n21015;
  assign n26027 = n7262 & n21012;
  assign n26028 = ~n26024 & ~n26026;
  assign n26029 = ~n26027 & n26028;
  assign n26030 = ~n26025 & n26029;
  assign n26031 = pi14  & n26030;
  assign n26032 = ~pi14  & ~n26030;
  assign n26033 = ~n26031 & ~n26032;
  assign n26034 = n26023 & n26033;
  assign n26035 = ~n26023 & ~n26033;
  assign n26036 = ~n26034 & ~n26035;
  assign n26037 = ~n25904 & ~n26036;
  assign n26038 = n25904 & n26036;
  assign n26039 = ~n26037 & ~n26038;
  assign n26040 = ~n25902 & ~n26039;
  assign n26041 = n25902 & n26039;
  assign n26042 = ~n26040 & ~n26041;
  assign n26043 = ~n25648 & n25787;
  assign n26044 = ~n25794 & ~n26043;
  assign n26045 = n26042 & n26044;
  assign n26046 = ~n26042 & ~n26044;
  assign n26047 = ~n26045 & ~n26046;
  assign n26048 = n8250 & n21003;
  assign n26049 = n8251 & n24596;
  assign n26050 = n9016 & n21288;
  assign n26051 = n9040 & n24428;
  assign n26052 = ~n26048 & ~n26050;
  assign n26053 = ~n26051 & n26052;
  assign n26054 = ~n26049 & n26053;
  assign n26055 = pi8  & n26054;
  assign n26056 = ~pi8  & ~n26054;
  assign n26057 = ~n26055 & ~n26056;
  assign n26058 = n26047 & n26057;
  assign n26059 = ~n26047 & ~n26057;
  assign n26060 = ~n26058 & ~n26059;
  assign n26061 = ~n25892 & n26060;
  assign n26062 = n25892 & ~n26060;
  assign n26063 = ~n26061 & ~n26062;
  assign n26064 = ~n25889 & ~n26063;
  assign n26065 = n25889 & n26063;
  assign n26066 = ~n26064 & ~n26065;
  assign n26067 = n25879 & ~n26066;
  assign n26068 = ~n25879 & n26066;
  assign n26069 = ~n26067 & ~n26068;
  assign n26070 = n11055 & n25599;
  assign n26071 = ~n25855 & ~n25857;
  assign n26072 = n25834 & ~n25841;
  assign n26073 = ~n25845 & ~n26072;
  assign n26074 = ~n25830 & ~n25832;
  assign n26075 = n3821 & ~n26074;
  assign n26076 = ~n3821 & n26074;
  assign n26077 = ~n26075 & ~n26076;
  assign n26078 = n3692 & n13161;
  assign n26079 = n880 & ~n13781;
  assign n26080 = n748 & n13166;
  assign n26081 = n3694 & ~n12786;
  assign n26082 = ~n26080 & ~n26081;
  assign n26083 = ~n26078 & n26082;
  assign n26084 = ~n26079 & n26083;
  assign n26085 = n26077 & ~n26084;
  assign n26086 = ~n26077 & n26084;
  assign n26087 = ~n26085 & ~n26086;
  assign n26088 = n26073 & ~n26087;
  assign n26089 = ~n26073 & n26087;
  assign n26090 = ~n26088 & ~n26089;
  assign n26091 = ~n25848 & ~n25851;
  assign n26092 = ~n26090 & n26091;
  assign n26093 = n26090 & ~n26091;
  assign n26094 = ~n26092 & ~n26093;
  assign n26095 = n25853 & n26094;
  assign n26096 = ~n25853 & ~n26094;
  assign n26097 = ~n26095 & ~n26096;
  assign n26098 = ~n26071 & n26097;
  assign n26099 = n26071 & ~n26097;
  assign n26100 = ~n26098 & ~n26099;
  assign n26101 = n11056 & n26100;
  assign n26102 = n11661 & n25853;
  assign n26103 = n11672 & n26094;
  assign n26104 = ~n26070 & ~n26102;
  assign n26105 = ~n26103 & n26104;
  assign n26106 = ~n26101 & n26105;
  assign n26107 = pi2  & n26106;
  assign n26108 = ~pi2  & ~n26106;
  assign n26109 = ~n26107 & ~n26108;
  assign n26110 = n26069 & ~n26109;
  assign n26111 = ~n26069 & n26109;
  assign n26112 = ~n26110 & ~n26111;
  assign n26113 = ~n25878 & n26112;
  assign n26114 = n25878 & ~n26112;
  assign n26115 = ~n26113 & ~n26114;
  assign n26116 = n25875 & n26115;
  assign n26117 = ~n25875 & ~n26115;
  assign po3  = ~n26116 & ~n26117;
  assign n26119 = ~n26110 & ~n26113;
  assign n26120 = ~n26064 & ~n26068;
  assign n26121 = n75 & n24562;
  assign n26122 = n9491 & n25605;
  assign n26123 = n10469 & n25336;
  assign n26124 = n11031 & n25599;
  assign n26125 = ~n26121 & ~n26123;
  assign n26126 = ~n26124 & n26125;
  assign n26127 = ~n26122 & n26126;
  assign n26128 = ~pi5  & ~n26127;
  assign n26129 = pi5  & n26127;
  assign n26130 = ~n26128 & ~n26129;
  assign n26131 = n26047 & ~n26057;
  assign n26132 = ~n25892 & ~n26060;
  assign n26133 = ~n26131 & ~n26132;
  assign n26134 = n7430 & n21006;
  assign n26135 = n7431 & n23833;
  assign n26136 = n7869 & n20906;
  assign n26137 = n7895 & n21003;
  assign n26138 = ~n26134 & ~n26136;
  assign n26139 = ~n26137 & n26138;
  assign n26140 = ~n26135 & n26139;
  assign n26141 = ~pi11  & ~n26140;
  assign n26142 = pi11  & n26140;
  assign n26143 = ~n26141 & ~n26142;
  assign n26144 = n26023 & ~n26033;
  assign n26145 = ~n26037 & ~n26144;
  assign n26146 = ~n26018 & ~n26022;
  assign n26147 = n5982 & n21024;
  assign n26148 = n5983 & n23033;
  assign n26149 = n6323 & n21021;
  assign n26150 = n6336 & n21018;
  assign n26151 = ~n26147 & ~n26149;
  assign n26152 = ~n26150 & n26151;
  assign n26153 = ~n26148 & n26152;
  assign n26154 = ~pi17  & ~n26153;
  assign n26155 = pi17  & n26153;
  assign n26156 = ~n26154 & ~n26155;
  assign n26157 = n26001 & ~n26011;
  assign n26158 = ~n25918 & ~n26014;
  assign n26159 = ~n26157 & ~n26158;
  assign n26160 = n5044 & n21042;
  assign n26161 = n5045 & n22199;
  assign n26162 = n5109 & n21039;
  assign n26163 = n5130 & n21036;
  assign n26164 = ~n26160 & ~n26162;
  assign n26165 = ~n26163 & n26164;
  assign n26166 = ~n26161 & n26165;
  assign n26167 = ~pi23  & ~n26166;
  assign n26168 = pi23  & n26166;
  assign n26169 = ~n26167 & ~n26168;
  assign n26170 = n25977 & ~n25987;
  assign n26171 = ~n25991 & ~n26170;
  assign n26172 = ~n25972 & ~n25975;
  assign n26173 = n3810 & n21060;
  assign n26174 = n3886 & n21318;
  assign n26175 = n3884 & n21057;
  assign n26176 = n4380 & n21054;
  assign n26177 = ~n26173 & ~n26175;
  assign n26178 = ~n26176 & n26177;
  assign n26179 = ~n26174 & n26178;
  assign n26180 = pi29  & n26179;
  assign n26181 = ~pi29  & ~n26179;
  assign n26182 = ~n26180 & ~n26181;
  assign n26183 = ~n25958 & ~n25965;
  assign n26184 = ~n25969 & ~n26183;
  assign n26185 = ~n300 & ~n353;
  assign n26186 = ~n362 & ~n520;
  assign n26187 = n26185 & n26186;
  assign n26188 = n514 & n1354;
  assign n26189 = n2473 & n2891;
  assign n26190 = n6430 & n13512;
  assign n26191 = n26189 & n26190;
  assign n26192 = n26187 & n26188;
  assign n26193 = n26191 & n26192;
  assign n26194 = ~n639 & ~n814;
  assign n26195 = ~n902 & n26194;
  assign n26196 = n369 & n750;
  assign n26197 = n933 & n1171;
  assign n26198 = n1243 & n1294;
  assign n26199 = n2561 & n2889;
  assign n26200 = n26198 & n26199;
  assign n26201 = n26196 & n26197;
  assign n26202 = n1121 & n26195;
  assign n26203 = n2008 & n2186;
  assign n26204 = n26202 & n26203;
  assign n26205 = n26200 & n26201;
  assign n26206 = n2796 & n26205;
  assign n26207 = n26193 & n26204;
  assign n26208 = n26206 & n26207;
  assign n26209 = n4225 & n26208;
  assign n26210 = n4954 & n26209;
  assign n26211 = n3692 & n21066;
  assign n26212 = n880 & n21592;
  assign n26213 = n748 & n21069;
  assign n26214 = n3694 & n21063;
  assign n26215 = ~n26211 & ~n26213;
  assign n26216 = ~n26214 & n26215;
  assign n26217 = ~n26212 & n26216;
  assign n26218 = ~n26210 & n26217;
  assign n26219 = n26210 & ~n26217;
  assign n26220 = ~n26218 & ~n26219;
  assign n26221 = ~n26184 & ~n26220;
  assign n26222 = n26184 & n26220;
  assign n26223 = ~n26221 & ~n26222;
  assign n26224 = ~n26182 & n26223;
  assign n26225 = n26182 & ~n26223;
  assign n26226 = ~n26224 & ~n26225;
  assign n26227 = ~n26172 & n26226;
  assign n26228 = n26172 & ~n26226;
  assign n26229 = ~n26227 & ~n26228;
  assign n26230 = n86 & n21051;
  assign n26231 = n4420 & n21797;
  assign n26232 = n4600 & n21048;
  assign n26233 = n4615 & n21045;
  assign n26234 = ~n26230 & ~n26232;
  assign n26235 = ~n26233 & n26234;
  assign n26236 = ~n26231 & n26235;
  assign n26237 = pi26  & n26236;
  assign n26238 = ~pi26  & ~n26236;
  assign n26239 = ~n26237 & ~n26238;
  assign n26240 = n26229 & n26239;
  assign n26241 = ~n26229 & ~n26239;
  assign n26242 = ~n26240 & ~n26241;
  assign n26243 = ~n26171 & ~n26242;
  assign n26244 = n26171 & n26242;
  assign n26245 = ~n26243 & ~n26244;
  assign n26246 = ~n26169 & ~n26245;
  assign n26247 = n26169 & n26245;
  assign n26248 = ~n26246 & ~n26247;
  assign n26249 = ~n25928 & n25993;
  assign n26250 = ~n26000 & ~n26249;
  assign n26251 = n26248 & n26250;
  assign n26252 = ~n26248 & ~n26250;
  assign n26253 = ~n26251 & ~n26252;
  assign n26254 = n5240 & n21033;
  assign n26255 = n5241 & n22674;
  assign n26256 = n5853 & n21030;
  assign n26257 = n5866 & n21027;
  assign n26258 = ~n26254 & ~n26256;
  assign n26259 = ~n26257 & n26258;
  assign n26260 = ~n26255 & n26259;
  assign n26261 = pi20  & n26260;
  assign n26262 = ~pi20  & ~n26260;
  assign n26263 = ~n26261 & ~n26262;
  assign n26264 = n26253 & n26263;
  assign n26265 = ~n26253 & ~n26263;
  assign n26266 = ~n26264 & ~n26265;
  assign n26267 = ~n26159 & n26266;
  assign n26268 = n26159 & ~n26266;
  assign n26269 = ~n26267 & ~n26268;
  assign n26270 = ~n26156 & ~n26269;
  assign n26271 = n26156 & n26269;
  assign n26272 = ~n26270 & ~n26271;
  assign n26273 = n26146 & ~n26272;
  assign n26274 = ~n26146 & n26272;
  assign n26275 = ~n26273 & ~n26274;
  assign n26276 = n6630 & n21015;
  assign n26277 = n6631 & n23190;
  assign n26278 = n7238 & n21012;
  assign n26279 = n7262 & n21009;
  assign n26280 = ~n26276 & ~n26278;
  assign n26281 = ~n26279 & n26280;
  assign n26282 = ~n26277 & n26281;
  assign n26283 = pi14  & n26282;
  assign n26284 = ~pi14  & ~n26282;
  assign n26285 = ~n26283 & ~n26284;
  assign n26286 = n26275 & n26285;
  assign n26287 = ~n26275 & ~n26285;
  assign n26288 = ~n26286 & ~n26287;
  assign n26289 = ~n26145 & ~n26288;
  assign n26290 = n26145 & n26288;
  assign n26291 = ~n26289 & ~n26290;
  assign n26292 = ~n26143 & ~n26291;
  assign n26293 = n26143 & n26291;
  assign n26294 = ~n26292 & ~n26293;
  assign n26295 = ~n25902 & n26039;
  assign n26296 = ~n26046 & ~n26295;
  assign n26297 = n26294 & n26296;
  assign n26298 = ~n26294 & ~n26296;
  assign n26299 = ~n26297 & ~n26298;
  assign n26300 = n8250 & n21288;
  assign n26301 = n8251 & n24584;
  assign n26302 = n9016 & n24428;
  assign n26303 = n9040 & n24494;
  assign n26304 = ~n26300 & ~n26302;
  assign n26305 = ~n26303 & n26304;
  assign n26306 = ~n26301 & n26305;
  assign n26307 = pi8  & n26306;
  assign n26308 = ~pi8  & ~n26306;
  assign n26309 = ~n26307 & ~n26308;
  assign n26310 = n26299 & n26309;
  assign n26311 = ~n26299 & ~n26309;
  assign n26312 = ~n26310 & ~n26311;
  assign n26313 = ~n26133 & n26312;
  assign n26314 = n26133 & ~n26312;
  assign n26315 = ~n26313 & ~n26314;
  assign n26316 = ~n26130 & ~n26315;
  assign n26317 = n26130 & n26315;
  assign n26318 = ~n26316 & ~n26317;
  assign n26319 = n26120 & ~n26318;
  assign n26320 = ~n26120 & n26318;
  assign n26321 = ~n26319 & ~n26320;
  assign n26322 = n11055 & n25853;
  assign n26323 = ~n26095 & ~n26098;
  assign n26324 = n880 & ~n13280;
  assign n26325 = n748 & ~n13160;
  assign n26326 = ~n3692 & ~n3694;
  assign n26327 = ~n26325 & n26326;
  assign n26328 = ~n12786 & ~n26327;
  assign n26329 = ~n26324 & ~n26328;
  assign n26330 = n3821 & n26329;
  assign n26331 = ~n3821 & ~n26329;
  assign n26332 = ~n26330 & ~n26331;
  assign n26333 = ~n26075 & n26084;
  assign n26334 = ~n26076 & ~n26333;
  assign n26335 = n26332 & ~n26334;
  assign n26336 = ~n26332 & n26334;
  assign n26337 = ~n26335 & ~n26336;
  assign n26338 = ~n26089 & ~n26093;
  assign n26339 = ~n26337 & n26338;
  assign n26340 = n26337 & ~n26338;
  assign n26341 = ~n26339 & ~n26340;
  assign n26342 = ~n26094 & ~n26341;
  assign n26343 = n26094 & n26341;
  assign n26344 = ~n26342 & ~n26343;
  assign n26345 = ~n26323 & n26344;
  assign n26346 = n26323 & ~n26344;
  assign n26347 = ~n26345 & ~n26346;
  assign n26348 = n11056 & n26347;
  assign n26349 = n11661 & n26094;
  assign n26350 = n11672 & n26341;
  assign n26351 = ~n26322 & ~n26349;
  assign n26352 = ~n26350 & n26351;
  assign n26353 = ~n26348 & n26352;
  assign n26354 = pi2  & n26353;
  assign n26355 = ~pi2  & ~n26353;
  assign n26356 = ~n26354 & ~n26355;
  assign n26357 = n26321 & ~n26356;
  assign n26358 = ~n26321 & n26356;
  assign n26359 = ~n26357 & ~n26358;
  assign n26360 = ~n26119 & n26359;
  assign n26361 = n26119 & ~n26359;
  assign n26362 = ~n26360 & ~n26361;
  assign n26363 = n26116 & n26362;
  assign n26364 = ~n26116 & ~n26362;
  assign po4  = ~n26363 & ~n26364;
  assign n26366 = ~n26357 & ~n26360;
  assign n26367 = ~n26316 & ~n26320;
  assign n26368 = n75 & n25336;
  assign n26369 = n9491 & n25859;
  assign n26370 = n10469 & n25599;
  assign n26371 = n11031 & n25853;
  assign n26372 = ~n26368 & ~n26370;
  assign n26373 = ~n26371 & n26372;
  assign n26374 = ~n26369 & n26373;
  assign n26375 = ~pi5  & ~n26374;
  assign n26376 = pi5  & n26374;
  assign n26377 = ~n26375 & ~n26376;
  assign n26378 = n26299 & ~n26309;
  assign n26379 = ~n26133 & ~n26312;
  assign n26380 = ~n26378 & ~n26379;
  assign n26381 = n7430 & n20906;
  assign n26382 = n7431 & n21294;
  assign n26383 = n7869 & n21003;
  assign n26384 = n7895 & n21288;
  assign n26385 = ~n26381 & ~n26383;
  assign n26386 = ~n26384 & n26385;
  assign n26387 = ~n26382 & n26386;
  assign n26388 = ~pi11  & ~n26387;
  assign n26389 = pi11  & n26387;
  assign n26390 = ~n26388 & ~n26389;
  assign n26391 = n26275 & ~n26285;
  assign n26392 = ~n26289 & ~n26391;
  assign n26393 = ~n26270 & ~n26274;
  assign n26394 = n5982 & n21021;
  assign n26395 = n5983 & n23220;
  assign n26396 = n6323 & n21018;
  assign n26397 = n6336 & n21015;
  assign n26398 = ~n26394 & ~n26396;
  assign n26399 = ~n26397 & n26398;
  assign n26400 = ~n26395 & n26399;
  assign n26401 = ~pi17  & ~n26400;
  assign n26402 = pi17  & n26400;
  assign n26403 = ~n26401 & ~n26402;
  assign n26404 = n26253 & ~n26263;
  assign n26405 = ~n26159 & ~n26266;
  assign n26406 = ~n26404 & ~n26405;
  assign n26407 = n5044 & n21039;
  assign n26408 = n5045 & n22186;
  assign n26409 = n5109 & n21036;
  assign n26410 = n5130 & n21033;
  assign n26411 = ~n26407 & ~n26409;
  assign n26412 = ~n26410 & n26411;
  assign n26413 = ~n26408 & n26412;
  assign n26414 = ~pi23  & ~n26413;
  assign n26415 = pi23  & n26413;
  assign n26416 = ~n26414 & ~n26415;
  assign n26417 = n26229 & ~n26239;
  assign n26418 = ~n26243 & ~n26417;
  assign n26419 = ~n26224 & ~n26227;
  assign n26420 = n3810 & n21057;
  assign n26421 = n3886 & n21825;
  assign n26422 = n3884 & n21054;
  assign n26423 = n4380 & n21051;
  assign n26424 = ~n26420 & ~n26422;
  assign n26425 = ~n26423 & n26424;
  assign n26426 = ~n26421 & n26425;
  assign n26427 = pi29  & n26426;
  assign n26428 = ~pi29  & ~n26426;
  assign n26429 = ~n26427 & ~n26428;
  assign n26430 = ~n26210 & ~n26217;
  assign n26431 = ~n26221 & ~n26430;
  assign n26432 = ~n159 & ~n307;
  assign n26433 = ~n319 & ~n329;
  assign n26434 = ~n380 & ~n446;
  assign n26435 = ~n798 & n26434;
  assign n26436 = n26432 & n26433;
  assign n26437 = n900 & n12975;
  assign n26438 = n1134 & n1669;
  assign n26439 = n2449 & n26438;
  assign n26440 = n26436 & n26437;
  assign n26441 = n26435 & n26440;
  assign n26442 = n1116 & n26439;
  assign n26443 = n4085 & n26442;
  assign n26444 = n4021 & n26441;
  assign n26445 = n26443 & n26444;
  assign n26446 = n5744 & n26445;
  assign n26447 = n14984 & n26446;
  assign n26448 = n3692 & n21063;
  assign n26449 = n880 & n21631;
  assign n26450 = n748 & n21066;
  assign n26451 = n3694 & n21060;
  assign n26452 = ~n26448 & ~n26450;
  assign n26453 = ~n26451 & n26452;
  assign n26454 = ~n26449 & n26453;
  assign n26455 = ~n26447 & n26454;
  assign n26456 = n26447 & ~n26454;
  assign n26457 = ~n26455 & ~n26456;
  assign n26458 = ~n26431 & ~n26457;
  assign n26459 = n26431 & n26457;
  assign n26460 = ~n26458 & ~n26459;
  assign n26461 = ~n26429 & n26460;
  assign n26462 = n26429 & ~n26460;
  assign n26463 = ~n26461 & ~n26462;
  assign n26464 = ~n26419 & n26463;
  assign n26465 = n26419 & ~n26463;
  assign n26466 = ~n26464 & ~n26465;
  assign n26467 = n86 & n21048;
  assign n26468 = n4420 & n22049;
  assign n26469 = n4600 & n21045;
  assign n26470 = n4615 & n21042;
  assign n26471 = ~n26467 & ~n26469;
  assign n26472 = ~n26470 & n26471;
  assign n26473 = ~n26468 & n26472;
  assign n26474 = pi26  & n26473;
  assign n26475 = ~pi26  & ~n26473;
  assign n26476 = ~n26474 & ~n26475;
  assign n26477 = n26466 & n26476;
  assign n26478 = ~n26466 & ~n26476;
  assign n26479 = ~n26477 & ~n26478;
  assign n26480 = ~n26418 & ~n26479;
  assign n26481 = n26418 & n26479;
  assign n26482 = ~n26480 & ~n26481;
  assign n26483 = ~n26416 & ~n26482;
  assign n26484 = n26416 & n26482;
  assign n26485 = ~n26483 & ~n26484;
  assign n26486 = ~n26169 & n26245;
  assign n26487 = ~n26252 & ~n26486;
  assign n26488 = n26485 & n26487;
  assign n26489 = ~n26485 & ~n26487;
  assign n26490 = ~n26488 & ~n26489;
  assign n26491 = n5240 & n21030;
  assign n26492 = n5241 & n22654;
  assign n26493 = n5853 & n21027;
  assign n26494 = n5866 & n21024;
  assign n26495 = ~n26491 & ~n26493;
  assign n26496 = ~n26494 & n26495;
  assign n26497 = ~n26492 & n26496;
  assign n26498 = pi20  & n26497;
  assign n26499 = ~pi20  & ~n26497;
  assign n26500 = ~n26498 & ~n26499;
  assign n26501 = n26490 & n26500;
  assign n26502 = ~n26490 & ~n26500;
  assign n26503 = ~n26501 & ~n26502;
  assign n26504 = ~n26406 & n26503;
  assign n26505 = n26406 & ~n26503;
  assign n26506 = ~n26504 & ~n26505;
  assign n26507 = ~n26403 & ~n26506;
  assign n26508 = n26403 & n26506;
  assign n26509 = ~n26507 & ~n26508;
  assign n26510 = n26393 & ~n26509;
  assign n26511 = ~n26393 & n26509;
  assign n26512 = ~n26510 & ~n26511;
  assign n26513 = n6630 & n21012;
  assign n26514 = n6631 & n23812;
  assign n26515 = n7238 & n21009;
  assign n26516 = n7262 & n21006;
  assign n26517 = ~n26513 & ~n26515;
  assign n26518 = ~n26516 & n26517;
  assign n26519 = ~n26514 & n26518;
  assign n26520 = pi14  & n26519;
  assign n26521 = ~pi14  & ~n26519;
  assign n26522 = ~n26520 & ~n26521;
  assign n26523 = n26512 & n26522;
  assign n26524 = ~n26512 & ~n26522;
  assign n26525 = ~n26523 & ~n26524;
  assign n26526 = ~n26392 & ~n26525;
  assign n26527 = n26392 & n26525;
  assign n26528 = ~n26526 & ~n26527;
  assign n26529 = ~n26390 & ~n26528;
  assign n26530 = n26390 & n26528;
  assign n26531 = ~n26529 & ~n26530;
  assign n26532 = ~n26143 & n26291;
  assign n26533 = ~n26298 & ~n26532;
  assign n26534 = n26531 & n26533;
  assign n26535 = ~n26531 & ~n26533;
  assign n26536 = ~n26534 & ~n26535;
  assign n26537 = n8250 & n24428;
  assign n26538 = n8251 & n24568;
  assign n26539 = n9016 & n24494;
  assign n26540 = n9040 & n24562;
  assign n26541 = ~n26537 & ~n26539;
  assign n26542 = ~n26540 & n26541;
  assign n26543 = ~n26538 & n26542;
  assign n26544 = pi8  & n26543;
  assign n26545 = ~pi8  & ~n26543;
  assign n26546 = ~n26544 & ~n26545;
  assign n26547 = n26536 & n26546;
  assign n26548 = ~n26536 & ~n26546;
  assign n26549 = ~n26547 & ~n26548;
  assign n26550 = ~n26380 & n26549;
  assign n26551 = n26380 & ~n26549;
  assign n26552 = ~n26550 & ~n26551;
  assign n26553 = ~n26377 & ~n26552;
  assign n26554 = n26377 & n26552;
  assign n26555 = ~n26553 & ~n26554;
  assign n26556 = n26367 & ~n26555;
  assign n26557 = ~n26367 & n26555;
  assign n26558 = ~n26556 & ~n26557;
  assign n26559 = n11055 & n26094;
  assign n26560 = ~n26343 & ~n26345;
  assign n26561 = ~n26336 & ~n26340;
  assign n26562 = ~pi31  & n94;
  assign n26563 = ~n12786 & ~n26562;
  assign n26564 = n26330 & ~n26563;
  assign n26565 = ~n26330 & n26563;
  assign n26566 = ~n26564 & ~n26565;
  assign n26567 = n26561 & n26566;
  assign n26568 = ~n26561 & ~n26566;
  assign n26569 = ~n26567 & ~n26568;
  assign n26570 = n26341 & n26569;
  assign n26571 = ~n26341 & ~n26569;
  assign n26572 = ~n26570 & ~n26571;
  assign n26573 = ~n26560 & n26572;
  assign n26574 = n26560 & ~n26572;
  assign n26575 = ~n26573 & ~n26574;
  assign n26576 = n11056 & n26575;
  assign n26577 = n11661 & n26341;
  assign n26578 = n11672 & n26569;
  assign n26579 = ~n26559 & ~n26577;
  assign n26580 = ~n26578 & n26579;
  assign n26581 = ~n26576 & n26580;
  assign n26582 = pi2  & n26581;
  assign n26583 = ~pi2  & ~n26581;
  assign n26584 = ~n26582 & ~n26583;
  assign n26585 = n26558 & ~n26584;
  assign n26586 = ~n26558 & n26584;
  assign n26587 = ~n26585 & ~n26586;
  assign n26588 = ~n26366 & n26587;
  assign n26589 = n26366 & ~n26587;
  assign n26590 = ~n26588 & ~n26589;
  assign n26591 = n26363 & n26590;
  assign n26592 = ~n26363 & ~n26590;
  assign po5  = ~n26591 & ~n26592;
  assign n26594 = ~n26553 & ~n26557;
  assign n26595 = n75 & n25599;
  assign n26596 = n9491 & n26100;
  assign n26597 = n10469 & n25853;
  assign n26598 = n11031 & n26094;
  assign n26599 = ~n26595 & ~n26597;
  assign n26600 = ~n26598 & n26599;
  assign n26601 = ~n26596 & n26600;
  assign n26602 = ~pi5  & ~n26601;
  assign n26603 = pi5  & n26601;
  assign n26604 = ~n26602 & ~n26603;
  assign n26605 = n26536 & ~n26546;
  assign n26606 = ~n26380 & ~n26549;
  assign n26607 = ~n26605 & ~n26606;
  assign n26608 = n7430 & n21003;
  assign n26609 = n7431 & n24596;
  assign n26610 = n7869 & n21288;
  assign n26611 = n7895 & n24428;
  assign n26612 = ~n26608 & ~n26610;
  assign n26613 = ~n26611 & n26612;
  assign n26614 = ~n26609 & n26613;
  assign n26615 = ~pi11  & ~n26614;
  assign n26616 = pi11  & n26614;
  assign n26617 = ~n26615 & ~n26616;
  assign n26618 = n26512 & ~n26522;
  assign n26619 = ~n26526 & ~n26618;
  assign n26620 = n5982 & n21018;
  assign n26621 = n5983 & n23205;
  assign n26622 = n6323 & n21015;
  assign n26623 = n6336 & n21012;
  assign n26624 = ~n26620 & ~n26622;
  assign n26625 = ~n26623 & n26624;
  assign n26626 = ~n26621 & n26625;
  assign n26627 = ~pi17  & ~n26626;
  assign n26628 = pi17  & n26626;
  assign n26629 = ~n26627 & ~n26628;
  assign n26630 = n26490 & ~n26500;
  assign n26631 = ~n26406 & ~n26503;
  assign n26632 = ~n26630 & ~n26631;
  assign n26633 = n5044 & n21036;
  assign n26634 = n5045 & n22632;
  assign n26635 = n5109 & n21033;
  assign n26636 = n5130 & n21030;
  assign n26637 = ~n26633 & ~n26635;
  assign n26638 = ~n26636 & n26637;
  assign n26639 = ~n26634 & n26638;
  assign n26640 = ~pi23  & ~n26639;
  assign n26641 = pi23  & n26639;
  assign n26642 = ~n26640 & ~n26641;
  assign n26643 = n26466 & ~n26476;
  assign n26644 = ~n26480 & ~n26643;
  assign n26645 = ~n26461 & ~n26464;
  assign n26646 = n3810 & n21054;
  assign n26647 = n3886 & n21812;
  assign n26648 = n3884 & n21051;
  assign n26649 = n4380 & n21048;
  assign n26650 = ~n26646 & ~n26648;
  assign n26651 = ~n26649 & n26650;
  assign n26652 = ~n26647 & n26651;
  assign n26653 = pi29  & n26652;
  assign n26654 = ~pi29  & ~n26652;
  assign n26655 = ~n26653 & ~n26654;
  assign n26656 = ~n26447 & ~n26454;
  assign n26657 = ~n26458 & ~n26656;
  assign n26658 = ~n200 & ~n278;
  assign n26659 = n654 & n26658;
  assign n26660 = n790 & n2548;
  assign n26661 = n5490 & n26660;
  assign n26662 = n26659 & n26661;
  assign n26663 = ~n116 & ~n178;
  assign n26664 = ~n290 & ~n416;
  assign n26665 = ~n523 & ~n685;
  assign n26666 = n26664 & n26665;
  assign n26667 = n301 & n26663;
  assign n26668 = n354 & n434;
  assign n26669 = n750 & n933;
  assign n26670 = n1247 & n1492;
  assign n26671 = n2170 & n26670;
  assign n26672 = n26668 & n26669;
  assign n26673 = n26666 & n26667;
  assign n26674 = n26672 & n26673;
  assign n26675 = n13670 & n26671;
  assign n26676 = n25945 & n26675;
  assign n26677 = n26662 & n26674;
  assign n26678 = n26676 & n26677;
  assign n26679 = n3163 & n5484;
  assign n26680 = n14114 & n26679;
  assign n26681 = n26678 & n26680;
  assign n26682 = n3692 & n21060;
  assign n26683 = n880 & n21613;
  assign n26684 = n748 & n21063;
  assign n26685 = n3694 & n21057;
  assign n26686 = ~n26682 & ~n26684;
  assign n26687 = ~n26685 & n26686;
  assign n26688 = ~n26683 & n26687;
  assign n26689 = ~n26681 & n26688;
  assign n26690 = n26681 & ~n26688;
  assign n26691 = ~n26689 & ~n26690;
  assign n26692 = ~n26657 & ~n26691;
  assign n26693 = n26657 & n26691;
  assign n26694 = ~n26692 & ~n26693;
  assign n26695 = ~n26655 & n26694;
  assign n26696 = n26655 & ~n26694;
  assign n26697 = ~n26695 & ~n26696;
  assign n26698 = ~n26645 & n26697;
  assign n26699 = n26645 & ~n26697;
  assign n26700 = ~n26698 & ~n26699;
  assign n26701 = n86 & n21045;
  assign n26702 = n4420 & n22217;
  assign n26703 = n4600 & n21042;
  assign n26704 = n4615 & n21039;
  assign n26705 = ~n26701 & ~n26703;
  assign n26706 = ~n26704 & n26705;
  assign n26707 = ~n26702 & n26706;
  assign n26708 = pi26  & n26707;
  assign n26709 = ~pi26  & ~n26707;
  assign n26710 = ~n26708 & ~n26709;
  assign n26711 = n26700 & ~n26710;
  assign n26712 = ~n26700 & n26710;
  assign n26713 = ~n26711 & ~n26712;
  assign n26714 = ~n26644 & n26713;
  assign n26715 = n26644 & ~n26713;
  assign n26716 = ~n26714 & ~n26715;
  assign n26717 = ~n26642 & ~n26716;
  assign n26718 = n26642 & n26716;
  assign n26719 = ~n26717 & ~n26718;
  assign n26720 = ~n26416 & n26482;
  assign n26721 = ~n26489 & ~n26720;
  assign n26722 = n26719 & n26721;
  assign n26723 = ~n26719 & ~n26721;
  assign n26724 = ~n26722 & ~n26723;
  assign n26725 = n5240 & n21027;
  assign n26726 = n5241 & n21306;
  assign n26727 = n5853 & n21024;
  assign n26728 = n5866 & n21021;
  assign n26729 = ~n26725 & ~n26727;
  assign n26730 = ~n26728 & n26729;
  assign n26731 = ~n26726 & n26730;
  assign n26732 = pi20  & n26731;
  assign n26733 = ~pi20  & ~n26731;
  assign n26734 = ~n26732 & ~n26733;
  assign n26735 = n26724 & ~n26734;
  assign n26736 = ~n26724 & n26734;
  assign n26737 = ~n26735 & ~n26736;
  assign n26738 = ~n26632 & n26737;
  assign n26739 = n26632 & ~n26737;
  assign n26740 = ~n26738 & ~n26739;
  assign n26741 = ~n26629 & ~n26740;
  assign n26742 = n26629 & n26740;
  assign n26743 = ~n26741 & ~n26742;
  assign n26744 = ~n26507 & ~n26511;
  assign n26745 = n26743 & n26744;
  assign n26746 = ~n26743 & ~n26744;
  assign n26747 = ~n26745 & ~n26746;
  assign n26748 = n6630 & n21009;
  assign n26749 = n6631 & n23851;
  assign n26750 = n7238 & n21006;
  assign n26751 = n7262 & n20906;
  assign n26752 = ~n26748 & ~n26750;
  assign n26753 = ~n26751 & n26752;
  assign n26754 = ~n26749 & n26753;
  assign n26755 = pi14  & n26754;
  assign n26756 = ~pi14  & ~n26754;
  assign n26757 = ~n26755 & ~n26756;
  assign n26758 = n26747 & ~n26757;
  assign n26759 = ~n26747 & n26757;
  assign n26760 = ~n26758 & ~n26759;
  assign n26761 = ~n26619 & n26760;
  assign n26762 = n26619 & ~n26760;
  assign n26763 = ~n26761 & ~n26762;
  assign n26764 = ~n26617 & ~n26763;
  assign n26765 = n26617 & n26763;
  assign n26766 = ~n26764 & ~n26765;
  assign n26767 = ~n26390 & n26528;
  assign n26768 = ~n26535 & ~n26767;
  assign n26769 = n26766 & n26768;
  assign n26770 = ~n26766 & ~n26768;
  assign n26771 = ~n26769 & ~n26770;
  assign n26772 = n8250 & n24494;
  assign n26773 = n8251 & n25342;
  assign n26774 = n9016 & n24562;
  assign n26775 = n9040 & n25336;
  assign n26776 = ~n26772 & ~n26774;
  assign n26777 = ~n26775 & n26776;
  assign n26778 = ~n26773 & n26777;
  assign n26779 = pi8  & n26778;
  assign n26780 = ~pi8  & ~n26778;
  assign n26781 = ~n26779 & ~n26780;
  assign n26782 = n26771 & ~n26781;
  assign n26783 = ~n26771 & n26781;
  assign n26784 = ~n26782 & ~n26783;
  assign n26785 = ~n26607 & n26784;
  assign n26786 = n26607 & ~n26784;
  assign n26787 = ~n26785 & ~n26786;
  assign n26788 = ~n26604 & ~n26787;
  assign n26789 = n26604 & n26787;
  assign n26790 = ~n26788 & ~n26789;
  assign n26791 = n19514 & n26569;
  assign n26792 = n11055 & n26341;
  assign n26793 = ~n26570 & ~n26573;
  assign n26794 = n11056 & ~n26793;
  assign n26795 = ~n26791 & ~n26792;
  assign n26796 = ~n26794 & n26795;
  assign n26797 = pi2  & n26796;
  assign n26798 = ~pi2  & ~n26796;
  assign n26799 = ~n26797 & ~n26798;
  assign n26800 = ~n26790 & ~n26799;
  assign n26801 = n26790 & n26799;
  assign n26802 = ~n26800 & ~n26801;
  assign n26803 = n26594 & ~n26802;
  assign n26804 = ~n26594 & n26802;
  assign n26805 = ~n26803 & ~n26804;
  assign n26806 = ~n26585 & ~n26588;
  assign n26807 = ~n26805 & n26806;
  assign n26808 = n26805 & ~n26806;
  assign n26809 = ~n26807 & ~n26808;
  assign n26810 = n26591 & n26809;
  assign n26811 = ~n26591 & ~n26809;
  assign po6  = ~n26810 & ~n26811;
  assign n26813 = ~n26604 & n26787;
  assign n26814 = ~n26800 & ~n26813;
  assign n26815 = ~n26782 & ~n26785;
  assign n26816 = ~n26617 & n26763;
  assign n26817 = ~n26770 & ~n26816;
  assign n26818 = ~n26758 & ~n26761;
  assign n26819 = ~n26629 & n26740;
  assign n26820 = ~n26746 & ~n26819;
  assign n26821 = ~n26735 & ~n26738;
  assign n26822 = ~n26642 & n26716;
  assign n26823 = ~n26723 & ~n26822;
  assign n26824 = ~n26711 & ~n26714;
  assign n26825 = ~n26695 & ~n26698;
  assign n26826 = ~n26681 & ~n26688;
  assign n26827 = ~n26692 & ~n26826;
  assign n26828 = ~n111 & ~n183;
  assign n26829 = ~n422 & ~n751;
  assign n26830 = n26828 & n26829;
  assign n26831 = n357 & n1186;
  assign n26832 = n3121 & n13513;
  assign n26833 = n13500 & n26832;
  assign n26834 = n26830 & n26831;
  assign n26835 = n2876 & n12690;
  assign n26836 = n26834 & n26835;
  assign n26837 = n7084 & n26833;
  assign n26838 = n26836 & n26837;
  assign n26839 = n2694 & n3629;
  assign n26840 = n12823 & n26839;
  assign n26841 = n26838 & n26840;
  assign n26842 = n3218 & n26841;
  assign n26843 = n837 & n26842;
  assign n26844 = pi2  & ~n26569;
  assign n26845 = n14099 & n26569;
  assign n26846 = ~n26844 & ~n26845;
  assign n26847 = n26843 & n26846;
  assign n26848 = ~n26843 & ~n26846;
  assign n26849 = ~n26847 & ~n26848;
  assign n26850 = n748 & n21060;
  assign n26851 = n880 & n21318;
  assign n26852 = n3692 & n21057;
  assign n26853 = n3694 & n21054;
  assign n26854 = ~n26850 & ~n26852;
  assign n26855 = ~n26853 & n26854;
  assign n26856 = ~n26851 & n26855;
  assign n26857 = ~n26849 & n26856;
  assign n26858 = n26849 & ~n26856;
  assign n26859 = ~n26857 & ~n26858;
  assign n26860 = n26827 & ~n26859;
  assign n26861 = ~n26827 & n26859;
  assign n26862 = ~n26860 & ~n26861;
  assign n26863 = n3810 & n21051;
  assign n26864 = n3886 & n21797;
  assign n26865 = n3884 & n21048;
  assign n26866 = n4380 & n21045;
  assign n26867 = ~n26863 & ~n26865;
  assign n26868 = ~n26866 & n26867;
  assign n26869 = ~n26864 & n26868;
  assign n26870 = pi29  & n26869;
  assign n26871 = ~pi29  & ~n26869;
  assign n26872 = ~n26870 & ~n26871;
  assign n26873 = n26862 & ~n26872;
  assign n26874 = ~n26862 & n26872;
  assign n26875 = ~n26873 & ~n26874;
  assign n26876 = ~n26825 & n26875;
  assign n26877 = n26825 & ~n26875;
  assign n26878 = ~n26876 & ~n26877;
  assign n26879 = n86 & n21042;
  assign n26880 = n4420 & n22199;
  assign n26881 = n4600 & n21039;
  assign n26882 = n4615 & n21036;
  assign n26883 = ~n26879 & ~n26881;
  assign n26884 = ~n26882 & n26883;
  assign n26885 = ~n26880 & n26884;
  assign n26886 = pi26  & n26885;
  assign n26887 = ~pi26  & ~n26885;
  assign n26888 = ~n26886 & ~n26887;
  assign n26889 = n26878 & ~n26888;
  assign n26890 = ~n26878 & n26888;
  assign n26891 = ~n26889 & ~n26890;
  assign n26892 = n26824 & ~n26891;
  assign n26893 = ~n26824 & n26891;
  assign n26894 = ~n26892 & ~n26893;
  assign n26895 = n5044 & n21033;
  assign n26896 = n5045 & n22674;
  assign n26897 = n5109 & n21030;
  assign n26898 = n5130 & n21027;
  assign n26899 = ~n26895 & ~n26897;
  assign n26900 = ~n26898 & n26899;
  assign n26901 = ~n26896 & n26900;
  assign n26902 = pi23  & n26901;
  assign n26903 = ~pi23  & ~n26901;
  assign n26904 = ~n26902 & ~n26903;
  assign n26905 = n26894 & ~n26904;
  assign n26906 = ~n26894 & n26904;
  assign n26907 = ~n26905 & ~n26906;
  assign n26908 = n26823 & ~n26907;
  assign n26909 = ~n26823 & n26907;
  assign n26910 = ~n26908 & ~n26909;
  assign n26911 = n5240 & n21024;
  assign n26912 = n5241 & n23033;
  assign n26913 = n5853 & n21021;
  assign n26914 = n5866 & n21018;
  assign n26915 = ~n26911 & ~n26913;
  assign n26916 = ~n26914 & n26915;
  assign n26917 = ~n26912 & n26916;
  assign n26918 = pi20  & n26917;
  assign n26919 = ~pi20  & ~n26917;
  assign n26920 = ~n26918 & ~n26919;
  assign n26921 = n26910 & ~n26920;
  assign n26922 = ~n26910 & n26920;
  assign n26923 = ~n26921 & ~n26922;
  assign n26924 = n26821 & ~n26923;
  assign n26925 = ~n26821 & n26923;
  assign n26926 = ~n26924 & ~n26925;
  assign n26927 = n5982 & n21015;
  assign n26928 = n5983 & n23190;
  assign n26929 = n6323 & n21012;
  assign n26930 = n6336 & n21009;
  assign n26931 = ~n26927 & ~n26929;
  assign n26932 = ~n26930 & n26931;
  assign n26933 = ~n26928 & n26932;
  assign n26934 = pi17  & n26933;
  assign n26935 = ~pi17  & ~n26933;
  assign n26936 = ~n26934 & ~n26935;
  assign n26937 = n26926 & ~n26936;
  assign n26938 = ~n26926 & n26936;
  assign n26939 = ~n26937 & ~n26938;
  assign n26940 = n26820 & ~n26939;
  assign n26941 = ~n26820 & n26939;
  assign n26942 = ~n26940 & ~n26941;
  assign n26943 = n6630 & n21006;
  assign n26944 = n6631 & n23833;
  assign n26945 = n7238 & n20906;
  assign n26946 = n7262 & n21003;
  assign n26947 = ~n26943 & ~n26945;
  assign n26948 = ~n26946 & n26947;
  assign n26949 = ~n26944 & n26948;
  assign n26950 = pi14  & n26949;
  assign n26951 = ~pi14  & ~n26949;
  assign n26952 = ~n26950 & ~n26951;
  assign n26953 = n26942 & ~n26952;
  assign n26954 = ~n26942 & n26952;
  assign n26955 = ~n26953 & ~n26954;
  assign n26956 = n26818 & ~n26955;
  assign n26957 = ~n26818 & n26955;
  assign n26958 = ~n26956 & ~n26957;
  assign n26959 = n7430 & n21288;
  assign n26960 = n7431 & n24584;
  assign n26961 = n7869 & n24428;
  assign n26962 = n7895 & n24494;
  assign n26963 = ~n26959 & ~n26961;
  assign n26964 = ~n26962 & n26963;
  assign n26965 = ~n26960 & n26964;
  assign n26966 = pi11  & n26965;
  assign n26967 = ~pi11  & ~n26965;
  assign n26968 = ~n26966 & ~n26967;
  assign n26969 = n26958 & ~n26968;
  assign n26970 = ~n26958 & n26968;
  assign n26971 = ~n26969 & ~n26970;
  assign n26972 = n26817 & ~n26971;
  assign n26973 = ~n26817 & n26971;
  assign n26974 = ~n26972 & ~n26973;
  assign n26975 = n8250 & n24562;
  assign n26976 = n8251 & n25605;
  assign n26977 = n9016 & n25336;
  assign n26978 = n9040 & n25599;
  assign n26979 = ~n26975 & ~n26977;
  assign n26980 = ~n26978 & n26979;
  assign n26981 = ~n26976 & n26980;
  assign n26982 = pi8  & n26981;
  assign n26983 = ~pi8  & ~n26981;
  assign n26984 = ~n26982 & ~n26983;
  assign n26985 = n26974 & ~n26984;
  assign n26986 = ~n26974 & n26984;
  assign n26987 = ~n26985 & ~n26986;
  assign n26988 = n26815 & ~n26987;
  assign n26989 = ~n26815 & n26987;
  assign n26990 = ~n26988 & ~n26989;
  assign n26991 = n75 & n25853;
  assign n26992 = n9491 & n26347;
  assign n26993 = n10469 & n26094;
  assign n26994 = n11031 & n26341;
  assign n26995 = ~n26991 & ~n26993;
  assign n26996 = ~n26994 & n26995;
  assign n26997 = ~n26992 & n26996;
  assign n26998 = pi5  & n26997;
  assign n26999 = ~pi5  & ~n26997;
  assign n27000 = ~n26998 & ~n26999;
  assign n27001 = n26990 & ~n27000;
  assign n27002 = ~n26990 & n27000;
  assign n27003 = ~n27001 & ~n27002;
  assign n27004 = n26814 & ~n27003;
  assign n27005 = ~n26814 & n27003;
  assign n27006 = ~n27004 & ~n27005;
  assign n27007 = ~n26804 & ~n26808;
  assign n27008 = ~n27006 & n27007;
  assign n27009 = n27006 & ~n27007;
  assign n27010 = ~n27008 & ~n27009;
  assign n27011 = n26810 & n27010;
  assign n27012 = ~n26810 & ~n27010;
  assign po7  = ~n27011 & ~n27012;
  assign n27014 = ~n116 & ~n415;
  assign n27015 = ~n1002 & n27014;
  assign n27016 = n799 & n27015;
  assign n27017 = n15079 & n27016;
  assign n27018 = ~n162 & ~n283;
  assign n27019 = ~n330 & ~n532;
  assign n27020 = n27018 & n27019;
  assign n27021 = n567 & n644;
  assign n27022 = n1858 & n1913;
  assign n27023 = n2234 & n2283;
  assign n27024 = n2608 & n3128;
  assign n27025 = n3325 & n4063;
  assign n27026 = n27024 & n27025;
  assign n27027 = n27022 & n27023;
  assign n27028 = n27020 & n27021;
  assign n27029 = n22547 & n27028;
  assign n27030 = n27026 & n27027;
  assign n27031 = n27029 & n27030;
  assign n27032 = n2166 & n27017;
  assign n27033 = n27031 & n27032;
  assign n27034 = n2867 & n27033;
  assign n27035 = n15054 & n27034;
  assign n27036 = ~n26846 & ~n27035;
  assign n27037 = n26846 & n27035;
  assign n27038 = ~n27036 & ~n27037;
  assign n27039 = ~n26847 & ~n26856;
  assign n27040 = ~n26848 & ~n27039;
  assign n27041 = n27038 & ~n27040;
  assign n27042 = ~n27038 & n27040;
  assign n27043 = ~n27041 & ~n27042;
  assign n27044 = n748 & n21057;
  assign n27045 = n880 & n21825;
  assign n27046 = n3692 & n21054;
  assign n27047 = n3694 & n21051;
  assign n27048 = ~n27044 & ~n27046;
  assign n27049 = ~n27047 & n27048;
  assign n27050 = ~n27045 & n27049;
  assign n27051 = n27043 & n27050;
  assign n27052 = ~n27043 & ~n27050;
  assign n27053 = ~n27051 & ~n27052;
  assign n27054 = ~n26861 & ~n26873;
  assign n27055 = n27053 & n27054;
  assign n27056 = ~n27053 & ~n27054;
  assign n27057 = ~n27055 & ~n27056;
  assign n27058 = n3810 & n21048;
  assign n27059 = n3886 & n22049;
  assign n27060 = n3884 & n21045;
  assign n27061 = n4380 & n21042;
  assign n27062 = ~n27058 & ~n27060;
  assign n27063 = ~n27061 & n27062;
  assign n27064 = ~n27059 & n27063;
  assign n27065 = pi29  & n27064;
  assign n27066 = ~pi29  & ~n27064;
  assign n27067 = ~n27065 & ~n27066;
  assign n27068 = n27057 & n27067;
  assign n27069 = ~n27057 & ~n27067;
  assign n27070 = ~n27068 & ~n27069;
  assign n27071 = n86 & n21039;
  assign n27072 = n4420 & n22186;
  assign n27073 = n4600 & n21036;
  assign n27074 = n4615 & n21033;
  assign n27075 = ~n27071 & ~n27073;
  assign n27076 = ~n27074 & n27075;
  assign n27077 = ~n27072 & n27076;
  assign n27078 = pi26  & n27077;
  assign n27079 = ~pi26  & ~n27077;
  assign n27080 = ~n27078 & ~n27079;
  assign n27081 = ~n27070 & n27080;
  assign n27082 = n27070 & ~n27080;
  assign n27083 = ~n27081 & ~n27082;
  assign n27084 = ~n26876 & n26888;
  assign n27085 = ~n26877 & ~n27084;
  assign n27086 = n27083 & ~n27085;
  assign n27087 = ~n27083 & n27085;
  assign n27088 = ~n27086 & ~n27087;
  assign n27089 = n5044 & n21030;
  assign n27090 = n5045 & n22654;
  assign n27091 = n5109 & n21027;
  assign n27092 = n5130 & n21024;
  assign n27093 = ~n27089 & ~n27091;
  assign n27094 = ~n27092 & n27093;
  assign n27095 = ~n27090 & n27094;
  assign n27096 = pi23  & n27095;
  assign n27097 = ~pi23  & ~n27095;
  assign n27098 = ~n27096 & ~n27097;
  assign n27099 = n27088 & ~n27098;
  assign n27100 = ~n27088 & n27098;
  assign n27101 = ~n27099 & ~n27100;
  assign n27102 = ~n26893 & n26904;
  assign n27103 = ~n26892 & ~n27102;
  assign n27104 = ~n27101 & ~n27103;
  assign n27105 = n27101 & n27103;
  assign n27106 = ~n27104 & ~n27105;
  assign n27107 = n5240 & n21021;
  assign n27108 = n5241 & n23220;
  assign n27109 = n5853 & n21018;
  assign n27110 = n5866 & n21015;
  assign n27111 = ~n27107 & ~n27109;
  assign n27112 = ~n27110 & n27111;
  assign n27113 = ~n27108 & n27112;
  assign n27114 = pi20  & n27113;
  assign n27115 = ~pi20  & ~n27113;
  assign n27116 = ~n27114 & ~n27115;
  assign n27117 = n27106 & ~n27116;
  assign n27118 = ~n27106 & n27116;
  assign n27119 = ~n27117 & ~n27118;
  assign n27120 = ~n26909 & n26920;
  assign n27121 = ~n26908 & ~n27120;
  assign n27122 = ~n27119 & ~n27121;
  assign n27123 = n27119 & n27121;
  assign n27124 = ~n27122 & ~n27123;
  assign n27125 = n5982 & n21012;
  assign n27126 = n5983 & n23812;
  assign n27127 = n6323 & n21009;
  assign n27128 = n6336 & n21006;
  assign n27129 = ~n27125 & ~n27127;
  assign n27130 = ~n27128 & n27129;
  assign n27131 = ~n27126 & n27130;
  assign n27132 = pi17  & n27131;
  assign n27133 = ~pi17  & ~n27131;
  assign n27134 = ~n27132 & ~n27133;
  assign n27135 = n27124 & ~n27134;
  assign n27136 = ~n27124 & n27134;
  assign n27137 = ~n27135 & ~n27136;
  assign n27138 = ~n26925 & n26936;
  assign n27139 = ~n26924 & ~n27138;
  assign n27140 = ~n27137 & ~n27139;
  assign n27141 = n27137 & n27139;
  assign n27142 = ~n27140 & ~n27141;
  assign n27143 = n6630 & n20906;
  assign n27144 = n6631 & n21294;
  assign n27145 = n7238 & n21003;
  assign n27146 = n7262 & n21288;
  assign n27147 = ~n27143 & ~n27145;
  assign n27148 = ~n27146 & n27147;
  assign n27149 = ~n27144 & n27148;
  assign n27150 = pi14  & n27149;
  assign n27151 = ~pi14  & ~n27149;
  assign n27152 = ~n27150 & ~n27151;
  assign n27153 = n27142 & ~n27152;
  assign n27154 = ~n27142 & n27152;
  assign n27155 = ~n27153 & ~n27154;
  assign n27156 = ~n26941 & n26952;
  assign n27157 = ~n26940 & ~n27156;
  assign n27158 = ~n27155 & ~n27157;
  assign n27159 = n27155 & n27157;
  assign n27160 = ~n27158 & ~n27159;
  assign n27161 = n7430 & n24428;
  assign n27162 = n7431 & n24568;
  assign n27163 = n7869 & n24494;
  assign n27164 = n7895 & n24562;
  assign n27165 = ~n27161 & ~n27163;
  assign n27166 = ~n27164 & n27165;
  assign n27167 = ~n27162 & n27166;
  assign n27168 = pi11  & n27167;
  assign n27169 = ~pi11  & ~n27167;
  assign n27170 = ~n27168 & ~n27169;
  assign n27171 = n27160 & ~n27170;
  assign n27172 = ~n27160 & n27170;
  assign n27173 = ~n27171 & ~n27172;
  assign n27174 = ~n26957 & n26968;
  assign n27175 = ~n26956 & ~n27174;
  assign n27176 = ~n27173 & ~n27175;
  assign n27177 = n27173 & n27175;
  assign n27178 = ~n27176 & ~n27177;
  assign n27179 = n8250 & n25336;
  assign n27180 = n8251 & n25859;
  assign n27181 = n9016 & n25599;
  assign n27182 = n9040 & n25853;
  assign n27183 = ~n27179 & ~n27181;
  assign n27184 = ~n27182 & n27183;
  assign n27185 = ~n27180 & n27184;
  assign n27186 = pi8  & n27185;
  assign n27187 = ~pi8  & ~n27185;
  assign n27188 = ~n27186 & ~n27187;
  assign n27189 = n27178 & ~n27188;
  assign n27190 = ~n27178 & n27188;
  assign n27191 = ~n27189 & ~n27190;
  assign n27192 = ~n26973 & n26984;
  assign n27193 = ~n26972 & ~n27192;
  assign n27194 = ~n27191 & ~n27193;
  assign n27195 = n27191 & n27193;
  assign n27196 = ~n27194 & ~n27195;
  assign n27197 = n75 & n26094;
  assign n27198 = n9491 & n26575;
  assign n27199 = n10469 & n26341;
  assign n27200 = n11031 & n26569;
  assign n27201 = ~n27197 & ~n27199;
  assign n27202 = ~n27200 & n27201;
  assign n27203 = ~n27198 & n27202;
  assign n27204 = pi5  & n27203;
  assign n27205 = ~pi5  & ~n27203;
  assign n27206 = ~n27204 & ~n27205;
  assign n27207 = n27196 & ~n27206;
  assign n27208 = ~n27196 & n27206;
  assign n27209 = ~n27207 & ~n27208;
  assign n27210 = ~n26989 & n27000;
  assign n27211 = ~n26988 & ~n27210;
  assign n27212 = ~n27209 & ~n27211;
  assign n27213 = n27209 & n27211;
  assign n27214 = ~n27212 & ~n27213;
  assign n27215 = ~n27005 & ~n27009;
  assign n27216 = ~n27214 & n27215;
  assign n27217 = n27214 & ~n27215;
  assign n27218 = ~n27216 & ~n27217;
  assign n27219 = n27011 & n27218;
  assign n27220 = ~n27011 & ~n27218;
  assign po8  = ~n27219 & ~n27220;
  assign n27222 = ~n14143 & n26569;
  assign n27223 = n75 & n26341;
  assign n27224 = n9491 & ~n26793;
  assign n27225 = ~n27222 & ~n27223;
  assign n27226 = ~n27224 & n27225;
  assign n27227 = pi5  & n27226;
  assign n27228 = ~pi5  & ~n27226;
  assign n27229 = ~n27227 & ~n27228;
  assign n27230 = ~n27177 & n27188;
  assign n27231 = ~n27176 & ~n27230;
  assign n27232 = ~n27229 & n27231;
  assign n27233 = n27229 & ~n27231;
  assign n27234 = ~n27232 & ~n27233;
  assign n27235 = ~n27036 & ~n27041;
  assign n27236 = ~n170 & ~n525;
  assign n27237 = ~n648 & ~n721;
  assign n27238 = ~n894 & n27237;
  assign n27239 = n749 & n27236;
  assign n27240 = n1012 & n2024;
  assign n27241 = n3122 & n3459;
  assign n27242 = n27240 & n27241;
  assign n27243 = n27238 & n27239;
  assign n27244 = n418 & n27243;
  assign n27245 = n4037 & n27242;
  assign n27246 = n14354 & n27245;
  assign n27247 = n1619 & n27244;
  assign n27248 = n5663 & n27247;
  assign n27249 = n27246 & n27248;
  assign n27250 = n2929 & n27249;
  assign n27251 = n1811 & n27250;
  assign n27252 = ~n26846 & ~n27251;
  assign n27253 = n26846 & n27251;
  assign n27254 = ~n27252 & ~n27253;
  assign n27255 = ~n27235 & n27254;
  assign n27256 = n27235 & ~n27254;
  assign n27257 = ~n27255 & ~n27256;
  assign n27258 = n748 & n21054;
  assign n27259 = n880 & n21812;
  assign n27260 = n3692 & n21051;
  assign n27261 = n3694 & n21048;
  assign n27262 = ~n27258 & ~n27260;
  assign n27263 = ~n27261 & n27262;
  assign n27264 = ~n27259 & n27263;
  assign n27265 = n27257 & n27264;
  assign n27266 = ~n27257 & ~n27264;
  assign n27267 = ~n27265 & ~n27266;
  assign n27268 = n27043 & ~n27050;
  assign n27269 = ~n27056 & ~n27268;
  assign n27270 = n27267 & n27269;
  assign n27271 = ~n27267 & ~n27269;
  assign n27272 = ~n27270 & ~n27271;
  assign n27273 = n3810 & n21045;
  assign n27274 = n3886 & n22217;
  assign n27275 = n3884 & n21042;
  assign n27276 = n4380 & n21039;
  assign n27277 = ~n27273 & ~n27275;
  assign n27278 = ~n27276 & n27277;
  assign n27279 = ~n27274 & n27278;
  assign n27280 = pi29  & n27279;
  assign n27281 = ~pi29  & ~n27279;
  assign n27282 = ~n27280 & ~n27281;
  assign n27283 = n27272 & n27282;
  assign n27284 = ~n27272 & ~n27282;
  assign n27285 = ~n27283 & ~n27284;
  assign n27286 = n86 & n21036;
  assign n27287 = n4420 & n22632;
  assign n27288 = n4600 & n21033;
  assign n27289 = n4615 & n21030;
  assign n27290 = ~n27286 & ~n27288;
  assign n27291 = ~n27289 & n27290;
  assign n27292 = ~n27287 & n27291;
  assign n27293 = pi26  & n27292;
  assign n27294 = ~pi26  & ~n27292;
  assign n27295 = ~n27293 & ~n27294;
  assign n27296 = ~n27285 & n27295;
  assign n27297 = n27285 & ~n27295;
  assign n27298 = ~n27296 & ~n27297;
  assign n27299 = n27057 & ~n27067;
  assign n27300 = ~n27070 & ~n27080;
  assign n27301 = ~n27299 & ~n27300;
  assign n27302 = n27298 & n27301;
  assign n27303 = ~n27298 & ~n27301;
  assign n27304 = ~n27302 & ~n27303;
  assign n27305 = n5044 & n21027;
  assign n27306 = n5045 & n21306;
  assign n27307 = n5109 & n21024;
  assign n27308 = n5130 & n21021;
  assign n27309 = ~n27305 & ~n27307;
  assign n27310 = ~n27308 & n27309;
  assign n27311 = ~n27306 & n27310;
  assign n27312 = pi23  & n27311;
  assign n27313 = ~pi23  & ~n27311;
  assign n27314 = ~n27312 & ~n27313;
  assign n27315 = n27304 & ~n27314;
  assign n27316 = ~n27304 & n27314;
  assign n27317 = ~n27315 & ~n27316;
  assign n27318 = ~n27087 & n27098;
  assign n27319 = ~n27086 & ~n27318;
  assign n27320 = ~n27317 & ~n27319;
  assign n27321 = n27317 & n27319;
  assign n27322 = ~n27320 & ~n27321;
  assign n27323 = n5240 & n21018;
  assign n27324 = n5241 & n23205;
  assign n27325 = n5853 & n21015;
  assign n27326 = n5866 & n21012;
  assign n27327 = ~n27323 & ~n27325;
  assign n27328 = ~n27326 & n27327;
  assign n27329 = ~n27324 & n27328;
  assign n27330 = pi20  & n27329;
  assign n27331 = ~pi20  & ~n27329;
  assign n27332 = ~n27330 & ~n27331;
  assign n27333 = n27322 & ~n27332;
  assign n27334 = ~n27322 & n27332;
  assign n27335 = ~n27333 & ~n27334;
  assign n27336 = ~n27105 & n27116;
  assign n27337 = ~n27104 & ~n27336;
  assign n27338 = ~n27335 & ~n27337;
  assign n27339 = n27335 & n27337;
  assign n27340 = ~n27338 & ~n27339;
  assign n27341 = n5982 & n21009;
  assign n27342 = n5983 & n23851;
  assign n27343 = n6323 & n21006;
  assign n27344 = n6336 & n20906;
  assign n27345 = ~n27341 & ~n27343;
  assign n27346 = ~n27344 & n27345;
  assign n27347 = ~n27342 & n27346;
  assign n27348 = pi17  & n27347;
  assign n27349 = ~pi17  & ~n27347;
  assign n27350 = ~n27348 & ~n27349;
  assign n27351 = n27340 & ~n27350;
  assign n27352 = ~n27340 & n27350;
  assign n27353 = ~n27351 & ~n27352;
  assign n27354 = ~n27123 & n27134;
  assign n27355 = ~n27122 & ~n27354;
  assign n27356 = ~n27353 & ~n27355;
  assign n27357 = n27353 & n27355;
  assign n27358 = ~n27356 & ~n27357;
  assign n27359 = n6630 & n21003;
  assign n27360 = n6631 & n24596;
  assign n27361 = n7238 & n21288;
  assign n27362 = n7262 & n24428;
  assign n27363 = ~n27359 & ~n27361;
  assign n27364 = ~n27362 & n27363;
  assign n27365 = ~n27360 & n27364;
  assign n27366 = pi14  & n27365;
  assign n27367 = ~pi14  & ~n27365;
  assign n27368 = ~n27366 & ~n27367;
  assign n27369 = n27358 & ~n27368;
  assign n27370 = ~n27358 & n27368;
  assign n27371 = ~n27369 & ~n27370;
  assign n27372 = ~n27141 & n27152;
  assign n27373 = ~n27140 & ~n27372;
  assign n27374 = ~n27371 & ~n27373;
  assign n27375 = n27371 & n27373;
  assign n27376 = ~n27374 & ~n27375;
  assign n27377 = n7430 & n24494;
  assign n27378 = n7431 & n25342;
  assign n27379 = n7869 & n24562;
  assign n27380 = n7895 & n25336;
  assign n27381 = ~n27377 & ~n27379;
  assign n27382 = ~n27380 & n27381;
  assign n27383 = ~n27378 & n27382;
  assign n27384 = pi11  & n27383;
  assign n27385 = ~pi11  & ~n27383;
  assign n27386 = ~n27384 & ~n27385;
  assign n27387 = n27376 & ~n27386;
  assign n27388 = ~n27376 & n27386;
  assign n27389 = ~n27387 & ~n27388;
  assign n27390 = ~n27159 & n27170;
  assign n27391 = ~n27158 & ~n27390;
  assign n27392 = ~n27389 & ~n27391;
  assign n27393 = n27389 & n27391;
  assign n27394 = ~n27392 & ~n27393;
  assign n27395 = n8250 & n25599;
  assign n27396 = n8251 & n26100;
  assign n27397 = n9016 & n25853;
  assign n27398 = n9040 & n26094;
  assign n27399 = ~n27395 & ~n27397;
  assign n27400 = ~n27398 & n27399;
  assign n27401 = ~n27396 & n27400;
  assign n27402 = pi8  & n27401;
  assign n27403 = ~pi8  & ~n27401;
  assign n27404 = ~n27402 & ~n27403;
  assign n27405 = n27394 & ~n27404;
  assign n27406 = ~n27394 & n27404;
  assign n27407 = ~n27405 & ~n27406;
  assign n27408 = n27234 & n27407;
  assign n27409 = ~n27234 & ~n27407;
  assign n27410 = ~n27408 & ~n27409;
  assign n27411 = ~n27195 & n27206;
  assign n27412 = ~n27194 & ~n27411;
  assign n27413 = ~n27410 & ~n27412;
  assign n27414 = n27410 & n27412;
  assign n27415 = ~n27413 & ~n27414;
  assign n27416 = ~n27213 & ~n27217;
  assign n27417 = ~n27415 & n27416;
  assign n27418 = n27415 & ~n27416;
  assign n27419 = ~n27417 & ~n27418;
  assign n27420 = n27219 & n27419;
  assign n27421 = ~n27219 & ~n27419;
  assign po9  = ~n27420 & ~n27421;
  assign n27423 = ~n27414 & ~n27418;
  assign n27424 = n27272 & ~n27282;
  assign n27425 = ~n27285 & ~n27295;
  assign n27426 = ~n27424 & ~n27425;
  assign n27427 = n86 & n21033;
  assign n27428 = n4420 & n22674;
  assign n27429 = n4600 & n21030;
  assign n27430 = n4615 & n21027;
  assign n27431 = ~n27427 & ~n27429;
  assign n27432 = ~n27430 & n27431;
  assign n27433 = ~n27428 & n27432;
  assign n27434 = pi26  & n27433;
  assign n27435 = ~pi26  & ~n27433;
  assign n27436 = ~n27434 & ~n27435;
  assign n27437 = n27257 & ~n27264;
  assign n27438 = ~n27271 & ~n27437;
  assign n27439 = ~n27252 & ~n27255;
  assign n27440 = ~n184 & ~n367;
  assign n27441 = ~n792 & ~n937;
  assign n27442 = n27440 & n27441;
  assign n27443 = n755 & n1171;
  assign n27444 = n1948 & n2042;
  assign n27445 = n3205 & n4857;
  assign n27446 = n27444 & n27445;
  assign n27447 = n27442 & n27443;
  assign n27448 = n5475 & n27447;
  assign n27449 = n12979 & n27446;
  assign n27450 = n27448 & n27449;
  assign n27451 = n22104 & n27450;
  assign n27452 = n4183 & n27451;
  assign n27453 = n2650 & n27452;
  assign n27454 = n26846 & n27453;
  assign n27455 = ~n26846 & ~n27453;
  assign n27456 = ~n27454 & ~n27455;
  assign n27457 = ~n14144 & n26569;
  assign n27458 = ~pi5  & n27457;
  assign n27459 = pi5  & ~n27457;
  assign n27460 = ~n27458 & ~n27459;
  assign n27461 = ~n27456 & n27460;
  assign n27462 = n27456 & ~n27460;
  assign n27463 = ~n27461 & ~n27462;
  assign n27464 = ~n27439 & n27463;
  assign n27465 = n27439 & ~n27463;
  assign n27466 = ~n27464 & ~n27465;
  assign n27467 = n748 & n21051;
  assign n27468 = n880 & n21797;
  assign n27469 = n3692 & n21048;
  assign n27470 = n3694 & n21045;
  assign n27471 = ~n27467 & ~n27469;
  assign n27472 = ~n27470 & n27471;
  assign n27473 = ~n27468 & n27472;
  assign n27474 = n27466 & ~n27473;
  assign n27475 = ~n27466 & n27473;
  assign n27476 = ~n27474 & ~n27475;
  assign n27477 = n27438 & ~n27476;
  assign n27478 = ~n27438 & n27476;
  assign n27479 = ~n27477 & ~n27478;
  assign n27480 = n3810 & n21042;
  assign n27481 = n3886 & n22199;
  assign n27482 = n3884 & n21039;
  assign n27483 = n4380 & n21036;
  assign n27484 = ~n27480 & ~n27482;
  assign n27485 = ~n27483 & n27484;
  assign n27486 = ~n27481 & n27485;
  assign n27487 = pi29  & n27486;
  assign n27488 = ~pi29  & ~n27486;
  assign n27489 = ~n27487 & ~n27488;
  assign n27490 = n27479 & ~n27489;
  assign n27491 = ~n27479 & n27489;
  assign n27492 = ~n27490 & ~n27491;
  assign n27493 = ~n27436 & n27492;
  assign n27494 = n27436 & ~n27492;
  assign n27495 = ~n27493 & ~n27494;
  assign n27496 = n27426 & ~n27495;
  assign n27497 = ~n27426 & n27495;
  assign n27498 = ~n27496 & ~n27497;
  assign n27499 = n5044 & n21024;
  assign n27500 = n5045 & n23033;
  assign n27501 = n5109 & n21021;
  assign n27502 = n5130 & n21018;
  assign n27503 = ~n27499 & ~n27501;
  assign n27504 = ~n27502 & n27503;
  assign n27505 = ~n27500 & n27504;
  assign n27506 = pi23  & n27505;
  assign n27507 = ~pi23  & ~n27505;
  assign n27508 = ~n27506 & ~n27507;
  assign n27509 = n27498 & n27508;
  assign n27510 = ~n27498 & ~n27508;
  assign n27511 = ~n27509 & ~n27510;
  assign n27512 = ~n27303 & n27314;
  assign n27513 = ~n27302 & ~n27512;
  assign n27514 = n27511 & ~n27513;
  assign n27515 = ~n27511 & n27513;
  assign n27516 = ~n27514 & ~n27515;
  assign n27517 = n5240 & n21015;
  assign n27518 = n5241 & n23190;
  assign n27519 = n5853 & n21012;
  assign n27520 = n5866 & n21009;
  assign n27521 = ~n27517 & ~n27519;
  assign n27522 = ~n27520 & n27521;
  assign n27523 = ~n27518 & n27522;
  assign n27524 = pi20  & n27523;
  assign n27525 = ~pi20  & ~n27523;
  assign n27526 = ~n27524 & ~n27525;
  assign n27527 = n27516 & n27526;
  assign n27528 = ~n27516 & ~n27526;
  assign n27529 = ~n27527 & ~n27528;
  assign n27530 = ~n27321 & n27332;
  assign n27531 = ~n27320 & ~n27530;
  assign n27532 = n27529 & ~n27531;
  assign n27533 = ~n27529 & n27531;
  assign n27534 = ~n27532 & ~n27533;
  assign n27535 = n5982 & n21006;
  assign n27536 = n5983 & n23833;
  assign n27537 = n6323 & n20906;
  assign n27538 = n6336 & n21003;
  assign n27539 = ~n27535 & ~n27537;
  assign n27540 = ~n27538 & n27539;
  assign n27541 = ~n27536 & n27540;
  assign n27542 = pi17  & n27541;
  assign n27543 = ~pi17  & ~n27541;
  assign n27544 = ~n27542 & ~n27543;
  assign n27545 = n27534 & n27544;
  assign n27546 = ~n27534 & ~n27544;
  assign n27547 = ~n27545 & ~n27546;
  assign n27548 = ~n27339 & n27350;
  assign n27549 = ~n27338 & ~n27548;
  assign n27550 = n27547 & ~n27549;
  assign n27551 = ~n27547 & n27549;
  assign n27552 = ~n27550 & ~n27551;
  assign n27553 = n6630 & n21288;
  assign n27554 = n6631 & n24584;
  assign n27555 = n7238 & n24428;
  assign n27556 = n7262 & n24494;
  assign n27557 = ~n27553 & ~n27555;
  assign n27558 = ~n27556 & n27557;
  assign n27559 = ~n27554 & n27558;
  assign n27560 = pi14  & n27559;
  assign n27561 = ~pi14  & ~n27559;
  assign n27562 = ~n27560 & ~n27561;
  assign n27563 = ~n27357 & n27368;
  assign n27564 = ~n27356 & ~n27563;
  assign n27565 = n27562 & n27564;
  assign n27566 = ~n27562 & ~n27564;
  assign n27567 = ~n27565 & ~n27566;
  assign n27568 = ~n27552 & n27567;
  assign n27569 = n27552 & ~n27567;
  assign n27570 = ~n27568 & ~n27569;
  assign n27571 = n7430 & n24562;
  assign n27572 = n7431 & n25605;
  assign n27573 = n7869 & n25336;
  assign n27574 = n7895 & n25599;
  assign n27575 = ~n27571 & ~n27573;
  assign n27576 = ~n27574 & n27575;
  assign n27577 = ~n27572 & n27576;
  assign n27578 = pi11  & n27577;
  assign n27579 = ~pi11  & ~n27577;
  assign n27580 = ~n27578 & ~n27579;
  assign n27581 = n27570 & n27580;
  assign n27582 = ~n27570 & ~n27580;
  assign n27583 = ~n27581 & ~n27582;
  assign n27584 = ~n27375 & n27386;
  assign n27585 = ~n27374 & ~n27584;
  assign n27586 = n27583 & ~n27585;
  assign n27587 = ~n27583 & n27585;
  assign n27588 = ~n27586 & ~n27587;
  assign n27589 = n8250 & n25853;
  assign n27590 = n8251 & n26347;
  assign n27591 = n9016 & n26094;
  assign n27592 = n9040 & n26341;
  assign n27593 = ~n27589 & ~n27591;
  assign n27594 = ~n27592 & n27593;
  assign n27595 = ~n27590 & n27594;
  assign n27596 = pi8  & n27595;
  assign n27597 = ~pi8  & ~n27595;
  assign n27598 = ~n27596 & ~n27597;
  assign n27599 = ~n27393 & n27404;
  assign n27600 = ~n27392 & ~n27599;
  assign n27601 = n27598 & n27600;
  assign n27602 = ~n27598 & ~n27600;
  assign n27603 = ~n27601 & ~n27602;
  assign n27604 = ~n27588 & n27603;
  assign n27605 = n27588 & ~n27603;
  assign n27606 = ~n27604 & ~n27605;
  assign n27607 = ~n27232 & ~n27407;
  assign n27608 = ~n27233 & ~n27607;
  assign n27609 = n27606 & n27608;
  assign n27610 = ~n27606 & ~n27608;
  assign n27611 = ~n27609 & ~n27610;
  assign n27612 = ~n27423 & n27611;
  assign n27613 = n27423 & ~n27611;
  assign n27614 = ~n27612 & ~n27613;
  assign n27615 = ~n27420 & ~n27614;
  assign n27616 = n27420 & n27614;
  assign po10  = ~n27615 & ~n27616;
  assign n27618 = ~n27609 & ~n27612;
  assign n27619 = ~n27598 & n27600;
  assign n27620 = ~n27605 & ~n27619;
  assign n27621 = n27570 & ~n27580;
  assign n27622 = ~n27587 & ~n27621;
  assign n27623 = ~n27562 & n27564;
  assign n27624 = ~n27569 & ~n27623;
  assign n27625 = n27534 & ~n27544;
  assign n27626 = ~n27551 & ~n27625;
  assign n27627 = n27516 & ~n27526;
  assign n27628 = ~n27533 & ~n27627;
  assign n27629 = n27498 & ~n27508;
  assign n27630 = ~n27515 & ~n27629;
  assign n27631 = ~n27493 & ~n27497;
  assign n27632 = ~n27464 & ~n27474;
  assign n27633 = n26846 & ~n27453;
  assign n27634 = ~n27461 & ~n27633;
  assign n27635 = ~n435 & ~n989;
  assign n27636 = n784 & n27635;
  assign n27637 = n1010 & n1685;
  assign n27638 = n1858 & n2168;
  assign n27639 = n2192 & n27638;
  assign n27640 = n27636 & n27637;
  assign n27641 = n2128 & n27640;
  assign n27642 = n6432 & n27639;
  assign n27643 = n7057 & n27642;
  assign n27644 = n1236 & n27641;
  assign n27645 = n27643 & n27644;
  assign n27646 = ~n329 & ~n362;
  assign n27647 = ~n370 & ~n698;
  assign n27648 = ~n894 & n27647;
  assign n27649 = n142 & n27646;
  assign n27650 = n530 & n1359;
  assign n27651 = n1430 & n2503;
  assign n27652 = n4167 & n4269;
  assign n27653 = n27651 & n27652;
  assign n27654 = n27649 & n27650;
  assign n27655 = n3431 & n27648;
  assign n27656 = n27654 & n27655;
  assign n27657 = n1668 & n27653;
  assign n27658 = n7016 & n27657;
  assign n27659 = n2330 & n27656;
  assign n27660 = n27658 & n27659;
  assign n27661 = n27645 & n27660;
  assign n27662 = n1607 & n27661;
  assign n27663 = ~n27634 & n27662;
  assign n27664 = n27634 & ~n27662;
  assign n27665 = ~n27663 & ~n27664;
  assign n27666 = n748 & n21048;
  assign n27667 = n880 & n22049;
  assign n27668 = n3692 & n21045;
  assign n27669 = n3694 & n21042;
  assign n27670 = ~n27666 & ~n27668;
  assign n27671 = ~n27669 & n27670;
  assign n27672 = ~n27667 & n27671;
  assign n27673 = n27665 & ~n27672;
  assign n27674 = ~n27665 & n27672;
  assign n27675 = ~n27673 & ~n27674;
  assign n27676 = n27632 & ~n27675;
  assign n27677 = ~n27632 & n27675;
  assign n27678 = ~n27676 & ~n27677;
  assign n27679 = n3810 & n21039;
  assign n27680 = n3886 & n22186;
  assign n27681 = n3884 & n21036;
  assign n27682 = n4380 & n21033;
  assign n27683 = ~n27679 & ~n27681;
  assign n27684 = ~n27682 & n27683;
  assign n27685 = ~n27680 & n27684;
  assign n27686 = pi29  & n27685;
  assign n27687 = ~pi29  & ~n27685;
  assign n27688 = ~n27686 & ~n27687;
  assign n27689 = n27678 & ~n27688;
  assign n27690 = ~n27678 & n27688;
  assign n27691 = ~n27689 & ~n27690;
  assign n27692 = ~n27478 & n27489;
  assign n27693 = ~n27477 & ~n27692;
  assign n27694 = n27691 & n27693;
  assign n27695 = ~n27691 & ~n27693;
  assign n27696 = ~n27694 & ~n27695;
  assign n27697 = n86 & n21030;
  assign n27698 = n4420 & n22654;
  assign n27699 = n4600 & n21027;
  assign n27700 = n4615 & n21024;
  assign n27701 = ~n27697 & ~n27699;
  assign n27702 = ~n27700 & n27701;
  assign n27703 = ~n27698 & n27702;
  assign n27704 = pi26  & n27703;
  assign n27705 = ~pi26  & ~n27703;
  assign n27706 = ~n27704 & ~n27705;
  assign n27707 = n27696 & ~n27706;
  assign n27708 = ~n27696 & n27706;
  assign n27709 = ~n27707 & ~n27708;
  assign n27710 = n27631 & ~n27709;
  assign n27711 = ~n27631 & n27709;
  assign n27712 = ~n27710 & ~n27711;
  assign n27713 = n5044 & n21021;
  assign n27714 = n5045 & n23220;
  assign n27715 = n5109 & n21018;
  assign n27716 = n5130 & n21015;
  assign n27717 = ~n27713 & ~n27715;
  assign n27718 = ~n27716 & n27717;
  assign n27719 = ~n27714 & n27718;
  assign n27720 = pi23  & n27719;
  assign n27721 = ~pi23  & ~n27719;
  assign n27722 = ~n27720 & ~n27721;
  assign n27723 = n27712 & ~n27722;
  assign n27724 = ~n27712 & n27722;
  assign n27725 = ~n27723 & ~n27724;
  assign n27726 = n27630 & ~n27725;
  assign n27727 = ~n27630 & n27725;
  assign n27728 = ~n27726 & ~n27727;
  assign n27729 = n5240 & n21012;
  assign n27730 = n5241 & n23812;
  assign n27731 = n5853 & n21009;
  assign n27732 = n5866 & n21006;
  assign n27733 = ~n27729 & ~n27731;
  assign n27734 = ~n27732 & n27733;
  assign n27735 = ~n27730 & n27734;
  assign n27736 = pi20  & n27735;
  assign n27737 = ~pi20  & ~n27735;
  assign n27738 = ~n27736 & ~n27737;
  assign n27739 = n27728 & ~n27738;
  assign n27740 = ~n27728 & n27738;
  assign n27741 = ~n27739 & ~n27740;
  assign n27742 = n27628 & ~n27741;
  assign n27743 = ~n27628 & n27741;
  assign n27744 = ~n27742 & ~n27743;
  assign n27745 = n5982 & n20906;
  assign n27746 = n5983 & n21294;
  assign n27747 = n6323 & n21003;
  assign n27748 = n6336 & n21288;
  assign n27749 = ~n27745 & ~n27747;
  assign n27750 = ~n27748 & n27749;
  assign n27751 = ~n27746 & n27750;
  assign n27752 = pi17  & n27751;
  assign n27753 = ~pi17  & ~n27751;
  assign n27754 = ~n27752 & ~n27753;
  assign n27755 = n27744 & ~n27754;
  assign n27756 = ~n27744 & n27754;
  assign n27757 = ~n27755 & ~n27756;
  assign n27758 = n27626 & ~n27757;
  assign n27759 = ~n27626 & n27757;
  assign n27760 = ~n27758 & ~n27759;
  assign n27761 = n6630 & n24428;
  assign n27762 = n6631 & n24568;
  assign n27763 = n7238 & n24494;
  assign n27764 = n7262 & n24562;
  assign n27765 = ~n27761 & ~n27763;
  assign n27766 = ~n27764 & n27765;
  assign n27767 = ~n27762 & n27766;
  assign n27768 = pi14  & n27767;
  assign n27769 = ~pi14  & ~n27767;
  assign n27770 = ~n27768 & ~n27769;
  assign n27771 = n27760 & ~n27770;
  assign n27772 = ~n27760 & n27770;
  assign n27773 = ~n27771 & ~n27772;
  assign n27774 = n27624 & n27773;
  assign n27775 = ~n27624 & ~n27773;
  assign n27776 = ~n27774 & ~n27775;
  assign n27777 = n7430 & n25336;
  assign n27778 = n7431 & n25859;
  assign n27779 = n7869 & n25599;
  assign n27780 = n7895 & n25853;
  assign n27781 = ~n27777 & ~n27779;
  assign n27782 = ~n27780 & n27781;
  assign n27783 = ~n27778 & n27782;
  assign n27784 = pi11  & n27783;
  assign n27785 = ~pi11  & ~n27783;
  assign n27786 = ~n27784 & ~n27785;
  assign n27787 = ~n27776 & ~n27786;
  assign n27788 = n27776 & n27786;
  assign n27789 = ~n27787 & ~n27788;
  assign n27790 = n27622 & ~n27789;
  assign n27791 = ~n27622 & n27789;
  assign n27792 = ~n27790 & ~n27791;
  assign n27793 = n8250 & n26094;
  assign n27794 = n8251 & n26575;
  assign n27795 = n9016 & n26341;
  assign n27796 = n9040 & n26569;
  assign n27797 = ~n27793 & ~n27795;
  assign n27798 = ~n27796 & n27797;
  assign n27799 = ~n27794 & n27798;
  assign n27800 = pi8  & n27799;
  assign n27801 = ~pi8  & ~n27799;
  assign n27802 = ~n27800 & ~n27801;
  assign n27803 = n27792 & ~n27802;
  assign n27804 = ~n27792 & n27802;
  assign n27805 = ~n27803 & ~n27804;
  assign n27806 = ~n27620 & n27805;
  assign n27807 = n27620 & ~n27805;
  assign n27808 = ~n27806 & ~n27807;
  assign n27809 = n27618 & ~n27808;
  assign n27810 = ~n27618 & n27808;
  assign n27811 = ~n27809 & ~n27810;
  assign n27812 = n27616 & n27811;
  assign n27813 = ~n27616 & ~n27811;
  assign po11  = ~n27812 & ~n27813;
  assign n27815 = ~n27624 & n27773;
  assign n27816 = ~n27787 & ~n27815;
  assign n27817 = ~n16364 & n26569;
  assign n27818 = n8250 & n26341;
  assign n27819 = n8251 & ~n26793;
  assign n27820 = ~n27817 & ~n27818;
  assign n27821 = ~n27819 & n27820;
  assign n27822 = pi8  & n27821;
  assign n27823 = ~pi8  & ~n27821;
  assign n27824 = ~n27822 & ~n27823;
  assign n27825 = ~n27816 & ~n27824;
  assign n27826 = n27816 & n27824;
  assign n27827 = ~n27825 & ~n27826;
  assign n27828 = ~n200 & ~n499;
  assign n27829 = ~n639 & ~n715;
  assign n27830 = ~n1034 & n27829;
  assign n27831 = n417 & n27828;
  assign n27832 = n501 & n635;
  assign n27833 = n900 & n27832;
  assign n27834 = n27830 & n27831;
  assign n27835 = n241 & n4829;
  assign n27836 = n27834 & n27835;
  assign n27837 = n1893 & n27833;
  assign n27838 = n27836 & n27837;
  assign n27839 = n3135 & n27838;
  assign n27840 = ~n171 & ~n235;
  assign n27841 = ~n243 & ~n362;
  assign n27842 = ~n459 & ~n537;
  assign n27843 = ~n597 & ~n721;
  assign n27844 = ~n944 & n27843;
  assign n27845 = n27841 & n27842;
  assign n27846 = n27840 & n27845;
  assign n27847 = n27844 & n27846;
  assign n27848 = ~n271 & ~n383;
  assign n27849 = ~n458 & ~n603;
  assign n27850 = ~n751 & ~n846;
  assign n27851 = n27849 & n27850;
  assign n27852 = n3868 & n27848;
  assign n27853 = n27851 & n27852;
  assign n27854 = n6874 & n12691;
  assign n27855 = n27853 & n27854;
  assign n27856 = n4190 & n27855;
  assign n27857 = n27847 & n27856;
  assign n27858 = n4062 & n27857;
  assign n27859 = n27839 & n27858;
  assign n27860 = n12961 & n27859;
  assign n27861 = ~n27662 & n27860;
  assign n27862 = n27662 & ~n27860;
  assign n27863 = ~n27861 & ~n27862;
  assign n27864 = ~n27663 & n27672;
  assign n27865 = ~n27664 & ~n27864;
  assign n27866 = n27863 & n27865;
  assign n27867 = ~n27863 & ~n27865;
  assign n27868 = ~n27866 & ~n27867;
  assign n27869 = n748 & n21045;
  assign n27870 = n880 & n22217;
  assign n27871 = n3692 & n21042;
  assign n27872 = n3694 & n21039;
  assign n27873 = ~n27869 & ~n27871;
  assign n27874 = ~n27872 & n27873;
  assign n27875 = ~n27870 & n27874;
  assign n27876 = n27868 & n27875;
  assign n27877 = ~n27868 & ~n27875;
  assign n27878 = ~n27876 & ~n27877;
  assign n27879 = ~n27677 & ~n27689;
  assign n27880 = n27878 & n27879;
  assign n27881 = ~n27878 & ~n27879;
  assign n27882 = ~n27880 & ~n27881;
  assign n27883 = n3810 & n21036;
  assign n27884 = n3886 & n22632;
  assign n27885 = n3884 & n21033;
  assign n27886 = n4380 & n21030;
  assign n27887 = ~n27883 & ~n27885;
  assign n27888 = ~n27886 & n27887;
  assign n27889 = ~n27884 & n27888;
  assign n27890 = pi29  & n27889;
  assign n27891 = ~pi29  & ~n27889;
  assign n27892 = ~n27890 & ~n27891;
  assign n27893 = n27882 & n27892;
  assign n27894 = ~n27882 & ~n27892;
  assign n27895 = ~n27893 & ~n27894;
  assign n27896 = n86 & n21027;
  assign n27897 = n4420 & n21306;
  assign n27898 = n4600 & n21024;
  assign n27899 = n4615 & n21021;
  assign n27900 = ~n27896 & ~n27898;
  assign n27901 = ~n27899 & n27900;
  assign n27902 = ~n27897 & n27901;
  assign n27903 = pi26  & n27902;
  assign n27904 = ~pi26  & ~n27902;
  assign n27905 = ~n27903 & ~n27904;
  assign n27906 = ~n27895 & n27905;
  assign n27907 = n27895 & ~n27905;
  assign n27908 = ~n27906 & ~n27907;
  assign n27909 = ~n27694 & n27706;
  assign n27910 = ~n27695 & ~n27909;
  assign n27911 = n27908 & ~n27910;
  assign n27912 = ~n27908 & n27910;
  assign n27913 = ~n27911 & ~n27912;
  assign n27914 = n5044 & n21018;
  assign n27915 = n5045 & n23205;
  assign n27916 = n5109 & n21015;
  assign n27917 = n5130 & n21012;
  assign n27918 = ~n27914 & ~n27916;
  assign n27919 = ~n27917 & n27918;
  assign n27920 = ~n27915 & n27919;
  assign n27921 = pi23  & n27920;
  assign n27922 = ~pi23  & ~n27920;
  assign n27923 = ~n27921 & ~n27922;
  assign n27924 = n27913 & ~n27923;
  assign n27925 = ~n27913 & n27923;
  assign n27926 = ~n27924 & ~n27925;
  assign n27927 = ~n27711 & n27722;
  assign n27928 = ~n27710 & ~n27927;
  assign n27929 = ~n27926 & ~n27928;
  assign n27930 = n27926 & n27928;
  assign n27931 = ~n27929 & ~n27930;
  assign n27932 = n5240 & n21009;
  assign n27933 = n5241 & n23851;
  assign n27934 = n5853 & n21006;
  assign n27935 = n5866 & n20906;
  assign n27936 = ~n27932 & ~n27934;
  assign n27937 = ~n27935 & n27936;
  assign n27938 = ~n27933 & n27937;
  assign n27939 = pi20  & n27938;
  assign n27940 = ~pi20  & ~n27938;
  assign n27941 = ~n27939 & ~n27940;
  assign n27942 = n27931 & ~n27941;
  assign n27943 = ~n27931 & n27941;
  assign n27944 = ~n27942 & ~n27943;
  assign n27945 = ~n27727 & n27738;
  assign n27946 = ~n27726 & ~n27945;
  assign n27947 = ~n27944 & ~n27946;
  assign n27948 = n27944 & n27946;
  assign n27949 = ~n27947 & ~n27948;
  assign n27950 = n5982 & n21003;
  assign n27951 = n5983 & n24596;
  assign n27952 = n6323 & n21288;
  assign n27953 = n6336 & n24428;
  assign n27954 = ~n27950 & ~n27952;
  assign n27955 = ~n27953 & n27954;
  assign n27956 = ~n27951 & n27955;
  assign n27957 = pi17  & n27956;
  assign n27958 = ~pi17  & ~n27956;
  assign n27959 = ~n27957 & ~n27958;
  assign n27960 = n27949 & ~n27959;
  assign n27961 = ~n27949 & n27959;
  assign n27962 = ~n27960 & ~n27961;
  assign n27963 = ~n27743 & n27754;
  assign n27964 = ~n27742 & ~n27963;
  assign n27965 = ~n27962 & ~n27964;
  assign n27966 = n27962 & n27964;
  assign n27967 = ~n27965 & ~n27966;
  assign n27968 = n6630 & n24494;
  assign n27969 = n6631 & n25342;
  assign n27970 = n7238 & n24562;
  assign n27971 = n7262 & n25336;
  assign n27972 = ~n27968 & ~n27970;
  assign n27973 = ~n27971 & n27972;
  assign n27974 = ~n27969 & n27973;
  assign n27975 = pi14  & n27974;
  assign n27976 = ~pi14  & ~n27974;
  assign n27977 = ~n27975 & ~n27976;
  assign n27978 = n27967 & ~n27977;
  assign n27979 = ~n27967 & n27977;
  assign n27980 = ~n27978 & ~n27979;
  assign n27981 = ~n27759 & n27770;
  assign n27982 = ~n27758 & ~n27981;
  assign n27983 = ~n27980 & ~n27982;
  assign n27984 = n27980 & n27982;
  assign n27985 = ~n27983 & ~n27984;
  assign n27986 = n7430 & n25599;
  assign n27987 = n7431 & n26100;
  assign n27988 = n7869 & n25853;
  assign n27989 = n7895 & n26094;
  assign n27990 = ~n27986 & ~n27988;
  assign n27991 = ~n27989 & n27990;
  assign n27992 = ~n27987 & n27991;
  assign n27993 = pi11  & n27992;
  assign n27994 = ~pi11  & ~n27992;
  assign n27995 = ~n27993 & ~n27994;
  assign n27996 = n27985 & ~n27995;
  assign n27997 = ~n27985 & n27995;
  assign n27998 = ~n27996 & ~n27997;
  assign n27999 = n27827 & n27998;
  assign n28000 = ~n27827 & ~n27998;
  assign n28001 = ~n27999 & ~n28000;
  assign n28002 = ~n27791 & n27802;
  assign n28003 = ~n27790 & ~n28002;
  assign n28004 = ~n28001 & ~n28003;
  assign n28005 = n28001 & n28003;
  assign n28006 = ~n28004 & ~n28005;
  assign n28007 = ~n27806 & ~n27810;
  assign n28008 = ~n28006 & n28007;
  assign n28009 = n28006 & ~n28007;
  assign n28010 = ~n28008 & ~n28009;
  assign n28011 = n27812 & n28010;
  assign n28012 = ~n27812 & ~n28010;
  assign po12  = ~n28011 & ~n28012;
  assign n28014 = ~n28005 & ~n28009;
  assign n28015 = n27868 & ~n27875;
  assign n28016 = ~n27881 & ~n28015;
  assign n28017 = n3810 & n21033;
  assign n28018 = n3886 & n22674;
  assign n28019 = n3884 & n21030;
  assign n28020 = n4380 & n21027;
  assign n28021 = ~n28017 & ~n28019;
  assign n28022 = ~n28020 & n28021;
  assign n28023 = ~n28018 & n28022;
  assign n28024 = pi29  & n28023;
  assign n28025 = ~pi29  & ~n28023;
  assign n28026 = ~n28024 & ~n28025;
  assign n28027 = ~n27862 & ~n27866;
  assign n28028 = ~n13688 & n26569;
  assign n28029 = pi8  & ~n28028;
  assign n28030 = ~pi8  & n28028;
  assign n28031 = ~n28029 & ~n28030;
  assign n28032 = ~n412 & ~n515;
  assign n28033 = n500 & n28032;
  assign n28034 = n1052 & n1948;
  assign n28035 = n2934 & n28034;
  assign n28036 = n1228 & n28033;
  assign n28037 = n1455 & n2333;
  assign n28038 = n12944 & n28037;
  assign n28039 = n28035 & n28036;
  assign n28040 = n12929 & n28039;
  assign n28041 = n28038 & n28040;
  assign n28042 = n2791 & n28041;
  assign n28043 = n1419 & n3457;
  assign n28044 = n28042 & n28043;
  assign n28045 = n27662 & n28044;
  assign n28046 = ~n27662 & ~n28044;
  assign n28047 = ~n28045 & ~n28046;
  assign n28048 = n28031 & n28047;
  assign n28049 = ~n28031 & ~n28047;
  assign n28050 = ~n28048 & ~n28049;
  assign n28051 = ~n28027 & n28050;
  assign n28052 = n28027 & ~n28050;
  assign n28053 = ~n28051 & ~n28052;
  assign n28054 = n748 & n21042;
  assign n28055 = n880 & n22199;
  assign n28056 = n3692 & n21039;
  assign n28057 = n3694 & n21036;
  assign n28058 = ~n28054 & ~n28056;
  assign n28059 = ~n28057 & n28058;
  assign n28060 = ~n28055 & n28059;
  assign n28061 = n28053 & ~n28060;
  assign n28062 = ~n28053 & n28060;
  assign n28063 = ~n28061 & ~n28062;
  assign n28064 = ~n28026 & n28063;
  assign n28065 = n28026 & ~n28063;
  assign n28066 = ~n28064 & ~n28065;
  assign n28067 = n28016 & ~n28066;
  assign n28068 = ~n28016 & n28066;
  assign n28069 = ~n28067 & ~n28068;
  assign n28070 = n86 & n21024;
  assign n28071 = n4420 & n23033;
  assign n28072 = n4600 & n21021;
  assign n28073 = n4615 & n21018;
  assign n28074 = ~n28070 & ~n28072;
  assign n28075 = ~n28073 & n28074;
  assign n28076 = ~n28071 & n28075;
  assign n28077 = pi26  & n28076;
  assign n28078 = ~pi26  & ~n28076;
  assign n28079 = ~n28077 & ~n28078;
  assign n28080 = n28069 & n28079;
  assign n28081 = ~n28069 & ~n28079;
  assign n28082 = ~n28080 & ~n28081;
  assign n28083 = n27882 & ~n27892;
  assign n28084 = ~n27895 & ~n27905;
  assign n28085 = ~n28083 & ~n28084;
  assign n28086 = n28082 & n28085;
  assign n28087 = ~n28082 & ~n28085;
  assign n28088 = ~n28086 & ~n28087;
  assign n28089 = n5044 & n21015;
  assign n28090 = n5045 & n23190;
  assign n28091 = n5109 & n21012;
  assign n28092 = n5130 & n21009;
  assign n28093 = ~n28089 & ~n28091;
  assign n28094 = ~n28092 & n28093;
  assign n28095 = ~n28090 & n28094;
  assign n28096 = pi23  & n28095;
  assign n28097 = ~pi23  & ~n28095;
  assign n28098 = ~n28096 & ~n28097;
  assign n28099 = n28088 & n28098;
  assign n28100 = ~n28088 & ~n28098;
  assign n28101 = ~n28099 & ~n28100;
  assign n28102 = ~n27912 & n27923;
  assign n28103 = ~n27911 & ~n28102;
  assign n28104 = n28101 & ~n28103;
  assign n28105 = ~n28101 & n28103;
  assign n28106 = ~n28104 & ~n28105;
  assign n28107 = n5240 & n21006;
  assign n28108 = n5241 & n23833;
  assign n28109 = n5853 & n20906;
  assign n28110 = n5866 & n21003;
  assign n28111 = ~n28107 & ~n28109;
  assign n28112 = ~n28110 & n28111;
  assign n28113 = ~n28108 & n28112;
  assign n28114 = pi20  & n28113;
  assign n28115 = ~pi20  & ~n28113;
  assign n28116 = ~n28114 & ~n28115;
  assign n28117 = n28106 & n28116;
  assign n28118 = ~n28106 & ~n28116;
  assign n28119 = ~n28117 & ~n28118;
  assign n28120 = ~n27930 & n27941;
  assign n28121 = ~n27929 & ~n28120;
  assign n28122 = n28119 & ~n28121;
  assign n28123 = ~n28119 & n28121;
  assign n28124 = ~n28122 & ~n28123;
  assign n28125 = n5982 & n21288;
  assign n28126 = n5983 & n24584;
  assign n28127 = n6323 & n24428;
  assign n28128 = n6336 & n24494;
  assign n28129 = ~n28125 & ~n28127;
  assign n28130 = ~n28128 & n28129;
  assign n28131 = ~n28126 & n28130;
  assign n28132 = pi17  & n28131;
  assign n28133 = ~pi17  & ~n28131;
  assign n28134 = ~n28132 & ~n28133;
  assign n28135 = ~n27948 & n27959;
  assign n28136 = ~n27947 & ~n28135;
  assign n28137 = n28134 & n28136;
  assign n28138 = ~n28134 & ~n28136;
  assign n28139 = ~n28137 & ~n28138;
  assign n28140 = ~n28124 & n28139;
  assign n28141 = n28124 & ~n28139;
  assign n28142 = ~n28140 & ~n28141;
  assign n28143 = n6630 & n24562;
  assign n28144 = n6631 & n25605;
  assign n28145 = n7238 & n25336;
  assign n28146 = n7262 & n25599;
  assign n28147 = ~n28143 & ~n28145;
  assign n28148 = ~n28146 & n28147;
  assign n28149 = ~n28144 & n28148;
  assign n28150 = pi14  & n28149;
  assign n28151 = ~pi14  & ~n28149;
  assign n28152 = ~n28150 & ~n28151;
  assign n28153 = n28142 & n28152;
  assign n28154 = ~n28142 & ~n28152;
  assign n28155 = ~n28153 & ~n28154;
  assign n28156 = ~n27966 & n27977;
  assign n28157 = ~n27965 & ~n28156;
  assign n28158 = n28155 & ~n28157;
  assign n28159 = ~n28155 & n28157;
  assign n28160 = ~n28158 & ~n28159;
  assign n28161 = n7430 & n25853;
  assign n28162 = n7431 & n26347;
  assign n28163 = n7869 & n26094;
  assign n28164 = n7895 & n26341;
  assign n28165 = ~n28161 & ~n28163;
  assign n28166 = ~n28164 & n28165;
  assign n28167 = ~n28162 & n28166;
  assign n28168 = pi11  & n28167;
  assign n28169 = ~pi11  & ~n28167;
  assign n28170 = ~n28168 & ~n28169;
  assign n28171 = ~n27984 & n27995;
  assign n28172 = ~n27983 & ~n28171;
  assign n28173 = n28170 & n28172;
  assign n28174 = ~n28170 & ~n28172;
  assign n28175 = ~n28173 & ~n28174;
  assign n28176 = ~n28160 & n28175;
  assign n28177 = n28160 & ~n28175;
  assign n28178 = ~n28176 & ~n28177;
  assign n28179 = ~n27825 & ~n27998;
  assign n28180 = ~n27826 & ~n28179;
  assign n28181 = n28178 & n28180;
  assign n28182 = ~n28178 & ~n28180;
  assign n28183 = ~n28181 & ~n28182;
  assign n28184 = ~n28014 & n28183;
  assign n28185 = n28014 & ~n28183;
  assign n28186 = ~n28184 & ~n28185;
  assign n28187 = ~n28011 & ~n28186;
  assign n28188 = n28011 & n28186;
  assign po13  = ~n28187 & ~n28188;
  assign n28190 = ~n28181 & ~n28184;
  assign n28191 = ~n28170 & n28172;
  assign n28192 = ~n28177 & ~n28191;
  assign n28193 = n28142 & ~n28152;
  assign n28194 = ~n28159 & ~n28193;
  assign n28195 = ~n28134 & n28136;
  assign n28196 = ~n28141 & ~n28195;
  assign n28197 = n28106 & ~n28116;
  assign n28198 = ~n28123 & ~n28197;
  assign n28199 = n28088 & ~n28098;
  assign n28200 = ~n28105 & ~n28199;
  assign n28201 = n28069 & ~n28079;
  assign n28202 = ~n28087 & ~n28201;
  assign n28203 = ~n28064 & ~n28068;
  assign n28204 = ~n28046 & ~n28048;
  assign n28205 = ~n235 & ~n242;
  assign n28206 = ~n893 & n28205;
  assign n28207 = n360 & n1053;
  assign n28208 = n2349 & n3344;
  assign n28209 = n28207 & n28208;
  assign n28210 = n3279 & n28206;
  assign n28211 = n14380 & n14877;
  assign n28212 = n28210 & n28211;
  assign n28213 = n5305 & n28209;
  assign n28214 = n28212 & n28213;
  assign n28215 = n13516 & n28214;
  assign n28216 = n1208 & n28215;
  assign n28217 = n2570 & n28216;
  assign n28218 = ~n28204 & n28217;
  assign n28219 = n28204 & ~n28217;
  assign n28220 = ~n28218 & ~n28219;
  assign n28221 = n748 & n21039;
  assign n28222 = n880 & n22186;
  assign n28223 = n3692 & n21036;
  assign n28224 = n3694 & n21033;
  assign n28225 = ~n28221 & ~n28223;
  assign n28226 = ~n28224 & n28225;
  assign n28227 = ~n28222 & n28226;
  assign n28228 = n28220 & ~n28227;
  assign n28229 = ~n28220 & n28227;
  assign n28230 = ~n28228 & ~n28229;
  assign n28231 = ~n28051 & n28060;
  assign n28232 = ~n28052 & ~n28231;
  assign n28233 = ~n28230 & ~n28232;
  assign n28234 = n28230 & n28232;
  assign n28235 = ~n28233 & ~n28234;
  assign n28236 = n3810 & n21030;
  assign n28237 = n3886 & n22654;
  assign n28238 = n3884 & n21027;
  assign n28239 = n4380 & n21024;
  assign n28240 = ~n28236 & ~n28238;
  assign n28241 = ~n28239 & n28240;
  assign n28242 = ~n28237 & n28241;
  assign n28243 = pi29  & n28242;
  assign n28244 = ~pi29  & ~n28242;
  assign n28245 = ~n28243 & ~n28244;
  assign n28246 = n28235 & ~n28245;
  assign n28247 = ~n28235 & n28245;
  assign n28248 = ~n28246 & ~n28247;
  assign n28249 = ~n28203 & n28248;
  assign n28250 = n28203 & ~n28248;
  assign n28251 = ~n28249 & ~n28250;
  assign n28252 = n86 & n21021;
  assign n28253 = n4420 & n23220;
  assign n28254 = n4600 & n21018;
  assign n28255 = n4615 & n21015;
  assign n28256 = ~n28252 & ~n28254;
  assign n28257 = ~n28255 & n28256;
  assign n28258 = ~n28253 & n28257;
  assign n28259 = pi26  & n28258;
  assign n28260 = ~pi26  & ~n28258;
  assign n28261 = ~n28259 & ~n28260;
  assign n28262 = n28251 & ~n28261;
  assign n28263 = ~n28251 & n28261;
  assign n28264 = ~n28262 & ~n28263;
  assign n28265 = n28202 & ~n28264;
  assign n28266 = ~n28202 & n28264;
  assign n28267 = ~n28265 & ~n28266;
  assign n28268 = n5044 & n21012;
  assign n28269 = n5045 & n23812;
  assign n28270 = n5109 & n21009;
  assign n28271 = n5130 & n21006;
  assign n28272 = ~n28268 & ~n28270;
  assign n28273 = ~n28271 & n28272;
  assign n28274 = ~n28269 & n28273;
  assign n28275 = pi23  & n28274;
  assign n28276 = ~pi23  & ~n28274;
  assign n28277 = ~n28275 & ~n28276;
  assign n28278 = n28267 & ~n28277;
  assign n28279 = ~n28267 & n28277;
  assign n28280 = ~n28278 & ~n28279;
  assign n28281 = n28200 & ~n28280;
  assign n28282 = ~n28200 & n28280;
  assign n28283 = ~n28281 & ~n28282;
  assign n28284 = n5240 & n20906;
  assign n28285 = n5241 & n21294;
  assign n28286 = n5853 & n21003;
  assign n28287 = n5866 & n21288;
  assign n28288 = ~n28284 & ~n28286;
  assign n28289 = ~n28287 & n28288;
  assign n28290 = ~n28285 & n28289;
  assign n28291 = pi20  & n28290;
  assign n28292 = ~pi20  & ~n28290;
  assign n28293 = ~n28291 & ~n28292;
  assign n28294 = n28283 & ~n28293;
  assign n28295 = ~n28283 & n28293;
  assign n28296 = ~n28294 & ~n28295;
  assign n28297 = n28198 & ~n28296;
  assign n28298 = ~n28198 & n28296;
  assign n28299 = ~n28297 & ~n28298;
  assign n28300 = n5982 & n24428;
  assign n28301 = n5983 & n24568;
  assign n28302 = n6323 & n24494;
  assign n28303 = n6336 & n24562;
  assign n28304 = ~n28300 & ~n28302;
  assign n28305 = ~n28303 & n28304;
  assign n28306 = ~n28301 & n28305;
  assign n28307 = pi17  & n28306;
  assign n28308 = ~pi17  & ~n28306;
  assign n28309 = ~n28307 & ~n28308;
  assign n28310 = n28299 & ~n28309;
  assign n28311 = ~n28299 & n28309;
  assign n28312 = ~n28310 & ~n28311;
  assign n28313 = n28196 & n28312;
  assign n28314 = ~n28196 & ~n28312;
  assign n28315 = ~n28313 & ~n28314;
  assign n28316 = n6630 & n25336;
  assign n28317 = n6631 & n25859;
  assign n28318 = n7238 & n25599;
  assign n28319 = n7262 & n25853;
  assign n28320 = ~n28316 & ~n28318;
  assign n28321 = ~n28319 & n28320;
  assign n28322 = ~n28317 & n28321;
  assign n28323 = pi14  & n28322;
  assign n28324 = ~pi14  & ~n28322;
  assign n28325 = ~n28323 & ~n28324;
  assign n28326 = ~n28315 & ~n28325;
  assign n28327 = n28315 & n28325;
  assign n28328 = ~n28326 & ~n28327;
  assign n28329 = n28194 & ~n28328;
  assign n28330 = ~n28194 & n28328;
  assign n28331 = ~n28329 & ~n28330;
  assign n28332 = n7430 & n26094;
  assign n28333 = n7431 & n26575;
  assign n28334 = n7869 & n26341;
  assign n28335 = n7895 & n26569;
  assign n28336 = ~n28332 & ~n28334;
  assign n28337 = ~n28335 & n28336;
  assign n28338 = ~n28333 & n28337;
  assign n28339 = pi11  & n28338;
  assign n28340 = ~pi11  & ~n28338;
  assign n28341 = ~n28339 & ~n28340;
  assign n28342 = n28331 & ~n28341;
  assign n28343 = ~n28331 & n28341;
  assign n28344 = ~n28342 & ~n28343;
  assign n28345 = ~n28192 & n28344;
  assign n28346 = n28192 & ~n28344;
  assign n28347 = ~n28345 & ~n28346;
  assign n28348 = n28190 & ~n28347;
  assign n28349 = ~n28190 & n28347;
  assign n28350 = ~n28348 & ~n28349;
  assign n28351 = n28188 & n28350;
  assign n28352 = ~n28188 & ~n28350;
  assign po14  = ~n28351 & ~n28352;
  assign n28354 = ~n28196 & n28312;
  assign n28355 = ~n28326 & ~n28354;
  assign n28356 = ~n15450 & n26569;
  assign n28357 = n7430 & n26341;
  assign n28358 = n7431 & ~n26793;
  assign n28359 = ~n28356 & ~n28357;
  assign n28360 = ~n28358 & n28359;
  assign n28361 = pi11  & n28360;
  assign n28362 = ~pi11  & ~n28360;
  assign n28363 = ~n28361 & ~n28362;
  assign n28364 = ~n28355 & ~n28363;
  assign n28365 = n28355 & n28363;
  assign n28366 = ~n28364 & ~n28365;
  assign n28367 = ~n28234 & ~n28246;
  assign n28368 = ~n274 & ~n422;
  assign n28369 = ~n838 & n28368;
  assign n28370 = n117 & n431;
  assign n28371 = n1035 & n1188;
  assign n28372 = n1674 & n1962;
  assign n28373 = n2207 & n3460;
  assign n28374 = n28372 & n28373;
  assign n28375 = n28370 & n28371;
  assign n28376 = n3398 & n28369;
  assign n28377 = n15077 & n28376;
  assign n28378 = n28374 & n28375;
  assign n28379 = n28377 & n28378;
  assign n28380 = n12924 & n14385;
  assign n28381 = n28379 & n28380;
  assign n28382 = n5744 & n28381;
  assign n28383 = n27645 & n28382;
  assign n28384 = ~n28217 & n28383;
  assign n28385 = n28217 & ~n28383;
  assign n28386 = ~n28384 & ~n28385;
  assign n28387 = ~n28218 & n28227;
  assign n28388 = ~n28219 & ~n28387;
  assign n28389 = n28386 & n28388;
  assign n28390 = ~n28386 & ~n28388;
  assign n28391 = ~n28389 & ~n28390;
  assign n28392 = n748 & n21036;
  assign n28393 = n880 & n22632;
  assign n28394 = n3692 & n21033;
  assign n28395 = n3694 & n21030;
  assign n28396 = ~n28392 & ~n28394;
  assign n28397 = ~n28395 & n28396;
  assign n28398 = ~n28393 & n28397;
  assign n28399 = n28391 & n28398;
  assign n28400 = ~n28391 & ~n28398;
  assign n28401 = ~n28399 & ~n28400;
  assign n28402 = n3810 & n21027;
  assign n28403 = n3886 & n21306;
  assign n28404 = n3884 & n21024;
  assign n28405 = n4380 & n21021;
  assign n28406 = ~n28402 & ~n28404;
  assign n28407 = ~n28405 & n28406;
  assign n28408 = ~n28403 & n28407;
  assign n28409 = pi29  & n28408;
  assign n28410 = ~pi29  & ~n28408;
  assign n28411 = ~n28409 & ~n28410;
  assign n28412 = ~n28401 & ~n28411;
  assign n28413 = n28401 & n28411;
  assign n28414 = ~n28412 & ~n28413;
  assign n28415 = ~n28367 & n28414;
  assign n28416 = n28367 & ~n28414;
  assign n28417 = ~n28415 & ~n28416;
  assign n28418 = n86 & n21018;
  assign n28419 = n4420 & n23205;
  assign n28420 = n4600 & n21015;
  assign n28421 = n4615 & n21012;
  assign n28422 = ~n28418 & ~n28420;
  assign n28423 = ~n28421 & n28422;
  assign n28424 = ~n28419 & n28423;
  assign n28425 = pi26  & n28424;
  assign n28426 = ~pi26  & ~n28424;
  assign n28427 = ~n28425 & ~n28426;
  assign n28428 = n28417 & ~n28427;
  assign n28429 = ~n28417 & n28427;
  assign n28430 = ~n28428 & ~n28429;
  assign n28431 = ~n28249 & n28261;
  assign n28432 = ~n28250 & ~n28431;
  assign n28433 = ~n28430 & ~n28432;
  assign n28434 = n28430 & n28432;
  assign n28435 = ~n28433 & ~n28434;
  assign n28436 = n5044 & n21009;
  assign n28437 = n5045 & n23851;
  assign n28438 = n5109 & n21006;
  assign n28439 = n5130 & n20906;
  assign n28440 = ~n28436 & ~n28438;
  assign n28441 = ~n28439 & n28440;
  assign n28442 = ~n28437 & n28441;
  assign n28443 = pi23  & n28442;
  assign n28444 = ~pi23  & ~n28442;
  assign n28445 = ~n28443 & ~n28444;
  assign n28446 = n28435 & ~n28445;
  assign n28447 = ~n28435 & n28445;
  assign n28448 = ~n28446 & ~n28447;
  assign n28449 = ~n28266 & n28277;
  assign n28450 = ~n28265 & ~n28449;
  assign n28451 = ~n28448 & ~n28450;
  assign n28452 = n28448 & n28450;
  assign n28453 = ~n28451 & ~n28452;
  assign n28454 = n5240 & n21003;
  assign n28455 = n5241 & n24596;
  assign n28456 = n5853 & n21288;
  assign n28457 = n5866 & n24428;
  assign n28458 = ~n28454 & ~n28456;
  assign n28459 = ~n28457 & n28458;
  assign n28460 = ~n28455 & n28459;
  assign n28461 = pi20  & n28460;
  assign n28462 = ~pi20  & ~n28460;
  assign n28463 = ~n28461 & ~n28462;
  assign n28464 = n28453 & ~n28463;
  assign n28465 = ~n28453 & n28463;
  assign n28466 = ~n28464 & ~n28465;
  assign n28467 = ~n28282 & n28293;
  assign n28468 = ~n28281 & ~n28467;
  assign n28469 = ~n28466 & ~n28468;
  assign n28470 = n28466 & n28468;
  assign n28471 = ~n28469 & ~n28470;
  assign n28472 = n5982 & n24494;
  assign n28473 = n5983 & n25342;
  assign n28474 = n6323 & n24562;
  assign n28475 = n6336 & n25336;
  assign n28476 = ~n28472 & ~n28474;
  assign n28477 = ~n28475 & n28476;
  assign n28478 = ~n28473 & n28477;
  assign n28479 = pi17  & n28478;
  assign n28480 = ~pi17  & ~n28478;
  assign n28481 = ~n28479 & ~n28480;
  assign n28482 = n28471 & ~n28481;
  assign n28483 = ~n28471 & n28481;
  assign n28484 = ~n28482 & ~n28483;
  assign n28485 = ~n28298 & n28309;
  assign n28486 = ~n28297 & ~n28485;
  assign n28487 = ~n28484 & ~n28486;
  assign n28488 = n28484 & n28486;
  assign n28489 = ~n28487 & ~n28488;
  assign n28490 = n6630 & n25599;
  assign n28491 = n6631 & n26100;
  assign n28492 = n7238 & n25853;
  assign n28493 = n7262 & n26094;
  assign n28494 = ~n28490 & ~n28492;
  assign n28495 = ~n28493 & n28494;
  assign n28496 = ~n28491 & n28495;
  assign n28497 = pi14  & n28496;
  assign n28498 = ~pi14  & ~n28496;
  assign n28499 = ~n28497 & ~n28498;
  assign n28500 = n28489 & ~n28499;
  assign n28501 = ~n28489 & n28499;
  assign n28502 = ~n28500 & ~n28501;
  assign n28503 = n28366 & n28502;
  assign n28504 = ~n28366 & ~n28502;
  assign n28505 = ~n28503 & ~n28504;
  assign n28506 = ~n28330 & n28341;
  assign n28507 = ~n28329 & ~n28506;
  assign n28508 = ~n28505 & ~n28507;
  assign n28509 = n28505 & n28507;
  assign n28510 = ~n28508 & ~n28509;
  assign n28511 = ~n28345 & ~n28349;
  assign n28512 = ~n28510 & n28511;
  assign n28513 = n28510 & ~n28511;
  assign n28514 = ~n28512 & ~n28513;
  assign n28515 = n28351 & n28514;
  assign n28516 = ~n28351 & ~n28514;
  assign po15  = ~n28515 & ~n28516;
  assign n28518 = ~n28509 & ~n28513;
  assign n28519 = n86 & n21015;
  assign n28520 = n4420 & n23190;
  assign n28521 = n4600 & n21012;
  assign n28522 = n4615 & n21009;
  assign n28523 = ~n28519 & ~n28521;
  assign n28524 = ~n28522 & n28523;
  assign n28525 = ~n28520 & n28524;
  assign n28526 = pi26  & n28525;
  assign n28527 = ~pi26  & ~n28525;
  assign n28528 = ~n28526 & ~n28527;
  assign n28529 = n3810 & n21024;
  assign n28530 = n3886 & n23033;
  assign n28531 = n3884 & n21021;
  assign n28532 = n4380 & n21018;
  assign n28533 = ~n28529 & ~n28531;
  assign n28534 = ~n28532 & n28533;
  assign n28535 = ~n28530 & n28534;
  assign n28536 = pi29  & n28535;
  assign n28537 = ~pi29  & ~n28535;
  assign n28538 = ~n28536 & ~n28537;
  assign n28539 = n28391 & ~n28398;
  assign n28540 = ~n28412 & ~n28539;
  assign n28541 = ~n13532 & n26569;
  assign n28542 = pi11  & ~n28541;
  assign n28543 = ~pi11  & n28541;
  assign n28544 = ~n28542 & ~n28543;
  assign n28545 = ~n283 & ~n307;
  assign n28546 = ~n364 & ~n846;
  assign n28547 = n28545 & n28546;
  assign n28548 = n137 & n942;
  assign n28549 = n1244 & n1672;
  assign n28550 = n3408 & n28549;
  assign n28551 = n28547 & n28548;
  assign n28552 = n5509 & n13055;
  assign n28553 = n28551 & n28552;
  assign n28554 = n2938 & n28550;
  assign n28555 = n5494 & n28554;
  assign n28556 = n28553 & n28555;
  assign n28557 = n2291 & n28556;
  assign n28558 = n1320 & n2276;
  assign n28559 = n28557 & n28558;
  assign n28560 = n28217 & n28559;
  assign n28561 = ~n28217 & ~n28559;
  assign n28562 = ~n28560 & ~n28561;
  assign n28563 = n28544 & n28562;
  assign n28564 = ~n28544 & ~n28562;
  assign n28565 = ~n28563 & ~n28564;
  assign n28566 = n748 & n21033;
  assign n28567 = n880 & n22674;
  assign n28568 = n3692 & n21030;
  assign n28569 = n3694 & n21027;
  assign n28570 = ~n28566 & ~n28568;
  assign n28571 = ~n28569 & n28570;
  assign n28572 = ~n28567 & n28571;
  assign n28573 = n28565 & n28572;
  assign n28574 = ~n28565 & ~n28572;
  assign n28575 = ~n28573 & ~n28574;
  assign n28576 = ~n28385 & ~n28389;
  assign n28577 = ~n28575 & n28576;
  assign n28578 = n28575 & ~n28576;
  assign n28579 = ~n28577 & ~n28578;
  assign n28580 = ~n28540 & ~n28579;
  assign n28581 = n28540 & n28579;
  assign n28582 = ~n28580 & ~n28581;
  assign n28583 = n28538 & ~n28582;
  assign n28584 = ~n28538 & n28582;
  assign n28585 = ~n28583 & ~n28584;
  assign n28586 = n28528 & n28585;
  assign n28587 = ~n28528 & ~n28585;
  assign n28588 = ~n28586 & ~n28587;
  assign n28589 = ~n28415 & n28427;
  assign n28590 = ~n28416 & ~n28589;
  assign n28591 = n28588 & ~n28590;
  assign n28592 = ~n28588 & n28590;
  assign n28593 = ~n28591 & ~n28592;
  assign n28594 = n5044 & n21006;
  assign n28595 = n5045 & n23833;
  assign n28596 = n5109 & n20906;
  assign n28597 = n5130 & n21003;
  assign n28598 = ~n28594 & ~n28596;
  assign n28599 = ~n28597 & n28598;
  assign n28600 = ~n28595 & n28599;
  assign n28601 = pi23  & n28600;
  assign n28602 = ~pi23  & ~n28600;
  assign n28603 = ~n28601 & ~n28602;
  assign n28604 = n28593 & n28603;
  assign n28605 = ~n28593 & ~n28603;
  assign n28606 = ~n28604 & ~n28605;
  assign n28607 = ~n28434 & n28445;
  assign n28608 = ~n28433 & ~n28607;
  assign n28609 = n28606 & ~n28608;
  assign n28610 = ~n28606 & n28608;
  assign n28611 = ~n28609 & ~n28610;
  assign n28612 = n5240 & n21288;
  assign n28613 = n5241 & n24584;
  assign n28614 = n5853 & n24428;
  assign n28615 = n5866 & n24494;
  assign n28616 = ~n28612 & ~n28614;
  assign n28617 = ~n28615 & n28616;
  assign n28618 = ~n28613 & n28617;
  assign n28619 = pi20  & n28618;
  assign n28620 = ~pi20  & ~n28618;
  assign n28621 = ~n28619 & ~n28620;
  assign n28622 = ~n28452 & n28463;
  assign n28623 = ~n28451 & ~n28622;
  assign n28624 = n28621 & n28623;
  assign n28625 = ~n28621 & ~n28623;
  assign n28626 = ~n28624 & ~n28625;
  assign n28627 = ~n28611 & n28626;
  assign n28628 = n28611 & ~n28626;
  assign n28629 = ~n28627 & ~n28628;
  assign n28630 = n5982 & n24562;
  assign n28631 = n5983 & n25605;
  assign n28632 = n6323 & n25336;
  assign n28633 = n6336 & n25599;
  assign n28634 = ~n28630 & ~n28632;
  assign n28635 = ~n28633 & n28634;
  assign n28636 = ~n28631 & n28635;
  assign n28637 = pi17  & n28636;
  assign n28638 = ~pi17  & ~n28636;
  assign n28639 = ~n28637 & ~n28638;
  assign n28640 = n28629 & n28639;
  assign n28641 = ~n28629 & ~n28639;
  assign n28642 = ~n28640 & ~n28641;
  assign n28643 = ~n28470 & n28481;
  assign n28644 = ~n28469 & ~n28643;
  assign n28645 = n28642 & ~n28644;
  assign n28646 = ~n28642 & n28644;
  assign n28647 = ~n28645 & ~n28646;
  assign n28648 = n6630 & n25853;
  assign n28649 = n6631 & n26347;
  assign n28650 = n7238 & n26094;
  assign n28651 = n7262 & n26341;
  assign n28652 = ~n28648 & ~n28650;
  assign n28653 = ~n28651 & n28652;
  assign n28654 = ~n28649 & n28653;
  assign n28655 = pi14  & n28654;
  assign n28656 = ~pi14  & ~n28654;
  assign n28657 = ~n28655 & ~n28656;
  assign n28658 = ~n28488 & n28499;
  assign n28659 = ~n28487 & ~n28658;
  assign n28660 = n28657 & n28659;
  assign n28661 = ~n28657 & ~n28659;
  assign n28662 = ~n28660 & ~n28661;
  assign n28663 = ~n28647 & n28662;
  assign n28664 = n28647 & ~n28662;
  assign n28665 = ~n28663 & ~n28664;
  assign n28666 = ~n28364 & ~n28502;
  assign n28667 = ~n28365 & ~n28666;
  assign n28668 = n28665 & n28667;
  assign n28669 = ~n28665 & ~n28667;
  assign n28670 = ~n28668 & ~n28669;
  assign n28671 = ~n28518 & n28670;
  assign n28672 = n28518 & ~n28670;
  assign n28673 = ~n28671 & ~n28672;
  assign n28674 = ~n28515 & ~n28673;
  assign n28675 = n28515 & n28673;
  assign po16  = ~n28674 & ~n28675;
  assign n28677 = ~n28668 & ~n28671;
  assign n28678 = ~n28657 & n28659;
  assign n28679 = ~n28664 & ~n28678;
  assign n28680 = n28629 & ~n28639;
  assign n28681 = ~n28646 & ~n28680;
  assign n28682 = ~n28621 & n28623;
  assign n28683 = ~n28628 & ~n28682;
  assign n28684 = n28593 & ~n28603;
  assign n28685 = ~n28610 & ~n28684;
  assign n28686 = ~n28528 & n28585;
  assign n28687 = ~n28592 & ~n28686;
  assign n28688 = n28565 & ~n28572;
  assign n28689 = ~n28575 & ~n28576;
  assign n28690 = ~n28688 & ~n28689;
  assign n28691 = ~n28561 & ~n28563;
  assign n28692 = ~n159 & ~n216;
  assign n28693 = ~n937 & n28692;
  assign n28694 = n1004 & n1755;
  assign n28695 = n2253 & n2839;
  assign n28696 = n3123 & n28695;
  assign n28697 = n28693 & n28694;
  assign n28698 = n2357 & n3661;
  assign n28699 = n28697 & n28698;
  assign n28700 = n12855 & n28696;
  assign n28701 = n28699 & n28700;
  assign n28702 = n26193 & n26662;
  assign n28703 = n28701 & n28702;
  assign n28704 = n13066 & n28703;
  assign n28705 = n14397 & n28704;
  assign n28706 = ~n28691 & n28705;
  assign n28707 = n28691 & ~n28705;
  assign n28708 = ~n28706 & ~n28707;
  assign n28709 = n748 & n21030;
  assign n28710 = n880 & n22654;
  assign n28711 = n3692 & n21027;
  assign n28712 = n3694 & n21024;
  assign n28713 = ~n28709 & ~n28711;
  assign n28714 = ~n28712 & n28713;
  assign n28715 = ~n28710 & n28714;
  assign n28716 = n28708 & ~n28715;
  assign n28717 = ~n28708 & n28715;
  assign n28718 = ~n28716 & ~n28717;
  assign n28719 = n28690 & ~n28718;
  assign n28720 = ~n28690 & n28718;
  assign n28721 = ~n28719 & ~n28720;
  assign n28722 = n3810 & n21021;
  assign n28723 = n3886 & n23220;
  assign n28724 = n3884 & n21018;
  assign n28725 = n4380 & n21015;
  assign n28726 = ~n28722 & ~n28724;
  assign n28727 = ~n28725 & n28726;
  assign n28728 = ~n28723 & n28727;
  assign n28729 = pi29  & n28728;
  assign n28730 = ~pi29  & ~n28728;
  assign n28731 = ~n28729 & ~n28730;
  assign n28732 = n28721 & ~n28731;
  assign n28733 = ~n28721 & n28731;
  assign n28734 = ~n28732 & ~n28733;
  assign n28735 = n28538 & ~n28580;
  assign n28736 = ~n28581 & ~n28735;
  assign n28737 = n28734 & n28736;
  assign n28738 = ~n28734 & ~n28736;
  assign n28739 = ~n28737 & ~n28738;
  assign n28740 = n86 & n21012;
  assign n28741 = n4420 & n23812;
  assign n28742 = n4600 & n21009;
  assign n28743 = n4615 & n21006;
  assign n28744 = ~n28740 & ~n28742;
  assign n28745 = ~n28743 & n28744;
  assign n28746 = ~n28741 & n28745;
  assign n28747 = pi26  & n28746;
  assign n28748 = ~pi26  & ~n28746;
  assign n28749 = ~n28747 & ~n28748;
  assign n28750 = n28739 & ~n28749;
  assign n28751 = ~n28739 & n28749;
  assign n28752 = ~n28750 & ~n28751;
  assign n28753 = n28687 & ~n28752;
  assign n28754 = ~n28687 & n28752;
  assign n28755 = ~n28753 & ~n28754;
  assign n28756 = n5044 & n20906;
  assign n28757 = n5045 & n21294;
  assign n28758 = n5109 & n21003;
  assign n28759 = n5130 & n21288;
  assign n28760 = ~n28756 & ~n28758;
  assign n28761 = ~n28759 & n28760;
  assign n28762 = ~n28757 & n28761;
  assign n28763 = pi23  & n28762;
  assign n28764 = ~pi23  & ~n28762;
  assign n28765 = ~n28763 & ~n28764;
  assign n28766 = n28755 & ~n28765;
  assign n28767 = ~n28755 & n28765;
  assign n28768 = ~n28766 & ~n28767;
  assign n28769 = n28685 & ~n28768;
  assign n28770 = ~n28685 & n28768;
  assign n28771 = ~n28769 & ~n28770;
  assign n28772 = n5240 & n24428;
  assign n28773 = n5241 & n24568;
  assign n28774 = n5853 & n24494;
  assign n28775 = n5866 & n24562;
  assign n28776 = ~n28772 & ~n28774;
  assign n28777 = ~n28775 & n28776;
  assign n28778 = ~n28773 & n28777;
  assign n28779 = pi20  & n28778;
  assign n28780 = ~pi20  & ~n28778;
  assign n28781 = ~n28779 & ~n28780;
  assign n28782 = n28771 & ~n28781;
  assign n28783 = ~n28771 & n28781;
  assign n28784 = ~n28782 & ~n28783;
  assign n28785 = n28683 & n28784;
  assign n28786 = ~n28683 & ~n28784;
  assign n28787 = ~n28785 & ~n28786;
  assign n28788 = n5982 & n25336;
  assign n28789 = n5983 & n25859;
  assign n28790 = n6323 & n25599;
  assign n28791 = n6336 & n25853;
  assign n28792 = ~n28788 & ~n28790;
  assign n28793 = ~n28791 & n28792;
  assign n28794 = ~n28789 & n28793;
  assign n28795 = pi17  & n28794;
  assign n28796 = ~pi17  & ~n28794;
  assign n28797 = ~n28795 & ~n28796;
  assign n28798 = ~n28787 & ~n28797;
  assign n28799 = n28787 & n28797;
  assign n28800 = ~n28798 & ~n28799;
  assign n28801 = n28681 & ~n28800;
  assign n28802 = ~n28681 & n28800;
  assign n28803 = ~n28801 & ~n28802;
  assign n28804 = n6630 & n26094;
  assign n28805 = n6631 & n26575;
  assign n28806 = n7238 & n26341;
  assign n28807 = n7262 & n26569;
  assign n28808 = ~n28804 & ~n28806;
  assign n28809 = ~n28807 & n28808;
  assign n28810 = ~n28805 & n28809;
  assign n28811 = pi14  & n28810;
  assign n28812 = ~pi14  & ~n28810;
  assign n28813 = ~n28811 & ~n28812;
  assign n28814 = n28803 & ~n28813;
  assign n28815 = ~n28803 & n28813;
  assign n28816 = ~n28814 & ~n28815;
  assign n28817 = ~n28679 & n28816;
  assign n28818 = n28679 & ~n28816;
  assign n28819 = ~n28817 & ~n28818;
  assign n28820 = n28677 & ~n28819;
  assign n28821 = ~n28677 & n28819;
  assign n28822 = ~n28820 & ~n28821;
  assign n28823 = n28675 & n28822;
  assign n28824 = ~n28675 & ~n28822;
  assign po17  = ~n28823 & ~n28824;
  assign n28826 = ~n28683 & n28784;
  assign n28827 = ~n28798 & ~n28826;
  assign n28828 = ~n14558 & n26569;
  assign n28829 = n6630 & n26341;
  assign n28830 = n6631 & ~n26793;
  assign n28831 = ~n28828 & ~n28829;
  assign n28832 = ~n28830 & n28831;
  assign n28833 = pi14  & n28832;
  assign n28834 = ~pi14  & ~n28832;
  assign n28835 = ~n28833 & ~n28834;
  assign n28836 = ~n28827 & ~n28835;
  assign n28837 = n28827 & n28835;
  assign n28838 = ~n28836 & ~n28837;
  assign n28839 = ~n186 & ~n196;
  assign n28840 = ~n199 & ~n481;
  assign n28841 = ~n499 & ~n511;
  assign n28842 = ~n512 & ~n989;
  assign n28843 = n28841 & n28842;
  assign n28844 = n28839 & n28840;
  assign n28845 = n444 & n527;
  assign n28846 = n1697 & n28845;
  assign n28847 = n28843 & n28844;
  assign n28848 = n28846 & n28847;
  assign n28849 = n390 & n2931;
  assign n28850 = n28848 & n28849;
  assign n28851 = n1025 & n3919;
  assign n28852 = n5658 & n28851;
  assign n28853 = n3199 & n28850;
  assign n28854 = n28852 & n28853;
  assign n28855 = n4246 & n28854;
  assign n28856 = ~n28705 & n28855;
  assign n28857 = n28705 & ~n28855;
  assign n28858 = ~n28856 & ~n28857;
  assign n28859 = n748 & n21027;
  assign n28860 = n880 & n21306;
  assign n28861 = n3692 & n21024;
  assign n28862 = n3694 & n21021;
  assign n28863 = ~n28859 & ~n28861;
  assign n28864 = ~n28862 & n28863;
  assign n28865 = ~n28860 & n28864;
  assign n28866 = n28858 & ~n28865;
  assign n28867 = ~n28858 & n28865;
  assign n28868 = ~n28866 & ~n28867;
  assign n28869 = ~n28706 & n28715;
  assign n28870 = ~n28707 & ~n28869;
  assign n28871 = ~n28868 & ~n28870;
  assign n28872 = n28868 & n28870;
  assign n28873 = ~n28871 & ~n28872;
  assign n28874 = ~n28720 & ~n28732;
  assign n28875 = ~n28873 & n28874;
  assign n28876 = n28873 & ~n28874;
  assign n28877 = ~n28875 & ~n28876;
  assign n28878 = n3810 & n21018;
  assign n28879 = n3886 & n23205;
  assign n28880 = n3884 & n21015;
  assign n28881 = n4380 & n21012;
  assign n28882 = ~n28878 & ~n28880;
  assign n28883 = ~n28881 & n28882;
  assign n28884 = ~n28879 & n28883;
  assign n28885 = pi29  & n28884;
  assign n28886 = ~pi29  & ~n28884;
  assign n28887 = ~n28885 & ~n28886;
  assign n28888 = n28877 & n28887;
  assign n28889 = ~n28877 & ~n28887;
  assign n28890 = ~n28888 & ~n28889;
  assign n28891 = n86 & n21009;
  assign n28892 = n4420 & n23851;
  assign n28893 = n4600 & n21006;
  assign n28894 = n4615 & n20906;
  assign n28895 = ~n28891 & ~n28893;
  assign n28896 = ~n28894 & n28895;
  assign n28897 = ~n28892 & n28896;
  assign n28898 = pi26  & n28897;
  assign n28899 = ~pi26  & ~n28897;
  assign n28900 = ~n28898 & ~n28899;
  assign n28901 = ~n28890 & ~n28900;
  assign n28902 = n28890 & n28900;
  assign n28903 = ~n28901 & ~n28902;
  assign n28904 = ~n28737 & n28749;
  assign n28905 = ~n28738 & ~n28904;
  assign n28906 = ~n28903 & ~n28905;
  assign n28907 = n28903 & n28905;
  assign n28908 = ~n28906 & ~n28907;
  assign n28909 = n5044 & n21003;
  assign n28910 = n5045 & n24596;
  assign n28911 = n5109 & n21288;
  assign n28912 = n5130 & n24428;
  assign n28913 = ~n28909 & ~n28911;
  assign n28914 = ~n28912 & n28913;
  assign n28915 = ~n28910 & n28914;
  assign n28916 = pi23  & n28915;
  assign n28917 = ~pi23  & ~n28915;
  assign n28918 = ~n28916 & ~n28917;
  assign n28919 = n28908 & ~n28918;
  assign n28920 = ~n28908 & n28918;
  assign n28921 = ~n28919 & ~n28920;
  assign n28922 = ~n28754 & n28765;
  assign n28923 = ~n28753 & ~n28922;
  assign n28924 = ~n28921 & ~n28923;
  assign n28925 = n28921 & n28923;
  assign n28926 = ~n28924 & ~n28925;
  assign n28927 = n5240 & n24494;
  assign n28928 = n5241 & n25342;
  assign n28929 = n5853 & n24562;
  assign n28930 = n5866 & n25336;
  assign n28931 = ~n28927 & ~n28929;
  assign n28932 = ~n28930 & n28931;
  assign n28933 = ~n28928 & n28932;
  assign n28934 = pi20  & n28933;
  assign n28935 = ~pi20  & ~n28933;
  assign n28936 = ~n28934 & ~n28935;
  assign n28937 = n28926 & ~n28936;
  assign n28938 = ~n28926 & n28936;
  assign n28939 = ~n28937 & ~n28938;
  assign n28940 = ~n28770 & n28781;
  assign n28941 = ~n28769 & ~n28940;
  assign n28942 = ~n28939 & ~n28941;
  assign n28943 = n28939 & n28941;
  assign n28944 = ~n28942 & ~n28943;
  assign n28945 = n5982 & n25599;
  assign n28946 = n5983 & n26100;
  assign n28947 = n6323 & n25853;
  assign n28948 = n6336 & n26094;
  assign n28949 = ~n28945 & ~n28947;
  assign n28950 = ~n28948 & n28949;
  assign n28951 = ~n28946 & n28950;
  assign n28952 = pi17  & n28951;
  assign n28953 = ~pi17  & ~n28951;
  assign n28954 = ~n28952 & ~n28953;
  assign n28955 = n28944 & ~n28954;
  assign n28956 = ~n28944 & n28954;
  assign n28957 = ~n28955 & ~n28956;
  assign n28958 = n28838 & n28957;
  assign n28959 = ~n28838 & ~n28957;
  assign n28960 = ~n28958 & ~n28959;
  assign n28961 = ~n28802 & n28813;
  assign n28962 = ~n28801 & ~n28961;
  assign n28963 = ~n28960 & ~n28962;
  assign n28964 = n28960 & n28962;
  assign n28965 = ~n28963 & ~n28964;
  assign n28966 = ~n28817 & ~n28821;
  assign n28967 = ~n28965 & n28966;
  assign n28968 = n28965 & ~n28966;
  assign n28969 = ~n28967 & ~n28968;
  assign n28970 = n28823 & n28969;
  assign n28971 = ~n28823 & ~n28969;
  assign po18  = ~n28970 & ~n28971;
  assign n28973 = ~n28964 & ~n28968;
  assign n28974 = ~n28872 & ~n28876;
  assign n28975 = n3810 & n21015;
  assign n28976 = n3886 & n23190;
  assign n28977 = n3884 & n21012;
  assign n28978 = n4380 & n21009;
  assign n28979 = ~n28975 & ~n28977;
  assign n28980 = ~n28978 & n28979;
  assign n28981 = ~n28976 & n28980;
  assign n28982 = pi29  & n28981;
  assign n28983 = ~pi29  & ~n28981;
  assign n28984 = ~n28982 & ~n28983;
  assign n28985 = ~n28857 & ~n28866;
  assign n28986 = ~n12996 & n26569;
  assign n28987 = pi14  & ~n28986;
  assign n28988 = ~pi14  & n28986;
  assign n28989 = ~n28987 & ~n28988;
  assign n28990 = ~n361 & n1421;
  assign n28991 = n2007 & n2682;
  assign n28992 = n28990 & n28991;
  assign n28993 = n1406 & n3256;
  assign n28994 = n4166 & n28993;
  assign n28995 = n13588 & n28992;
  assign n28996 = n28994 & n28995;
  assign n28997 = n1946 & n7067;
  assign n28998 = n28996 & n28997;
  assign n28999 = n13334 & n28998;
  assign n29000 = n2233 & n28999;
  assign n29001 = n28705 & n29000;
  assign n29002 = ~n28705 & ~n29000;
  assign n29003 = ~n29001 & ~n29002;
  assign n29004 = n28989 & n29003;
  assign n29005 = ~n28989 & ~n29003;
  assign n29006 = ~n29004 & ~n29005;
  assign n29007 = ~n28985 & n29006;
  assign n29008 = n28985 & ~n29006;
  assign n29009 = ~n29007 & ~n29008;
  assign n29010 = n748 & n21024;
  assign n29011 = n880 & n23033;
  assign n29012 = n3692 & n21021;
  assign n29013 = n3694 & n21018;
  assign n29014 = ~n29010 & ~n29012;
  assign n29015 = ~n29013 & n29014;
  assign n29016 = ~n29011 & n29015;
  assign n29017 = n29009 & ~n29016;
  assign n29018 = ~n29009 & n29016;
  assign n29019 = ~n29017 & ~n29018;
  assign n29020 = ~n28984 & n29019;
  assign n29021 = n28984 & ~n29019;
  assign n29022 = ~n29020 & ~n29021;
  assign n29023 = n28974 & ~n29022;
  assign n29024 = ~n28974 & n29022;
  assign n29025 = ~n29023 & ~n29024;
  assign n29026 = n86 & n21006;
  assign n29027 = n4420 & n23833;
  assign n29028 = n4600 & n20906;
  assign n29029 = n4615 & n21003;
  assign n29030 = ~n29026 & ~n29028;
  assign n29031 = ~n29029 & n29030;
  assign n29032 = ~n29027 & n29031;
  assign n29033 = pi26  & n29032;
  assign n29034 = ~pi26  & ~n29032;
  assign n29035 = ~n29033 & ~n29034;
  assign n29036 = n29025 & n29035;
  assign n29037 = ~n29025 & ~n29035;
  assign n29038 = ~n29036 & ~n29037;
  assign n29039 = n28877 & ~n28887;
  assign n29040 = ~n28901 & ~n29039;
  assign n29041 = n29038 & n29040;
  assign n29042 = ~n29038 & ~n29040;
  assign n29043 = ~n29041 & ~n29042;
  assign n29044 = n5044 & n21288;
  assign n29045 = n5045 & n24584;
  assign n29046 = n5109 & n24428;
  assign n29047 = n5130 & n24494;
  assign n29048 = ~n29044 & ~n29046;
  assign n29049 = ~n29047 & n29048;
  assign n29050 = ~n29045 & n29049;
  assign n29051 = pi23  & n29050;
  assign n29052 = ~pi23  & ~n29050;
  assign n29053 = ~n29051 & ~n29052;
  assign n29054 = ~n28907 & n28918;
  assign n29055 = ~n28906 & ~n29054;
  assign n29056 = n29053 & n29055;
  assign n29057 = ~n29053 & ~n29055;
  assign n29058 = ~n29056 & ~n29057;
  assign n29059 = ~n29043 & n29058;
  assign n29060 = n29043 & ~n29058;
  assign n29061 = ~n29059 & ~n29060;
  assign n29062 = n5240 & n24562;
  assign n29063 = n5241 & n25605;
  assign n29064 = n5853 & n25336;
  assign n29065 = n5866 & n25599;
  assign n29066 = ~n29062 & ~n29064;
  assign n29067 = ~n29065 & n29066;
  assign n29068 = ~n29063 & n29067;
  assign n29069 = pi20  & n29068;
  assign n29070 = ~pi20  & ~n29068;
  assign n29071 = ~n29069 & ~n29070;
  assign n29072 = n29061 & n29071;
  assign n29073 = ~n29061 & ~n29071;
  assign n29074 = ~n29072 & ~n29073;
  assign n29075 = ~n28925 & n28936;
  assign n29076 = ~n28924 & ~n29075;
  assign n29077 = n29074 & ~n29076;
  assign n29078 = ~n29074 & n29076;
  assign n29079 = ~n29077 & ~n29078;
  assign n29080 = n5982 & n25853;
  assign n29081 = n5983 & n26347;
  assign n29082 = n6323 & n26094;
  assign n29083 = n6336 & n26341;
  assign n29084 = ~n29080 & ~n29082;
  assign n29085 = ~n29083 & n29084;
  assign n29086 = ~n29081 & n29085;
  assign n29087 = pi17  & n29086;
  assign n29088 = ~pi17  & ~n29086;
  assign n29089 = ~n29087 & ~n29088;
  assign n29090 = ~n28943 & n28954;
  assign n29091 = ~n28942 & ~n29090;
  assign n29092 = n29089 & n29091;
  assign n29093 = ~n29089 & ~n29091;
  assign n29094 = ~n29092 & ~n29093;
  assign n29095 = ~n29079 & n29094;
  assign n29096 = n29079 & ~n29094;
  assign n29097 = ~n29095 & ~n29096;
  assign n29098 = ~n28836 & ~n28957;
  assign n29099 = ~n28837 & ~n29098;
  assign n29100 = n29097 & n29099;
  assign n29101 = ~n29097 & ~n29099;
  assign n29102 = ~n29100 & ~n29101;
  assign n29103 = ~n28973 & n29102;
  assign n29104 = n28973 & ~n29102;
  assign n29105 = ~n29103 & ~n29104;
  assign n29106 = ~n28970 & ~n29105;
  assign n29107 = n28970 & n29105;
  assign po19  = ~n29106 & ~n29107;
  assign n29109 = ~n29100 & ~n29103;
  assign n29110 = ~n29089 & n29091;
  assign n29111 = ~n29096 & ~n29110;
  assign n29112 = n29061 & ~n29071;
  assign n29113 = ~n29078 & ~n29112;
  assign n29114 = ~n29053 & n29055;
  assign n29115 = ~n29060 & ~n29114;
  assign n29116 = n29025 & ~n29035;
  assign n29117 = ~n29042 & ~n29116;
  assign n29118 = ~n29020 & ~n29024;
  assign n29119 = ~n29002 & ~n29004;
  assign n29120 = ~n184 & ~n296;
  assign n29121 = n366 & n29120;
  assign n29122 = n1006 & n1947;
  assign n29123 = n2108 & n2608;
  assign n29124 = n15037 & n29123;
  assign n29125 = n23087 & n29122;
  assign n29126 = n2322 & n29121;
  assign n29127 = n29125 & n29126;
  assign n29128 = n1016 & n29124;
  assign n29129 = n29127 & n29128;
  assign n29130 = n6195 & n13635;
  assign n29131 = n29129 & n29130;
  assign n29132 = n5507 & n29131;
  assign n29133 = n3457 & n29132;
  assign n29134 = ~n29119 & n29133;
  assign n29135 = n29119 & ~n29133;
  assign n29136 = ~n29134 & ~n29135;
  assign n29137 = n748 & n21021;
  assign n29138 = n880 & n23220;
  assign n29139 = n3692 & n21018;
  assign n29140 = n3694 & n21015;
  assign n29141 = ~n29137 & ~n29139;
  assign n29142 = ~n29140 & n29141;
  assign n29143 = ~n29138 & n29142;
  assign n29144 = n29136 & ~n29143;
  assign n29145 = ~n29136 & n29143;
  assign n29146 = ~n29144 & ~n29145;
  assign n29147 = ~n29007 & n29016;
  assign n29148 = ~n29008 & ~n29147;
  assign n29149 = ~n29146 & ~n29148;
  assign n29150 = n29146 & n29148;
  assign n29151 = ~n29149 & ~n29150;
  assign n29152 = n3810 & n21012;
  assign n29153 = n3886 & n23812;
  assign n29154 = n3884 & n21009;
  assign n29155 = n4380 & n21006;
  assign n29156 = ~n29152 & ~n29154;
  assign n29157 = ~n29155 & n29156;
  assign n29158 = ~n29153 & n29157;
  assign n29159 = pi29  & n29158;
  assign n29160 = ~pi29  & ~n29158;
  assign n29161 = ~n29159 & ~n29160;
  assign n29162 = n29151 & ~n29161;
  assign n29163 = ~n29151 & n29161;
  assign n29164 = ~n29162 & ~n29163;
  assign n29165 = ~n29118 & n29164;
  assign n29166 = n29118 & ~n29164;
  assign n29167 = ~n29165 & ~n29166;
  assign n29168 = n86 & n20906;
  assign n29169 = n4420 & n21294;
  assign n29170 = n4600 & n21003;
  assign n29171 = n4615 & n21288;
  assign n29172 = ~n29168 & ~n29170;
  assign n29173 = ~n29171 & n29172;
  assign n29174 = ~n29169 & n29173;
  assign n29175 = pi26  & n29174;
  assign n29176 = ~pi26  & ~n29174;
  assign n29177 = ~n29175 & ~n29176;
  assign n29178 = n29167 & ~n29177;
  assign n29179 = ~n29167 & n29177;
  assign n29180 = ~n29178 & ~n29179;
  assign n29181 = n29117 & ~n29180;
  assign n29182 = ~n29117 & n29180;
  assign n29183 = ~n29181 & ~n29182;
  assign n29184 = n5044 & n24428;
  assign n29185 = n5045 & n24568;
  assign n29186 = n5109 & n24494;
  assign n29187 = n5130 & n24562;
  assign n29188 = ~n29184 & ~n29186;
  assign n29189 = ~n29187 & n29188;
  assign n29190 = ~n29185 & n29189;
  assign n29191 = pi23  & n29190;
  assign n29192 = ~pi23  & ~n29190;
  assign n29193 = ~n29191 & ~n29192;
  assign n29194 = n29183 & ~n29193;
  assign n29195 = ~n29183 & n29193;
  assign n29196 = ~n29194 & ~n29195;
  assign n29197 = n29115 & n29196;
  assign n29198 = ~n29115 & ~n29196;
  assign n29199 = ~n29197 & ~n29198;
  assign n29200 = n5240 & n25336;
  assign n29201 = n5241 & n25859;
  assign n29202 = n5853 & n25599;
  assign n29203 = n5866 & n25853;
  assign n29204 = ~n29200 & ~n29202;
  assign n29205 = ~n29203 & n29204;
  assign n29206 = ~n29201 & n29205;
  assign n29207 = pi20  & n29206;
  assign n29208 = ~pi20  & ~n29206;
  assign n29209 = ~n29207 & ~n29208;
  assign n29210 = ~n29199 & ~n29209;
  assign n29211 = n29199 & n29209;
  assign n29212 = ~n29210 & ~n29211;
  assign n29213 = n29113 & ~n29212;
  assign n29214 = ~n29113 & n29212;
  assign n29215 = ~n29213 & ~n29214;
  assign n29216 = n5982 & n26094;
  assign n29217 = n5983 & n26575;
  assign n29218 = n6323 & n26341;
  assign n29219 = n6336 & n26569;
  assign n29220 = ~n29216 & ~n29218;
  assign n29221 = ~n29219 & n29220;
  assign n29222 = ~n29217 & n29221;
  assign n29223 = pi17  & n29222;
  assign n29224 = ~pi17  & ~n29222;
  assign n29225 = ~n29223 & ~n29224;
  assign n29226 = n29215 & ~n29225;
  assign n29227 = ~n29215 & n29225;
  assign n29228 = ~n29226 & ~n29227;
  assign n29229 = ~n29111 & n29228;
  assign n29230 = n29111 & ~n29228;
  assign n29231 = ~n29229 & ~n29230;
  assign n29232 = n29109 & ~n29231;
  assign n29233 = ~n29109 & n29231;
  assign n29234 = ~n29232 & ~n29233;
  assign n29235 = n29107 & n29234;
  assign n29236 = ~n29107 & ~n29234;
  assign po20  = ~n29235 & ~n29236;
  assign n29238 = ~n29115 & n29196;
  assign n29239 = ~n29210 & ~n29238;
  assign n29240 = ~n13908 & n26569;
  assign n29241 = n5982 & n26341;
  assign n29242 = n5983 & ~n26793;
  assign n29243 = ~n29240 & ~n29241;
  assign n29244 = ~n29242 & n29243;
  assign n29245 = pi17  & n29244;
  assign n29246 = ~pi17  & ~n29244;
  assign n29247 = ~n29245 & ~n29246;
  assign n29248 = ~n29239 & ~n29247;
  assign n29249 = n29239 & n29247;
  assign n29250 = ~n29248 & ~n29249;
  assign n29251 = ~n29150 & ~n29162;
  assign n29252 = ~n307 & ~n437;
  assign n29253 = n413 & n29252;
  assign n29254 = ~n126 & ~n168;
  assign n29255 = ~n510 & ~n1086;
  assign n29256 = n29254 & n29255;
  assign n29257 = n1359 & n1488;
  assign n29258 = n1579 & n2253;
  assign n29259 = n2658 & n2801;
  assign n29260 = n29258 & n29259;
  assign n29261 = n29256 & n29257;
  assign n29262 = n29253 & n29261;
  assign n29263 = n806 & n29260;
  assign n29264 = n3223 & n29263;
  assign n29265 = n29262 & n29264;
  assign n29266 = n498 & n29265;
  assign n29267 = n2075 & n5645;
  assign n29268 = n29266 & n29267;
  assign n29269 = n29133 & ~n29268;
  assign n29270 = ~n29133 & n29268;
  assign n29271 = ~n29269 & ~n29270;
  assign n29272 = ~n29134 & n29143;
  assign n29273 = ~n29135 & ~n29272;
  assign n29274 = n29271 & n29273;
  assign n29275 = ~n29271 & ~n29273;
  assign n29276 = ~n29274 & ~n29275;
  assign n29277 = n748 & n21018;
  assign n29278 = n880 & n23205;
  assign n29279 = n3692 & n21015;
  assign n29280 = n3694 & n21012;
  assign n29281 = ~n29277 & ~n29279;
  assign n29282 = ~n29280 & n29281;
  assign n29283 = ~n29278 & n29282;
  assign n29284 = n29276 & n29283;
  assign n29285 = ~n29276 & ~n29283;
  assign n29286 = ~n29284 & ~n29285;
  assign n29287 = n3810 & n21009;
  assign n29288 = n3886 & n23851;
  assign n29289 = n3884 & n21006;
  assign n29290 = n4380 & n20906;
  assign n29291 = ~n29287 & ~n29289;
  assign n29292 = ~n29290 & n29291;
  assign n29293 = ~n29288 & n29292;
  assign n29294 = pi29  & n29293;
  assign n29295 = ~pi29  & ~n29293;
  assign n29296 = ~n29294 & ~n29295;
  assign n29297 = ~n29286 & ~n29296;
  assign n29298 = n29286 & n29296;
  assign n29299 = ~n29297 & ~n29298;
  assign n29300 = ~n29251 & n29299;
  assign n29301 = n29251 & ~n29299;
  assign n29302 = ~n29300 & ~n29301;
  assign n29303 = n86 & n21003;
  assign n29304 = n4420 & n24596;
  assign n29305 = n4600 & n21288;
  assign n29306 = n4615 & n24428;
  assign n29307 = ~n29303 & ~n29305;
  assign n29308 = ~n29306 & n29307;
  assign n29309 = ~n29304 & n29308;
  assign n29310 = pi26  & n29309;
  assign n29311 = ~pi26  & ~n29309;
  assign n29312 = ~n29310 & ~n29311;
  assign n29313 = n29302 & ~n29312;
  assign n29314 = ~n29302 & n29312;
  assign n29315 = ~n29313 & ~n29314;
  assign n29316 = ~n29165 & n29177;
  assign n29317 = ~n29166 & ~n29316;
  assign n29318 = ~n29315 & ~n29317;
  assign n29319 = n29315 & n29317;
  assign n29320 = ~n29318 & ~n29319;
  assign n29321 = n5044 & n24494;
  assign n29322 = n5045 & n25342;
  assign n29323 = n5109 & n24562;
  assign n29324 = n5130 & n25336;
  assign n29325 = ~n29321 & ~n29323;
  assign n29326 = ~n29324 & n29325;
  assign n29327 = ~n29322 & n29326;
  assign n29328 = pi23  & n29327;
  assign n29329 = ~pi23  & ~n29327;
  assign n29330 = ~n29328 & ~n29329;
  assign n29331 = n29320 & ~n29330;
  assign n29332 = ~n29320 & n29330;
  assign n29333 = ~n29331 & ~n29332;
  assign n29334 = ~n29182 & n29193;
  assign n29335 = ~n29181 & ~n29334;
  assign n29336 = ~n29333 & ~n29335;
  assign n29337 = n29333 & n29335;
  assign n29338 = ~n29336 & ~n29337;
  assign n29339 = n5240 & n25599;
  assign n29340 = n5241 & n26100;
  assign n29341 = n5853 & n25853;
  assign n29342 = n5866 & n26094;
  assign n29343 = ~n29339 & ~n29341;
  assign n29344 = ~n29342 & n29343;
  assign n29345 = ~n29340 & n29344;
  assign n29346 = pi20  & n29345;
  assign n29347 = ~pi20  & ~n29345;
  assign n29348 = ~n29346 & ~n29347;
  assign n29349 = n29338 & ~n29348;
  assign n29350 = ~n29338 & n29348;
  assign n29351 = ~n29349 & ~n29350;
  assign n29352 = n29250 & n29351;
  assign n29353 = ~n29250 & ~n29351;
  assign n29354 = ~n29352 & ~n29353;
  assign n29355 = ~n29214 & n29225;
  assign n29356 = ~n29213 & ~n29355;
  assign n29357 = ~n29354 & ~n29356;
  assign n29358 = n29354 & n29356;
  assign n29359 = ~n29357 & ~n29358;
  assign n29360 = ~n29229 & ~n29233;
  assign n29361 = ~n29359 & n29360;
  assign n29362 = n29359 & ~n29360;
  assign n29363 = ~n29361 & ~n29362;
  assign n29364 = n29235 & n29363;
  assign n29365 = ~n29235 & ~n29363;
  assign po21  = ~n29364 & ~n29365;
  assign n29367 = ~n29358 & ~n29362;
  assign n29368 = n5044 & n24562;
  assign n29369 = n5045 & n25605;
  assign n29370 = n5109 & n25336;
  assign n29371 = n5130 & n25599;
  assign n29372 = ~n29368 & ~n29370;
  assign n29373 = ~n29371 & n29372;
  assign n29374 = ~n29369 & n29373;
  assign n29375 = pi23  & n29374;
  assign n29376 = ~pi23  & ~n29374;
  assign n29377 = ~n29375 & ~n29376;
  assign n29378 = n86 & n21288;
  assign n29379 = n4420 & n24584;
  assign n29380 = n4600 & n24428;
  assign n29381 = n4615 & n24494;
  assign n29382 = ~n29378 & ~n29380;
  assign n29383 = ~n29381 & n29382;
  assign n29384 = ~n29379 & n29383;
  assign n29385 = pi26  & n29384;
  assign n29386 = ~pi26  & ~n29384;
  assign n29387 = ~n29385 & ~n29386;
  assign n29388 = ~n29300 & n29312;
  assign n29389 = ~n29301 & ~n29388;
  assign n29390 = n29387 & n29389;
  assign n29391 = ~n29387 & ~n29389;
  assign n29392 = ~n29390 & ~n29391;
  assign n29393 = n3810 & n21006;
  assign n29394 = n3886 & n23833;
  assign n29395 = n3884 & n20906;
  assign n29396 = n4380 & n21003;
  assign n29397 = ~n29393 & ~n29395;
  assign n29398 = ~n29396 & n29397;
  assign n29399 = ~n29394 & n29398;
  assign n29400 = pi29  & n29399;
  assign n29401 = ~pi29  & ~n29399;
  assign n29402 = ~n29400 & ~n29401;
  assign n29403 = n29276 & ~n29283;
  assign n29404 = ~n29297 & ~n29403;
  assign n29405 = ~n12787 & n26569;
  assign n29406 = pi17  & ~n29405;
  assign n29407 = ~pi17  & n29405;
  assign n29408 = ~n29406 & ~n29407;
  assign n29409 = ~n168 & ~n435;
  assign n29410 = ~n459 & n29409;
  assign n29411 = n567 & n1843;
  assign n29412 = n29410 & n29411;
  assign n29413 = n2003 & n23083;
  assign n29414 = n29412 & n29413;
  assign n29415 = n1889 & n3435;
  assign n29416 = n12799 & n29415;
  assign n29417 = n29414 & n29416;
  assign n29418 = n1595 & n29417;
  assign n29419 = n4491 & n5286;
  assign n29420 = n29418 & n29419;
  assign n29421 = n29268 & n29420;
  assign n29422 = ~n29268 & ~n29420;
  assign n29423 = ~n29421 & ~n29422;
  assign n29424 = n29408 & n29423;
  assign n29425 = ~n29408 & ~n29423;
  assign n29426 = ~n29424 & ~n29425;
  assign n29427 = n748 & n21015;
  assign n29428 = n880 & n23190;
  assign n29429 = n3692 & n21012;
  assign n29430 = n3694 & n21009;
  assign n29431 = ~n29427 & ~n29429;
  assign n29432 = ~n29430 & n29431;
  assign n29433 = ~n29428 & n29432;
  assign n29434 = n29426 & n29433;
  assign n29435 = ~n29426 & ~n29433;
  assign n29436 = ~n29434 & ~n29435;
  assign n29437 = ~n29270 & ~n29274;
  assign n29438 = ~n29436 & n29437;
  assign n29439 = n29436 & ~n29437;
  assign n29440 = ~n29438 & ~n29439;
  assign n29441 = ~n29404 & ~n29440;
  assign n29442 = n29404 & n29440;
  assign n29443 = ~n29441 & ~n29442;
  assign n29444 = n29402 & ~n29443;
  assign n29445 = ~n29402 & n29443;
  assign n29446 = ~n29444 & ~n29445;
  assign n29447 = ~n29392 & n29446;
  assign n29448 = n29392 & ~n29446;
  assign n29449 = ~n29447 & ~n29448;
  assign n29450 = ~n29377 & n29449;
  assign n29451 = n29377 & ~n29449;
  assign n29452 = ~n29450 & ~n29451;
  assign n29453 = ~n29319 & n29330;
  assign n29454 = ~n29318 & ~n29453;
  assign n29455 = ~n29452 & ~n29454;
  assign n29456 = n29452 & n29454;
  assign n29457 = ~n29455 & ~n29456;
  assign n29458 = n5240 & n25853;
  assign n29459 = n5241 & n26347;
  assign n29460 = n5853 & n26094;
  assign n29461 = n5866 & n26341;
  assign n29462 = ~n29458 & ~n29460;
  assign n29463 = ~n29461 & n29462;
  assign n29464 = ~n29459 & n29463;
  assign n29465 = pi20  & n29464;
  assign n29466 = ~pi20  & ~n29464;
  assign n29467 = ~n29465 & ~n29466;
  assign n29468 = ~n29337 & n29348;
  assign n29469 = ~n29336 & ~n29468;
  assign n29470 = n29467 & n29469;
  assign n29471 = ~n29467 & ~n29469;
  assign n29472 = ~n29470 & ~n29471;
  assign n29473 = ~n29457 & n29472;
  assign n29474 = n29457 & ~n29472;
  assign n29475 = ~n29473 & ~n29474;
  assign n29476 = ~n29248 & ~n29351;
  assign n29477 = ~n29249 & ~n29476;
  assign n29478 = n29475 & n29477;
  assign n29479 = ~n29475 & ~n29477;
  assign n29480 = ~n29478 & ~n29479;
  assign n29481 = ~n29367 & n29480;
  assign n29482 = n29367 & ~n29480;
  assign n29483 = ~n29481 & ~n29482;
  assign n29484 = ~n29364 & ~n29483;
  assign n29485 = n29364 & n29483;
  assign po22  = ~n29484 & ~n29485;
  assign n29487 = ~n29467 & n29469;
  assign n29488 = ~n29474 & ~n29487;
  assign n29489 = ~n29450 & ~n29456;
  assign n29490 = n5044 & n25336;
  assign n29491 = n5045 & n25859;
  assign n29492 = n5109 & n25599;
  assign n29493 = n5130 & n25853;
  assign n29494 = ~n29490 & ~n29492;
  assign n29495 = ~n29493 & n29494;
  assign n29496 = ~n29491 & n29495;
  assign n29497 = pi23  & n29496;
  assign n29498 = ~pi23  & ~n29496;
  assign n29499 = ~n29497 & ~n29498;
  assign n29500 = ~n29387 & n29389;
  assign n29501 = ~n29447 & ~n29500;
  assign n29502 = n29426 & ~n29433;
  assign n29503 = ~n29436 & ~n29437;
  assign n29504 = ~n29502 & ~n29503;
  assign n29505 = ~n29422 & ~n29424;
  assign n29506 = ~n177 & ~n303;
  assign n29507 = ~n703 & ~n792;
  assign n29508 = n1480 & n29507;
  assign n29509 = n479 & n29506;
  assign n29510 = n1575 & n1652;
  assign n29511 = n4687 & n29510;
  assign n29512 = n29508 & n29509;
  assign n29513 = n3352 & n12716;
  assign n29514 = n29512 & n29513;
  assign n29515 = n29511 & n29514;
  assign n29516 = n1290 & n3261;
  assign n29517 = n29515 & n29516;
  assign n29518 = n6842 & n29517;
  assign n29519 = n27839 & n29518;
  assign n29520 = ~n29505 & n29519;
  assign n29521 = n29505 & ~n29519;
  assign n29522 = ~n29520 & ~n29521;
  assign n29523 = n748 & n21012;
  assign n29524 = n880 & n23812;
  assign n29525 = n3692 & n21009;
  assign n29526 = n3694 & n21006;
  assign n29527 = ~n29523 & ~n29525;
  assign n29528 = ~n29526 & n29527;
  assign n29529 = ~n29524 & n29528;
  assign n29530 = n29522 & ~n29529;
  assign n29531 = ~n29522 & n29529;
  assign n29532 = ~n29530 & ~n29531;
  assign n29533 = n29504 & ~n29532;
  assign n29534 = ~n29504 & n29532;
  assign n29535 = ~n29533 & ~n29534;
  assign n29536 = n3810 & n20906;
  assign n29537 = n3886 & n21294;
  assign n29538 = n3884 & n21003;
  assign n29539 = n4380 & n21288;
  assign n29540 = ~n29536 & ~n29538;
  assign n29541 = ~n29539 & n29540;
  assign n29542 = ~n29537 & n29541;
  assign n29543 = pi29  & n29542;
  assign n29544 = ~pi29  & ~n29542;
  assign n29545 = ~n29543 & ~n29544;
  assign n29546 = n29535 & ~n29545;
  assign n29547 = ~n29535 & n29545;
  assign n29548 = ~n29546 & ~n29547;
  assign n29549 = n29402 & ~n29441;
  assign n29550 = ~n29442 & ~n29549;
  assign n29551 = n29548 & n29550;
  assign n29552 = ~n29548 & ~n29550;
  assign n29553 = ~n29551 & ~n29552;
  assign n29554 = n86 & n24428;
  assign n29555 = n4420 & n24568;
  assign n29556 = n4600 & n24494;
  assign n29557 = n4615 & n24562;
  assign n29558 = ~n29554 & ~n29556;
  assign n29559 = ~n29557 & n29558;
  assign n29560 = ~n29555 & n29559;
  assign n29561 = pi26  & n29560;
  assign n29562 = ~pi26  & ~n29560;
  assign n29563 = ~n29561 & ~n29562;
  assign n29564 = n29553 & ~n29563;
  assign n29565 = ~n29553 & n29563;
  assign n29566 = ~n29564 & ~n29565;
  assign n29567 = ~n29501 & n29566;
  assign n29568 = n29501 & ~n29566;
  assign n29569 = ~n29567 & ~n29568;
  assign n29570 = n29499 & ~n29569;
  assign n29571 = ~n29499 & n29569;
  assign n29572 = ~n29570 & ~n29571;
  assign n29573 = n29489 & ~n29572;
  assign n29574 = ~n29489 & n29572;
  assign n29575 = ~n29573 & ~n29574;
  assign n29576 = n5240 & n26094;
  assign n29577 = n5241 & n26575;
  assign n29578 = n5853 & n26341;
  assign n29579 = n5866 & n26569;
  assign n29580 = ~n29576 & ~n29578;
  assign n29581 = ~n29579 & n29580;
  assign n29582 = ~n29577 & n29581;
  assign n29583 = pi20  & n29582;
  assign n29584 = ~pi20  & ~n29582;
  assign n29585 = ~n29583 & ~n29584;
  assign n29586 = n29575 & ~n29585;
  assign n29587 = ~n29575 & n29585;
  assign n29588 = ~n29586 & ~n29587;
  assign n29589 = n29488 & n29588;
  assign n29590 = ~n29488 & ~n29588;
  assign n29591 = ~n29589 & ~n29590;
  assign n29592 = ~n29478 & ~n29481;
  assign n29593 = n29591 & n29592;
  assign n29594 = ~n29591 & ~n29592;
  assign n29595 = ~n29593 & ~n29594;
  assign n29596 = n29485 & n29595;
  assign n29597 = ~n29485 & ~n29595;
  assign po23  = ~n29596 & ~n29597;
  assign n29599 = ~n13283 & n26569;
  assign n29600 = n5240 & n26341;
  assign n29601 = n5241 & ~n26793;
  assign n29602 = ~n29599 & ~n29600;
  assign n29603 = ~n29601 & n29602;
  assign n29604 = pi20  & n29603;
  assign n29605 = ~pi20  & ~n29603;
  assign n29606 = ~n29604 & ~n29605;
  assign n29607 = n29499 & ~n29567;
  assign n29608 = ~n29568 & ~n29607;
  assign n29609 = ~n29606 & n29608;
  assign n29610 = n29606 & ~n29608;
  assign n29611 = ~n29609 & ~n29610;
  assign n29612 = ~n376 & ~n503;
  assign n29613 = n431 & n29612;
  assign n29614 = n1452 & n3444;
  assign n29615 = n12962 & n29614;
  assign n29616 = n12820 & n29613;
  assign n29617 = n29253 & n29616;
  assign n29618 = n29615 & n29617;
  assign n29619 = n4471 & n27017;
  assign n29620 = n29618 & n29619;
  assign n29621 = n4933 & n6885;
  assign n29622 = n29620 & n29621;
  assign n29623 = n1607 & n29622;
  assign n29624 = ~n29519 & n29623;
  assign n29625 = n29519 & ~n29623;
  assign n29626 = ~n29624 & ~n29625;
  assign n29627 = n748 & n21009;
  assign n29628 = n880 & n23851;
  assign n29629 = n3692 & n21006;
  assign n29630 = n3694 & n20906;
  assign n29631 = ~n29627 & ~n29629;
  assign n29632 = ~n29630 & n29631;
  assign n29633 = ~n29628 & n29632;
  assign n29634 = n29626 & ~n29633;
  assign n29635 = ~n29626 & n29633;
  assign n29636 = ~n29634 & ~n29635;
  assign n29637 = ~n29520 & n29529;
  assign n29638 = ~n29521 & ~n29637;
  assign n29639 = ~n29636 & ~n29638;
  assign n29640 = n29636 & n29638;
  assign n29641 = ~n29639 & ~n29640;
  assign n29642 = ~n29534 & ~n29546;
  assign n29643 = ~n29641 & n29642;
  assign n29644 = n29641 & ~n29642;
  assign n29645 = ~n29643 & ~n29644;
  assign n29646 = n3810 & n21003;
  assign n29647 = n3886 & n24596;
  assign n29648 = n3884 & n21288;
  assign n29649 = n4380 & n24428;
  assign n29650 = ~n29646 & ~n29648;
  assign n29651 = ~n29649 & n29650;
  assign n29652 = ~n29647 & n29651;
  assign n29653 = pi29  & n29652;
  assign n29654 = ~pi29  & ~n29652;
  assign n29655 = ~n29653 & ~n29654;
  assign n29656 = n29645 & n29655;
  assign n29657 = ~n29645 & ~n29655;
  assign n29658 = ~n29656 & ~n29657;
  assign n29659 = n86 & n24494;
  assign n29660 = n4420 & n25342;
  assign n29661 = n4600 & n24562;
  assign n29662 = n4615 & n25336;
  assign n29663 = ~n29659 & ~n29661;
  assign n29664 = ~n29662 & n29663;
  assign n29665 = ~n29660 & n29664;
  assign n29666 = pi26  & n29665;
  assign n29667 = ~pi26  & ~n29665;
  assign n29668 = ~n29666 & ~n29667;
  assign n29669 = ~n29658 & ~n29668;
  assign n29670 = n29658 & n29668;
  assign n29671 = ~n29669 & ~n29670;
  assign n29672 = ~n29551 & n29563;
  assign n29673 = ~n29552 & ~n29672;
  assign n29674 = ~n29671 & ~n29673;
  assign n29675 = n29671 & n29673;
  assign n29676 = ~n29674 & ~n29675;
  assign n29677 = n5044 & n25599;
  assign n29678 = n5045 & n26100;
  assign n29679 = n5109 & n25853;
  assign n29680 = n5130 & n26094;
  assign n29681 = ~n29677 & ~n29679;
  assign n29682 = ~n29680 & n29681;
  assign n29683 = ~n29678 & n29682;
  assign n29684 = pi23  & n29683;
  assign n29685 = ~pi23  & ~n29683;
  assign n29686 = ~n29684 & ~n29685;
  assign n29687 = n29676 & ~n29686;
  assign n29688 = ~n29676 & n29686;
  assign n29689 = ~n29687 & ~n29688;
  assign n29690 = n29611 & n29689;
  assign n29691 = ~n29611 & ~n29689;
  assign n29692 = ~n29690 & ~n29691;
  assign n29693 = ~n29574 & n29585;
  assign n29694 = ~n29573 & ~n29693;
  assign n29695 = ~n29692 & ~n29694;
  assign n29696 = n29692 & n29694;
  assign n29697 = ~n29695 & ~n29696;
  assign n29698 = ~n29488 & n29588;
  assign n29699 = ~n29594 & ~n29698;
  assign n29700 = ~n29697 & n29699;
  assign n29701 = n29697 & ~n29699;
  assign n29702 = ~n29700 & ~n29701;
  assign n29703 = n29596 & n29702;
  assign n29704 = ~n29596 & ~n29702;
  assign po24  = ~n29703 & ~n29704;
  assign n29706 = ~n29696 & ~n29701;
  assign n29707 = n86 & n24562;
  assign n29708 = n4420 & n25605;
  assign n29709 = n4600 & n25336;
  assign n29710 = n4615 & n25599;
  assign n29711 = ~n29707 & ~n29709;
  assign n29712 = ~n29710 & n29711;
  assign n29713 = ~n29708 & n29712;
  assign n29714 = pi26  & n29713;
  assign n29715 = ~pi26  & ~n29713;
  assign n29716 = ~n29714 & ~n29715;
  assign n29717 = ~n29640 & ~n29644;
  assign n29718 = ~n29625 & ~n29634;
  assign n29719 = ~n13050 & n26569;
  assign n29720 = pi20  & ~n29719;
  assign n29721 = ~pi20  & n29719;
  assign n29722 = ~n29720 & ~n29721;
  assign n29723 = ~n245 & ~n332;
  assign n29724 = ~n361 & ~n512;
  assign n29725 = n29723 & n29724;
  assign n29726 = n628 & n1186;
  assign n29727 = n1242 & n1268;
  assign n29728 = n2078 & n29727;
  assign n29729 = n29725 & n29726;
  assign n29730 = n429 & n994;
  assign n29731 = n1535 & n29730;
  assign n29732 = n29728 & n29729;
  assign n29733 = n3223 & n14117;
  assign n29734 = n29732 & n29733;
  assign n29735 = n14971 & n29731;
  assign n29736 = n29734 & n29735;
  assign n29737 = n1938 & n29736;
  assign n29738 = n4879 & n29737;
  assign n29739 = n29519 & n29738;
  assign n29740 = ~n29519 & ~n29738;
  assign n29741 = ~n29739 & ~n29740;
  assign n29742 = n29722 & n29741;
  assign n29743 = ~n29722 & ~n29741;
  assign n29744 = ~n29742 & ~n29743;
  assign n29745 = ~n29718 & n29744;
  assign n29746 = n29718 & ~n29744;
  assign n29747 = ~n29745 & ~n29746;
  assign n29748 = n748 & n21006;
  assign n29749 = n880 & n23833;
  assign n29750 = n3692 & n20906;
  assign n29751 = n3694 & n21003;
  assign n29752 = ~n29748 & ~n29750;
  assign n29753 = ~n29751 & n29752;
  assign n29754 = ~n29749 & n29753;
  assign n29755 = n29747 & ~n29754;
  assign n29756 = ~n29747 & n29754;
  assign n29757 = ~n29755 & ~n29756;
  assign n29758 = n29717 & ~n29757;
  assign n29759 = ~n29717 & n29757;
  assign n29760 = ~n29758 & ~n29759;
  assign n29761 = n3810 & n21288;
  assign n29762 = n3886 & n24584;
  assign n29763 = n3884 & n24428;
  assign n29764 = n4380 & n24494;
  assign n29765 = ~n29761 & ~n29763;
  assign n29766 = ~n29764 & n29765;
  assign n29767 = ~n29762 & n29766;
  assign n29768 = pi29  & n29767;
  assign n29769 = ~pi29  & ~n29767;
  assign n29770 = ~n29768 & ~n29769;
  assign n29771 = n29760 & ~n29770;
  assign n29772 = ~n29760 & n29770;
  assign n29773 = ~n29771 & ~n29772;
  assign n29774 = n29716 & n29773;
  assign n29775 = ~n29716 & ~n29773;
  assign n29776 = ~n29774 & ~n29775;
  assign n29777 = n29645 & ~n29655;
  assign n29778 = ~n29669 & ~n29777;
  assign n29779 = n29776 & n29778;
  assign n29780 = ~n29776 & ~n29778;
  assign n29781 = ~n29779 & ~n29780;
  assign n29782 = n5044 & n25853;
  assign n29783 = n5045 & n26347;
  assign n29784 = n5109 & n26094;
  assign n29785 = n5130 & n26341;
  assign n29786 = ~n29782 & ~n29784;
  assign n29787 = ~n29785 & n29786;
  assign n29788 = ~n29783 & n29787;
  assign n29789 = pi23  & n29788;
  assign n29790 = ~pi23  & ~n29788;
  assign n29791 = ~n29789 & ~n29790;
  assign n29792 = ~n29675 & n29686;
  assign n29793 = ~n29674 & ~n29792;
  assign n29794 = n29791 & n29793;
  assign n29795 = ~n29791 & ~n29793;
  assign n29796 = ~n29794 & ~n29795;
  assign n29797 = ~n29781 & n29796;
  assign n29798 = n29781 & ~n29796;
  assign n29799 = ~n29797 & ~n29798;
  assign n29800 = ~n29609 & ~n29689;
  assign n29801 = ~n29610 & ~n29800;
  assign n29802 = n29799 & n29801;
  assign n29803 = ~n29799 & ~n29801;
  assign n29804 = ~n29802 & ~n29803;
  assign n29805 = ~n29706 & n29804;
  assign n29806 = n29706 & ~n29804;
  assign n29807 = ~n29805 & ~n29806;
  assign n29808 = ~n29703 & ~n29807;
  assign n29809 = n29703 & n29807;
  assign po25  = ~n29808 & ~n29809;
  assign n29811 = ~n29791 & n29793;
  assign n29812 = ~n29798 & ~n29811;
  assign n29813 = ~n29716 & n29773;
  assign n29814 = ~n29780 & ~n29813;
  assign n29815 = ~n29740 & ~n29742;
  assign n29816 = ~n136 & ~n145;
  assign n29817 = ~n370 & n29816;
  assign n29818 = n2208 & n2451;
  assign n29819 = n2502 & n5299;
  assign n29820 = n5678 & n29819;
  assign n29821 = n29817 & n29818;
  assign n29822 = n1279 & n29821;
  assign n29823 = n2478 & n29820;
  assign n29824 = n29822 & n29823;
  assign n29825 = n4171 & n15042;
  assign n29826 = n29824 & n29825;
  assign n29827 = n2545 & n13643;
  assign n29828 = n29826 & n29827;
  assign n29829 = n4491 & n29828;
  assign n29830 = ~n29815 & n29829;
  assign n29831 = n29815 & ~n29829;
  assign n29832 = ~n29830 & ~n29831;
  assign n29833 = n748 & n20906;
  assign n29834 = n880 & n21294;
  assign n29835 = n3692 & n21003;
  assign n29836 = n3694 & n21288;
  assign n29837 = ~n29833 & ~n29835;
  assign n29838 = ~n29836 & n29837;
  assign n29839 = ~n29834 & n29838;
  assign n29840 = n29832 & ~n29839;
  assign n29841 = ~n29832 & n29839;
  assign n29842 = ~n29840 & ~n29841;
  assign n29843 = ~n29745 & n29754;
  assign n29844 = ~n29746 & ~n29843;
  assign n29845 = ~n29842 & ~n29844;
  assign n29846 = n29842 & n29844;
  assign n29847 = ~n29845 & ~n29846;
  assign n29848 = n3810 & n24428;
  assign n29849 = n3886 & n24568;
  assign n29850 = n3884 & n24494;
  assign n29851 = n4380 & n24562;
  assign n29852 = ~n29848 & ~n29850;
  assign n29853 = ~n29851 & n29852;
  assign n29854 = ~n29849 & n29853;
  assign n29855 = pi29  & n29854;
  assign n29856 = ~pi29  & ~n29854;
  assign n29857 = ~n29855 & ~n29856;
  assign n29858 = n29847 & ~n29857;
  assign n29859 = ~n29847 & n29857;
  assign n29860 = ~n29858 & ~n29859;
  assign n29861 = ~n29759 & n29770;
  assign n29862 = ~n29758 & ~n29861;
  assign n29863 = n29860 & n29862;
  assign n29864 = ~n29860 & ~n29862;
  assign n29865 = ~n29863 & ~n29864;
  assign n29866 = n86 & n25336;
  assign n29867 = n4420 & n25859;
  assign n29868 = n4600 & n25599;
  assign n29869 = n4615 & n25853;
  assign n29870 = ~n29866 & ~n29868;
  assign n29871 = ~n29869 & n29870;
  assign n29872 = ~n29867 & n29871;
  assign n29873 = pi26  & n29872;
  assign n29874 = ~pi26  & ~n29872;
  assign n29875 = ~n29873 & ~n29874;
  assign n29876 = n29865 & ~n29875;
  assign n29877 = ~n29865 & n29875;
  assign n29878 = ~n29876 & ~n29877;
  assign n29879 = n29814 & ~n29878;
  assign n29880 = ~n29814 & n29878;
  assign n29881 = ~n29879 & ~n29880;
  assign n29882 = n5044 & n26094;
  assign n29883 = n5045 & n26575;
  assign n29884 = n5109 & n26341;
  assign n29885 = n5130 & n26569;
  assign n29886 = ~n29882 & ~n29884;
  assign n29887 = ~n29885 & n29886;
  assign n29888 = ~n29883 & n29887;
  assign n29889 = pi23  & n29888;
  assign n29890 = ~pi23  & ~n29888;
  assign n29891 = ~n29889 & ~n29890;
  assign n29892 = n29881 & ~n29891;
  assign n29893 = ~n29881 & n29891;
  assign n29894 = ~n29892 & ~n29893;
  assign n29895 = n29812 & n29894;
  assign n29896 = ~n29812 & ~n29894;
  assign n29897 = ~n29895 & ~n29896;
  assign n29898 = ~n29802 & ~n29805;
  assign n29899 = n29897 & n29898;
  assign n29900 = ~n29897 & ~n29898;
  assign n29901 = ~n29899 & ~n29900;
  assign n29902 = n29809 & n29901;
  assign n29903 = ~n29809 & ~n29901;
  assign po26  = ~n29902 & ~n29903;
  assign n29905 = ~n256 & ~n259;
  assign n29906 = ~n365 & ~n443;
  assign n29907 = n29905 & n29906;
  assign n29908 = n431 & n533;
  assign n29909 = n702 & n799;
  assign n29910 = n2043 & n2208;
  assign n29911 = n29909 & n29910;
  assign n29912 = n29907 & n29908;
  assign n29913 = n12718 & n14903;
  assign n29914 = n29912 & n29913;
  assign n29915 = n29911 & n29914;
  assign n29916 = n24361 & n27847;
  assign n29917 = n29915 & n29916;
  assign n29918 = n22118 & n29917;
  assign n29919 = n684 & n29918;
  assign n29920 = n29829 & ~n29919;
  assign n29921 = ~n29829 & n29919;
  assign n29922 = ~n29920 & ~n29921;
  assign n29923 = ~n29830 & n29839;
  assign n29924 = ~n29831 & ~n29923;
  assign n29925 = n29922 & n29924;
  assign n29926 = ~n29922 & ~n29924;
  assign n29927 = ~n29925 & ~n29926;
  assign n29928 = n748 & n21003;
  assign n29929 = n880 & n24596;
  assign n29930 = n3692 & n21288;
  assign n29931 = n3694 & n24428;
  assign n29932 = ~n29928 & ~n29930;
  assign n29933 = ~n29931 & n29932;
  assign n29934 = ~n29929 & n29933;
  assign n29935 = n29927 & n29934;
  assign n29936 = ~n29927 & ~n29934;
  assign n29937 = ~n29935 & ~n29936;
  assign n29938 = ~n29846 & ~n29858;
  assign n29939 = n29937 & n29938;
  assign n29940 = ~n29937 & ~n29938;
  assign n29941 = ~n29939 & ~n29940;
  assign n29942 = n3810 & n24494;
  assign n29943 = n3886 & n25342;
  assign n29944 = n3884 & n24562;
  assign n29945 = n4380 & n25336;
  assign n29946 = ~n29942 & ~n29944;
  assign n29947 = ~n29945 & n29946;
  assign n29948 = ~n29943 & n29947;
  assign n29949 = pi29  & n29948;
  assign n29950 = ~pi29  & ~n29948;
  assign n29951 = ~n29949 & ~n29950;
  assign n29952 = n29941 & n29951;
  assign n29953 = ~n29941 & ~n29951;
  assign n29954 = ~n29952 & ~n29953;
  assign n29955 = n86 & n25599;
  assign n29956 = n4420 & n26100;
  assign n29957 = n4600 & n25853;
  assign n29958 = n4615 & n26094;
  assign n29959 = ~n29955 & ~n29957;
  assign n29960 = ~n29958 & n29959;
  assign n29961 = ~n29956 & n29960;
  assign n29962 = pi26  & n29961;
  assign n29963 = ~pi26  & ~n29961;
  assign n29964 = ~n29962 & ~n29963;
  assign n29965 = ~n29954 & n29964;
  assign n29966 = n29954 & ~n29964;
  assign n29967 = ~n29965 & ~n29966;
  assign n29968 = ~n20910 & n26569;
  assign n29969 = n5044 & n26341;
  assign n29970 = n5045 & ~n26793;
  assign n29971 = ~n29968 & ~n29969;
  assign n29972 = ~n29970 & n29971;
  assign n29973 = pi23  & n29972;
  assign n29974 = ~pi23  & ~n29972;
  assign n29975 = ~n29973 & ~n29974;
  assign n29976 = ~n29863 & n29875;
  assign n29977 = ~n29864 & ~n29976;
  assign n29978 = ~n29975 & n29977;
  assign n29979 = n29975 & ~n29977;
  assign n29980 = ~n29978 & ~n29979;
  assign n29981 = n29967 & ~n29980;
  assign n29982 = ~n29967 & n29980;
  assign n29983 = ~n29981 & ~n29982;
  assign n29984 = ~n29880 & n29891;
  assign n29985 = ~n29879 & ~n29984;
  assign n29986 = ~n29983 & ~n29985;
  assign n29987 = n29983 & n29985;
  assign n29988 = ~n29986 & ~n29987;
  assign n29989 = ~n29812 & n29894;
  assign n29990 = ~n29900 & ~n29989;
  assign n29991 = ~n29988 & n29990;
  assign n29992 = n29988 & ~n29990;
  assign n29993 = ~n29991 & ~n29992;
  assign n29994 = n29902 & n29993;
  assign n29995 = ~n29902 & ~n29993;
  assign po27  = ~n29994 & ~n29995;
  assign n29997 = ~n29987 & ~n29992;
  assign n29998 = n29941 & ~n29951;
  assign n29999 = ~n29954 & ~n29964;
  assign n30000 = ~n29998 & ~n29999;
  assign n30001 = n86 & n25853;
  assign n30002 = n4420 & n26347;
  assign n30003 = n4600 & n26094;
  assign n30004 = n4615 & n26341;
  assign n30005 = ~n30001 & ~n30003;
  assign n30006 = ~n30004 & n30005;
  assign n30007 = ~n30002 & n30006;
  assign n30008 = pi26  & n30007;
  assign n30009 = ~pi26  & ~n30007;
  assign n30010 = ~n30008 & ~n30009;
  assign n30011 = ~n30000 & n30010;
  assign n30012 = n30000 & ~n30010;
  assign n30013 = ~n30011 & ~n30012;
  assign n30014 = n29927 & ~n29934;
  assign n30015 = ~n29940 & ~n30014;
  assign n30016 = ~n29921 & ~n29925;
  assign n30017 = ~n21223 & n26569;
  assign n30018 = pi23  & ~n30017;
  assign n30019 = ~pi23  & n30017;
  assign n30020 = ~n30018 & ~n30019;
  assign n30021 = ~n278 & ~n460;
  assign n30022 = n593 & n30021;
  assign n30023 = n898 & n3664;
  assign n30024 = n5495 & n30023;
  assign n30025 = n2369 & n30022;
  assign n30026 = n14890 & n30025;
  assign n30027 = n5307 & n30024;
  assign n30028 = n30026 & n30027;
  assign n30029 = n3654 & n30028;
  assign n30030 = n3845 & n30029;
  assign n30031 = n12323 & n30030;
  assign n30032 = n29919 & n30031;
  assign n30033 = ~n29919 & ~n30031;
  assign n30034 = ~n30032 & ~n30033;
  assign n30035 = n30020 & n30034;
  assign n30036 = ~n30020 & ~n30034;
  assign n30037 = ~n30035 & ~n30036;
  assign n30038 = ~n30016 & n30037;
  assign n30039 = n30016 & ~n30037;
  assign n30040 = ~n30038 & ~n30039;
  assign n30041 = n748 & n21288;
  assign n30042 = n880 & n24584;
  assign n30043 = n3692 & n24428;
  assign n30044 = n3694 & n24494;
  assign n30045 = ~n30041 & ~n30043;
  assign n30046 = ~n30044 & n30045;
  assign n30047 = ~n30042 & n30046;
  assign n30048 = n30040 & ~n30047;
  assign n30049 = ~n30040 & n30047;
  assign n30050 = ~n30048 & ~n30049;
  assign n30051 = n30015 & ~n30050;
  assign n30052 = ~n30015 & n30050;
  assign n30053 = ~n30051 & ~n30052;
  assign n30054 = n3810 & n24562;
  assign n30055 = n3886 & n25605;
  assign n30056 = n3884 & n25336;
  assign n30057 = n4380 & n25599;
  assign n30058 = ~n30054 & ~n30056;
  assign n30059 = ~n30057 & n30058;
  assign n30060 = ~n30055 & n30059;
  assign n30061 = pi29  & n30060;
  assign n30062 = ~pi29  & ~n30060;
  assign n30063 = ~n30061 & ~n30062;
  assign n30064 = n30053 & ~n30063;
  assign n30065 = ~n30053 & n30063;
  assign n30066 = ~n30064 & ~n30065;
  assign n30067 = ~n30013 & n30066;
  assign n30068 = n30013 & ~n30066;
  assign n30069 = ~n30067 & ~n30068;
  assign n30070 = n29967 & ~n29978;
  assign n30071 = ~n29979 & ~n30070;
  assign n30072 = n30069 & n30071;
  assign n30073 = ~n30069 & ~n30071;
  assign n30074 = ~n30072 & ~n30073;
  assign n30075 = ~n29997 & n30074;
  assign n30076 = n29997 & ~n30074;
  assign n30077 = ~n30075 & ~n30076;
  assign n30078 = ~n29994 & ~n30077;
  assign n30079 = n29994 & n30077;
  assign po28  = ~n30078 & ~n30079;
  assign n30081 = ~n30072 & ~n30075;
  assign n30082 = ~n30000 & ~n30010;
  assign n30083 = ~n30067 & ~n30082;
  assign n30084 = ~n30033 & ~n30035;
  assign n30085 = ~n145 & ~n245;
  assign n30086 = n164 & n30085;
  assign n30087 = n292 & n528;
  assign n30088 = n782 & n1087;
  assign n30089 = n2108 & n2501;
  assign n30090 = n4325 & n30089;
  assign n30091 = n30087 & n30088;
  assign n30092 = n14081 & n30086;
  assign n30093 = n30091 & n30092;
  assign n30094 = n6925 & n30090;
  assign n30095 = n30093 & n30094;
  assign n30096 = n3643 & n30095;
  assign n30097 = n912 & n30096;
  assign n30098 = n14901 & n30097;
  assign n30099 = n24524 & n30098;
  assign n30100 = ~n30084 & n30099;
  assign n30101 = n30084 & ~n30099;
  assign n30102 = ~n30100 & ~n30101;
  assign n30103 = n748 & n24428;
  assign n30104 = n880 & n24568;
  assign n30105 = n3692 & n24494;
  assign n30106 = n3694 & n24562;
  assign n30107 = ~n30103 & ~n30105;
  assign n30108 = ~n30106 & n30107;
  assign n30109 = ~n30104 & n30108;
  assign n30110 = n30102 & ~n30109;
  assign n30111 = ~n30102 & n30109;
  assign n30112 = ~n30110 & ~n30111;
  assign n30113 = ~n30038 & n30047;
  assign n30114 = ~n30039 & ~n30113;
  assign n30115 = ~n30112 & ~n30114;
  assign n30116 = n30112 & n30114;
  assign n30117 = ~n30115 & ~n30116;
  assign n30118 = n3810 & n25336;
  assign n30119 = n3886 & n25859;
  assign n30120 = n3884 & n25599;
  assign n30121 = n4380 & n25853;
  assign n30122 = ~n30118 & ~n30120;
  assign n30123 = ~n30121 & n30122;
  assign n30124 = ~n30119 & n30123;
  assign n30125 = pi29  & n30124;
  assign n30126 = ~pi29  & ~n30124;
  assign n30127 = ~n30125 & ~n30126;
  assign n30128 = n30117 & ~n30127;
  assign n30129 = ~n30117 & n30127;
  assign n30130 = ~n30128 & ~n30129;
  assign n30131 = ~n30052 & n30063;
  assign n30132 = ~n30051 & ~n30131;
  assign n30133 = n30130 & n30132;
  assign n30134 = ~n30130 & ~n30132;
  assign n30135 = ~n30133 & ~n30134;
  assign n30136 = n86 & n26094;
  assign n30137 = n4420 & n26575;
  assign n30138 = n4600 & n26341;
  assign n30139 = n4615 & n26569;
  assign n30140 = ~n30136 & ~n30138;
  assign n30141 = ~n30139 & n30140;
  assign n30142 = ~n30137 & n30141;
  assign n30143 = pi26  & n30142;
  assign n30144 = ~pi26  & ~n30142;
  assign n30145 = ~n30143 & ~n30144;
  assign n30146 = n30135 & ~n30145;
  assign n30147 = ~n30135 & n30145;
  assign n30148 = ~n30146 & ~n30147;
  assign n30149 = ~n30083 & n30148;
  assign n30150 = n30083 & ~n30148;
  assign n30151 = ~n30149 & ~n30150;
  assign n30152 = n30081 & ~n30151;
  assign n30153 = ~n30081 & n30151;
  assign n30154 = ~n30152 & ~n30153;
  assign n30155 = n30079 & n30154;
  assign n30156 = ~n30079 & ~n30154;
  assign po29  = ~n30155 & ~n30156;
  assign n30158 = ~n30149 & ~n30153;
  assign n30159 = n3830 & n12765;
  assign n30160 = n2959 & n30159;
  assign n30161 = n3630 & n3638;
  assign n30162 = n3821 & n30161;
  assign n30163 = n30160 & n30162;
  assign n30164 = n24524 & n30163;
  assign n30165 = ~n30099 & n30164;
  assign n30166 = n30099 & ~n30164;
  assign n30167 = ~n30165 & ~n30166;
  assign n30168 = ~n30100 & n30109;
  assign n30169 = ~n30101 & ~n30168;
  assign n30170 = n30167 & n30169;
  assign n30171 = ~n30167 & ~n30169;
  assign n30172 = ~n30170 & ~n30171;
  assign n30173 = n748 & n24494;
  assign n30174 = n880 & n25342;
  assign n30175 = n3692 & n24562;
  assign n30176 = n3694 & n25336;
  assign n30177 = ~n30173 & ~n30175;
  assign n30178 = ~n30176 & n30177;
  assign n30179 = ~n30174 & n30178;
  assign n30180 = n30172 & n30179;
  assign n30181 = ~n30172 & ~n30179;
  assign n30182 = ~n30180 & ~n30181;
  assign n30183 = ~n30116 & ~n30128;
  assign n30184 = n30182 & n30183;
  assign n30185 = ~n30182 & ~n30183;
  assign n30186 = ~n30184 & ~n30185;
  assign n30187 = ~n24464 & n26569;
  assign n30188 = n86 & n26341;
  assign n30189 = n4420 & ~n26793;
  assign n30190 = ~n30187 & ~n30188;
  assign n30191 = ~n30189 & n30190;
  assign n30192 = ~pi26  & ~n30191;
  assign n30193 = pi26  & n30191;
  assign n30194 = ~n30192 & ~n30193;
  assign n30195 = n3810 & n25599;
  assign n30196 = n3886 & n26100;
  assign n30197 = n3884 & n25853;
  assign n30198 = n4380 & n26094;
  assign n30199 = ~n30195 & ~n30197;
  assign n30200 = ~n30198 & n30199;
  assign n30201 = ~n30196 & n30200;
  assign n30202 = pi29  & n30201;
  assign n30203 = ~pi29  & ~n30201;
  assign n30204 = ~n30202 & ~n30203;
  assign n30205 = ~n30194 & n30204;
  assign n30206 = n30194 & ~n30204;
  assign n30207 = ~n30205 & ~n30206;
  assign n30208 = ~n30186 & n30207;
  assign n30209 = n30186 & ~n30207;
  assign n30210 = ~n30208 & ~n30209;
  assign n30211 = ~n30133 & n30145;
  assign n30212 = ~n30134 & ~n30211;
  assign n30213 = n30210 & n30212;
  assign n30214 = ~n30210 & ~n30212;
  assign n30215 = ~n30213 & ~n30214;
  assign n30216 = ~n30158 & n30215;
  assign n30217 = n30158 & ~n30215;
  assign n30218 = ~n30216 & ~n30217;
  assign n30219 = ~n30155 & ~n30218;
  assign n30220 = n30155 & n30218;
  assign po30  = ~n30219 & ~n30220;
  assign n30222 = ~n24519 & n26569;
  assign n30223 = n30220 & ~n30222;
  assign n30224 = ~n30220 & n30222;
  assign n30225 = ~n30223 & ~n30224;
  assign n30226 = ~n30213 & ~n30216;
  assign n30227 = ~n30194 & ~n30204;
  assign n30228 = ~n30209 & ~n30227;
  assign n30229 = n30226 & ~n30228;
  assign n30230 = ~n30226 & n30228;
  assign n30231 = ~n30229 & ~n30230;
  assign n30232 = n30099 & n30231;
  assign n30233 = ~n30099 & ~n30231;
  assign n30234 = ~n30232 & ~n30233;
  assign n30235 = n3852 & n3881;
  assign n30236 = pi26  & ~n30235;
  assign n30237 = ~pi26  & n30235;
  assign n30238 = ~n30236 & ~n30237;
  assign n30239 = n30172 & ~n30179;
  assign n30240 = ~n30185 & ~n30239;
  assign n30241 = ~n30166 & ~n30170;
  assign n30242 = n30240 & ~n30241;
  assign n30243 = ~n30240 & n30241;
  assign n30244 = ~n30242 & ~n30243;
  assign n30245 = n3810 & n25853;
  assign n30246 = n3886 & n26347;
  assign n30247 = n3884 & n26094;
  assign n30248 = n4380 & n26341;
  assign n30249 = ~n30245 & ~n30247;
  assign n30250 = ~n30248 & n30249;
  assign n30251 = ~n30246 & n30250;
  assign n30252 = pi29  & ~n30251;
  assign n30253 = ~pi29  & n30251;
  assign n30254 = ~n30252 & ~n30253;
  assign n30255 = n748 & n24562;
  assign n30256 = n880 & n25605;
  assign n30257 = n3692 & n25336;
  assign n30258 = n3694 & n25599;
  assign n30259 = ~n30255 & ~n30257;
  assign n30260 = ~n30258 & n30259;
  assign n30261 = ~n30256 & n30260;
  assign n30262 = n30254 & ~n30261;
  assign n30263 = ~n30254 & n30261;
  assign n30264 = ~n30262 & ~n30263;
  assign n30265 = n30244 & n30264;
  assign n30266 = ~n30244 & ~n30264;
  assign n30267 = ~n30265 & ~n30266;
  assign n30268 = n30238 & ~n30267;
  assign n30269 = ~n30238 & n30267;
  assign n30270 = ~n30268 & ~n30269;
  assign n30271 = n30234 & ~n30270;
  assign n30272 = ~n30234 & n30270;
  assign n30273 = ~n30271 & ~n30272;
  assign n30274 = n30225 & n30273;
  assign n30275 = ~n30225 & ~n30273;
  assign po31  = n30274 | n30275;
endmodule
